// VWEAVE: BEGIN PERL
//
// matrix off;
//
// module;
// ports;
// wires;
// instance "RdmaStack.v","uRdmaStack";
// instance "ReceiveBuffer.v","uReceiveBuffer";
// instance "SendBufferV2.v" , "uSendBuffer";
// endmodule
// VWEAVE: END PERL
// VWEAVE: BEGIN GENERATED