`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zp8/YA12WOvJT0xWa6E4DOsKCCv5n6T0k+uU3m0kHAuwyNFpqKZeNmkaWAu27oVC
2Rne78O/CWZ7O43mdiYaezxZsJC39TG/3nOf5P749PSuqvOkaH80a/dgc/IgsMxI
89oj8gP2lPPJ/SNxQksnyo6LdBKlf0z9rjkE9iyewF8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36304)
7Va+cX3a2KMzqxQW7aG9jwdzi6qaDMyqUhvvnZeodIdn5PsZejGTZIZgJzkhbeNL
R7oN2EI+vzux7pTgTZa233GskAzxXg/on5KZ7IGdpSdGltk5EGeospcwgJe016in
xyGIJf4LM1K5SagTAAJL9BRFudP/NpW1EUsDrdcBkRlQ6+SCRMd2mvRsIxlsO7+4
JCtz1iegvykh2I2f24JWPKka3sFXyXkt7jUkPDPCC9kunFXbVRaKFDB4IqBd0N6j
cUlluVJq8anP/xWOQqS2+u4Yuge4FY6Q+tw115q8fZcmJO/HXoWS3zbCwf3WdBHE
Xsfe2hKOzldbOb1cBrD/4Vzjc5mNmuMWWiQToNf4sQFceA0SXosA/gom+hZ1F0F6
gpPllCOC0CBxdM9Qy2Huu2uqrrZMkI5rkodl8W+iZoZmif7ZqjmcpEr2dlPM/Q54
ADYwxUcEnUamJstgOrPn2MIsy32ApzWxaNmC6BGYqtfNDYAsjRxjFQhn4bqBiav8
+MsMqGCqxpRkO6opYYWLrk8+1MjS5QALxNUgalkE9cojYM1XQVluZFQFL2KiN20K
A+HMCY/Re2rq+dyK+mldnW73sjuTVjzonpMjC5p0MK15ZPZ930WbYDFB8KlmcBqh
Py2j56y2VbA1zLWimGAlYXbAXa5z6oyXetv5BtJeGCN8lO0UruFu8idERvj8NMii
n7lE071klxoFZw/K9EKWHB/5cvsrgGvRDgASqeh+kc/lRCDOnDwYRWg4cqxhRu2L
WPCOXtF3YPMl7lb4taEtGRxczaXPgXvgllgicFkPoU1TtsMuneuQ+MzmJntBvNiM
t3HdPM2eCNC6iwR/fiJZkAkLIfQ3owCb7UcvipnOlXc4tFWXGguTGbGx0YBS+IES
j7/TcfvtmxuR5KGjFNlJZK34gBELwpb+VoYwmuWedFcGDMAXTHgOttspDsLo/JW+
0R1BO44rfnuEUurpEFAf/dzfd5DBADvX7WNRSsTXSN5XWsRNze3mesgZDaUC9ySI
YNKC95F6wIBz0rJpbgTuA+t3exAGCPGTPsF4ZjsC2gQ33eRWePwm7BEKaSW37/UI
VRL30SgBeoJCcQI0IEG1aQTxpyamv6F5GGrvyiANFfah4MbgEx1lTcXMBAj89uiR
zR+MJqkggC604A6GW7os4rW0c5vDLGt9RvdmUm8XRlMSOLOnYfda+1K/UjaRPjpy
NmktHR2WewOldhyk7+X+5xAOmljkY5m4ssXq/i37FVcaglwQxUO0PKw19Jup/rNv
Xs4fs4MoS7te0j780kQVgr+8m3G6aRBy3YwC5drhv9tYk+0BJuk1uTlbSMDIECiH
GfZQ0qrFaCqFNxUyJg+X2chqekskaw8nSzaRF9CkcHC27yhAeGOiDpD2X5V7VmTa
ZZINaBUfI8+FKMjwLf6CN4XvLdRyjJAx+pTy41H8iQ83deUNb6AmfCjNDYM3J2aW
OJFlSpyyezmJeWfBr9mmIiTc2RMYb3AK1grJREJ073yXgBc0yCsGUO+ME9qXtU4T
tnrc7O/On9vh+msNOpsxXQDVWFT4uzoR1EI+90K6JF19bXXZWyeveYJBLDZ2E60U
zDbxf89eLB4fq4mt4k/GCKX0f5XfF1NOFbI15+N8vjTi7/QVyZBiCtCSpQhq7c+b
XRllHmzzmD8Iv6BUkQs0xmQAeGCy4l+HJtmdVAUWi0iZlFE2fs2HNAwqJaLf71/p
IevXnNf1/JlfuOo2JJPLNwjILP7SkLooZ7DXOZHLd4Xp1bwl7osD6AltRjFxPkyQ
BdeP1X3Hd7pNaoHhCqAaeWgCQfSRCvyGTaXZc2GqADJ6srIpiLA9TKhHTPLG4F9K
oMCPRZgAWtkohR0aSW0jzRn0JsLX+jiF38av5RUnE9lSeuSJjsYQ1HoC2d2mhNpF
2eApXmB7ckCdtL5C/gyTBbpgslzjuI7ralKHloNjW3+3V0MsqnOmS5wMphMf0YfF
4x9UIBC4BdKRphoyAbLhiZYNnMb8mfW5k05G7as3LyZ6freBN1vuaK7qWuYMgJcZ
XwxZTetTu8++GwiENqZM0EDJ3yELwl6wNRu1RPDZIS+rYqRPpyjw8uI7ji48zzqF
c183glqZ+2FFgJ8BpVTBm/91bp/zj5+Ot8gePPsjzAAmyNUQ5ZHvddjV98G10vZa
8Ml3nWkOXt4E8N/wdMGL7h+rcfUbizqYXLRaMjVCulSKrNDqfx34yQ+S0deolx4t
fF6L3gz89NK3J6SA/6iEKzZgay6JZ4SdnaBkcVyTCAALI99l+AdBwHj/U9DWtGd5
EtYDtheYOIKkkAVc7HEJ1AqRe+nrpvtUFTaSJifSbTHVHCpz7CDkw11lEzyqzDHZ
7PQmSBVv8WTLR+cibKBwFVexPeB7tTDLLJ9LHl7gw3sZp6ViUGu+Yo+s/N+sY6zC
shiwi3noUwTy7g0WVIV3XIYH9x0OfTmlbkPRzYusCNaMV6KugDSK+6BWdVF6N80y
5appfRRU8wlRrtgIBdHVdcjg+JQzYctv+063XtXX/mpn2rtTjugFUcgqSiTok/B3
OnXBjdXElKDJoSVUCKf0RbOQC730z05jNksslQqLZY+qeUK6yzgqMudboBRftlpB
cH8cK1O3S5Kd3bmiWfSpR9PJZm5qkg0TvwTW+/tlSBty7PFIyQnJx9VQuNdm2CGK
vlILRjmq3CIROssUvSNrOTx5Ud3LWfzV4vLgcAVBwfY0sb+sXg+0YCKLoxsaMzND
tFn96XOgzxDyPHB/T/Ke20Dxo7hpomOm1VkCJt2GeF9uE2cyZRK7GrK4zv2B0dHI
Jpv2yjtx6Te8+IDEz+E5U1/ZXxkmxc/Ck6oYqUZx4BPDoOwWvv2w/D77/K7tjiEm
Z40zp655jFqQmybEpRhvuJCTtXn1flO6ZlrD1+9Nu27LXE+95GJDM00mXQ98ECPj
YF0nP7k1pKaDP/zyLs4U9zJWuwMVN5zwXyWLc/E2Q9bu4PpGTj5HWZRv6rVf4PAh
O1Eh2A3ST4KUZi2l5W750OqS+sjtPYCKXmcqWbkNHY5ZK3FWFFr4dvL2MSHjgKGn
iYvbxa4PPcVnsxSnn5H4+p773/Y1ewTEJKTNcHMLW6jXEvZ4U9EUjtQDgh1mO/pz
qpfL0c/0YbrxWdeNQrvsgKQmvtrrKjvMKv4Jfa19pTIOYtd9YupSi+VoCNhhpPZd
AtqEG2Q1vqbjOY1+JqtHgB4+ZtWAUlBAe+mJVd5A/4c4zBn1pluSucpbmRj0lh2s
vc0ZBiTfs+QRnrvaSjWOnDFJLquUjSsieUSHe6r6S4TQdo4E7QJ15JCPukBfclxf
5XaYKQcSiQYVOmOaTtjH3lBw//ay9T84yF44xqXE8MPTvwWcNgoQ9v4xwUpy10cs
MevAK1qadh0dFzaWy0fyQ1EnWB9KDLZt/H9+ni/nCkV+30ylD7QzB7yqqR2R8fWp
eZbPHsM7rTrtq/fD8t5PR0wo5hOwHcD2+hzcf+pJYvRRttD6fx6VC3LH1g8S6z6E
py1tfFHrewLSJYdwl1lvyX1Nc5HCm9S8DBo9FAcpZLhknxG2PRs+AW0iXDfu2fmD
POm4zMPnrlocqGIzGooC1TEUPV5XC8XNaMrtleEnP4Jy7u4u6ipVeL3ONrv4+cGD
tPRJTdmVu5jMjGkz7eAr21DSlyZLVfx1aT9LScejQhUK/3V0eMT9kviF5OooWZsS
+dW4T+gu0Mcs4y/2C/qSaqI0ZSKUrU7FeyCr5HY3EouzvkQXiC8/xOSDBbMQaHAq
ppx+ierOC7+04+n/xSXRWNMWN60Jcl4aE1Y14+F5IbpAVkUCjJ2JaBtvyhI87MFQ
0r/kQZGzTt6geNVInuHQ6buz1pmqncJaCn1xjZn20+RP2Cbjz3/iMVZD0+jzhubT
tP7G7B6DZibAad70mz60KgJz4QJh1ZF8FBn/bTT6+K91eiXp8AuhOjk+Bl+D5Ntc
CKbvknSPGDdz6p0OuddGUC+nzSXpvOKQfgnB3Zu7D1LTOdIi4oS9wQfAMxIQLPC3
XQ3a1hAygLsLr9FcVUc9mUS41JWu9Oo5EOuOFyEVwX6ohGDiPaFAbZRqohjCfWjA
a6bhn9nxqO10xxz0vK3jfvhQAPmJWeYu99kFQG2sLyk/ELuiDS1LFVRoi3qv57uJ
mhHJCsAy9XkxCx0qUaUycuYSknvC6qgkQo49iGzQygMfuOqkE+GfR7o08EfdRGlX
XkpYBhtrAi4NHP/JL/mcdczdh9kDkxadwUv+WTYhl1lwG/oYKGL8mTAdFx/oZpgC
pzj1hawx7MZycSYzvRTPN2AGY2Li0pvtFDzJpWPLPeX3+pHMK86iqJLGKBabVMvp
1tE5ol+zexZuv45EUMNrJ4J4hhyX9QaUOf7yqRB/VCP3XdLURW+/ucjucZSllQnw
byBxTf1aiblMCJVj+oYAo+fAenkQGwtqhQRjCyjjT3axGfUBesTBiFilOaDzSAoi
Q66a2lZH7FMEvdstb4uhYlPic+qCzVJVGpC+AKS3BlTHgyJK2sKhkfPj3Wh5jYjZ
QH24ZsnoXc31q+JxE7MUvpoZ6Kx5+5y+wf1cYyozxjlglWh6U4/tegEFWzoyQUch
tiumQPudyjFIfC67kQyJUOfS6ltONIJL7iluprlJW7j/x7DgnGT8Cp9cmayPLp8l
BQQZwOWMoFQlWEHrphv53p+ybm4reYGuZh+8oEP5jYw/XI4B4ldtpB/xstc7me4x
LHpxZj2/pyccgzjj6DQCKvHzelT1za2z5mnimb2PkpWS1GBhGgCdAhTcQJ5dGo1o
ABcvppQtvF1qnnOp1uPCjHHMsrW1tZodUntm6bfz9zxobsxuQ/JWc4BwEDUEANUa
N3kyVsvu4DAZmNUlFcI917A+SSo0mEKXpbcHISTX4wYrZb30aur2rBSQPnbLSKCB
Cx4mExymWqcGfsGru0Kb8VaDExoCR/ZC/wQjgVcSw/S33rQsJew7tqL3ICDX3vdu
VgDdEaL6rbiUdjEgYNgRXSWa0vDiPVeFfiZMiRcSfaYmnFOQHOgWJ84xybQf1kVk
U3/GPZQZgN1vXsaHezIQlLBu6uUXu2dYdPuQijoS31RY64WKwA7xKA9AHAvH83hD
xHaTBW+x5muzv1Lel+m8fkSoLEiX2zVFa99jt8I8XoRsMyml3s9A+bMSCpUe/6G8
vLPhUaUKU8EPzgRRCA+WICAFEKLVzPK3BcZKzEMncrsao65Z+ggWqYyZAnCveH3R
SuaGvwRet+W66G7IDHTp697yF6abQGSX0QAznbYaxMX9q9ftNyFaSDW9vkJvdClD
t9d5XRN/LQx1sYPCu1yVinPk46VsdrnvGMjkDfV3n/+fGkwiVhZafJWJXq7eKOYe
fgUIlvDXNg9BMC+xpM7a8BUJinNUxtGe5VHDe68+Cry7X2feUWeq9MlQAXN2xlIK
JqjMtL3OOt8c/BB7R6SKhWQZapX7bw3RBPs7Udqh6V03LO5VKbIELoVFjs/P6NIP
HbPaPb7o4/JT0N7hz3fpd01IKfFturM5Uf3m35/gXzsk+89EB35HKd7Ef//q7g3D
KKuUxnY/7QlXHjbX6D/mNXfOJlGZkq0e1wTES2BY6tcXIQl6hLsLbsM9AnWv09IQ
+I9DsAuUMHb5QDR+0ePx/ZVh7mpbscmsYlkkIkxGd0nFKB4Laom3mDE2Mi7/81KG
ccw4LOE7nHx/0dkqGIVkE45yHI0XmsO5dtKwPxIMq7bA7OB5UqJIT1Hxhed8W/w1
9B0jKl7Ba42trvAmf0oJVcLXFMEv1nuB8u8felFPBUsaDdLME0daX2qKv7ZraV8/
bLO28+xnVgGIk4jEMEU+I/L9RlCuFCFPPFBmTbcpY81ZPoH/Q3Tn0ipjSUaNht42
+alo1KXxUjvP5O9I9sgPasW5c1VQVOsdaFBdxEImQi3Ha9lEadpMk6HqiPjy2Ey7
/hlTtCNIjWPU+t23CqFI+CVsPMI3C55UturdM06Qjy7j9UvDY4YUH0cedxC3ZMvs
pZigJPgciOlpvhJsYNal/k8LnGMZF5JW5wKYa5DVvhXgc/td69Mlq6/0xRZ9L4J7
b0K4Ctwt/oSatV1JEAAZaxM+DDP2TfmAFrgNtyOHbGXhJjAdfvKD1pr+pLVumygb
F3oVWo1pF9ofuTF0NVhktmGgzJ8JTvdzzTpV9OOvJbhTiVv9cYBnDVrdIjNAkxgx
RGUNsUsD7YVDtkjxy3MMJHnO4izZlJW50P6Vg5wlyC4IwH6gI3ar3CStQEDukw08
ocSUVcCPgMss6kxTWIBFhdpDuA1AuI/H+6nQx7BSDiHWc34LTEG+d4zfR3lL6GB5
b9IVGBid+7Cgdnm5htCl11ICPaWMkCFNdt5a3SQJYX2dw8C6CQK25VzDly3JNpeX
lyY3H+TpvN2a92Z9jVq+vYYykigYHaBYakRv8NXxsAs+rHyZ1FIb9dx5yKi29viE
0+T72dTn7Y1uT7XHXPAwuadQvfEfrsZnwY124NjYlguwWJJ7AmlbBgcTDfQiYJBd
R4Xt4v+sJW1tiapRu8h51qYyOX2aosjgp1gBG1gGn2yEKp9IDp/f2i0GWY98JA3G
/oAVk60LuRWWdtBZheBboPWDIoIquoZtXIu/Id9cn4+mNjaw2kzTdNN06BKp2y4C
IIk3NNXr2JhTAMPXELA8IrVxaZk+JEMFQMFvGDfpScLRebkFSVlpO750n+BFicW1
ijRagPwD5J9Gra7ZDn1uJSWMErR+w/hVbV55+fRdeYDuF/943WdPBUB3iFLa+2HK
945QePxHCj7Mnc7PAmGeH4/DSazU3dhCvhrw53bsK8LGhqNXMcGJq7HXFhyIlLAG
sIfGYJCQsAtVoUuqupTjEEPsnHW3ST2Q3h34GkXJeEP86y4FxpPhPZgUudtLWfbd
+EwS3J8KTbRx+Piq66QVpliNo6Elcq3CKcpw9OgntkhKEutiVXDVR8gDBsl83I7/
rjvddPS7S+8DVzWVoN8jRN30257yVZkZajNsRDLkDKfaSgc2KiK+mTECcwgox3HY
D5hqK4kSWtIZSWr1gT3yYU6NaKMB/8j4TZ5463MfCQ+bTjPpZJJu/XixB2GP4SLT
Q7yzhmdqLYe4bgBuMRKd7Ql/gEEjJqSFQdctZCDRHf7Ov2DDTprH0mzy5F4Z/iIi
l7RHCyE5PQLb3R6NsWPIN6YyhbqO7AZoPkJBRrDtMoMvD7GbFHae1JnS6yq9rPHP
pOixdQHIigeKcRrDz5/PVs0MTUmlLfMINRf1pyJJN+ThYhbADxmijc2521S1sYPp
D0HUrYqeljH0JLjt0bJyxQoaVOgJPTOeykBJbxc+5vEnwIUqdH999FmjDRishYUb
R+Yy7/mLewXWiHDcXLq2k3c5kshjbLpnwUImAuVLwMiRmjxxXFONwatZKGFRvjV9
YH9U2mGygbsJxdBW9QsZoHMA2ZXo0tDPWYJKnuVzHoTkTM95bv2xryed0dXjNXdU
ncTK6Md6j2RREtLFsWdq9G7M7JjhyQm6MqO5szJvjrh3Yzrp/T/qLKTYH0ybJdSF
oRP9J/30di0Ng+FsISHXEMFqlsXlSShUJ/PyE02mkOoV4FA/zP7BYR0EHkAajf0O
0tgj5hA8dtgTpmpPAJBg+QuF8NFtg2ETU40lm19wTRrp7ba7YMuyG7kMNowUwNpt
KSoiQtZ6K8xk61oDGtDXE8zIWpIvVNhQdmYuFyesOmARglCmn57zwt8Uf0O2oI0I
y++D055aoHs2d8b0N2IktJ+eu84o4XoqVvICcFJhsO/h461/mUi6VAf3MZ+klza4
lf25jovsw6Od2wSYfuuk8PZ2r5NXn0YIrQ3wHx50LCi5LoxjpuzwyKdC/+nFQkIU
7jIwNc65FhVOt1383a82uP89d7qBPnHfNXehoe7JIypouqDVvQtI46hsXh6SAatX
Pj24WH2KGy96N677mtaU5182g0d2Q/FBJDEK+lWtTStib0//DMMnrlw3g7u6F8bX
hdl/iDs1txmiQjMo5gZruJJfMBKTJJ6/Jj3pa5emjmKvJ9nuN7w+4vF1RT14T9WI
eb6RBszDcQAs3B7ixfMp3HkLEJ7SFBZlbdIebht6HVw1L+PQuMjw+b8102YBJukc
2dYwKFiSe+SvsSaHgDfamaET+cfrHgWLTzAcY8unPdLJbwL9WXYZ8imSBeLykIFy
lIQMPnuX9GDfEpcU4SaI91vECjpmdZ8SSAqLRnrcWM6/X5oCOXbha+rHfnAvvkdB
n3CB382wyLCx/bKU1O72JEwAYidaZoq2rorZITcuGDR+pKwppTOkit/YK12NtGLZ
tJ/0Zyp7UoqdrKRrWRguTLmRBdV7Kmk/alNGDAsWELcMOHy3bipyd/7Sa1EMQvST
HsP9mZ5aTUJeKb4dScDMICzdjhXDeg2UktgX8GodRuq66F1LbiDVUMxxkxqXd34o
3oI4I7V6i2EQ7nFZhfNb/R3DPT0Bz/1mmq1craDZ9sz1ZfxPI7PkPpKDKeF13bde
E40PGbNGys5Vf6spLpaehQH2A39FUoX7s65LcmZD3TmStLN79GWL6qH28+0UwrbT
ZMHAsyvHTiOL60kX7yQVgSLBFsz7Ra2U+NwSKw9hqqfXq1VLisEyBKr4xEE3ms7T
cdcQSJIARP7xZ6z5vLhf6USvT4OqYji9wvY7waeVxkHtaBkCFWfbR+2n6CeIBXnd
5MAfu2+b95JZe/EgMsngHUElFzff5e/+vDi2I+6cenSPMh6aBL1uSb3a/3sz/KV7
V24iUObWUKDKNztA+R4DFCHufGJvFzCe/scHtySCkzIz6Q1NjEBNCsR4T8O2Lcsp
njWhsyUflVyW32Dpu1UZ1tcDVKz7EHbwsPRzBliDBaToVG83LMk8Ko+Tx8PzSaqz
ivDajsSbL7tYDjkCG1a+yJiT/9FvoW0sXPhmax69Ro5097TpYBUm3uoNlQeiDGNt
PjdFkwgJQb1P1YN0hMECoPR/bMPYgFu81LfYSX0yd5JrXuAUQhmm6wg7Tm8hDiUh
+rh8DSSZXiX7FvC97wm3Y3ZXHm+3rwDZm74I4aUnkw/A0HaMxcD819NG5L/maNGW
eZvYJuvIbMN5cecK2rsVf/ymaJFSQU71HEClXwA8qakjopthg0eH+x5UsJiUYma9
KyIoNP1hZab/CQl2EMOCOYasBrOGAatgjRFoDZ2SFkXtfXArSAkiPuiVp9TGhrNf
wpyQPjcUcB442YnNdDeZbpRBO2FL7VxspnzZ5iiRi5jc3kGZyJZi5wX+d1IQCOQ1
lsFFhYDkoozO0Ijhg070ihLomuFGnnhjrEwrdcvZtNowPhFprSTP3HtAQTI2U1q0
9zFaDh7DjWGBjQ1n6BChAgGahM68JM7LAhW312ietBtw7kxadb9+x1zHcShWbmnZ
ZWi66Ym5HsryWnb0JFkt0XXzSI4hGCJR2Qj0WmztEPhcBpbC1SMLqV2rvf9fW385
St9oz+qyPB6H3Neo2zomHzbQCmrmQ8o8VoVXNYNmpd2NkEs2ydjSzGysM/rqOFGr
UlCCgqDZIH94IjYSHUdnv4r4ZBFB5b9Iuwf7tuHP0TSoROI56t543Fubx3pRg1oc
+k96NdwvLaarTi2n89YpFMsPkrAbDbMR6bfcSti7HYEbsBIbi1V4RGXQmd4yQb2w
pEkrTN7KgSkOQfstpr7Z/9Z/EtWauMRAB9rtQgD4U+P3+HobwsKizpG5+mwyVZc1
1N3uEqgffT/p+XjB4KdLmQhUf498h81O3BTg8a36cctOK+feiP0OCJ1X3RW2SbJE
IKkydomLPPYoq85UsziPnhFKQoU3dvVXFLmI2iTzDzXvFS9iqS7UPjmUVh/Sb4s8
930QySnvGoYq/qZzFqvq1kcAAQ5mw2msk6007m3SuMz5zwu4g0NVm9K9+Ks//kL8
ff+luRL1+umqOJLC+CdXGAzrnjI1h6XipEkcXJdaWkA9jbtLUt12qxyAFzMe05QA
NBYlnVYzDW2v9d0QAmLsyqKoY5bPELKurW7i815QmqTuU6EXB9X4/kTWEnwfYGw2
X/+RcRSE49SJz5Ot+QA8uQ1e7E7jSDM6mnxUKe1vz5LnwRYuPcbgNAKV4UIrAzC6
xTjoEAbPLQKrW/EsYAcvjTwNq0Gs/RAyICJqEpDIs4SwOG+zDZKxgrCW2+AvBV/F
ex6W7uLz4hjZDYSpePNFH+A1YlfCG44y5fZ1kgz/MWezyWVDrhCw2aL/qBWKoUWY
uXFdG/5x+jJ/akiW7Q0nFVokihybJ+A6PzUDMqXVTPCAnrPdFYTBSybVRHG98Qfa
nwJohYOG/4z508mrQMJCtiGYMyZ/n93nWJAxWUCECce0ef3O9J1to7vHEt8ar7Me
UPO2Dnl49DVUvKRt1E+yPWTsJ1RpND52QI0QM1v9SwLfFv8PG+HeTLwBbTejJeEb
F/4JeBNzIdEEwkh7LdItruOEJZYNOeYAqX0n0GlE9eI2Ea9Q/SWw6aAzmmeK8GGD
3/3KijlhJYBPdaRCNsDYBOeFmpwd2cMeI0apcUCHt21rPWjpdsSDfCpaKNBdf6J4
9sCk9TiI0vi9fRq4hxg4EBAbOl0dtC0E2SHMr9nO0uAoVg+YoVy5M80/g93Szi+l
FKfafZEFXIb5cCyKbO8AJND7PMWhjc3wRK/Gd8M45DHNHODOaeqdbYQTiraURGii
zgIGTleTTZ9mXJbZlkcy36jbPeZXgaMjJTBQGiWSr4t8ont+Wfc1KEyHo+McI5lL
twRC1FaOAej1LsA/6hx5hC8Le8zc1lyGFUJJvtyBIm2+WpewkkK88ILrpt6CgoN4
jwvKpCerhWQ9jnD41pOEOeuOBJuoRfvKNExYoGM2N/a+rLTp+fmyWpf6B88Qxtl1
JHbAggmvWI49SRe6YhVOjFOLFx3tzljJXdY804PuFWHQV5dJesk1FNOseviae2av
+yyHHK+kHrhVFYbLe5IknOqlOX5/+CTMILuujM6FGLHvNXb2uWO/Oyx3qacXWt+I
eEtefnOxITcuzIpBL89ZSlhGYZRoEhxwz8UiwIcA/kqd1JIJXXBRPwTRGZwxId7v
kq9bXsWfLHx/CqhtM7hu9q+IyVpJocbLYUsDnXQAjGMwoe8XCLnzrD9RHWmBCyoP
t/D9fM+9uhq6nX/J5vh3F0agSCo3aw02vING58h0DxvCgpXRZ/nOV24EYeGJjDaF
nV6YDb2tuXzm7CA8sqll1Q1v1IMtO3bwWSlOe0QRn6syYYpbV2AFSyuYQAAJXa24
DmWfehO07gbTGWhcSl/Mfyz4zo3VCdPZOrp1gcm7Xm/505kpRqzGs/0wNCI3FfHz
eBXFZ19s3px4S3MRLpbg1TfrbiBa4lm1V1LEUIXGJENCh39qrJ46A14P1mdyXmM/
/rnbrYPQMufEwzd1lG43KigurCJ2VvYTAOq2nxMh/OKo2XL5qP3WJMUO1o2MhYpD
cpc41BzbfyRU/1TGeU9VXJfHXbPGAOhwL5DGblkcxaHpCPyLgT7eeoOzk5kglvfk
PL0UT7XD+936SG3FICPxoM90ynNWA0UWvwZysqkAvc4YJ7q3PCJIV2+dIiEAVjNY
5Q7t1AhLmJHTB2oXSAIKmG+kBBTy3j1L2KzMyJQyj1vjV9I9hik+5jfrhd1KFjlF
D/bnijgjarx2zX43Vr/4oGAFfkmhjKpOZNvrEaBZwDGg6SskdJRakm0j375eMKhi
o+Exqhq9wCp2Rf7Bz5cL57x1khDBdPrw6oRUTquTfhN7yfm8mpuxRDd+DAsPK0fl
PZ7bxNXZqRs7vXWX2BSSTopRkoM+cXdThACUQ3Wf8t+PH/XStgDZLTTcV2MjPKKz
Hbde1Y7GCNQKMKQrlfnkMA5qJk/pdBnsmyy9HIgjGKQm6cIwL00EtvoTAkMDKhLI
4g8XlcUyN6CtTlBbVKFrL9jEPI3r8GJ2fZd2ogXH6Ap/N+hy2Ohwqz6yJyDVWtnT
qE9fM6Pvl0ssRIbmlEKywjNzZHVgwJMqbOEDNgekEraB0P2pn3hJR1SPR+2JT6IB
oi9H+kI8K+7CuzuQ9VzQcuRT9wLMNRJsU6iNBqOUkHkYEoGWBi6Rc2BNoYmNpmZ/
uLHXsbq+Un5thhT9HhP8IXlG72DSRd6b3Vg9Va2WlNXQOHhBfiOvyQhfDa2/WXFq
mOV2uXwWP9HQE1IwA7ImrIiToflIwnse2VP9vkUvDPFX5v+jXplL6DoPxLr0P3uB
stmLZc1L87uCakdGgYLIWZYlpSInVwmaTP+I2Z5TnaP8fFTEiHoskgvmg6oWdV3H
19WLKmiC3DWqM3OFvWhLultfD8XdeGaq4l/V4JcGYm/JEoYHmTP0v1gckdwZKm+8
btDFLBEjrlvCTmf+P6Zvgw+fboNE7JQ1DkqdC7m+1blwd2zjoH6/qwOjSc1hXMnJ
zN7FODf91V4xzwUa+qHHqyJWyHxBfJ6UzSM3bmJdmI2VmNQI1FDI9dFTqJkw44t3
mLMugqIdEPxFzNz8n93BPjuX5y1MZfqEomZe3yzEDenY0oOmc49zMnS9DT+7+iuP
gzgzFsXrywSRWP/r0wRqKxj4hXEAnbw4No7u7srcRmEiBgz7STMN0Vp0nlBA3+Cf
hjjCOJ31kwI5Er+UoeM63dJ6mu7NRmW04+Kp8Kb1WNDksnnReMDdHLgN1xdMMdHO
TJ/FiiykEo0URUXh+Xftoh8OlISxTNXKdBRsdrBHEdqzjkplWfN3ZZY8LcpkH2Rq
7gm2GJWIcMuXLmq/TzGvrxB22aDnE13ZyF3gz8OFeyDrkwTOvG4QLRHCfr5ArCha
p1owWdG3sJS0gBk/fxrke3Gzstz504QpGK2KJGHegWsFGCSCM0gmIsIM3u8zBLBV
IlntgQc50m7/4k4VPUO6AZsn4nywaA3QD9MQ5CvD5MjyS5SUPkjeekOILdxN7EWu
xtEt/L9jF10T0ITsoZAqIxOQWb8SHGCp9cWrL00p79JUq/S9b+hCs0nt0drI54Sa
f0Mta16llC8QmPU3z88/uuYwDijyJ6UY28TfNyqNEmjm11sTJPAlPf4SVp735m1G
sf6F04x5O8rPyG1cXTq0QbGHpdQpdoDIuVW6qDsx2Alj8n2BD7j5gYuLBN4I2h9l
HxNPVxsaMEO9KMH050aTsex5X3eSfLIELGBje1e/IiU0KafPHifiTdYvgRcFJHPB
RSnmLTH+B7Wv13GrtgfyPFFWu+hFn8qgzZ6tXQwK6ZQI1iYzpEAFcw0AGmC0njzs
HwG2xq/Ngt14wZ2GHbBxTMRkg7mG0zbR+WCsTH4bH5/PncjmYjgzr/2O2JP9iqfw
InQgesx62GDWOKs5qH4YdQ7eu7SpMbLiaJn9OJC9e4WLcUcg+2v5357y7PxuQ0E6
Cf2jeLZY27A6RrjuIrHJ57u/gEBRkCD7uLwHuHzVzpQsHJCon1UhHWB/2bMxnI6U
uDv2wEIWKlKsTnqPrKj+y+aVH5g8HdCORkydQGFGRWx4HGkd4u9CbS4l9FgeQY8L
rDPYGjxgWAyNfmQ/WeciZY0wfcF3TI6++dp94++yGC4MrpVT1HT4fsuLNmUcA7EY
R12FEDbcLehVDstpPlPSZabJqCykDCAhaasGBk8iX8M4n2nRVtxmfLRvD2MAv5xl
MjqmKsdYZbA89UEazuzxrX8Qkngno86i8PuBjUkaiG0EB4OOpcctfE6+OeqOxvog
eksNOrJ+Bi0D6J8hLET7HXzDd3ZdXISlNltM0jBdtUPAlSGLh4nBlL6goRbQmD7p
h4TFW6N2HAmZvqrNXshbhUKUtc2N0kB0kzzdSfFqMPTOWAPXMXvdojj1KL+I0aEg
Qc1u94pC7nR089J1HcUnr2BXRPUXc3p1YXozIcEDx6BQI1BSC68f1HkO1tZNxuMR
YlllY2l+LpTtkJCzhz9IfvkFqv6eyfPdNWP4GjMGhQNYQTtu+xk2ZPtY7pHCNt4A
DSN86gy1YdeZI5Qg/fz8cqGFzaw7WSROieGSk5jcsDBH7u+IEBMyBrsJqawod275
BAjkcR/M3o3bDFifgSDFRCmxlpusPIavBE39J+PykU1yaYXjYhK2lS3BCcS/qplJ
QkIWh/Q+KdRKL1itSgV29ojSFyM1dKQWu4xnXZKdYz5qgxhFZTq94sdfYc6svkIC
eNCyvpiq6/Dlp4othBizg4OjEDeYPZzuMutcj0P6NAkw3FRnTmDpZviYaXnIzYRX
B/yNDcJcpLO/vIeYyBYeClx0YtFH5mrgogO1PvbzYWn4LHOaCZ1nOYvobhgahBae
LRs3I1M3rajDdrDDDBRuTScK8DX4j4mfG8aVC5xwT0VxRDJU5UUxkZ/s7ZN0gPLc
+pt3Xbc9YB3u9clxcwzwG/AqvZWw9A9XzscBmXXAld9rZyIHhkNjmSEi6JOX5VML
werzGSN49Yo7MGpYzuh+ifEFopylL+VPtcc/1YEmZar5zqd0F4njCXoFzBWK/EUI
c5H98FuR3cP1nJqBE+rI8GP2vdEEhDb0BSgoTQ5AL3SL82kcM5xDBq2+8Mr3dOVh
Bn2b2EzlD87ng5Wpal7bRtkRQKAt9lkxyVgFigOEnBh18dcFt/WhEcmgX1cnTT6z
gmvish9U6oKAmcO99WCqi27LnepWz+bt5Sql9WZIk5xSu5xJB7Bw4wTKmbP8n/WB
LW4u3tHVY3lokkJu2jv8DAOeGhGlKzBYsCfy8H0hka2TJljsOk4r4NbSpXv1mDCe
L1lJczYXId0XcA9QlWv1OiD+RUr3SKEyQIVdKT1jGL03cP2mTUBOLcxidbr+aHNP
zdYpvQ4kMwVwWrgXkviPjmIqeG/svIDU3rjivp/mrn6jabUlLAt8foOU4VyrHI3i
ZYK9lqkC365oDDbhdWB75C0jdINYXSS6J05m5YfN95HL+QYHiwjMfK18o0BuLPnD
bH+x20hagQqiTZMfg8pSjhdSvP3RihtnsIBlnbgd7ieIyU2+3hUEfeMFFne6fc+q
i1Pzcdgo9oM2ht2I0yTqWtO90ad5gyUi07n4tlEBjKEUqvoCS+11ao0iaPoyI63W
PunDvjYg4dnTfb1AneCDvLDw681RN2MowMgEQ0F0OrhEUuMmYgq/xgSXBtv+M4Xs
ysvbIcXcrVX0W1mqRIUATJW0MbqV6AfGW/IY1dPKM7O2UNwQBlSBiX0UG52hUcjG
Mxq3YI2n3I1BH9ZujeOzOo1t9ttBctXF/1OLFNNiVtnrzYp5r1YiDx9C2a2BK+VS
JOwU0ks7Olj6QwEvZy8nnGsLPooBv8KF51UYPVW+JVKZQSzBjyivJaWvEuybc3jH
EbtQOaF3apBDWxwbjVtTQAtAk3FtHOZPWrtii6ZqnkS+/dPzSkRC5RZEHehCsdwX
etmMkBi4RCusSqAVVVku2PNMoPcLpCAMbI6LWoaG07akdzT8RY+pwE01339u9Bw9
/0+tADtR7Xv9nxxo3v8WsBKLogHkMGUcT/aPzsHBDXu3FfV2Bq+1MWR2umMDv/Nk
dMpxgiQ8TjkeMrh9TtmHSxaZuu0c1Erfi+Dt+cZGizZkpwpQfyjTNE1ODmopF9dZ
2O3aac7BVYhdIJTyMfWlPsHiniqHwHsuPbscZP9KvWV+PXsRlpb+cL6qrwlhlVfn
QdQgpl70DLtTNsVZPqbG88y9hnfXlD+mbM0KyGD/pUQn50n8uwRS+DiRc3fZOxTj
pWJwHGT5hPYgI93mcW73MD9Nf9ZL6Lpq6ksCaw3hf4CXnTM6ioLNmRoKaFLvQNje
giRpPMe4oVS3JMsbzDWUPWUyP1aE6IEk8NXSSOnZ8dJSoDNKQJCCj7+nL/BOvlT1
h5dfWv3/eCyeNauyS7Qe/rlhJ0pKwENCNPiJujLmdY+MtW6s8+zhJQjFqveVtjFZ
g3b994uxDnFB/WEBEA692SpYFYbl9TUVhuGLPsjS+a4f1oe+IqUYZB8/F7CFjEdb
xEpkvkRWu2c3mcAO6b5VC4P4wE9F/Xw71iT/mpvf/0VAvwPisw1xyPZecjDNWHzF
3ukLMGPVHvoFu3Hn6VNXbY3faiznahiMzTYVEJefZqN895txyCydsjbyWeCwoY3S
77B4hx+tquaiacGNMrzB5mdQycFf0OARl10u73h1mzaehprD/CXl3M9x3d1pw0K/
3puKfAcUQ4oHMj/tLU0EtMi7N9DEMSR6SYbmnb9yDppwhEqunCMpnsmxbP+DV+n6
263uKIKI1YJQQVp1dM7edfcWoFq43SM1yD4qYCE0IcL4THG0Cwi1YSDdnAYu2qg1
z9Ou4sPXjlymqjBGFWaLChaZhbt5ykG5a9G7UFdprffzqtm/kQxT9Pk9P+wONsBm
66QJtm8N7zjVapGpPhJbt2LVPH0DmfNXj3ZO0mAa2viFTS+61WT5lrFet1tCp84m
NThnXualNluvYJNp1HddBun1M0QP3pWaLc6QXnXmhzWsRSiJzx4LewYtaFEXfKGD
155XOJ8duo3wuXYgq2R4S8mCNOCMlKOQzySFOIJNAhEoYq/WDxqM92VHI2HUbkWB
e6/ngL0OfZTHgi1f5HiWlRS+ypCi1kAyhdOzd8+QuoPixFYY5z+gC0f+BQWmvJxt
o/Nszl+RZ0OPVzaFH53UJ4D+JbfgCW2JeIb0QWGa6kDHW6R1H9OIA1YBrgh/+AVy
VceSTM7HoO9KMOzmRZAMOnNsEIq5ETZRmOHV8jT0+4APjWwoGY55ARXUrYRJzwl5
kl9SQ2mHMo/VihrudU6EhOClSC5i93Sy+0HkI1uNGwQTp+BpvpSWh0EZYSkvBD7R
Ir0SYDnQBaYDhurIDi0A8fSTmRzw+erTO8JiB/jXTWz1ltNQCW6vieJ7oaaGw2a6
Nk+25s37GH3fO7jmcZIcc2fAKqZn4aQ8XmZXfqnMveR28wPlJlpQ3T9O9dRjoe3p
DO5TX/xL6AD4Zkou+/FGtGbP7bpPOB0q3QARkjHrTOnR+LnxKaemKXUxN5W5C9Mv
a1g3Zn1NsQc/eZ5jbGk0UREZmwMpfPbeYgjJfrEVJnrVNP6mQd8jWwm7B1X/razQ
CmDwUXj6HAqTqZj97PlJDfX6XaS3KeR806NbprclK6Whwx7pnsOtU2q1w8fgT8kl
tGf0eN+U8P8B10Eu/CZu6k7amrgBVAY8R5TZ92vFZsLv5XMPG/dGCoYRS80lsx9c
UObGltSsqmwq5T65IIqKic2+THTw5BPBWHmro5ciRXFAh1x7dLMKWWnRTzrOt42g
pn8nCS3Y2cCA1CNdZdTsFE8BXpXGD/x4F2RZ/OywhlsmHLWK5B+DjgWwhINn5Nwn
C/Tso0Opht9GLG7B0N2tyNZb7x6lz+uudCxs2MZgsvX0/94Y5gMc+EmuU3v36i56
m4kG4iMpSwKc7rh9lzW9wbTdMQijhJ7Ig99Y5Y7rJMUocVPSc0w+px9mjtki3Gyy
reaueI30pnwj+2+d+6Vb9FAlKzUljTYmUtar/BV+y6F3sclKO96Fl2S+vSaBtrJD
RSJ8EmZKzIbHzcu4hcgYg1tocGteVE5lkOmiS/i4MRx4JprtQ0bsdxXFpL4VFT3S
Y4LAoI7NWgH+duNqFe0SKLhBEBoPPiMeG840u7EPOzJe9TfEbPb7R1giJHMVC13j
gp4ecMYOg3ext+KwSYvBDtpNmFVNQ0btwd6MZlmMbGKEjShfmIRhdVKXDLIhOTy+
xk54SNxVM2MNBXYUpeTM+wet2SlW1OpMLQWsWoLKood2dyB8GeQk6VcZZOH4grjE
cL1NY7lcpRV+Cl1eJShcwn+gS2GdOyN/1GlQYHgixSuCADLEGAzxGp1LPWnoA6lb
8N1QAXeDZli9ICZltsko73CFGTVUVKbpLOXGOi0R5Uk9NGzflMl+viUUfPzHoIKV
4krSGvoRUQrQoKMHGG4hLZ/lDoM3EeFAjW4eJ6Ya1ZEqDC6j9X9VvhRRJJmsmPHR
CLdq3mF8t2FNDuckTo0EI6kGBRsoQyrcw4Pbdwx1cB6FUn4kpVxSsVZN6htABvzb
lkqVlFv0xWPEQpVbWa4ryQU9nAT/h803pXD0I61n1BL5CjPx1VqKCEaczZ876VYU
W7UYtQcR6dQU4Yj/uNJlv0IzAHg+SVpYwA8K15ivHo0BdoYvVXzb5d/HYGWMbnwq
EswTNxSsPslFIOI6UCj6XLGFhy7j4STdSqSHQUnctY25DqcYUPQ2LHZr7AloYFCT
+5IZEzTUstYA153yg0ujfqelzC78gz6XwGJL80EmD7QXr1OKm//q18FD/WHuKiiS
0exOV/6b/TRlbKfn7W0vuv1sNKl/JrkDvVfWJoz6V4T5KQ7yHZbRhA00ZKKApak6
ker86H+Tu+xMxbfj4OaB3AaZX6pu8My9GY01mBSdgrzNPwcSWnWlpZkYjtG7o/w4
huKgri4v7hYKF5cgeeXzft3OtCUN4vwzwoQG0QE5aRDMqQXfueaMSIbnb1CF2sku
tCCEZkBk0yT/FPwIspYPEjwysYm+dUBaFeWrtFBvQBti63wID4acCKnsPlSvyHNq
7ZsBRkszyi0hEm0ophl9vAs86XXQ+FDjMZH8cmNm2tDoK/JjvAnFdk3ZKznH10A9
a5WcKyaKzehr+zkpatS8+41g49cmbbQstQwGTll+/6wetPFZ2HFBV0RRxVefh2fh
Knx7zXC7hXEJmSlv9s4c6ZCH2aBod2wXLpVaX8fquseyAyKtNb8aG7gong/t91H+
BFL7gvquqAlr2f4ifUdwmrxcTA8SmgySnffC7+jOIuCb0Ik37oZ8pTpH1k0c6FtO
0A3Z7aHVQaz/aWSgkeiJYJBNgLUqfqTyLfr8ZCTn+hiqdGqiiUCCNkLcpH/kPGFZ
zbdcrURX0RB0+yyc5E5IbvNwTukVZhs00CwScwx7oy47kz5M8JZIV0goLJNSuio5
/XobkQYhTBI4jENOS0CEn2z6e4F2Y0TvRt5HgZO/30RsgehNZHKTr9ZimE4mD01v
DUMzMGNT877JKrcx67r6DEJFwXEnWdz2+fGdb4sdLKZ7AEdSnB66oKUyOIKc0xsE
jj+FLYLeqPt0tDAK1T6bQ7/e9B0Ya2P24Sx7IwIdiZvRjm10uRh4qnlsRoPffLd+
VYH7BZkgStHiLIQVrxg4wPLU6hNgL35qnjS7d+szmg4cJ3WRIcuY6WXGeG8fqW3j
3WQjCq4tbe8WYZ7bCutBNx3eDLeeuotBaOVAzZ+KeMtKC9B6MwFSyXS2n+0a8YOK
sB7mF2WGyLV65dHrCJlWBLouIgFDHnPTX/9EWL/8PUZ9BBS+lO+7Tj9HI//5fgnX
l3ID2nP/2DWdeSN0+huRfqvkRwlncWligSqqGql5+OOsP6vR7O5mUOCdRL78mbD/
6+zTEcr9cAJiasQSuUvqgIslidQ/yco8Xcgf1FFsvoBefDufjSKjdDRkHp+6yj91
M44f+kZVAvSZdDgfeLNZkvK68gp9Xzv4Hv2AjLE0zoYWAAdeofv4GJL7UGjXWayD
cAou2p6pe49jHi4VDXt+dXoeT5uuwdL4eoau+AoRJ883NU0WQGAvLx75a5uV++HF
qlmUc5UO7iNZ2SNLPuz4MxtKpxh2jx8TGTJ9wrbB4vDjk78pKoTr8c5DYor4JkX3
xqkNnOLLwqGIl+H9f/vo/Z3iA+aEX9p+XEuo6m3G8ALnO1+AGV8AAZRJNpz4yBxO
W4qKd9EbDZqWTCZFcgqYdqMpo2j+cUl3W9Ku/Yx21+/Ftws0izBAxl9nud3OZUjJ
Mxph43Bio9equoxkso91Z/t0e2AwE8ZDt6/nBMrOCN/2cSr1iqxOLyL1H/81wQTG
iGDKwzTW/44wZlJKbsd/3pECrgpHHET0PjyMdQTdzriW9iiGIofzLF+pgNh3oXGL
wROzRNOIodLGKj6aCgipZwp00m9hMq9zSvmlIt7ZiAQANBcDoIBZZzspohe9My6R
qknW/lbclov0ifKQpAyrTnY36iuBCULo0kpWVaTQ2fqluE7AOmEDFcW47TmcGU1P
BnzhURUQ/o1zi0Nqq8wXKhxtsJQOyl3zJXLrGtDy0CtStPjtbLFEyBCXbqKK/e+8
86M3QAaHZKuY35H5stkWtywflaAC27UI/y6496ea/4qyOplkU1R5DoFSOdzAz7RA
3P2/9jOBIOW56O8Af5oyki8kgMFxfJoi+JhHx4TBk8wUhSzFSmii4qYVgf6t+b5p
tLkIl5MYLuo9HvsUEeGdTKIvmDfI3LAqvNZYipo8BlqYoo1jataTULv0un/uiHY7
HvbU4naJuRMmX5S9ZBe4vSPb7jSZ3SKtbBJE/ztuolABtr9exgdiQWWXMGTJrJIp
EFjg0jbyJEMF1qZ2SYuz7BaML9ZYR6L1ft3VY7ZXm2bSJ+CKjukriiPlyMcP86A+
5HSrvPfRG+2Vmaa0CCC9TnKchCURlLq2uES4+dmKPUIN9V/6GMEn0Kf689FUUuLD
bzodJ9Uu+ic43zYVlsF1hvqvcVPWvsF1S2zYjQIoeB0Sdkg8f8yEPCrkCerJogVg
B1KiDEYvq0wX2OYEOhpBzRd0y9A6aj9/aSdnzwi6/LHzXExyKTjNi+YEqQifPdzL
LIo8EJ8a13iapb1ccrcSXuAXHS/bo3UU274bUYYL1hqXFHy3wYrTFUeqKpQ4d2Gc
nyose9qtXkSXFy1Zl9KtUVl4/pEbqpb50VRholNw3Oh8mkLtSOt+qKj9XhS+9Wf3
QQb7mstxFugID89RJbBGkHmuOGud9f6kMNEdVynAeAi1eIuXGMfc8Pm7DcjiIB81
aqSOUNAjqAifkb27lxrVMKv2F7TH30l4JSRnVTyF3V+JI02mtpnEowk89PNnKwjJ
O0bPmJk9T20dVH6xL3XaJlIPcGZECtXXeXx4HcADZb2tQYIQ/wDoiBly0R48/X1Z
pQidRNWEXPKZ0CBkcbL8f6TyL9Src4MfSIj8RYKX3KzrZiE1IdKdugwjYZSEM71J
pTjMPV9iP/jMgfLHF/uIDjB8gaie4vNphY0uJtP+eOz2mfLvy0pQkgXoXE3zTlsL
gNF57jbl6niB0nGIdg7vBOReS/7w9NcmTpZcAWH7udp0KUzHFX9KnXawf0Rig+Vh
zmYqQySy+TezyEt2zQkEoibRu/L8GfhGjoSlzARk+JOBKbr3NP/ISkTuSmdhas0Z
HjpKZ0sGvPrS5qJD13zlKaVptKM6Hy92VLOKjRbQkDH8fD5OqL8vFy5RhRkv04eT
1kDZWQkwUFE0B749VbsIffarg0dZ2RZagn0ZOm/UuTjPTeMCgnJp1LaSAL1St+n6
YFyi3puf4pKBTNsQcyFJQpeD9iZRGzOKFq53jloZ05ZEYc7WuQXrqAi8Yxj3oCLl
RuoRWj+IYlafpKUNr5b9VWLHMtQaGsNI2JtuAvc1B3J7lqg0BS7iR+FXODAJBkBm
cXMtB0DmlR6hbOQmHV0S8wWp9ae3GNN6xo+FmjIQ+Wd42+uWwBzwgrUGlUxfzjZ+
Ut/00T3N4u5z4nrE2QLQ/58V13BPJBTRL1l/VUuTUWF0kR60G0o9vMxsI2zbFLRR
rybyeHwcNBSD/Ao2PpqCJAK0mqCqlZVl6Od4LOqeOcwRk/h6XRvqkwrpBQlzXKtn
y17WipviTYrTBm8fm6OPVmwHLAvgnXqhy23GXFJ1u9WmveToagaRM6u5y5VzNpQ6
TFbFs/gJUGHGhFkx3stuwDeLmhd71nlTrzXOnt41ZUa9enBL4u5RrUuNDjue7wZV
QykMOcCVyUa9xPk5AIlo7S12w8QGljS3jdUGHZK4MZDLqIMTaToQ53BJM6PPCCSV
FUbdR7mBwu9xKtw6Ux9//4VqTUspEUXOh6WgEqHWjaN1kbuvOBiHi4WlaOd3asDm
3xvP7GE9LiCi0IMUpVPmc0TGt6bzcHQ2zodId7yObDXgn3w8uJ6P4UkysIisb7Wq
dGHK99cnChzylAvYtN7gvH7nJCUrgcYuZcW9spqbODT/TUJZcoTLSqxAio5YD01N
KocXaYjwkC0KMClflh901p/6O8W6NrFNLqLX3SMCEyayEQGIMAVGlmtQqcafnG8z
1UmCqflIRT5mnZ8y4n+W0nBe6ByeCeQYCM6P58rW7fpiQpj6d4HcZX/fL7SfXZHQ
WsmOJd27ITdq3/L+VvsU+enE8LkThh2YNznkBSF46DM6eJzHvNs8aT0+AI6dm3WG
wpMVrLq+wF8hoVM++a20nVrYpyhVIctudmkvKZATZuq8hz+SFfm47M0vD9heVS31
hxEnAH0uACqM/1nKJLzLmsgGI5Sv+yQYje37U4071EtNFVUW2W/JI+NvYQ1cMY0W
4MkEDHwffVq+yK0wr1AQ7QLYMN6y5QdYJIa84ga1bi4BY3EU6RynnIM13ulHbnQD
u8SYoPK0H31UVAwStMKX1icZvJ5Ac3yMNM7Z3W9+SpRvAKZ8X2bOpoKjgHEWRiCw
aTxKnNEofOIwNdGpIeDMSNisufwIU+oYqfW55i4RYYuNwY7ppzQ/WYB0fS8DvJR5
wdjjTfWeQc7SqqIO1TnkZw9Mp/Hp+oC7IdUhyT07MjLO7AdZdzue9T5+QXwu7uH9
vp9z9yO5sUxqfgDOcma+un/hBhd8FctVh6JImH/v8Hgf67AYamUdnOW8oSZCI57Y
StPRTR2bNYQJ1ldnTxWMujZzChe+AA1SUpm93mdbtw2/YNjP2juwwUqhcuSZ42Nw
MNUthJ+mL2j3kd4MXiZiA5Fh+T4+nPNTpKhRPkJybxUW8u7jfoeGMNCQjboz3f8y
4MkDgeTSSaQFGN6cvX2tsMvUmCrWEaoiogj938Eji5HJqBJ2pGMBysFNjEnSR+6v
Bh0t5NUzs6IIeBtAGOIXbTQcnXLnOK4pK9rLf9Wefywpji14CZp3TUvA6t4OPtK2
b3ZImhpSco+jNnYPbsz2ava6qZgFllVtim+YMqAfslWucRLIjknltww61nRmlVpN
cdy/5S7rKYNJGMHzv4NzbiRqMYdsKwC7tI7qoPJpsJItYqr0wi0O726VvLQHxlbX
ucqTd+3M9oV22v6B/mtkDkrfkadxwR5tnIMHef0pYsc3CeJ0GkBmGjuGhNg9IJBF
1iFTqagIwxQh7YJbAj9Ntkmg9hMa7P318bJQerZPIUwJvZMaErBIZY42Y69OJHcv
QcpB+778pmEEzv89IMnWNG+dyBCPw6oVH8HyTCBW1fzRQMsvWX7UJDCYqkLVha6F
213gtkZvZFlhs9/kfXbIN0mweLLT6I09FkTGRJapcpTbhPc0j3j6MKdo8q3EygHJ
rtY0TwHVayLsFDbl2aZ4beBq/uEmtGbv4Co6xSwR5GFrd642i0ui9qGxI/iwIDXM
EzcEr0DRWQ5W1aCumaWdD9zQV1TDZ8Rye8nNRkd5d91WnoG43P0hCD4Qt6uHEvub
wE4jVrdbUY5Dyt8EPG8jCXUnwCtX7Z8o7ebOl8R7q+iKTSkAa1OZvVyZnVdJgnel
Hoe6SwOp9fl1gxpl7u2/tY9wHEo96e+hRWPecBXcYhAP+mkwVAHW9+ciYijkxdEH
L3yXJbjQhyv32WNEXIXrVy6gTim/Dff4k98EtYJ7h4CK89PZ59+w2Y9mav1TXZvl
S5uSOlx6AD62v+i5+QxqDE09Ory/bxQlg8NlEOBRp8JP+NC+DtevOLAGZuGCE7nW
xPyL0Zz0prjWRXUmh9GuJNPhbZYFKkslqIdKSsE6mfNwnHAuBEHGifIzOMq08Jb/
kY9YcS1qU0SLNwpP5XSJOyWnv1XHBSPx5r9NWYNCFFpl1a4IdslCJPQKg6Gjrcmu
BvS5crr1udv3TJVkG70J8ywVh6bdpjDBMjw+NOdKhg9sPICm1b6EPpIHLGVszgb+
f52RV9b4hBSYjRBYlUoVhOdHfgYEh16RCLrV2Ic67PZO6oqC9v0hiyMfMvI3EsF+
Bfx9Q0ZgM+kKck2RFd9AyQ9knNTgLkUcz2xzAGvpE/PWbb128mHkQ6Il3GEMQB+q
zzamiONtyp+F0a1X4hNNetV0DOxNMPOkIgLtaP5/G6vpuyOthpDEb5ZR2oRHUVcW
nNeb8r74oY53Q3FsjHey/k37G1nhkC8dyX29VsRUC7Le2Uedd4zARiOVcqxpkNIk
bJt+jrrpWnMGgfMlGA43ak7i2J6Q1Zt+63Na3avUBaB386h7jjZvopY6X7cp0arE
pmARH4vMibr5+BgNAfM4vqF0+XqiZhTKPhBVaF0IbFzHLTkj4advM3SPKVpoXker
WrZT9jJMfYFXGaVrNESPxZFozelpNvVEjtDHHo1n6h+38CguWlWvA3GG3LVG6nFN
f9hVC31/d/CSH3/qYjOdrW23RMmAVzTcvBXYZN6Fljc7gtiSCJ60CMu+4+NZR1Xm
HN7MdyjTEQvYs5cO8J4VMa8qsJ7by/668OLnmCleAJ9Pj+1M3S6japFbp72JiWUB
HTAMS+dSdsboKDq6Y4fbFjqq0CF3oukO+jshZt/sKD/79FqgxLz3oyUVw03zPE/v
/DZVBM/fI70ayCVt1lBfIUpV03rLJKgE4wOwdnJIAuprjDHM46Kk7XQfiVaa8zcc
4t37atHa198F2cEiBkbOYnb1G/bofbz0ZejVfv0pRkLWRwmGXPkdBaDXE5PYhrRB
rQO1eby1RLNSuNp1RX5aQy2fH5tF0ccOf6aOhjJ/Or7sD+kW+8DsLYaShqHFLx+m
fG+8a9AX6otJx+Bj/ts22zDFZNIZJPDSzTyosoSmNNkC1vpIFrIJ4ZybudIAdKUq
js0X0fYyMB1rFUwz0PsEmb4oM7csV2E9seKJLizXJIOolzVHomPWfu/071YRNzOV
hUcXo9Dc0LlutQtNS4OUfNk0EBLYZ19UBF6RyJhbOnNkzsfFpmEdJ7ISYstslXU3
U7sRc0EMS7RGezB6Tl1cOSU8uK14/Awqd2UNomQbPJ6mykbsUBLm0Wzm/iTEnmvG
rP4b8Ru055QKdHCarzjdmOLMtH7yHN24aEO44mcQAiTOtxoxH89GlEsl+4r7p30y
uVDU9O8AeI3PKlvtd8KBK2gTE+/8AQkKBo237Aortl7V3kXDXGy+Frv8qVm8SKX+
FiDONbjNEAd494nYjZv0932bZ/WF65P3pFc81XJf7pop1a5T6pi0x3sji3swprQe
ut/L0kEud8nCX6LYSEBjHTzg83Uuta1ZquACK+Sqz3jyOrp6VZFtMXYJO0dr1L+D
mQ/7lf6rb/j4s88veZ8wnvBv5f6HXsmdiUpV/kwQPxhMF3kXYdBT3HSwJyltQawW
80FQ/FnO7S1awqsE7Q6lYt62m3zIwkdM3v0BlaSy6UanVF5JwyqQCrLQUVaBpRrZ
HAnDkQuyftuxxzMAa1c+qpD34dHiMBZdkJa0ZaJSfFw7CCXBmIgLDzXedFJaQ0sg
HZNkiLU8/mjV/SoWIsogvAvLIMel3loetoVKKvHMXevJUESNuIrwNxJ48Qx2XkYN
LKrp+Jt72VcJFMpIDPkokD0NOLQa31e4lA4JhvmO6rf+OuHuvEgFttbUbyjOTWCk
KPvR8jmzmFsAo8dSG5Ie97dc2EulEaksJ316uB1gVZgZishr2lBrsYyTcG8XXyxi
/LvUllKc5YMo9F7mrtM9doHxSkX9UExrA1QuhRsaYPAPF7ZofJ2WP6mOnMPMpJRz
obywn5hKXDY2yWMpSpWS0j6UEA8uXhWYj2QySwoQWOX2WFETjv1wK5yNJAOmvBb+
e9jkPG5mFJbjCtLc2cC+djFlssgQVcTrKIUHBUk+5923LyVx2DV4OjLJU5i/Phk/
ZSSOZrnbhkqeOQYYHPFvygCMUxtjgU2HLM+2OTm60XffOw1OVqZVEoQ+n/Z5fCyf
BqLBCc/kbSdpjU+xQlS7akh4ifmxalIDuo3YDrsbFv4LLu+TPIoDXSAjtDZA1p0t
WwM/4j2ks62qxjrHhD4IEceEeT45aiOgFLdNl68JHc3+YZ/Qlo2VGyH9p8aXUcSy
3FygCoXo/8Ad4UVTUXHHMlqGLeVjYy0F9NUpyae+Fci4M5quVccedu+IO6XovRZK
ClctrStev92UOezGYApRur6PjWELmjE2I3MAHioQXB6nVmb8GQyUNQOD5B/pFO5S
LpQxmDDnT/x91WaEeF3HINX9qj69ZFYSnfhAVkI1kKyVMwWC1juvdb8o6WlyQxCm
Y2Ni5gnr6zoPYSkPJRc67w3C4TROZEVeZGRZ+ECZsVkShdYjfT3dvQNydYYdJEWa
mDiu7khWaNZ/OhsCro4JFdApN7yUQpYyDz40tle3qmEgatB6/m1os9rDjEc00oCE
ku9piofvu4e3+2BJDCI2LnkJ6/t4SOeb4DzjSy52QtKA4RfwzM7EwELD2+oLIxck
XeTmjaykvBFp9DrwkH+CIbQaOtz4prOra3MEi+Vjywd4+kOEsAkfd+GlwDzTcpw4
l6ov4rlGaOoCuVclhOCbfPPqLlG65vMoT1lUh5nGUT7o16a7xFBdcrtilYXaU5/+
voSCh5KEILLpxc+31If7k7oz5/C8hzGlomxewxuwNEVSI6fzaivLe6IshS/wJKvB
uiPG5lR6hn5NP5fWk7b7jEpQlwkbIYznQnICDGE7FGphOEZYplk7w7Uh91LMlhtF
fMpjTkMCP8QldYvYRoqkFvx77bHA0WAf8+k/+1A7Tk6Qx8sBCe70Fo6n6pXB1MBk
eS00XLuGoj+c9HCL04KkLXIYDz/CbZyJGialQ8HDnqy5e/OC0Gcu136cIebYtiZE
W5SryF0sCvz9wTKyMJppXBzqaP/hvWvFNmQAUZlkA0xv/ESw+tAiKxeeqxQRgR5q
tpsxZeEH3Ki8+ka2ZvNoJkogx2COCNCFH45/RVxZ+RukTAzqHko9Fva57rVQoj1e
U38NPQSihXCrYqbGcpOIWfiPAM6UtXqlQeFA0k7PB5btuH5X5912yI3/+1B8DLxG
c0G1Z0b3GcncU9Lr3qgZ92I4W87vuWjGkCT0XxUPDL5FfbzWrysGf3BD/TXUvrnZ
CTjGdynlWeib6QDKB9Xat4f0W5NwfKLKn8mca3HbrkgZTTCcCvVPChuoZmt3W8Nb
drc0leRLGPMhyx+l+dcR7fmVmH1RVfRHtTPurDsKTnsdph7DMZjRx0+tJ7MpOu2S
uMnA29dt0Jv45gCqtLhdIB+M6nRMqM2LZW2j52ouDo2n6S1SdMlv1t/YZz5W2eF1
/kITDbht8iq57f/KzXExPk5s7mpEwfvvt+GlZ79mKtJkbxhqXMnvGXgvXvgmgK5i
IlQUh0qTgZ3hsbOKH/MT6YRtBQk119Xz7bLS3TP4WxC6HGGqYsrft8zvY90iDFZz
chOtSKxgiwpy8ttQdKcRxqhaEGbtH2at4knC4r21oRtemmH///PuLHBLMThzu5Ye
+Wr9EGWFltxNVoj1sHGUdfQ4RK4Fgr+gbAoRh/5xYRCGcWJSiFtvybCHJiCTVm9N
4Wr76pj6LwfxPiGGmgVY9x091j8dRTiy4aVZp7JaKhP6A/Iq9z2uwonJZSb7kgdL
oWkfoUGusQed6Re2vHTcJv2tcmXMOiMWfXtZDhTboKYhYNEtdJbk7hJ8nXUC0tyI
yAvm3QrXplBu/UiUWihWN5+7mgePXzpd1bsivZItU4usxAacY3IBjLqsL0aF8rZR
HHRHSJorvzXtUZKgZmt8MElipCUzkjXyVPS45eyAp0QEQ78N2c4PurM90r3cu0RR
DsTkfBDwQVt1RGsjIzx+gZLSHVvm9zL4xn/Xe14vIZSFdJJL8z1pxrIjYtPEjcFR
7WO8+uDJEeTJYQ5xxcxxVP3rair+tqXAXVqRAraHFYbxuthPliqO/dMXWXx3MyPX
96Z4afFY0Rz26ViZBc9ThDAEZbAhwzriw0iXDJDym18K/9F5RKg1gRTdnT5QPi2Q
bTz1+QKQ9dVKvI84t1OCZLxDr4mtg7ly7b9cq2sd/M682/QKUxZ/G5NRZI7IWfdt
UiO0q21/VsAXPcXPER6w6cIDUsmALxAwB/By16f7uZJXVCyLXYIGmz1kg82ETBZw
dYemwzoOe8JKA5i8aZ9Ab5c17gd/4Z1ijHiZrFGfzXBoiRPKo1+IXhu3bu8R5jaM
NmabayJf34EEP3pGa8h/oyKbg/zErkNUr0I0trmsp2umZnLddHnpEhSYOpGh6i19
xXkTNctPOiy/4Bw7JnQ9/i//YLL++9Jb0g0z4cSAQl6kpykro6z1qVe+ksf9VtFh
9Tj2rgZbOAt2DNCrv3qbKMEdKRRW+/rbePo4MCmYkJkM7vw/jl0wx1nLfP0RaBBX
AB9cZLVSfDrw0WAB3UwbejFnEld5p+/8gOlsfHwMkZ8Qdcg9rn+fqEXbVNelxrAR
lnV+pkCEmOjTnnHcGPknpnB+XkMTFigcEdZvGNEdwGbPzZHGGZdG376IDQY11FlV
a1Dg0+nC5mX4k5neyekJsW/f4zxnSCqm1FIqlnpniz1ZrDi8wWUia6kIvewdZrU3
N/NSSQFP7ha/2q8SSh93LFCGN5xZgRHhrBamep54ZXUhzebtAitBZqr0H5YtpTie
TTfLvi3+ONUS9aeqvD7eJgeQxyyW7W8qVfV7g98zDPvj2v5LHHKTIJJ/raHhKYlR
0S64m+QbPtmYNtdLaCj3OCR7XU7NznPPpvoF05Cm+rD0uSq0lXNctVw5wbGR1B/R
6ji0RO2yntb/9JHCO01M1foU1YjU2WwPuNJoXM4sxCCSu7gdPlYzqxfaqTczpGVk
xZkgeD/SSHKOziZm6hCjoof9In39S2pHeeeT1hBuh+tP7MDTq0HIlpT8go9Dssh/
Rob2vMxCB0KFqXbimn7dYDs5isS2IJNSFdpcIeBuoitNyO7bArxK05LUgM+/LeyZ
ZN6o8+XlTPj80Npgi31L9PwgwbQ0ZRzxZ8TN04sslle19DUIJ2ox3imvCaJ0/HaB
6c4OFjrWg/bVs92vcRaxNDDh6OMXPAiAdYDja4ek+QJsv+nNCQ4Y8xjglrt/8D2g
e5oqZa/GVQC51JQKxUyR1p67aUbOv+mGB6VfVQG2lrhyDDk9bXcrdv50aCPUtd90
EjftM7izj/BeOBCzgef0uqoBYg23jJrFZkYJakOZkdpPWktQQL0/0gRhQqHMMCYv
n1qLlZIuI0w+TApVW8HE3sQgP0OWrpYqJEB2cbxfN0MSYeoogf1WfT6/KbWcrkbA
TJr2h8KvB7/ddH2Bds+c1pHSaVVmyurRid9NIlKvj22p96apxGbdmUZuUidbQcLV
0fPmoYl41+Z/NfUTIXnEBGYFHQJcNDHeIxnmyDH0hoi+yxZzCTaoTbZcAMhFXMGY
PCjZoWVcRdPQc/n/z1qYKAN8JaDe+FFD4ArlxUQPhPri6GJIQOpvmB1A7iGmKyc5
lVu59iqvuzWRvQRfyPDYh3W3i2EyKNFd23MXJF83Wk2vVPG67R6YnjC5o2QwhxoG
tBLEzQyxeucL/5EmjI/LukP6XTk4E4IqKBOWQqsBZUGc1hhLGpDJD5VGwIUOeiWY
L4mwfvDnFf78Reec5bnPVPE+zhnVebC8ADTNwFJHZErSbgJUJ+RxccbvBmx7fP3z
Z8y/iz9RkN52fuH9VPyGWLfYnC3z8MMVZ6AweWeLqafgCZOp1F1Uf49b0kuxW1GS
FULme8e8wTlqGFW7dXOQF+vRcp6dXBBAlvE5gaKe2hKk62i5EH9DZ/oNDqueSqpT
T22fAuY4ACMbhqFmGI6gjQYr2B4EGWo+Nwuc6rjdjmSD8UNTJ82sibNlW9LbDhPU
Ha7mfcgqs3m1Xh7/DmuZ/5AN5ffBKwbMNimgtojdBMs5qv3SYQRMJtyJ030BgZsr
SnIdgX+Wv0j3O59O73We9qbhY0vDQk11OCftsaod8PvPJiqqOpai2BgDQIbOqiQc
5dUzvMyUGQcLsYQsRrRbuK/HyitzT63egY5asVnnDHQzS/VgWLHMWppUv1ofbpXZ
z9ow78TESDEPvn9OXZlAKiq/P3lnnJNSLrlPr1Cw12A7yOju8scNG9jK1Qwom0kj
j5DUm+jVoEruPhumb+ztj4EDpttiPRFFO9e99G9HYoltCgHhW9Z8tdYcl7X2z6zS
r9+YlnTRoI8J8/MP6DxrDMFNXPjUIXJAn5bSdw1dMC3yBSNAfELRfULPnuhLvVR4
c6ykz8qAJHzFSGRVcorKT87t2DhmL1GYDwJw2eUVEtWTy3jecLYbsv+XdnA1jsHs
PwpXm1BsxVaMpYUFdEhV/ol5kYPcoboYKGc9MCpDlwK/ybXvxy6PTPehbdSNnS9f
u0CBVT+A8986ozSOTi5p/Un+lSWtv6uE3KxtvHP6Ywf4MT34hmItg6iNyOBL/4A5
/BP2jF7V964mUx6dh0fjWgDG2WZM10B8/Y0aQPkXlifeiId+tUSdKHksFN651pD4
DQxBV7wywkAv/fDX1j3Az+X0+Qdlc653ZgN9X93IGxJ3KZtQSe+9P2mNEY1iuLSd
aMwnysnv1REiiJqQN6CCybV9r851pKC14ZSnTjZp9Q7OgTd+6FEHEnExBhLoHuvX
NLrYb1NZHFRz6PeSD5Ru5RyAdJHRgnyDJo9xEnR6qrrL9tDh9K7gSBqvXR5TEySi
/Bu2xtmBzUqwB4zfLEM3nqEQs0VXiA4IRAFam3GftvgiOfvSHLHvM9U/2GK+uHCM
eva8aGyRbQzNkXZV/UlktQlqAXFBBZXCz33b4yjDPPvn5h9VDll3J/g+Af/SSZ1s
5/TM8N6DVNscLyAb2obrbxowslM1cw2jusrmst1F15qcSraqFmWuxHjbkCcYx1qB
3R3kmkJMlsngVcMfDVJUfWCQxPRfKrs9XsGpoVSGjD6gnGdPgz75Qxh1FlTvS2Ba
JiErYaDeoAk8IbZvcq0fRYIfoglsJo845Ke1dTwWOrnLIhweFVxXv8pvVJDwrAMP
67xUpaoGWxf9dEE+sbnpPtH4cdp8hzgMVE6MutF6rER6Nyji9ztPNLbeT7PBM702
oWYYMj2IU61LTGfOcUHipRqqk9aMeWTyTfL1/dOuEnE8ZC90zA3B2cvXtoFX0n6H
QDq7vuWjn2b3sccgu8hAhL8Cy6gqIOUKYbuBu64CRY3K2iYWj2Xt2TdjnPiRHIKH
4ZMSr3DByY49XlbFfy0WTg0FoF5LzMmtzUH4uo21AtQKsw+XGhft0oUcbv/74i0X
XiSZarqIGSef1Uhv4wxHjZNE39wum0LeQqB5BrHu/dH8p/SG3GzRbxDqJJkbNd2d
ZKk8N3AtPeJpZ3Uqt8G1CqSxJZ6b6jR03g5woBSoUhoN0n3dFrEn705jOSFfJtm/
+3cQZTcYowEuqkc3BH3QaeqD852VjUxDDhUPU5Na8h2/+qBE5nhaZDSSMJ0EIonX
pJC2AhAGYkl0PGLqm/ANTVrYwfAzNZJoFYIG5/htXW1Fg8ItrygtoZVIG4jf1QuP
V7fLUFxAX59tgOpvF3nat4Plr3Q+G6+t5HFIB4b836eXDeM2Shapv5/CBvAP1TGS
Wk4+VRrBf+q3rfY80uVNi7nLCv1j5YAWoOzp492Wl25210NaEpIqNJ+76WCWNKNk
kUEp8CSTtAj7bJZZmspe1toPdc3TFlbgwZmbl+oDYRxCaXlvj859fG3SSIeG3Qdd
jRKXQtZuXF+dJFN0fyhSQ1Ds9iHRtj9s05rUrQKeNvCHG8QmgpzVTcdxyTiqe/c8
9k4GVf0JCUnVv5JskGz31sUaM71XLw934duo0u1U6HsAJ6U6WEl9nQ/9jXGIf3HY
trXWlUSLV/W2myxPODbJ4xFj1WXSrwuQu6QjItXP/RD10QeaLdPka2Xu4E7B7gNI
EogOHMZnsdv4z0di/cGGYlsY5PlUS0D6dmUvJXKjWWlCkpTnJUFoXRUWqCkNbiGW
+t7oFEuBkU4u1OKjUzkZpO65l5QvNynIIDzJOEd/X0fAGWe9axhHs2lHT75bqkOC
3mEqj5xe40fTiLeawtXntgqBqn+HEY4KkkYR3Y42xd049gShPftO/jjHtT5psUvu
JXTK2ufSEwYN5nqKZ8Vjpht7SBaeZRkB0LMT8Twmy+B6qYCdJTiV52iptn8rQ6+l
Nh1W0CyVCc0VWwlj6APkYqOdWntkhjXt85cUNETF2B41GYb537Po/BAavq30kcLS
aBNVmj3x/cviAPGrvFKiwj22k+wKG/nIA81HB4i6dRxid1DuiFeHFDMj1Bsu280L
bULo4fd5K1ODtgFTcDVt2HKjux9wYN8U3DZYSh8ZtdC45fIHiJDmccDIP4kw5yWk
hq+jhaoWx3k2Ak+8GUjABrIXLMJRUDlgdamupB1tPOzFCffIfPe51B8S0YX1dk6Q
t3dBpTDQxH59nj8yZZFxhsHhCiiNr9gQ8hKN0ObSCDTUATgF6TYzvUvFAEjOaGTk
/tzvYhBxisIF0wsbPyTBmhrHy0dN+k+h/sGV0mFqo5Mq1veMaF91fP7roTUr/tOb
BqENca30m/57dLF8fJhKHpAGuaJfXXGFkJldY6sDmFiN/8mTVY2gg8ibZssCkgHS
b/6XeV+lx8zr6x6LTeaN+MeOngwKOc65A11UCCXH51lr15WuqIMo5X9ui8a39aLd
BpBUxb1hBLOAaEfnLOp1+ptgnfMuswV2Ibet3dO6h0aOBMhcjwNRUA38vkhqcyFw
9sJNIxg96m72YMbJONNl9/xWDdQm38rArno/9C0KIKBzQV5YNhlJb22PO1tUkhKw
B9R4itik5pb85hKhOhP6lfCBfsXO2GV3xpQn9E25CDXDEThBQBYUyjuiIl3yVuTa
eUvtk42igJwu3iwLkYpjOHrGvSnCRVS9I6RfM0Y0lY/s527gI4i1L3GqfGzJpR/2
r3Tn7MvcpaPKsQvmMw7qA2d32//ghvzyNh15G+NhDS1P9pn/L4c6x8sC3ymOkgv1
VC7F9sDvVBVHXpquQ+Z3OX/ssm1JlAD4MyXCT9bWhKMRz3GRrO72ewVcrTfZZy6i
qAl20omW3OhoZ5gsQ70gCsFRzEoQjaR6RE3QnFJ0Sl0t/hXiV6ADKu8ud/OCWYcB
pqqOoYM+wFMMXGbn44TWN5Ntw2PLZiymsagbSEjAaEE7cngghWocqGMuZbT/euBG
ek55e8H+XP9NK0q9ECduHbvvvHPSlAGuauUkGm/8h0/GcgK1AwbEVqHniER/NxTn
RMk0O5xqesSnW45+n1dy8kRloy1MyCqbkRoGph1qlTCFd+uNZjnnXDXEGb0kt6T4
OsbfLjYicIgzLdVj85Y5WRXBiIEYxtXaOpelofDa21H8LNLhMGrjGUlKR23RzlXy
xDSfxU0Yi1JNqMnZEdKmMXxo3F3mwmJaf2zR/hRK6X4Rct6nCzZM6YefZSKTTCVK
NmV9qnefLwsjyPgXegBnvaoyGa4GAakXld8cRp2D7WN942+O0MoYd9/nk8nA+mXx
wacTOhydgeynsrx0QatS/ckxnMKVCG/G5zQrl9c004HaIRnbeStOPOK5wov3w/lv
KeLiLFBcJK49HXzvvihK5XFko4DDQNcDx9pzQ99a9iW49KVAKcCxD1mEfkyGpJR5
/NBKOk27fDU40gptEOPBtflZI4X6Zo1F7R1fO3p0EAL5jVgR+IWbnoqA139KiuD1
hrsX9FONxPhp3ATcqAJr3CEZC9Z65ixD09KORYgklUmmsU++YWEmTPWXOuiOWkVG
o1Whvf4fn0ObMTLYnTjJu9lRIZVKa8iyi4xL4Jv3ZubjwW4O1x4fteJ842fRbGUi
DPzPO5oaK004gzG2SPlOG7O33BERAQqme56xLl1SLsQ/7nNMRPTpHSLiLwmWP39g
ra+gB3ZPzlsa1P7KiJP+G8m6CG4U2VzeraE0U0ZfwqCSRuQI+ib8nG1PbiEIbCn1
ALix9CrpXDvHBqPbiLUDGEJfCPYFb9M2VpljbnU0EsLAXi+TS+88jOCG/gGZDkKd
QpXwDIrX6HXLnntWZByBaQgkfepWnWEsl+gZaPHy+fWIOankZfBhNZzcfFZnuP5a
EZymD1qBxUgdSQRMAHSDZlc47VuY1gHxXfpe9o5O6sFV/EL5qhm6YtRgrieKVTbD
DbwNw5YaVByyuKViWEpYpfbE+uSj0Cc6OriyAQCB8iS5CtSNsbEmb/dfsP3Dw6gk
ASSXBzd6znlEj3e7GLM5TtmLu+Q7ZPp/QfsooTzqB5SUg0KYe1pQxpye6xUmPUQx
InYG1L3Gz3w308qtRNx6F0nzyLZUjPWL4Qtd3xZ8VsvEgSy4azWKybSxt+ynbOLk
xiEu0P1kb6ltIebOhhzG8L4HbPdfBgH+nUS4B6+foEOJ07F6EmjmX1ZNBekGPIpn
sJsvCRmbNiurhQL+JbonbAzx98dXzVLZkIt15AZR35bWPT9FycWXTQPq/LY3+Pk2
5B/4FSDyHPQDdrdr25CPNmud9D9IqYAZqPeyuXI2ffJ8ANOrWdmoHjn6saTTqxiC
gakrhqoSpvyeYI02CnfsHoBGtIyR1T7u9dOwt0bC8n9r/UE4LVKNALRk6pj2UhHv
xg88o7eg1/zW61pBcNYy8sfdeqcQBIcl1NtQzDVQpv9kj30b5jeecJNqpmnV6ZTM
OXUezf0KI6W/+so3gYqqVzDwCA+yuWYywEnWKHVQLewFVtim6880xeuK5/iJ+khT
TsMDTZmvQTQyLqWN4Kk1kiqpYtdl5SlC5/Q9Hp6erPn167D6lG5pOmBvhOcE9nwt
xOhinTOpSXWRhMUbOqmso0etx8ox/0/fnI8OCdYa28znPCDU09hinIfhI2DA0EKN
YO0u0fL3q9FVwQNuwQOPF+KoGzcBMozTfvSOQItrig8wrk2VPb3pZBQOzdeT1ybD
ShppI/iPdxZ2I0mE7aX9oKHKakQ44OpI2uSDhnH1v+IfcBdIKdC8XY7iPnm17S6S
mcgBk+rle/43DQseSl1M21vhBwT0/YSBiVx4QHaaH2L4Chyd+a78aYWLYOjHlKJ9
+ntPf8jaA3z4uRpu2lmkW3xCKobdA39mtJZqpzVWHHLuJ3k6EbJ8mX4VRkptO0Cp
52RWW8CxvPSB2pAwWQZ0xE4NQXWs16aoo05X8OA620SEDi3poil/wjhvWSnzLbEu
hcpe1ljHC+sbuTNallovX686RpTN1ky5ukl0IKFxZDqmc1K0kgZaRC9lvqnAX4bJ
hVEwgll+vuhE94mO1oFCBu9Gi9osKdcgJk1Yt6w4fXjOoJ4fzSLG9UdG8jfoKzGi
Oi7kF0RPBZGOxzvj6fj1rzj+5cslVLcrUcc2An2xRW0QSHol5IHJW/2spw7hyMFO
wPA9U412NJ3CiXyPWU50eM4QQN+/brbYkAo2VxBRvUITRwHbwHm3prRVLknuhwDl
RjVrQotRpXW12kLC4FyKpCHqDu6utkpHsnNNcP3/TssUDpLOrgodJ9Rh9g0HBOPs
9FDE2NRf2uH9GxOry0KTy4GmclEUO5Jjxq2xOlyFEAGe+d87HvkOXbDCuPW8MXNU
eSZvUILT2XBCvUU1wwdS6WyFnq7fR3zc4dHNMxEtNNOi3rcK6fVLngosgmCf0YYA
xOtWrmEaPkpjwjwmmkDEIDWbEyDSGR5ggIUVyHXsQJc6emp4NCIC1951RJ1TLYNF
8y/pH6rgOz2WGke8XsqzJThAEMhv8mVAHcm9jP1Pk+kocKEGdZAOWc7U4oKIisES
pwihAjnCUtLxE0S9Sx3FeRizlr9lLeeG0eWiSPkPoo4IbZmD3z0O0HQlBZ114sx+
JQoqNAy2t8SIboo6lsHZnxoYnVU+pYMcJ7Mg5nSftOOjv8Sea/W+k6+UQXNsEtUm
Yc7AkOKF5E/Vj6XGFgfBMhrTe8f82lGQo2iuE/ABie7PWFzG4t/EsZrfSDOII3b3
UT8kllGs0JjQeDPYvBJJSjGipl1lj/tgRA4AM1ufyOMwGy2kfBq7SIBgaYCrMfPt
h6DivFucXLo9N4JT1FAgkaZN1p1qH1XJrmCw2hykMBXeaDuGALIdeV0lORWzsNyx
NekEvDQYhhz6obFebscBXPnlLhPJ2jhNn4T7xUmH0isr/JnXhDLWAFxuV+I2rVkP
SydyXDj6TSvFZX/OhJUhdL9648hXy27KA9laZyelyPP4i4F6PfEAY+jKR6HfJHGt
4u6BWcuoVXWH1j0nMEO8K3zOnneyrhU0/nXSLrIc7uGEBLjwQEhsHILp7g2lfqHj
kEuYL4jEq7dL+Ko+JgGRsPp4mSl4ceHqzLrtEV9UpskWMCYzf1umbL4+h1L+JGU2
V4T0kUWTDZQoOp4sV7JlRMGfh0re6VnNj0Cr6H1J/OxtpqPRdM9LCS+hHOfyAuWI
9zzHVDcsviWugN0/Ob0n6Yq8WMopyAROsz5FFVUggY4Gcw7bRbR4OFjiGneb2LFz
VYSzGtB5KSvIagQxLpukZXAzuhzOuD4EHF3kIcfxYbvxm/ctNTpU8BevhFa9l2Y3
HfTlgqylwPBv1u6lE5TMBqkGglhIeTgWhfTu1icFWS4aSpR/k++ohfILQ450Lp7L
5Fo12+AeZAsZSaIz69NHbfA01N89dAwO99gqqcO+SmNUrnpad9FJHZ08X8M7uEqO
wet92/WFQKkWpHgD3eN8gnd7ywFQm5BVGe2mC3hyl9yQqJLTQk+0FK9xnmHHOHS2
+xgba6wvp19UR+mY9KaCbEte7o0vF4mc9zhsXuqmSP1iLT1MaaWQsnQRnHvX3Jpp
CBuhy3jQpNAgEir3ko5aeYh7EhIulvQhvoHPaCoz9kg7OGo9uyPN8msA4GoRxkt6
ucA9rKxJXMT8wP2a9tzSo2tPEs+42RMBZB4ml607CFhRn8yw6N6JoD3v6Nvc5Ip/
oCJjkY3nBZOQKVLC3e5LDERBiq8dLnpqPC+d4GOJXFllkxnx4FFeXbrCV+lw+OGY
6oaeczMFzkyvRXpEPCJ8trJ06gpmN/6oBGb6p8nEhF9SKUG4aqkmTRP7IqUWjtdP
mr15uOEut2speQavdV7ptmGWa2VO4FOw+aQFz5Xo12iuTXbAv7U8UdZH8dNg1FTl
jgqs8sEizH/9DoOFndYd58z0HDXg4yEL/3MY6X3jE+mipC4k6GjP8CyhaZQXGDqJ
OqAVhTTcc4+ky+6CcMMbjd+2xURqvyS+FfoqnNElxEvp6GUNqXIRGdyD4MI5Ru0g
OKO/7iyoQU4pFNgBNp/yoylyiIjaB1Le78oj1HcCZ/815wm5+Jj22qD9CHKaN55J
LNUHDSOwvtCL/TJgFp/KmbHwPHz5VkhmrOxVQ9xzBcSp3Rc0Bt0Z4nKdgNHQTD1N
lTSrV03f2xu4XZR+04flOLa01RTWVf9pBaHPqYc1cSdFpFN0EqqttL1pTMxbZcBZ
tIX0DGzze4376O00Wtt1XDzlsZQPQjJG24Mc6ijFB4JX2zP0VkInTTCjRO0KgEO3
Ct3hHrKiHpO7zs0m5jGyplCCvSWVGg3G4QrbhPpsBvoudry5BmAnxyGFmJATauRv
4DJPxcNHoObQTn5avZW3baL5Jah3wdVyR0AWUT6KyFZdMicD45B8ecP6hrMTT3eB
e+WgrqLIz21my2WQvvyOlIreMDzPEGvNTLLfJrkSPh8FBoHCEV7iJ/PNdWO04FkO
pHvC0QFIo3k5mWJ/t9YltYEiaFvO7RBrfz1n3DDkrjOHnWrnfW1Dq3jCXsaibZuw
OcpUno+pmr9oSn/XXqJM8pp47t72liZbHZQC3Aqm9Z3OEjcEKSCCC4TyizpMy7UX
FLoMGhNKJEUoiAHz67tsUm6Dbs8rGG1I06mDzsqQwbPig8jU1Bt+1hNJefyHCmmo
xTVnygUyS9/4FS5BHAA0oVhtaf+fu2siXKiWWxWGIWchyTq/g1I2Lx4/G96Udgqc
l+poYRX34RP3MBoxpQJCQxLn2pRFYgMnMPZpIPdbQeWEL06Z+LuzUDE6oZEgzFvW
PnwB5I7c9Y1FFjWK6GnXi2aspFPHFrgc7QuW203a3i/j2QTpQjHLp5HnfLxIquZm
Xn0CCMlbnlc8V86EqwMYco5eZZhhoQPdY5Ys+xM3oE8pOlhzh5CxQqkkAavhBhfg
PU1RGG5u2iGt5L0jZGzTEULy7zIa3eEK36aFSsmibDPP2oQgAKaJ2DGFnY9LwmAZ
2ql+QVvYOgfkWxoSIk8tjpy2kPz0KAxozPRJikqsMXaS7TFBLhlTbqB9/xn6/WKt
0ko0SEvAv2Sdvu4mRpzOZNurzNNyxcjFdDptHXgnLVclMERkUMKzxcDC72XGycc8
H7Kbdkt6vobSsSE8z/gIzn7+2rZhoIcUyOxJpIBO4B0iAqcYg3cR09PRZHC5m0JE
ZZU3GYwAkgPoLpvAAsjgj4Mpzn6ESwHJUjGEv8K8Zj5ts2J7KFKPSGflXnCs18CC
3hQm0UbEIXQHI/kVh/kUk6UZPvLQGGxziZIgYy1+fnDMVhT8B9HTM8Zty1xSpKWj
XV2HBCVMEBTCy4nx1+NHuf/TJYspkeBc1L3UPpHCPYMYELdrQe8IvwxCwNt4THSZ
Qp0hKemk3N3RCeV+aZC29JHDWg9z/ayKVGh68NP3SpOP35iQbdqVb9e/2wOHsbm1
zer8xbcrFZ74wqnntc24HQeobadXzC7YKUixZrlVj+FKec1QcmmgPc6xEZJdL9B4
w4/3LZW/cweZyHbgZ2xpVs0ofbyc3Mm+bF4nYCZOZ4Nm34llLllKSdQ8EVyq7Vbp
M/51nXn1vuJypyjlslmzJm6tK0OyjmU4sOUD5IaqvWA80w0qxYgRQuCQ9gZYD09+
XJA8KwIRlynZI8S4NL8loO6zaw+pdnQaXjEHnom8VctioZdI+D68vP0cW/2hMLxw
ETovjheKasZRVozNAJLT9xfq3DcQZMiuSPzlUusCQ1LZPpitpcsKyykamn3dglIc
MnhuXDIkvyTXQBtK9NVtMaILNy69a52xdJKFQFrXzl+GN4/3jIzxDa/a/GQBcjTV
3e0Xa1aGlyW9eaczES15dmKReB5Eym4JzgVTTRH2v4D8HyN56/9gpSVuTll79OvR
qtBIDxOYsW0edgxeXBsum2TlNNRMwHk8Khx+EViZKKchzuWgIMOCt99PLTN0oTLL
HPFP2FAtdEbyGhq7eCMPidnqxKMfPDYeoLELKeJ6czcEsMX3OXG/eLdRHHKcS+mr
SOsXw46vA8FEDOJkKCA1HSeZt49Re/Fh0Eg4LvFagsyhvzB7eQGno4dfrwyjN9Yn
bInN9FXixF1omkr+15buCo6U2hYHzoeSnX/Vf0Y6RLdrvLyi4/TF3sWnXl4/NEUl
YPbtNXNgjxuJPym4kontoLv4LmDMfWHOF2vHL1a6t14KFup/P51ZG4fWhKHsWFrJ
YX9wP+qLsYQOgwDZKFitqnuGZdPgYITPBn3limw95aMKODn5hP7XscHHrshFtaUj
knxTktLUCvPZPGjm4+/ek8mjXxnVlF0qKwFdndgp47wTLDMGoWje+f80tbEwM7YW
52NmnAwq6gXGiZ1EvM7ymsQJOk6Fd3QuPwMgfGeaKIP8h02Q1YHCrVh7bfOy/nU7
FcWZsf9Y0eEWAHcZWzQN2H1jRfP6D80DBLAVXy1o05Q7f2oky+6hVZSP7F4syMnB
p4oUFa+h2bzcXzdRykfpPCelLRV0mmrKbxwtY5zpaG3v4Rv0pQJ9NKFDzgrXn0Li
eHk3Hpzss3dzhru51Y9kfcyUWSC01ZXR/UmKgc6XA2ffM/3ZKniul3HNwNrGXSh4
FT5DP8TBS1SvmN9cuOMwzFpC/meusTyisM4FTnzZFDUpj/5DAgQ3Hr2B3UF92wKq
9sfM8p2mc3dwthhFsUq8BVhlELa4dqUVslC0LwSvHwqapIiFnf8qghlFCFuKVBQd
cs5zCmiBuNISLZQAgS9Z1lnL6cpUi9+RtauvL4IOsaRGf40ZeiNAvbxFHvQqEe4F
clCsFtC09tUxM3bzpDNEsKgurOX/iZtuxPhE1tGJphKY3aCZezMiu/sPeBi/G5Q/
cePo+5h9iqV9KyM4fY69dmhTNr3b9tmtZjAP+KiZhQti43tOMmf1ocDcNis/LgZ9
g/IzrDSfvqBbPTyglYMXiDOdk+8hajFSFVm+Woid/7CA0RbidDvMLcBen9TWGQXd
BVFbItQApKERsEi3DFbsYUhyFuba0Lyt7i46lSIiW6fT8w2ZcQOjyGh496iGo9n2
9aq/rLHUzFj/auWSJ6ctDg8mFBlhinl7oHKSw+Pwddj8ZI0DMeQohyDCCNLPoYEx
pKbwlJVYAvAdqpzV17kwI4nhYRqEl8rB7CnxrU2uPuRltP3Fu/mzWBdmlPffWD/9
Dj6fVeZRDglRZWfUgoFKtnNm17J9/YYkBaICWAhkD/DVllQtVwRD0KhBshGrQxVb
TitEPLWv9VUX1PrvOkMQ56+4Sq+0STMmwrAfC3eKaHqEouUtRnfqJnmiuB1faALo
M8uDmhKlmWOdwbBYQ/Tao6kVpRbnOYtdu3zczo2bx7xHS4VR1r5qg94uQGgCk1me
se7Zmqyz9RLJ188gIAj585JrS/FoU7ssaoD8wPejGAi7NgoSfNc4607qQDxgogJy
YwPfSmbG1E8EzvKs0FJfCaD81s5mG7Kl93DEV1RCCxNaIQoMW92R0Zr50hGp7eeN
N7DEXpE8xsgAyqQBKN6aNlTArQM9RuheQYdHwXv9D0aHcDSCWeEnY65BzdSpCdzO
xlTTjCKkutaXZMLE44M9yB3R3CvDJULVqw0JleklhOO3QgdG/fRYYXIAgtxzwV71
vf853edixMkpDn8fbm4bRM+qJv9NKH1spu1B2E1fKpkzZkfcfegL+hsBX6/wBaAd
pc0OD11C/hw4vTr5swbhYr06Sya+qpljNWzm175j+r1DEaMsDQlO2uRq9VA6M7ux
xWwD5pOTW94OWLq9WGrMQaVfXCShc4xpxU02+QNWs69xQ2V6r4PihOSZjiJBegQn
HnEoCKMqrHx7uWchZMnmlNS3F8RSPkTbfbqePyQs7y9N0Kx9W5A3ozWNG36LpdYy
147De3MYEP6nK/LpLBem4uTBEZAu4Ae2JXx36putzzcFiIqu7s9nL24trbiu5gMW
H0s6UkxYRmdQmfkQ9q6hcHqHp5f67OK3718LkkculwToQxHAx3M4k/RWRA8/1Anp
hkivH0VBsa3LLwNNQeXu2gflXA8uhA3zP5NVWlU262+d1fh/JoY09VWwojm6u5Fn
vHlkQKjb0NMjR35E2sIgFA3Y3/IW6CHSpA+BbURXtWcgLDaGukFzVsLmlDL/imlH
seRNXasoSp64vnc1YM9SQQf+DrGn9xb/SxNQiGay8Li3O6ZerBGk8+j8i0a1Bckf
5xOHGBjTRH08husrEdwPAx3AlX0IgpsO9aW8RjL1gJliBOXzTYN0U8c0LK2yGDu9
6ge5K1PncXuVoXCEwI6xo+qpW6HHUqVxLmTKXXXCH7njBzvFewqCFRTK9c4eFtwL
7CKH6EoNpbJX6bVGtLu6KWFP9Cw04anUq6OO5IiWfz5Ho75m1SlK0UWaRkI+cgpz
p2nxP7i6xpA83tyQl2J7LF9so2eRxzSq20hbmxkwyoDOUiyiuGe+67HHBoXTUPrY
DRwhCVfZWrQamOxZzv1vIP4TAPaO1wlI0rdkOjBe28QVGg78rqw/iBe/B4/Y+CG7
Ge4iMRQDThqSCfwnXLHghtbAkbAK96rt56aDmqBWMTAfMv146Hh8JgMYrO69DY/6
DZJ7jiWKGroCGE95jWVapigpJoZnkKouBZFmw+VjFglhZjkWJKEtmxBGz/qd6Nly
XYRxiiIrKb03M+YMNsxtPaSaa7p8c18LUsx1N3U+Co71UrsmAhLAlt85cJOQeGCi
pHt08SdeTbZu46Uy0TxQ2CbV3OyG3Po92JEOHCJk1X5AIjL/HzKr1ENe1nn4Ogmt
lkW3+dlUJmnCqACzKUyc8oVRlhosKjXcpJDqq5AmFrbcnYdVXvL11ysBcWO3I+bP
f81BTK5e1GOMaQLXUnIrjdynhBpzqtukLqVrBM7/hiwS8xolqxWPnMTQXeau6QXO
SojGYQtDL7ipd9XCRPGdah3o9ugcnUCpnJFZ9ybE8kUMH203RfUiKiuYSxZeGJOZ
l+26S9dUZFUNJc/KFFw6ONvgxAoIZb+lexTP074DJabEMEqFfBlTarGS71ndLh5L
3g9Wck9nQu5smWYSRCLHcFmj4QgJQUmusMCJ4RM7rSZ82/ibFBL7AYfWfAjysXkK
gP3A5SeqbmtI4thKscz2+CQm1tTGUjU29txmKP1WPNrcxe8iz2Q83R7rc+3AYfnv
CmhTrsjJeEyGJTTDaoUA/KH5MUDfxNF/uMTxPOVpX3my+A7aO/9b7YZdzB0Yt0Rt
ihpOOPYSdUhp2O6GUIzqlpicOsuOmmF/5GSewVp8gpVigdA4eH83+YmUkE9Ik7k7
ncyo+KFQPDoINC6SIUHUZMUK1/SRQeQyRMt2C19Y/TZ0ZJ2yaQGZuUeGOg5Rm0+y
cdlc2DQDQ+FFuQZRVC1YvgBQMYuvV5Qy5Xb6rZ9zRt0m1jpWZzMRzCNy8poRKydG
FM4QYvBwe1ICoJ4kJMVBPV3A1LmyMTC5Ra0c2ebBsmgT7M6rJ7a69rZmuAO0JR9E
jEReumnPtRq/2Hmtu8bTC49j7ar6ulsBGfNJ2y0XCTrpobIIaQzcfcQcGdEpKflg
pG6cegc1ISCwwHECywljNEeJXqr67oye83cK9emvygL6hdxYjZKn1Iah+kLNICkr
tpS09HgqMGpyDC37OVXIb5mXtB2W/ccpH4CgLbCfUdwe6aWKKfg/OgY3NfsBTaWi
sqwWlHTDzRBEfENJwam1iGj3R/xHgvtEDfbqRaBQ3/XilfMunY5tJJvCDrxtmlzP
nrwmUXNM1bl54JyYyDwljfj+efLeAKJcKKHVJFROEF6zgOZDIag+ERTIma069MxJ
JZy3HyWIi8qj6yaC/iDfvTTov/XHwfTjKAyL3xULLnAWvVbNYVuCItAzZ9XrFsCN
FYGLd5C6+EHwVS4RWWR9+5am1IzEbZBLvCnF/iAAnofu28rg5SsXdtjSbj28AA+R
hLGipz5FSKbvTGcOhI662RLbY7S+le/VrsyNWc0oR0lMOFYKH0Wf+qgMJpYXCcl9
mlKgMvDk6IqBGqrHJ6oNaABPlI6iZ+z4GsBoBEOZJFYuZa/4EkJKQVHNyJOktukC
H77jGW0zxzef+XmjS2lHM1l1i7xxhRADVDNblTPTaAi8uiDyeT8ceJ9QhRW5OlMR
WHJotVCIHqz1PM+OEObKfmWeUuVspRoBRKDqi7ZHmVjC1yYMv8W+sTrB72reFORA
os7q5aey0jdVXY7fHmGkm6PPPyj8g6GKIE4Vi9GBgHydbxP/VsTqDkuWtROMxRmL
pZlQdS1NI0f5Zb7kcENPnm8+0/bSbieD6un5V/b5IZwDU18REv1EiBYEfNVQEsHx
lUudVA3xug/OlXvw3muLidNiOT0Wo8TjBsBmBa+zGwowHCaUR6wiMrAEhWegrOV4
dy+UAQkVFy1Ir4sC21PnaozHj01o0VPgBIOBARnTFlmBdtM1PsNGP8HxHwhxKdwx
G+l/6+UU0Kn7GwLA94GWH6arvlhutZmNGFYctEgQec6+wWv6/C5O3b96rmnbfpz5
HW7Co56s0U6c5HbvKRq0R0nlEVrD3ojvFQ+BItE+CoCd00+p4c4DUOCqc035ZgEu
7F415eRDoCpmkwi6HPt0p7XhdfzqsMnpjEYTNZ+zuKfmtN1k8CCW7DNiB6FOHMhe
05zrkrdXJw9Jr5OeFJNmlC5nBTPzBCMGR7jezM4Td8lTFYL4iWFtd2NPwU5b7WP0
ERuFE+cijpmQo7koRKQ7AygCfBBeJx5KYmyvnsW+BsgHVY9f5J99HPP6QxW126A3
ZYp2LtRMGO5bt8IrjzT1kG8l4Wq2s+FydyVGGyIWLi9WTueFa553wjFo5qe53a8L
X3kgc2Mue4I5TWhqqaMvOeAO8JRSoyGq011xqWlMiC3/YAB4mH/L4E2nOjbnVDO0
jrAlZoEkTV0Lp/vje98v0ACuadKtFZsZCw0LYXGgM76MZ5rLoevimPBOatiT3aZI
YbgUUTO3z66k2Vbsh/3gTEsq3WsQgU1dEUReMC4428ljojXa9OVEeqcrwY4s+Qpp
J+L0XQvcpYtdcwxCU4J9dJaiyvq+ju6zyjHSrX4QBCTkKm/C9y2YHFZH/5T3xxuE
/HhNdF2FwMyMYuiNuOQbve1EdBPpQnLEMHRvWoOSAnV6btakgL2eKbyB/wwUUI+z
iBgNEKXOSTW86OupG9VyjUXU7PxNXxNjTOnjo+vph6T4FdWft8Td0E+U3+wr1DQs
+A7UJKgGKhhb26wH2zsIgFy1Zq9G1xbDRg5omapj5Op0TmGi9fz0FVCdp/rbQ+DR
dfEpEE44cdoxUQ46Bi0zzEocHmHKfnv4f0gz4ZU8T5tpR8DWGbKLWfCWna77Sb+X
wTvW0AjmXmgr5Kx/l21KRgk0Vq/h3+Gq5BpKe5rjf/sHdEGFIRR6JHS49gPAWhQy
nqTeHvHoNeTvs/w6lEFelC3KbOQYr1/zfmevb4Khi4/Uf2wUT2wlZX4tS20b1q4O
9+5JxoJ1BMz9XRztE4Bzua4mhfm3Cuokt2u7wWhMt85wlBFOXVqp2wfteEufgx5F
2/svprAMjEErmvZBDnL72mXbuBdpE5DzN48uTpB2RnAAp1HoHfObXAvfKKgDgZl7
wjA+N9O9riS4rHOhSlRnhQwvV4XKAlQ6IxFV+3qOzW5O2GYPDcLnYf9Z8nRWg17M
hoYFu+xorW6g2pjBbKeA7TUXLJN7WfM2ETAlhZE27u1Ssq+h2O3qJ9bl8RNvwGXj
XG+/FIpMzrSjtFLu4R2DwfhYb94iaNS1amIf1U4wCMBz+oMgeLg6uVm8hddD4OwV
ROQaeo4zntRPz8ShsZlxO6vik9s1C4qJ7qVmnnj/oXxGrI3ip/clTWybJ3g7wYVe
/uDZhLiZ+e6KrBEDL3IKeVGpAkDsgYC06TN8XkNmGCfTBLOJ7wDwXqJLuibdD/OJ
I58wA3XuPAfgErXW1VkhMcyMKp0CihZurkWkTzjpIJp7vysMRrmq6uNOaY51Jmlc
XWVSr+WpkHSXcE+JXb7zBq+sin+W6Xyp3ff8cCHVt+mBgYR+8wY8KdHchkuaI6Sb
cwrYnQsCX/c28XxGXvCFVMHMWf6hHUSc9lQH5XM/AEHBf+PS9KWNyC3agbbkkA/F
tSWZ0hKliPLS6tSt28prBHMA8aIdAxgI59bhbnP3EqvVoI1oYYJ3e7cVO+/mmpi5
k80+IS+WtiEyxxPNHluwJeEGRr/pjHVcCKYYROkOj6xcfUiy8NnJTItyhRptTjVq
3Cj2f6sQ+0vgSF0uQSnNR6DABNe73ZIJ2H4AWldRKatyzgt5ozLlMCFEIIJtjz0z
B6T0DYdaM8lwgNMVpPblkD2zIZHfoHgiZYNAg0xDdgZ9+XHWpz36VM22rMqZHXX3
mL6maovQqSlWVUW/FyNB+4kg8JfxjcbDa2OzM+kHKHsPNEx+1hD14UcqZmG4T6JM
0+q79zpSp5yMOPM9rLItIVBIqTXNQYZvVfZldqE6d0HgtfsyLfUZXxYPV56q4+wN
DW72e4BwrOX5xtfHlsMErgkLIQL36h2zXVYDOq9M9Xjdyn5L3NBTwM52qpWdJ8OP
S4qwIPYe4GNfRVNOBmw6nA6I82L6bg7X/jVsmTm5Na48Xxe2fw1n3ETWaODtdN5F
kpUAgEDAVJYrAywIFAO+JA+XaRTidCeSgdFxfsGpi8yNO9KRRSARX+1T2V+jxz0B
fby+EHvlUHqFoamCRrYu5ox6KItGD2P7LfoMA3KZfe+5QlYNKZGAdjIJW7lT4HY5
8N4YpLj6JQzPcVgLoJfSQ/YmR5fH8svLBTfAnywHXoKOQ5u6W1Y/gWncPKLzPYoj
Hl8bIz8JtqD8ozzzuK4MRKizDgk9TQng4iw5AA8J/g7K0t9zjf2dDBhEAYpB8Q17
zh6eU4q2sGZZqKCQFIi7xioSu5InLVimbvR0avOhSMSFEPAgmGoGFiQy8yPiM/IY
8xZCTWYjNP/FqeVwGUsyoClskXFADudXxsnQn1q8CDFmFFoG4RCqqlC7w/9DsuWm
3mH54JwU7agaBoyl9iq0e3PJteT1dpOu6uySTOzp0npplgBv/DO47VZgRunTHbFe
0KHkro1MN3y0dsXjuVPU8HJZuo57fz+3Or17/IEwbORE9rjp0Vd1UIgnrI5aRv8P
x2tD4YSdmxV7DgnXB08JuFHVNodUbJguL2SKueuKmefsEv0eo0dQ7wPkYEHidrOg
UP1xwb1IehgT8V4Y5kWUFVXn1ljKU5clX9naylharwSUnLVBQavDPXio+EenNKh5
fKvAStF9MKZYr1OIOk5SDgnGKtnQXMvQDqJuLSVE30D4sutuUxNkP1FcrekCAEl8
WBcAvxRuu/+gUVawSWe3eTYf57xoKV4RWX4hZe+WIo3QHMCfZw+YqGBZRghh0zGn
o+5CdAxI++ba2XnXYPyJfm36zSCNQ3udEj5SIMmB2UAzMYbxa3jVC7Mp6Qvb6sSH
KQ9hOc0d25OfN1HfdVvQnvuXNNL2iiey9Dz+y13UmSN6uUSE/Wx/OfPutvC0brEs
flcXTwlqTUhf4EJaPHTVKIqzB9yqIuRv0Kq62jNL+64klqLBZNeGoRl9FiWp6xwI
cnCLLInGIM3Gk9rjgQOmL68Busep+haakZ6PTo9GZ/MN5WJ6wwUq7R0NQs7XX64M
y2IB2ozSjuKbqYeTHHMGAX3Hw7Hpd0AfwwDCMXD5YL3FeQ9J2gdhwvbkRN0o4Ilp
bs6WVrcgut6CWa0J52p28YaVOO9T6zi9lG1a/uDAa+YkoRliaZsC5w9aqy0k1IJH
gPR9Sun7rm12LFn4zWhaVDHeo+1P+FFdAcfeHnWMxufcLoFQ2b4mAt7mLFyNnSCQ
s8rt0nkXxsVgM5IB1kd8px6qgCidHO2RMVgwQ2pq+TR8QOjGJal45inWa5ad5ahH
kfxKexPE4D3Qg6M2jqO/NyS30kufTkbENmI0lavLKO5a2dSK+YZdugc8Q3QTwn94
57jBSXpY7A2LYJWZ6kmX2LoAgSBhLe+Sh5j1PLeolfQZgQEi6FZBR3u8O/6YGPVs
h05aQp9ATp8JUZ7tKCQLf0RmV8Dv6mGB1lnu7KtUfWL1ckZvmLYCJO6SNIP+AF6M
na8gVho5VB181szPNtZ8Gqb41eqpI5/OB7YFmUaNjaTFy4dVEUSlf8ehuy/VJvCf
lAj3v3sYMcK+rmiuLXc8TX5Ru05ynjWlQeZkTOhsr4+uuX/VgULCMQi6eB65tMwr
AkMysRrhjoh75kJ2/d1AF9dRzp3/flQEVDqh6RGlTAMzgAmbo7SNi8HwdGmvvqcL
5s5Jw0WYci9q5bPAjhmIs4b2bl6DjGl68XMiuFyas1OvsvRt7UXTtOrtykjPQxtl
0r6z8E3a7hVt4yvy9whXZzXKo3hMpjMEZ6aubyVQC436BFrcgmVQFIEyWNciZas0
/mz3Yk1/jrpC37DXGP70fsm3BKs0JuGRxWzONoXeEzaf1W7UFC38Go1tp8AX2Tlf
vVA1RbeHNsj0aKxx3C+5kwpbvcOyDkPPsZT62b9qH4i+LNu+5X4Vm70Nd5Kib8cE
n0cj1bz9g9Ok/rW686qZ15y1r0ybZZtEoGvG21S4/s492DQNwmIHGBEQvJ/m+9u8
girgytonrCRBVwDkXodecSSw77DuSNVLY3b6fFD8PzwAwaU3kdYdg0NWqjKU3f2V
s9FBsF8gVg6fAZ2TUFmU8GHQ1+BUHgLQMeno8edbUMUoVVN77+xLtGRxKvk0tstO
s08DSL36f2+QlxjH4SSzExQ0Fa4TC2sTXsbVXwxORke3kNPXTG5IE5krzRzwD3NF
7NB/dZ/nrgUFCm+ShEfSYsa/UoJp9gWO+xz4aFRxC3iLMSs/B9eFaASQe0jt714f
Wz5uy6LcapqXbds4LHiHunHE0Y1e0myFiVt/op8umbnC7igzik5KyTEXHcBzxLUo
wCl0IFZKNvdq2x9zao0sXMTYaLEZR9Z+X5oAkZopYLS3/QyO7tnGwwYtz3Qe040J
eBoTUWPlKECF0tnu1w/3gjOWdRGEzX5Qq/XTm+1EHvXyhSi5d6fBG+u87Vatw8Fz
UpGo1F7p+JNVPOXkpK7T6vnYSxxZK7Tk8thYtlVcOUG4I8bHbgZpdEH8T4L/UF15
uIR0AjLVh6nYtShN/11ToFfiuLFLLNa5Hfp+RPG/mHvZjTnzvQKWMihzDkGRE7YG
d1FXnkBVSlPObMcm7MRgEZc/xOTY+ZDA9gskZhLiIojJUOvCVOGc33s1IUOjdaDn
j+4Ya8AGc+dY7gtYDExQjHAu2pz2BeJ3+JAQUEaRAKDPjgPsJ85bR7LR0fV9RH74
dOH/D4lmWSPQVSAmNeMvO3U6KugOb6cJzLUtuwuJnok1+OAWo9ZRufVdYJMm0PEb
uaoXViS84orqLrM7ZfSWJA==
`pragma protect end_protected
