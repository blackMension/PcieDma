`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
isCvUTIzSJ8yecmnKrwzOHGAzCwtQAr9YkHhtgteGVixtd4AWqcbCkJFOTe5BQ7Y
V4240Qw9NQ24GhhwyPf5EM3i1MAMU8WBw1ctvbHUVBAKhcYhyLCDUMWJYxavrK/o
hkSCUR9LYRsguC5nzHIWtEV7ATzoA0j6SCSZ7Vc/5Ck=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34464)
Z8WR7jY+tx961U0LxMCu8HxoCjh1/JlHKecnAOUlXmne9H8fKUovSzrJKr2wBK1S
c69dBjPnTemV+WFNjVzlubX6T/UsVZkZ1tICqf2z6HyFK88UYrvVTIhBs28DJ7S9
+oOHJtfEYnib/kVa+CldsO0q2zWwd+EPD9AqqhrNxNAzu3fmJerrao59n5/On7B9
YNzERVDtqVinozLgnz2zkthdgowNddtkOeU7td1y6fCrvSC5BJ0VN5Cb/23SSfiQ
qWOcfvb9R0M5u9KZdaeMoKZv7fPgLInfS4CF9GHnlSdEyb4seFuN8St/KiwpmPpv
Wi3+dY22fVlh5tpKeofeI+I1OxJmkPeQB9+zfCoEWJRQBGLuqDl2MK9xTO31bP4x
ta8IC22/LgOEpzFFWwEsvpsNjmYOo/u0lNqLnWi65B2gVOWNUGj4ocZPS8W5xcCc
pBjcv76Gf1IkmVHJvik4MyLr0Vf8xQpDotLSrw1Rl7ymyU3T+j6O1ZVkoI7in7ZU
hcWSQQSDEK2YVd8ACTOuS/o3PILAWcGSR+R3oJ7Nzbstr+M3oC3CnBqtO5M1pUb+
UBOUsisARnxCmNAe1I65E+ijr0XmhLtDr1V/uZol6ENe8bJ+YqiS3i7IPpIAdGBc
n3nTpLG0FMoNObmwrLEPCxEb8nih/hbl63t193PTaxU7CvTUnxeLsyGW0pRRU/re
2Y7Zc4w19L22v60F88qba6MqqUcm4L/0Sc+pY8CXXpvncQ4s4p8bdM2sYm0TCjlW
r/KL3L4VOuNWJRbgBe9gc0fBUb838ptIUSY/f3DzyA67uknNCmTX/Z3k5GLml7zy
OA7bfNEjgihWuLdtFBxZ7OoN7goC4vg+bcUt22BPbnTVNcdyAsvSurpJFxZPzz05
8BGnvI7ZfuhwCmJRpQlOe7FoCga9IJR4fprtmjE1Rvo2SwPYnACSmEs1G345BRSH
1dyIgB9DEQx/h0ZlBMeZr7f92uSQu1/ds7NcTUTeF1CKA9fP+uQ1G9Mgjn1c24q1
Am+G9YDMXnrf3L/FXsWA1jbFGqvYV9GNKlvmu0PHP++6XTEbHWLSUNY1XLcm3jHu
ZiXS2am7PiZLGlp2n/wL4a7SCJTQ7JpBZ5hjQ+QRzrIS7+fMAmPNGmokvuulmSrg
nDG0j1WOGEblbLDCpHKUFLlJ0pvKnVjO2Lv25TIlOEe9LR3QqUn1NfiBQofk5R3c
uey6CGbGktLVZFfrp9VGRrmhQM2d2Nx+D6GMUPkOF4uVK+0/zrqiZbud3l7F8Exa
kowFtU0MxcPcK+a53otNDwsjZM8YhDpj0ui7KoN1IVGJEj5GPPwRwVS/NXwSi7PG
EvMl7+kSfBqB8IgB6zfvkdHZqNDxzo2rGJwOaicSlSwy2FCoGr9hIQ6VANz6cex6
EnLVuLY5jb7HV0Ra5hgIvdYycvSaON5+F7BMb9Sg8kivj068/W9hCqcHCxWFbO1d
2NUGUsPu32KB5YM1/IA73E96u6uV9N4aEbfoiI5RF864TAFbyLaJNYlAipJcxFpN
NvLAlI7RV0iMHVat25+FV7q/+jWoZBsHKoLAq+4y+kUEGEvfcBdrz4qNkxevtlk9
sfGkpGDfcIw/uTtdh9TAgwIFmcRPbxKP6II1G/uhvQ891W0WJs23iKJewLGWGZur
DPnePJWQzIfIXo4gYIGRJqBdMZxuIrzl/OuCbJHR6gY58BaDSgNQKQnPultDeztJ
pXANGALsaOBNLo763rHWdaEsNuN5h8MmDe5s1I8VNlX2667xy4+q/rBRXpnyPRh7
Q+YrOZRQMC8bcXOcpTah+jBI0K5tHt7iFoH0F054Tg6bcCqi2VCDl1u0BIhsSZ5I
JGp6gp46UP3EE+twBaLP858eABtOS4Isi0LIDfjMaSzK8ysrvGJOUzJCVivv0YFJ
q75jR+QctqhR1g/VOhDJffumQkyToLhg2S7s+GFJWr/LVdsGXE82zNSXX/84PIV5
mruz5+QNnQT8CGzYYR4405pE40ecFIR+0fL1roVX7PCdqDzNGRZD6Tft439VA6wz
Bsg/WwaGpft38CpWjFEJPaefVZjuToYlxo+G5nHMpljN+URb1sJY3ujjzYlYD/gP
+Ne6dC4mFqH6DaysLva0ugxeuk1O/Ut/Pe2tM/dpO8Is/7gdiNCG5ApQ7vNyL3Cm
0Q1WM2f6VCtDtPdGezHxnMlTYCiGTRV2U7pJHarE/xJ8Ugsa3DAV3FyRd+CUM1P5
Rexerxso/YDokIfPewLTCRj+Dzm9J7qXhgXu9McPwLROIrfb2igpZQCR/T5SpGVF
nwp1xa3VRCPvI4t5V7/CfTPIPyGHGOGBXu4GvH34pFHOk755kEeSexTBC6Nrxhri
uGOhDxGv9SSkA9gFc83Pt5/csigIjEUJfiV4EL3RObtw8Ds50+xwkUbZ2Nto36mY
VGbKmIe7UWYhy5XL6ePyPUYorvqleSzW5TDnWjZC8BMrUdVZRgQJO5b90w0tiLGf
vX9fK6zoN25XBJEtYmOCRR9BPGJDKdwK+CE69P/QyaAmr0UTxIEPStIlAZ9X7sSy
2az+xMXsFLoC8FmtcI2Mz0ELfpz9LVb4aEPEh0nTKltebIebyf0nEv+eqEwspwkx
GvmTtYJs2ZcSknwl0Brlw+ukkdou7gnNj0x3AHfYvEweSmPvCvfl78jeJReKVSeI
9RNteQL+5DeTc13aWQUuxzVjUJjzzhnCysvY44LbdLBL+1WH3l8lG8WScOdjCWAA
m1daxci7WEIGbO7kcsPlvn+lHw25IJYsqcnfeFKby+j+vTLLCos2YwSHMblx4HHP
UvLQM1buJjFAxUA8DBOja5fRTiL3FQfom+4+uNjG8d1sGdrFTZV9Dj42tczkRN5u
/+SSTG4NHBQOvkfIZyofF6Dhr7BO5JbRhzkehG4r37zjgy5q0ejNcfmbq4VQ1SE9
7UbAsUpakbuHHh7c7QkHbWTx2FICVvQSdF2YNJQUNX4EO5mrgeJJk7gVQHr9udwb
NQjZ7+KK5AnbNz2E0DmNWNQoqpqTVz8Qgq0MFdfseRMUFzJ9eEQnoPKR/1OuMQEG
Ms4on0wWIvgwHWbj6cEy/N9f2aTvBtsSZeLG59Ybso5dcn4SOPJ0FxGd94Cbldjd
1yto/leKTYCn6UulbS3549HG+Eipa8H6POzrctBnSemIZGIlu1SpeLzQyPZsknD2
YiMcbhlV4FGPZRpPOmhqKtim7Fy7/bxZV+CjqiqQIdAYscQI5MgoSCHHcAtulNAT
90gVAFinWb+iSDEVvgdyNbP4yNSqq6bxIYscc29KnuhFOt8sqpsA7EZn9cubR4RL
YtJ17DXTFnsiF3k/YxIgwOJhOta6QJMRJcacJI1u93EidzLVTTimV8mN8buslFNC
LIXm3kks5yVi4DTBUVMX29rKXuhIUWAtIF+0Ui7NhRC96fF+CfI5tBbyiumdP/XI
dU/xOw7dDyaNyieQrtcnF4whAY5uTQcEcgicdnTxdfklftbWD9Vc9N3wsdQyjnMI
PRDao5TIdBjzmvnEmX6gkzOkIoGQA3tJER5mkq8sVO35/w59anqyED/vGfclz7aZ
+4q3/IIeGjd0y/0g4rJWYPwngU9A71mHt12c9H3KH0MnorCflgkvaR3qIlxAaFjz
QxEn/FA/QO9Om1EaIVoGHbJySSTChNNZO3FfxbXPrE58s/nKUyBVPCTFMC/C64R8
MQP9v2A0EjVq6wfJaK5mL36isNAoc3kCVYvQ6hhtBmAfK86pIR1gkQwSBtZyt5Fe
WPBqcA7rAh0dZxwJTA6t/M+q2yLO4WXozmsiOamJGOtrmj5yWEkDelB1lphM+yG4
E+zkWOLTlBheHhca2isE4zSWUEiXgE1ZvOjNyTqAGnmhWFYfB1DIQCA1alWdbK5S
biSquMyvvewTWbwlarVWKXJlL1GZh0/PB5jsCmmc8hz2pt1/mmh9kr31cSSbXoRc
u9hdUXDl8ndOTm5Fq2yvsSC6fj7OXfTEekHgkZBO43xkOtT1n4Qv3Xkmri+5NBAL
+2Ya9yUwuBNprkywL0Al2ALqBZ3EYUZTguuJNd2l/swZ9ydPkxMFpeFV0stmu463
0q97XhgrI9HmIbZDwgqC0J1Qlt8aRuGHY0CQB5WdYsgdjOUY6O4yQm1vdx7yPyNt
KgnUefLPG9+tfrvf+jR2RIg2tODcvSYiEmwhxy+DcshZU4L62xrIgrFuhNIh5//J
481tPjcY+VPN0YH3nJbSt/5kfJh+VfHVRTS8wO5/S2sgFVF9uNnVA7+DZOFTfV7o
xSjTK/d3WqJeoApDj2kH/pDbqkjox/81RSWXYZMgmNWqsqnvn6jsE1CPjjmeMQKo
wwAeQ4m4fa+TB5UpiyN7mH8utlHR9nuKok/k/MS7q7qB/un/0GtlUqslgEz/p8yQ
wQM9MB0M08rW198ehP9PSV1nHPJMpLLQ3rjrhSUcbEfIhgHbMCByBnDxRKXSbPL+
JL18AApu5ewESeHfdrZMM6c52FKJVv1Ksk9ghBzNi41Gbkl3ETMkkNV2O7ASr360
hr4hMg+T1na3FrUaUAAkgfAHCO6hdtUlFHIjHmr8TN0a/RtWndT9bX/KzH3nYWUg
gSNC09KxAsU0I+7P54FskZtpE/Txwi0cnKmRVDyb48sXPhh0fy4DYGsw6fIb7/ac
bpgVYDvSFRRsJ2Llp0XSs4en/UGA+xJYNEMXkoFKF0wodoLLB+TGbT+vFjZ5gEld
JHH7i45+j8FiSJHKmnzeBGw/HL+IzVgyd+J2SN01F/kbmFNxG//8hujiym5HVBir
ZC7Q4PtZ9jHGIq6MbecnESdXfj8EdZ6pwY6V3L65g3ouwCVXTbxXjVTeedd2jzte
K+zQk50lEhF0ZRfp3V4yYLZou8xij4cAnkkXRZKJxmtKKHbO1TVHjN3HF6cllgXK
TuntsA/pRRLSJpLZobg9zaVtvzHUFfRQsPUgP3wB4FZkxcIi5l6qbD0mWXLVaRur
Pol3JWs1eSYwCQL8WpCouUdmP6836vwD+sqHax9fAFH+9Q4+rS/vPGJtSbUYl04x
i/8oFYQ/4qgh0GxmcT1HMQciGD3gjA0OWqFgdscvptjyOS4pCH5tWZ0feQNtrWxd
cp85DxV7Mw090Exns5eKMWD4BErV7P+xn6i/ll7X+1k5Dz5a5j9oPvImKhhQP+FB
JC6FZSHMi91wcpw184s07HN6tjUOPc+N+Dm72yz/XlAuD1J0qW1JQ0x5pAWMAY5j
qJZn5tIW5w+nbeSXooz6ykt+bZC+iKsc5LNX+8KNalffeBLViNEW3XpSuZZDphgq
t/NITid+KPxP7iKXfF5Pwhz8FjUvhlukV5uO2g+XCU7SU2OlRqw7PENmU8hAAjY/
dc1tj7hWi9LTGELQ3JUgyWBDfwq0MoF/YDdavQvdvvxTk38e++/Mc1LU7UOVRAG9
oClhnCOIjAi5pUbjr2ohqhECF+2ZgWPPEeux+IlITWKJey1R//oEYESBvlM+JiPf
aOqVqMi862PWMYbq4T+mtWT+mU35v2uw2IiC5zNJRWCpugs15QemiZd5ghnPR3OK
siXdPsbVLx4tJ9jb/Fa2XSyvA+T9ZBxyVnnbeY+DILn6iSDBVtCBgS0YTmMVqxwI
T6KiCAKQfcAFf5XT/Byuqg2VHh6duh/EWWbY/rDS8qBEOLo6G4wYXtxTA/ZpdDIN
3FadXaac/zxRMAXb/7F7ePfNY+oBKClNxDxbeLl7Cjd5LPqzpc/MBvX71NG/ZBvB
LsWve1jDReyUnQuK2xjWU6cdTrrfANwwx+1BM2n8ZwJaf30uMyNknhoKBbpRRyFO
40Ujn8uSLLo9j6sF3lEkO991R+cRlJcyEOmkpOnxmRrEVgXGi/HsgUrxHsuJ1FJQ
FbhyiKq0Op0fwI34JBK2tyVJciKe2Qt4lNITEPiFBSZEFEWYOmsY45s+g1Jo1fW4
tHLser6bslbvQ9+qokX/OQTYCY/iaiRIMAN/EvNppDhPmeO+51sA18t39sWGfsOt
AST3AN8eywSRLBEJDMQGHnvPeWqjzv1LUCCgv7k5IweJi53clnG/owxcz6NQGr6D
iHK29/EBuifCYWQjlRPJD9gC33J3eZsWGgKJTfT5x4YAYkIoGhawgacyOsOSAEr2
z2gI93ejIhfq0TmKY+h/1RLRT8G9SP96yEfUeR5e3r+7qtS6b+x47l+IQ6i8QouO
NLZQALL11GxtiCO0NyF8LLEnQqMmmQ+9qewN/GqePHbrb0lCIneR7sF1qduiexUs
Sm/zSb2cMMfGcmMCtfe+3q+3341Ny/7D7QBUBDYhBgtf7kFa54sflYyY7at/lZrN
1yIRtQNeCjpLN3tPV9MgKOAjpkMdcUig1QzYBD4IITJ3PYJb07BXNTnIECEZAygr
GTRpqn2zxoJgkrJXQcI831d7qtEiPytzSYqBCmUsaBjWODlHfpiD0BZiIkVf2LKL
UBAF10jp1lLSEHYKjICbD7V2b2WqEBxz+Yk0q5oLEF8JjfjcHKFC1VS8CsBbv47N
8TB4mJ78Rlef3HAI70ql+7Xo5/q5Lycf3B7wd+d/JoLGlCW+HUUGRfQ57/8GVmqJ
BGq3ZbtXOaUWrT9yEl330xNKiBzRcR7wL/NByGBjkSpahKAMsiguEx0gsLM3XcHp
rPSF/Z6cFhMBNedU74OMwOdt8HHbvV3F29zrNShI3jbC0irvGb4zplf+0pR7Y0Xl
Dz7qe2JQQIEJIwti7e+PhgNfZZncTaN4qWQEB3RLIgy9HvWSEbyiNHe6y8l5pGwD
7aScEJJK5E3HnnpXFyIhcSrXbyYO7ss/eUYv2MlxaW4BzNTRq/tqiMUlyY/vnczs
h6K0b0NPIhchSiKTwIHaCA7QCiumIEpwJrjILYfCQbZmAB7oLf1DOIu/jPnA4+WM
jeXnU1sPTGUJie7A7BWIYF+iMky+D4GSmoBaUpkSEETPR+shg9XMI2cH+k81KDT7
KDitoJ8AL88i8432+WHL0f2IDK3rCIi2B5iPPBi3xJlqegeM6lPEaPlIr0fe6ME3
jUDTDgRBC7GdWqwX1eU2u6wVkokCL+2THMT/VJSnajnaU97OYm9tBeUj8aBHkQsx
zK4rfggknywP5ApB4rYlrchk9/FYuE4jnI4CTlWKam5HxiH4N8ScAt/gXhRoJWS/
OPjMaM2VhVwic+2AX9TClZ9xHteKRxRdtcRSogi8t10nQ6D7W99KGL31EpLP4aig
qqeTaHS3ewITJYHCHns6QwfnUH0u8sealBIrx8ORyTu+FsY2mPEyG2SR8C0ZFbFd
fi7TkmgO/Jf8dU4Dx3iDXFs0CjUNx5yrYLtBSSElWvEkolSWmfllS2IzNkDFjxsT
4B8miqDoKgQIXaILFzhVumoA6rzRM2HMn5sWmwV4wrFVEdJswLn/zuCiPzFBp8D3
6/lSOHcPXstVmXt5PyjNypX+L11ZeFlYX6GBaS1i2KjvtUdBWi0hY8coXJ5wxd+M
umXYO3KWekSnCn9KnmU5SWat/orq9fSqVJXnjx/rSAXiPopNqGQDP27uDgQgtigA
dOm8N3NMF9utsnvPJRob7DNqHQS8NKmWadIFKe6rtmw21MM9AP19l49SM3LVwEpU
UOWtQh8zZJY2Gu95aRw4CIXT60crQbIHzvvUGiy2MgZ1KvFb3BR/Q2Zd5hR3YUIg
jDgvTKhdeIYUlYrBLwpR9/zPWozbu3tfCod5dVzZ0/WSDWK0upDSFul2f2hlovkA
RwO4SDo2/psqvY4lRFbmYBDFudAovaMz4jiVMMoHjCyc+UCgP2JYpaEaK7WGHD6G
0kOiJAnS86FZYesP2DuMOr3GMVsw6rIhxFyhk02Lm0hInXhAfvLIDejjYpV/LNfB
xuTNZtNp9r0Sb4BBMOX8nge2Nnim9vwIcvEht25r196k3Hmnt877lGd6Y5SekO4I
el9Pud99v9nT26CYPhaCOStdQ6Rgk6smAyDlfgo7qqU2lEM5RACsIw7zkumgBlUn
xMISE1V0JmDktYDv+ZGZRpVOAF3+ZzSgyUWAIikFycZiR71FQy3Xy2N1kg1ZJfs1
q5axaEZL2NBcOSnbbTkntU/TWUBu3qCPhYcATKJsbjutn6eA/x3aAo6fG30Oc9J3
Ci4QJ0Iv+ukXR4+3Z6lo46BCMVNksHCZBZ1DKx8Vbloilq3Tq43Kv9nYI5JBYkR2
jacnZHUd8KxmUnaTG8yukRtH1mtsFUtN6FumR96qTdawwA2GHxVoQz+/lKZw3/iC
jgm7C0gvrLSKx0CR91hCDNn/f92U7U0qxMnmVZg5P5XNHzyKjtEw9zXjVLjjXaA+
ZOBmpVpqaCDk+G60i/zsFnV8GGJrBMBXTbHWik4tzRKBtTaAl4c0p5GtNXR9JEpQ
RtDGiF3vrLbONeSsMkyxX+pSFxF8fq1QMjF1LOVbh3s4khQgvtF9C+nk+Sk2SHH3
CHQaCFsikDmLCUV3sTbYMGwo8SZwJbFKEQvEh8MvGdCrrzLi4df/kNGwvEw2Vrgy
oZ4U6cb8e970ng2+Z4c4RvI7peh9qQPyrPDYDKMmg61sbwIh+6TQWFTPWhRcGt12
4RXcQW2zgD4auT1zvuxyQEGkoc7U5YKZb+LZbbkcgiYTMlOE53KDwvX/hcJQyo+s
IidATM4eRGWCVq/ZPe/TPWt05iRioqSjk/EdgbMH8wpSRdockfxxNavzdvoGiGRU
R0kaCrgpy6mdZkggXM+eQrGx1M1dkHBnYovXepjQl4ZceM/SHg7PZSxQc/7r3YMW
4KZKbqjEdj8i418GaCCpo88hiksW160OHGo6/67eHmpmkSRnCzLxzpyIyTCHf+8/
JLBnpbm2NPuuJwvw+4q+3HYioBqzg1M+dKUYSu0LLnLfPEKYnw6eWwEN9WbKL7+2
dZ9N8/NoUsHsIMt2XY8ZiWfQ5FBJ9HGI+H3j60CeSuhy0rB1WzQTDvzP3EoXZ3pO
unzy11IJK9FOCOZ7Xh0iP0FaBtJSe/StMvz0qK+QihU45q06imlZBPOND1mC9Hn1
J664qnfGAyZAuIOrcCzLxM4SBsMKi0VzEYr6MxOtm34Li/d4FrqOkGHE9YwG5URk
bq6w81JTkYpQFEeTaVeCCAg4dMNYA7r9mlskmx4CFEkm5WQNrLyWpNjgy30R3IL2
hkJjTSCCrZAdRigSkp4SsQrLMlqvhSmxip7sUbWZDF4i75oku7JfKOiZw1L2euSN
UBdngv9bnpmLonpVFgAf5DqakvnYiR+29cl1kB1t61pNRDc4oohfB3zuPo+ZSzgu
bufAjAf7fGO0BxHqzGDeflNK8oTv9uBAGmwqkTukhEHCeDYh9odHC6YAAm9MBm+1
IQDQHMCJBSi9npleA9RqjjJEdtV63QR03XaUnf1Z9pBIezbL++JpegI052DZgcLh
53CjYFmepCb0iN9C3M4gx+w/3psHxmzvaIHJNt9OjzkN6eYvPhXRTL8A8pQfGIWo
5F3oda2VIE6zsevP/1f5CjiajopJ3gk3rFZnaBmqhsiCZ/v4Xswl5KFjxjJgJjUg
DuPCh/ueAssmBlsnY+aMvzhtkDE88zavLNKmsItIuHSTzw6FOQF0sgAsuNJ11geN
dTa0JHJY4kJUKoyHrME9ECvrzyvFhD7+sYNH0C1a3nwbNmxT9kxrEOKE1rNsQ0QG
Ctmx09VGP0J7mkfIqFtc5Cys2AH6rWRnmBhprPaOTu1h1/e1oOkCdIJYLG5VTapw
vNUSvCaI6yq8CBzzxqVAP+LTzAQx72Rmcz8j67qh+Ilq8fTOts4Xr9AX+9TZxqka
LRmnMzxyIdBExLwKemqPgBUcToB/7ac81XST7qp0icsruxGNbJJz8ZFLbwIoP6Aa
JMTV4dp5Aym+62NCtUVG1upbB3sfVshBN1HwZhsoF5L5xh3U5PzTkprjJsgnIldd
Hq3KmiUScrR+m5XGbTPAz4zF0yO5w7m5wIK2mYIYAf3zk/dtzM+HV9ZRrrlqldBb
G5CtKYFdPcVLM8b3kn831Xnwb6pyLFYXzW29tcyNk8QRXIdsfAed1jpWKre0q9Iu
B57JQVZoCDlproEwnzCAjsgrtRugxtIG9ZcQqCX7Q3Q6+ZmWye12+nSzJ1duuA00
6athcOiGX994+AmIsWAjKLyrl8UMq2d4BkLk4n9tTaqNNqLCHionFOhZBVX98uwU
Hx2hPhRiFkDq0s5KwXIOoq8jY/1N+GmJBgXXUxpCw3+pR1dS1n0geYlyNnMxNw/q
A2cm/ZoSWR7m8Co6iohLcLPDRaUnPgt9AnBhI861en6r/vR+e4CosnmkPh0k2eFs
2KHguhbMxlbh1Hhqp6kxxW9zcQJA4uXO8tURvQag/7y9iMmGkDA5LRIWa8Pptro9
yVCV56gWwEBx+iPhvn5OokqR0I0A4nBUeNRTDwm5gzpX4qDSFM3IlHdTxDyPrqN/
w7UhTZPtL4xtNuTZ7qN6flmv/wsgAisvOI++06/WZPDYEPY49vRA9E7gkYGwU+c0
/bWYUgSkiBxVu0GDcVstJTNAM+gtB6JpIQcp7LmXWdOk8DcdagTtxxac3QK9WFVC
k4Oqqju7Uh3k+CWCga/Q0sNPIPgI45g5ztNMvlPw+likjnFjgeuesGziHyfCuLnV
LbfgvY+op9YQm3+BPknmr+BhUGU1F1mJqzvYBHqUNzv6tTnOc7Z22ENDQDBFnIip
wnbvrxL1nXhL4CDRbeIvQE1uq7CzrD9JCWcv1GsbYvDWUG0pXMqtcPiDX0uUezMn
INS79mp5RfN/Iba8h/0XBAgtgSuVGIjpS7zEHZQTC0RF96hAyssAf0IwNTQIHdNR
PTprOhkZ97JCkCyOh0mPkjhtN1j91+7rKJsEv37ryaOh2nxQt4Epw/hzQG00aMDz
cFA2EgwlGLkDbWG3h9lIkWgbHkzmIBLPStMgZFndKO1sMHszLSADliCgtMMvgUZ5
Qz5Yj2dBcacKmWmt7Mi1eMplDWELDBkUJL4rDoa7NyPKLJX4EXXUSW56H7coWAmY
zFVZD3qyFZSUaLcPp1VVtv/JVgqrpMeltst93tn1lLj6WeNtglxOe+4vjsxrEHA6
IUX9aW1MWD+rFLh8LYSlmvf9+y7MD6BcrB0zR8EP32M4jH0E5zxjH5Ucd8pGgKCG
udmYFBF/X51uJdvMRwQcuCcCkszNR/FR+N9A5arBhTQqSDdQ6WOp4XoK3gfk+ZbA
CJQzygL7LlDeXiXdN8f4Ed0kS+Bk4J0hNIeNHDypZGpANez7cyvs9rSUZf/J8jt9
gQcVs5vPQrvzrJHlHgoV3kXJnGkZI81r+kcKB4YZbOj460jDcjD/kCdRiHvJKLng
vTYNP0xQaPxhRAWBZPt/rE29ikvWeV2sr8kgwpu9UCOvIhFRFqAQFObckzi/s/Sv
JOgSuo2GIu6ST7iopELSzWqqboDlL7h50YRRqMbb9+WbrGC+9YshG/xRiFGXTBdl
tBNypGi4wicFXdusVp9Fg3mzMDwIRiGuAIpFwrrmeNaK5JEnW6VNrXZt+keBBU3o
G4omgy2xsXuY21hpF8e2Zq30d76Ury380HhNg0q19sge1/MKa/7OipkK41MPokXD
a3NLl/o89zm124M18Qwlqm0HVC/M31QEAC8lWNHOIc6vBgWiwPqsL0kcMZFdzMq5
1zrQTHiBTQHXwUtF7IZid5T1fmIrHx0uj7wNWQJ1MnvvtHWJGUjjSLiCn2eV/bSX
OgGjRe0pczCkVjxa6THRSDzrYm+yvaG5D44UHJYF9ebpjCYSg/W+IE+6dcsxnJ0j
MRFw50EIeeNCsfN6ZsbWCZy/DaAZT2GWHWBEmFyhDa7CxEW+jkjdkkRpMVr6k8LA
TwUar8JAOufZS6YOAATIyU5BpI/eUwtlVHZapCf075XSfNLQ3xEVoauuTuncgVrX
qOvl7xNv+u6SakQHk80Enk5wZOmH32ORtfDTC23HDsMbgi6uhrAgXE+OignSFB9z
Cmv+iRfegFuqCH8XF4oDk58p4XIwE0QB/5bwHz4S5jo48b1FGs5QdPRY0VXkXC9D
7WywFHex5PTnahBsyvXzWuyIRgYoew6zJMJYCQ1vnarDGZray2Nnik5T7ljTTML2
aL9l10b1onVTVVAMISZXJNwseE2/fSVzXKraQZUFJ9VhHzWXiuwDvaCcSzL7j87/
68gbsxJKgihUx9HLgS1N6n832RtWw0kdDmY38Jfb0yZ2fYbMx8ghFiOOaBBmDzC+
ZLpUqLx1uBy4QSTAT3LbHUJZr2LcUwp9Dscfs1JXfPD6xZlRQsEnBw6icIa8ZUir
4iE0fMrcncZr69Swq9o3eW9wPju9yxNhiBKF0S98r2tJA77en+p+XovqHhv7t863
Ugi9E7dT1aJ3PHb22xfE8WEv1s6qBZwAUeZEmKkjxYCSofpu4yBKO2GylEBuvkZT
lvqYgMs0iJOQQGQ+mGLFMfgvhEOoqsZzdgExFNRWlj09+HpMgCRTbwjkEOYg23a8
pU+BOTc7C/tkYFsabGoE3lJp1kwu+YMM9qDpCWRLZ+Mi0inkYuDBABQiyyFRxb54
vIHdQheDRJBlR8UwO7it8byJVA36pKpN+FbmwxZLtx/3C0trME/CRcus1SwKcTUj
Bfyc293s7y+1LNsbCBWvYB1QJpJMQWB0Jc5jDum51+z65Q43siBideFFXQXO1Odt
HPzIGndZf0/AIK33Izm99V230YntGVE9GnW0jaihzygrRZSkDlvWU8/yS6HdLclf
TMkFc0k2YJTp1e5mZC2lUkMOr0MRVQDIn3o9VtNsg4MHgm8nLLHnav957IKCF0f5
yA7zQfDM4MGHL0hW8j7rKj+x7rNiqo0wXtxhlmSHx0nUo7R5OyVvCdfEj09CC9/F
2HCUtdxfqRlTh8fdBPcFF0N/Xz36lmH5VR/XuLq1sL0flWMJi75b8D4SGlZYAv+3
bVYkaRD60j4lPnlB7pCSM03GuXu6+Jg5wH2QQIz6/U3D6iG65x9Nj2FcSjOza6aR
GPag+owPTu3st//BD0ldpgphv+WZydWWFb12/ZNcDfuLzrJibD21/bFwSuacChBE
Gwl9RFMSCiyC9IICSyyWUKp32hoyb/DoqG/A03O6cSRW1XatY/pDhg7jVBkEmXUy
v/0/+ANeU3LJd+f4mJ8DRS+8Nb3uI3u4FsC8lEby218sL+X1W9/zR69aqHcqbIyl
sP55BksPCrnn/MYmx99kYXQTN4yzDSOHSg8dDS3pwtRlFSe2QYGZY6nq7a4X9BVV
rkoYTDdyLyIWsZJmZo7LfV9d0Qa5ngJQdKzPL8dvHjwDtQqD7W7Sle/78lWo7mvM
/TmgDwIm5f1ONPuWDFDCkNzeXx+XMEkpgUs56+D+EfheyQ+a0pUIJvHroRSKuzp+
bUPIdWtJDp9Oo8vi0Renq1/rA67L5M9wkIr/W/GVQhjLXkdEx3iFvaqOEINmdobD
VgiXbzMLbTyhQAiAuF1xte8BHllQ2TbH0gTgbjMZSiGqrzLnSsAD2Kis/q6Z9fZ1
VkAX/j96yMAA2o+wlsuYsh/A/hZ3XbGcLsEa7SlrqyHgmWlfrC/4nIsJS1AoAhda
93krG/2LsNHjBPnhWZnpjl+AuEoH5trNWqE4qoLacRkL9bBKENNJLz6+Oa46g/cI
HBDnIMfkT9JhUZIA6WvKB3eeyv6RctYjZBQ34lC3tAYsLmY+5SXggCqK3IO7R5lo
4O6GpUPQ6bVY9092DAWN7d1EyR/o+rqw4XuMXEceT0Y67g1fcu0gevXKfAgxolOB
4Ok2UhmkZBFGg5IAzuTkG56ZSNgVDgQ4bQt6SFIYMW+RHahCvmHmD2O0NG7NxfFw
CXyAdkYi12ZIOH1HyYqU6FJtDg74hDsPaNipM6vsGtrMj0+bDbhHW3RmUDu+wo2C
tKkTA2bUMnzwgNoGH0IYCFO9g3xWjFnMFcaDg+iKwoRiuWb64VdduH98Zaoe8pxt
Sjcn7a2AZaLulwymOf9b3lpcMPguzCYlzGCZaV2VFUbCJrOQco++tLepC5fKyrP5
DYd/XwHQL6dvd3XTIchBHyP574Dw4Rvnl7ME/qQcksRZgESS4Y4XcjlPPWGyyt6l
5IKCDiQQm9Vu3ZrJcSjwgeQL7ekazX2FIRG+W0FSVaMF1VrOnF5rfooJZWrL0QUb
okCOSZu9v5mFpfDAAsz/DuvR6q4VNNL/SWrNYZ29Uspjwju215eBKG1K6HlvPl+/
XlciNfvW0/FSeBVMJTu9q7KO3E8VTHS4ASrWB7c1FAiM1bM2OpjPKOMmQkW/VjAl
BpypdaibeFWS1ZX/Znt09N8mJdHcqm3qkQ+d/ZaDnat8nx/JezgznUw9rLvFyzG8
Laqsuv6rK4Ei/fjxaR6T+qA+AOXAYfpo2UMIZHCX2uo/kbymnSLKdLwt/Wp6iXmu
S9GupAzD7mQCP7abvO2ifYCB3WA0I87iqtFzf+oii0itShyziMkzl0sE6nWQ8rjo
4yOcCbl7vc7DOF84YFhWOh45EDrGh2nULAnVX1nzX77m8QVl1yJ66jYZS7SY5L+R
J/ymiu6RuBkHP0fg9WHj7blExr3XzlhzAcL+Weg/GcflKYrFZPuq9P+TS7VvqEFd
nEwCR55/c1M87Kp1flE9jOAtn53EFsM9DoxKDc8kjSN0R+7VrfKk8EnKI/2tv7vS
TuATv8PAw+gqilOrpt8glCkcQ0Iban9K30KhKpCg5M5wJXyezCyjb3NTfig209/N
5368ymw86o8+IMpQnDhgMB4iuNMBfT6eR+RdJ9xmYeRYWPNUrYy8FIOt9fYJw+Nf
QOM68ZRO5QYtOCo27K3EGhAE+YLmVkeeSg+BJeporBOfjQ1n9zhEWhKYTTLRUs0x
xSexzePeqH/ZHKcYnNtk1PD1upixXuGg+gpRtOe6buUqF/m/5Rsu64+H+X+9Lhrq
5nPEqsb/ca42Sd8KYBpkijWRbqv4jOG5jjKaFcjgU8/RUVnBpGMHkBBwyAYHUYFN
Aj5ke+2/YbmHeOluRxFLEwH7z6pynMYV/00rrzKlF6GInqUwdq6KBBrEeJ/tAKa0
iRH3kr3McGD3G80eO8BiCDvpqrvV1eg4H5WHOXuvQGo44hje57XKfdnoGd+O7taP
XjQwnWIGXp24ArOvp4TGnj2X387WraAYWRfvUkD++17FVxV3o1oRb9H0xO8xWFU/
bDQn180PjqWmjQlp/B23BGh1kzl+QvcCCgY49uSvTTD1j50Y7J59JoMUmKb57ZT6
3GrCuVRi3kGQulkJZkwU8VcqUBDJEGuGfADXElypyLQ7ZXyms+VBU7+L8ZgaCttu
dxGwR+S89snNUjpW9DoOdNckv+w8ke9NI8U/5Qja/58Oze6T9QorevqkquxMsqD+
as0vkSZJTVvJHvkpGDg7ylH2PbMT9jgJ5+Y57Gq6d03ggCW1VyZUEPYjYKaz2Si4
9Q5gb9qjz5/SOYFnXAZSAWgbSRquH64aJtKWOMg11q32/RHbxBALs2a+yK0Q84CY
nRQB9HiXrzy6gXVJYKi/XkbcseUjjT0IfifcmuXqGk3fLJzp/iLqyvgw4LAj2hm4
z5jd7yjQeqiXGemAoC2ZpVcONYAicQd4Pi+UfM4gaRaEJ9tgx3ON2AuDBPE5nMgG
9Ogn1MARK1KzzEzu+DTwCIs9I6AjU2E7g7Q8V8fr/8xu2TU84qU0RnmSINHaw6nd
sktGv3YB+u273/44F27AIR8WaiBH54d51PRUbgVCwuqor3q6MaNybk32tQYC5HSj
6mi1GqLB+wtH/Qww4UzwlWWnm1pQ80fXmSpS7NECw6PGmQH0tIWXCA0t1CXekkR3
OIManpaPDFN9wuoOY2XBdGM/eVCHLWE1h28oPyU6qFvs9ABqZq15XzfTVIPl29XV
7ID9qMBgySeXxlVPGxKynSvtDYKg+B6Es8KkktIcPRKw2wsPWodBP3Ndth80KwKQ
EC4YWvp7YBcO/gNdZUMBVL6ExgjcmDF9dv0Dp94lK26Odjw25IgcZIoSA3Y6U5pG
r50jbc9LcCr43yvrcOPLe2fRwFw4TdETsEHuIMO99f1T4VwkZndlFR8vukVDUbfT
B2nuswjgmlZ0Nz/M9+hCtRp2Tiyj4udui5RwZe2HWGbR9jS06CDb05n/Cv29SIID
ccSdQqnefqS/4+T1rvkkrXsD3kMmUEQrZ9Nvg29uEIgRsxgvk/JIMvBlujz5IoTZ
auLdcJUyIR6DB3a1botIX4KbwtO+6JRcsHSnWVfkDCWDvV90uMYEEAx25W8OW1F3
JssBeH/gw6VseNXO8nlzwVxH1vquv9vWxSb9TFeCDB0DEXLACt+4Yme1/PELlhbt
Ml7lJ62OZJDQHa3rlm639waI6UUQA15FvP72GcfrEPxLPWumqv5iLoJRNPMPfzhx
Jod8q1994J0Rf/ZLK4QxEgyHtZl+9RPYN8uvHCqknZ3rnxgKhEQ4SCnG336Z+ux/
XqcJ3UgXA/3/V82JZoD8jAN77rLb2nLnmGYOcLp7+BGqM38s3E0Qwq6H5AmEWrLq
sYJ8RDyCZ1H/QCydgQjCXPogz5JlwnA0+5xOEum+s7/scfSUWdi1sWZfZhlVU32J
OLNJcPqkCgGV1+5cxPbTvUjISIFOwgB71WfErrU3XM/u9ZNo+MVTIoVPTGZiUiCU
gMdEB1Fgq+0qLK76O3pkOXIGW21GSKkQ9bAj9TFoWkid4hec96F43nzmDa6t3cW3
grvd69fMF+u1zs+yKY2N+JyGAn7FAY68hakY02n0vYwEbJcxO7kbpxNAHVtXyaTh
+ZaaelTqS7OO0OSG8w5Lsi4T0AD1GY34kQdHxrI0mZ05wpFTITiGMZyWP2hrfFfI
MxxXlOKHZp1MKOE7FTU5VqjQRBYbEtGZenwhguKfizmlm/RWrkGGkj34WQRunOeU
5xaX4tfaqqQSqG4Xt8DIXv/UwUYTqvW+bTZz/SlAYr7nt9zJrnr7ocQZwPTIYTjd
0pht6o83/AXxFx+9S7HdW/LyBm/1ImjhhDs38CKl4caRHulJGnZ1jahipIuDFmZm
p2LuKGLjTghTIrHPZXgEEHVd/PHl6cp1Mdi5FUX4mxN8KA8uuPj8Q9+QG3ElNU/J
1EpTttgDTMt3uEUqEvnhTax6rDwS33otdCBkfU+G8iCqEgBsFheMbdAYhFdhieth
eLpcQ8GLv2HtVwqunfMQJwKfZ1zDzZJlQ9Q8ZC7IuWehYLAXo4XflIumWV26wQSE
VGvlsJ1ow9samDpAqPTiaV33euiLbJP0elEzDUAREv+sC210m9o7JuOnGwxsG3fY
PDHCy0bYwpU5O6s1cjSqRT/4wBVH2I/1R5ACGewjkCNaqzKsuUjME/06XHucl5ru
+ZwQBkwK7i9lPLDyZf+HOWRFPfr/UxsuvhCBI+6P9UGQ4l9fA9oyowpcKYxKkh/b
mO4qrrOZcQ/bOcHwryqWs/k7Yo4ymycRVco6F61LXWL/Rw+DuAfTKjVjAs5gw/vM
JpAnmn1eS0i/k+xZ6d4GwFpmvMQJvZgzxq/U8uE1x22zQRwJ/67V3WNTT35csKIE
FoGG3ilnF2pjbEWFnOoJMp4Msvb8zMgtFx+l+BdBBAEprq7JdR4ZVq+wdZiNEKZu
1zqMmfDO7tUAUa+mbkbtOAQHCYrN8C3RdAt2UN9zFjTKVVZ86S6TfJSERLQDPcNK
eqQpaDm7sOnOR23YHYKdm8gOR5V3P4mEq14Yk9G+HaxSjANBPED74GiW0N3kdXLt
rIy1Ri+U5e58Chqygq4Of/W6/cRyGb/SUF7L0bcbNJjN4XTVJejqMsEwGr3gsIqc
Cc2LRtpW18P0xhtwbUc87xhcsj+LPN+lMGbkDG9d8ugKRPrRt5gbR9IRP4LbJPll
5O7FyPPdHABer7fYf7WTLWIZu+V7iWjwEfabLPf6LPFBaEvv4wXHxhRx7mZv6TMG
8ZXJi/0gRc+q9GjahjWULFDB8eS3kODcF9b2PDn557Q5vFXe/lV6n6jcEu0600VO
XLsdfWyYhR/In7kBv5rCqarbOxvZVfhk2zYPqItI4TRNraRDOESTJVGK/FDp7IWk
2PKCaE7idN1Ms2FU+IxXipNcvIJbYBIe1D5cmy2HNQnZyfb09Gz/Yibm2kgdLqre
VcD/Gt6puBtjUrT18pM1WKyRiiJt9M/6fTg3aseCqQkewxcVDlb+8IuZBcDmZhYB
IVtv97LPr3UJWxHrk/GvzmUjrnRA38YCllRVYwZqpg7mhEQk2HeKwQ9dwKwz4ipb
31p3e1C8MlcLjy9yrJgJ3RaeMreqKy0qJqFVZLj2Q7diTjdTBxH63yBc2xhYBtOO
0vxFuqEw1jip02HAV7ecjXnus8AxOp9bkP149yjUV1QBaxTUrQZjNFrcgWLuA9Yo
Ma0WFzb8bT3UzSnDA7w6HW9cNxiFkg+xX11lmVxupZgBD7DmMcda1GYgFdYbUu39
nHVs8ZIsAEzoILjsP0uFEB+4PXydfDvl3SstyeKV/GHYu8dcGVPYCUQM0l+M6zQa
nD1itx1H4vrWxUycN01vYhcp6q7w4CALX9RSa28Dm2ulHcUAUET9OjnXh0uKLUj8
BBcML0rWfb5B5WhpMRNP8KbSyLkQSyiIAANW4A06LarKBVgwTxO6jb+k9HBat1On
Me3YEAvbko20SqHtDuB0wlNt3xVmSOpmrY/X2CvEMyumwmZ0muU8MmyUetrlPWMd
aT8tzubYN645xfOW+FvT/K/YsKBxEO6wqGNQYb5VE/gv9fdTa4Quhf00ViUHrXEE
URD23mC/M/wulRLSnPernG4FU9r2uaI6P1ZMF4tPqb+Ht2EWC9PV8QADk+DoTk9o
CGiX0X4GleOLru2GUNM7QBunWYYY2oCea6rEDcSQqp7yZQDhTpRRTng5kGuwXBgb
chT6IxQXPYGGh9hEuEwjrcHhERBBAl9L+2g8xRqSO9NPdfrzSBZnxS5o3/dlSvyq
J+hmdOBiPqO4ksGcI/nRci4HBTQAGnJtC4RtzkSy+D9hqtxRBDohc9gzAtCcnu+S
LThNTBGBrynUaeX5hOcvO1pkzTFQfUD9JSbRPrlGYAs0Kf8kbrnDRJ0SIgk/ghm1
q2wbIKMYhsqBdgw4fDnpPdLpMIP/x1gzYFVzO0eCCjTjB97LTwDooEKVTFo0weV7
C4ojIsCo4VLyHqOJ/RagXp1PjQNDXZ/EcJhhFWq1gj0rN7Q3DreAixsZ6e+9HEuG
IDwHeYerWA1CIewuvPB+7raBFu25LTQFsar924kOOCxUEolx4SiFK/kAUVI69VHo
C6PjJY7KrG2azR+IcI+wNqrTAyi75ATumnHMLmdASdJY4U81oA5xSuX3NGFs4AsS
JS6SqUHRcIuEXAqsJvWea7VcZf0GHW0OtjAxdJsb3dA2hXr37sK4EFs5MYFXZvu9
ZaDEVufaSCYL5Zm4WaXufwiu3TWqHdrQPhYLks2C0rTXXt31XhtM28fTKkD2rU1T
lQDg2cA9AOjIZuOeufYIzEBqMktIMX62di0tgVBwiTHZkDaQfoyxTLJJnAIG+Svx
4ZaiBCV1tgUlTK/iljwWYcOg8k1BBEnDGsG0e7oBqsd7d8ugPYoQM5RP9FPeZckp
xCGXrWWDTHKRzQhqTVVK+YbzdZfO/YNg1naRntCTrmToqM1htQt7eoj+6RHbJiCI
wr5BRUMrRGyv/fZC7wZmdPq1PpZzBOHLYX1tUwNWtqRgetgXR8JSmhTEgVnU2ePU
nF6xy33pk5yO2dWAdpNgYm1wf6EnHLUp3V83CswXTFb/ycc7o0pkPhiEajYpRycC
53LzQ7SnAGn60TE9nD3hmrdmhxdzkzqkIRtGpo+f9TuiK9brARDwe2gJklhwJxDg
O2/argXhwxGeC1Jg/wvE5ujlpLfBOhJZPaLKfCCKUi8CteoPykSQVMD7EKAx3WV9
0Ck7MxhR4QNtCv9QHxKoA0TagKOpGjRt/hlAvX1gGuLgic3I/p3aZDaqEgicXxmr
9peKWslsJlDOBaRovIaJGjUkxQ8QCTxZM98dhG3Nc5k2kDdVzdNBfcgaX7sS9gor
dWtpvCXuj7s5dhwgCNWr6gUYeimNml/IcLrO2zsOw45S8UzC5buQgzOwGVi+ZZy4
HsoHm1+B2m7VmpXRNjk/t7w12xWbYtZc7PX8jobqH7wxwBE9IXHrx0TtodxdE0x8
y0opGnH9yDdKd6hgCQBBNbM3AHlBfyTp+2XduYK4o9ZgBwGuvViB0qVB0yLf5kRF
wwDFOwYi5SsdCEoBjNi4CprYSBYrBfx2QEwSJ4sV7PthRZH0O9XDz2kRbsL07D0A
tGTpldnts2ScaMBRvS3u6J+w/P0X8F3MBE2Ur7M12QulWaOfjyLzpLS33VUNZVa0
Md/HgaMdD06e//YAUT2wZbTiswhosjRhiEnCd3E32/Yrn3qzN8yOpdFMmeOf+G5H
nomqvLzECkIbzIWDaBE9jFc0hjazs+qCkbB5Ugc4A/QZ9F3a0QmX2Aw3mHM5T8RB
W2NfDFGw3ZpL839jYg4Tfj7Aigeeqrn8UVBfujkM5AHS7gdfVlF0Ey8XXUixEvMj
Yv3tZSUa6hi18MFpF+9MBJTiqqyfJYYVp8NVw7y6d445ENcrJh76y/UY4nZOcW0/
Bx/gv+qenKMvS1qIWGWcNO22FECPtyoh3WLFgdwRmxET/au9ketYtk4pjY8/+lk2
z2ctHvbTK9PifaTYSiF5OxssS5SFGKtQEWniZ1fQIsFoLBeVOJ7TCoYNBCpulibP
DEu65NS99tF4bVOPFptQmDSD4C0H8PnNB2Eg9Khyse/PQsKnLq5dDl3JXElU5IaE
WmXHUWgFAmSDPXNKxSB+B7yYcGXVOeQdkH5g8doys1DfbhH6b9kiXn6rzyD8OsNV
CteUD7PfN18YiNSmC83xegzg8IQuzmOGs5w7gF4Mf0uL9hISBs+MZBhIcdaT/WLO
xEAP/fM25+Nk+u07ybIyl9iIP8eTUC9HW7iyfFaNGe/q+/DEM3TMlVdL71cRxl7Z
KhmdOjxegVDQMtFe7lP6XsoC8l8fBhHIY4UpY3RVgRwEelrSRoDyel1Fg38/3Uy9
yUWYJkjVy023ku2FpLIYmpbzWWmbwqqRFJ0rAhQkDq/BTrW/Z9Ivu6LA+/pxBEZj
+yGnqOFrB0pbFbtnjaFOV6iaeGbmec0+v+jKdYEJ9xGmjSmX4On+QRm39OltloPR
Vb5xpnCCeYvjCXaSfw2QgTKSNfq+ZTZ7RZbYu2z+Dfsz1JsyOb5s60DPafZLXUVP
3pvG+AIdh2QlsbRSqqN/rdIOOlSPtBWcTqDp2Mot/X5fVNDRtQYSYL+DQfyxuKtr
0TyzoZtglZHJ3eVl4ZFc2mMx8P8MYC+oBsjcGLlB5xmQ2NyIgkEQ83LrwaDQ0vEL
ws9Lhulnku7RZaJem9Y2j1Ogllo72bgkrGj5bgOgfeq+9lIbpYkFn1qzh5xz6FkN
GoGC4a50mhg5n+w5HZjz8FrHOPzTa8kU8ufhqItyFK9w25D+cNROhcUXSUNp66st
qnBts7v3fDWAkzZJfCoWsvtngrvQU2veI21HcUMYjKCLuBkQo4q8pIIuZIH0DHOy
I+KCNwzeZFxfFBiXh5keo1BYJsL2i6taYGwdYFPs1q5eRBdQJE0zQoWoOc+4LFno
Xfakz05y7v+19SjUodnWmXDGg7GNDvABQpNnz63eCVLzw/bLRiSbU0w+Kv0JCIgV
dAWzs3LodzZhG26F+VyLf6jXN/G85KGddTXvKvLahhmQ3Td2krGE6B6JwivBa9U8
oU17euCinF0M7UakJHRYz4CIKsmZSEXa/9BrZGVDi/HN8aKimNwqdBYBNquYmoyL
HAEsGE3PuowURaAGiwzDS5wkztOI25sd56Qh5db9zr2HhM6r6Q/aKrW3dqmfB0X5
NsS2Ypd0WmZsx6478ZliVaAJACwchHgVvnwTgTX0CbIeo5zuOv8JfPYuCQTiRHB8
ipL8kI2lM+/kqf68oBq40vCTXgDU1X//DjXKCzj/SH3rGNYI18gUFT+avuF+7Vn8
5sb7/8WrZ8IeilbCKFtnKNdy6vuOVAc5slmC6KogJu9Xz8m/PZxITsgYk/fZmvXV
qqLCmoNL04V2VbVJt9bxt173/0PtwXPq7USpBpmG1K0YgLqr1lsLuaBzcWjghEHE
+ApKM9r+0lRQ+dWzZX1HyodaEh0LMOOdmMkXlKA2nKkrfvLHSlWV4by3MQxLzMm7
UH2ethMVcrTX1xtEK/IslMGA5KR+Grquk+FP1+uLmmHrbNNuACRdo71XsKBRKMKI
AIVKbwVkrnBXtTMdRD/3CPFihNafo8W5/ULk03ZsS5wkdeN4kXmPEErYXvD6k8OE
tKCjESPapWVUkxVzBRMPNRCngTlCg7URmwAqq2XO8OyuHPT5Z4vlLoXFX/Ob9C/O
xs2pBtWpCSPbDDzIhpVCcPsk2Nh5yxNFv4KEf6N1y504Z3jCxFsi0c60cXCq3wUO
4A8UgIdZIMhRggxiB2FlpdctKtapFlQlDqRx70IuKa/Hfbs4r6MSnmut25TFQ3dE
vgdLH0A4TDuBCbZzdCRHAQ0ZqPmkTAQ3DbZWzS2BhO0f4xEa+UIWZnIqFmbE8KiQ
Ihx3JvJpHt4s+tncC+w3mKwFREqj0tRTpIxw3TMTNDkl/LqMzyCruKCJ21EE6hEO
bPdWOxsKxGR6hVwXqcvlFU7POFi2Q9Yh997EuiLVMA5cZvi+iXrxJlcvU2gAeA0I
6nb+F9d4ZH/q/NoVnpfKxZb/b/lLEHuguCb3g1unondYhfG2DHlRWJiLFANj31av
EtR5sXCzOjcwUQ9HHOoYK6RbLrCOlJeSuqqtgwPGq7k7rL0R76Cw9sjSz+hFKd7u
scP7Njj4IAiPF9FsQk9KPDQje1YYQtSs5xiSiduk1qMKEBl1CyF3b89XJzh3Re+9
0vc44hrUCqQ9nBJIjjD9scfNXHhRq900EQpkI8mYRVBRpuHbZf74ehxkf03sCJla
WTWIwAmFqKI/IwC0fugW7EkCfkKeK4XmdKpz9YS5jZ/zY/PK+H45nAL/9ohl6ZRp
HIOODTXXZL6DLOygjWHuUlFYdjJ97jdJxBSFhrDBHFcZytE61VY5VYWEwhVClEr2
MRokaYJ8LBs3dpGvWd6e1Dnto2Ab+gNEbZ5gPj9hW5ckFNJrglqFBUILekNXom2i
DqwMIjPjgdujcDnLt+xdqVJ0oOzK4EcM0PAKWVoaDp3xiBd9p0pexW5srzuMuNFl
JpwpQwDA3TtITTEaqKVC/inSopxYx4oqJ0L7sqqIjL3uiwppGaUX/aOZqweBteCY
nm67IplcBHOuHH3zvdntq1tDoHX2X2VnDfD7h58AuCdDuqVS5gqcd8vHTUuHciu2
OpbQPVWbufcEysCDmzyrwiemAPaoxr+atnY1xqr9A0XmH+GwfKxVXHqDuz4EdeVK
EQzOtkJkdbyq5o1/cKy2WHaWcwZ/Zw0PjNh9cFfru1cCMhs80iWqMVr70uUMK6+t
7RXTW1Kp1otwhjBYc8a0Mf7uzM/ypkSlnvfxX2KM4TkXWm4tH0q6THid0YkJ0ut7
L4LVQYKEezTfo96q8O+fJQxT46P9RZbL8UDT0WSdvmswT/ZokTvzXI6yVrpBLvxj
xlpZIymn1oUTWIhUeagwwE1FPqpCI+zOTlL74Vv2lRRinwpHpiuUfHEba9BdKf91
SxxubbjadxjmWjCLedPVRKWyMnj/3AhAkdOmwyNBd3fgX6GjmSlImcWupR8RAC7O
wnAD9sCAN1EOKRuB3fcYRAolNjsDGpscfBV4qiBsieCLzzCWntGQ/2qndSYqWSSm
ceTYCDSbPqkiYfQS7oMssJFF6xmxW7imPU2eNrKUWiD4vvFC9Si/iAL/0KriEoNF
blwXReQ29WKgwC5NHReM5zi9E+CUljq5oLvfpp+3tdgrrNRFw2YVy3YcwRroEoEF
ilLf4nwpfeYrRKs06CNAG/bKsmHkTg07VXY9DdpH3UIY1l8R+BYQOhS+dQkJhtZ3
0/pAjuJfF2oN8+iMgTAbbd7R79/hD0VRxeqUKHO/JDRli165zn8/45xq2xmaVOHS
zct6wvBodkUMGUFVjszyAVaH4urechP3SajQN9ebaNNTebrXwZbsu87FJOUWZX1i
a474mJqLHPB5FZW6mMdO88/v0Rb4gZOfwh73nXe+0/NWxy4cHc1RxCT7Ta3B9OtL
v8ntYBXcfI/pOOYpG3WXkbO0lJZG3iDahCS/e4wmv6B5MOihYbAuCQNYwi+NNwX9
dbLGFuNlPpIOG6DZXt1ahjSiJE9JKBUdr2Kc4VrKzUubXESxE5kNFV/hME5Y4czo
C9VrR1QtS3ATLXaCbfIJveWgPYi3sqWyMrGBsvq04G1HO4qUXa3Sxt16TrN+UwK4
efjkuprFze8Rev/rC75+V5ctDaYnfNIXraTLDOQl5rK614mSzXLyIry23kwnuaqC
yz012Z1j2+C5bgOivaEYjhSqGVWR8k+8st7SqzLP1wssRcQgBdWkEsQwwuMMKcGH
+eBJXGvR5W8JS9HW9a58euRy1O4PiOo7djGJJHWq/fk13J6ay2vtutVJIY1WtDfE
9CNs2K1DLrsNIRFvAiEDboeH7IDrXskySO8v7bRWC5Vi6Pe+Ft+IELITPkoLZb5w
4BYWreB08k/SSF+9FdU9HJf2tFqWdSJhy7rHbo6eiXoxMDATj58HPYCyij2imdlL
1+VvODjVuajBNrX6xOEyhxXV8x5ZvIMRzIco7RdEsAr+4T2n6DpBSqGkXvzVIuFV
utx1byLqzquIlnsvFTypfNIl4DHjeR2IuZJKqvCNcYmDPwXYwIwq/ZiiHNqT/lj+
ptHV86FQJgwutdVVNADFwuTd4IX+KaOvUrRZiLbAxFiq0Ff40CpTzcmv/Jy173AQ
uRw5n52f8mFvxNKG/koqGZ9LeI0kfPhbgUXkyAH8AWmMbO+z+tD2ke1fUVzF8TnY
dBKGIZRLpBawkb+GrDIk8R8ESCpmz+vPyjjKiVOtsA42coO2OIJGzKplCp4Rwtj2
QpB5bN8/3k8tVOBJ6wbXJtsfz1A+9NtHug6u1cO15oPw0CgPQS+qaLxaJw/48ufg
3MgDWOEY0vGQl84xEc8r7kwDjpaBkrUl3D0BjRax5fgYOA5updBwhv4URdNt96ue
ycZNWPnwtvpaiG6hAUqXpT4gFApL4w2CbSjBX4RsOAUAueNNfbgj/RMnfvsSIYpA
V5UGyVVaX8EtQhRNq9Xlrw9ZXnmbD+Ew4tRQn3KiX5bNuPG/5F5cJ0hMabatORH4
eD2avzbSFtUPyu+7rrTRfiQv2jYuwYeEdeIwVVdT9KsqBYzql8MsUcXz5AmsEoEL
2U1y/rx5rF8MZzKR9Tcdhn+pGeNsGuy5wCzJREgHKZV3KIUCnP2i9iAvCUj7L6PP
X45oD6z63zexJOrn5tIX3ckAD5u6LAzni6wZnFoUwrgC16UeD3NsttqNaGglQeVy
CUEYmlZjPtHvc2Z0YsvfEZbEvzyrnvRQzL5qlurF957lRL4X0QBFZqbGR9FLFqpk
xNubtb0nH0crS6+4gdYThhSBoiB5RCV4gsB0pn8MiPcsldoWCUkaGU2A/FGta05O
ybBNtWdAMq3NDjQzx2xukf8u4Zo86S/wUpCmIEXmLOH6evS38BLXcpNQSR9vPj+R
NfSUoiHqIthlvtSu+e6tjvmcHiwOhogNEu5qGjpQn3h27BDjmHDEs6R9BNd+AMdK
NwSVh/sFWqSThrn6jdTBhf0nchJc9ChJ0ZcKWGBbm60CmB+kgoNj7iC847IlySiK
Rb5RO/KVTWbXt2ejez1rars6vCXdubdEYQEsm1fW984iW1MrPgAiUGxzY1P9HI3q
Q3+jwQRiaSPNcd18JTlgj0pWZRcM9MhKEBP+NQqlvbmPLWATQqP0R0zgW8sjLDjH
TEuQIF1YKnlsRfK47B/7gjogP7u7ZDCUqeSbqKd6HqSpLG+vZCyDBm+AdJh7/ynw
Kbl5eQrUQt3IbkUgZnAxbPiAot6iKJ+NGgPcbdU8xCPbPFtyO1DpGMA20xc/GBTT
/1f1FTH4gPnW+4cGh1HH6FlmgjuwRVoHucziwfpf2MVH7ZXlIRUea7sTokUyKePJ
LHPReI0/qnVM/3kt1fJpCumqhVCcpqtnJPrAc4KcsZ/ePeVdWKHOEKDcczE0T1X1
TrFC9QNlMnQrmGMK0jVNQkKsCHZ6SNhiHT3+UaZrv9tCmx/V8cw0dr2w4tjjBP5c
4QRLhTLOo0A8d0j86ZrlR2EYKOAhqCLC7GrwDpKhKMSsIV/81IMR1jyQBN1Ez7lz
113NjJy2+6LKdGOFVqfFGI6JgTBDCucWxWHkRqyMQ0/d2ABvioN5D/QNYgFBnJXA
yI5G8WGB+tnC2n1cT/5GLUyFgcEJMtP//lIzZGoCr1VG5HwVFXFivIVDc8qzX0Ge
vVyYZTk2NbrxD5URrxKYLon6KemKmkjP4bvWud7BZ8yxsq8wOwj19bmxeA9u7XyJ
lHQ3cnTBSM6N8IvR3F8B5184axkv3JpG8RT10VqABffCUV9QB9tukV0yG+zYw9AT
RhImpWiRkNHINClFf0/YbjXEd+rsMJDryrmOUfi8453m+HShKkhvNtKZSPixzIRq
Ut7ALPZkCDv987mT28W5ttJyel2MUdHZ9TAC4WxZE+tsmL1dQwN/MGOQWW3qLh9Z
Q10E4hk+asp9jO0sByBW2ZGAev/mdpY18yA5T12vynSG7INh6MQAQHZCMgvmlF37
lT/KRSjRqPvi2gSlrFhqJgU5YwOelFPpPlCBttPIouzK4MW9fwHsEIFcRdhRJxOy
sg4o0XYfRVh/QHkIXC5oDOL2zRKXE0RJAdorfC/ujRtqP8PSvBnVBlx2FN8jN0mD
V7s5vow7MC+ohJ8psLHlt+MWdRK5EGRE3d4M8Hz82KRqGwPLQheLKRrSIz2S+wcu
a+RaFtb7xzV3Vs7pk/ddZxNqU9urpKDrDEApIk1jebEDzDIYw9j/hxebU8MUE3eQ
ACCjYht6Wp15Rg+q8wlRoZVAFzU6aQh1o/MfrcxNiKa8RrUzNds6eM1aBFXLCG4w
kFwj5P/9iJuzcSwzPAbrdWOvGUIfREZ8Rb/11dn+LMVRoxmwNbwDl/DS7Ea95XNV
frSXEIVtd1isWLAkTFos45CYkvJAqhl5+rfjFJC/1G/sL3PFYJ1QwLleSS1NHNLd
nhNgFAI8TEPgBTTTpU/A12f4+ZwfMY1/ZnvGh0P6aW/NJv3xfuRBTRbc3yL6J0pu
wwpvfZv9GwKKDOFTvFO0h1NCBokR8lDfSUwlo1B6wn1jjmZvepFNssDeYbcCzors
xWvJ26cZrZSOyGr0n8XUPrP4d6n9dTt0wwRU6oym0/KHXN/neEwczhRxSqXgj1sX
YtENL6ydvc46/AztSvSvU7+BV3DzsP+gLTS0LwoP67Hn9CNO7i7CTRTYS+EbtvsF
lSg0B1cYgQ/RHwquiotpeyL6Ixs/fb3N1jZ9F15RjCiR+rS9jnE3Yvu5wCCSDWdZ
lLemw7fx+dl5IkjcWuGe2lyr22TCIM/dc98bjZV/gCVrIAweeXFpBaZvEhuaSAd2
hkll8AIB39mpeqbe14z6QzmJ/yQVq3IBKBvDAEcHqoyiozx7SU1ZxryK7XSjyt55
zBNhmo3zWwS7X164O8iBXBxrQb+7tIrb0W13OJvRMp8r+xYu0+rIthkyDBHXjhNp
hWgpmzRxj+X+JBe/yC85l5yYUvGDT30Bg5cIFwUBKy7/kc2IuRhz5vf5d1h3l4wT
QQk22RpGPrvfzcu6T9EEIyTk9yqXmdmz3fdjXqhI/Qdig1lTzu6NvjYc2DyKrPUA
uQLEKNX0osZygzc5g3nOkov0Ax7DEE3LwaTpyoRQWfEXKl4AeHrYe7obmewfy8tb
cOTIg5nEhdc6Chy/LbSvTBkMxsY9FIPwH3WWdNfjsmpUNcP9fUcHxjquD6KES+sG
7Jut1ub77SS0mMq5RTXawvfsvu2L1lBbo85UztIX9HH6ozQ9BbOUlvxHrTra26A6
dn9mhl2tV5CUl8jLJHnyVUa2eJsX7yiGS6ETKBlEC3PNVTRR+cae2c8j6pSSV2Fw
1id2xb+SVn0ez+tXBTQSnp3Gu96TFJma8Ex3jS35Tg+I18nn3qdVOu2UnMmQ26YZ
WeMBIPO4ejef+Z1qw8DMM+SZ0YUXxUCuyWOOMfqjrbkm91rKPRdyldukjriRBUI2
OQ2o9676am9rL0m8RFzBY1eigJuZceNgjjHF2VwFQYh5Sb9abZknqR1epGDCo0Wk
jFS78w8Akd/VUI3o2tjEmVPUKUAyB7VF4mL/w90/N5pUQJk3xm0YUjNtx8zL2Bta
YKKIyjY2/CqGVvT+a89dmZ/MUss2lxiwIb5hN+mZYzNzBfkRxzs46ktpOvUuCLzZ
rRQFpVjKZkqLGHb2GGJgucT1xtHoPz6P4WSSPX3M1KJUPzD92H3oziyKE54oYjhr
IwnmdT0tWtSI2Gb6X30vc0WzUYB+lwbjvgZLfOAxiyNpcGfwFsqlZjq8qMVmQuHJ
V9yN/coLjUSLYzF9JAELOSj8vtblVZhJgK1u05YL2T0iIqegCoIt8lVvh2AGViGq
JoWape7Ul2Mledf18YCAO5TXgO3e7oiFu6VRzIJZPfr+s+kEZRsDIS4OdjumBgNE
aisnHC+FBdW86+yYwWgvyf6gGAjT14UItnk1JMMb3fxdgPaQrHA1VrxLds7KWona
0ok+GITddXdgEaxeNKBiDZIb/3JsQvY8EbMiiCbMoq4ZRJxvSLVqt0OMQ0S6Dju3
2o2a47/01CvaGhC4DO7dGZ+298EqZza3p7j2/gG26bcLrqhOnRg4cXFGNCSDcZZa
9qa6T2tVNOXoBDObRueHNXr0IMM7DHDNHCINBzaUnOsUFSeXIh3JdFdKf8lHypHg
HpyZplgqTDg/mIoJPlfFtu6MvV66fNbkeL63Z1Ue2daO8tDkitYtO3Z/S+QuJD2e
JfJB8rs/T8v7oY5C/Q1XypKz+MGh2981CX1fpv1PahRNdLyUIJkmNrAPctzbAofL
oMKD8QYnwFqj79bdI9vggmjnC1PeHl0j46caaNtlbiZpMkPjBgVV3hOYo38Q0fPD
rpdhFgkROSG8W0An55Lc6uX3JW179w1TRKBk1Nx1P6bcb65HMOpgBHNG4a9CzGZU
HNlIaLRtFqGmGeGYaF7OiOHoC2yf8KLkFZVAH7KM5mbzIQj5VQGS2sYsb3cgFIei
81uypUpREcfcnjtpffUeBg9jarx9h2lnMTDdb5mBjaGrUTIDObIeHYOLpCWU3VJA
H52pXr5/UN+JhrwKD1JMTpNaVTmD5n86kHSpyHWkVSL3OACpjS7Bdw7OIjlBvRqN
WCzoM4WAv+uLAogZ5hP/zOuyUn8/ZIf1KRpm1IM0bVrjn5/ibUzimGiH20J1znOm
hPIUDKzozJQ/AG4EQxBOc31AAOzNWiLS2AgTVdRM6YrJy8XzXdnZZvuMZ1r9Ns9l
+91IJOBe9LIEG/q12LQtb+DJQh4Oa7xfb3R3pqj6YbEMDdjLTTmqObEh5Xpog9LO
EGX+4HJjynkonOgcuqIlKcTYWPotbhl64TdwQdLiIDhier0XhZ5OH0QTKtPZo2c9
mNWPnlnVfRJW+vEjj5fKf3OG4cBzddjJ/PFw8fBfkSu66Yg8dnGKp8/qa8SKP8L9
5xG4Z30jHObnjo1bEz8gwz90YfUv1VhEivoB3a2Qq+jluvmz5w6b7T5O92AqxvMv
kd8Gm1Z4eaypVtEn79Wxbr6Vd66DKf2+JGVs+pLapoyPL2Kvb8rm5w4ndOGGRYfJ
X9jH5S+VF/iu/R7grAUD4R71AuHpW7Bns2xTzg2Er2SNtRraxkEmczaoQ4ERf9ho
rjxuwC9L+rMnH5jGKJbp73P9+S4UeBXyxlovrjsF15iREKXD2UmuAtUtMNASX62c
TVPvVnKu0/jMrg9D7hb05M+1O0hI4UesRpcwNIcFVDTcOj/lj6jLqcCKi7J4tkNp
jH9Z5nQTII3I4QJaJ6rHYXo8ToUFLqODn3UGQbW104j37iOPLyyovxAZXQf1zFmJ
z7U1kDvVW6kjUOow83KC6OfHGAniYOhjPZnDqYU7g/pknzhIQ/vQiPxIdVYPU0JW
VTowD2cmIIkZ5Q+e+yyj66/Laa+qZ8T6I/wutJ14Z0BODA9ruzcJ/OWaEPShDxO4
duiOXnU1ItX+OpdgaKQRgJSJBR6Dehhh4GpZMxnm5ocft6gsOufxr41o3qGVfrS3
Ka1uOyuglOIlA800ZrFISBi3s2fdOUm8pHkDhhbjBmaHw2WV5ieOzi79YcGdUmop
xmMoZVPB6X3ttbYG0copn9otL9O9sDqknLNAjmvYSx7qTrwEheK6vN2GvEFeBr/r
WECG7kutn9jucdWCgbPac4igMyTQDfnOR8sQqwvcBmay0rQ38OAb67Q212Pr2ENy
950Rt39KZjVAwsC4NYrnBhA/nrNIM4okyzt7iVk+39IxiPKm8yGtlnlwIqbS1bx4
kEp7HLz2AFXmPjmtspIW1+c/avuDTihiy7D5v+B/UthRIaJN6fegbJwF8B+Y+oIm
nc4H+lfhKE9fZcxvI3X/Twuy5zurw6pHE9TGqgWPN/d5+9Bvowwh6nmdKXHWssNW
OfLhRIDS1vq71SWWO6nJU6SsX6rUtQEYMc8lR+OM5TcrNSg/fbkS3a+VZpMeJtGx
GebOrFdktN43OeRr4D8PYVfVreCGpxpNLde61g5Ywhr4u0oBgfXMp2KmDPuxRi90
kHTv3VuhPaEHCFXASDnz0YeTuBvpo2zapLeZsM+MoymvYS6vboVTqQRD9Xc2BoaV
EZltjOZOyu7XNiQ0lBCgpVluTgEAZ+sBz9MuuMRzDyVu1cWCV0xrS/S0lcR8tzcP
sDSaQf6tQl65sRMVPAUSldr2sXtuGO4b/xN9tyhFsxu388CJj6xq0scjfS8sPJa5
QpW+9BqZES6myP1IRaoJpsV0sLfBeXi4rGJFQTF5yqY0sNOVSeIP1Mkfhy9wB/qu
AkHa9dc6v1fVLVQcs151MS8StqysnQX8c7cn7xsvRGdnA5LwXOKl2cawmAcSRfNb
D8hkRGyv8KgRMPshSWgOOjf7gU3WDtfqFjGts6/q0n+JOCPP+8lF3YBBrr9+vfna
/efvYgQdD8axT+xJUeu+MwIajVVZWQDPXJdKGazXjgVG9fCMFKMr0TZfo2zfQ0a5
PApNxkz3C1pg9oCRXB/qQiK8R60rTg5jZnkFqF/WTNLk14uZiKjq6dMhoqYb9Qoy
NhSahmJCJRGEdAXP+2wJk23Kbk8pM0qJQj8uO//CJof/oX3QcSonHRBtliLbNLZm
+uOi0upWlZmNOE/10T1FUHbha4p8dlBscTfG0+0CiYK5C/hi81sKuRkhmoAMKIlh
573oNbTF4z3OFjYL3f8xQSMYWcCtQmefTmtx3Kui2aBNAeVAQqGbaB4usbjvbjKE
8XZtbBuJ8RvWZZQ5I5xPyLu0PZsaaN0QlrZN4EBE6HrWhd+5kuWekhc6RLBvMgic
Psrd3IhXehi0Xd4qrHNvz57knC0Xe95GfWgejP2FGHGtAFkS+9H1qp25cavy74N1
Mlo+On2NkwnWY10oDtEWlvvjG1IM+8eUBJem4/wW4NFZokmugMwyoR4TBgKeR/Cb
yeAHcfjMZDvWGt498wi7LZMVNOxSqKjzQP3frPhRUa+gY+Cfx5QjbxNy1Hljq2Hj
9+9WzUYRw2ka4BQ1tYavvHx7NpjaiDgdJPCusnjYBj2UFgKfrar3AAApVXTBLDgi
OLltF+EWMoJc5gtPw9/qy4MCxxGx00td7b2UbpSpmdpIgvyWu4hkQEpLCPMCJUS2
a/ON//5HbEmSQQaCt28uU+OdN5yljiSyRpIcJ1hFcp1AdrFYGKgDoStg1Z2+x1wY
Gy+SlREHu31nzO2Wk6MK+P7lnc4RQcPwMLFHNxbPzGCfOqd1QI/Sic/9SYBlER8A
c2HEjEVAGJbPXpf5Rq7pY8vjP/VWwZJTn5EgYEL2t2qH1bb6tDpBXQhmtvklGqwI
UTleavsWRh1Xf6FJrXitLzV7qvHhO8eCo0ssyypT4NLOrpO+1qgnQ+IuGCKOQoEk
wGXKsBgQsI0PgsD9SIVhjGVigqpkjaGfUo1SoizAhTxdLailIw+NDful5QPTui/z
62R3HtuWtXQysUsLCY4UxPYFyHfRXo0CQnlgsEVELRwxZBDYCKQ/03idxQH7BIeH
/vWdm2lakSajTn+qYazHj+JOlLqILFO4TrTx4Z1e0Rk2GpMwkWiH2YI+wMRHzN20
qz3i3w3RP0rmHLuhHug2DDz3XLSN231A/v1jnqG4vzRvQpf1dsqXSr8SyNl5MQZD
iqZmXvNK9tUdfTmFpPS2/KnaDVWmO8gVog/G3utOHq3PuzUvBZ83CLqmkUrgclze
xAl00yJlqefsEy9RFRuit7C+eOtdIKKLAfdp09gByHYDoAlprZ0DmG1WhBZgJwfs
roHVUr5kiuMs6T2omsdw1/IySR2uUbu/yvgZPncfWvK3IBgSWRw2sdcgJ+KyVhu9
gJn4L/pv0YFUXWakQJrK4ZAsZBAcyGhBcr/El+Tq8rL6oXu6gmr/AR3Aqn4muC1F
731JhmLb1bFGPddUubcG/ZjNqokU5vg1N5MWP31juF0js+ypbNUYVDbrIBv4SefR
QJktuUy3P6pWIK9oEDEolzFuXbnIHUvn8Y+SiFMxQ0ZYBONOCXZR1jym+rbt4VhU
fCnfJiOWabS+eI0nt7vW7CQPrDqFxuWurJWo7AORXVYxPb3o6MY37zD3eJtqUm7z
/oe/9bGebIePwuJoCYO2KjnemAZo+IUrLNITZJIVv9LWD3wqPcFemxgly1PFB8h4
3Rz+siXrBM+y6YC5T85Re0FCUGUnKeT8KFZ5rprv0ybfVI4xC++H0HgOyfHIsnI2
Wa3Wd1sHSv557LBcZCkYjpOaZQOnXviqfBToQnBx9TrWosK3b9Wg8nKG/9uhn+19
SRhS5rgYya6AW+VmdbgecjgDfSnqcPd5aoKGLvH9oxNJ2iBmI4A/hT+hU7TPdTWR
BaRdLjBS/RctL9X1aJvgEzSm+i2e/gs7Up8JqIMOVwgQw+kr0agDfHMd+GZ+GBG0
3DHHu8ZtfO40MY0WgsM8SubJ31Mi759LqrMRrSMgUWQH71tJ8+2DYj6mSHT2+QA8
QKeDQjxLZCL/GuOV5SH6va8dw6A29y5hflfflp7Z/xjOOuZwiMKC0yPdH89cr/jK
60DQcp1Zd+wXYldz/Uj1omaYWbQ0wZGw98/D1aKBAgA7ql8Y/fItps0YKuLyMxqh
v0bHdQTx6tkHhkIo6LJnqoRgVLA7eDKuz28eP1sSKt0UVE/ad57JZmHHDh9bKDfx
2AeNtzhG2OeGH6gbmc8FRnI1P0iWvgo5MLr1qFXm2KqBVpncpL4Ay7zUry6Egv63
DX2SSVGyGdjrkKG3Z2jMUqTUGhBR/WgQynfrHZ7YRWgJhv8wz6S4SENnTuNf380j
m8qB4cpxFrv8JdaXYszc91cZtAcuKjak4REYqsd8S/C9I0izYS3OHYsPHlqOa3+Q
f5YTLhY8iiLS+bamOjQ+mV89fEGaCsnNQzppB2Xy/f/Ji4GC0cjiY0bZYz5F9HI9
MKPEMiVlOhyL8UJ6EiEcidwKQy2x0CnFZRdCIeqj22CwCsrx2tMeJDaUgUt54qFi
gK2Qak11XLVpjjMelyBDkW6pO16xG9MhqfzyouIy+azmKKgGCVn3NyFWzoyJFz6A
99zd+SoMcwAMjULJAkWr5rFJO0mgrFidd+5eudX8H8Rj5ai5Ugw1Z5ibn4piDoXw
GcJtEVrTNVhdHKMOETYeNj7Rv81zAvfOsAO98+ZegyxLrXovwIdQmYG54U66d8N+
fZym3qWC2Ytp1NDFupHWH3StCfGZNznfCxh1FyuaXNnNvJHGMvo/Vx0t7Hk7Psgh
0c998nyKr4IK3LKm9kxusAuTLT6WKge6T/mw246vCyy5R7AbSS1REfb+aSd3j8nf
1KY64vg2EwRjowVPxjyMmRrvLRPcRBeEZUq2MSBJxz+Zf6kgP7wJR7t+4jHS0HEc
ziI0SSQ5oSYrRyXEaHw0psAJJortzl0AQu2+3rUwqoUgb3SdfJJI8JQfEsizHzi1
doFxSBBwtMFYFuiKY/w8Z7dDLDNSZblVscDReEmzd30F4rZvbxueJZVjXayQnDNO
JP6rJQLE3yGZzqHCKCWYgHFMWbGy+gt//vPUsrJehe8PpHttG7gXeqYDsj5Z1msh
n9QLtt2yUhjxB2CIuux205jzNgmOO7vEAK4G2P/ssODxdd+TaiPNnyapCUUj0SZq
qME3QNcFm7ETdpfcm8bYZkb1mRdEJoWcdjKd4+32wQrrIneaH8HWNmT+RxjFCh2Z
4l8u8mYoeL7ZxeZixV3qTEs+NBCDV6K/3f1DfTMJJ9QNBsuxZiiTVmnQExT8gELE
e+smoNW9vZTEYXpC4r8ujwMP9ugJ0pjnVyK3PsEvW/A76Mx9KVZFNwIiapqtGiyK
f4ZAbKj+z2bLA4ELUf16oAzK2WA488VromMzBJDtdHZVlLN57Ny18yOA2XKNnc5e
hVeOKoDOnZ+xExnkwKPsBaDziiwTr1v8enCgwGTz/16Vqxi+Gu9OLRXGzII+Z0+X
OcKXxEtre7acmAhjqPsU6CxRGEvwmBs6nNdqZb4nTXsSb1elCSzb8B5spE3GQ0dD
MjK9J/oJpP5Zax+S8ushd9sFKMuPQNTpfZqd2J4F+EO4+c5jpn8NL1PhycJfEKG5
d73zFhxvgMi4DEN7iBC7wGfPVq3Op+fktcbeUHSIjeMOSYn1/CqeQ69bTr0XahB4
fXEb5+QvnmRCFbrYnZc/rHRqk5H81GDiU5ljd5KsloRJo2YLtnWUxXZU9H8eluah
rd/BnFmU6DGp8sB/SXUAUCBzE3afWUyj3CTdU7b0kE5nR8jJbhwQStf+C1ckme3M
mE8jvz3CYgYFP4WkPGTF7l4/XEOE7G+rsbddRYcP/ThOOgcweLTKdtjdjNJuUjuI
6Hy52jBBZ4aZNP2Glo8qsU8GmS1ZqptvNXaeK94A+nq9rE4GgQUwRWOEYLBCQUrw
J5GpkPYTZ7IwxdwchuHjiYNMWC0elrC2RPJSg2/cfAYeH1vacq38jHNlJr2IhxEd
Xf5WDUfSEdAJ64dZdorJ10IKxr1fmFobqUcJFC7gGV+3RLwlRghM6imCtD5dYeeg
9htBs5qFO2kBxoexF0uq/NOUiaAbjz/et9G0bCid/V3BS1oWyPUnbVQ9hPJCFkqx
6aXWdmuUHVgeCf3rbul5yCWFp9csc6iX/FTW5H/9Qu1BoNb/WIrBiQ4x+VGG93Pw
6Rsl4217xwdv2Z5RIyRrrEz68/mWSt2Q27QhHQrdvCWIXKHe6asmHcNG7Z7aQ6i7
SRJKb4zIHbUmsXiN0BEcYvhea3IASltnUeppL5nbSK4E8zlxwVUEA73EgmBE9SJ3
kadYmfE3cAYY6175N4pUpevpTAQR9e3mJZ0VcOp5eB+4CzTI6fg5a2wetVP+mg/5
qCKXsf9w8oJB+RRSOFoPms8Hed6niy3kA/Sgx7LDXEBtSolt2Rp7fDIp2CvV3RVh
v1EhgdZ1ZtKphMCLhis3usqRZZU8V8i6mL/ZViBusr/C1qQhz802VexjE9jb41hY
2znXnLr1CRLfyjAugPC637k7ixy8REON3jNF/wL9ZNiAuNxCvRbaaTJgSMOIGdKB
cg7k6LzkEgsM4o/UwVTfbqQDjFkq0VkjICK/9KUEVWAkam5UXQ5HWetRHMo7pniU
cTq5sD8HRYoGLAdBOu5uuLR2dCZ8ZuiVupB3+eKCuzhxMBg40QNe/vGgjsquZEKA
rn23+kCU398i0GDhoSsbQqd5Iz5yj7YyuOr5VplWQiQc1g/DVdGJLTOCFRUsFSRb
Cp7qllLB7mozBOW40VkqzdAsBcpN/51HTL3PPSt3UZstf2kFN1f+ZYGwoEVI+CJn
PjgIhlel4UGau7QfjdC51Us7R1nQW4hzbvzliGRJCCmsGWpw6lxHQd3MWc1Bnw0r
DDN7lvypGUqmJ+hEkfOWFN19spB6jzTImNdi4BUdGaDnbJmNcvKmJ8xtL2kacvNg
ii67SJ8kbmCkA2fG6y8xXGi2uZ5she/SfmSzUF8a2mzVdL+D0VDAV2gZPcEr7n/E
dkIlZYhVS5T8weCDt0qXXgIKZB4XO2HfFGA2ZmIu/0mO0dyh0Q2v6rLqSvBJiFQ3
CGaPYMtTicdtO5ZXJ1nJwSnwUoDybZPXI+QCIr9dvZ6H69IOUCWIRahBafYt+JrQ
urua2RXEr2ss09FSPuvfhVazgw5NAo8VD1qFr9SjoFSS/zH8wSviYCW5thPusEaG
83kZchQ1OtShPtn8bBD2yoSpcURgM5lBjxgJISLs1NS9XFGPzmrfx3tfERFuZ0nk
cht+Vde4mWsGyxFhfM2a9zYWZamnKJ+6Cd6aWQ4Vjj+VYmT+16RoHThpLVl6lpSr
g1L82D00NzmXMKuHGiBSvVoy30kMGllV73UDD+3BA7YIjMzQuWfG4u2pC6kHDmWG
SCscFIeRXxcx+NAUDfoQweEiZfg59JO8Anp1GhwslRgsge1ZzzqlnMXKfahVXWVB
esqgCHog+NKubDEhL169EfqaXzlPyy9AkaE3e50S3Ul/ymGFEjqRuvFdyroJmI9I
lSlQdzz4GmJl65+94HbTaiGlUn0jKnrLLvBBgwhu2WHRb5xvRYXAWlNEksM8vgQr
nYKIuz4HoYMqqkTU4u93pGt1VfaMbJtTxRyQIXUirqkzkpq360LPJIlpFCniVpJz
yQy/52TH6ktgRCdHMEgP1NYg4DZT6DGJyOdTB8Gv7PvAQ0Lpc/Oy8sm2Ew3UYlAk
6i0+FWTGdVq32OJEN8Q62y6nz/1aVnArW0oxzEQKgtE2PwjlgNGfxuaPKUHlbwX7
hjAgORkVuw3tysJ1m8tWof0ctX5xDGcA7hJDKbZRMLx+juETNNNOAC9iBiFZCOuT
cGJ7d8D3dg9zjYS4gZCx6kDt+nmMQwNXULH7iBIj26AsahLjqv95O3xR4WQsIvn5
WCm4YEO/vMraS8nXHIMRmyGeZXae/AbcENXgQLS5YZ8zWC9B+cKoDvY6aYknXGb2
VBp4sOf2eDsivCwaAWqLS8f91fjK4oXkDPQMPxg3d89JQRNIzhzgPvnDPPOpvnvV
0M57L6gCajut6CHU8iHzePe6a56jj5XjN+B6ZdNr0To8fdNLisWnyA/BiO4Cw5+0
ISUgZf+LQQtZZRprQ75ejZ0f9bgHEYBAaypIb4KyS5QxIsopsBXnytWhk06Ga18o
+fennb8njpaOF3IE89Dme7BDxYZOPJ0N1ttCk3fB4S1Et8LwgG3ky6rP2w4LNQoP
o1wylF0LIjhS1xXHdnB3JsRGZM8qW4BndVRUXU9ebzpltwlYDWuiGvpmb1hl9ttX
B0MBzX6MH6wAsNBLkAutZ9o19/O247VLM50MPLHPhF24C6nhPI/gkkzHDK40UsEu
ZFLbB7jO4q4SD1PgwhebyHUDpOlWNqSrVHn4d/hna+nkn0HkvLAolMDMIaf15NPK
0SgeBz7nkeM91FAsYyomlnL5XqnFD1Z4HyAL2GvqTja1RpsSQQ7xMuw311jw6jLc
JEwhMziRcEGY60JFU2tFJpTVAcSWoJVzlwZCmZGPno+oar0AtiRbWFRFcVVo5r4g
TRyowIE8MRVvRwSsRrGwspfT8hAZe+rluyGtx0Ny03R/NijtI4j3MHtaVnSAiwhI
uftvrpNDUDOoDzRq8JNh1jHoOBczBPtDUzkI9uySm4fkyHS2LMWOSXnJfbQO0XH8
quU0IcdPfjysaaSaoGrLgGl+wLXv3eht+v81vB8Edu6X6IsZ/8Ho2hNZ55SRmA+Y
Ii28T8cU/qik4PSSGNbLnndU6gKarbYa7Vti6lZcN+Dduwc4mwl8TUSVSt9I10IL
YfZvfDofKbLs5v6TMS9kB5XkTbJWs3kj6L22r4hU1bDnuifvNRZ7K56Wfed4f94a
mSN1z4njEL4JFvda2iYwq9YBpPLiiNZR2TxYsJOQLZZ8DoAfu00IH8V5bf06Gklm
GG9FJezAGoqVNFXx7Ktz1mY6BhHVEkMUPkVy2BKxOYkkyfgDoZSrkJH0AcNS16AK
Q+W2DUMIyyAl4AXZ5JIXcb0Bl94FnhKBXFqJTpQkaV+zno/WMKocuUA4h9GxAozB
TWjnqE/nMntjTDnb/mDY5gd8AbWDeMXvufCBSWbfHDpTBusNkOFxQkYeYJkey8NN
Vu4vf39ZXTVJoE1BRA/Zfjb4Jp+Lcph59gW22YU+rm43R3SL/ASR4PerM4yg89wQ
JEes0AYUZEmbx/akZyFXjxTNlCcNjhJNXuN7LkZuMh54t4N6ItcgMPyzVlQHWiKX
wd/GUPjMHUfz4c75uj4nufa4jmsXdJaJbXDRjtCSw9gKLnr5vDr05TtQqO2Ersu2
K4CiN8cIw4jF9gVoeXT5MnQ/KgN7w1tDYRsHWtjVV/dNa7wUmDTtwKQjqBjMUeBp
y/BCWg1vjWPmc+vi4R0IL29j4wKcWV0Pi+KK+PVRbcn7A//NrVcd//e1vu0Prk1u
gPFSJ5RxeiqfXe5x41Wrcj9pV8L3Ty7hyXj5QeN+YQzx7qvmWt674kd6yIxoht44
s4a7ZvW67tosMtEvZUi3maAy08AXmZ1iQySM+Z79ZCAZvYXkhyHaHjSTUfhFnZqc
2xVWcbZnpKyjDmO9KPeCRVHYP3uaYseYqH5BzJfWQyemS1/29i4gi99M3VTCCfJa
JOuUDUcIdKVP+NRC/7E9frrHGQ5dIJQJV5qQS9Eyk6HDOq1anl1Y3ftVMaU/1BEm
Mk7sJg+LiT2KHyVG3f483PceFc4F45I38bkU1FsuFHJY/2m/38lLiS22/M2SlcTD
S2lbj8ffhoBSRCrZnysCg00WOGtuJ1u/+bF7orc7bQVi/WKTMuGWjepUG7rq+dSK
sesI6Qx90qqi9qh2DQ55Y2BwAYQeTWbSgnMfqB4MdJVF6qc2NWUH+Kqf2HfXkSBL
MzzzlZYhlmqQedypPqBtydzvbR0fX8+IgVnJuBwLHK3pI4zh4cF7s2JZmzeCAoUu
LVbK0eArJDKWXskDVqupLnpD3Gphv4JfMDm5zGMqq2MvtmXPYtrrQkqGofE65HYe
DnSZTu2kqBtEzflcldMiQtCWydQTWYXlvrAqUpRXUCmc7pYHEve06pfNq/teTJrS
TRPYifTeezaZKuuAGeVM3JmOmU0/r+CmlMg2HPWHE06ClIRLE928TzUSbwzsfhN0
NII8xvRsfC9QPZhlMmn4uoyoiKeLKY9C+rh8ZlhbORfvcPSGxH6fI7H8VRUaKnol
WZUHpounKRg6hASBYft8ZKh3qPe9ve+fV4TvezWcMIyfCuEYMzJtQJp1STstSIPo
UsMIr0fqHjIOFtNVTQntexv/S9wWqXCm0Pu9dCqallIUkFvcUT37PHKWcBRQ4HSm
qtell5OHQedvxwOhjh+SxxBhTB2Q3/uVbioi1aOlfHafJG3+iHy97kz2Dz+4gQBx
ZuDi9PYGirPxfJjhHtuDHNpCumni/KC8LYK7X01PH6eJXLnhAfwaSg5TQexu1xDI
r4132SM5bBsu0cIK6BBV3I9LNL6MM63Vs0Oajcwv9KuKVpMXY9vEUqogUYdw1Smj
3SSFfMuQ1xRFIIqHZkdAv2VAZxwG8TwLPUoKHXHFMIeD0olhBbQO9NSoa1c5MlZw
6LKZ0vPz/Pr3f63KR4CNUI6YjOAE5D/ilGT06HQjr6Xsz5rhhYQi0ORcun/hS2vx
+0s59xNRGXuqcuVI5iDiUzKeeScRleLqBl0vte0YnBuleDX7Glw77TT9ZUqrnwbV
0Fzouep5q9ot3eBef4yFHZMMvFqsIlpyVpDlSCY9kUCYaO6FOCg/eDng7TPL47K2
8tJ9y30uLtmADfgxa/9xbrkJM7errglBvWUel5U5HLE0gew0hHLXxcvNrXFyLJGc
Jy+kVLllwRd5Y8+xk6mcEzzjFtZFTPePbiWU7CvfjHrEdjLnogY94L0lMJgULEPK
VFV7VaWgWSoNyVVEA+rrPfEE3nFXT2Siusgnk5sxTkI+BGdzIFInZ8cMOH7b89+A
vRPS+cz69p6745m+Oa3XAup4O1CkJwNGdqjcmBVfs23m5bLKuIpxtJZN/RBHGNHL
4cBfGcE7bjqgLX2b1VXd60fjh/w/PLUosArn+RpIPs9IAZJl+4ICpf5Up+e5IqFj
xDDmRQ2LZ9CQ64pHNdG31JjzKPak/WNZwMyUOXk0P4aazEN6BzjZ66jDaVzi+hgS
a9Y1oNrOrkztHzngsYv/8Jb+J3mkwCF7oS9Es36xNkgbKfqUC9RnwZnHde6QHlgF
9nT+U1BFOClhY3DcZC5QFfNCONy6eqsBPLGBwnxWv6/5tMgEYn2DWB+6B9vFrtDU
vOZdXIJWqmrA/dJTfyoRKbHSB8F9vI1aAnDoa8f2ScRWUfObhXdDU5JEDPzO4nRy
1t8KlyTXKizWSfZ3gKTYjQlRKTuPd/n0jFDlWB6v6ZXlIfEQCwzwyis0+sG2Ev5f
7I0ZxD2aZ+xCpsSMDVGXbLzEmzdwJr5isw7FW3D/mcIetVeLN7/oPjHJwhWt/0/J
LHUwv+7EI+iXTnkrLNLTFymizuRzmgou/uCNepyXeoRjdiy7SF9MhRVKpKCEXvCb
PK8aBbohgttq3o2v46jT1V6uj4+hM0e1R2qjhfLJ7FUjZJVd0ThTTjOaJY1cx+8P
YBct9qH7aNHPjHcLGpiK1VqXqdVxWw8hx4nJIhloMDnsXATgtUqS4ZCbp9NJ8fJ7
iCNr5p0oVCl4+J4VzE8p20DO0Avaca8lr+S6EIBNbId6e+3C+E3qtkBvBN1QO7cq
00JXxFTyGfnVsrk4PuzXIRuNzKpi8PY8Hcq2WMMFScjwvbOK51HBnhiLixrITjOp
bqwkl4qMfUmtv1rcPUBXV6nWwunICYmrtWbokrN8h1ap95B1sFuz/ONOwbVfmvaw
1z4NBxWuud6FMRYdmlDAd6vJXbY7ZCv1qc/IaoQYq205KYb4d7PbW58Ma52x9OxK
XaThiWMEVZACMBfYDzHG5EKQu4eGuSGpslfgjWYQM7HEAaeSdSbcpeCH7cfButCb
0M+CSZQ0DhUCTuhy/5Ihc2IInmgNqrXD7yszpuS/0530xvOGdtB3bqcdZ5VhJErE
Ja8UG7SA4+3KbNDb0G4BOlJzLw9tFZbSEy8+lp6T55WPkf5mtOnVAozTqUQbvlZH
QzmLW74EiSVr51edaaXq4WAFNRw7ZS6abN3IW20aeMZu3jzTcyVPJicEgLiiCl2I
f0yDwCCuh6dTmucgYga/vX3Jd3wCXmDo5YBeeKQmooMhM+KIFndsHwfeBCeBqGPa
9CEOZz57JLhVIhpO6zKdhJxABGT93f05LmSEV82GPWsyCPjrQvdeJ1rVeabUMquI
OWwmL7ANZDib3aSzS/dChV+620lpUTkrmL3n3ao7PmTE3hWq4CTRHgyhX7dYVcHD
C/jAuV/qbGXAz7C8Ir5sLTiggBLnX9LV6CRjLYors6TNfcRnt5/srq1lIfSOMCIr
H49ByoZdavdokjUs2dQzrnoulTgoUbTbyL4/B1GBRwDRVl6CRRsW82pQto1Wzaez
/iKziAiGX1DbV8NiN9cg1mzSW06YINb/1+Q6UHO3kKG5MnfI6eCtagd0fzOwGYqS
B+seLvQOUWlG+CwsdQdpRdvyULP8MWwppIjud5JRZU5zkNhcGgSnszbVN+V/kif0
N+dNKWT1jjqvwzfE5zs3lMuUa8uhp4chxHam2dAH2pH91IMsFUEkm0MwJqaiFg9M
tZB488UtmNgH8WA4QNgNPacH45mn1LW7g8dyTtN8Whg8FKwuvPhIlCW7Gh7ihO4B
7aCn4MBK+sZYk7dw0h+uzKAB3fY94zexRk4uWgvno8x33EIaBf5n2d+Ar2m7vU/p
13Y68++qrIzZ+kEkTC8xsav2YpevQR4CUQjB+GLnpkLIUxIFG2U84o1FXijt0MEN
LrnQL4rSseGLNTSl0I+fpx45hr6ypZb1708dUbqn3zfvYN73SiAzLjjIm665uGK1
9FmyFEzWTXpL1dfyUjioeyj3St6bcDI91IdVWqM6GdHrQpAI+WNR5e5C6Qo3rz5F
Ih2j3MFcb8CLm6eJpzrFnFo144zodbI35PzwQ9QhtHahDw8/SE6b4RLZzF7VmzDb
h6+87G3L37SH99MC8APIkQicvOHMzr7lAtkyJamMfRIlS/jZxjogpDWoELjk7dkR
Z1MrVC0F27KWr2sDn4Rr+Yc1o9O63AkugHDCvbvmD1YNCsxBIWrGZhI8vQSdM/a3
r2XIHWt6KhU3ySBWA3xY4jCC60o1MkkodtcMNyd3L6vO7g1eG7TdY9xRUm7dCXew
cXgOvG2DvI1rXQqfc8AUKLYKMm7kdgubbmCIRsY8HHxjlVdqFgbwk0joWLHMk+3W
8pp/jYvq5wopN0aeTB3LjO/foxmhSqzuz3bPfGq3yt513amUCL2nBeLZ+EW09hj9
kd13Zj8VkTsKtZh8RiwEoke/m5fRoClK6aSjcMbDUak6BKAWAwsIXu7spaz4Nwyp
jIAKJTspNgEfhUSnNBFBY5L5sdCRneT4qWraIHADE3VcCEmaDVH6gtHb3+OD/NMC
Hyd3YJPon+e6fnuDnI1mrkpZ4kbooqqAp31BtCl8elJQNCTmeQlu48KPEw6Wf0jX
AXLjNtlXU2gk50zWsFyn5Q5cmZmqZ7FR3sMApxlB4LPP1q5qygDDXZgRA1G+vpPx
uObMYDUavzWGB2PahiJGZINyEBeIVqqEWyVvkCuQClXEoR/0GeuVLsuFhwfEqPpc
mZ8Td+g7AEJqnnO1OodXI4dQ5kaEVOvep9IbqXxd5AzZUBRhWcO6pjTT1sM999W9
t89BW3HBMIwbJujR35Tc/Y7huSJUYqj67ZLgDXaGsUYqOH3oe2sf6Iq5c4B10n3a
59v888RT7lX6H9KWjGBli26UkI9w5Kzo9hgfvsn52FClfijjYpzpM+ASKPYpZGUS
dfGS+2sIa2twx+GqTylgESM28+ssJXbaYNtxgO+F8+Ks9nOrTHOus1zbMvdeCcgP
99YN6Kls2dIJ86vATGlotAVsvAyFEyAcY22a7NiPl3fyw07KacGN+w4X0yv/Upy6
dRtjyhxLGO15MRxdYeOiD7U2m2hXAa05ScMx6DZxtt1Dj45WPcIJxcazt+pgHYMx
KDBOIvJzpVjQ1MmK4rVstUypWSUPzHr0d4BaTiWWRAvkobXYjvJEeu/5FYDwNkDl
rpqIZqZNhsuVribymOFbpWO5LnAm5332wtB4w1nh/Y7H9igbvS8Q4HQAFAk/PrEL
BbOBVnZkDBdEdWXF2lfqjqZ7xj2C828Rq/PE48e0BuOUkQCvOOTGXjyobpE9pxT7
nM0L4GtwRmTZxIpC31gQV4vchTrQxBh3cOqFA2ltR1H8g/m9oCb9zuzqZqvVJN52
7xT91iaojPgnHPIgrX0vrVQ2sED8/zJEJM/hXLD6EKw1zRk80yKFE8FSot/4wunz
SeT1ImMtIwpHnWet+ImX9faERR3q4gzQy9tsEVyE1KoYyCt1c7dBrABa3OxQ8F29
BkNq7HOi0zCFyMyDp101ml7rIu39LCawrXSLF/XZ1N5DP2vIEuL39BlmZ6PDjdJ5
gQzzZdtlsNoi0G8om5zlhOGKZ0aXMHTU+TZ6P/l54hrbyJUE5lwhzV+YfBGGq1Nj
biRhwSS51O6maXN0XZKQkBlkCmMtD6l29KdrCFLwxpJOeo+nHUyVzqUrhVEkus+Y
GWAOiyhCuUB8Yij2pTSCq3vKytoigB0pygMz/MB7pgkjusdC/KzkSJv6XPQDz78A
Cn39Pfh0gx/l0EDCl792efEy6dbAQVRfO8CV8kMNcEAVBbK6mkDTctkNnTz5qjtW
qexKZXCXMRzciy5UnA/SMIZn2s0qG1aksthgxv4ZSRiGMbkAoSdTi+JKKavS1iyG
Kvs7hhX3GUxdf3P5vZhe+QbrWlDNF1gNyK89YGgrSPFyzebayc5+R6vPVr8X2X+N
9PltQ9WNrtJd3I9oTcVSQ4PjsSKVJhWp9OqBQ9eDzIJpUn8eNFTgIQJyVadNzxop
emJu00kBYwXH19vhad9rygApjSOW2rLbJv7eVvYRHW4PdhjRyZMD9l91eFIY8/Qg
CyIqmJzBsZweAmMgA6AOmY8eGHuDdvIFoEwvRi91dqaq56fWN3qOY+NZt7xi15zg
jXPtKjJx/tczMoA/4H7bSkEC7C9EiVsT+2q4+S1/gDynyyOfSnbMl/0QL0f+DKVY
fv/HN0EGx5Wu7QQcBolhUg7IDYDnYSUCZ1bcp7MBFs96pRK0xnfkBS44PDULoDLW
5a5yrE5u1pXhGAtsUMDvaQNyPzZAqsQwLd6bUZED2JsHGSCTBBmYCr2+Te4iCX/5
WVVCitveObPURvavj3WIOJOye6EMlOlzcl1wrYgz0G8tsXJUq2TidvrbIJiL8QTE
t585DHsCor6GmnBpCdZI6P0gKi4rFlgLM3boGgP3fjMtpQp+xZHkTr2+6Z5ulokj
3UggJM5KJj9XeNXW80L4xTlsRJLRIFPggeeDUmjXH7mgBtDzml/t/3ZP9vBv96D/
KFUtik3IWitVb6fPlCHATc/pQw9aQ+1Ce4DcEUaNSaaXFmDImUpo0e1SmTyKZ0PJ
rCLMsfQKPJHU0qBWc6RVJHjOCvbarTqdeKBmVRo7W6BE6jv8qkEAeeulwkq/KiTk
Xoi+x0xtTX6p/jNwhbzPMt75y3XMWkGh/I68X6Iu08yGi26Wf3fpb+Cxn40VpXsl
aQRU4vzbqwhIqdjNP3HAT5i/HCC06ENzniCQ3vfX20CxENKJBsYo+E+2RLF0j0Qu
iNGB3wr2MOiLq5OmxbYmvrPkPMkSi1znirfKXTwNR4bfHcls5c2NT9F3rP/0uqqt
uShFxSSAUJLqSIyXSSRFcUNoEVgukkPviQGWETkr6sa/2wN6i9si7VDD8onmh1JQ
9lOPvmfJfLHI9NLD4mwOdWT2UGoQbXYbMQWnxEEh0uKcShdr1+UOMJRDkRIliGaF
CpbtHsQ6gD9N2mY9zs5udnUVJoQybP9k17rOGeoKJhfxRSmBQzc/mQE7olr/NtgE
ne8upMNHLlCBkc0efguspR/bsWzIm74op/UMlzQk+78t8xGXEfXxRC7PYyhC9t1v
GXWrql/ls+cw+3peUvlrIM0bFp9ZBhMOVOws+Fd208uz46B6N3m3nl32cLvFRUU6
/nXLZWlYTCYrf9Vq2TryEz9JVLfxnpl6xMHdPfMUWaqsbMuqENTBNHTnoMELcYO5
2D3mn3lq7BRakS6ib26T0uaDBFYTENN69wgrPU1vAiwZtJcIcAWGNAilRQs1eYK9
4xQR01Er4DBDj72i+4mVLYDdex2ZKds39dYwZzRH0K+j17pSooivkLCGJxttylao
vv99yoiLeN1pC4WK9GMBVogNPIPtfBc5tIllTOFNx7A0cXfRXD51DqDwi4Krxt9V
OcTtWNKT5xUzYIZep6/3RobAB8SOl1dmcjVMpiobdkfoc7ejp2leF5QiZ2fBL36k
rYVSmsS8CrYk2hi35mzyPFT732OKe/+IEJpjR0xCy5vZQv0fKyCWwuYIODpZPz25
kAbN8AuMjo9Qfb/JbKF4MsbNq+5UEUg9n6RJG6PmRljm8bN9a5w+pHEA08cRu80q
iv1FQSyvDKi1KhmHT4DdJKFfAIu6tBoR++SbEN9AfYGmWducVBnUeNeg3iizvMRP
TEDQ6ricAZRnPhENedM9NCbZJkcHlUrZkplbEKoeRVfWDfI6UoyuitGzCV9VS3WS
`pragma protect end_protected
