// sc_fifo.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module sc_fifo (
		output wire        rx_sc_fifo_almost_empty_data, // rx_sc_fifo_almost_empty.data
		output wire        rx_sc_fifo_almost_full_data,  //  rx_sc_fifo_almost_full.data
		input  wire        rx_sc_fifo_clk_clk,           //          rx_sc_fifo_clk.clk
		input  wire        rx_sc_fifo_clk_reset_reset,   //    rx_sc_fifo_clk_reset.reset
		input  wire [2:0]  rx_sc_fifo_csr_address,       //          rx_sc_fifo_csr.address
		input  wire        rx_sc_fifo_csr_read,          //                        .read
		input  wire        rx_sc_fifo_csr_write,         //                        .write
		output wire [31:0] rx_sc_fifo_csr_readdata,      //                        .readdata
		input  wire [31:0] rx_sc_fifo_csr_writedata,     //                        .writedata
		input  wire [63:0] rx_sc_fifo_in_data,           //           rx_sc_fifo_in.data
		input  wire        rx_sc_fifo_in_valid,          //                        .valid
		output wire        rx_sc_fifo_in_ready,          //                        .ready
		input  wire        rx_sc_fifo_in_startofpacket,  //                        .startofpacket
		input  wire        rx_sc_fifo_in_endofpacket,    //                        .endofpacket
		input  wire [2:0]  rx_sc_fifo_in_empty,          //                        .empty
		input  wire [5:0]  rx_sc_fifo_in_error,          //                        .error
		output wire [63:0] rx_sc_fifo_out_data,          //          rx_sc_fifo_out.data
		output wire        rx_sc_fifo_out_valid,         //                        .valid
		input  wire        rx_sc_fifo_out_ready,         //                        .ready
		output wire        rx_sc_fifo_out_startofpacket, //                        .startofpacket
		output wire        rx_sc_fifo_out_endofpacket,   //                        .endofpacket
		output wire [2:0]  rx_sc_fifo_out_empty,         //                        .empty
		output wire [5:0]  rx_sc_fifo_out_error,         //                        .error
		input  wire        tx_sc_fifo_clk_clk,           //          tx_sc_fifo_clk.clk
		input  wire        tx_sc_fifo_clk_reset_reset,   //    tx_sc_fifo_clk_reset.reset
		input  wire [2:0]  tx_sc_fifo_csr_address,       //          tx_sc_fifo_csr.address
		input  wire        tx_sc_fifo_csr_read,          //                        .read
		input  wire        tx_sc_fifo_csr_write,         //                        .write
		output wire [31:0] tx_sc_fifo_csr_readdata,      //                        .readdata
		input  wire [31:0] tx_sc_fifo_csr_writedata,     //                        .writedata
		input  wire [63:0] tx_sc_fifo_in_data,           //           tx_sc_fifo_in.data
		input  wire        tx_sc_fifo_in_valid,          //                        .valid
		output wire        tx_sc_fifo_in_ready,          //                        .ready
		input  wire        tx_sc_fifo_in_startofpacket,  //                        .startofpacket
		input  wire        tx_sc_fifo_in_endofpacket,    //                        .endofpacket
		input  wire [2:0]  tx_sc_fifo_in_empty,          //                        .empty
		input  wire [0:0]  tx_sc_fifo_in_error,          //                        .error
		output wire [63:0] tx_sc_fifo_out_data,          //          tx_sc_fifo_out.data
		output wire        tx_sc_fifo_out_valid,         //                        .valid
		input  wire        tx_sc_fifo_out_ready,         //                        .ready
		output wire        tx_sc_fifo_out_startofpacket, //                        .startofpacket
		output wire        tx_sc_fifo_out_endofpacket,   //                        .endofpacket
		output wire [2:0]  tx_sc_fifo_out_empty,         //                        .empty
		output wire [0:0]  tx_sc_fifo_out_error          //                        .error
	);

	sc_fifo_rx_sc_fifo rx_sc_fifo (
		.almost_empty_data (rx_sc_fifo_almost_empty_data), //  output,   width = 1, almost_empty.data
		.almost_full_data  (rx_sc_fifo_almost_full_data),  //  output,   width = 1,  almost_full.data
		.clk               (rx_sc_fifo_clk_clk),           //   input,   width = 1,          clk.clk
		.reset             (rx_sc_fifo_clk_reset_reset),   //   input,   width = 1,    clk_reset.reset
		.csr_address       (rx_sc_fifo_csr_address),       //   input,   width = 3,          csr.address
		.csr_read          (rx_sc_fifo_csr_read),          //   input,   width = 1,             .read
		.csr_write         (rx_sc_fifo_csr_write),         //   input,   width = 1,             .write
		.csr_readdata      (rx_sc_fifo_csr_readdata),      //  output,  width = 32,             .readdata
		.csr_writedata     (rx_sc_fifo_csr_writedata),     //   input,  width = 32,             .writedata
		.in_data           (rx_sc_fifo_in_data),           //   input,  width = 64,           in.data
		.in_valid          (rx_sc_fifo_in_valid),          //   input,   width = 1,             .valid
		.in_ready          (rx_sc_fifo_in_ready),          //  output,   width = 1,             .ready
		.in_startofpacket  (rx_sc_fifo_in_startofpacket),  //   input,   width = 1,             .startofpacket
		.in_endofpacket    (rx_sc_fifo_in_endofpacket),    //   input,   width = 1,             .endofpacket
		.in_empty          (rx_sc_fifo_in_empty),          //   input,   width = 3,             .empty
		.in_error          (rx_sc_fifo_in_error),          //   input,   width = 6,             .error
		.out_data          (rx_sc_fifo_out_data),          //  output,  width = 64,          out.data
		.out_valid         (rx_sc_fifo_out_valid),         //  output,   width = 1,             .valid
		.out_ready         (rx_sc_fifo_out_ready),         //   input,   width = 1,             .ready
		.out_startofpacket (rx_sc_fifo_out_startofpacket), //  output,   width = 1,             .startofpacket
		.out_endofpacket   (rx_sc_fifo_out_endofpacket),   //  output,   width = 1,             .endofpacket
		.out_empty         (rx_sc_fifo_out_empty),         //  output,   width = 3,             .empty
		.out_error         (rx_sc_fifo_out_error)          //  output,   width = 6,             .error
	);

	sc_fifo_tx_sc_fifo tx_sc_fifo (
		.clk               (tx_sc_fifo_clk_clk),           //   input,   width = 1,       clk.clk
		.reset             (tx_sc_fifo_clk_reset_reset),   //   input,   width = 1, clk_reset.reset
		.csr_address       (tx_sc_fifo_csr_address),       //   input,   width = 3,       csr.address
		.csr_read          (tx_sc_fifo_csr_read),          //   input,   width = 1,          .read
		.csr_write         (tx_sc_fifo_csr_write),         //   input,   width = 1,          .write
		.csr_readdata      (tx_sc_fifo_csr_readdata),      //  output,  width = 32,          .readdata
		.csr_writedata     (tx_sc_fifo_csr_writedata),     //   input,  width = 32,          .writedata
		.in_data           (tx_sc_fifo_in_data),           //   input,  width = 64,        in.data
		.in_valid          (tx_sc_fifo_in_valid),          //   input,   width = 1,          .valid
		.in_ready          (tx_sc_fifo_in_ready),          //  output,   width = 1,          .ready
		.in_startofpacket  (tx_sc_fifo_in_startofpacket),  //   input,   width = 1,          .startofpacket
		.in_endofpacket    (tx_sc_fifo_in_endofpacket),    //   input,   width = 1,          .endofpacket
		.in_empty          (tx_sc_fifo_in_empty),          //   input,   width = 3,          .empty
		.in_error          (tx_sc_fifo_in_error),          //   input,   width = 1,          .error
		.out_data          (tx_sc_fifo_out_data),          //  output,  width = 64,       out.data
		.out_valid         (tx_sc_fifo_out_valid),         //  output,   width = 1,          .valid
		.out_ready         (tx_sc_fifo_out_ready),         //   input,   width = 1,          .ready
		.out_startofpacket (tx_sc_fifo_out_startofpacket), //  output,   width = 1,          .startofpacket
		.out_endofpacket   (tx_sc_fifo_out_endofpacket),   //  output,   width = 1,          .endofpacket
		.out_empty         (tx_sc_fifo_out_empty),         //  output,   width = 3,          .empty
		.out_error         (tx_sc_fifo_out_error)          //  output,   width = 1,          .error
	);

endmodule
