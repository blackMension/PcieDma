`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qMqI3eSmdXO3tlge1uYoAHt7v55BIeQ/eyA9GLwfdf8KfISc/DdiM1CiekJy57YQ
IldcaKoEE70ECnjgyTMBjFzwCLo7v+ODLLsZC1mqgpf58uJ0IBFprTynCHM+Iy8H
EW0cC45j8AeSxDJfqpK0c1rW1W0ntjUJHsZRvMKq4Pw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
3pv0ppFWKgPZcMnQDhcObLDGENduLcboOHVkZgs1HO6DYbeUb0guXCVfTyuSKgn6
/b3SvnoGbMkvrqIzfVYLLRsnlyDqcXPW+QOtk+EEi/mafP3s19hkLVuywsM0f7iw
5o02AB3LipB9bcuM8hsn7X7AegvxZDgZacoTu13jz+13ic7eDcUKSqNyjow54o8E
xZRKTz+WEkItxTAC49SVqWTZDVjYvxiBx+LUTDtH9QqVwmQJnzA7SQfksQ7K31hM
tzREdbQRzcRSP3rMwh4zGCBoO2nZB+g1/GxSLVQQh8btROeSzabVh8GUnV3wTbiV
y0XU8MIJBd8D/KGkD8r+9NgzaVRbPLMaQnAp9LihbpOQIFTKe12K7n0khliq/mQ6
mzgjnD2KkGlZayAtMIh4kD/N5w9eOGqkuOwbtIkvtbZTw7BAo3rMU/BkzX3PmNtj
rzhadNBcN6hCuKubbO3W4l1k47B69vFYCcLhb3QwjsR6NxoD5FZc2f1ns3VWv5xe
kqhAYn8yqnQg4a8RrhaY3JwMxkMpaVe4S3I8g8Y4u7ArbFM36RyAm2mMG8iG4QLm
BGM/pJr2L09Xl1bOALRbk/8XU0p2y7xruElRYPIYj5g4JHgTOPrhulAOZl1Rnwfa
kb1X7oep6K7pScN++QAh+pI/1JqJCSeolnhNbGJLAajB/iiYvcGWSkCjZhsFQ5vR
y39xpYPn4W1ATpYBFm9vcE0qWzcm8x4+6bv/5zrF9+nhGjxxuJLjgq7T90iOO5Fb
Pm+xpcZrqlvgKl/rei4aSusKKBLnZybj8OiiZ6eo8Kkea9OdZS4+9S58Zhb2ddKU
GAVE1ifejkXqt3miOrpwT9yzJK1KBabNhl/sOVBHUbtsH8vFFzg2lpkeNScJ+R4n
sQB2b0lz/PAQmYB7RsHSP5gUo7QEd15AWPohhAxtxvPihFkmB9hA6gM+D6MuiU+D
aJsvUZdu8WJGwZaxdHRzaIv2X1gxxh2Vs8VXGlCFid+sdOjBAOXazED4pHLAJlCR
/j6BwGGAJG3DK0gS6k+zBw90kDgiE5cBXh+RN8EXOwi2Hueu/zTxjoyWYZamA9g2
SZLcSeVIAWXNuajqL/pj75SlVzC8tEuU76dB4H0S34bVnuJSlxOEozVIoQv2lL2+
JE7LjflKmGeo5I+y6CPyxcLCiL3qZqIa8lNJkg/7BWKoagCAwvjtvaOHPsSJoBX2
kLmXX31I5nlkfEwm9Lt52v6maNFs6vbjlqEd6fqfUhxF+fd27qg9+bE5KogSHcGE
CS1S8bAWn+HiW8Z2QzVF//+qenezvrXwFK7KV9+a5rdFQO1AnG+/m3p61URU85NX
1ge98E5MPoYDpWJC9qbucvjuoXbmc8NTG/Ijmz14sSYOb8adNZT8QwiAocGTKy6+
G2SjoDr719aAoY9WkjtLznAC0Kt05leyozvVblQ8Oyey9CjtVLJhuxrTyStm5iuZ
vH9xkLwxUg0zYNRUFyTlE5A99O3pcrxofFbJlIlJpkUSskjg+Y8F+RgxnlSYx9pQ
iPgCKkOpYrHc7p//e7qWlXKINe8I3gqjzM3zxdvVxGzrMRt4ZVu3HDmI8TaGtup6
V6DRDGZYV/W/DErg0mKYLL4TV1XixDueCx7GiWAHqpgkrFodyrQ941iFH1wVQGb9
nQ/tIsUQI3pWSLxhQKvYSu0HNI+CfoLvIiJhRSSkjkUA9wu7rILoW6fjrXgdYwQa
RC4hFdNoEodsf67bBRE1H8KgopfTtVy4tCb0bW1qmmEnTC5qxjYW9/PHanjRYGaI
tS0vYDN7DUKGVY/8eFjzCN+vjeFOyzo5Axh5EFhZ/IMdEX7pqKe72INk1KliekwL
fHARgObwakfPUvtKrAN9qTW79ZsVS0tQ6TgWdslEjCzVz41GQaykjNyg+bvATQNI
suy+Q+SUvd4xTQR0Ecxlpn6jidEzIZKzQ1mXI7lJTy19uJJewQV8ClKqla7dwRWV
4ccn61Tyz04U80FoS0D5OhYyh/Eqh7WFVHXebMxEbbaiL8r48mGS+pshMIfB4eg0
bgcHi9w31Uwm/HDu/nTTKAc/M+5LpnC7rhBE/IHMR5vRBaVTWNaCvIc254Si98c7
QU+n1X2NeP88m484kRFP2KsC/c9FBmldwmCO20tvoBVCaedQEW1mIPxfH+TBKAbM
OT4Uup7jaYMwTeYCfcVgOhJvZnoxd3lwtgrao6n+F2/UFQaHqRr65zwVEo1QFjDk
sK6h9dyvsEzZNKrZp3sUozE79Q1+PcbOoSLyf8AffhozbF8m2Bv3gQs4R/WdfxiT
lUb+joGPBx2U1lHHtP3nUqchj5MSPFGrvsnMYTdpHBTTGD5q8IDOkxpD5YxgfiZ+
rqofV/mEW8c2c7eszcVm0En58PJOL0//4NJMcT1w5ndFIGaQP6rgDL2F7yHNr5TQ
1jaYxRb/KFR9WOzxv9ZhhUaow9iRboxeyeX4QQn03SyvfeNbMTUA8FDbVkvfFptg
6WFkQJYbs9Knk+Kmg3EsLapAPbhbgIzVANRmZ1vwyWfhw9hu8lqx8yzMEbNVSbbn
idatiq5k8sAZPTWMuVWOtB1afTqNGv0R6NJGK+PAE2zwQG+ui+owBTPDnfwIt4tp
ywhq4ufVumL616qscMgL/190SR4lvfGgoI5IvQms+lDrt6Z6vVHrPFELSNgLJD2y
VlxUqaCAs5+uH/XGNZS0sDHPfxhreJ1Cf/jgpqd/Iv+UT5BS8j3zGBnVj2Ytu2LV
11JJdLXIc8LOk3M7CqhnCxDyXvuYMBTByUsDngUPISf6a+VpiOuRps8g97yRHqJz
K0ovcnvmgx+P8tGlZCVcTjeo7jRQ9aF1gvSdRiuDM/u8x4QPwF8/hGFLz/oWWAKi
Tnk7lM2uT3DkwPewrWMcmKKvPxNk9hCFecjYfjcdTDot8OnBJuBZ17naqSDEQLze
ZeVnsGWYcs54eZLlHaZCo09fcD5JZpOmkDEmfKQzIKlq/hIz8e44lPFH/yc/SG4U
W6A84L3KXcRf+P111DhK5hHgR5+X01SqbfOhk1ljGgL/42x2mYHtufpfQMB89gxM
QMWj81E96IrbRm7/JBYu35mJc6StxQ+1miLd6HWZRdgUt7DLdxNUPhdN1F9AHHq2
LL6dg1Njp+LVZoqq9K18nYl/rlmjhwAJN/ZVlnM8/sQ8PqM9+qJ4zEua2Od5bML6
mJMGyTWGwGQ37o8y/NOyI6MLN3zBbTQXcYGz1jv1LHU+K5+pCTpnTUfuXrsu16tX
PV3AWhhTTODis8fDefNMZXra4N8VF+tMASDlKh7OcMquibJxwWUayJl8CWpYYnJC
gpZCsE9yqIaoaVpvy6lCX9zGD+k8E6d9casmv4SXM44SeNKLW5ApGUUu6M4wHKkn
NGzoDZ9NGya0T5GcxdiAUzjisGvhxaKiP1KUIf/Uyy2CNedHIi4R5KVmsfAJjprE
vkSZVmRwarj+rrjFxhz3aHHHwrzgHt9vPl/k9gTJjp+U/atvnInZ9r8B+C1gRqtK
WzYAWca2OjlcTgBT/jYQAJmlXhuYBrLCDlXI/7V9HtlhYxXwPO3xByle0poXymuX
G/l2mQ85IFphtPiTPnmogJFTPDRVif+G4q+o7QwlHkZkl2N0sRzJ9S+l9t3rltkW
MVfpTBO5tUNqVEtmvhty667pOezFG1BsDHNT4wb5vwZlV77spmO4p/I7PlcEIWt9
V9uxcSEP7OA3GRXU08Nwvo3tY1ytP6MWU+c69G761qA6DtW0qVeUSSAXFzYiu/x6
7j0XBhO38dbnnuDO0NRpEu6B+mRgyhQrYiO6stM38DBqxrXjaaBalTWzlY8pIDcV
YcYOMl4nHBwfuRNdimF2r4ja39IG+ARjPkae5D2i6ojEcG1+1ed+yW8uOSiVbhq0
epYPqT4bv79K5HSdon+MSGyS+iiUWREtnzD1MMSLZuDOh2O3v55hbc03fl6rkwWO
OoWg/DyazLkUYdKttfNYtg==
`pragma protect end_protected
