// XG_tb.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module XG_tb (
	);

	wire  [31:0] xg_inst_csr_bfm_m0_readdata;                 // XG_inst:csr_readdata -> XG_inst_csr_bfm:avm_readdata
	wire         xg_inst_csr_bfm_m0_waitrequest;              // XG_inst:csr_waitrequest -> XG_inst_csr_bfm:avm_waitrequest
	wire   [9:0] xg_inst_csr_bfm_m0_address;                  // XG_inst_csr_bfm:avm_address -> XG_inst:csr_address
	wire         xg_inst_csr_bfm_m0_read;                     // XG_inst_csr_bfm:avm_read -> XG_inst:csr_read
	wire  [31:0] xg_inst_csr_bfm_m0_writedata;                // XG_inst_csr_bfm:avm_writedata -> XG_inst:csr_writedata
	wire         xg_inst_csr_bfm_m0_write;                    // XG_inst_csr_bfm:avm_write -> XG_inst:csr_write
	wire         xg_inst_avalon_st_rx_valid;                  // XG_inst:avalon_st_rx_valid -> XG_inst_avalon_st_rx_bfm:sink_valid
	wire  [63:0] xg_inst_avalon_st_rx_data;                   // XG_inst:avalon_st_rx_data -> XG_inst_avalon_st_rx_bfm:sink_data
	wire         xg_inst_avalon_st_rx_ready;                  // XG_inst_avalon_st_rx_bfm:sink_ready -> XG_inst:avalon_st_rx_ready
	wire         xg_inst_avalon_st_rx_startofpacket;          // XG_inst:avalon_st_rx_startofpacket -> XG_inst_avalon_st_rx_bfm:sink_startofpacket
	wire   [5:0] xg_inst_avalon_st_rx_error;                  // XG_inst:avalon_st_rx_error -> XG_inst_avalon_st_rx_bfm:sink_error
	wire         xg_inst_avalon_st_rx_endofpacket;            // XG_inst:avalon_st_rx_endofpacket -> XG_inst_avalon_st_rx_bfm:sink_endofpacket
	wire   [2:0] xg_inst_avalon_st_rx_empty;                  // XG_inst:avalon_st_rx_empty -> XG_inst_avalon_st_rx_bfm:sink_empty
	wire         xg_inst_avalon_st_rxstatus_valid;            // XG_inst:avalon_st_rxstatus_valid -> XG_inst_avalon_st_rxstatus_bfm:sink_valid
	wire  [39:0] xg_inst_avalon_st_rxstatus_data;             // XG_inst:avalon_st_rxstatus_data -> XG_inst_avalon_st_rxstatus_bfm:sink_data
	wire   [6:0] xg_inst_avalon_st_rxstatus_error;            // XG_inst:avalon_st_rxstatus_error -> XG_inst_avalon_st_rxstatus_bfm:sink_error
	wire         xg_inst_avalon_st_txstatus_valid;            // XG_inst:avalon_st_txstatus_valid -> XG_inst_avalon_st_txstatus_bfm:sink_valid
	wire  [39:0] xg_inst_avalon_st_txstatus_data;             // XG_inst:avalon_st_txstatus_data -> XG_inst_avalon_st_txstatus_bfm:sink_data
	wire   [6:0] xg_inst_avalon_st_txstatus_error;            // XG_inst:avalon_st_txstatus_error -> XG_inst_avalon_st_txstatus_bfm:sink_error
	wire   [1:0] xg_inst_link_fault_status_xgmii_rx_data;     // XG_inst:link_fault_status_xgmii_rx_data -> XG_inst_link_fault_status_xgmii_rx_bfm:sink_data
	wire   [1:0] xg_inst_avalon_st_pause_bfm_src_data;        // XG_inst_avalon_st_pause_bfm:src_data -> XG_inst:avalon_st_pause_data
	wire   [0:0] xg_inst_avalon_st_tx_bfm_src_valid;          // XG_inst_avalon_st_tx_bfm:src_valid -> XG_inst:avalon_st_tx_valid
	wire  [63:0] xg_inst_avalon_st_tx_bfm_src_data;           // XG_inst_avalon_st_tx_bfm:src_data -> XG_inst:avalon_st_tx_data
	wire         xg_inst_avalon_st_tx_bfm_src_ready;          // XG_inst:avalon_st_tx_ready -> XG_inst_avalon_st_tx_bfm:src_ready
	wire   [0:0] xg_inst_avalon_st_tx_bfm_src_startofpacket;  // XG_inst_avalon_st_tx_bfm:src_startofpacket -> XG_inst:avalon_st_tx_startofpacket
	wire   [0:0] xg_inst_avalon_st_tx_bfm_src_endofpacket;    // XG_inst_avalon_st_tx_bfm:src_endofpacket -> XG_inst:avalon_st_tx_endofpacket
	wire   [0:0] xg_inst_avalon_st_tx_bfm_src_error;          // XG_inst_avalon_st_tx_bfm:src_error -> XG_inst:avalon_st_tx_error
	wire   [2:0] xg_inst_avalon_st_tx_bfm_src_empty;          // XG_inst_avalon_st_tx_bfm:src_empty -> XG_inst:avalon_st_tx_empty
	wire         xg_inst_csr_clk_bfm_clk_clk;                 // XG_inst_csr_clk_bfm:clk -> [XG_inst:csr_clk, XG_inst_csr_bfm:clk, XG_inst_csr_rst_n_bfm:clk]
	wire         xg_inst_rx_312_5_clk_bfm_clk_clk;            // XG_inst_rx_312_5_clk_bfm:clk -> [XG_inst:rx_312_5_clk, XG_inst_rx_rst_n_bfm:clk]
	wire         xg_inst_tx_312_5_clk_bfm_clk_clk;            // XG_inst_tx_312_5_clk_bfm:clk -> [XG_inst:tx_312_5_clk, XG_inst_tx_rst_n_bfm:clk]
	wire         xg_inst_tx_156_25_clk_bfm_clk_clk;           // XG_inst_tx_156_25_clk_bfm:clk -> [XG_inst:tx_156_25_clk, XG_inst_avalon_st_pause_bfm:clk, XG_inst_avalon_st_tx_bfm:clk, XG_inst_avalon_st_txstatus_bfm:clk, rst_controller:clk]
	wire         xg_inst_rx_156_25_clk_bfm_clk_clk;           // XG_inst_rx_156_25_clk_bfm:clk -> [XG_inst:rx_156_25_clk, XG_inst_avalon_st_rx_bfm:clk, XG_inst_avalon_st_rxstatus_bfm:clk, XG_inst_link_fault_status_xgmii_rx_bfm:clk, rst_controller_001:clk]
	wire   [3:0] xg_inst_xgmii_rx_control_bfm_conduit_export; // XG_inst_xgmii_rx_control_bfm:sig_export -> XG_inst:xgmii_rx_control
	wire  [31:0] xg_inst_xgmii_rx_data_bfm_conduit_export;    // XG_inst_xgmii_rx_data_bfm:sig_export -> XG_inst:xgmii_rx_data
	wire   [3:0] xg_inst_xgmii_tx_control_export;             // XG_inst:xgmii_tx_control -> XG_inst_xgmii_tx_control_bfm:sig_export
	wire  [31:0] xg_inst_xgmii_tx_data_export;                // XG_inst:xgmii_tx_data -> XG_inst_xgmii_tx_data_bfm:sig_export
	wire         xg_inst_csr_rst_n_bfm_reset_reset;           // XG_inst_csr_rst_n_bfm:reset -> [XG_inst:csr_rst_n, XG_inst_csr_bfm:reset]
	wire         xg_inst_rx_rst_n_bfm_reset_reset;            // XG_inst_rx_rst_n_bfm:reset -> [XG_inst:rx_rst_n, rst_controller_001:reset_in0]
	wire         xg_inst_tx_rst_n_bfm_reset_reset;            // XG_inst_tx_rst_n_bfm:reset -> [XG_inst:tx_rst_n, rst_controller:reset_in0]
	wire         rst_controller_reset_out_reset;              // rst_controller:reset_out -> [XG_inst_avalon_st_pause_bfm:reset, XG_inst_avalon_st_tx_bfm:reset, XG_inst_avalon_st_txstatus_bfm:reset]
	wire         rst_controller_001_reset_out_reset;          // rst_controller_001:reset_out -> [XG_inst_avalon_st_rx_bfm:reset, XG_inst_avalon_st_rxstatus_bfm:reset, XG_inst_link_fault_status_xgmii_rx_bfm:reset]

	XG xg_inst (
		.avalon_st_pause_data            (xg_inst_avalon_st_pause_bfm_src_data),        //   input,   width = 2,            avalon_st_pause.data
		.avalon_st_rx_data               (xg_inst_avalon_st_rx_data),                   //  output,  width = 64,               avalon_st_rx.data
		.avalon_st_rx_startofpacket      (xg_inst_avalon_st_rx_startofpacket),          //  output,   width = 1,                           .startofpacket
		.avalon_st_rx_valid              (xg_inst_avalon_st_rx_valid),                  //  output,   width = 1,                           .valid
		.avalon_st_rx_empty              (xg_inst_avalon_st_rx_empty),                  //  output,   width = 3,                           .empty
		.avalon_st_rx_error              (xg_inst_avalon_st_rx_error),                  //  output,   width = 6,                           .error
		.avalon_st_rx_ready              (xg_inst_avalon_st_rx_ready),                  //   input,   width = 1,                           .ready
		.avalon_st_rx_endofpacket        (xg_inst_avalon_st_rx_endofpacket),            //  output,   width = 1,                           .endofpacket
		.avalon_st_rxstatus_valid        (xg_inst_avalon_st_rxstatus_valid),            //  output,   width = 1,         avalon_st_rxstatus.valid
		.avalon_st_rxstatus_data         (xg_inst_avalon_st_rxstatus_data),             //  output,  width = 40,                           .data
		.avalon_st_rxstatus_error        (xg_inst_avalon_st_rxstatus_error),            //  output,   width = 7,                           .error
		.avalon_st_tx_startofpacket      (xg_inst_avalon_st_tx_bfm_src_startofpacket),  //   input,   width = 1,               avalon_st_tx.startofpacket
		.avalon_st_tx_endofpacket        (xg_inst_avalon_st_tx_bfm_src_endofpacket),    //   input,   width = 1,                           .endofpacket
		.avalon_st_tx_valid              (xg_inst_avalon_st_tx_bfm_src_valid),          //   input,   width = 1,                           .valid
		.avalon_st_tx_data               (xg_inst_avalon_st_tx_bfm_src_data),           //   input,  width = 64,                           .data
		.avalon_st_tx_empty              (xg_inst_avalon_st_tx_bfm_src_empty),          //   input,   width = 3,                           .empty
		.avalon_st_tx_error              (xg_inst_avalon_st_tx_bfm_src_error),          //   input,   width = 1,                           .error
		.avalon_st_tx_ready              (xg_inst_avalon_st_tx_bfm_src_ready),          //  output,   width = 1,                           .ready
		.avalon_st_txstatus_valid        (xg_inst_avalon_st_txstatus_valid),            //  output,   width = 1,         avalon_st_txstatus.valid
		.avalon_st_txstatus_data         (xg_inst_avalon_st_txstatus_data),             //  output,  width = 40,                           .data
		.avalon_st_txstatus_error        (xg_inst_avalon_st_txstatus_error),            //  output,   width = 7,                           .error
		.csr_read                        (xg_inst_csr_bfm_m0_read),                     //   input,   width = 1,                        csr.read
		.csr_write                       (xg_inst_csr_bfm_m0_write),                    //   input,   width = 1,                           .write
		.csr_writedata                   (xg_inst_csr_bfm_m0_writedata),                //   input,  width = 32,                           .writedata
		.csr_readdata                    (xg_inst_csr_bfm_m0_readdata),                 //  output,  width = 32,                           .readdata
		.csr_waitrequest                 (xg_inst_csr_bfm_m0_waitrequest),              //  output,   width = 1,                           .waitrequest
		.csr_address                     (xg_inst_csr_bfm_m0_address),                  //   input,  width = 10,                           .address
		.csr_clk                         (xg_inst_csr_clk_bfm_clk_clk),                 //   input,   width = 1,                    csr_clk.clk
		.csr_rst_n                       (xg_inst_csr_rst_n_bfm_reset_reset),           //   input,   width = 1,                  csr_rst_n.reset_n
		.link_fault_status_xgmii_rx_data (xg_inst_link_fault_status_xgmii_rx_data),     //  output,   width = 2, link_fault_status_xgmii_rx.data
		.rx_156_25_clk                   (xg_inst_rx_156_25_clk_bfm_clk_clk),           //   input,   width = 1,              rx_156_25_clk.clk
		.rx_312_5_clk                    (xg_inst_rx_312_5_clk_bfm_clk_clk),            //   input,   width = 1,               rx_312_5_clk.clk
		.rx_rst_n                        (xg_inst_rx_rst_n_bfm_reset_reset),            //   input,   width = 1,                   rx_rst_n.reset_n
		.tx_156_25_clk                   (xg_inst_tx_156_25_clk_bfm_clk_clk),           //   input,   width = 1,              tx_156_25_clk.clk
		.tx_312_5_clk                    (xg_inst_tx_312_5_clk_bfm_clk_clk),            //   input,   width = 1,               tx_312_5_clk.clk
		.tx_rst_n                        (xg_inst_tx_rst_n_bfm_reset_reset),            //   input,   width = 1,                   tx_rst_n.reset_n
		.xgmii_rx_control                (xg_inst_xgmii_rx_control_bfm_conduit_export), //   input,   width = 4,           xgmii_rx_control.export
		.xgmii_rx_data                   (xg_inst_xgmii_rx_data_bfm_conduit_export),    //   input,  width = 32,              xgmii_rx_data.export
		.xgmii_tx_control                (xg_inst_xgmii_tx_control_export),             //  output,   width = 4,           xgmii_tx_control.export
		.xgmii_tx_data                   (xg_inst_xgmii_tx_data_export)                 //  output,  width = 32,              xgmii_tx_data.export
	);

	XG_inst_avalon_st_pause_bfm_ip xg_inst_avalon_st_pause_bfm (
		.clk      (xg_inst_tx_156_25_clk_bfm_clk_clk),    //   input,  width = 1,       clk.clk
		.reset    (rst_controller_reset_out_reset),       //   input,  width = 1, clk_reset.reset
		.src_data (xg_inst_avalon_st_pause_bfm_src_data)  //  output,  width = 2,       src.data
	);

	XG_inst_avalon_st_rx_bfm_ip xg_inst_avalon_st_rx_bfm (
		.clk                (xg_inst_rx_156_25_clk_bfm_clk_clk),  //   input,   width = 1,       clk.clk
		.reset              (rst_controller_001_reset_out_reset), //   input,   width = 1, clk_reset.reset
		.sink_data          (xg_inst_avalon_st_rx_data),          //   input,  width = 64,      sink.data
		.sink_valid         (xg_inst_avalon_st_rx_valid),         //   input,   width = 1,          .valid
		.sink_ready         (xg_inst_avalon_st_rx_ready),         //  output,   width = 1,          .ready
		.sink_startofpacket (xg_inst_avalon_st_rx_startofpacket), //   input,   width = 1,          .startofpacket
		.sink_endofpacket   (xg_inst_avalon_st_rx_endofpacket),   //   input,   width = 1,          .endofpacket
		.sink_empty         (xg_inst_avalon_st_rx_empty),         //   input,   width = 3,          .empty
		.sink_error         (xg_inst_avalon_st_rx_error)          //   input,   width = 6,          .error
	);

	XG_inst_avalon_st_rxstatus_bfm_ip xg_inst_avalon_st_rxstatus_bfm (
		.clk        (xg_inst_rx_156_25_clk_bfm_clk_clk),  //   input,   width = 1,       clk.clk
		.reset      (rst_controller_001_reset_out_reset), //   input,   width = 1, clk_reset.reset
		.sink_data  (xg_inst_avalon_st_rxstatus_data),    //   input,  width = 40,      sink.data
		.sink_valid (xg_inst_avalon_st_rxstatus_valid),   //   input,   width = 1,          .valid
		.sink_error (xg_inst_avalon_st_rxstatus_error)    //   input,   width = 7,          .error
	);

	XG_inst_avalon_st_tx_bfm_ip xg_inst_avalon_st_tx_bfm (
		.clk               (xg_inst_tx_156_25_clk_bfm_clk_clk),          //   input,   width = 1,       clk.clk
		.reset             (rst_controller_reset_out_reset),             //   input,   width = 1, clk_reset.reset
		.src_data          (xg_inst_avalon_st_tx_bfm_src_data),          //  output,  width = 64,       src.data
		.src_valid         (xg_inst_avalon_st_tx_bfm_src_valid),         //  output,   width = 1,          .valid
		.src_ready         (xg_inst_avalon_st_tx_bfm_src_ready),         //   input,   width = 1,          .ready
		.src_startofpacket (xg_inst_avalon_st_tx_bfm_src_startofpacket), //  output,   width = 1,          .startofpacket
		.src_endofpacket   (xg_inst_avalon_st_tx_bfm_src_endofpacket),   //  output,   width = 1,          .endofpacket
		.src_empty         (xg_inst_avalon_st_tx_bfm_src_empty),         //  output,   width = 3,          .empty
		.src_error         (xg_inst_avalon_st_tx_bfm_src_error)          //  output,   width = 1,          .error
	);

	XG_inst_avalon_st_txstatus_bfm_ip xg_inst_avalon_st_txstatus_bfm (
		.clk        (xg_inst_tx_156_25_clk_bfm_clk_clk), //   input,   width = 1,       clk.clk
		.reset      (rst_controller_reset_out_reset),    //   input,   width = 1, clk_reset.reset
		.sink_data  (xg_inst_avalon_st_txstatus_data),   //   input,  width = 40,      sink.data
		.sink_valid (xg_inst_avalon_st_txstatus_valid),  //   input,   width = 1,          .valid
		.sink_error (xg_inst_avalon_st_txstatus_error)   //   input,   width = 7,          .error
	);

	XG_inst_csr_bfm_ip xg_inst_csr_bfm (
		.clk             (xg_inst_csr_clk_bfm_clk_clk),        //   input,   width = 1,       clk.clk
		.reset           (~xg_inst_csr_rst_n_bfm_reset_reset), //   input,   width = 1, clk_reset.reset
		.avm_address     (xg_inst_csr_bfm_m0_address),         //  output,  width = 10,        m0.address
		.avm_readdata    (xg_inst_csr_bfm_m0_readdata),        //   input,  width = 32,          .readdata
		.avm_writedata   (xg_inst_csr_bfm_m0_writedata),       //  output,  width = 32,          .writedata
		.avm_waitrequest (xg_inst_csr_bfm_m0_waitrequest),     //   input,   width = 1,          .waitrequest
		.avm_write       (xg_inst_csr_bfm_m0_write),           //  output,   width = 1,          .write
		.avm_read        (xg_inst_csr_bfm_m0_read)             //  output,   width = 1,          .read
	);

	XG_inst_csr_clk_bfm_ip xg_inst_csr_clk_bfm (
		.clk (xg_inst_csr_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	XG_inst_csr_rst_n_bfm_ip xg_inst_csr_rst_n_bfm (
		.clk   (xg_inst_csr_clk_bfm_clk_clk),       //   input,  width = 1,   clk.clk
		.reset (xg_inst_csr_rst_n_bfm_reset_reset)  //  output,  width = 1, reset.reset_n
	);

	XG_inst_link_fault_status_xgmii_rx_bfm_ip xg_inst_link_fault_status_xgmii_rx_bfm (
		.clk       (xg_inst_rx_156_25_clk_bfm_clk_clk),       //   input,  width = 1,       clk.clk
		.reset     (rst_controller_001_reset_out_reset),      //   input,  width = 1, clk_reset.reset
		.sink_data (xg_inst_link_fault_status_xgmii_rx_data)  //   input,  width = 2,      sink.data
	);

	XG_inst_rx_156_25_clk_bfm_ip xg_inst_rx_156_25_clk_bfm (
		.clk (xg_inst_rx_156_25_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	XG_inst_rx_312_5_clk_bfm_ip xg_inst_rx_312_5_clk_bfm (
		.clk (xg_inst_rx_312_5_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	XG_inst_rx_rst_n_bfm_ip xg_inst_rx_rst_n_bfm (
		.clk   (xg_inst_rx_312_5_clk_bfm_clk_clk), //   input,  width = 1,   clk.clk
		.reset (xg_inst_rx_rst_n_bfm_reset_reset)  //  output,  width = 1, reset.reset_n
	);

	XG_inst_tx_156_25_clk_bfm_ip xg_inst_tx_156_25_clk_bfm (
		.clk (xg_inst_tx_156_25_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	XG_inst_tx_312_5_clk_bfm_ip xg_inst_tx_312_5_clk_bfm (
		.clk (xg_inst_tx_312_5_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	XG_inst_tx_rst_n_bfm_ip xg_inst_tx_rst_n_bfm (
		.clk   (xg_inst_tx_312_5_clk_bfm_clk_clk), //   input,  width = 1,   clk.clk
		.reset (xg_inst_tx_rst_n_bfm_reset_reset)  //  output,  width = 1, reset.reset_n
	);

	XG_inst_xgmii_rx_control_bfm_ip xg_inst_xgmii_rx_control_bfm (
		.sig_export (xg_inst_xgmii_rx_control_bfm_conduit_export)  //  output,  width = 4, conduit.export
	);

	XG_inst_xgmii_rx_data_bfm_ip xg_inst_xgmii_rx_data_bfm (
		.sig_export (xg_inst_xgmii_rx_data_bfm_conduit_export)  //  output,  width = 32, conduit.export
	);

	XG_inst_xgmii_tx_control_bfm_ip xg_inst_xgmii_tx_control_bfm (
		.sig_export (xg_inst_xgmii_tx_control_export)  //   input,  width = 4, conduit.export
	);

	XG_inst_xgmii_tx_data_bfm_ip xg_inst_xgmii_tx_data_bfm (
		.sig_export (xg_inst_xgmii_tx_data_export)  //   input,  width = 32, conduit.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~xg_inst_tx_rst_n_bfm_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (xg_inst_tx_156_25_clk_bfm_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    //  output,  width = 1, reset_out.reset
		.reset_req      (),                                  // (terminated),                       
		.reset_req_in0  (1'b0),                              // (terminated),                       
		.reset_in1      (1'b0),                              // (terminated),                       
		.reset_req_in1  (1'b0),                              // (terminated),                       
		.reset_in2      (1'b0),                              // (terminated),                       
		.reset_req_in2  (1'b0),                              // (terminated),                       
		.reset_in3      (1'b0),                              // (terminated),                       
		.reset_req_in3  (1'b0),                              // (terminated),                       
		.reset_in4      (1'b0),                              // (terminated),                       
		.reset_req_in4  (1'b0),                              // (terminated),                       
		.reset_in5      (1'b0),                              // (terminated),                       
		.reset_req_in5  (1'b0),                              // (terminated),                       
		.reset_in6      (1'b0),                              // (terminated),                       
		.reset_req_in6  (1'b0),                              // (terminated),                       
		.reset_in7      (1'b0),                              // (terminated),                       
		.reset_req_in7  (1'b0),                              // (terminated),                       
		.reset_in8      (1'b0),                              // (terminated),                       
		.reset_req_in8  (1'b0),                              // (terminated),                       
		.reset_in9      (1'b0),                              // (terminated),                       
		.reset_req_in9  (1'b0),                              // (terminated),                       
		.reset_in10     (1'b0),                              // (terminated),                       
		.reset_req_in10 (1'b0),                              // (terminated),                       
		.reset_in11     (1'b0),                              // (terminated),                       
		.reset_req_in11 (1'b0),                              // (terminated),                       
		.reset_in12     (1'b0),                              // (terminated),                       
		.reset_req_in12 (1'b0),                              // (terminated),                       
		.reset_in13     (1'b0),                              // (terminated),                       
		.reset_req_in13 (1'b0),                              // (terminated),                       
		.reset_in14     (1'b0),                              // (terminated),                       
		.reset_req_in14 (1'b0),                              // (terminated),                       
		.reset_in15     (1'b0),                              // (terminated),                       
		.reset_req_in15 (1'b0)                               // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~xg_inst_rx_rst_n_bfm_reset_reset),  //   input,  width = 1, reset_in0.reset
		.clk            (xg_inst_rx_156_25_clk_bfm_clk_clk),  //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
