// ep_g3x8_avmm256_tb.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module ep_g3x8_avmm256_tb (
	);

	wire         ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm_clk_clk;            // ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm:clk -> [ep_g3x8_avmm256_inst:reconfig_xcvr_clk_clk, ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm:clk]
	wire         dut_pcie_tb_refclk_clk;                                        // DUT_pcie_tb:refclk -> ep_g3x8_avmm256_inst:refclk_clk
	wire  [31:0] dut_pcie_tb_hip_ctrl_test_in;                                  // DUT_pcie_tb:test_in -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_ctrl_test_in
	wire         dut_pcie_tb_hip_ctrl_simu_mode_pipe;                           // DUT_pcie_tb:simu_mode_pipe -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_ctrl_simu_mode_pipe
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity4;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity4 -> DUT_pcie_tb:rxpolarity4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity5;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity5 -> DUT_pcie_tb:rxpolarity5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity2;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity2 -> DUT_pcie_tb:rxpolarity2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity3;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity3 -> DUT_pcie_tb:rxpolarity3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity0;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity0 -> DUT_pcie_tb:rxpolarity0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity1;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity1 -> DUT_pcie_tb:rxpolarity1
	wire         dut_pcie_tb_hip_pipe_rxdataskip0;                              // DUT_pcie_tb:rxdataskip0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip0
	wire         dut_pcie_tb_hip_pipe_rxdataskip2;                              // DUT_pcie_tb:rxdataskip2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip2
	wire         dut_pcie_tb_hip_pipe_rxdataskip1;                              // DUT_pcie_tb:rxdataskip1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip1
	wire         dut_pcie_tb_hip_pipe_rxdataskip4;                              // DUT_pcie_tb:rxdataskip4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip4
	wire         dut_pcie_tb_hip_pipe_rxdataskip3;                              // DUT_pcie_tb:rxdataskip3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip3
	wire         dut_pcie_tb_hip_pipe_rxdataskip6;                              // DUT_pcie_tb:rxdataskip6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip6
	wire         dut_pcie_tb_hip_pipe_rxdataskip5;                              // DUT_pcie_tb:rxdataskip5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip5
	wire         dut_pcie_tb_hip_pipe_rxdataskip7;                              // DUT_pcie_tb:rxdataskip7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdataskip7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph7;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph7 -> DUT_pcie_tb:txdeemph7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph5;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph5 -> DUT_pcie_tb:txdeemph5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph6;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph6 -> DUT_pcie_tb:txdeemph6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph0;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph0 -> DUT_pcie_tb:txdeemph0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph3;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph3 -> DUT_pcie_tb:txdeemph3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph4;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph4 -> DUT_pcie_tb:txdeemph4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph1;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph1 -> DUT_pcie_tb:txdeemph1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph2;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdeemph2 -> DUT_pcie_tb:txdeemph2
	wire         dut_pcie_tb_hip_pipe_sim_pipe_pclk_in;                         // DUT_pcie_tb:sim_pipe_pclk_in -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_sim_pipe_pclk_in
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_pipe_rate;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_sim_pipe_rate -> DUT_pcie_tb:sim_pipe_rate
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip7;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip7 -> DUT_pcie_tb:txdataskip7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip6;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip6 -> DUT_pcie_tb:txdataskip6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip5;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip5 -> DUT_pcie_tb:txdataskip5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip0;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip0 -> DUT_pcie_tb:txdataskip0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip4;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip4 -> DUT_pcie_tb:txdataskip4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip3;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip3 -> DUT_pcie_tb:txdataskip3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip2;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip2 -> DUT_pcie_tb:txdataskip2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip1;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdataskip1 -> DUT_pcie_tb:txdataskip1
	wire         dut_pcie_tb_hip_pipe_rxvalid5;                                 // DUT_pcie_tb:rxvalid5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid5
	wire         dut_pcie_tb_hip_pipe_rxvalid4;                                 // DUT_pcie_tb:rxvalid4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid4
	wire         dut_pcie_tb_hip_pipe_rxvalid3;                                 // DUT_pcie_tb:rxvalid3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid3
	wire         dut_pcie_tb_hip_pipe_rxvalid2;                                 // DUT_pcie_tb:rxvalid2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid2
	wire         dut_pcie_tb_hip_pipe_rxvalid1;                                 // DUT_pcie_tb:rxvalid1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid1
	wire         dut_pcie_tb_hip_pipe_rxvalid0;                                 // DUT_pcie_tb:rxvalid0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid0
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak2;                                 // DUT_pcie_tb:rxdatak2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak2
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak1;                                 // DUT_pcie_tb:rxdatak1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak1
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak0;                                 // DUT_pcie_tb:rxdatak0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak0
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak6;                                 // DUT_pcie_tb:rxdatak6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak6
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak5;                                 // DUT_pcie_tb:rxdatak5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak5
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak4;                                 // DUT_pcie_tb:rxdatak4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak4
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak3;                                 // DUT_pcie_tb:rxdatak3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak3
	wire   [3:0] dut_pcie_tb_hip_pipe_rxdatak7;                                 // DUT_pcie_tb:rxdatak7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdatak7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing7;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing7 -> DUT_pcie_tb:txswing7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing6;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing6 -> DUT_pcie_tb:txswing6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing5;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing5 -> DUT_pcie_tb:txswing5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing4;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing4 -> DUT_pcie_tb:txswing4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing3;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing3 -> DUT_pcie_tb:txswing3
	wire         dut_pcie_tb_hip_pipe_rxvalid7;                                 // DUT_pcie_tb:rxvalid7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing2;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing2 -> DUT_pcie_tb:txswing2
	wire         dut_pcie_tb_hip_pipe_rxvalid6;                                 // DUT_pcie_tb:rxvalid6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxvalid6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing1;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing1 -> DUT_pcie_tb:txswing1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing0;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txswing0 -> DUT_pcie_tb:txswing0
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff7;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff7 -> DUT_pcie_tb:currentcoeff7
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff6;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff6 -> DUT_pcie_tb:currentcoeff6
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff5;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff5 -> DUT_pcie_tb:currentcoeff5
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff4;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff4 -> DUT_pcie_tb:currentcoeff4
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff3;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff3 -> DUT_pcie_tb:currentcoeff3
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff2;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff2 -> DUT_pcie_tb:currentcoeff2
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff1;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff1 -> DUT_pcie_tb:currentcoeff1
	wire  [17:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff0;    // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentcoeff0 -> DUT_pcie_tb:currentcoeff0
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel5;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel5 -> DUT_pcie_tb:eidleinfersel5
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel6;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel6 -> DUT_pcie_tb:eidleinfersel6
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel7;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel7 -> DUT_pcie_tb:eidleinfersel7
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel1;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel1 -> DUT_pcie_tb:eidleinfersel1
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel2;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel2 -> DUT_pcie_tb:eidleinfersel2
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel3;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel3 -> DUT_pcie_tb:eidleinfersel3
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel4;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel4 -> DUT_pcie_tb:eidleinfersel4
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel0;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_eidleinfersel0 -> DUT_pcie_tb:eidleinfersel0
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata5;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata5 -> DUT_pcie_tb:txdata5
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata4;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata4 -> DUT_pcie_tb:txdata4
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata3;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata3 -> DUT_pcie_tb:txdata3
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata2;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata2 -> DUT_pcie_tb:txdata2
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata1;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata1 -> DUT_pcie_tb:txdata1
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata0;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata0 -> DUT_pcie_tb:txdata0
	wire         dut_pcie_tb_hip_pipe_rxelecidle7;                              // DUT_pcie_tb:rxelecidle7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle7
	wire         dut_pcie_tb_hip_pipe_rxelecidle6;                              // DUT_pcie_tb:rxelecidle6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle6
	wire         dut_pcie_tb_hip_pipe_rxelecidle5;                              // DUT_pcie_tb:rxelecidle5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle5
	wire         dut_pcie_tb_hip_pipe_rxelecidle4;                              // DUT_pcie_tb:rxelecidle4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle4
	wire         dut_pcie_tb_hip_pipe_rxelecidle3;                              // DUT_pcie_tb:rxelecidle3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle3
	wire         dut_pcie_tb_hip_pipe_rxelecidle2;                              // DUT_pcie_tb:rxelecidle2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle2
	wire         dut_pcie_tb_hip_pipe_rxelecidle1;                              // DUT_pcie_tb:rxelecidle1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle1
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata7;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata7 -> DUT_pcie_tb:txdata7
	wire         dut_pcie_tb_hip_pipe_rxelecidle0;                              // DUT_pcie_tb:rxelecidle0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxelecidle0
	wire  [31:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata6;          // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdata6 -> DUT_pcie_tb:txdata6
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd7;                                // DUT_pcie_tb:rxsynchd7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd7
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd5;                                // DUT_pcie_tb:rxsynchd5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd5
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd6;                                // DUT_pcie_tb:rxsynchd6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd6
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd0;                                // DUT_pcie_tb:rxsynchd0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd0
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd3;                                // DUT_pcie_tb:rxsynchd3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd3
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd4;                                // DUT_pcie_tb:rxsynchd4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd4
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd1;                                // DUT_pcie_tb:rxsynchd1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd1
	wire   [1:0] dut_pcie_tb_hip_pipe_rxsynchd2;                                // DUT_pcie_tb:rxsynchd2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxsynchd2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst1;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst1 -> DUT_pcie_tb:txblkst1
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate4;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate4 -> DUT_pcie_tb:rate4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst0;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst0 -> DUT_pcie_tb:txblkst0
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate5;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate5 -> DUT_pcie_tb:rate5
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate6;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate6 -> DUT_pcie_tb:rate6
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate7;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate7 -> DUT_pcie_tb:rate7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl0;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl0 -> DUT_pcie_tb:txcompl0
	wire         dut_pcie_tb_hip_pipe_rxblkst0;                                 // DUT_pcie_tb:rxblkst0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst5;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst5 -> DUT_pcie_tb:txblkst5
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate0;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate0 -> DUT_pcie_tb:rate0
	wire         dut_pcie_tb_hip_pipe_rxblkst1;                                 // DUT_pcie_tb:rxblkst1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst4;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst4 -> DUT_pcie_tb:txblkst4
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate1;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate1 -> DUT_pcie_tb:rate1
	wire         dut_pcie_tb_hip_pipe_rxblkst2;                                 // DUT_pcie_tb:rxblkst2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst3;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst3 -> DUT_pcie_tb:txblkst3
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate2;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate2 -> DUT_pcie_tb:rate2
	wire         dut_pcie_tb_hip_pipe_rxblkst3;                                 // DUT_pcie_tb:rxblkst3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst2;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst2 -> DUT_pcie_tb:txblkst2
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate3;            // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rate3 -> DUT_pcie_tb:rate3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl4;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl4 -> DUT_pcie_tb:txcompl4
	wire         dut_pcie_tb_hip_pipe_rxblkst4;                                 // DUT_pcie_tb:rxblkst4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl3;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl3 -> DUT_pcie_tb:txcompl3
	wire         dut_pcie_tb_hip_pipe_rxblkst5;                                 // DUT_pcie_tb:rxblkst5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl2;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl2 -> DUT_pcie_tb:txcompl2
	wire         dut_pcie_tb_hip_pipe_rxblkst6;                                 // DUT_pcie_tb:rxblkst6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst7;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst7 -> DUT_pcie_tb:txblkst7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl1;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl1 -> DUT_pcie_tb:txcompl1
	wire         dut_pcie_tb_hip_pipe_rxblkst7;                                 // DUT_pcie_tb:rxblkst7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxblkst7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst6;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txblkst6 -> DUT_pcie_tb:txblkst6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl7;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl7 -> DUT_pcie_tb:txcompl7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl6;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl6 -> DUT_pcie_tb:txcompl6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl5;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txcompl5 -> DUT_pcie_tb:txcompl5
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown3;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown3 -> DUT_pcie_tb:powerdown3
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown4;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown4 -> DUT_pcie_tb:powerdown4
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown5;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown5 -> DUT_pcie_tb:powerdown5
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown6;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown6 -> DUT_pcie_tb:powerdown6
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown0;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown0 -> DUT_pcie_tb:powerdown0
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown1;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown1 -> DUT_pcie_tb:powerdown1
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown2;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown2 -> DUT_pcie_tb:powerdown2
	wire   [4:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_ltssmstate;   // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_sim_ltssmstate -> DUT_pcie_tb:sim_ltssmstate
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown7;       // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_powerdown7 -> DUT_pcie_tb:powerdown7
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd2;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd2 -> DUT_pcie_tb:txsynchd2
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd1;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd1 -> DUT_pcie_tb:txsynchd1
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd0;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd0 -> DUT_pcie_tb:txsynchd0
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus2;                                // DUT_pcie_tb:rxstatus2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus2
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd6;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd6 -> DUT_pcie_tb:txsynchd6
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus3;                                // DUT_pcie_tb:rxstatus3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus3
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd5;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd5 -> DUT_pcie_tb:txsynchd5
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus0;                                // DUT_pcie_tb:rxstatus0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus0
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd4;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd4 -> DUT_pcie_tb:txsynchd4
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus1;                                // DUT_pcie_tb:rxstatus1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus1
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd3;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd3 -> DUT_pcie_tb:txsynchd3
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus6;                                // DUT_pcie_tb:rxstatus6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus6
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus7;                                // DUT_pcie_tb:rxstatus7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus7
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus4;                                // DUT_pcie_tb:rxstatus4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus4
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus5;                                // DUT_pcie_tb:rxstatus5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxstatus5
	wire   [1:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd7;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txsynchd7 -> DUT_pcie_tb:txsynchd7
	wire         dut_pcie_tb_hip_pipe_phystatus0;                               // DUT_pcie_tb:phystatus0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus0
	wire         dut_pcie_tb_hip_pipe_phystatus1;                               // DUT_pcie_tb:phystatus1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus1
	wire         dut_pcie_tb_hip_pipe_phystatus2;                               // DUT_pcie_tb:phystatus2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus2
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset7; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset7 -> DUT_pcie_tb:currentrxpreset7
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset6; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset6 -> DUT_pcie_tb:currentrxpreset6
	wire         dut_pcie_tb_hip_pipe_phystatus3;                               // DUT_pcie_tb:phystatus3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus3
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset3; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset3 -> DUT_pcie_tb:currentrxpreset3
	wire         dut_pcie_tb_hip_pipe_phystatus4;                               // DUT_pcie_tb:phystatus4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus4
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset2; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset2 -> DUT_pcie_tb:currentrxpreset2
	wire         dut_pcie_tb_hip_pipe_phystatus5;                               // DUT_pcie_tb:phystatus5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus5
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset5; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset5 -> DUT_pcie_tb:currentrxpreset5
	wire         dut_pcie_tb_hip_pipe_phystatus6;                               // DUT_pcie_tb:phystatus6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus6
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset4; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset4 -> DUT_pcie_tb:currentrxpreset4
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin1;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin1 -> DUT_pcie_tb:txmargin1
	wire         dut_pcie_tb_hip_pipe_phystatus7;                               // DUT_pcie_tb:phystatus7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_phystatus7
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin0;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin0 -> DUT_pcie_tb:txmargin0
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset1; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset1 -> DUT_pcie_tb:currentrxpreset1
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset0; // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_currentrxpreset0 -> DUT_pcie_tb:currentrxpreset0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle5;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle5 -> DUT_pcie_tb:txelecidle5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle6;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle6 -> DUT_pcie_tb:txelecidle6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle7;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle7 -> DUT_pcie_tb:txelecidle7
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata2;                                  // DUT_pcie_tb:rxdata2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata2
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata3;                                  // DUT_pcie_tb:rxdata3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata3
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata0;                                  // DUT_pcie_tb:rxdata0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle0;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle0 -> DUT_pcie_tb:txelecidle0
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata1;                                  // DUT_pcie_tb:rxdata1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle1;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle1 -> DUT_pcie_tb:txelecidle1
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata6;                                  // DUT_pcie_tb:rxdata6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle2;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle2 -> DUT_pcie_tb:txelecidle2
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata7;                                  // DUT_pcie_tb:rxdata7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle3;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle3 -> DUT_pcie_tb:txelecidle3
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata4;                                  // DUT_pcie_tb:rxdata4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle4;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txelecidle4 -> DUT_pcie_tb:txelecidle4
	wire  [31:0] dut_pcie_tb_hip_pipe_rxdata5;                                  // DUT_pcie_tb:rxdata5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxdata5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx2;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx2 -> DUT_pcie_tb:txdetectrx2
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin5;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin5 -> DUT_pcie_tb:txmargin5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx1;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx1 -> DUT_pcie_tb:txdetectrx1
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin4;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin4 -> DUT_pcie_tb:txmargin4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx4;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx4 -> DUT_pcie_tb:txdetectrx4
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin3;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin3 -> DUT_pcie_tb:txmargin3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx3;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx3 -> DUT_pcie_tb:txdetectrx3
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin2;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin2 -> DUT_pcie_tb:txmargin2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx0;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx0 -> DUT_pcie_tb:txdetectrx0
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin7;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin7 -> DUT_pcie_tb:txmargin7
	wire   [2:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin6;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txmargin6 -> DUT_pcie_tb:txmargin6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx6;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx6 -> DUT_pcie_tb:txdetectrx6
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx5;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx5 -> DUT_pcie_tb:txdetectrx5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx7;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdetectrx7 -> DUT_pcie_tb:txdetectrx7
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak2;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak2 -> DUT_pcie_tb:txdatak2
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak1;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak1 -> DUT_pcie_tb:txdatak1
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak4;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak4 -> DUT_pcie_tb:txdatak4
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak3;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak3 -> DUT_pcie_tb:txdatak3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity6;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity6 -> DUT_pcie_tb:rxpolarity6
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak0;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak0 -> DUT_pcie_tb:txdatak0
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity7;      // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_rxpolarity7 -> DUT_pcie_tb:rxpolarity7
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak6;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak6 -> DUT_pcie_tb:txdatak6
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak5;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak5 -> DUT_pcie_tb:txdatak5
	wire   [3:0] ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak7;         // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_pipe_txdatak7 -> DUT_pcie_tb:txdatak7
	wire         dut_pcie_tb_hip_serial_rx_in0;                                 // DUT_pcie_tb:rx_in0 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in0
	wire         dut_pcie_tb_hip_serial_rx_in1;                                 // DUT_pcie_tb:rx_in1 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out7;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out7 -> DUT_pcie_tb:tx_out7
	wire         dut_pcie_tb_hip_serial_rx_in2;                                 // DUT_pcie_tb:rx_in2 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out6;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out6 -> DUT_pcie_tb:tx_out6
	wire         dut_pcie_tb_hip_serial_rx_in3;                                 // DUT_pcie_tb:rx_in3 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in3
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out5;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out5 -> DUT_pcie_tb:tx_out5
	wire         dut_pcie_tb_hip_serial_rx_in4;                                 // DUT_pcie_tb:rx_in4 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in4
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out4;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out4 -> DUT_pcie_tb:tx_out4
	wire         dut_pcie_tb_hip_serial_rx_in5;                                 // DUT_pcie_tb:rx_in5 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in5
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out3;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out3 -> DUT_pcie_tb:tx_out3
	wire         dut_pcie_tb_hip_serial_rx_in6;                                 // DUT_pcie_tb:rx_in6 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in6
	wire         dut_pcie_tb_hip_serial_rx_in7;                                 // DUT_pcie_tb:rx_in7 -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_rx_in7
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out2;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out2 -> DUT_pcie_tb:tx_out2
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out1;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out1 -> DUT_pcie_tb:tx_out1
	wire         ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out0;        // ep_g3x8_avmm256_inst:pcie_a10_hip_0_hip_serial_tx_out0 -> DUT_pcie_tb:tx_out0
	wire         dut_pcie_tb_npor_npor;                                         // DUT_pcie_tb:npor -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_npor_npor
	wire         dut_pcie_tb_npor_pin_perst;                                    // DUT_pcie_tb:pin_perst -> ep_g3x8_avmm256_inst:pcie_a10_hip_0_npor_pin_perst
	wire         ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm_reset_reset;      // ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm:reset -> ep_g3x8_avmm256_inst:reconfig_xcvr_reset_reset_n
        

        initial begin
           $fsdbDumpon();
           $fsdbDumpfile("./PcieDma.fsdb");
           $fsdbDumpvars(0,ep_g3x8_avmm256_tb);
        end
	DUT_pcie_tb_ip dut_pcie_tb (
		.test_in          (dut_pcie_tb_hip_ctrl_test_in),                                  //  output,  width = 32,   hip_ctrl.test_in
		.simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),                           //  output,   width = 1,           .simu_mode_pipe
		.sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in),                         //  output,   width = 1,   hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_pipe_rate),    //   input,   width = 2,           .sim_pipe_rate
		.sim_ltssmstate   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_ltssmstate),   //   input,   width = 5,           .sim_ltssmstate
		.eidleinfersel0   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel0),   //   input,   width = 3,           .eidleinfersel0
		.eidleinfersel1   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel1),   //   input,   width = 3,           .eidleinfersel1
		.eidleinfersel2   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel2),   //   input,   width = 3,           .eidleinfersel2
		.eidleinfersel3   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel3),   //   input,   width = 3,           .eidleinfersel3
		.eidleinfersel4   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel4),   //   input,   width = 3,           .eidleinfersel4
		.eidleinfersel5   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel5),   //   input,   width = 3,           .eidleinfersel5
		.eidleinfersel6   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel6),   //   input,   width = 3,           .eidleinfersel6
		.eidleinfersel7   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel7),   //   input,   width = 3,           .eidleinfersel7
		.powerdown0       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown0),       //   input,   width = 2,           .powerdown0
		.powerdown1       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown1),       //   input,   width = 2,           .powerdown1
		.powerdown2       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown2),       //   input,   width = 2,           .powerdown2
		.powerdown3       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown3),       //   input,   width = 2,           .powerdown3
		.powerdown4       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown4),       //   input,   width = 2,           .powerdown4
		.powerdown5       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown5),       //   input,   width = 2,           .powerdown5
		.powerdown6       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown6),       //   input,   width = 2,           .powerdown6
		.powerdown7       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown7),       //   input,   width = 2,           .powerdown7
		.rxpolarity0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity0),      //   input,   width = 1,           .rxpolarity0
		.rxpolarity1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity1),      //   input,   width = 1,           .rxpolarity1
		.rxpolarity2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity2),      //   input,   width = 1,           .rxpolarity2
		.rxpolarity3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity3),      //   input,   width = 1,           .rxpolarity3
		.rxpolarity4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity4),      //   input,   width = 1,           .rxpolarity4
		.rxpolarity5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity5),      //   input,   width = 1,           .rxpolarity5
		.rxpolarity6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity6),      //   input,   width = 1,           .rxpolarity6
		.rxpolarity7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity7),      //   input,   width = 1,           .rxpolarity7
		.txcompl0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl0),         //   input,   width = 1,           .txcompl0
		.txcompl1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl1),         //   input,   width = 1,           .txcompl1
		.txcompl2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl2),         //   input,   width = 1,           .txcompl2
		.txcompl3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl3),         //   input,   width = 1,           .txcompl3
		.txcompl4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl4),         //   input,   width = 1,           .txcompl4
		.txcompl5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl5),         //   input,   width = 1,           .txcompl5
		.txcompl6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl6),         //   input,   width = 1,           .txcompl6
		.txcompl7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl7),         //   input,   width = 1,           .txcompl7
		.txdata0          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata0),          //   input,  width = 32,           .txdata0
		.txdata1          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata1),          //   input,  width = 32,           .txdata1
		.txdata2          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata2),          //   input,  width = 32,           .txdata2
		.txdata3          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata3),          //   input,  width = 32,           .txdata3
		.txdata4          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata4),          //   input,  width = 32,           .txdata4
		.txdata5          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata5),          //   input,  width = 32,           .txdata5
		.txdata6          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata6),          //   input,  width = 32,           .txdata6
		.txdata7          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata7),          //   input,  width = 32,           .txdata7
		.txdatak0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak0),         //   input,   width = 4,           .txdatak0
		.txdatak1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak1),         //   input,   width = 4,           .txdatak1
		.txdatak2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak2),         //   input,   width = 4,           .txdatak2
		.txdatak3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak3),         //   input,   width = 4,           .txdatak3
		.txdatak4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak4),         //   input,   width = 4,           .txdatak4
		.txdatak5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak5),         //   input,   width = 4,           .txdatak5
		.txdatak6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak6),         //   input,   width = 4,           .txdatak6
		.txdatak7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak7),         //   input,   width = 4,           .txdatak7
		.txdetectrx0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx0),      //   input,   width = 1,           .txdetectrx0
		.txdetectrx1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx1),      //   input,   width = 1,           .txdetectrx1
		.txdetectrx2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx2),      //   input,   width = 1,           .txdetectrx2
		.txdetectrx3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx3),      //   input,   width = 1,           .txdetectrx3
		.txdetectrx4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx4),      //   input,   width = 1,           .txdetectrx4
		.txdetectrx5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx5),      //   input,   width = 1,           .txdetectrx5
		.txdetectrx6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx6),      //   input,   width = 1,           .txdetectrx6
		.txdetectrx7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx7),      //   input,   width = 1,           .txdetectrx7
		.txelecidle0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle0),      //   input,   width = 1,           .txelecidle0
		.txelecidle1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle1),      //   input,   width = 1,           .txelecidle1
		.txelecidle2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle2),      //   input,   width = 1,           .txelecidle2
		.txelecidle3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle3),      //   input,   width = 1,           .txelecidle3
		.txelecidle4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle4),      //   input,   width = 1,           .txelecidle4
		.txelecidle5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle5),      //   input,   width = 1,           .txelecidle5
		.txelecidle6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle6),      //   input,   width = 1,           .txelecidle6
		.txelecidle7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle7),      //   input,   width = 1,           .txelecidle7
		.txdeemph0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph0),        //   input,   width = 1,           .txdeemph0
		.txdeemph1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph1),        //   input,   width = 1,           .txdeemph1
		.txdeemph2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph2),        //   input,   width = 1,           .txdeemph2
		.txdeemph3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph3),        //   input,   width = 1,           .txdeemph3
		.txdeemph4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph4),        //   input,   width = 1,           .txdeemph4
		.txdeemph5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph5),        //   input,   width = 1,           .txdeemph5
		.txdeemph6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph6),        //   input,   width = 1,           .txdeemph6
		.txdeemph7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph7),        //   input,   width = 1,           .txdeemph7
		.txmargin0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin0),        //   input,   width = 3,           .txmargin0
		.txmargin1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin1),        //   input,   width = 3,           .txmargin1
		.txmargin2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin2),        //   input,   width = 3,           .txmargin2
		.txmargin3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin3),        //   input,   width = 3,           .txmargin3
		.txmargin4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin4),        //   input,   width = 3,           .txmargin4
		.txmargin5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin5),        //   input,   width = 3,           .txmargin5
		.txmargin6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin6),        //   input,   width = 3,           .txmargin6
		.txmargin7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin7),        //   input,   width = 3,           .txmargin7
		.txswing0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing0),         //   input,   width = 1,           .txswing0
		.txswing1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing1),         //   input,   width = 1,           .txswing1
		.txswing2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing2),         //   input,   width = 1,           .txswing2
		.txswing3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing3),         //   input,   width = 1,           .txswing3
		.txswing4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing4),         //   input,   width = 1,           .txswing4
		.txswing5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing5),         //   input,   width = 1,           .txswing5
		.txswing6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing6),         //   input,   width = 1,           .txswing6
		.txswing7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing7),         //   input,   width = 1,           .txswing7
		.phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),                               //  output,   width = 1,           .phystatus0
		.phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),                               //  output,   width = 1,           .phystatus1
		.phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),                               //  output,   width = 1,           .phystatus2
		.phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),                               //  output,   width = 1,           .phystatus3
		.phystatus4       (dut_pcie_tb_hip_pipe_phystatus4),                               //  output,   width = 1,           .phystatus4
		.phystatus5       (dut_pcie_tb_hip_pipe_phystatus5),                               //  output,   width = 1,           .phystatus5
		.phystatus6       (dut_pcie_tb_hip_pipe_phystatus6),                               //  output,   width = 1,           .phystatus6
		.phystatus7       (dut_pcie_tb_hip_pipe_phystatus7),                               //  output,   width = 1,           .phystatus7
		.rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),                                  //  output,  width = 32,           .rxdata0
		.rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),                                  //  output,  width = 32,           .rxdata1
		.rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),                                  //  output,  width = 32,           .rxdata2
		.rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),                                  //  output,  width = 32,           .rxdata3
		.rxdata4          (dut_pcie_tb_hip_pipe_rxdata4),                                  //  output,  width = 32,           .rxdata4
		.rxdata5          (dut_pcie_tb_hip_pipe_rxdata5),                                  //  output,  width = 32,           .rxdata5
		.rxdata6          (dut_pcie_tb_hip_pipe_rxdata6),                                  //  output,  width = 32,           .rxdata6
		.rxdata7          (dut_pcie_tb_hip_pipe_rxdata7),                                  //  output,  width = 32,           .rxdata7
		.rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),                                 //  output,   width = 4,           .rxdatak0
		.rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),                                 //  output,   width = 4,           .rxdatak1
		.rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),                                 //  output,   width = 4,           .rxdatak2
		.rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),                                 //  output,   width = 4,           .rxdatak3
		.rxdatak4         (dut_pcie_tb_hip_pipe_rxdatak4),                                 //  output,   width = 4,           .rxdatak4
		.rxdatak5         (dut_pcie_tb_hip_pipe_rxdatak5),                                 //  output,   width = 4,           .rxdatak5
		.rxdatak6         (dut_pcie_tb_hip_pipe_rxdatak6),                                 //  output,   width = 4,           .rxdatak6
		.rxdatak7         (dut_pcie_tb_hip_pipe_rxdatak7),                                 //  output,   width = 4,           .rxdatak7
		.rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),                              //  output,   width = 1,           .rxelecidle0
		.rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),                              //  output,   width = 1,           .rxelecidle1
		.rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),                              //  output,   width = 1,           .rxelecidle2
		.rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),                              //  output,   width = 1,           .rxelecidle3
		.rxelecidle4      (dut_pcie_tb_hip_pipe_rxelecidle4),                              //  output,   width = 1,           .rxelecidle4
		.rxelecidle5      (dut_pcie_tb_hip_pipe_rxelecidle5),                              //  output,   width = 1,           .rxelecidle5
		.rxelecidle6      (dut_pcie_tb_hip_pipe_rxelecidle6),                              //  output,   width = 1,           .rxelecidle6
		.rxelecidle7      (dut_pcie_tb_hip_pipe_rxelecidle7),                              //  output,   width = 1,           .rxelecidle7
		.rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),                                //  output,   width = 3,           .rxstatus0
		.rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),                                //  output,   width = 3,           .rxstatus1
		.rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),                                //  output,   width = 3,           .rxstatus2
		.rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),                                //  output,   width = 3,           .rxstatus3
		.rxstatus4        (dut_pcie_tb_hip_pipe_rxstatus4),                                //  output,   width = 3,           .rxstatus4
		.rxstatus5        (dut_pcie_tb_hip_pipe_rxstatus5),                                //  output,   width = 3,           .rxstatus5
		.rxstatus6        (dut_pcie_tb_hip_pipe_rxstatus6),                                //  output,   width = 3,           .rxstatus6
		.rxstatus7        (dut_pcie_tb_hip_pipe_rxstatus7),                                //  output,   width = 3,           .rxstatus7
		.rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),                                 //  output,   width = 1,           .rxvalid0
		.rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),                                 //  output,   width = 1,           .rxvalid1
		.rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),                                 //  output,   width = 1,           .rxvalid2
		.rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3),                                 //  output,   width = 1,           .rxvalid3
		.rxvalid4         (dut_pcie_tb_hip_pipe_rxvalid4),                                 //  output,   width = 1,           .rxvalid4
		.rxvalid5         (dut_pcie_tb_hip_pipe_rxvalid5),                                 //  output,   width = 1,           .rxvalid5
		.rxvalid6         (dut_pcie_tb_hip_pipe_rxvalid6),                                 //  output,   width = 1,           .rxvalid6
		.rxvalid7         (dut_pcie_tb_hip_pipe_rxvalid7),                                 //  output,   width = 1,           .rxvalid7
		.rxdataskip0      (dut_pcie_tb_hip_pipe_rxdataskip0),                              //  output,   width = 1,           .rxdataskip0
		.rxdataskip1      (dut_pcie_tb_hip_pipe_rxdataskip1),                              //  output,   width = 1,           .rxdataskip1
		.rxdataskip2      (dut_pcie_tb_hip_pipe_rxdataskip2),                              //  output,   width = 1,           .rxdataskip2
		.rxdataskip3      (dut_pcie_tb_hip_pipe_rxdataskip3),                              //  output,   width = 1,           .rxdataskip3
		.rxdataskip4      (dut_pcie_tb_hip_pipe_rxdataskip4),                              //  output,   width = 1,           .rxdataskip4
		.rxdataskip5      (dut_pcie_tb_hip_pipe_rxdataskip5),                              //  output,   width = 1,           .rxdataskip5
		.rxdataskip6      (dut_pcie_tb_hip_pipe_rxdataskip6),                              //  output,   width = 1,           .rxdataskip6
		.rxdataskip7      (dut_pcie_tb_hip_pipe_rxdataskip7),                              //  output,   width = 1,           .rxdataskip7
		.rxblkst0         (dut_pcie_tb_hip_pipe_rxblkst0),                                 //  output,   width = 1,           .rxblkst0
		.rxblkst1         (dut_pcie_tb_hip_pipe_rxblkst1),                                 //  output,   width = 1,           .rxblkst1
		.rxblkst2         (dut_pcie_tb_hip_pipe_rxblkst2),                                 //  output,   width = 1,           .rxblkst2
		.rxblkst3         (dut_pcie_tb_hip_pipe_rxblkst3),                                 //  output,   width = 1,           .rxblkst3
		.rxblkst4         (dut_pcie_tb_hip_pipe_rxblkst4),                                 //  output,   width = 1,           .rxblkst4
		.rxblkst5         (dut_pcie_tb_hip_pipe_rxblkst5),                                 //  output,   width = 1,           .rxblkst5
		.rxblkst6         (dut_pcie_tb_hip_pipe_rxblkst6),                                 //  output,   width = 1,           .rxblkst6
		.rxblkst7         (dut_pcie_tb_hip_pipe_rxblkst7),                                 //  output,   width = 1,           .rxblkst7
		.rxsynchd0        (dut_pcie_tb_hip_pipe_rxsynchd0),                                //  output,   width = 2,           .rxsynchd0
		.rxsynchd1        (dut_pcie_tb_hip_pipe_rxsynchd1),                                //  output,   width = 2,           .rxsynchd1
		.rxsynchd2        (dut_pcie_tb_hip_pipe_rxsynchd2),                                //  output,   width = 2,           .rxsynchd2
		.rxsynchd3        (dut_pcie_tb_hip_pipe_rxsynchd3),                                //  output,   width = 2,           .rxsynchd3
		.rxsynchd4        (dut_pcie_tb_hip_pipe_rxsynchd4),                                //  output,   width = 2,           .rxsynchd4
		.rxsynchd5        (dut_pcie_tb_hip_pipe_rxsynchd5),                                //  output,   width = 2,           .rxsynchd5
		.rxsynchd6        (dut_pcie_tb_hip_pipe_rxsynchd6),                                //  output,   width = 2,           .rxsynchd6
		.rxsynchd7        (dut_pcie_tb_hip_pipe_rxsynchd7),                                //  output,   width = 2,           .rxsynchd7
		.currentcoeff0    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff0),    //   input,  width = 18,           .currentcoeff0
		.currentcoeff1    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff1),    //   input,  width = 18,           .currentcoeff1
		.currentcoeff2    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff2),    //   input,  width = 18,           .currentcoeff2
		.currentcoeff3    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff3),    //   input,  width = 18,           .currentcoeff3
		.currentcoeff4    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff4),    //   input,  width = 18,           .currentcoeff4
		.currentcoeff5    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff5),    //   input,  width = 18,           .currentcoeff5
		.currentcoeff6    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff6),    //   input,  width = 18,           .currentcoeff6
		.currentcoeff7    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff7),    //   input,  width = 18,           .currentcoeff7
		.currentrxpreset0 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset0), //   input,   width = 3,           .currentrxpreset0
		.currentrxpreset1 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset1), //   input,   width = 3,           .currentrxpreset1
		.currentrxpreset2 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset2), //   input,   width = 3,           .currentrxpreset2
		.currentrxpreset3 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset3), //   input,   width = 3,           .currentrxpreset3
		.currentrxpreset4 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset4), //   input,   width = 3,           .currentrxpreset4
		.currentrxpreset5 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset5), //   input,   width = 3,           .currentrxpreset5
		.currentrxpreset6 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset6), //   input,   width = 3,           .currentrxpreset6
		.currentrxpreset7 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset7), //   input,   width = 3,           .currentrxpreset7
		.txsynchd0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd0),        //   input,   width = 2,           .txsynchd0
		.txsynchd1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd1),        //   input,   width = 2,           .txsynchd1
		.txsynchd2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd2),        //   input,   width = 2,           .txsynchd2
		.txsynchd3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd3),        //   input,   width = 2,           .txsynchd3
		.txsynchd4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd4),        //   input,   width = 2,           .txsynchd4
		.txsynchd5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd5),        //   input,   width = 2,           .txsynchd5
		.txsynchd6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd6),        //   input,   width = 2,           .txsynchd6
		.txsynchd7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd7),        //   input,   width = 2,           .txsynchd7
		.txblkst0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst0),         //   input,   width = 1,           .txblkst0
		.txblkst1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst1),         //   input,   width = 1,           .txblkst1
		.txblkst2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst2),         //   input,   width = 1,           .txblkst2
		.txblkst3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst3),         //   input,   width = 1,           .txblkst3
		.txblkst4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst4),         //   input,   width = 1,           .txblkst4
		.txblkst5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst5),         //   input,   width = 1,           .txblkst5
		.txblkst6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst6),         //   input,   width = 1,           .txblkst6
		.txblkst7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst7),         //   input,   width = 1,           .txblkst7
		.txdataskip0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip0),      //   input,   width = 1,           .txdataskip0
		.txdataskip1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip1),      //   input,   width = 1,           .txdataskip1
		.txdataskip2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip2),      //   input,   width = 1,           .txdataskip2
		.txdataskip3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip3),      //   input,   width = 1,           .txdataskip3
		.txdataskip4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip4),      //   input,   width = 1,           .txdataskip4
		.txdataskip5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip5),      //   input,   width = 1,           .txdataskip5
		.txdataskip6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip6),      //   input,   width = 1,           .txdataskip6
		.txdataskip7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip7),      //   input,   width = 1,           .txdataskip7
		.rate0            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate0),            //   input,   width = 2,           .rate0
		.rate1            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate1),            //   input,   width = 2,           .rate1
		.rate2            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate2),            //   input,   width = 2,           .rate2
		.rate3            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate3),            //   input,   width = 2,           .rate3
		.rate4            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate4),            //   input,   width = 2,           .rate4
		.rate5            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate5),            //   input,   width = 2,           .rate5
		.rate6            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate6),            //   input,   width = 2,           .rate6
		.rate7            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate7),            //   input,   width = 2,           .rate7
		.rx_in0           (dut_pcie_tb_hip_serial_rx_in0),                                 //  output,   width = 1, hip_serial.rx_in0
		.rx_in1           (dut_pcie_tb_hip_serial_rx_in1),                                 //  output,   width = 1,           .rx_in1
		.rx_in2           (dut_pcie_tb_hip_serial_rx_in2),                                 //  output,   width = 1,           .rx_in2
		.rx_in3           (dut_pcie_tb_hip_serial_rx_in3),                                 //  output,   width = 1,           .rx_in3
		.rx_in4           (dut_pcie_tb_hip_serial_rx_in4),                                 //  output,   width = 1,           .rx_in4
		.rx_in5           (dut_pcie_tb_hip_serial_rx_in5),                                 //  output,   width = 1,           .rx_in5
		.rx_in6           (dut_pcie_tb_hip_serial_rx_in6),                                 //  output,   width = 1,           .rx_in6
		.rx_in7           (dut_pcie_tb_hip_serial_rx_in7),                                 //  output,   width = 1,           .rx_in7
		.tx_out0          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out0),        //   input,   width = 1,           .tx_out0
		.tx_out1          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out1),        //   input,   width = 1,           .tx_out1
		.tx_out2          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out2),        //   input,   width = 1,           .tx_out2
		.tx_out3          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out3),        //   input,   width = 1,           .tx_out3
		.tx_out4          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out4),        //   input,   width = 1,           .tx_out4
		.tx_out5          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out5),        //   input,   width = 1,           .tx_out5
		.tx_out6          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out6),        //   input,   width = 1,           .tx_out6
		.tx_out7          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out7),        //   input,   width = 1,           .tx_out7
		.npor             (dut_pcie_tb_npor_npor),                                         //  output,   width = 1,       npor.npor
		.pin_perst        (dut_pcie_tb_npor_pin_perst),                                    //  output,   width = 1,           .pin_perst
		.refclk           (dut_pcie_tb_refclk_clk)                                         //  output,   width = 1,     refclk.clk
	);

	ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm_ip ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm (
		.clk (ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm_ip ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm (
		.clk   (ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm_clk_clk),       //   input,  width = 1,   clk.clk
		.reset (ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm_reset_reset)  //  output,  width = 1, reset.reset_n
	);

	ep_g3x8_avmm256 ep_g3x8_avmm256_inst (
		.pcie_a10_hip_0_hip_ctrl_test_in          (dut_pcie_tb_hip_ctrl_test_in),                                  //   input,  width = 32,   pcie_a10_hip_0_hip_ctrl.test_in
		.pcie_a10_hip_0_hip_ctrl_simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),                           //   input,   width = 1,                          .simu_mode_pipe
		.pcie_a10_hip_0_hip_pipe_sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in),                         //   input,   width = 1,   pcie_a10_hip_0_hip_pipe.sim_pipe_pclk_in
		.pcie_a10_hip_0_hip_pipe_sim_pipe_rate    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_pipe_rate),    //  output,   width = 2,                          .sim_pipe_rate
		.pcie_a10_hip_0_hip_pipe_sim_ltssmstate   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_sim_ltssmstate),   //  output,   width = 5,                          .sim_ltssmstate
		.pcie_a10_hip_0_hip_pipe_eidleinfersel0   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel0),   //  output,   width = 3,                          .eidleinfersel0
		.pcie_a10_hip_0_hip_pipe_eidleinfersel1   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel1),   //  output,   width = 3,                          .eidleinfersel1
		.pcie_a10_hip_0_hip_pipe_eidleinfersel2   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel2),   //  output,   width = 3,                          .eidleinfersel2
		.pcie_a10_hip_0_hip_pipe_eidleinfersel3   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel3),   //  output,   width = 3,                          .eidleinfersel3
		.pcie_a10_hip_0_hip_pipe_eidleinfersel4   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel4),   //  output,   width = 3,                          .eidleinfersel4
		.pcie_a10_hip_0_hip_pipe_eidleinfersel5   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel5),   //  output,   width = 3,                          .eidleinfersel5
		.pcie_a10_hip_0_hip_pipe_eidleinfersel6   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel6),   //  output,   width = 3,                          .eidleinfersel6
		.pcie_a10_hip_0_hip_pipe_eidleinfersel7   (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_eidleinfersel7),   //  output,   width = 3,                          .eidleinfersel7
		.pcie_a10_hip_0_hip_pipe_powerdown0       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown0),       //  output,   width = 2,                          .powerdown0
		.pcie_a10_hip_0_hip_pipe_powerdown1       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown1),       //  output,   width = 2,                          .powerdown1
		.pcie_a10_hip_0_hip_pipe_powerdown2       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown2),       //  output,   width = 2,                          .powerdown2
		.pcie_a10_hip_0_hip_pipe_powerdown3       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown3),       //  output,   width = 2,                          .powerdown3
		.pcie_a10_hip_0_hip_pipe_powerdown4       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown4),       //  output,   width = 2,                          .powerdown4
		.pcie_a10_hip_0_hip_pipe_powerdown5       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown5),       //  output,   width = 2,                          .powerdown5
		.pcie_a10_hip_0_hip_pipe_powerdown6       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown6),       //  output,   width = 2,                          .powerdown6
		.pcie_a10_hip_0_hip_pipe_powerdown7       (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_powerdown7),       //  output,   width = 2,                          .powerdown7
		.pcie_a10_hip_0_hip_pipe_rxpolarity0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity0),      //  output,   width = 1,                          .rxpolarity0
		.pcie_a10_hip_0_hip_pipe_rxpolarity1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity1),      //  output,   width = 1,                          .rxpolarity1
		.pcie_a10_hip_0_hip_pipe_rxpolarity2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity2),      //  output,   width = 1,                          .rxpolarity2
		.pcie_a10_hip_0_hip_pipe_rxpolarity3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity3),      //  output,   width = 1,                          .rxpolarity3
		.pcie_a10_hip_0_hip_pipe_rxpolarity4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity4),      //  output,   width = 1,                          .rxpolarity4
		.pcie_a10_hip_0_hip_pipe_rxpolarity5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity5),      //  output,   width = 1,                          .rxpolarity5
		.pcie_a10_hip_0_hip_pipe_rxpolarity6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity6),      //  output,   width = 1,                          .rxpolarity6
		.pcie_a10_hip_0_hip_pipe_rxpolarity7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rxpolarity7),      //  output,   width = 1,                          .rxpolarity7
		.pcie_a10_hip_0_hip_pipe_txcompl0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl0),         //  output,   width = 1,                          .txcompl0
		.pcie_a10_hip_0_hip_pipe_txcompl1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl1),         //  output,   width = 1,                          .txcompl1
		.pcie_a10_hip_0_hip_pipe_txcompl2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl2),         //  output,   width = 1,                          .txcompl2
		.pcie_a10_hip_0_hip_pipe_txcompl3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl3),         //  output,   width = 1,                          .txcompl3
		.pcie_a10_hip_0_hip_pipe_txcompl4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl4),         //  output,   width = 1,                          .txcompl4
		.pcie_a10_hip_0_hip_pipe_txcompl5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl5),         //  output,   width = 1,                          .txcompl5
		.pcie_a10_hip_0_hip_pipe_txcompl6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl6),         //  output,   width = 1,                          .txcompl6
		.pcie_a10_hip_0_hip_pipe_txcompl7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txcompl7),         //  output,   width = 1,                          .txcompl7
		.pcie_a10_hip_0_hip_pipe_txdata0          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata0),          //  output,  width = 32,                          .txdata0
		.pcie_a10_hip_0_hip_pipe_txdata1          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata1),          //  output,  width = 32,                          .txdata1
		.pcie_a10_hip_0_hip_pipe_txdata2          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata2),          //  output,  width = 32,                          .txdata2
		.pcie_a10_hip_0_hip_pipe_txdata3          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata3),          //  output,  width = 32,                          .txdata3
		.pcie_a10_hip_0_hip_pipe_txdata4          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata4),          //  output,  width = 32,                          .txdata4
		.pcie_a10_hip_0_hip_pipe_txdata5          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata5),          //  output,  width = 32,                          .txdata5
		.pcie_a10_hip_0_hip_pipe_txdata6          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata6),          //  output,  width = 32,                          .txdata6
		.pcie_a10_hip_0_hip_pipe_txdata7          (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdata7),          //  output,  width = 32,                          .txdata7
		.pcie_a10_hip_0_hip_pipe_txdatak0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak0),         //  output,   width = 4,                          .txdatak0
		.pcie_a10_hip_0_hip_pipe_txdatak1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak1),         //  output,   width = 4,                          .txdatak1
		.pcie_a10_hip_0_hip_pipe_txdatak2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak2),         //  output,   width = 4,                          .txdatak2
		.pcie_a10_hip_0_hip_pipe_txdatak3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak3),         //  output,   width = 4,                          .txdatak3
		.pcie_a10_hip_0_hip_pipe_txdatak4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak4),         //  output,   width = 4,                          .txdatak4
		.pcie_a10_hip_0_hip_pipe_txdatak5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak5),         //  output,   width = 4,                          .txdatak5
		.pcie_a10_hip_0_hip_pipe_txdatak6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak6),         //  output,   width = 4,                          .txdatak6
		.pcie_a10_hip_0_hip_pipe_txdatak7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdatak7),         //  output,   width = 4,                          .txdatak7
		.pcie_a10_hip_0_hip_pipe_txdetectrx0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx0),      //  output,   width = 1,                          .txdetectrx0
		.pcie_a10_hip_0_hip_pipe_txdetectrx1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx1),      //  output,   width = 1,                          .txdetectrx1
		.pcie_a10_hip_0_hip_pipe_txdetectrx2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx2),      //  output,   width = 1,                          .txdetectrx2
		.pcie_a10_hip_0_hip_pipe_txdetectrx3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx3),      //  output,   width = 1,                          .txdetectrx3
		.pcie_a10_hip_0_hip_pipe_txdetectrx4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx4),      //  output,   width = 1,                          .txdetectrx4
		.pcie_a10_hip_0_hip_pipe_txdetectrx5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx5),      //  output,   width = 1,                          .txdetectrx5
		.pcie_a10_hip_0_hip_pipe_txdetectrx6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx6),      //  output,   width = 1,                          .txdetectrx6
		.pcie_a10_hip_0_hip_pipe_txdetectrx7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdetectrx7),      //  output,   width = 1,                          .txdetectrx7
		.pcie_a10_hip_0_hip_pipe_txelecidle0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle0),      //  output,   width = 1,                          .txelecidle0
		.pcie_a10_hip_0_hip_pipe_txelecidle1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle1),      //  output,   width = 1,                          .txelecidle1
		.pcie_a10_hip_0_hip_pipe_txelecidle2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle2),      //  output,   width = 1,                          .txelecidle2
		.pcie_a10_hip_0_hip_pipe_txelecidle3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle3),      //  output,   width = 1,                          .txelecidle3
		.pcie_a10_hip_0_hip_pipe_txelecidle4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle4),      //  output,   width = 1,                          .txelecidle4
		.pcie_a10_hip_0_hip_pipe_txelecidle5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle5),      //  output,   width = 1,                          .txelecidle5
		.pcie_a10_hip_0_hip_pipe_txelecidle6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle6),      //  output,   width = 1,                          .txelecidle6
		.pcie_a10_hip_0_hip_pipe_txelecidle7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txelecidle7),      //  output,   width = 1,                          .txelecidle7
		.pcie_a10_hip_0_hip_pipe_txdeemph0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph0),        //  output,   width = 1,                          .txdeemph0
		.pcie_a10_hip_0_hip_pipe_txdeemph1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph1),        //  output,   width = 1,                          .txdeemph1
		.pcie_a10_hip_0_hip_pipe_txdeemph2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph2),        //  output,   width = 1,                          .txdeemph2
		.pcie_a10_hip_0_hip_pipe_txdeemph3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph3),        //  output,   width = 1,                          .txdeemph3
		.pcie_a10_hip_0_hip_pipe_txdeemph4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph4),        //  output,   width = 1,                          .txdeemph4
		.pcie_a10_hip_0_hip_pipe_txdeemph5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph5),        //  output,   width = 1,                          .txdeemph5
		.pcie_a10_hip_0_hip_pipe_txdeemph6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph6),        //  output,   width = 1,                          .txdeemph6
		.pcie_a10_hip_0_hip_pipe_txdeemph7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdeemph7),        //  output,   width = 1,                          .txdeemph7
		.pcie_a10_hip_0_hip_pipe_txmargin0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin0),        //  output,   width = 3,                          .txmargin0
		.pcie_a10_hip_0_hip_pipe_txmargin1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin1),        //  output,   width = 3,                          .txmargin1
		.pcie_a10_hip_0_hip_pipe_txmargin2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin2),        //  output,   width = 3,                          .txmargin2
		.pcie_a10_hip_0_hip_pipe_txmargin3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin3),        //  output,   width = 3,                          .txmargin3
		.pcie_a10_hip_0_hip_pipe_txmargin4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin4),        //  output,   width = 3,                          .txmargin4
		.pcie_a10_hip_0_hip_pipe_txmargin5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin5),        //  output,   width = 3,                          .txmargin5
		.pcie_a10_hip_0_hip_pipe_txmargin6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin6),        //  output,   width = 3,                          .txmargin6
		.pcie_a10_hip_0_hip_pipe_txmargin7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txmargin7),        //  output,   width = 3,                          .txmargin7
		.pcie_a10_hip_0_hip_pipe_txswing0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing0),         //  output,   width = 1,                          .txswing0
		.pcie_a10_hip_0_hip_pipe_txswing1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing1),         //  output,   width = 1,                          .txswing1
		.pcie_a10_hip_0_hip_pipe_txswing2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing2),         //  output,   width = 1,                          .txswing2
		.pcie_a10_hip_0_hip_pipe_txswing3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing3),         //  output,   width = 1,                          .txswing3
		.pcie_a10_hip_0_hip_pipe_txswing4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing4),         //  output,   width = 1,                          .txswing4
		.pcie_a10_hip_0_hip_pipe_txswing5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing5),         //  output,   width = 1,                          .txswing5
		.pcie_a10_hip_0_hip_pipe_txswing6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing6),         //  output,   width = 1,                          .txswing6
		.pcie_a10_hip_0_hip_pipe_txswing7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txswing7),         //  output,   width = 1,                          .txswing7
		.pcie_a10_hip_0_hip_pipe_phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),                               //   input,   width = 1,                          .phystatus0
		.pcie_a10_hip_0_hip_pipe_phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),                               //   input,   width = 1,                          .phystatus1
		.pcie_a10_hip_0_hip_pipe_phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),                               //   input,   width = 1,                          .phystatus2
		.pcie_a10_hip_0_hip_pipe_phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),                               //   input,   width = 1,                          .phystatus3
		.pcie_a10_hip_0_hip_pipe_phystatus4       (dut_pcie_tb_hip_pipe_phystatus4),                               //   input,   width = 1,                          .phystatus4
		.pcie_a10_hip_0_hip_pipe_phystatus5       (dut_pcie_tb_hip_pipe_phystatus5),                               //   input,   width = 1,                          .phystatus5
		.pcie_a10_hip_0_hip_pipe_phystatus6       (dut_pcie_tb_hip_pipe_phystatus6),                               //   input,   width = 1,                          .phystatus6
		.pcie_a10_hip_0_hip_pipe_phystatus7       (dut_pcie_tb_hip_pipe_phystatus7),                               //   input,   width = 1,                          .phystatus7
		.pcie_a10_hip_0_hip_pipe_rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),                                  //   input,  width = 32,                          .rxdata0
		.pcie_a10_hip_0_hip_pipe_rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),                                  //   input,  width = 32,                          .rxdata1
		.pcie_a10_hip_0_hip_pipe_rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),                                  //   input,  width = 32,                          .rxdata2
		.pcie_a10_hip_0_hip_pipe_rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),                                  //   input,  width = 32,                          .rxdata3
		.pcie_a10_hip_0_hip_pipe_rxdata4          (dut_pcie_tb_hip_pipe_rxdata4),                                  //   input,  width = 32,                          .rxdata4
		.pcie_a10_hip_0_hip_pipe_rxdata5          (dut_pcie_tb_hip_pipe_rxdata5),                                  //   input,  width = 32,                          .rxdata5
		.pcie_a10_hip_0_hip_pipe_rxdata6          (dut_pcie_tb_hip_pipe_rxdata6),                                  //   input,  width = 32,                          .rxdata6
		.pcie_a10_hip_0_hip_pipe_rxdata7          (dut_pcie_tb_hip_pipe_rxdata7),                                  //   input,  width = 32,                          .rxdata7
		.pcie_a10_hip_0_hip_pipe_rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),                                 //   input,   width = 4,                          .rxdatak0
		.pcie_a10_hip_0_hip_pipe_rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),                                 //   input,   width = 4,                          .rxdatak1
		.pcie_a10_hip_0_hip_pipe_rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),                                 //   input,   width = 4,                          .rxdatak2
		.pcie_a10_hip_0_hip_pipe_rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),                                 //   input,   width = 4,                          .rxdatak3
		.pcie_a10_hip_0_hip_pipe_rxdatak4         (dut_pcie_tb_hip_pipe_rxdatak4),                                 //   input,   width = 4,                          .rxdatak4
		.pcie_a10_hip_0_hip_pipe_rxdatak5         (dut_pcie_tb_hip_pipe_rxdatak5),                                 //   input,   width = 4,                          .rxdatak5
		.pcie_a10_hip_0_hip_pipe_rxdatak6         (dut_pcie_tb_hip_pipe_rxdatak6),                                 //   input,   width = 4,                          .rxdatak6
		.pcie_a10_hip_0_hip_pipe_rxdatak7         (dut_pcie_tb_hip_pipe_rxdatak7),                                 //   input,   width = 4,                          .rxdatak7
		.pcie_a10_hip_0_hip_pipe_rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),                              //   input,   width = 1,                          .rxelecidle0
		.pcie_a10_hip_0_hip_pipe_rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),                              //   input,   width = 1,                          .rxelecidle1
		.pcie_a10_hip_0_hip_pipe_rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),                              //   input,   width = 1,                          .rxelecidle2
		.pcie_a10_hip_0_hip_pipe_rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),                              //   input,   width = 1,                          .rxelecidle3
		.pcie_a10_hip_0_hip_pipe_rxelecidle4      (dut_pcie_tb_hip_pipe_rxelecidle4),                              //   input,   width = 1,                          .rxelecidle4
		.pcie_a10_hip_0_hip_pipe_rxelecidle5      (dut_pcie_tb_hip_pipe_rxelecidle5),                              //   input,   width = 1,                          .rxelecidle5
		.pcie_a10_hip_0_hip_pipe_rxelecidle6      (dut_pcie_tb_hip_pipe_rxelecidle6),                              //   input,   width = 1,                          .rxelecidle6
		.pcie_a10_hip_0_hip_pipe_rxelecidle7      (dut_pcie_tb_hip_pipe_rxelecidle7),                              //   input,   width = 1,                          .rxelecidle7
		.pcie_a10_hip_0_hip_pipe_rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),                                //   input,   width = 3,                          .rxstatus0
		.pcie_a10_hip_0_hip_pipe_rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),                                //   input,   width = 3,                          .rxstatus1
		.pcie_a10_hip_0_hip_pipe_rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),                                //   input,   width = 3,                          .rxstatus2
		.pcie_a10_hip_0_hip_pipe_rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),                                //   input,   width = 3,                          .rxstatus3
		.pcie_a10_hip_0_hip_pipe_rxstatus4        (dut_pcie_tb_hip_pipe_rxstatus4),                                //   input,   width = 3,                          .rxstatus4
		.pcie_a10_hip_0_hip_pipe_rxstatus5        (dut_pcie_tb_hip_pipe_rxstatus5),                                //   input,   width = 3,                          .rxstatus5
		.pcie_a10_hip_0_hip_pipe_rxstatus6        (dut_pcie_tb_hip_pipe_rxstatus6),                                //   input,   width = 3,                          .rxstatus6
		.pcie_a10_hip_0_hip_pipe_rxstatus7        (dut_pcie_tb_hip_pipe_rxstatus7),                                //   input,   width = 3,                          .rxstatus7
		.pcie_a10_hip_0_hip_pipe_rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),                                 //   input,   width = 1,                          .rxvalid0
		.pcie_a10_hip_0_hip_pipe_rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),                                 //   input,   width = 1,                          .rxvalid1
		.pcie_a10_hip_0_hip_pipe_rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),                                 //   input,   width = 1,                          .rxvalid2
		.pcie_a10_hip_0_hip_pipe_rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3),                                 //   input,   width = 1,                          .rxvalid3
		.pcie_a10_hip_0_hip_pipe_rxvalid4         (dut_pcie_tb_hip_pipe_rxvalid4),                                 //   input,   width = 1,                          .rxvalid4
		.pcie_a10_hip_0_hip_pipe_rxvalid5         (dut_pcie_tb_hip_pipe_rxvalid5),                                 //   input,   width = 1,                          .rxvalid5
		.pcie_a10_hip_0_hip_pipe_rxvalid6         (dut_pcie_tb_hip_pipe_rxvalid6),                                 //   input,   width = 1,                          .rxvalid6
		.pcie_a10_hip_0_hip_pipe_rxvalid7         (dut_pcie_tb_hip_pipe_rxvalid7),                                 //   input,   width = 1,                          .rxvalid7
		.pcie_a10_hip_0_hip_pipe_rxdataskip0      (dut_pcie_tb_hip_pipe_rxdataskip0),                              //   input,   width = 1,                          .rxdataskip0
		.pcie_a10_hip_0_hip_pipe_rxdataskip1      (dut_pcie_tb_hip_pipe_rxdataskip1),                              //   input,   width = 1,                          .rxdataskip1
		.pcie_a10_hip_0_hip_pipe_rxdataskip2      (dut_pcie_tb_hip_pipe_rxdataskip2),                              //   input,   width = 1,                          .rxdataskip2
		.pcie_a10_hip_0_hip_pipe_rxdataskip3      (dut_pcie_tb_hip_pipe_rxdataskip3),                              //   input,   width = 1,                          .rxdataskip3
		.pcie_a10_hip_0_hip_pipe_rxdataskip4      (dut_pcie_tb_hip_pipe_rxdataskip4),                              //   input,   width = 1,                          .rxdataskip4
		.pcie_a10_hip_0_hip_pipe_rxdataskip5      (dut_pcie_tb_hip_pipe_rxdataskip5),                              //   input,   width = 1,                          .rxdataskip5
		.pcie_a10_hip_0_hip_pipe_rxdataskip6      (dut_pcie_tb_hip_pipe_rxdataskip6),                              //   input,   width = 1,                          .rxdataskip6
		.pcie_a10_hip_0_hip_pipe_rxdataskip7      (dut_pcie_tb_hip_pipe_rxdataskip7),                              //   input,   width = 1,                          .rxdataskip7
		.pcie_a10_hip_0_hip_pipe_rxblkst0         (dut_pcie_tb_hip_pipe_rxblkst0),                                 //   input,   width = 1,                          .rxblkst0
		.pcie_a10_hip_0_hip_pipe_rxblkst1         (dut_pcie_tb_hip_pipe_rxblkst1),                                 //   input,   width = 1,                          .rxblkst1
		.pcie_a10_hip_0_hip_pipe_rxblkst2         (dut_pcie_tb_hip_pipe_rxblkst2),                                 //   input,   width = 1,                          .rxblkst2
		.pcie_a10_hip_0_hip_pipe_rxblkst3         (dut_pcie_tb_hip_pipe_rxblkst3),                                 //   input,   width = 1,                          .rxblkst3
		.pcie_a10_hip_0_hip_pipe_rxblkst4         (dut_pcie_tb_hip_pipe_rxblkst4),                                 //   input,   width = 1,                          .rxblkst4
		.pcie_a10_hip_0_hip_pipe_rxblkst5         (dut_pcie_tb_hip_pipe_rxblkst5),                                 //   input,   width = 1,                          .rxblkst5
		.pcie_a10_hip_0_hip_pipe_rxblkst6         (dut_pcie_tb_hip_pipe_rxblkst6),                                 //   input,   width = 1,                          .rxblkst6
		.pcie_a10_hip_0_hip_pipe_rxblkst7         (dut_pcie_tb_hip_pipe_rxblkst7),                                 //   input,   width = 1,                          .rxblkst7
		.pcie_a10_hip_0_hip_pipe_rxsynchd0        (dut_pcie_tb_hip_pipe_rxsynchd0),                                //   input,   width = 2,                          .rxsynchd0
		.pcie_a10_hip_0_hip_pipe_rxsynchd1        (dut_pcie_tb_hip_pipe_rxsynchd1),                                //   input,   width = 2,                          .rxsynchd1
		.pcie_a10_hip_0_hip_pipe_rxsynchd2        (dut_pcie_tb_hip_pipe_rxsynchd2),                                //   input,   width = 2,                          .rxsynchd2
		.pcie_a10_hip_0_hip_pipe_rxsynchd3        (dut_pcie_tb_hip_pipe_rxsynchd3),                                //   input,   width = 2,                          .rxsynchd3
		.pcie_a10_hip_0_hip_pipe_rxsynchd4        (dut_pcie_tb_hip_pipe_rxsynchd4),                                //   input,   width = 2,                          .rxsynchd4
		.pcie_a10_hip_0_hip_pipe_rxsynchd5        (dut_pcie_tb_hip_pipe_rxsynchd5),                                //   input,   width = 2,                          .rxsynchd5
		.pcie_a10_hip_0_hip_pipe_rxsynchd6        (dut_pcie_tb_hip_pipe_rxsynchd6),                                //   input,   width = 2,                          .rxsynchd6
		.pcie_a10_hip_0_hip_pipe_rxsynchd7        (dut_pcie_tb_hip_pipe_rxsynchd7),                                //   input,   width = 2,                          .rxsynchd7
		.pcie_a10_hip_0_hip_pipe_currentcoeff0    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff0),    //  output,  width = 18,                          .currentcoeff0
		.pcie_a10_hip_0_hip_pipe_currentcoeff1    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff1),    //  output,  width = 18,                          .currentcoeff1
		.pcie_a10_hip_0_hip_pipe_currentcoeff2    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff2),    //  output,  width = 18,                          .currentcoeff2
		.pcie_a10_hip_0_hip_pipe_currentcoeff3    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff3),    //  output,  width = 18,                          .currentcoeff3
		.pcie_a10_hip_0_hip_pipe_currentcoeff4    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff4),    //  output,  width = 18,                          .currentcoeff4
		.pcie_a10_hip_0_hip_pipe_currentcoeff5    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff5),    //  output,  width = 18,                          .currentcoeff5
		.pcie_a10_hip_0_hip_pipe_currentcoeff6    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff6),    //  output,  width = 18,                          .currentcoeff6
		.pcie_a10_hip_0_hip_pipe_currentcoeff7    (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentcoeff7),    //  output,  width = 18,                          .currentcoeff7
		.pcie_a10_hip_0_hip_pipe_currentrxpreset0 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset0), //  output,   width = 3,                          .currentrxpreset0
		.pcie_a10_hip_0_hip_pipe_currentrxpreset1 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset1), //  output,   width = 3,                          .currentrxpreset1
		.pcie_a10_hip_0_hip_pipe_currentrxpreset2 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset2), //  output,   width = 3,                          .currentrxpreset2
		.pcie_a10_hip_0_hip_pipe_currentrxpreset3 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset3), //  output,   width = 3,                          .currentrxpreset3
		.pcie_a10_hip_0_hip_pipe_currentrxpreset4 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset4), //  output,   width = 3,                          .currentrxpreset4
		.pcie_a10_hip_0_hip_pipe_currentrxpreset5 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset5), //  output,   width = 3,                          .currentrxpreset5
		.pcie_a10_hip_0_hip_pipe_currentrxpreset6 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset6), //  output,   width = 3,                          .currentrxpreset6
		.pcie_a10_hip_0_hip_pipe_currentrxpreset7 (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_currentrxpreset7), //  output,   width = 3,                          .currentrxpreset7
		.pcie_a10_hip_0_hip_pipe_txsynchd0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd0),        //  output,   width = 2,                          .txsynchd0
		.pcie_a10_hip_0_hip_pipe_txsynchd1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd1),        //  output,   width = 2,                          .txsynchd1
		.pcie_a10_hip_0_hip_pipe_txsynchd2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd2),        //  output,   width = 2,                          .txsynchd2
		.pcie_a10_hip_0_hip_pipe_txsynchd3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd3),        //  output,   width = 2,                          .txsynchd3
		.pcie_a10_hip_0_hip_pipe_txsynchd4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd4),        //  output,   width = 2,                          .txsynchd4
		.pcie_a10_hip_0_hip_pipe_txsynchd5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd5),        //  output,   width = 2,                          .txsynchd5
		.pcie_a10_hip_0_hip_pipe_txsynchd6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd6),        //  output,   width = 2,                          .txsynchd6
		.pcie_a10_hip_0_hip_pipe_txsynchd7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txsynchd7),        //  output,   width = 2,                          .txsynchd7
		.pcie_a10_hip_0_hip_pipe_txblkst0         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst0),         //  output,   width = 1,                          .txblkst0
		.pcie_a10_hip_0_hip_pipe_txblkst1         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst1),         //  output,   width = 1,                          .txblkst1
		.pcie_a10_hip_0_hip_pipe_txblkst2         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst2),         //  output,   width = 1,                          .txblkst2
		.pcie_a10_hip_0_hip_pipe_txblkst3         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst3),         //  output,   width = 1,                          .txblkst3
		.pcie_a10_hip_0_hip_pipe_txblkst4         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst4),         //  output,   width = 1,                          .txblkst4
		.pcie_a10_hip_0_hip_pipe_txblkst5         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst5),         //  output,   width = 1,                          .txblkst5
		.pcie_a10_hip_0_hip_pipe_txblkst6         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst6),         //  output,   width = 1,                          .txblkst6
		.pcie_a10_hip_0_hip_pipe_txblkst7         (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txblkst7),         //  output,   width = 1,                          .txblkst7
		.pcie_a10_hip_0_hip_pipe_txdataskip0      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip0),      //  output,   width = 1,                          .txdataskip0
		.pcie_a10_hip_0_hip_pipe_txdataskip1      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip1),      //  output,   width = 1,                          .txdataskip1
		.pcie_a10_hip_0_hip_pipe_txdataskip2      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip2),      //  output,   width = 1,                          .txdataskip2
		.pcie_a10_hip_0_hip_pipe_txdataskip3      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip3),      //  output,   width = 1,                          .txdataskip3
		.pcie_a10_hip_0_hip_pipe_txdataskip4      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip4),      //  output,   width = 1,                          .txdataskip4
		.pcie_a10_hip_0_hip_pipe_txdataskip5      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip5),      //  output,   width = 1,                          .txdataskip5
		.pcie_a10_hip_0_hip_pipe_txdataskip6      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip6),      //  output,   width = 1,                          .txdataskip6
		.pcie_a10_hip_0_hip_pipe_txdataskip7      (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_txdataskip7),      //  output,   width = 1,                          .txdataskip7
		.pcie_a10_hip_0_hip_pipe_rate0            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate0),            //  output,   width = 2,                          .rate0
		.pcie_a10_hip_0_hip_pipe_rate1            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate1),            //  output,   width = 2,                          .rate1
		.pcie_a10_hip_0_hip_pipe_rate2            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate2),            //  output,   width = 2,                          .rate2
		.pcie_a10_hip_0_hip_pipe_rate3            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate3),            //  output,   width = 2,                          .rate3
		.pcie_a10_hip_0_hip_pipe_rate4            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate4),            //  output,   width = 2,                          .rate4
		.pcie_a10_hip_0_hip_pipe_rate5            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate5),            //  output,   width = 2,                          .rate5
		.pcie_a10_hip_0_hip_pipe_rate6            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate6),            //  output,   width = 2,                          .rate6
		.pcie_a10_hip_0_hip_pipe_rate7            (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_pipe_rate7),            //  output,   width = 2,                          .rate7
		.pcie_a10_hip_0_hip_serial_rx_in0         (dut_pcie_tb_hip_serial_rx_in0),                                 //   input,   width = 1, pcie_a10_hip_0_hip_serial.rx_in0
		.pcie_a10_hip_0_hip_serial_rx_in1         (dut_pcie_tb_hip_serial_rx_in1),                                 //   input,   width = 1,                          .rx_in1
		.pcie_a10_hip_0_hip_serial_rx_in2         (dut_pcie_tb_hip_serial_rx_in2),                                 //   input,   width = 1,                          .rx_in2
		.pcie_a10_hip_0_hip_serial_rx_in3         (dut_pcie_tb_hip_serial_rx_in3),                                 //   input,   width = 1,                          .rx_in3
		.pcie_a10_hip_0_hip_serial_rx_in4         (dut_pcie_tb_hip_serial_rx_in4),                                 //   input,   width = 1,                          .rx_in4
		.pcie_a10_hip_0_hip_serial_rx_in5         (dut_pcie_tb_hip_serial_rx_in5),                                 //   input,   width = 1,                          .rx_in5
		.pcie_a10_hip_0_hip_serial_rx_in6         (dut_pcie_tb_hip_serial_rx_in6),                                 //   input,   width = 1,                          .rx_in6
		.pcie_a10_hip_0_hip_serial_rx_in7         (dut_pcie_tb_hip_serial_rx_in7),                                 //   input,   width = 1,                          .rx_in7
		.pcie_a10_hip_0_hip_serial_tx_out0        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out0),        //  output,   width = 1,                          .tx_out0
		.pcie_a10_hip_0_hip_serial_tx_out1        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out1),        //  output,   width = 1,                          .tx_out1
		.pcie_a10_hip_0_hip_serial_tx_out2        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out2),        //  output,   width = 1,                          .tx_out2
		.pcie_a10_hip_0_hip_serial_tx_out3        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out3),        //  output,   width = 1,                          .tx_out3
		.pcie_a10_hip_0_hip_serial_tx_out4        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out4),        //  output,   width = 1,                          .tx_out4
		.pcie_a10_hip_0_hip_serial_tx_out5        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out5),        //  output,   width = 1,                          .tx_out5
		.pcie_a10_hip_0_hip_serial_tx_out6        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out6),        //  output,   width = 1,                          .tx_out6
		.pcie_a10_hip_0_hip_serial_tx_out7        (ep_g3x8_avmm256_inst_pcie_a10_hip_0_hip_serial_tx_out7),        //  output,   width = 1,                          .tx_out7
		.pcie_a10_hip_0_npor_npor                 (dut_pcie_tb_npor_npor),                                         //   input,   width = 1,       pcie_a10_hip_0_npor.npor
		.pcie_a10_hip_0_npor_pin_perst            (dut_pcie_tb_npor_pin_perst),                                    //   input,   width = 1,                          .pin_perst
		.reconfig_xcvr_clk_clk                    (ep_g3x8_avmm256_inst_reconfig_xcvr_clk_bfm_clk_clk),            //   input,   width = 1,         reconfig_xcvr_clk.clk
		.reconfig_xcvr_reset_reset_n              (ep_g3x8_avmm256_inst_reconfig_xcvr_reset_bfm_reset_reset),      //   input,   width = 1,       reconfig_xcvr_reset.reset_n
		.refclk_clk                               (dut_pcie_tb_refclk_clk)                                         //   input,   width = 1,                    refclk.clk
	);

endmodule
