`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LCR2MnCRkjfWr/Vf9MUl+9b0TJDPPCW5qM7EkwiHp5FDFJbXEZD+QaBdf/NFoQX9
Hzx+USN/zIEl0J8HZW9pyzZOrpRrnnetYoT79F3yTYAwvJZVY5N35AXx4tcg97/C
XslM8R5TCBI5n9JlUOPoaDfWJOsTd+QA1oaqikmLEco=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
ar1yX5D4kw0gq5l4w8Mwmi8BD8Xlry17WlnHKNpJsuDH6Z5xIuFh+PCZxMhzHznP
jn+QC4ipsSsdzaQ0ymEUSQskFavlL8nZoG7Q+kYyypmyO0fRkYx21Vg/RXkfa93+
kfeTUckxQTWTbEMT2HNZhThgbjzGfN2EdN8ZtNv1oL7pjCGMYnx5YxVyfcsvGX/+
yA2jKtdwIdxKXzgrX4BJU5eETif2Fc2XhULN1dfe1XIfM+Q+ajIvEJUL9nhm++/j
e4q/+llEA/DqmhhjKuhQsrMYeaO5urUqt9QDyjEDSp55eNeMIl9+ffnRuA0Ziq8u
5rgECUcfBEW3b4rzr3GhP3SmHv+rpRG7uU5gvwiHM0V9OdoIc7do1BO+HAr/+CLR
nBIehnNVDsaGJd4RS6g8N+j76J4lu6+2xoh6RiQ6Wg7kkmm5kb0/9R+lYgeoeBes
2eo3qH+5Q9eNzNARDypEH+z6YFSddymBwPlI83N2Y7eMkVNwOhvPc/8kl/yqzTTu
JOyn2Zmry2R4ww5Y3Yi937lE/J2XUnkAAHn/42SCHSTP7JmkCq6ufq4DwiQpjRJc
hK96A0o6WSkKA/8nPuyWVdmPQBbP6OERMJf+27oaniOhU9i/9URjFqeqCMflne3d
IJWxyDU5OXgR9j2yxfA71HsKV8j6/DhWp+y0H3pPt71wiIXgHaro04q1qP3XhY5v
GM+Ei0GYyIm/3ALNQEuvf3qlSET9oyh4So0hJ0WMhTzKKmFotBJvUbT5uAFZiBxl
nYaPN233HXfwG2hCFMUESURThr9hpdn1IkJwW9/d2TZV3gmGqtx8nxfY0G7OIJo5
AD3km7Q6q4cypl5WQ+dOWecsK146pOnrjNrpwkMSOS/qqf4B4UE2gptFoALj8f8E
R/JgxH5Ucedqr3Yd0+hcN4YOQmxVSvhSrhVYNFZCxfe7dTmBD82Ng4VT84bDvsFn
WJyoUk2+NHZUi5wvSqyyKMkwx+GsqlV8rzuCqQLWiQVuifdRo9IHWB29h6Avu/oO
QhBeKjnG0bVebQSssHAcxqZwaB8bu2Ga5rLG4V2Gm6bmnJH3gC5wDHLJLJlhfY3P
Q0ITDsoZ7XrDC98oDQ1DLCI76cHQlrrlqs2ChwEl7NpXQZP7pMaUKeB6cxIneMej
90wCAhwz/yY3xI/MHoIapeGziVbORyn04QqmTSjlFRtA8QJs+OuFPmLJWU7xw8UJ
UgcLp4JHomlAsmuwN1kblKfmPSJI8BA49IF0MkVSKhLPLyfdy5PLttGFx1gdXlV+
/qc7eNX1dhDWwT82vlizfNwUJLtEatDoHQcQ0PvzcDcUKSTG5mVF9X6En28GZFVf
KmWvutLBAhBVQthk3gNgaXVWX6O9waQSnSTOBe8loG9TthLtQvOrmEBZBLWbDQrQ
SEvrfZH/FrKw2/SxorfpLBY2nG1jWflbINPAy6id8P2ktZIhZ38uOZpZToIMwiHS
jABJbRfu4XtlzkG/p3//xpvl03UklU53w6nBn1MEYCtdrPWvtoM+XiElBgMTjIBP
wdgH+g2WmrWwRGVcPWxMNrQi7Bmtr/LbEu3VIFXOmBMW8opQNv5vfc1Jiuyw7LXn
5KAFyrAjoA0BAQCQPCEFJ+Ur0LpXqwVBS7tfSOjrAdoT4JNxcBPUB7wiwut/Sg8L
Oojb9o5rmEirobBV88wj+v74hH9SHFt/Pqh61FU0hxVwFRRMpH3XtLCEci2l5hYp
tsdyxd0Ff4hNZHDPRQ7j/xauxTpCDReY6JVH/BEwUSFgwHle5PSf0742mzBTipEW
1VjzdPo6gpSYLl/y27qJNVzC7rf/n6Qq+nYmuKLui2FwbTJrWs1vNXEnKgjzcvLE
61MtbgQsa8polgZq1ek5tgMw6+H0QDW0Bv925NLhiSiWHSbphQr4goZfICfcv667
40GLiD8jHp68xqTdtGo4Yt1JXSREPbI81M/Mbw+GTZRNYId1VRntVwhaeU/D3EVO
BwfxY0LYuiNzRybjJwOCa2ABx4Wep73g37+JEGYeM+ERfguvudOEkd1QUf+xB18A
6T1RCC3Nt6HDxVjJlUGgVVzu8u2CxhHHyrLyviHwrtDwbBH9gv32fjBedPzT7SoM
Sl6rzouCy+vSO8dKSGuV2zUomZTiK5nQv7riEoKHdpSnLKAg1dWW53EzA+ozlfYQ
THkpaCh7ynpXk1egvweCUBAvL/7ChGanfltEtA1qCyIrGA6U6nDJSd+gyDfOaTtQ
jMcYS2FRNySj5Y1a8l9c2+Gqeb6aG5gAHLdsEVAQURQqrHqaG0PmTHO/0YhTR8PH
oQr6TTRXN7pumsd3/ALtkUJhavIZNQqW3XxQys6VfN75Z/DiA4aY8NYUJr2BKx6x
iPgLuZAFhXtTSvt3tRWLVL6uo0r4Y4bd8PEKWDHGg7gXgbNSawjc5hy3eUgrtXjK
6maTuR/TJFz2jA+iWOOG7zVcXv6l0bMXjjOkOfDj2gfeHdScVnJGy+jy2l9l8jku
nHIpesyDeroir9rEZGf3mol0P+JDDQZUpBho6F6ewzM57cOzPKPJY6eJr4DROlUm
MwSfeCuoXXgkgtO1PmaECbSXlfzbQSB3mpda6jj5I6II0hNUWqvAIJZG1594a2pM
SzhYeIJPQn6uteYr6qwlt8aZsQ62LTnY4xpTCfJ0UkmOjDbTwpliVHdWG23ex5KT
k2LOK4ZpF2WJbQeBSBU9TyB1ACSnFCwacw21iV4CLW+BIZTfnOPlBTaoaWcNQC9Z
vnpUBVtam108G0OgdcyPl58LtJARaWKZdi0pj0UFDqIjBtn5772351vcF+c7Smig
j00ZPtTWnYvKh6fxUW0K+w+WPSHkMWIj6tyvyVOMz5wVvPOq/2EGFQFcwtYnIsE7
LR1u1hSnCXzBtFfaW9OqawB1tjoISNeqoy6Su/PP+RkvKhhHpCzLP3mpOK1u5XL8
4RgnPdPf9ky1I00AjB0ykdF2JYHYUBe5UXOX7/fBKrZIGUIXXNygVzRMuSeU+ZD5
xlrgdE0RqumPEp3nKmIqRPHjXME1g30lRLCnzS2N0skT3A94qVLegyMzerXt9ECP
4XHasyWhmlmid/53SefzxfoCNgjVSbs//ocPsWxle4fIhDSEj9gTyh3gc7yP3tXj
VBitvKtJE03o62ZXKqmPLqQ0+XyV0LPSmTDsRcpS6VMTi//ctEMLmhzA/Qn2Oek2
anaippfiyKphp/6quoYktdYEwNjyEjA5Uypz7D6c6gaLt3FyR/0UcuBOjZj4eb2E
8BrfVX4WnXG2b3uy608BWlGOMRFHIzYFmeU4RhaEREMl37p20uZ+/jSulz3GlQz+
iCumUquFgMHuoEHcb0/TbC+VQc0Fzutpf4VaQmIoam/wRZ+s69DdJb3Pua63BQ/X
YvdyAa1suTxBwgofU1xkRzUadftHVCMe/prDmy0EGSDunjNQQ0l+h9q6cs14k1zH
tRxXAf/JJ0Nk3UhVfKv4VuiqvBKVz/KFG+tciBfsAsg+kb6sy28M9tH8UxPZS9A3
15ZpK0vprs9En9nUVLdzeWMGIk4cUfx++UKxJ8BpqSZiKMbjeoIEYCNbf8KVnZkK
enbqlApAuxEMgACoj8F49/kPHJwzhiN+i6nZD5R1KAxe/nq9cAs/gG1vd47YHcKo
bZBZJR9Ux6RLgi26AHysxqmf4gAL0mlmE5wy+Eq/EM+7rREwyN5tmg0J6L0dJPpT
RhE/MNVZVkzkJtuYXFU411UCzZWkij5Q4DEiuYyxqjpSWH6AWOk3jsxDpCE0xP+h
1LNtj42muI13PIMsKf6XGs02sr57gHsjL7mgz+nlEtkiAP2Hj7AXi9NWFtQ8AX9C
ovDVVq1gKdWFIXivZts/a7ivLQfQiwCUJDsntDNa7pB6aZJFP9HzdMd1vU2mw8jR
VlhXQfIDouhpwG7Xrec9w9mr5Yj4ds90RQR/ZypyU7kotqNB2wtVEtZexnC1WscJ
/3kUp+aMl6IiFy0jWR9cgT1gq0uGNqJey9yRd45ZloRymkBUDFAjeqE3YiEdWA/u
eDgrHbp2F4WCOzWVqMcInR6XGsCiQu+EKxQyWNb2HKg/8w/H0j5R3jZDbH01uOcU
tdSOEaRn6MtIJzBCG6LCsVzNO9Gp92ggh787y7K8MpfGYK5RQglEnhYSSt1YmgDp
jiw/lNto5zz9aB1iJMfhsAz5+3Zqpep4SH3uN8uG2VH/6VKzmQklSAh+dmGNwAkH
UPoHyZbEZow330j7wSXkyJV440wpQXm/H7R6rFaMMeAjVhkrEcZWlUThYHz6hfsa
R/Xr9Fthzw2dfRW6Mw3uH+7nihD6v9oTpHuBSmT5113k0LfqGZDX7FJUwico+QC0
0oiteUU9L2FnswrZV7gQOXvq56mdR1aHCHZg/DDuw54Ds71H8Vq46+UwIzVDxYYB
OnbeBJBrXh48Am1Vib2I+cg5Y7bTqJik4UExu0NTztdkdMxZ5nquMOz0UY07+okq
v7JEzKXJrflvSc15+mQXopk/5JvBO4ozQO4ZrNtbdCo1PpS/3kncptyMZd0Sibsv
DvdsJjTbnn9ditnEe9GIPCcXeOxeTplt6pZisx8MyqZCIha1geIRfqIfjA+eUhsZ
rbiSWBjH+rwRMhAizjUWzzN7s0LZdTQ9N+wPe6o2CYFNDrCCu9l3eI8IVTzeKUHp
GfmamYeje9Xo1zzTeSTmtRkASWINvTu9K2MZqMTCc4Nmsbk4u0Z3g/gmdiqG+W8S
fTbAUPCDOlwH0p/p6u5KGJG14Bn+1P5WxUQ2oaZWwNb3S/d6dPejqfT6Y0SoJU7a
kQDdxkyPuZeNe03J3V/dlRYZRUBRDPZgi4ck+ayBi1jPtq5Uaxc0uaVZivVa7GPg
B+uDonZLFczFqD6YkYIAwJxxKvZX2C69MTUp3rjG6maPZv5MpM1Gi53YAwHWCkfy
9jPw4y//+IYjHXBJOumJu5/QjEVvIqxfCJFctaS3ktNb5yfwBYU0O/g9A+vZ2dBA
jr43YNpwR7ctn0ANDp8VkNMCIFOPDGyD2r7lROjqqVX+Vx/4sTFr1pzkqbouDYYi
0d4cNCUD949I38wPs9iZmtzdGLP5hl/1Ko8UP/O+3awvbcmED7acAVBAa92YwIuJ
sWIud2kBvCU+xAdHMIvE+PnBxf7g609SSAVDuyVlTYCjZ3e6e8Nk6AdND2/NEcBe
Pv/ETnnygqgB4ybbYqIJdM08tT8SCMtcmvYM4VWuC7E7HPTLqNFjj9a10VlNPZkv
3zWIx4MrOlHa1yoNb7+TmCU33FaBFxZ+2Zgki7TB46YGIEZ8xH2Qemdhd8UChdL0
64KSONc1UGdjp1RGo2tFWs5CuMWi2iBt4ytaZ8aHzX+0N2iKecRXzEsm2Kzkoruc
hOX5Je2l2sHv/5czdkG8vC4iQATkMuSQRqoj1C8BIsxqpOD6X8kL88HTk+L8fqbe
eRpTT+xlmrajiwJFWe+otlSI5y0PyqKxMQ2C9oyPyi1nZ7Vk6WXO8D0pYyfIYC6Q
YpHH+hEMpO7Aoxij5f1RFme/CYcMwBQEJEcK8GzTtlXPLgrk+oeXwmFKrJro7jep
ZpwAy4wEkvfnRNNSXKKWKcjIfsONUa8qY2XOlB2Tz0aO1yeLZQJ3UPDbaYAib0Sa
TCG0n4AjN5iVNytrn0SRJ/ZcE4TYbUjF8wKcnRbNsSIPgkGwas9p/oUC4CapothI
krXcgm1ybMWAKv9t6DcW58Tq0NXYoFdL9BNEHhXDbj6CztJa57c126VLkQ2aOlmm
D+TwaoYUrGTUGEaia8NPSsatpKnLVgXzJsWyVMgeE1/L4qaM3c/mr3z7yC2oI9gK
qHA5B6EM9rEk4pbTXaCZ3Ub8p2kLyeK3vGazWI6X93ZwRaYjde/dq8bFz+tGh2UL
POOEx4Ry1AboIP1JYa8U2wm4BV833aqIIFsiKxQdRzp0hLRwKqcqsEypwS/XXNbG
7f2uTJZc/BZSzunSY9HPYjdwmnF0piBUIgp6j9CJY4Xgu5h/uwJS8shIHSk+p9WN
78I9YgeN8TdTkhkj108SKnsFSDHXfD01m7T5UUUIjMjJqqIE9g1CAWb+hJrb7kWR
LF4zQzZbpTvjJ7xz81qaoRhoMccxpmKjmhwBcTZVhccLsUtqZ8fTcB1XINkyKq2n
8jYxaN5gJ+Qdk+VNYGpFyG6W6lbiM7fl//APP4Y3Qzs1h4LPeCVWxOdFgDaWuyQf
WqxeMyLn2JRRxzXxiqsFOqm5HeV48uXVXCeAXGjUlH9wtHHNIrU8TClhVvd8U/tY
1gGHP6R7YT/5aegfsmWvRe199tbA6rNbPgID3oF2Wlp6VFmFJ3w/5oILEatm3xUJ
1iYUgZgoHPW+hm070t39nYkF1T8OgAwb+rlTzIN3Qikp30dSGYswOjGi12gdeilf
sVZe8uHNQMJyghhTIiGmxx1qxiX3CgEGCgRtKloAVb5eUFKiIG4D6PiVYdUV/oxt
kEa26vJ8+GtlCIurx1v9ryQmVDvcSOPiY7uSFgmUyehF0DU3JSoAnWHspbdu87lG
uzbhrzX+/rDCw+1mfA+Dy+/5ItmlqRJPNMymhvyxAHQDNMseNlB6vYKSSgXtmo2/
GSUacw1hTXUTgzF3hXoHJJBqJKesBYDSEJHSDa53XIQSWeARHBDTUAlYEg83+hzC
4on0kln5d3YpMa5M7oAHHFdwZwkChCV/zGo3tuGBpN3jhSd4IVgIpbvaFe83RwwY
MICNmu3wafH/f2GuXp/Vmo5FCNm9HNnbRh0bI67+fnxpHhg6/pWvSC8gAeSuAk7e
QG0VQ6OPA3fBBiBYLOrkcld9UV8mORDK9HWkvmsCFq4s0IXosmdDxSVMVlLfr4ui
kM0BAVMx19vF8UJNsHeMMyEgYU5T5YUQT+WumLVqVpRa6OiNoW1go7XBTN0WpAdj
O1CbPmDDeTb7qbJFAAYDVEwpmoE/y5+InYf4fv3xx+XAynXZJkePbXjpVgQHc0qg
hABs5LPL7boJHloKbh0sN5W96XlTTx1UPUd3UCVIog/lx+6fHk0jum+qvofwNDDW
BLb5AhVer+2Vz36KXVZml4IZTW+1chTsFYLpfzTW8eiaK/yVmTlW+KaK/+iJrESM
YUfM9VwdIR5+3u7r7JoV1QJnWuPcTxA1dUbrVzilgx6t4JzlCBfuyb5RoQkbOYH9
T0sfcz652Frb6ZwBkZOmFoC2Z1TDl4kg6AQxCsepOSzaHY6qAAtQ62y2Rs60Q4Wb
MN8FRZUwv7GNiD+opkxyflEjTWQAIO457tAzR0F4ylQTFNMQpL6xcK8l4KrBlC1/
4//4WcaOeiZxy2HifG71oJG4R/xxme/oAwE+RlOw5J7YW0uc8NCQ+tNluuRugW6n
4U4VHChFO4ZCKOoX5HQOIXaaJL4SIPHi5hHB9X/pZumw6mbCstxagtWlN3KZRk/y
5/pqz81uQK8nijp16jp3VTmxv/8hF0C3otpHR517QkSgHm7a2aXVXK7zeUdQmPl5
7EazlmQbxxzjgRc5TdYVzyYeUBxuUlkr6n2s3WDKzJmgR2FCwrA2HNrUH6hz4uzS
wMlqq6015hldVAKuBowfegE9wKkkt1NphGbFpHZQFpX1vU6d4/0zACMh/MpErVhh
IKvb+4iGDJOMZNBmHj3jV7tiYDh3naIdb263QjMMXi8bC17vxxhAjyI3oHRu8FBU
Cxs6awfSjrFp1jP3Gg88Y0v29Vuhanwb1N75sj2lX7RC5rzLlYkvvUDDpV5LBhXh
NqvQ33omJPIaIGoAgZoLH5PURhtv2T0L4i3roJx9MTzA72uJPPy1iHD474IwwMrj
F0kG276mv7dXT7D6tmGs5Ucs189L/9qw/9UQMN1yRpgSFmv4N9TWJTzX5pGQqx/r
6CY7K09aFvVqKLwT5iXtl8hwaEvB4is9e1wnxHapN0VM76TRAc1JOD33p+nA3v6q
utztLR4GuL3syOoS8HvH6JDrEw8QFYSiGFIBXAI27Op//HyPLMZyrt8RFslBFajE
+z88AldqR2Ur9YXbjvlYmTaxYfLiQoXnyse4NS2+RlRKwZMByFKiPTYq26zZwwh7
kvDerwoSJH96Q4eVxkKpl4W1t5oOJAI0BBzynkytxA1eZPaeX5VvBH3w6epH6Jnf
ErBYUgY+l/c8P3MEHO+/bj34wRWo+Y2lydJX/n0wf20gJqGO1RpaEK4KyVB7sQ7m
8nghgX1shm8oxPmDhoOQEmiVss1g35drtxE3HRm3OWfGm7hmLTtlMJu4QRoP5da8
WAQgIesK036YS8orM/fz3w==
`pragma protect end_protected
