///////////////////////////////////////////////////////////////////////
// File:  CRC32_D128.v                             
// Date:  Fri May 24 08:39:32 2002                                                      
//                                                                     
// Copyright (C) 1999 Easics NV.                 
// This source file may be used and distributed without restriction    
// provided that this copyright statement is not removed from the file 
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose: Verilog module containing a synthesizable CRC function
//   * polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
//   * data width: 128
//                                                                     
// Info: jand@easics.be (Jan Decaluwe)                           
//       http://www.easics.com                                  
///////////////////////////////////////////////////////////////////////

  // polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
  // data width: 128
  // convention: the first serial data bit is D[127]
  function [31:0] nextCRC32_D128;

    input [127:0] Data;
    input [31:0] CRC;

    reg [127:0] D;
    reg [31:0] C;
    reg [31:0] NewCRC;

  begin

    D = Data;
    C = CRC;

    NewCRC[0] = D[127] ^ D[126] ^ D[125] ^ D[123] ^ D[119] ^ D[118] ^ 
                D[117] ^ D[116] ^ D[114] ^ D[113] ^ D[111] ^ D[110] ^ 
                D[106] ^ D[104] ^ D[103] ^ D[101] ^ D[99] ^ D[98] ^ 
                D[97] ^ D[96] ^ D[95] ^ D[94] ^ D[87] ^ D[85] ^ D[84] ^ 
                D[83] ^ D[82] ^ D[81] ^ D[79] ^ D[73] ^ D[72] ^ D[68] ^ 
                D[67] ^ D[66] ^ D[65] ^ D[63] ^ D[61] ^ D[60] ^ D[58] ^ 
                D[55] ^ D[54] ^ D[53] ^ D[50] ^ D[48] ^ D[47] ^ D[45] ^ 
                D[44] ^ D[37] ^ D[34] ^ D[32] ^ D[31] ^ D[30] ^ D[29] ^ 
                D[28] ^ D[26] ^ D[25] ^ D[24] ^ D[16] ^ D[12] ^ D[10] ^ 
                D[9] ^ D[6] ^ D[0] ^ C[0] ^ C[1] ^ C[2] ^ C[3] ^ C[5] ^ 
                C[7] ^ C[8] ^ C[10] ^ C[14] ^ C[15] ^ C[17] ^ C[18] ^ 
                C[20] ^ C[21] ^ C[22] ^ C[23] ^ C[27] ^ C[29] ^ C[30] ^ 
                C[31];
    NewCRC[1] = D[125] ^ D[124] ^ D[123] ^ D[120] ^ D[116] ^ D[115] ^ 
                D[113] ^ D[112] ^ D[110] ^ D[107] ^ D[106] ^ D[105] ^ 
                D[103] ^ D[102] ^ D[101] ^ D[100] ^ D[94] ^ D[88] ^ 
                D[87] ^ D[86] ^ D[81] ^ D[80] ^ D[79] ^ D[74] ^ D[72] ^ 
                D[69] ^ D[65] ^ D[64] ^ D[63] ^ D[62] ^ D[60] ^ D[59] ^ 
                D[58] ^ D[56] ^ D[53] ^ D[51] ^ D[50] ^ D[49] ^ D[47] ^ 
                D[46] ^ D[44] ^ D[38] ^ D[37] ^ D[35] ^ D[34] ^ D[33] ^ 
                D[28] ^ D[27] ^ D[24] ^ D[17] ^ D[16] ^ D[13] ^ D[12] ^ 
                D[11] ^ D[9] ^ D[7] ^ D[6] ^ D[1] ^ D[0] ^ C[4] ^ C[5] ^ 
                C[6] ^ C[7] ^ C[9] ^ C[10] ^ C[11] ^ C[14] ^ C[16] ^ 
                C[17] ^ C[19] ^ C[20] ^ C[24] ^ C[27] ^ C[28] ^ C[29];
    NewCRC[2] = D[127] ^ D[124] ^ D[123] ^ D[121] ^ D[119] ^ D[118] ^ 
                D[110] ^ D[108] ^ D[107] ^ D[102] ^ D[99] ^ D[98] ^ 
                D[97] ^ D[96] ^ D[94] ^ D[89] ^ D[88] ^ D[85] ^ D[84] ^ 
                D[83] ^ D[80] ^ D[79] ^ D[75] ^ D[72] ^ D[70] ^ D[68] ^ 
                D[67] ^ D[64] ^ D[59] ^ D[58] ^ D[57] ^ D[55] ^ D[53] ^ 
                D[52] ^ D[51] ^ D[44] ^ D[39] ^ D[38] ^ D[37] ^ D[36] ^ 
                D[35] ^ D[32] ^ D[31] ^ D[30] ^ D[26] ^ D[24] ^ D[18] ^ 
                D[17] ^ D[16] ^ D[14] ^ D[13] ^ D[9] ^ D[8] ^ D[7] ^ 
                D[6] ^ D[2] ^ D[1] ^ D[0] ^ C[0] ^ C[1] ^ C[2] ^ C[3] ^ 
                C[6] ^ C[11] ^ C[12] ^ C[14] ^ C[22] ^ C[23] ^ C[25] ^ 
                C[27] ^ C[28] ^ C[31];
    NewCRC[3] = D[125] ^ D[124] ^ D[122] ^ D[120] ^ D[119] ^ D[111] ^ 
                D[109] ^ D[108] ^ D[103] ^ D[100] ^ D[99] ^ D[98] ^ 
                D[97] ^ D[95] ^ D[90] ^ D[89] ^ D[86] ^ D[85] ^ D[84] ^ 
                D[81] ^ D[80] ^ D[76] ^ D[73] ^ D[71] ^ D[69] ^ D[68] ^ 
                D[65] ^ D[60] ^ D[59] ^ D[58] ^ D[56] ^ D[54] ^ D[53] ^ 
                D[52] ^ D[45] ^ D[40] ^ D[39] ^ D[38] ^ D[37] ^ D[36] ^ 
                D[33] ^ D[32] ^ D[31] ^ D[27] ^ D[25] ^ D[19] ^ D[18] ^ 
                D[17] ^ D[15] ^ D[14] ^ D[10] ^ D[9] ^ D[8] ^ D[7] ^ 
                D[3] ^ D[2] ^ D[1] ^ C[1] ^ C[2] ^ C[3] ^ C[4] ^ C[7] ^ 
                C[12] ^ C[13] ^ C[15] ^ C[23] ^ C[24] ^ C[26] ^ C[28] ^ 
                C[29];
    NewCRC[4] = D[127] ^ D[121] ^ D[120] ^ D[119] ^ D[118] ^ D[117] ^ 
                D[116] ^ D[114] ^ D[113] ^ D[112] ^ D[111] ^ D[109] ^ 
                D[106] ^ D[103] ^ D[100] ^ D[97] ^ D[95] ^ D[94] ^ 
                D[91] ^ D[90] ^ D[86] ^ D[84] ^ D[83] ^ D[79] ^ D[77] ^ 
                D[74] ^ D[73] ^ D[70] ^ D[69] ^ D[68] ^ D[67] ^ D[65] ^ 
                D[63] ^ D[59] ^ D[58] ^ D[57] ^ D[50] ^ D[48] ^ D[47] ^ 
                D[46] ^ D[45] ^ D[44] ^ D[41] ^ D[40] ^ D[39] ^ D[38] ^ 
                D[33] ^ D[31] ^ D[30] ^ D[29] ^ D[25] ^ D[24] ^ D[20] ^ 
                D[19] ^ D[18] ^ D[15] ^ D[12] ^ D[11] ^ D[8] ^ D[6] ^ 
                D[4] ^ D[3] ^ D[2] ^ D[0] ^ C[1] ^ C[4] ^ C[7] ^ C[10] ^ 
                C[13] ^ C[15] ^ C[16] ^ C[17] ^ C[18] ^ C[20] ^ C[21] ^ 
                C[22] ^ C[23] ^ C[24] ^ C[25] ^ C[31];
    NewCRC[5] = D[127] ^ D[126] ^ D[125] ^ D[123] ^ D[122] ^ D[121] ^ 
                D[120] ^ D[116] ^ D[115] ^ D[112] ^ D[111] ^ D[107] ^ 
                D[106] ^ D[103] ^ D[99] ^ D[97] ^ D[94] ^ D[92] ^ D[91] ^ 
                D[83] ^ D[82] ^ D[81] ^ D[80] ^ D[79] ^ D[78] ^ D[75] ^ 
                D[74] ^ D[73] ^ D[72] ^ D[71] ^ D[70] ^ D[69] ^ D[67] ^ 
                D[65] ^ D[64] ^ D[63] ^ D[61] ^ D[59] ^ D[55] ^ D[54] ^ 
                D[53] ^ D[51] ^ D[50] ^ D[49] ^ D[46] ^ D[44] ^ D[42] ^ 
                D[41] ^ D[40] ^ D[39] ^ D[37] ^ D[29] ^ D[28] ^ D[24] ^ 
                D[21] ^ D[20] ^ D[19] ^ D[13] ^ D[10] ^ D[7] ^ D[6] ^ 
                D[5] ^ D[4] ^ D[3] ^ D[1] ^ D[0] ^ C[1] ^ C[3] ^ C[7] ^ 
                C[10] ^ C[11] ^ C[15] ^ C[16] ^ C[19] ^ C[20] ^ C[24] ^ 
                C[25] ^ C[26] ^ C[27] ^ C[29] ^ C[30] ^ C[31];
    NewCRC[6] = D[127] ^ D[126] ^ D[124] ^ D[123] ^ D[122] ^ D[121] ^ 
                D[117] ^ D[116] ^ D[113] ^ D[112] ^ D[108] ^ D[107] ^ 
                D[104] ^ D[100] ^ D[98] ^ D[95] ^ D[93] ^ D[92] ^ D[84] ^ 
                D[83] ^ D[82] ^ D[81] ^ D[80] ^ D[79] ^ D[76] ^ D[75] ^ 
                D[74] ^ D[73] ^ D[72] ^ D[71] ^ D[70] ^ D[68] ^ D[66] ^ 
                D[65] ^ D[64] ^ D[62] ^ D[60] ^ D[56] ^ D[55] ^ D[54] ^ 
                D[52] ^ D[51] ^ D[50] ^ D[47] ^ D[45] ^ D[43] ^ D[42] ^ 
                D[41] ^ D[40] ^ D[38] ^ D[30] ^ D[29] ^ D[25] ^ D[22] ^ 
                D[21] ^ D[20] ^ D[14] ^ D[11] ^ D[8] ^ D[7] ^ D[6] ^ 
                D[5] ^ D[4] ^ D[2] ^ D[1] ^ C[2] ^ C[4] ^ C[8] ^ C[11] ^ 
                C[12] ^ C[16] ^ C[17] ^ C[20] ^ C[21] ^ C[25] ^ C[26] ^ 
                C[27] ^ C[28] ^ C[30] ^ C[31];
    NewCRC[7] = D[126] ^ D[124] ^ D[122] ^ D[119] ^ D[116] ^ D[111] ^ 
                D[110] ^ D[109] ^ D[108] ^ D[106] ^ D[105] ^ D[104] ^ 
                D[103] ^ D[98] ^ D[97] ^ D[95] ^ D[93] ^ D[87] ^ D[80] ^ 
                D[79] ^ D[77] ^ D[76] ^ D[75] ^ D[74] ^ D[71] ^ D[69] ^ 
                D[68] ^ D[60] ^ D[58] ^ D[57] ^ D[56] ^ D[54] ^ D[52] ^ 
                D[51] ^ D[50] ^ D[47] ^ D[46] ^ D[45] ^ D[43] ^ D[42] ^ 
                D[41] ^ D[39] ^ D[37] ^ D[34] ^ D[32] ^ D[29] ^ D[28] ^ 
                D[25] ^ D[24] ^ D[23] ^ D[22] ^ D[21] ^ D[16] ^ D[15] ^ 
                D[10] ^ D[8] ^ D[7] ^ D[5] ^ D[3] ^ D[2] ^ D[0] ^ C[1] ^ 
                C[2] ^ C[7] ^ C[8] ^ C[9] ^ C[10] ^ C[12] ^ C[13] ^ 
                C[14] ^ C[15] ^ C[20] ^ C[23] ^ C[26] ^ C[28] ^ C[30];
    NewCRC[8] = D[126] ^ D[120] ^ D[119] ^ D[118] ^ D[116] ^ D[114] ^ 
                D[113] ^ D[112] ^ D[109] ^ D[107] ^ D[105] ^ D[103] ^ 
                D[101] ^ D[97] ^ D[95] ^ D[88] ^ D[87] ^ D[85] ^ D[84] ^ 
                D[83] ^ D[82] ^ D[80] ^ D[79] ^ D[78] ^ D[77] ^ D[76] ^ 
                D[75] ^ D[73] ^ D[70] ^ D[69] ^ D[68] ^ D[67] ^ D[66] ^ 
                D[65] ^ D[63] ^ D[60] ^ D[59] ^ D[57] ^ D[54] ^ D[52] ^ 
                D[51] ^ D[50] ^ D[46] ^ D[45] ^ D[43] ^ D[42] ^ D[40] ^ 
                D[38] ^ D[37] ^ D[35] ^ D[34] ^ D[33] ^ D[32] ^ D[31] ^ 
                D[28] ^ D[23] ^ D[22] ^ D[17] ^ D[12] ^ D[11] ^ D[10] ^ 
                D[8] ^ D[4] ^ D[3] ^ D[1] ^ D[0] ^ C[1] ^ C[5] ^ C[7] ^ 
                C[9] ^ C[11] ^ C[13] ^ C[16] ^ C[17] ^ C[18] ^ C[20] ^ 
                C[22] ^ C[23] ^ C[24] ^ C[30];
    NewCRC[9] = D[127] ^ D[121] ^ D[120] ^ D[119] ^ D[117] ^ D[115] ^ 
                D[114] ^ D[113] ^ D[110] ^ D[108] ^ D[106] ^ D[104] ^ 
                D[102] ^ D[98] ^ D[96] ^ D[89] ^ D[88] ^ D[86] ^ D[85] ^ 
                D[84] ^ D[83] ^ D[81] ^ D[80] ^ D[79] ^ D[78] ^ D[77] ^ 
                D[76] ^ D[74] ^ D[71] ^ D[70] ^ D[69] ^ D[68] ^ D[67] ^ 
                D[66] ^ D[64] ^ D[61] ^ D[60] ^ D[58] ^ D[55] ^ D[53] ^ 
                D[52] ^ D[51] ^ D[47] ^ D[46] ^ D[44] ^ D[43] ^ D[41] ^ 
                D[39] ^ D[38] ^ D[36] ^ D[35] ^ D[34] ^ D[33] ^ D[32] ^ 
                D[29] ^ D[24] ^ D[23] ^ D[18] ^ D[13] ^ D[12] ^ D[11] ^ 
                D[9] ^ D[5] ^ D[4] ^ D[2] ^ D[1] ^ C[0] ^ C[2] ^ C[6] ^ 
                C[8] ^ C[10] ^ C[12] ^ C[14] ^ C[17] ^ C[18] ^ C[19] ^ 
                C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[31];
    NewCRC[10] = D[127] ^ D[126] ^ D[125] ^ D[123] ^ D[122] ^ D[121] ^ 
                 D[120] ^ D[119] ^ D[117] ^ D[115] ^ D[113] ^ D[110] ^ 
                 D[109] ^ D[107] ^ D[106] ^ D[105] ^ D[104] ^ D[101] ^ 
                 D[98] ^ D[96] ^ D[95] ^ D[94] ^ D[90] ^ D[89] ^ D[86] ^ 
                 D[83] ^ D[80] ^ D[78] ^ D[77] ^ D[75] ^ D[73] ^ D[71] ^ 
                 D[70] ^ D[69] ^ D[66] ^ D[63] ^ D[62] ^ D[60] ^ D[59] ^ 
                 D[58] ^ D[56] ^ D[55] ^ D[52] ^ D[50] ^ D[42] ^ D[40] ^ 
                 D[39] ^ D[36] ^ D[35] ^ D[33] ^ D[32] ^ D[31] ^ D[29] ^ 
                 D[28] ^ D[26] ^ D[19] ^ D[16] ^ D[14] ^ D[13] ^ D[9] ^ 
                 D[5] ^ D[3] ^ D[2] ^ D[0] ^ C[0] ^ C[2] ^ C[5] ^ C[8] ^ 
                 C[9] ^ C[10] ^ C[11] ^ C[13] ^ C[14] ^ C[17] ^ C[19] ^ 
                 C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[26] ^ C[27] ^ C[29] ^ 
                 C[30] ^ C[31];
    NewCRC[11] = D[125] ^ D[124] ^ D[122] ^ D[121] ^ D[120] ^ D[119] ^ 
                 D[117] ^ D[113] ^ D[108] ^ D[107] ^ D[105] ^ D[104] ^ 
                 D[103] ^ D[102] ^ D[101] ^ D[98] ^ D[94] ^ D[91] ^ 
                 D[90] ^ D[85] ^ D[83] ^ D[82] ^ D[78] ^ D[76] ^ D[74] ^ 
                 D[73] ^ D[71] ^ D[70] ^ D[68] ^ D[66] ^ D[65] ^ D[64] ^ 
                 D[59] ^ D[58] ^ D[57] ^ D[56] ^ D[55] ^ D[54] ^ D[51] ^ 
                 D[50] ^ D[48] ^ D[47] ^ D[45] ^ D[44] ^ D[43] ^ D[41] ^ 
                 D[40] ^ D[36] ^ D[33] ^ D[31] ^ D[28] ^ D[27] ^ D[26] ^ 
                 D[25] ^ D[24] ^ D[20] ^ D[17] ^ D[16] ^ D[15] ^ D[14] ^ 
                 D[12] ^ D[9] ^ D[4] ^ D[3] ^ D[1] ^ D[0] ^ C[2] ^ C[5] ^ 
                 C[6] ^ C[7] ^ C[8] ^ C[9] ^ C[11] ^ C[12] ^ C[17] ^ 
                 C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[26] ^ C[28] ^ C[29];
    NewCRC[12] = D[127] ^ D[122] ^ D[121] ^ D[120] ^ D[119] ^ D[117] ^ 
                 D[116] ^ D[113] ^ D[111] ^ D[110] ^ D[109] ^ D[108] ^ 
                 D[105] ^ D[102] ^ D[101] ^ D[98] ^ D[97] ^ D[96] ^ 
                 D[94] ^ D[92] ^ D[91] ^ D[87] ^ D[86] ^ D[85] ^ D[82] ^ 
                 D[81] ^ D[77] ^ D[75] ^ D[74] ^ D[73] ^ D[71] ^ D[69] ^ 
                 D[68] ^ D[63] ^ D[61] ^ D[59] ^ D[57] ^ D[56] ^ D[54] ^ 
                 D[53] ^ D[52] ^ D[51] ^ D[50] ^ D[49] ^ D[47] ^ D[46] ^ 
                 D[42] ^ D[41] ^ D[31] ^ D[30] ^ D[27] ^ D[24] ^ D[21] ^ 
                 D[18] ^ D[17] ^ D[15] ^ D[13] ^ D[12] ^ D[9] ^ D[6] ^ 
                 D[5] ^ D[4] ^ D[2] ^ D[1] ^ D[0] ^ C[0] ^ C[1] ^ C[2] ^ 
                 C[5] ^ C[6] ^ C[9] ^ C[12] ^ C[13] ^ C[14] ^ C[15] ^ 
                 C[17] ^ C[20] ^ C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[26] ^ 
                 C[31];
    NewCRC[13] = D[123] ^ D[122] ^ D[121] ^ D[120] ^ D[118] ^ D[117] ^ 
                 D[114] ^ D[112] ^ D[111] ^ D[110] ^ D[109] ^ D[106] ^ 
                 D[103] ^ D[102] ^ D[99] ^ D[98] ^ D[97] ^ D[95] ^ D[93] ^ 
                 D[92] ^ D[88] ^ D[87] ^ D[86] ^ D[83] ^ D[82] ^ D[78] ^ 
                 D[76] ^ D[75] ^ D[74] ^ D[72] ^ D[70] ^ D[69] ^ D[64] ^ 
                 D[62] ^ D[60] ^ D[58] ^ D[57] ^ D[55] ^ D[54] ^ D[53] ^ 
                 D[52] ^ D[51] ^ D[50] ^ D[48] ^ D[47] ^ D[43] ^ D[42] ^ 
                 D[32] ^ D[31] ^ D[28] ^ D[25] ^ D[22] ^ D[19] ^ D[18] ^ 
                 D[16] ^ D[14] ^ D[13] ^ D[10] ^ D[7] ^ D[6] ^ D[5] ^ 
                 D[3] ^ D[2] ^ D[1] ^ C[1] ^ C[2] ^ C[3] ^ C[6] ^ C[7] ^ 
                 C[10] ^ C[13] ^ C[14] ^ C[15] ^ C[16] ^ C[18] ^ C[21] ^ 
                 C[22] ^ C[24] ^ C[25] ^ C[26] ^ C[27];
    NewCRC[14] = D[124] ^ D[123] ^ D[122] ^ D[121] ^ D[119] ^ D[118] ^ 
                 D[115] ^ D[113] ^ D[112] ^ D[111] ^ D[110] ^ D[107] ^ 
                 D[104] ^ D[103] ^ D[100] ^ D[99] ^ D[98] ^ D[96] ^ 
                 D[94] ^ D[93] ^ D[89] ^ D[88] ^ D[87] ^ D[84] ^ D[83] ^ 
                 D[79] ^ D[77] ^ D[76] ^ D[75] ^ D[73] ^ D[71] ^ D[70] ^ 
                 D[65] ^ D[63] ^ D[61] ^ D[59] ^ D[58] ^ D[56] ^ D[55] ^ 
                 D[54] ^ D[53] ^ D[52] ^ D[51] ^ D[49] ^ D[48] ^ D[44] ^ 
                 D[43] ^ D[33] ^ D[32] ^ D[29] ^ D[26] ^ D[23] ^ D[20] ^ 
                 D[19] ^ D[17] ^ D[15] ^ D[14] ^ D[11] ^ D[8] ^ D[7] ^ 
                 D[6] ^ D[4] ^ D[3] ^ D[2] ^ C[0] ^ C[2] ^ C[3] ^ C[4] ^ 
                 C[7] ^ C[8] ^ C[11] ^ C[14] ^ C[15] ^ C[16] ^ C[17] ^ 
                 C[19] ^ C[22] ^ C[23] ^ C[25] ^ C[26] ^ C[27] ^ C[28];
    NewCRC[15] = D[125] ^ D[124] ^ D[123] ^ D[122] ^ D[120] ^ D[119] ^ 
                 D[116] ^ D[114] ^ D[113] ^ D[112] ^ D[111] ^ D[108] ^ 
                 D[105] ^ D[104] ^ D[101] ^ D[100] ^ D[99] ^ D[97] ^ 
                 D[95] ^ D[94] ^ D[90] ^ D[89] ^ D[88] ^ D[85] ^ D[84] ^ 
                 D[80] ^ D[78] ^ D[77] ^ D[76] ^ D[74] ^ D[72] ^ D[71] ^ 
                 D[66] ^ D[64] ^ D[62] ^ D[60] ^ D[59] ^ D[57] ^ D[56] ^ 
                 D[55] ^ D[54] ^ D[53] ^ D[52] ^ D[50] ^ D[49] ^ D[45] ^ 
                 D[44] ^ D[34] ^ D[33] ^ D[30] ^ D[27] ^ D[24] ^ D[21] ^ 
                 D[20] ^ D[18] ^ D[16] ^ D[15] ^ D[12] ^ D[9] ^ D[8] ^ 
                 D[7] ^ D[5] ^ D[4] ^ D[3] ^ C[1] ^ C[3] ^ C[4] ^ C[5] ^ 
                 C[8] ^ C[9] ^ C[12] ^ C[15] ^ C[16] ^ C[17] ^ C[18] ^ 
                 C[20] ^ C[23] ^ C[24] ^ C[26] ^ C[27] ^ C[28] ^ C[29];
    NewCRC[16] = D[127] ^ D[124] ^ D[121] ^ D[120] ^ D[119] ^ D[118] ^ 
                 D[116] ^ D[115] ^ D[112] ^ D[111] ^ D[110] ^ D[109] ^ 
                 D[105] ^ D[104] ^ D[103] ^ D[102] ^ D[100] ^ D[99] ^ 
                 D[97] ^ D[94] ^ D[91] ^ D[90] ^ D[89] ^ D[87] ^ D[86] ^ 
                 D[84] ^ D[83] ^ D[82] ^ D[78] ^ D[77] ^ D[75] ^ D[68] ^ 
                 D[66] ^ D[57] ^ D[56] ^ D[51] ^ D[48] ^ D[47] ^ D[46] ^ 
                 D[44] ^ D[37] ^ D[35] ^ D[32] ^ D[30] ^ D[29] ^ D[26] ^ 
                 D[24] ^ D[22] ^ D[21] ^ D[19] ^ D[17] ^ D[13] ^ D[12] ^ 
                 D[8] ^ D[5] ^ D[4] ^ D[0] ^ C[1] ^ C[3] ^ C[4] ^ C[6] ^ 
                 C[7] ^ C[8] ^ C[9] ^ C[13] ^ C[14] ^ C[15] ^ C[16] ^ 
                 C[19] ^ C[20] ^ C[22] ^ C[23] ^ C[24] ^ C[25] ^ C[28] ^ 
                 C[31];
    NewCRC[17] = D[125] ^ D[122] ^ D[121] ^ D[120] ^ D[119] ^ D[117] ^ 
                 D[116] ^ D[113] ^ D[112] ^ D[111] ^ D[110] ^ D[106] ^ 
                 D[105] ^ D[104] ^ D[103] ^ D[101] ^ D[100] ^ D[98] ^ 
                 D[95] ^ D[92] ^ D[91] ^ D[90] ^ D[88] ^ D[87] ^ D[85] ^ 
                 D[84] ^ D[83] ^ D[79] ^ D[78] ^ D[76] ^ D[69] ^ D[67] ^ 
                 D[58] ^ D[57] ^ D[52] ^ D[49] ^ D[48] ^ D[47] ^ D[45] ^ 
                 D[38] ^ D[36] ^ D[33] ^ D[31] ^ D[30] ^ D[27] ^ D[25] ^ 
                 D[23] ^ D[22] ^ D[20] ^ D[18] ^ D[14] ^ D[13] ^ D[9] ^ 
                 D[6] ^ D[5] ^ D[1] ^ C[2] ^ C[4] ^ C[5] ^ C[7] ^ C[8] ^ 
                 C[9] ^ C[10] ^ C[14] ^ C[15] ^ C[16] ^ C[17] ^ C[20] ^ 
                 C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[26] ^ C[29];
    NewCRC[18] = D[126] ^ D[123] ^ D[122] ^ D[121] ^ D[120] ^ D[118] ^ 
                 D[117] ^ D[114] ^ D[113] ^ D[112] ^ D[111] ^ D[107] ^ 
                 D[106] ^ D[105] ^ D[104] ^ D[102] ^ D[101] ^ D[99] ^ 
                 D[96] ^ D[93] ^ D[92] ^ D[91] ^ D[89] ^ D[88] ^ D[86] ^ 
                 D[85] ^ D[84] ^ D[80] ^ D[79] ^ D[77] ^ D[70] ^ D[68] ^ 
                 D[59] ^ D[58] ^ D[53] ^ D[50] ^ D[49] ^ D[48] ^ D[46] ^ 
                 D[39] ^ D[37] ^ D[34] ^ D[32] ^ D[31] ^ D[28] ^ D[26] ^ 
                 D[24] ^ D[23] ^ D[21] ^ D[19] ^ D[15] ^ D[14] ^ D[10] ^ 
                 D[7] ^ D[6] ^ D[2] ^ C[0] ^ C[3] ^ C[5] ^ C[6] ^ C[8] ^ 
                 C[9] ^ C[10] ^ C[11] ^ C[15] ^ C[16] ^ C[17] ^ C[18] ^ 
                 C[21] ^ C[22] ^ C[24] ^ C[25] ^ C[26] ^ C[27] ^ C[30];
    NewCRC[19] = D[127] ^ D[124] ^ D[123] ^ D[122] ^ D[121] ^ D[119] ^ 
                 D[118] ^ D[115] ^ D[114] ^ D[113] ^ D[112] ^ D[108] ^ 
                 D[107] ^ D[106] ^ D[105] ^ D[103] ^ D[102] ^ D[100] ^ 
                 D[97] ^ D[94] ^ D[93] ^ D[92] ^ D[90] ^ D[89] ^ D[87] ^ 
                 D[86] ^ D[85] ^ D[81] ^ D[80] ^ D[78] ^ D[71] ^ D[69] ^ 
                 D[60] ^ D[59] ^ D[54] ^ D[51] ^ D[50] ^ D[49] ^ D[47] ^ 
                 D[40] ^ D[38] ^ D[35] ^ D[33] ^ D[32] ^ D[29] ^ D[27] ^ 
                 D[25] ^ D[24] ^ D[22] ^ D[20] ^ D[16] ^ D[15] ^ D[11] ^ 
                 D[8] ^ D[7] ^ D[3] ^ C[1] ^ C[4] ^ C[6] ^ C[7] ^ C[9] ^ 
                 C[10] ^ C[11] ^ C[12] ^ C[16] ^ C[17] ^ C[18] ^ C[19] ^ 
                 C[22] ^ C[23] ^ C[25] ^ C[26] ^ C[27] ^ C[28] ^ C[31];
    NewCRC[20] = D[125] ^ D[124] ^ D[123] ^ D[122] ^ D[120] ^ D[119] ^ 
                 D[116] ^ D[115] ^ D[114] ^ D[113] ^ D[109] ^ D[108] ^ 
                 D[107] ^ D[106] ^ D[104] ^ D[103] ^ D[101] ^ D[98] ^ 
                 D[95] ^ D[94] ^ D[93] ^ D[91] ^ D[90] ^ D[88] ^ D[87] ^ 
                 D[86] ^ D[82] ^ D[81] ^ D[79] ^ D[72] ^ D[70] ^ D[61] ^ 
                 D[60] ^ D[55] ^ D[52] ^ D[51] ^ D[50] ^ D[48] ^ D[41] ^ 
                 D[39] ^ D[36] ^ D[34] ^ D[33] ^ D[30] ^ D[28] ^ D[26] ^ 
                 D[25] ^ D[23] ^ D[21] ^ D[17] ^ D[16] ^ D[12] ^ D[9] ^ 
                 D[8] ^ D[4] ^ C[2] ^ C[5] ^ C[7] ^ C[8] ^ C[10] ^ C[11] ^ 
                 C[12] ^ C[13] ^ C[17] ^ C[18] ^ C[19] ^ C[20] ^ C[23] ^ 
                 C[24] ^ C[26] ^ C[27] ^ C[28] ^ C[29];
    NewCRC[21] = D[126] ^ D[125] ^ D[124] ^ D[123] ^ D[121] ^ D[120] ^ 
                 D[117] ^ D[116] ^ D[115] ^ D[114] ^ D[110] ^ D[109] ^ 
                 D[108] ^ D[107] ^ D[105] ^ D[104] ^ D[102] ^ D[99] ^ 
                 D[96] ^ D[95] ^ D[94] ^ D[92] ^ D[91] ^ D[89] ^ D[88] ^ 
                 D[87] ^ D[83] ^ D[82] ^ D[80] ^ D[73] ^ D[71] ^ D[62] ^ 
                 D[61] ^ D[56] ^ D[53] ^ D[52] ^ D[51] ^ D[49] ^ D[42] ^ 
                 D[40] ^ D[37] ^ D[35] ^ D[34] ^ D[31] ^ D[29] ^ D[27] ^ 
                 D[26] ^ D[24] ^ D[22] ^ D[18] ^ D[17] ^ D[13] ^ D[10] ^ 
                 D[9] ^ D[5] ^ C[0] ^ C[3] ^ C[6] ^ C[8] ^ C[9] ^ C[11] ^ 
                 C[12] ^ C[13] ^ C[14] ^ C[18] ^ C[19] ^ C[20] ^ C[21] ^ 
                 C[24] ^ C[25] ^ C[27] ^ C[28] ^ C[29] ^ C[30];
    NewCRC[22] = D[124] ^ D[123] ^ D[122] ^ D[121] ^ D[119] ^ D[115] ^ 
                 D[114] ^ D[113] ^ D[109] ^ D[108] ^ D[105] ^ D[104] ^ 
                 D[101] ^ D[100] ^ D[99] ^ D[98] ^ D[94] ^ D[93] ^ D[92] ^ 
                 D[90] ^ D[89] ^ D[88] ^ D[87] ^ D[85] ^ D[82] ^ D[79] ^ 
                 D[74] ^ D[73] ^ D[68] ^ D[67] ^ D[66] ^ D[65] ^ D[62] ^ 
                 D[61] ^ D[60] ^ D[58] ^ D[57] ^ D[55] ^ D[52] ^ D[48] ^ 
                 D[47] ^ D[45] ^ D[44] ^ D[43] ^ D[41] ^ D[38] ^ D[37] ^ 
                 D[36] ^ D[35] ^ D[34] ^ D[31] ^ D[29] ^ D[27] ^ D[26] ^ 
                 D[24] ^ D[23] ^ D[19] ^ D[18] ^ D[16] ^ D[14] ^ D[12] ^ 
                 D[11] ^ D[9] ^ D[0] ^ C[2] ^ C[3] ^ C[4] ^ C[5] ^ C[8] ^ 
                 C[9] ^ C[12] ^ C[13] ^ C[17] ^ C[18] ^ C[19] ^ C[23] ^ 
                 C[25] ^ C[26] ^ C[27] ^ C[28];
    NewCRC[23] = D[127] ^ D[126] ^ D[124] ^ D[122] ^ D[120] ^ D[119] ^ 
                 D[118] ^ D[117] ^ D[115] ^ D[113] ^ D[111] ^ D[109] ^ 
                 D[105] ^ D[104] ^ D[103] ^ D[102] ^ D[100] ^ D[98] ^ 
                 D[97] ^ D[96] ^ D[93] ^ D[91] ^ D[90] ^ D[89] ^ D[88] ^ 
                 D[87] ^ D[86] ^ D[85] ^ D[84] ^ D[82] ^ D[81] ^ D[80] ^ 
                 D[79] ^ D[75] ^ D[74] ^ D[73] ^ D[72] ^ D[69] ^ D[65] ^ 
                 D[62] ^ D[60] ^ D[59] ^ D[56] ^ D[55] ^ D[54] ^ D[50] ^ 
                 D[49] ^ D[47] ^ D[46] ^ D[42] ^ D[39] ^ D[38] ^ D[36] ^ 
                 D[35] ^ D[34] ^ D[31] ^ D[29] ^ D[27] ^ D[26] ^ D[20] ^ 
                 D[19] ^ D[17] ^ D[16] ^ D[15] ^ D[13] ^ D[9] ^ D[6] ^ 
                 D[1] ^ D[0] ^ C[0] ^ C[1] ^ C[2] ^ C[4] ^ C[6] ^ C[7] ^ 
                 C[8] ^ C[9] ^ C[13] ^ C[15] ^ C[17] ^ C[19] ^ C[21] ^ 
                 C[22] ^ C[23] ^ C[24] ^ C[26] ^ C[28] ^ C[30] ^ C[31];
    NewCRC[24] = D[127] ^ D[125] ^ D[123] ^ D[121] ^ D[120] ^ D[119] ^ 
                 D[118] ^ D[116] ^ D[114] ^ D[112] ^ D[110] ^ D[106] ^ 
                 D[105] ^ D[104] ^ D[103] ^ D[101] ^ D[99] ^ D[98] ^ 
                 D[97] ^ D[94] ^ D[92] ^ D[91] ^ D[90] ^ D[89] ^ D[88] ^ 
                 D[87] ^ D[86] ^ D[85] ^ D[83] ^ D[82] ^ D[81] ^ D[80] ^ 
                 D[76] ^ D[75] ^ D[74] ^ D[73] ^ D[70] ^ D[66] ^ D[63] ^ 
                 D[61] ^ D[60] ^ D[57] ^ D[56] ^ D[55] ^ D[51] ^ D[50] ^ 
                 D[48] ^ D[47] ^ D[43] ^ D[40] ^ D[39] ^ D[37] ^ D[36] ^ 
                 D[35] ^ D[32] ^ D[30] ^ D[28] ^ D[27] ^ D[21] ^ D[20] ^ 
                 D[18] ^ D[17] ^ D[16] ^ D[14] ^ D[10] ^ D[7] ^ D[2] ^ 
                 D[1] ^ C[1] ^ C[2] ^ C[3] ^ C[5] ^ C[7] ^ C[8] ^ C[9] ^ 
                 C[10] ^ C[14] ^ C[16] ^ C[18] ^ C[20] ^ C[22] ^ C[23] ^ 
                 C[24] ^ C[25] ^ C[27] ^ C[29] ^ C[31];
    NewCRC[25] = D[126] ^ D[124] ^ D[122] ^ D[121] ^ D[120] ^ D[119] ^ 
                 D[117] ^ D[115] ^ D[113] ^ D[111] ^ D[107] ^ D[106] ^ 
                 D[105] ^ D[104] ^ D[102] ^ D[100] ^ D[99] ^ D[98] ^ 
                 D[95] ^ D[93] ^ D[92] ^ D[91] ^ D[90] ^ D[89] ^ D[88] ^ 
                 D[87] ^ D[86] ^ D[84] ^ D[83] ^ D[82] ^ D[81] ^ D[77] ^ 
                 D[76] ^ D[75] ^ D[74] ^ D[71] ^ D[67] ^ D[64] ^ D[62] ^ 
                 D[61] ^ D[58] ^ D[57] ^ D[56] ^ D[52] ^ D[51] ^ D[49] ^ 
                 D[48] ^ D[44] ^ D[41] ^ D[40] ^ D[38] ^ D[37] ^ D[36] ^ 
                 D[33] ^ D[31] ^ D[29] ^ D[28] ^ D[22] ^ D[21] ^ D[19] ^ 
                 D[18] ^ D[17] ^ D[15] ^ D[11] ^ D[8] ^ D[3] ^ D[2] ^ 
                 C[2] ^ C[3] ^ C[4] ^ C[6] ^ C[8] ^ C[9] ^ C[10] ^ C[11] ^ 
                 C[15] ^ C[17] ^ C[19] ^ C[21] ^ C[23] ^ C[24] ^ C[25] ^ 
                 C[26] ^ C[28] ^ C[30];
    NewCRC[26] = D[126] ^ D[122] ^ D[121] ^ D[120] ^ D[119] ^ D[117] ^ 
                 D[113] ^ D[112] ^ D[111] ^ D[110] ^ D[108] ^ D[107] ^ 
                 D[105] ^ D[104] ^ D[100] ^ D[98] ^ D[97] ^ D[95] ^ 
                 D[93] ^ D[92] ^ D[91] ^ D[90] ^ D[89] ^ D[88] ^ D[81] ^ 
                 D[79] ^ D[78] ^ D[77] ^ D[76] ^ D[75] ^ D[73] ^ D[67] ^ 
                 D[66] ^ D[62] ^ D[61] ^ D[60] ^ D[59] ^ D[57] ^ D[55] ^ 
                 D[54] ^ D[52] ^ D[49] ^ D[48] ^ D[47] ^ D[44] ^ D[42] ^ 
                 D[41] ^ D[39] ^ D[38] ^ D[31] ^ D[28] ^ D[26] ^ D[25] ^ 
                 D[24] ^ D[23] ^ D[22] ^ D[20] ^ D[19] ^ D[18] ^ D[10] ^ 
                 D[6] ^ D[4] ^ D[3] ^ D[0] ^ C[1] ^ C[2] ^ C[4] ^ C[8] ^ 
                 C[9] ^ C[11] ^ C[12] ^ C[14] ^ C[15] ^ C[16] ^ C[17] ^ 
                 C[21] ^ C[23] ^ C[24] ^ C[25] ^ C[26] ^ C[30];
    NewCRC[27] = D[127] ^ D[123] ^ D[122] ^ D[121] ^ D[120] ^ D[118] ^ 
                 D[114] ^ D[113] ^ D[112] ^ D[111] ^ D[109] ^ D[108] ^ 
                 D[106] ^ D[105] ^ D[101] ^ D[99] ^ D[98] ^ D[96] ^ 
                 D[94] ^ D[93] ^ D[92] ^ D[91] ^ D[90] ^ D[89] ^ D[82] ^ 
                 D[80] ^ D[79] ^ D[78] ^ D[77] ^ D[76] ^ D[74] ^ D[68] ^ 
                 D[67] ^ D[63] ^ D[62] ^ D[61] ^ D[60] ^ D[58] ^ D[56] ^ 
                 D[55] ^ D[53] ^ D[50] ^ D[49] ^ D[48] ^ D[45] ^ D[43] ^ 
                 D[42] ^ D[40] ^ D[39] ^ D[32] ^ D[29] ^ D[27] ^ D[26] ^ 
                 D[25] ^ D[24] ^ D[23] ^ D[21] ^ D[20] ^ D[19] ^ D[11] ^ 
                 D[7] ^ D[5] ^ D[4] ^ D[1] ^ C[0] ^ C[2] ^ C[3] ^ C[5] ^ 
                 C[9] ^ C[10] ^ C[12] ^ C[13] ^ C[15] ^ C[16] ^ C[17] ^ 
                 C[18] ^ C[22] ^ C[24] ^ C[25] ^ C[26] ^ C[27] ^ C[31];
    NewCRC[28] = D[124] ^ D[123] ^ D[122] ^ D[121] ^ D[119] ^ D[115] ^ 
                 D[114] ^ D[113] ^ D[112] ^ D[110] ^ D[109] ^ D[107] ^ 
                 D[106] ^ D[102] ^ D[100] ^ D[99] ^ D[97] ^ D[95] ^ 
                 D[94] ^ D[93] ^ D[92] ^ D[91] ^ D[90] ^ D[83] ^ D[81] ^ 
                 D[80] ^ D[79] ^ D[78] ^ D[77] ^ D[75] ^ D[69] ^ D[68] ^ 
                 D[64] ^ D[63] ^ D[62] ^ D[61] ^ D[59] ^ D[57] ^ D[56] ^ 
                 D[54] ^ D[51] ^ D[50] ^ D[49] ^ D[46] ^ D[44] ^ D[43] ^ 
                 D[41] ^ D[40] ^ D[33] ^ D[30] ^ D[28] ^ D[27] ^ D[26] ^ 
                 D[25] ^ D[24] ^ D[22] ^ D[21] ^ D[20] ^ D[12] ^ D[8] ^ 
                 D[6] ^ D[5] ^ D[2] ^ C[1] ^ C[3] ^ C[4] ^ C[6] ^ C[10] ^ 
                 C[11] ^ C[13] ^ C[14] ^ C[16] ^ C[17] ^ C[18] ^ C[19] ^ 
                 C[23] ^ C[25] ^ C[26] ^ C[27] ^ C[28];
    NewCRC[29] = D[125] ^ D[124] ^ D[123] ^ D[122] ^ D[120] ^ D[116] ^ 
                 D[115] ^ D[114] ^ D[113] ^ D[111] ^ D[110] ^ D[108] ^ 
                 D[107] ^ D[103] ^ D[101] ^ D[100] ^ D[98] ^ D[96] ^ 
                 D[95] ^ D[94] ^ D[93] ^ D[92] ^ D[91] ^ D[84] ^ D[82] ^ 
                 D[81] ^ D[80] ^ D[79] ^ D[78] ^ D[76] ^ D[70] ^ D[69] ^ 
                 D[65] ^ D[64] ^ D[63] ^ D[62] ^ D[60] ^ D[58] ^ D[57] ^ 
                 D[55] ^ D[52] ^ D[51] ^ D[50] ^ D[47] ^ D[45] ^ D[44] ^ 
                 D[42] ^ D[41] ^ D[34] ^ D[31] ^ D[29] ^ D[28] ^ D[27] ^ 
                 D[26] ^ D[25] ^ D[23] ^ D[22] ^ D[21] ^ D[13] ^ D[9] ^ 
                 D[7] ^ D[6] ^ D[3] ^ C[0] ^ C[2] ^ C[4] ^ C[5] ^ C[7] ^ 
                 C[11] ^ C[12] ^ C[14] ^ C[15] ^ C[17] ^ C[18] ^ C[19] ^ 
                 C[20] ^ C[24] ^ C[26] ^ C[27] ^ C[28] ^ C[29];
    NewCRC[30] = D[126] ^ D[125] ^ D[124] ^ D[123] ^ D[121] ^ D[117] ^ 
                 D[116] ^ D[115] ^ D[114] ^ D[112] ^ D[111] ^ D[109] ^ 
                 D[108] ^ D[104] ^ D[102] ^ D[101] ^ D[99] ^ D[97] ^ 
                 D[96] ^ D[95] ^ D[94] ^ D[93] ^ D[92] ^ D[85] ^ D[83] ^ 
                 D[82] ^ D[81] ^ D[80] ^ D[79] ^ D[77] ^ D[71] ^ D[70] ^ 
                 D[66] ^ D[65] ^ D[64] ^ D[63] ^ D[61] ^ D[59] ^ D[58] ^ 
                 D[56] ^ D[53] ^ D[52] ^ D[51] ^ D[48] ^ D[46] ^ D[45] ^ 
                 D[43] ^ D[42] ^ D[35] ^ D[32] ^ D[30] ^ D[29] ^ D[28] ^ 
                 D[27] ^ D[26] ^ D[24] ^ D[23] ^ D[22] ^ D[14] ^ D[10] ^ 
                 D[8] ^ D[7] ^ D[4] ^ C[0] ^ C[1] ^ C[3] ^ C[5] ^ C[6] ^ 
                 C[8] ^ C[12] ^ C[13] ^ C[15] ^ C[16] ^ C[18] ^ C[19] ^ 
                 C[20] ^ C[21] ^ C[25] ^ C[27] ^ C[28] ^ C[29] ^ C[30];
    NewCRC[31] = D[127] ^ D[126] ^ D[125] ^ D[124] ^ D[122] ^ D[118] ^ 
                 D[117] ^ D[116] ^ D[115] ^ D[113] ^ D[112] ^ D[110] ^ 
                 D[109] ^ D[105] ^ D[103] ^ D[102] ^ D[100] ^ D[98] ^ 
                 D[97] ^ D[96] ^ D[95] ^ D[94] ^ D[93] ^ D[86] ^ D[84] ^ 
                 D[83] ^ D[82] ^ D[81] ^ D[80] ^ D[78] ^ D[72] ^ D[71] ^ 
                 D[67] ^ D[66] ^ D[65] ^ D[64] ^ D[62] ^ D[60] ^ D[59] ^ 
                 D[57] ^ D[54] ^ D[53] ^ D[52] ^ D[49] ^ D[47] ^ D[46] ^ 
                 D[44] ^ D[43] ^ D[36] ^ D[33] ^ D[31] ^ D[30] ^ D[29] ^ 
                 D[28] ^ D[27] ^ D[25] ^ D[24] ^ D[23] ^ D[15] ^ D[11] ^ 
                 D[9] ^ D[8] ^ D[5] ^ C[0] ^ C[1] ^ C[2] ^ C[4] ^ C[6] ^ 
                 C[7] ^ C[9] ^ C[13] ^ C[14] ^ C[16] ^ C[17] ^ C[19] ^ 
                 C[20] ^ C[21] ^ C[22] ^ C[26] ^ C[28] ^ C[29] ^ C[30] ^ 
                 C[31];

    nextCRC32_D128 = NewCRC;

  end

  endfunction
