`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hQykim29IynKQNLJGHNP1nO4iSRI+HDJ2HJQHF4ZRdjA469XtOc1teMiBGo3Vmdc
vv0STnAH7K8h0kqdJdEgCiHNpBTdXGWCMzNAsNfSVrcWM5ZnpJfHx8ZC0JbUznot
WZ+AZBCYmVHWc4Uskwy3+002g8eQ5IoGLqA7IDJzlgI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
t9Lepwt1imjy/t7oFYqxPhp9UgCL6/86dZTpxhlXewXEqRYncJI0jX8utNb410aK
4D0euCahkuxMmq3rhpBScrHtNEmpBX2CDYkLXjTtBsqWzO9w+V7K5vWOsJQjINpt
703ugYlWR4cj4hIR1m9+UV9F5oY/TQm3bS8GheKriUtcG5rG/4i3YaFQZgnyHzYA
mJmOQlWlD8eItWcVZv9T0RQBGYDbiLJCER6opTGnMZUXpYp4MgBqBsl6uzGkPO+e
Zo9UMOSLz+Suah6mDguW9ps1H58P9VLiVO+xdKiW4BPcXG6tGdpJTSROWEMlpTe3
REsAMrHwWIhk1QpC85dBITNyYG2S0sATSoOnlt7o/IbtU8RMKylmTIkzHbpdQCtQ
FKS7v1PaA6GLig/2VC8DyEDOPkv6CLJmKJcwu+Cf5SE44LoXQ2pTQ7H11S0HTCeM
chn4TO5ZIttCUVW/OxRe6/xPsluR/EgNQpvaW22EFvWJCvt893RrXMpaA4vxU9fg
/y5Z8S8f1qbRfMKCPrCyYA2z6qyqEdH/UMcGAOYUoranXN8TbD6BxdMc9qvvHA9Z
jLHRvGXu5QDly6IoI5bWTtNxnf3UsNk/TlcX+W0BTWl598MCkbkVdgE5mb8mTyoM
0OSzzhe2CIam+3dfOHSMS5L549tkz38H+zj4H4ZVzQJpnE5FKf7tLOtYcl3LHl1u
e1mxgGe99vUoN92cWLPIsM/uhE5MkpgcsyYxn07b9DoYUUU4cXxi91jCX9msgfYb
upS6vwVAB4nCGgmoep/CpiaWW623LuMA1HWHmW+1D4e5YGPkd4sztJFb6Gl2fnuW
I8RYQWgT7p5jey3R/qx4iAcR1PTzFc5oW+AbAtSH9bWYW/InjOHoTDoghapFwhvI
VPHRBa6wuRFQV9f0NH93Er0pT7gvXLqNjY+OK38HWQptvDPfoOZM4QTS26n+8WgL
OYPFAzrq/eNKeDnl8HO8rN4WWs9Qni1jKvdndU0M99qXMTiDJJw95gTHjQLbJwkd
OwQqdnedAwIjGVGCIcKVFVBwzOje/Gq85FzeSWsDGU+p+IigYfPucPOqk+ufa5HU
kErZ4PA+kWr9mVzOw86W7M4VwSZEnE/Bwi4R/QJIjEimktyc2KKxodj/jxhmd5uO
8uHWgEvV9XvkaObDV6IOtVaVEgz7IMbG7lixJeYesFrWkp/ju9W2zX42OF3Nt0L5
7k6qJwuxKf6jM3zWZA8B9hWaid5f1d711xNy+LPt+pWETnlGRj+cpzuVNCnUxoHb
hztZ7DHiySOavXyN3DEOI2nVHm2K4B7RiqIM/ljzwGauR8PfO20zuBEwSOet5M8V
ufJB0xcWIx0YyJA+rRqV7XsYD9ksqjXhQF6eGbBs2GYWu8JDxMDOBjvmvI0iefD1
UoB5e4eAZO5Ox44IT+kWN9u1eOyNyGWbZNVdIN/bVTUZgJ1nlDfmibJsH8sC3KYd
sd/Y1W8kOCrdjAiUO3zjMU4AsP6GKvSkgqRSID59uAaEvcEC3ubutmIPbzQ+vJIh
lSJx0owXJpkkH7AJ7zDC/Dhzpoen3CzgIYt6ossuqFEEKPT6sdUgSkLotrjQiu+E
nr0fS2QP1hfXZOOO5Ny9oG2Pi1LBeOhlLcqZI/qIsuB01LxJmwWkN+SgnidwaMcJ
stHOKk0BJKsxhT3TzKCiMUfhkmr1VFByUgQM618P79SQJ7O6Yk0bg9gETkGMhjSD
1HGIXQE28iqzBG1Ax+dJsZm/EimnFQCnbO88TZPCtV9/0KbHQU5n1UhpDEaqhrRZ
vu9KvYDGoaobGuuWYFM2D7ebtf7vuyK1CJjLDBs6nkRfogH0HDOlUC08Na7jz/wh
0OFXhqpyT5XSdCIx257pcxo5OmE/Wx/3C7SEt0C2l3JKq9MNipch21XA6EKlT3mz
hwmcKfjbVxZN2ylEa+jb41GNHFcGjbI2g9q4XvWEZN2qJ86rJZYTJvFWgu8Rt6A4
c5y5TZcDyQJvxlEBR0er34j/aLrrkVk9bkCQkGhRakhZvrbyGhEM8mQ1toz5tcTz
mh94u2FENU5/csxXbqsHluQpdtnBjsgkLyUmU7uosCZ58deGyNkgQ2R/WHxOhEST
pnG0oRYsB9tXVDfTe7RpRCzEaxm4XoaB5syhLzZcEZnNEqRQIBjT3sRFwh0ZOL8c
t1wUM+Q5tYlpLbVZOnKrGUKJfwuyYCRk0SAR2eD5CAEV38B5z95B+OMaCHu/Tl9O
A4STVoz14YEs6wNxuupe891Y7v/6zPZBAv0jHhaAPTQwU35QajcMQEqVV29Q/mV/
4LDxYETbslyTBr94dPEcPZOAB/EoEfVO1e+5NdHZTa5b6SvRXeJ0vK5Pp6btdoa7
wplS+YOpjAb0YG0VEj+UwEH89PsuTjhukkLM7Q9xNYDH2O1Yp5pwPLjXzApuJWT5
rX2GQvXC/7VsFf5/sud7yM+lfmRoEYdFs3N+erVNeoTUab+325yYmCZw+O6MTno3
kDIeaLCo7t8vYmFl7es/A8XxtK1N2g3f+kapOd2Q3N6jeQ6tJMuAgti+BMNogO+G
fuftPa7H1RkpdYEZoT3RM0SAWTDshqmTONxYK4eKQIDTg74hUENhuAj+TyaMb4Ug
K+6aREyToml/zswr3pvK7D7RAWI93IxQYmGJNa3GLMpzRW3P86ZoVS7IqBRHalYc
jwopN3ifwTEbse2xp2r41zIMcr+l1hV3niEvEkarCK1p1tbzV8MyYDsXJMNsnREM
9b1U5S/z0fX3oACGYlU42mvhYN2wKt2U2gNSnotirQBrrQ+NY7J1c4mSSQwg3Ub2
MoeJK+FRjDUAtKkYGcqQghxqvuX05iZGhJGOtBaebFKCE87kCJUa2AiTFVm0IX5f
G1Tqzbm1NusZ/FpT/PigBUmSSlTgXi7CqU+FEWREOI3mRszGU8KozvgwnXoqFyAx
Dt/yGaW0aD8tON+eLosA9AkgEU9frDcMx7uQ1dq8S7veGMLQsB2+XcIH+5d+xUkm
eQPHDJ8mofkKbl4q64PhM5O954Grx9XpM1gvpeKM5+nrfjLG/UWJbC9oQrj/HFdj
JDw6SLElob3yz7srEiXDPq5gBTIIMIa+W9XW/DIetBNau7S5Xa6dy8f2++aTNVrD
MZm7tJLB4M+faF3H/8tnFRmmT7y2jI2k0xwrmmI8B/mUvPtCSKT1740iq/DtpfVg
+zr82P+vIvg6WZrQaDlkFPoPY3+aXsupRaI7WGlImU4UZjL6ZG51w/Hbunfdymob
6C5Q98YLJSTHBuTMokMDt0Hii4JTkVBbmPO4mJtzJKNp5Hpajz0m90aYDhV85Zu9
fwemC/XEGBXEDmUsD6eSHOxZjRQcxZDVLpUOcyOl+VmNbiJ7kSk4LgLWuN+VwDzQ
4PKXKBcxvSpi16MzCQvFHBh1Yk6+/h85/thqFl4wPBKWvV9KCM0MLKs6q3P8FP4A
jQ2wEwX7gtIs7hWdeul8g9a37vx02puB7JXbHFUtI7j58PtdJZNaSTYvxyCNkY54
+/aOX7VpJt25zdJxiXAf+IcU46AVF03cdAOuPI2xeCaI6I6GUoZfjCMR7fzPA1hR
Up1m8/WSOsiArHtgsdt7qNlqVzUB5VPNGrEvw1355/8AV7thO48IQrylWoP+FPgq
gJgfdtDk5t9BKrCuN7YJfCjFmiwmc/+AJIbjQHur6/rXmmG2hoLAiBxEOqDyk4hH
+j7rYtJ4g4fTDqudVqhhDya+5s3HgyvkBYD+P8dwOoKC11E9Oevw8cfu7CdXtoDd
EUsf2QuM0G4l5l/ZA2Rec2utpm0/IM9uvo6T29adphLQGCtFTh+KIO9PBPJcETA7
XdT5iWsyFXLvIa7Gecr0+xdJX2kUrMIlR6843cJl0ioulro2HrVV0AyWyi6AQVwe
SLS256VTewRwPkwrUykNPIR3UEbv814cblFtBTZIfI9o0mN9I0gVlSPp3H9Tpicx
4sCjeQ+ZmZ4SZAqc8Kr5MUzMzGOtniqt8GxznyMun12LjxRIBS/oVw+HwUmFIMeY
zCK0j8Wd5L2qT7hmP5f0FHWen7sIhk1c1nO2K6WU302Ea/JwrHMwZkyQ5UXiCSaQ
YaHaS6dSZn6ZndR0HmuIjBRHMz1jWGqpF6xLT9teQ7zbgq0eO8v30yBfTZ0EaJY2
oc3fnwcaHyuslJqu3mmvbLa7JfhAQipTCB4p0XJe3KmZ4FdonmD9ADeMRWmhJYmY
n/PaRDcFWof6Xu+sFq3p2IW8vsG+GZJjTdBvmHj6c2RrXtx3n/+IYedMn0rXbWyX
FNcvtA/vLZW2YCf/O75Z0XWENaRyP5f08VviesSCZe5IsoM67QtrxWo1RA2+k3VK
Fqg0oT/AdorNOOPZuN1JeDOocd9E7Ogf0BCySl5jwLkITAB2djrY4tqwrVzfxCCz
fh/DO4YBsA4iRgDTCL8JOVFxEbMK5rSNVZpy+UvGhl6Vg737TLtlHYeEkqt6VqwO
kplCaa+LIdQ+eF0SOdi6Q4LPqgrLv7WbD2mvAneBZFSev5YLMRrnUiZndpIVpmF6
bUaTO41plQtUONLoI/mkDDf100H2CTHg6nFxIuTy5SCdoJG81dw+yj3m7WbNAO1C
8S2hguxdoMxyxLZoyho5JmQt1TFObQwxY3umUg6axK1gwE+HRjm3IQ+UkS5t8KzQ
/VTlq85tFAUKbMvWJQn6H+WaFT0ohky+TJbJcgtPufdh7aWpq3lW72cX1Wk0JXdq
Qz8fjRTmKMgLAHiTj3UQ9F3tGPw4MjlSZ2fRe52d/PijLkdGSN21KzDkyFPKR47b
8Sbdd7AzLpohUisui+Ly836MhCYsaMFUAxUZzwYVhemPOv2qgTY849yHTMjcJIFy
3Cn9d4XJjdE+AUGQfPaoWOk36Deq/VbiN9uN0dvf2UcITnwHoZf9Huga/3Ql0Hfi
gNfpHZ4YwzYUZGhCjgCIvUv8X4JWwqtSinjjFEsSunmc61w36GreUNgKcr5G8YaS
UaFMtX33/UXhhc/6qk7+HU+SqKKwWGzc6Ui9UwVWMLx/6tpm5+gzHKSKLTMn6v/8
AHz7RN3C5OfRiEuFLx4Gbh0IB+S9g5gvqfVgRl/yA3mcO9WKmctwzIt1G4Yi2ppm
4bgH+H8OkOnhoxMM6SD+6NsD4vTKzyjqXvFtDrpu9CUR0SccCB564lM2H+M0fXtj
qfCZeqZ050C2v1y4phBTHS6xYp3P1HT3PqcPftAkJQy8uyd3W2vZeuJ+FfCD9ReC
YXw53JoCz5YSaPyAuHaTiNReO511NG5XVLU7wLBh1p5CUQlLHcLT1pW8eQf7oeKL
AB71faOyAYXp9QRiSElIKSpQDCAcEc0vJgcszlbVHe4MFy+C6vQYy/Z/YiMBQ6EL
jCEXYFmpOWmcqRC9MdEXp4rT1ZBJD5nIDAqE8ABN7H9zUFLE6K0Z1GeDU7zbR9OH
Y+u8YQ8wqgFyao21vVOzL7c0FBCS1GOzR3kGlrcOcDmlO3THS6RgAQH2F7cxhntj
R0urXr5x3Wsn+JA5IaDzVk7T2bBl4E45f+CGiiDh+xpM5fD81gv7vCh8QaGzUbGN
xxv31huQAiinWlZGwZXhQshThPBosit0Rf2OOv4cALNiNp+LtJCEV4gVq8NvUaGU
xtT6guMBE+6Kgha8MMbDdSKu3W3MxQPoBG4DekEwhmMVu47VSlorDqykzxIa1J4l
t5qGBoQroklFTbozjk6SqBm84A+M2wtXM51l5b8/rZLszJQEjWEk4tEpN4n25VBQ
DnjRuEhHp5VbrlTGao3XBAcRvjnNIKayAQ5T8AtDbNgPJG7dyY9YODd7/jGGkRvK
Xuj0ovMOCEKFHizABQy2eJHZp/rJUxAeZjmCB8Nkj20HwN+60lV1GyWNQouWlE2x
5M47IoXjVWdkhczDrdkIvp1iPlEyANbRaBqQoJsiD+2OTqVZ3niet2pyTWD87bRS
6HUJRnt3iPX+gIfWbzKVAZRqERsyBmSYwB4vZY2Jwgur1XywnqoSmpmsVWTOusle
7oskzXmAXVFYpd6zBBMU2k3NXXMImbOXHsggBiOjeVXFaoKZAcri+f/7E/dpMQQq
RwD3NVOIVU0O91UEsuCsA8cx0thInEjYlaecgXmRwoOJuQeIDzS9S15EZoafbv3M
SC/wss2PdN96mHtyzCTHlrMWNOiMmO3ObP/XJAf7NclFPdOyAD/QZgALONXiJwfn
dWejy14wMPAb2h8vYvdwga2uA24FvEVAO2GY2jeo7e3Q2w0Utv5sJNC5uD8dWP0+
L6HgkGBtig7fUclwCy2WXAXDIExwzMQk2cVTziVD3QIwqK9xKLFds6Sj8GJXg+P+
Jet2ubNBiIxhekBAPYHKQPIJtzeqPk1xsxBQN0LDceEycUc7XQiB8aG4snmPBu8D
4yPnOwqH5bo13x8JjM5skCl2qglDf7sXDKesOwB12ov+TFf+J4cCTF9eo/NM0W8J
XF7NRIQ/CJZVrNpU0Uy5gJ4nlD7GjeRzeAkTOoTayMX8RUr6tn+vDItnpEjAMZ4Q
O0ChF2jJEKhx4TfAUf5i243aZerQyYWQOAUoMJqX2LNAUZvDrQi+PsKCT36l+XLc
XytlO6kDW9AyN/CAprdDrE01topNpdo4lO9wK2Xog+JDeM06IENL6wMcAwkbw1u6
YFhl6aH0o1Xo/6ex3dZNkEnzcRhd25Ze9qIxfEFS74aG32yP7ZXHkW6hZassBhXM
l85t0wj6EImdHmPYJh3625e6YuNrYjKLZs/SSdy5N6mVcejQ6rrqELogd3+n3dO1
G3q/295AMxgGOJCD6xDFuswoukgVUq58w78PefRY5xV/+3VyVC4wdHGduiqZ4Jy3
hAmJoK4jJCpHcUv8a8pPVcswXRB2m5ERUusbcMUT9OgvptYkvNuCyZocEaQ0olOY
aPXPQmKVmbvDn40OV4Lya7QGnsSKYDkml/K7vBORSTGdn+5Oq/60QjK/Y/765iTl
twFaKPWAmvTkVNNEJ4cBXfojeWTpvx6PZz/AJUAwmMSP5dzEHrPKE1FBmMJ/MhW8
zTA9qKbUKXRotwjKaBXzRxpzTpeH0Kyz7qcBppYa8g1SlgcfBOwqutZRDrNgCKtE
H/D1I6yZ31RPTyvN2pCHYv44TyeZq2Il9c/SCYe0H05jPUtf21cWXZr6+QdjN7un
7/J6AFSL5lFhclTZa6azRyDWDKxcqEknYe75l4GT6gfAogvvF2LDfA5J/wyYisIp
z7hBbIelxvVz/UPBOqW3+H0IiCIwih5VT65tXJZkgTPhDHDanzHcd/Qm1ah9KqUU
O7HnC2RFX1K8kEgHe3itKRq5odq07As6ragbn/smxbBF3psK6hvyeQza9Bbsp2IQ
NGz2DmVHFo367IyNtx6QOasGZHsfbPSqrFz59A3hANNRzZuMqrjUvp5+zAAajres
+SfSO5WP1pQ7bgSXF6TzWu2hT5S6cRKPE03AkOaMu79t+Haz2mN+TjtpA8rrvJUR
iA2Zb5kSlzinzeEGRyZYsyak2IijL4r86lSrwMaL1XaJvytVVnEFAPINLrPlDi4O
GnGEbs9GDsOgZxGSE2+8SfYrJFYcdrutsKZkSwVeo21IExLlhkWUfxU69nT8wJBj
NCn9Yylvsu39U8UtnnkFP/0zls/wmUIT+tfVLNiMULgwqeDP01UZmTNixB4VTkvm
CaTUsbbZ5RxZgt0Nzaehu3xjI7RWk1GnWL1B/fQ7MbRS1Us5bLX5EI2piziMfWlu
mOeUdEdEDiFXDtjFm4xklwlyzvkJFLKirKWI2ErO7DEffIg0MpklfNUC0Dr52xV0
bAC6GcTDBjOlRIj/3BfiVNmOkCI0uIdu5TZInHwjlVoNtcOHKoeE8LQpXEFGbfCF
SPR8FSBHzHP9Vfr2FSwje6Ql7xkHWQHhmyOAs16vWdEJtXgI1NZVr0igrOuCXRvh
K9y+SCdzrXnHJS0w1MJaRD8jalrAZ4ys9W1y9MkYCAAKY4M0r7ye5U6lV+BF8k9z
YF5D7uoRfkhAqfgecsYXivYr/lKe8v8aTof5fFIlKGySME49K2pYjXj1RkFTp3Co
qG+Ww8e3hX1r8B0n+5OTQTz8MXftAHjJ+vIZXUBA5RjI8rRtSVQNPnVYCOEWyxPQ
o/RvSbCTVbywwIySF+SsAlsMIH1+1SdQ6dqrL9JDjh6F+L7J4Mz2mAENVwXhzMcb
TZJg7kJz2Q0LtozwQfnF02dMkd5x7apVi9euyLDCozsu0Z2tixQfxIMaf7nQa41m
5R7Y5pHvUJyY13PZ+hMz6j1eEvig4cE34m/W4Ixf6FJbHv7Swwb9XyxVi4cvEojK
tDAJgna2JE7rnM8ohsPx+bvAIhGDhvC/u4cFtVrbuxilc/005VQOgZQeHTgguU8D
0UaYK9GYbcDzsg4A0mCCuZGZIbDg/rWQLSdqfAWu6kNEnnh5mPvX6A6eiPCyt89Z
FmOJnX1Oa7mN4yGhN+74OXpOOfdWe1qkkPOuzN2Jh9rs42hdW7yTVo8VuQ9Mdrbm
rW71YG6uXaPVcwntyWDyLn9M9+dHyVe5pfv7AgVzQPb6niyS65489neHIgxpW/QJ
jWCd0f320Y66YwPFGQGUSyjstfl6jh8/9eSpx8Yt1GlhqNg8rYC7UwEQ8oyo5HDk
i2v1hguNkJX1btR6KPUIN76FlD/s9BQT5u+gWKTUrXf3dtS/wh5u8Zp1BNlZdaij
EttdCLPqxjfmzYgoRRVFayInMQ70loXhYlpsIII5qPHoB4KoBJqGTl5joMhiYqNm
49DnbnuyV6YL7jQRuDrzTxTbIDc9daPvKq+wJnJvJL98qfED7eAcX//Drh3l6CUm
MDoadyxZGsuQLAybELRwCJHNCiRQWi/+jeq7+iBkdHXVxKdhCZeV8jfD/x99kRW9
T5XzudENXKu9I556rPJkAcL/HsXLQoO9vXBluiXSrtq46KsYqf1nEd/1wjl+ITuh
dzJgiqsOWh6l5UFqKMJulw06U0/Ak2RP4+WFsv6Bk45edeaT1z2gAry+toG5RNaN
Cau1tnk/twoWcrfWf5+U9F2sDO65rh7Q/MLTZmPLDV6Wxt6llCmsm42PZPhen44Y
1CGABrGXvk1S9rUkr6Nev1go/9yaCmYRTWyvs133xJmIrHR1lfaPN8kJjpD+mvyH
LRXslmWI1aVndIzCrrRXmj7TMNlU1y9PkVDe7iQHkn1ge/0GNrDru8n6RhyR7LnO
N+QWjaib7DWDRrEyppuM/beWrhuDj/shxTMyurz50pLfcMQOY1rEK80B9X6zt1Kz
eg224R2PyVwehaNRrncqddPsU51mUNh8cDiM36J7Fb1GhaCi5fHFcfQRNx0xOyx7
EIqcpJPi30UJ3zSAwDPwu+zvmIdlbXJiFfL1fMz0Lz+ycaAD09UDWS7DLz5g2+NN
zK8wYSs5w/AoW4t4YtoWvV8eTOtJ2xWfP0QGbw5f8N37aPDF++6Pp20ZbLClnt6d
EzVmEMmUqB+Ay6MvWxMoV6QWOn+Zcw/CMfAP9JzL11HvLzbHDQLckzy3Y8xW/kIi
YQXQ+tTeU1MQCBmq0qF2vN90O2zda+YPWfOBHK8SkLO7zc6V+U6/BUh6dgJ2taLu
M3IU4k7dfO6MJltJqpRQml5I9RW3tTau3DywiGhLb/Dt4qJOdquyHoxRBLJQchQQ
hQbdxyqwJcEuFZANnoMQVG/VroFwGIXmw7tFayMtM4n/xkfICqAduRK7fh8FDnAC
NPG7EZ3ANWPLAIZiCoIJCZpgDIU+t6dz6D1brrKoLiLeLVlytY8yaEd/QatS1c4j
C5L3XVZZJwjybGFue/PyV2LKb/pdwFkZnPPuT1bt/WZMC6jhtBYuvgqAJY1px7zG
j4ZRHpkaS0Bmf4Ubq/SfLte1i0bBbnmSU1mMlXfi7Z005i1pW2GInsAVo05TLUm0
Zeyc5+cJQHX6WWQN0TZdZCSMJ5X1tPy/QjagnJKabAzRsK0zDZ6j0ulKrlX3EszW
bJZKkOq6IXQzdGRxh7vzxbtfemGAyJ49RMIZaBmNpP5fKhoYXHS3Uqkwl+6/Uapu
ktrSFNtuDsc5TUux/dJXjuYmv65lu4m1QcFhH6/wfOUPMJIDzGh3IgkRhmy2tD3S
xfMpRaCUOmofijvaIkARI579RcXi7Q2+p/sbggAwIaHU+R5LNF/Rrv3cCUZxlr8F
1AVvdmFiTlbIg8nuYr86McZMwzajjIo5AbFKgYN6moGhzGO9VV+iJUh/Yt5vi4KJ
WV8giezKUpEz9JysWP61ncTOYmLbGGp1lvRLQiqsgWAzNdMBgjuK8h4+eLjWxBqa
HM9pVXNzat78/O6jxQW5GErB6/oEJ5Vg34FTixpFGca0a5iZcEJENe6ofMtwhdjO
nmg2iMNSIc4Egulw7M3Hy3OZ4QCy2SVygN7485iSwiHdmkSPlM5+JlXlkp1g6w3t
Ozxe89Z8y5NS3f2IK9thSJ76quQpI7926LGle14FtdgmFGaQ+/R398lzDL9IGFP/
B5dyhv795unZyBK0bw/ZP48eWfxJNXLzWJtF246SJ0UGUPX8KriNaH5F9y+t2tcJ
0lJ0qSOp0zf7cs1F6OkH6ndWt7lhsfoBmT6T4F+jxr56oaXt86lZTxhFG3hhSuQ2
0ntUsBSmfvRC2Hegz7p+SbyphT1cCc90IahtP+81pll8c2yBdgkwbx0FB2mrlCyx
Pbll4whptdrZb9guACZXUJwJnLFNfCIAk8qsyok4QnIgOC8J1fvidDnDjFOGnYkX
5Jzne7ScutyzZHyZT6X1Pvmu0YWt9xeewyBL03OxrZCpzPr74yJSCwFKxs2OYVZb
gyQACE6VYJQvwGs4+d3iJEfXJCwXfee72aVeKvHIMyBAoC8XoN4ZFuhWhTSWMhmc
jcQCeqv05qaVA9mzCZPulIbjJ0a3BgmqQ59A/Dfyhneqp0OUEOYQn9mvKktOCpFS
E8SQpcwP0ozMLUH7abKEHWm9cPjZCS4qZldf2UnAaYdfqkpjHvwKIx9Zaj4hwSQO
M73XY+NCXID5CbkmQwpTkdNpdAcrGUgaRuCpaTohd3ST/vwXXSRzCgSUUVOKIFEw
WjZfTUrkg1k8Y01sn5X2cquuRghonGpM2EnohTsDKA2onJJCouQGPmffkvJZAfoP
+GPbwUiL1tXy8oZ7jOFO5T7gI0p8v4NAmMU/yXtKGecpM1IcEm+2VsSyRrKRFXFx
5zPQh+JectAj+iOJytZ+3SgItXxFyGlScyHYhQeT2vnFlaZSfj2RsesqUj1lZtXl
GucszjdQ2C/13EIyu6pizjpzmTr/lk2IIgjtg3QZNB6jU1q5w/LJxx2F5hWvODgG
qFA2rjrqGesk+TBny5fTrSZewGqAiGMe8vAmSBjJP9UZPP1kw5Ulv0INlZiUc72a
h4F/eVOAWDSFk8apfTXefqm4dD3KkgGG/yzepLVCXj5MfhSnJe5Ie/gVc9bU/6Hj
ls8bo+RHQpa2FbNhGgI+sP76voR6i+HCfdrBNQ5GNNRjIhdX34UjrpYo9wLLJOkt
yBI4+O6BT3nYzAUGRkreyvuZo1BLvimjdJIuTop2VVFFN20sM0qXf/BWt/G17U3E
ztDA2jhdncVhrjHAN5qkrZ7SqEvsRw47J8JqYy2JJUFfiXDNvRZLIfVOL1v0b+PW
NT499BEHWV4BnftJf6XKlvJp+izws7jDwSEjRSVWWvSV1l61nxR2EHj7C8YehEzB
zmKFgzx6c6T/Uw9a65V0LyiGD5VL5ow+rbnEGTLAZ0pjXLXZHrYyKQZIjjh6rzcJ
972qisuZclki1qNSRrNC3U8DMSFpMGW1H70YAvqPrpjiTxKTQj3eII6YliVU9PIH
weBmiRD5B1VAzqAeaEbRBV9MkRFP02ySqpioKgMJq7XKbA2k2cV/lerk+uF2dhDD
ftVG1V80SzFn2xPnFZ+scMgL4K+4F2atfbesuiSmH31yA/RAiV2PlhVaOo9tGxCI
nP5F/UUtSlMzAcgQM+7tHgt1h/OGk82WvWLKM3AnG0Bq+OAxC2wXoi6oEVfslAM7
3575L/JGUc0hME6gZ/nH5zlzoG2h20SFm0ExBF+2Wj0gC+Q4b3PDG/APmBVzj2xx
D8bfJDlXbdynE7gCmCxiPC7lelHIkjnG/0ZvE6g+wQQ+9/Vz6NKan0fMSYS0pbSu
i9nT7S77yQ3rgokTdos0lSSfqBJKOuitVKIkrSvxgVeiNGspPFakddQ5MEPOiz0J
WPRVMbWMa0ljDNULvjVkloFqyiC9mkbyNe3QRpMo2nbfrjxq7BeBYG0WKiXz+m5R
H4SAPMk5hXwKE7UcFApTPevvVbIdHDj/did17hMo+8SsGBuC4TQq7NggJvEZ4a+T
3TIy8BGxHT2NrjDTkPxlIBRWzMf0o9yZuT2bZVbM1Ea4suaYUUJH1Zq7yHSg3wE0
U0/l0aSLdzuB5ogh3dcKrY0/D27X5tuieBEORU+qISBtyFaYWLIxUFAVLH/oAYSD
wriR00VlKvxM0zPwzpuUae9SaUI3mNwUs3Rfy3K6Qa2AvrKydyqKFP68AjtW2p33
u8qpNZjU1DWgZ/Wg3PgSREaIiYptRx6cS76yoYQB7lXfP9qC2dkl3xYyJD7DLAls
b8zQD+RgSGqq6fFYIeKjCJA7yyR41HFDajLQ/H9utShWeK8ydu7hxpFbXkiGpJq/
vRXiykBQsivaVf0t15hZyEnKyRlbT144NnxyXzfgFvU0ti+IhRUAP/nFC2JjgMGB
p1BDcgEhL1e3zmNGU94/2rqPbF4uJux0d8WwlWck5KYTn1aPQD5ffI67YnyZ6uyR
gJDqNBBbM03xxuzMm3adYZlJpNs05qkDOO4PoyrvgSFbede8i9TWTRhE533GuhJk
dB/Cvjm0X38vMLbY2qHQ2W8gaoBJIc6HPlt3/+5P7S3JmYJB1RE8hBGSgrbLu897
6GZ2iyNDJR0i/UcMfjWFvU67jr2+1cpRmpLtIetB/UQPAZv7qa6dp6tlkCQ0sZlB
TvJkq+jwz5ZwI2ClHQMfdMk5XKOGg83/2OKyLtNVFbVTcOQHjpUqwDknPWakF6kM
/mST0ggZkAVM0ZuDAR27jJl7JwwDQ4mt4JLDK5UTIvURWCUZlf7N9XiTcaxwC9mg
vf7xe2SNEcTgxZwIrqYq/SrJyKMKnB/D5eqHdbmK7/uaRsnIFgqt7b2uiLc5V2Um
NxtFIcXMhGtBe9x/M0+Dz/A+typpJXaW0T5TwtfYPFoskT68qRdoMOiuVBAP/opD
T7MoLYDZ5o9wAIKu51HksBGo2tVHerwbnlSZyZls8BmDs0T4g+KYaRTd7402shPd
UZKphoFuO5FGc9S2Hp5dDO64pSkvEkx6REAmaJeUsKBw3UyP4w7xQ+TvwCEUEEWt
Ai2k2fwIhrXZc/6qiv7BN+cveCy/JcSQyTglWTI6xjNnPvcrCzcPwk/FWxSMnw5C
kzjwwAJ3gVE0cV1uP0xMlPtFCifpOqHdYc5MNw48n/Sft6u8TI9kafxwSH6Wt3ky
ZiKmgEB68xIkNSjJ2BbSPYm10/918CDVXb2iHKP+/9CRBA9qBHLEPeiDKbojSBEc
/Cz9m3BQbORwcm024lqI+NMy1umXbFvPYiwh7g2O6HqKzpt+dJiYDE5599Ugpve0
+1JX6jzGPXkRZcH193QqLyyXlq7m00BxCzKNNDaq3hn4pi1BzFJu+yxoCWlkIT6I
5ybO5QdtPsCa8Ij6qvi72u6or2PBL+i4FDU4DFXgVJZcwJQEuhbBPeBMLRo6WJh5
XlI4eTY+in6F+B5+siYEenePByXZyRvb8WzQVTTI4phCOfJxnYH7JEVarEOZVnxz
32K3rszW37BabnYgrcNvZvVgGUZ9N8F3N2AnWMs/EMYhCLPbUemVAfUMN8fx9wbn
jJPyGO48BZ0tbYBKqei3ed8l2qq+6v3v6gDZECjN0gPMiwHL/4Lfqg7VsefZ6GJL
SY9R4KpFu6UhgpSIFrvDNayWVSgsHUxHqKbNQJ4g0f8EL+N1j4SgDPG39J9/oVfp
nI9ifDNZ4jN82EKhdzzQzQ==
`pragma protect end_protected
