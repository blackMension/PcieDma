module pll (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1, // outclk1.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);
endmodule

