`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QNR+NynscvcfNotB90UgBcWHea/YBGE+UYjLkja61W+YEq7AcWbbmZ9ZdnM9gY5y
Kd3RBSp93tzlEwIQT8Mra4E4cpUcRjD01h0q8Dms/ENWNhLuP8vcN8lqPcFCi0Vd
KMsPSaHVmHdMLMS8NkUjSt9brJ39b1FVc/1MNPqkyKo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809888)
TynGTnWFeHLzgjivgSTRlDfOkT293MsP64L91QdDc1WDYVn9aEB1q3IYlqPpN2o2
IIAAUfzsaHaCaw6xDqeK4YSPt7wZANkkVFLEqd7NUPLcgMHuh/Zz25+4dChzvYIA
nZOCIluZJ91zVlca14Ej5Ma4hq8ftpQt/qrulO33BKnX0O72QsA3Cg3XIaRuJfZ/
mFQjAbTagnxHf8HcfzchND5HlQFkrnsiUVlOXtoBr85ancONPySN+tI1B4xlWBDg
EXxfZQcfJK/OwqcrtCNsPJQClCuu09UpFZ4FRCZLTbYhn+Rgp8/zL0USf5IZNveH
jpm0lbIZQilB7jEF6W5l746jTLf9DUPoTgfQYZWJNYVi5QpZamiTmMOQOMnn4nCl
CGPWrsQKMbNpiunaTfToN4NGfMXsiSqsBjz3hp3mSvC4esh9bkdfmBBN61N2FXl6
w2dZWnHEAAnDb+5e0vziC1t/IH1sSTZL9VI9kl+nwBUXR9QgPE8BT3GZUZGCv/rD
smuJKUWWAqJHC40iw0ShZQ0lDTvVdLxWBYvb522qeH7+F0qSUhFAC6I724bYMcZp
u5VQ/br6emwFJZw+sbivs1XSHbRjffjdvTX+lBMVOqdi0c6xTt1XmNoQH+uEl12E
WILkB2Y9ZSb3uDnr2pfonxqPAWvy+t4z2kvUfbvdGIUdlMLssJ6xYZJYSsoS1599
0ePTj3No0RkVL+Pp3FDlcC6ZmVoNAVZhX2WNKltveTwFyFg/EPQ/aNtx++zbCKAF
ezJpoa10E41O7fdRwamTxL6hP8OWU9/7kcFpiUzIBf4MGNZGIawRnBgpn9VtD4a7
Wm9LsPQGDh0fYAg2SvCeDgtGDiUu3j3n0KCClmWtNyCftp61zIhAVVbwEVoNxnwo
SCHRVVfysTU+nqHydAf5VD3O1Zu2xnBzVJf6E4vOdgQj3JzwjkIqp1WMu8XawMpw
4QaQS41MACj9v1GOH8kp9WF9/inL3o0TtczdUDq47qws8JD2opRPDPxsFgrU2/EA
VdKHv2LpLWzD3uEi8dxgEnISGx+zQcy4ea2oWKFUtxC5uwNAvwPDOvcTw4far1mu
tLCxjI+ParbkgOSc9UE8CYc9mvjx1xPxMH9fWpAsJv8iCA4xCvh3UQxwmbXF7A39
3i6XjzAFDAbOd06RdTQrDzgisdw30IZvGNAhPIkg4ub8r8MqRZrAh7T+t+TCqm7Y
nNDMQs7L/H8OP/qwz+/hcEL8nz5qGRxxHscc31Sq73YdaODuzEBDi+0L2cDSC9mN
JDj/FD6FHagCR3/Uyh7D2KBQmEX8DmrfIs9cRAwpHdAHmtJy/HyYr9iaGjkvklMN
XK0M6jpxG4aT+IoVmKcOb4rDpus/RI9xsOFVjKmxy0Vm9ejAreZr5VYymsJbqQaE
IwY1PD4dFjPUpKfXUbuzaQuL9JR0IMQbmLcmXeGjE4hNRVBa44D8pQcDgGlGKNnB
KTu3IRmdtIjYHpS2DmqLem/5TGJSfBSfh2nvIOQkZE7A6enGIvrX6z+dSajxrvur
mp2IsR2tzRXLRfO/mbdu49KU2G0rC2rRCwX48Nj/SlBiNxpCWvjrZ/b7lIBKcV7K
3wV1BPLknjfEfygsijz+sZDKg8mNfpVCWlbKYTBZT1xM2+TvGEL6+IcASTw2iXZq
QCYYtQKUbbT+fuE5/pLTJhMTid0iadyPS+N0t5c8uy/xXhz7UnFmWcRGU7FmSNJE
ONAvTWXD2a5klPnBH11zpwupqKxOZEOfMq2k79cPu4XN2XcCBRBivY7HIjmPx/NJ
eelt5GlxZ2dXz6c8eEQ2rEVd05MOWyzZeUSR4CeajgpK7jS2Hs+l1W4rsYQfYvfr
FZHCw2x0FzoIfSoKeDwE2LdBXUoBPQr/nfi/IgCGrK0bd6jYsMvwDZP43Q/icE0/
XgbPCoG+j5p63PgsQV9rZvuLdEPJyaklC3KzAMvtPamo9e4B2vgyY4130z+Lp8dj
BYWKv+UuaRD7qo/5zQCBk8G+QS2F7z6J9Ta0sHL9AIvSZndlt/ciDE7RyWgOTIs5
ztLiNLwQjNhHraBUGYaE2XAl9S6Kal7VgvOpwSntwJP5yuFZ6FJpf18Aocni4sdA
JzYa4ZH4kRoeYjiBgWRwQ+k3iPWdmvPpWdphQV9XnavlPLv1pyqB51/uZmwP0BhR
pIs5YctZYr4+7LpV5yUWhEQYndPx7PWWHJ6soqdfS5i7N/EXc7Tm4/O31oazIGrG
gtj8uhcZQdiCGolvWiVet6iLZ8D3FKYnrTxctbGD2csePPxF+mZXCpmp46zzqNGS
zZaEpfisGjkoieDPcZ4Lsx+gB3w1aG+AOFeC5BdCkX2DOWw3i6RFaP2HLzrCmaVJ
WEufygC6MxYnOzfpl/KnjZoswlY743snPKtT/Etip1ob4oAkV3tQDqrVOujL5t+z
yBQEAWupnnBihSr5puEtNwgnyWcRTOYtsYSRdXyUCO/hy8Es0EtxXedsx63Es/wy
ZczOYHWaVsz7I+Xmtrp5hTBiA4cMqQuazLjcJutn9pvqsQ/xPp5JWf219lQeXsYa
cjqCoLRkiAkaMbL36aDzGbTlgX6sH98dd++6G6Q7gpJNPWR3N/n9RFn7EFk/bgbV
5HYhl71n4AoFsZZfxZqDzNYSRWdyl6rzz1Lw7KG1ObeQhHOcr7WDhK/HuPYHiwLM
jD//4NJZly0gimNXwClQ2HFtJLuXqPKieOxpWyCeyzSlrzc8xBHoxGJpzfwBp/Ls
uQ3fX79EYjjdLxbNPkVUU6nIMjEEXSWoNDlupmluueiSypNHC0KL8J8eTtgs6b9J
AwAW/g4NQdExM8kgM1EFOi/y8JzSeHtrqAQZOEguQ3noFdVDqJ/X6Eo2H+gzkv/c
DZbMmvf14oBXevowNYEB8J1pWa6iHfT7uIoZXFT4g1IPZkWV95mRdPQh6PzGA9bh
hLEa0GxIO6P+vzhaVvUUpltM5EIJcXQzlEyPeqIXzNxZ7ThVxSGo+2BNHD1cyv3C
YvKT6g6fjHxuPRepu18prsXFknDUVIxYFGlwWoFC4sGoCneAFOKNMS9BYysMVoA7
OC8F1som2k3SlESI336y+4CfY0PcByO7NQHnUfAQbMrsy23ThH9udknZUWr8aveg
nziTROdRVFtv72s3P9PQTZacoc1C7OWCSY7njkjo+1nlDfJ+hJfW+6PisyawonGB
ZdhgqD49FsIZ2GOlsaj595nmavUUA/GK3scfRJMdBHOqcFWnknZenvlCFOT7sKw1
JZ9yb/fElzZVZZPF4Wq0cVaUvhoH9c2D8+xvCUFB93YiR5RbA4M+qKhCUcB9tvVE
XifMlsdQkOibjV8vjnMV+JIXzBTiFwhsfyN3ksctZp1Qq5bjQQPIVNunC3XqHrs+
6plxHkaFVGVURuCCRhERjEWV7EbkMqcJT6VLSpF8Oo78sYNe8pTa6FBfeJ5r3FJS
e8eejfNSQxyABquZoN0CW6SBBcKmxyTE9Rxb7j5jXDTISq9gqg4qIPev4IGEIuXR
9e+Zw0hB311N7heYWuuUIPfXz/Fy32L0Yo8sLVGX50702+rmOapTaoqMaSNhz9Rc
yKSdYQCcY+OAWrg6x6H6vC2gBiDGpNiLB2x0iMtnO5kWXK4vfMcORZooSLYu+sbJ
nLqIR81fW95VXf/FE2tjD39NBWp6TVvjdKNu4S3figcveOt2kCJTpK15hXuhqvGa
9TEKuO0Rl4ENIeX6HS1GXHelNRdpAnEaR3hGy0mUhykZe7QVoByAUFKNWAxIbney
DZRw2PMgs7VMYE+TNSQunfyv0PDRKwGSkfaXO8UIUWfvwYe2HQbJBeWd2fxamcic
MWTI0omZCeNvM3x3G2jIN4Gn5mCRLWy2OvenLgQ8HWKXYvqQkcXol11uatMr7k6u
mTopGckp2xDvq6aM5tzivYYXzTUi9GSY+TJX/KfI3ELIqjLQupGDDhK8RltWrlqf
/6jxaRcV1Lm9upU7jkMdGdUlP055ydWxS0aQCods3Zv6TsnQvOAYJq1Z1uaa4OK1
9xUhb/Dk0EHPbrkYPmJtB88qFb+snKMiqWurQSlQ4ZlWrciovGqc97rxluNfvziD
yrSWdlUDXdceSzR9hfgUFBLYiQX/E5xwEAtl4B3fPu084WyZOl7k70Rj2SvEtpzu
iube7vWo99D7RVWuzb5V+tvI3yMjqfbO73kvv7wH6yvEqhmW+nOImffJLjZw0CVJ
dGJ5rLxIcPtOVVMJqe+nzZyckmgIWvzozvr3ZSdBuZSADsRZxKybQ/l5pOxl1QJ0
mizTILs9GJYRI+U64cs/hnkDqtRy/T/UDiGcnfqlj0pXNwCUYGmbmAM8dMCROhn4
ZjnQ/ZMkGs/baX83M5GNYptrSxEH4FqXGlHZvzNBKgSTeR5VcqlYubZ0t7/JGQzu
ZLdziO1SB11A1yBYw74pqI+erH/SS3Z+lq3ioKIdf5ka4I79WtdK2E8uXkTyQf5i
a0E2IS83Vo9bVJdhJ0LWQ6MV3cBvmLNey+OtcztqIyzJPdBlGmhvWXHnX2KRq2Xd
sgS7Swo/iNaRgZtIEuepzuOSacwtzRnrWmN22BB0aTyQnPYgQXb45zX63VBbFNlz
xAJyvzDFEslenu3jRMqRN++qGJkg/0drLvNXqad/dPmjIkMtM+9woF4KUSuMStiI
ClR8FqTOPUjSMxcFpQEkpG5RrItp47dRg0pydjSnXvRi8TI/ZLt4LmCIHLffRWYP
BY0v4gdIIbE0dO6DC9pzG3ERugjuY1jBpYJLwFm4l3XSe6vUZfjtskNmEMzZbiA2
eikch2+WaTGuJMo10WHuZod63828BPzDb2yNN8Mx+LcBr/Fxnh4GGOtBy8loEz+E
CzCSPr9u2r7kF5Q32FOh8/ny8Cov2Ffti9j7L0YC2aN2dQb2+WgEyL+VvuzXyuND
6XrHa7QSpV0VKaE4ms3l3YXLb4FpBHHMvrqtij5qqkdXBN4oDw2P4S3YlUwkLf65
lK2b9cqJMOXjwqlcircqq4iXh767mzRG6NGyOJXQGbVVRlxaERny+iHZZwJu/aiz
G/JHpnQHiwjKlM6TgA49FP+0ZIyinW3tV3tK4be6SDoJICv8/sDbD11vjNZ5UhnS
SpEQrm6/ScWJma0deyKyleED/Csztrla2d0LxwLxTgQx7o/YSe4CIB7W5j1xn01x
R9Sgd8w7o6XQMvoG7/tRnGivR+by4XyxwQyUY08jplXi4KeRl7Bf7UV1q9ZEFcqH
4eTbcKiUNhlluqT7bwoosAEEucatk3VJbk9uk99BuXEDDSpw81wAp6/wadsWP5WD
LLioO/0gFjDapQKmPjf2ourcWFqIf+d1ynos1EK6N0u59IbwpwyejVzfXRRvETzk
OWClf1L9qy0n2xMGAjnK8mrYdcKBcBQj+X7t2rmNw9EtORcJD1vjjDjwUPXLeXi7
qG2/Wrg63VRsm1iVHbqwqK+MsUjMe3yOqf72o1dQrJWPLC+H/med29FaJTwmsfg8
7iIcvsEN2JhFS5F0bDNp9aeyrUwjkw1VEE8BmYG4tPqMJNfqoNmf6iEdmKWY/V/h
bw7CDd8o1p0ooEjanJR2Ex5GppLxNMkuugDcXIrldiQEKNndlupU5oWp/sB26ScQ
ESGzhZno5StuOKNeu2QFCBglAviLxFx62RSJLzBbUtgNAMiNdpnBGH2ODUSDLzJK
P5YNOY43ESWOTRXLD9dJThg8lSdxIWbpAkPirMZMA8GsDagd+9Xr57gTiHq4fAGz
30EC26WyM15OXhgcbzwQ5ix3t8wB5Db6epUinkz/xtBBJwvZanyu6e7uRsnc37pe
5y5sPj+ldOeorvBV2YgzM963Y6IYvNZj/mUMMCd3bEwYYn8oIyOgk0AX9nEkWgqE
skKou6SzfK+yEUxa7zccD5VODw0z6llWDI4b1gnAFN5iEpc7YAh0ETDA1XhlpDL+
rU3LgOSXcZANdlejl7Xfwlx4tsA8O6/JKIPp2MQXJBd6bxz7J6N4VfQ+F7Rn6JMu
yKNhhDYb3dr+EtciEutDOfTs9nDBZrSAHkO3871pFfDDAAm/PHHtAdUHn672upzD
DZeNf6XRcSuIhOLYaBgetPSEgqHaNCNw9gxRhP23M8GmpeoHtnM4KF4d+dZDOXMa
PhUy05k+LxjaciTJwPqWEUYwGtOjssTZc3D36E+2i1hTdhExZLNxTLgBJb0l+EgY
ovOjQMVt4tirCI5Ts3y/heQD8xqO1Mj22HNUdlwbhRWXlHEdqIUmBObvEEDUeurq
gdY4acE8JKP6l8xKJfQPJyqliTAJSk4OBjLwI6kvyQTxC8I8p0xqzUzz6cfOP+qx
hOxJbpw/vY9uP5JAe1SeJZ0SI9TYMRgzVFSoXLPzMevnJWL0lmbcAW5ShcgmEYat
eqitEv7p+1LPmcMAqwo+YvlL/II/YJ6X/k78RxWbRYP8EOI/Jk3qjWebiTSHx29I
/cGR+BTlGFi9QRwBWKBbwjBUA9kFDaruJC68gUTc9h+oVVDhSLRc7+i07Brlfx1g
cAf/6jEBuOIxCm6KlbQH6W3/0wVBWSZTHZxmliivmLx/2qZVcGCLfNgNNLXl8Sm1
N3Na5GDOuMHpvErNtP9XmDydyplZsFbrsE3DJCBjXkslE2otaUPI7BNxlr37BRQ/
RjVmvgF5OtlPiMxdCCAppB4HNBOG0bGy2+FXuN4/qFx+vELIKPp3RV85YcSn6eLE
rPV+C2ou7cAzZk5/m9DuieYBJ+Rf1tPWt8zGlcekkLt4PfLK5iH7B4X9xy0sWzrq
V55PP153v7YC4/aZr0IKuZXkYtVmB2sfS6PrkRrAYtykF6OWfkjo8YtI6f+YmfQL
GsbieUsy09rBxc804kP7G+Ad6FcSs29vve+QHJnjCQum+vd+Fhc3b/3X/H1Bu+4u
GxZXEjmKw/F5V9kAncvKY0AjHXhZBPU7nfiSDo34MCFOm97z/rzXpCtzGwtQ7ecJ
73vZ4Zf6G6WGGtI1DDXLwQdFpBQw8GIHOG1D1zh1edpFkhz3yyBLxvDtrywRk29u
4LfA6mBlPcI6ApEbFeaT3z2YTASs9f4qw56Eg2Vm/D4xwQPzEnLdCaMmbz0ehkXt
cp2LbJbPnp8+GqRgbiQrJyjn+2ZnPwqZO5xZby20xP88tjLDPLfu+oMM5CzDNttn
u6qlnokAk3B3ev7Mk74/fLXJYzgc45hJpKflzczEIKpLnzDoY4ndgKRSfKhmdMaQ
t13tqFQEka7oG4mwyHsezZAAYQOwo61Ni3fnpIeqoTSn8Yi87aPOmq97aNENYEDm
yvfaWVOWfUp6H5d0b5kfL1LhieTQDaFwTBbYUtRLT6EkfufrgG4OVm6PEbsfThJ2
30zJxOO4hzp3uZofu1S/TlpH20vCcPvplkyPv8/AX4gNV2+7czu5q91V7ooj0Npn
xMSsbNXL8qoLlh7Xck46yRVRHsv/mrzgGLUTHVre70/seMv9Xjv1rf8NVLlI7wub
uLNTAzN1VXzUe6GSWcyzqB4qZPkZPLNvR7mjD9Lwq8V6aGNKRflmb0MgVRdjE7bB
MMDK31koG0sHFm3iPClmi3jejjZSiiLptDMjHxYEU9EfOmc9qc708e+igJ1fIIDI
REXt5q0rs0hPTfHvAjcvoU9xq5LWd0DtOKTXdaFBr3+DjZXH40POd/9BoIEfUDkD
vIK5X3zP7geS6ocW52zAeyNcWQDKGlW5H0HAKIH2zxs96WWJYlT39hffwx8wZD1B
MR95m3xxgyuSXbXJQJAjtrCit7JLWeoE2UEDFUe7dDMf5CGnyNXMTfskqzo4m5A1
IICW4AS0ZvAAwFunDdZIw6Nk7mYFw1CXVcP9M/zd1GbFbyqzqRfuD6ckDx/PJf9l
6OXqjiVl1b25CsGtpXV/+KQvdOMGhFQKKCd+2spspHiEcdlNWr7Csq5GMx9UlmCN
Zoz0/53RotuKTWtM14OIqKwCnrndghRMo6Ht0gIGT+oUe1PLP0hMEN7ZYPtpzVri
yI6e0Q67yNAuo7iZbQv88Kg9wXV6jWKK6TNOuuClAcHGz9hMp50aO7g6cZv02AWZ
1xzT/x6l+uxNiK2Gc460u92fzgJHEY6RU63uRpe4FKBNwtW81eMQyuI3ffsgVNfe
vjwbj6NDbcHcZmeRAHvTuDEMGN9WsBzhytSV20rkU2lpoGnKLrzy/WaFp9W26Bve
NG9smSkaSy/cU9Ha2YXB91ZYWWttKO0OGY5ykVJo5Sgni88yZRkpj5wP4awz6DUS
Ke0SVSS5lkeBPXrDXYycF88GjIOSo6llQ5j91kCNBA0LF8nuD7ciFLQOR8vZUtjX
jZlI9H2CAHtqO4AuYDH+JTC1oX8hzOxYV+kRdelMDRFD1MXwD+xUtWJayGrMpGue
CfGqHN3k8XEVBU7eWwcHjJUfi4V8ZOrhAEi/1oaScKQH4DLg5LuNruEHMoIIwoUv
gENY0ayp0MWOPuy/QFGhXfbOF08xhQkKW8idjVNY3ngZP1hc8xMYO+9VUdP9pwyr
FNma84i6B0jMAg/jfBNArO4uNy7E7m8ESL7wv7GwAP/sGkJFECN+5oLwd4LQdb1M
9zfdjsQ8rrgN3b373kU8DlUNfi6untMfYngWI70j/rCH1YJ8tNS0IzB6c9/NPWVX
WtZVQ0H8mMvqGU+PNpp1Ph1fQKcYJErfqU8B//tDGtCk9H+o7Lp1eAkoob1GHdmJ
e6EA89Y4AD2kMgtdzM6+xIZu8o6Nrl7mWHYwJcN9DdTl7npAFKcKjOmH9YVNFrlL
VunV5YM9U0wsD2Nx1w2HwyX7xZAR9dVHuePH1ekxfdcDq7m06vXe+JN/poPB1t+F
flbILgVhfhQE72YKpnmAmYKACqihkOcu9xe1JSH8bpMt83HCHnJrEfhanSkW/2vJ
9GzqCDsMdIMGAY+3dDkCNCTJ79LSxUaTU3o8KYeGVmWnRBMb8BHmWSmA0LQ1x8Ds
Gk5aLagvNtgnj3jTyFLJj9+hrS7R30Nn/0yRNY1PuoTPvnMSLGDDNmXlNZkcVFzf
+8e4r6pg+1czYPWNm4LB6L1UMcVFA/MOU2jq1z35weiVE6sFFNxm3R0Hk8AhNHXK
MvLeWOHrNu/+Nd6i/Yf4EPUVn8gWgpJ3l2hIrWevSCxTrut5SJIr6VKDuOQgXUe8
uuAEhm7uV2V9JGu7x1iwixZDvbet+Jr6fFseK1q8G/UFFijiZ7S5EJpn0Z50/n3I
DfGb9i/AbvDe/CKh6t/Qly/vi14T+tUJI0qbgikS/RxZQr7yZXnHwQAFZAUoeaIj
3+yhkwifdtPrluXy7ARojHMdSasFwBeQS6OS+4Wqp7/2lR53eoDrbSqzbm6VKwws
Gf1nDKmrmgAXtzIgCMknqSWfjZuoxjcutr1RIdEP91f8JT+e6zL7kDYZxwcRGKkk
JmRgo8vn4hvLfTo8BGb++VbyAVRvsn9cr9PSaCditFfNqdk9rMY4bsnJ2jOovDsx
8DdI6Sf7mvFvEb520CkBDBGf8SA1tJw84xSImWpXwF5y/iLSvtvkLScgwb/mrwo7
8xCxVNRmJJtu99HOg94d12KgxiGFLq6reKNheYlvLreE0AlL5pLdfIaQItRE8ORA
WQJwGuQup4q2+efKSHhLS83M4Vqa6G57Hf0KneFAx4+yrL31vnYe7EYrxasnu11G
UrpzqxMiIlSr9Pa2Tpnrs1wVTqzN+3apVwePKpUjx/jfHqPJ1WPg8MgMldUh9lYT
t3ubOMoSyAHxaJ0ASYVfQbJTH6bQIM78ksU6QgkWs1aIjgsrZAdLrD50x93JqANH
Vs5ku8aTfgK9sXxMjGld+MDgO6NjGNB3dQ9RUv/tOaZV/77+WbEFDZPzVdwwNagu
NulLDg1X7K3LxzLfrCdu7xR2lrKAAxc75Ip8+RGJVo4g1VS/Soj6fMSWHBv9e/QT
5rVnoapHHGoI3BIpOQustJ3KsZVpspuzHp7I23Ix8juoBqLY9FttUEcH0pwuVGkj
xkURoNmoyRxHdiP7DECUJKygZSCS9yw7Y0ibAt1VXm6AB3Brscn9FGzC/B1vAxEL
j5WH9dJHUseJuORTVSDtd3IOuJ0bMMeyFhVj1g1SdUa+ZN7znNMXSpfeuATOrnxG
7f0/g9htEEkHoCY6uLFEx2Wnktpcp25hMMThgfSdpmrrszTC+P08vC3gDnTt2oow
XsHs3bnsuiNq11JyTAVr50T93qZ9q6lQAGl9ukJ6SXg86eKprllHP0WNQ4UWUVBD
zEjtsAckBCF1PrR0cnXgAra3bBv/rIiigaAXRRHCzg+IqhKBpv93b7a/rKUQj/xj
tDqfhncFttd6h+RXwuWGn3tqBClzLc0wRuWsFntKXmkL1w0dzfXJi0S+hy5EJ08B
6swMcGD1nDNtmVyJqAI1Ki+zATHeDAcN2oj/1HypddjqzYpuGrtmPYXaflwIeB6Q
Q1OiuP0i2vIbwIJyMA00wXQJn8eIitNZq2/wsFmM6xdqoNX0uiaX/QhfEgxi1ym9
sX/VRr9froaEHGrhnv5icPQKPJUfz84MiiSAhd2yjPEtar7qUVnVcK9aEx7YY/nw
Q7VKt2qgYpR6hNgifHucPqoj0mE+HAYhapnl2kXKQcKZqvmaMNmZ+1XOH69T/kUL
wAEyzJ3HvVqvDr0EaJ1JRPlJjmF8gJoE89IVC2phPxGlX7P38wcXD/Pun4fJZeJC
rUGKffYYroHkhnZCERX0rci4HHDbGBmjVn+E/8OHB18ZK3p3MFm0QvQnxlN7IzUo
FHgD5PC2ivNUwZbbOt1lh6CoVkTb9FuuDZ3K0+HLJeMXVO64pgF3pd1YbWmvLJGC
fk35APhBBk467RIP2Hka4j23Hk/8biikqFT/KaBzws+nBE8T9PVZmZ9FWQoAvftp
M7XDmnxUApxSQHaR0rSC9WoT4sFhgGqRwkuZdEdt7z4e3bO8vpTQIqTy8p4sEIM/
RCk1t1lGWB4Q/yh0S6+/t1Ev4vM7ooQZUytYiwDhNvuhlVD8iSCPq4TIJMlspEFc
OaXQ5k6MvTUxN9P0TVzRS0RNgkEu6+sqNX05hWMHwKtP+5sv4W7SZGPwl81wTtVa
4K32AmO6DR/GRq74Q0gG/ja7V3F26byMRl/ZF+YVrimz0AU6Bj2g9bObqwFrfIu0
VT86z/xopxpBY+UpbM5l/Zd8PtMRM5xZZ60hTFQDNxe4Zf6jiW1LlogplLUbkrQD
kUrOZEOzWj6wq6J5oe4m2TfsOt0WG3G6YcX+vp6WAx2YvxXTMwNQ3dJh4qpuvpLY
e6Nk2LIcCFQnQMDhGc34bpQorAUHV8v8eDrBgDPvlR9ai9YRjc/zXMZVwjPr3RNG
YXNZ4D7yyILipuzxHrZB9Jx3XlEzSkTEVu5eazVA5YmeO8zkAw/aTOlCHDGfB9Vy
GaLoCRgN5D/xCCEJz1EKY+mvqgxflJ+NbTzYMa9tUhcUi1k/QmEZOTtTBY8bQN7Y
8fv+KubtGI0J5No9Ud1P+llmYWLf2prIffYOfmp24wG9G1J7SN3RwMYxk4f+0bE4
o7JX06z6VvgrdB3AMO8YhORieAtQrFSINTPGK1rV2Jdcy9dProLJwNY9hVb7ahbo
r/1ibliZ5b/BpTU+1VYXWJNPJrx60uV/g9sX0QJkFjuPfViHdPZs/GnHs86FUXHo
DtYaWLTKdjHeJJ9cLqly1xMv41HhKns4+6eOltsyQthOhDrMVYVOikzP1vIBDhm2
mSJc3hExLiH5qvZKCx61FV5qA3jpvu6JteVd9XcehtYH9dPwKTVzGqIOeB0VBBYo
LzBY5sf6Gq/OBkudXTIYI8y1xHFKcPzpEW3t3C1Zkb31RAFD3FcsmTiWhh3PuV8D
z4Ymo2Y+UYA5aQXRzmI2LlLl+2hrh3Gsff++KpX/RM9BREi7dGIIz6JGRtv3npXd
hYHX8L+k4BeLngVtCpGXxy9JhxjiRVebDsjOAAajYQyObfegYzLEX9zk94pCfgiY
6pAinNBUMr5xwCWufNYy3jLdyrqVaG2j+kXHULOcgAh4In/MDqM+GDZP8yXmq/d9
0E3JX500j8lxbpHezr32+3FOSCwdFxXLA0E4Nfgyb8SHory6eeb8b0qjliFlRQj5
nae94sYdGxpjp1K2dMCD0+4WKuImX1M4HlTSvNLpwfywBPJ7PccDr2qFHkj9XvM/
bYnpMcukzqHLMvWgt3z+ToHXogs0F2cE26xcNZOrQT3Y8/lt4aVXO1Zx1PtuSppw
oQ9oglcFdc7cJ/YcRB7A3C1eIUhvxQhRUy9Aiu0ORyqOLplfdS0k/oM9xMCSsIXQ
zv/z8TLy9iGqXwxrTMlYMKLnnok/W7/lhp5RDoAf6QcYbKc9W2vXvtmB8do83o5c
Qkw//oZppGDE7D6SjreR/sTIgBNc/1b0Ev4JgHrRpAEhzCVRq83I/bp+c82bIj2h
uQjj2eoW5fc8pSBgjDuj1tbXOIx8j1CprjN+4u7kV8COB3TBbigRJ+15R5MUK10B
k7YY4zY4qbiPwo8Rzu0OvTi5Y21Xun3TGgMlHY3AnuLR6Ttdg3kLNpkkgXo602Ar
RunE05KV4Us+MlxAN3vy8vct8eT8jvpkG1WbuGmE7B+mjXW3ZZ+cPx9uFKBWv5gj
BcEM0nkCN3BpB2UABWi7vx0o42dABY7OeHoac9pfj5j0Wtdtyhw8Y/KwtDrVt8A3
GhimcUSSjcQtBVKkdEiiJZf3pNvdaT0uptcVshOeiDtA3bxxyZpSo/kb2lvtUFUX
9jcvrB/8CwobTxxIsF3qiNJfI8HH8R6C56OLYxLtwcKy4TvWdBXuvCxzYpSeCEI7
3RyM19ZuSbO8R8jjWOz3iGmOf36EyXMLRkecEeqKoY+JaSuX/ptioNY0FuDnJ3ty
g1jWQ1CcH6V4Dp+6rkYYSymC4DOrvsik1sr8Z0fmooNOCa43yDk4nasr/+pMgNHo
51NDtk0ve8p2MAhDkPPjFWjyGjrJFsVTtDil0ietRIvsjnMSBWTRdMV1K2WITCkV
icBZ27diXdgGCTws1sM4pz0KSCSAYhZtijjXfqqUavRJcY5lE/C3eJo0SVgaOPFP
FazDu06SN4Q8uc/qMw2JSjitVFCJSYITADQTPqp7YXniOFjtDeAZjWUWvHOn1f2d
rUrm31c/UpwR5daOV9dm6q4+Gsd2P2aQKNPUfH5uphzuAzBaHQtFEywDnKWLj5XZ
xtLHSOXM+Z1mb8KRAzGoD67wWmU0AFOyLQaMTEWS3S+xboJjTX8XXwA8na6aRbEn
zOGOVhZ1c+UO9AWJq9ZDhTd32TNAY+wegtnpd+nir2UYyebHw1BIJxhRktGN5ZZR
wHmrqVe3lfvMZhR1o6q93sBEvIF1BdPnqPyo6/gzVZGLf638vQ1tyzzjAshilUqb
mbZ7IdzODz7UBmYxpPpPndOGeS4NA3fwBrXEFKQ8Niq77PH1gQ+DzY6gSeQYNBVM
Hz4JFIbEAt/hTG4uI0PzvF0J5wPeORDlF02vj/bxg2zb2NUoGmFc9ezdUpQZuYn8
xnhoiLeUX5Ni3A7/HvBB63zD3w78aX4qAUK2ZO9sw/JicxX8rQenNA71WAHrCwBN
rkmsFTg0TCy/3LtVzBj7UF0bbaNcHGEjnwSQSCKGBo3UHz5y6ORlZNduLtpuiY2k
Lt487/mn9p9JjENgeXrMghNaTRRqmCf8zirRBu3mOSFi5iuihAETQYvGVIoRKtBw
F9AKY3S6HGN1/wdj9kKxYv4v6ZP0T7ezLWlNYGsRSvmKDP5AMILy10GmgIA/tnvp
cAK4GckTM0mZcvVQYskpawDKtXdNfK7EK9qv43eqe1mE10mf2jPRPsXy0elqZxBT
XxD2Wh+jqx5tB6GmgMFmp/bUWX/+Dwf+MngX8kE1p86o4mDwUn5nM85AY8kkh1AC
KEzl94Kt67BVEtSfxzRGG0yzklBpSzYnoqeDgh4vJfXo+R1vpI1q9QCu/Erx1pi5
D3J8NVCkQg+MxfmDHlG5r6PR4m9+2rfPu0kQ2v0/LNDNJzpLcjk1lB+XA62mnnsj
QMSv8Hw5fVUX+4G/jAt0YI+Ru9dPS/9DixwT6JGg9Lhe+pg2f60h/3yipdY738E5
1Ug5j7x5B80byDiN10Y+vYAk6OV1DA0LEh0OMuxBjIaZdX0mhw/q3jEacahEc5Vp
7UNb67wMGesc22BcQQ0CafcjmsxAgaIure29Oa2eyc0AQrKzPUoV5aVlE1+u9GVh
KG7fHt8squknyEIOtZWoY6803jEtqWxsCOhOfigV/KA2lnjhGe+ACUUZZS3/k/gS
rN3ynUd/u8+lUKp4A5J8+O0PP3+DKgQRbcKgJAgJ90IDRFDd3sR3glf9hRy88DjB
k3h3DqxU+kKH1yV4iRiaeWhHmR2hEqO/Qu53NE2pcacVnPURuu6xl5LO2iUfEFKL
B6jasycaVASvaQTcDNEpd21pTD1lgiIiW53oJyR/w6w7/nyzNx6NLPNy6uCeaqIy
nVql6j+tdy80hvIPgpuyIsOvp/GpuMc1EDniFN7BCvJbKZUbyEwIxNzLUOmhVrCZ
RWyj+OprbrGsF60Fm3zik0IP/96x2ylIX6H91S0ZFWA+j/IWRn2apVFSCsotZQjf
EpYzIvSYY2nXwW1/IzFMF/qFt9vwFgIEB6TwJ5k59umTrGw2a2uANHmyFJsC24sQ
mRd/McnXqDyXlT7u/KHW2zl0wCH4+HsIzuRauN0LFsPfUMA0OCdKWkgrQccf87g6
9lN0RPb/oNs32q3oXDZOVkJXiKZJ/PKefi19qsGjsXDIOj5BsbWVISfm2vxsdzXb
mvXnPFGEutvtP9OE+i6Bn3uEU/d9AK1rHs076PwyLVDPxwe4hEXXemOADgMf9GcQ
mdIxTpO+hrOtPAhbWj5l6pRETTToGco7trWqSUt9RhBxKxCoGHNsv8sEZ2jMk20H
DKdWHX1VcPV1gIG91e+UrxqA7i0pTi8MCY+jXqfaIaeAJnPhb5edFbEkD1gTl83J
LlSqnVKgO71VTHgndBpAKRFgApFOGiP3/+e7jVdQqM74J66siYgze9QoAJXLhCGj
xiTBwpb/WXOgCcaoXp9ZrHQcemD9LGVsypvp+TKMg60ZlcA/AWSdKf1O/9n5jHBR
Hte8GCtJOySrrYiYDEfDfXDvqwBGLh21HphqV62C0luMNtr55SyUjZuEYTQjP01J
WAZMbqfHf6OvzLq3ut3bKMCq1nGqsSldFw++x7Pq660hymh56MsYHVwN7WwJfTlX
8nOoWPChTNXgFmPaBEL8yYCPP6Z3thwzu6kJ1um52ubU7DqwFL/z+M/LZFdup/Gx
wnTR2nlxQs2THk7I+EC9+U07t1iQ+AZ0pzYtTiCPjALWzsi4Z7PKDcmsDTaMVA+Q
8Ik/sjHGlacbXK8A9NyjeWL+70FlnuSbgwtjMMfdCgizrcDzwGNk/fTzZ4MdzUUF
u/5znft/KhfK0eKMay4gs5s52Us6xw7GimAkSFmOg9YE64RoVE0c4USXlmSBQA+L
8Uxf1MypUZw5Jazw+hJ1tKv5SSbmVXuQX4HAsJVxSIuygrmTFcdkQefVZNH2I2/J
YxVTC8etqZ19KT0H5lw/lM8LmKdvqpU14zeRxgPkGhjsYQcPpDOUg7IwjQcGVQpN
3eQlb2FBs5oAKR9P2bjp/tUNALE/V0EoEIemNjAgexPZieF8tKylxPtpPgPPNpLi
/xmM0LoYGJdprub9CF7+eOWYeTpQtFrc/nlXR7zpoS5XhMnL3aD7z3P0SASOn07W
AlJ4GP5WIcgsqVzMzPSObj8lrKLljXSy+BjsxxQn1Ttyh3839q7XbCVgdVF5+EEH
X6jUQBugtd+LqXlSoinGn8wMYLkHXqPImrcxqJ8Q5sv4GxY1HxWXOjPDLO7b1GBa
tJiM7k3ibycLsrj0ghPCEI94I6EvIkjAu6DbHVxxp0EKJsDUpBYSFbKKjpAMQt9u
wZXZj3JDyRvt4KgWAJi7+2tu9tfMr4Cc8n5nMzDNvhr4VUoODxPIjQpNanRZLyXM
Hco3ihgREbCm5c2wVCqC4qpHCWztH153idgT4qbJbqmYChi2/KjzhUVAyoA3KAOv
FrpyB10LDU+Cq0WMjrcxKC6j601sHLgfUgdu13EO2+fLgXFrLGS2gtZiYF+Hv2y2
ulyIyYKUgOMGpL/1G21mx15ZuOfweOuEV5esD3i+RYWh5RZDjX7Z9ELlUd9FLOEx
dFQd+J+yiZm3DUrprbRy8xOHwJnRJysCl5DaotFquiuBEe21/mX31AZz5IAtala0
rDxsKdmKX2//q9E/CS3mCzVn6UQsvCgUsCuTRZp0gK9iAbw/kTk3DvLDivCXm6na
PFKstoNkJlBjfUuDGx3EacDuZW8XZcCUPjppdK+xQpLlMrX2MS1G3VgZYCQVQuvx
lQAyyRg/Me1poK1tBftI2u2J9dFdV75YtjR1wMgspgMZ+hHSiixHz7kdezk2FZWb
MAvXy/fgR3o+in2NVDLFoBrA/1nWorrTn2qO0x+nQaqxzNl5LG1XCk6PSD0Rbc6h
nsPj97d8boW26ZhPbfLIRMy5cY5XgqIw3lf/3t/XYGt/gFVbSVjReRbpwt43m7RV
prcG1UYUGUHjbsVBU3dOj6fCEXhh0CYI4XQ+bStdAT3yAaIPcGghMxUz7V7jT7HW
2ZC4AESBuN7suAWcj+GFezBLh2SXWsau8dZ/fHq1lhFGnsnmlfy6giKPTx3dlyy+
bSCDxClHwY9EUmNDQcCiOPIlBAektZJAkieqFCCpjm0XTAOmyixodggzHOMBxMhc
9XDj87OujTpHOSyA8p4Fah4kULQ9UHq0UAhbykSnGLdtJOrAYHBdc3wX1LUC69AL
C6YY6Ea3AW3PkNoI53ZtjopaqP85Ozgf/e4CagReJU0ABzH6dCB46QsktnUxgLV7
wxlv+xR3p2rRrfUkbUpLShvyCeu/uM3DfivL/4egcxO1WRwOrChIXqk6yO7MFnbD
nb5BE3jCiFy6jGyH/XDPmQa5/KjMCXJKF7wIjaAxB2rDBzzumx9gZSE24Th+EBZa
pUWNS7e3mt/tcgBaihkluXniyQE8OhXWTfVJwU5PkZtoSFkt6N1KNzwf2X4j6GdD
uwnxzp7okGVslLQL4IMMMO/bj/XR/RYvDmyMy2ObcYc8mbJsJlEr3PBJVwm5SK+i
elKuays8yCzCd0jw0Y/FQEENwj1PAS+qfr1jBAfn6e8DrBKTQM6mRL10+bTEVgsi
pXMopXHxHdM6gkyft759OMdfiyoDSs3m2uYNGjTTSsAmjsKo+qU9L1vJfsEARNWC
HkfZrvX+JOA4x0p2yDjtChaKcjLH9SnvpyNhYOlVSJNONQxenRfR4HMfWandioO3
8VQH/4QIPN3r+TlFJAVy8xioFHer5/sAnnBaJT1fkkQ4GHHYa68NigWbIyob2Yi3
TRQsW8GAI5gmXZbJhFbQwiDApL6KmfcQcPT+5eOMh9cq1hb+p5nOQM8gXZckl1kU
wG/FcIExTq03EuMWZCFnfkFNQWTU7tbF/WD7izg4Laa26q1BnCRlESAlavhWvyFu
CUhOYgrvoaAR9LeAZB/qAAgbi028nkZto1J7s2iLq3w1RMEFBcRhZWu37zHVkFVB
7XrLxYQimpT4+Pee565ySV3IBG5HE0YxNtLfAak6LLWomUvvRqQ8/t0XeeiiA8ds
QLcTd6EgTnK+XAqu1MIZNrh4EhtQOW2WXe3Z5l54PadMzTAEqP2wwprBy3XzZWqt
iGmc1TqjTCDwxDv9q8HGxp1Hq/bV4BiUdsy6SEi/EIuZfINrtFpjKaOiMlqpwCs6
cFwqdxMz5HJ5ufkNzmpVK9uiRFwEg6GqZR2GnZycIq45WVPZ/ng3pula3zneXonz
hzD+AbyHS5DEgm1C/HH5SgzpEXP8JBfdBmlmoettStURhsdjd9SmutaBcauZJJPr
5XW3wZbbnwg7bOrjvmyZtyZeGha2tsX3rTwn5+BKAOKTNnikE00Tv04Mb4xFJ5hM
CttoFd8I23O99GclT+1Mf82gOy7LGadYAsJyVPFGFQbxAKeSt12t2JCi51XBVm7E
z5hxk7+pPv1oCJcI5qJQZAzB1rBTEdCocKWJ22lZr3TexYpXRaJe/M073lCn8d3f
204CF+55EIWxodFsUR7MRGPbHd41c3K02U2f45U5zK826DCZylZOwk89qYkhHfqx
ZT6QAAyW9Fzm7aBfrsiFnW2ycOiy1DUWS0Pa62X7TyaSS5EQLQo7RjuMVoeWkLLm
QCWWKm8z/ZgMfEZhK3xCHwEJmiT9AWxAR5XDhrZZZGjcn6pCKOEGesUh0u6j5PKW
CV/XTIka2IbWhy0yMG8sRQglZFnSkwIhyh5Hh4PdMX7AOJ6kr7gNKi9kVCYyIt9h
boEoxKf8AdOId6etsVinK2QHJEHzDI2tJf3JYpaxlIefptEk/vW4a9KB7Gte8GYI
zq2Hs4MtTWwF8DxpWIrKylqkokgtnZ9Ht8TE8y4eT+zj7yfsyT8XAYjtN+AKzJEH
xQTCrNsNzESKE8YHPeQntwkHYssUgLYKbfmL7RfPfy+z6nmSDjvwjjAtxgyl5rJh
9z9ZL/O6cpMIHmGGbuf250J40xS0ud/EGUd8cJAX80QXtIP8A/SsrUeT064hcDLK
NZwrqIQ8bYXdEi3MqTB7Owg1E4l285QCk8OfxXtCEZ4I9A2TMOS1Mpet3VBGXQve
M8Ov/guVaqTWskGEF4IeXjr6pJXSy4cYIdYQf1ap9/CG9IdVncxmVrKPn2ELbqPB
ysNRSOjV8N/MGUz8XTXcFWl+37mlAY23Ln2eVVSP7qR/G4+hU7J/ZwO8fA4vlWXN
Y7oqD3WqTjl/MAgZAhXGOkUZ9mWh75HnrhyvOa5+X666/zQHsw5tUe1sZNZqEQ9f
SraPXDFO03crCAJ70DP8MvDn3V6X2Ls/a1s2Lf7cjtEjTrvoC4qu6tNKGAb5ixF5
eNRkCzmC3o6DlBMQn2zqLO8bAGUA8230BhaF1Eg+5hA+io/wHndYp8LzGiJ1Fdy2
MHBxS5Xy2E0qPlaaKfUb+XOB2kkldQAiK0z1CYnBX91FuLzl5lYFpq5ONUJmY9zo
YlLkvCThKT0go/Uj3um/lmyS+Fo7VbfF05Reqmqh7N2x/FmrhhN1ng7G6fDqyGaC
TriauyNaeHJjuPZE/Xa1pMv/pY8OHcUsq0ydDfk0Ta5fHqj+bXXqs7iM8uCfHK7r
MMijtskBGm7TlXt3Q9rQidgiIzjduDTunzYR5YCNTSP3UftFv/NwwxdAsHfWXIWF
w62ixRMVlLz3yEtPsBAEOYyhhSlHL67w5FG4ndjqNcR8APIyElmbzo5PINbhfZ8D
jKl7EFf50hqKMoEF5GzHGhnTXzx1r3cFcCXm57UkqBS78G4Hunj/Jv0Gps2sK+vH
Aoyzk4O/mVS6+OvjEgvPoxho7TzmQRD9G2z0LKol93Iox35vXYqJkrXiUMCUfYly
Cx28nxJ/S9sQHndGHIRNfjSIQN2KOxwadMQxfk1iWVFXu5Co8cl+VnKi9QUc3+vv
+XbzHZ2cqd03r9H700jIDvW4/kdrvNy+93KpBkvf5HyjFDOkw9Ld1lSDSdqsQfLd
nY7NIZsemy5ipZ/HadFNS/DJR2U1YHmB//RB2GAI4nhIRaYPHY7NwXSaY4tw97bm
VK64Bwpxgb5lqDEcjE89b6k/8ar749aF80Ntd8M+lN3dSXkauU5hVwZwN7zhj2e2
+RfwxQFhVJUw5iiSdgMEaIcFfVYxUuGTtDzSJTI7+SRKiukiN2XPKUbVJ9+i6w9B
iC0NV8iSXz4sMqHF1ke84TDVR84lBQe4fiGEroPkr4FsSQy9m26U7i0usUB7hCts
/bn1RXPQFYPDGMBnecoGqdwHCmc2UVN/WBOJ/X6N7fsthBahKf78mpm+sgGbAUZh
WFgQXLQc1x6aQmfP14Q5U++K82YLKvcxG+BNiZOAmU2XojhHmtk5YRDjBxqkfVDc
IhgGFTT8vKabE6GppYIqdnyqwIZvmBQ/oVcIMvvkkGc8AhVMvcxQwKGln8B1pEGd
f8ST0eN//tymcNl91tGqWHEdGHj9zvuIQRzAOMd1GHsCdrrSl2gcargx+/YjJKl+
N8R0Ew9j2OPKyOpKWUbJcXwKCcJjdBylOAgqwdfB9morjMY2Y5cXejgm4bGMrF0i
PdgcF0DZ1fgsIgaRnBA33MvmffA7cmiKu3DadJOJvLVBl4eng+dRO3WBJBgXbY/i
dk5sB2VrFmD2dNAjhbG9Rc6qu/l1QjEV6pAY1COgh4OkhK/sdhgAiXRl2yrBlnbL
TCn0Ye6E/wzwAXgOZdxBRjdI/50I+CEjeGJS61swrvuN9eNVO+9zLCpL/m7vE9wv
pOP0TGm2tXAQuKkrHjoYXXpqYGkgFjN0plc02v0DH03XoSyITqWI1d9DKKelftTx
KMvtsg1QVWAP2K6ToKN9g4SadS5qUeQF1OpF1Eb8sn5YcRb9XKfcEiQW66VZsn6t
R8hU75qXjabkGfMV7E6M7hiSvFRcOBSAKdcgp5+tIpuj2KpSmb9AxXa2zFEDKVPA
WxSsASLEsLVXdyvRwXPDcizXMxCfYOyTgYjn133z81DKtHz9LrxNJnykgPkZUa2+
k/DYVH/fPfc+ucToBDnoAk4PUTf5+BQyBWfHpm2/xhM7AtPqGDUbeiOD5MvDfKZS
AxyCMpCvPzx8ehKoRV86PdSmr2A7/isjvAt830+hs2q2+n9aAdf24NExdejgycNM
Zk4QHHC+vEng7DD/X+5njgBp6F+CUq2qJojdebtX6iepiSH3F0tHCu50OvEyJi2E
dQvFQwM0nTeYPeqM6qoLCH5wTKygEAGgySSw4dEqlpJfcraIJwh15WzTc9oadscZ
e6j0sTCmc4AsPR5Yol2xWSARLICGfTuUerbdutTjsn1zrQwHA27JjfJD2PuWcydP
Qxw7u0udSB4uumi7I1ejV4n9vO4vaged8pSYmaXXU7353LkuiECNd7+efANwuD+n
0RIAr++7BXId6ZeSNCCtyvFnTgXF7KTKvdzdR1K973HFI+Gt/J1r85MEJFIu80qD
SS2hpnTQ11r7AmzaypHTazwqCyMew/wxd+OIKYJz/uBiK2P+xfoMMPUGGHWXU0a/
df4FFI9rZCoE5AMGxHSsQCQvcBrDYZWuLE9fGSeDeA9MFJ7peBYLnXzj1Rh4A7YT
duBCsulA6NdBMpBuMwakoX7Fb1u2xLY6gbe2QsehsRfMrUIIZ5qqO2mlQunEI4f/
7lKh7Q4NkhQqh+gadzS271KVJ6m+95Hpyllg9MRyByfLVQwUcGiHOm5zVLoIx2TP
cHdMO/n+I24HRGxPpfwDUOnRlYeALTPc5TIeR/Ri34mArsr2F31A363pezCr9hO7
55CdmYl1OT8P9dIfXpNFmNm+ZoUx89UJNyyYesLTlZWHNDgbHAIYdEuSSjyWmUM8
iiiAvI35zVS6FKo/CXk2L5pCcSXClyx6AnZXR1SWKJ9FYstb3UEtAi0T8ySkElEk
Gwr1uvv7KYC2puTZftcC4df7F6q8Kl+LQMmxrDhhSlqhIvoUJmujpjobsNSNgYyx
iXLX3+/Lq4zNU0KS8Phvx8uD7XHTquYPAxyLIwp+Q2XxFqQM0p5b/os6ybDge7HN
PXM+pypqmUbk2NFpCbPdrP+aDjBx2/u1Qkr7x9yj4plFleL/nBBcuzNx/7giDT88
uEgtKw1GRib8P4dS2rLi5IXLk2d55okokZUomVNDqbDQS7+L7sjrMdau6Z14o9cO
0nlPGYIeURRfYL+6cAXINIvRvWebqTTfaOy3G/icYEM8WHfzkJIQDb6kKQWcAcAV
IMVj2+3xPLbM2/al8UBrjYHmHGrZ6gWk6am6oqPfLjOB03ZfwEq/3eNMfy0MJEXs
lGB770QjadjM7uqTyJ77an64i7gkS0BhU5JYzEpLXMVdtmJONGs9Q6jgEH6Tqq1P
AE+sMtRkcvXQGKCn9LYbDr0b4QSmGgzIr9kQYYfUmRZX7ZSdbqE1WX/UzeDPgs7E
yLqh8Vlsgnog0ear+aEnpc2kaXuIMNAZqfDVPaoIovEhbkNSW2asPKbak8bF9XWW
98edlxfie1FJ3voX/RXK6hkFBMpEPNGKk/lqAu1QG6G6KT4HZQazJ2I7GnH8lxWW
nhIeuV9lx9yBRVoxHLe/e1z5/MeFNmiQEuFGFkeRT7C4vJ0gILglIkdvmPmkoW7m
LafeYH3GeIyJ8cDO0KOHHfPi4CcDetxqQs6JqQxATgtbI8bdzodUTw8ejLmfdDwP
uJ7Y9KpXuvyBVi7wfp4ESXTpf7rXLTJJANys0ayZN2G9PIeLZvf93NioUdmgGBme
QLns/CVyiihm5POzrfX80k6gZF9lAYiB9TqnRu+ZLvmPzTdnPvkxF474ljvxDe3G
NrTc4Z7oTY5Y37Lv58OU/mEobZ8fyNfrQUWJ7M/tVbxqaBtU5BwgP/uyHnL1YYQN
IRhiD9Yqfo7jee4/6RsaDbe9JezEjGKwwEuoKuXQmB9CU/l/3KMU6mFVeWhuxd8G
FnGjmWHlwasu/yTSF/VToy4FuRF7Y6Enboo52qSXi3IQ8RPUyJRNHRQCnjPKyex4
Rkl2t+xBcTDkf2IbUqU49Qc1iig1a0dCnrsz9jEyxKAh4SzjfIkWk8eLIAkOYHnB
dgQuZkmASkUPRuXZoozoz7QZsYvL7ooGZMsDtcHZmRfGdkXvd663DzjVsSUspOiP
PMz5ocEAJzJQx/2CFL5uVeh12/EK8mgK+wJlkBiN5kjAfkBGz6GL1GmHt4XzN022
q+L6TxhCG0Y39KQtHBLAAEfWG9zOBognsLnkiY5la3vxIOqmsWJ+lXycj3i+YtiK
bYrxbxNBW2XPE+GeeLdzmDu8J2zWgI6EaFtV7S3kqiTSx8cUg5Z0oTHDzcONqwy5
jOQY7xqNryZ/BbLFyLC3n3C2gLzHxrlP33fRWTmkpQhZd/hCp1kKWu+hRLP/O/9/
M1PFyT/3q0JadAFbBLffD78C81z1hCXg23TU6P+av2BQlVPi7UoLsVgsytEspPgo
+vrMRIOdk8z0ZYO8urpDYZiK13eSM58zdXrPQq1qidzdtiPK4Sg+Nu7EPfPggnkC
pk3muiNtpcdGF39CNL4J+Am1VHNxtQEHMTgwFHnD99f58eoH7UCTtjkCniqi4Tve
9dGLcqA9yV4JzZWtxyeFmdvuB84yfW2I2G+xa1szBmbA2efJun0Mye3Qidp+pnfS
sDMjY/RQUE5UupTI7MQMjla7XRvnITbe8DHAYOwHL9m5M++NnYyqjiWIpavFfjj0
lDS+C0KKaJIOHAFOhL2GeacfwQlsfwXr7zK9VxP0FR9ebOsZBSA1JBickuW4L2uw
bwh0bDbVMEch5FffMsux7zRosmnaV1K35XucBUhrUzmTLC3YFyQ6xiXlE2b0xip8
9DbUgHlmxLv9jMjMo3SqsdiuHM1j9ZIizf7f+IqELoc7OoyQqlbTeX1wltew4OwJ
3qs6nsXqS0IuFffNtwHHaU18+4akKOxxtriCDt79U+5gm4mH8zFUzo690RPzAVni
nmVlGUZGQw+qDKAsrcyJKLzqwL6iofLcfCXEn5vPfbFlJGeLxedG9dzSM5pVP4TV
GQlqOdE+MWoyWwhlkSvw9pvJ+RZ8u6ELAm5Uq3lXXiiqLmXcNpMqfeHlFiavYPHg
qOcMDSOhRNhWcQGRM9lHal2tScZfCjAv+4m6gwnNUjZAnNXq3egUYtUZeHY/tKcq
dMTBnMJEkts1Zp8lYlOhmRG3vQ5yqIXDqjlM5qq7tf4e0MnP0uZ0pDzvATjMCMb/
xl3S1acb/YxIwhrwxOC0BPbN+y3d68RP7bW/utXfYcaZMMm3oBMJLLKNgg37Ivnj
1O2uBij6gq7oh9h38cyCS4+6I/fZ/UclG4+tpJdp1FWx7iLDuuFpL5Nly5WIjsg0
WnHQOIj/83HtJGaNOujxDq90RpLduR16kKecUZCA46onhQMJYJAYpC6RGzhyU3WU
ZfwHjLdZiAvzh1ZceRmewLhMQI1SsPb288Ukh2f+UfPOzYWZFeh8RLE8fq4qM4e3
pUgsQbWM/FclGOORFannSRQEzBU/4LD2We4cxSdQm6qSTGCU0qCnU9RaNyXnOFex
/x9yosQ6OrPY8ubkykoiQxcZCedW5Tfp2iMflHZccElEj6nTfkNeTDHEB1SiggrY
+AxMyJqvn13MRIND0p7bYZER6ok429bpeqcQz322tmT6bud9mJOZhkEW4JeV0qjo
+bW1uO1rs3BQi6klcu0kIqRI6BFzW2hS6unlZa4BeRHzkXu3rWElsOCQAIihU68Z
wDKjKjhjHmAXlT68CtdjRu8tUvAPEMyDfm5Ic+N9ldA9ml9Fomtia1S5PIQq63Sv
PvyoarGKMcigkcTbAynjnxG+kcdqoTf02X0BtUuOHOtq8voM2XSo36Tr2F2rhz0M
VnqCGfo9phsDdoUAuZs6SVW5N0dNL8I5u38MZK8aT0MmI9SbJvbJzPN0pPcK1b9F
NSslaRhBNw9tLsA/6a+dRlOAVfpyldPcOSw5cgpMjkndFBMgT9YlZm0LLi4oWrQ/
Js+9RSUaDFGmVVoUzW0ZKumJl4QqFFfPgXMQ47ygmIyO1Zc2ZzWpKJQJwLHk1smC
pqUx2CcYHSlG7ySoJwrSknoZeiKOCJU8lLpHAmcYPYfi8XaNZf5IWqcPRiXpeLgf
MoLyz5ZrGU4kwfo4vXa3RJuYuTix0MyQ1Y1fLlvUHR0HCCL7C5upURurSPvEoXuf
XxqKvd8cc9ImlhUpJmtXbuW79Ts4joKdOEHnXidONF4uMZYUzUtJ2S9VYK8o2FFf
L7SogS6U5EXvKWAGd7BkwimO8yC4nfaACvXvYh8cEFbsKDOWAsTZ4SFOHCzVIHBn
6t2uXIurdpkk0wYwG0ZvKBYI5vJaJuQqtwvgkTGCJLnAQ4GVLw8ZIsjPj2dDG11V
8e+3IhmosWV+JsYUIF9Q1Np0Sgh5S9B+XpSUV6MP5Cf/vpN9mI4WgCcAkCvofuqX
SRmIPYWvVvvoXpjRjvoGXdG2ZiCx6mBzE6VR4V6V1t9YcrXngpQJCBCb6YvFORwG
tl8EUGEEfIa+HD0denQwPiVz/9Y1UrjLCEwwrNvQheYCxsf5Kzd6Kiy0Mc20EU2i
I/ezsrVqmpYBedlrZvNaBEHcRReYCOffbD5Q3x+TgDogbpRKkuLYfL2LwuIE4Va8
Erbbf6f6XxbAPpmxHMwuGJK5xSdjW5f7MgfHKBt2gf+QKAOD01khJkIaMCx9Usmf
NKHhJSdRL3MLJ0rFK2JzO4vgySfMw+dHESZY39M/4HhRpacvGFHY5nwS71qtFJrW
u8GHmLqXR0QG+AqeOj4odLf1UGsXbbK5PDSwXbfKiWNDvZ9uAJ91RGfSJuOOuGHn
iKNY9vfJQb8CSXki5nZD4h2pKBgUXjXwTXpA0xuBxatRGQQzbpM3dd//aI5bsfzO
HHyyFdA7UNP8UuM4zh3MjQ0uvDmJWGZv9oTkBo3DUl/ehfJshqrnYBWtBt+uFU48
SrYI9oWRz+g9xAnV7R8xRdDIaU0JiXHZfuUbNUnNmRrC/X0NvPbXTtXmn/J5162U
np2EDAjxAhmyihC2Pr1IEzMpwrkkoVwL53gYP38TG6uHXNknn6E6sBnSdhIm7mf5
arvt/b0R6BC0q+3MQa65z1jvErk1c+eKocbUzkabRh0of9qR/E1LhlGXFyw5Qmct
iojfghAswDP9hV+dFx7cOQKYSKDHDIDQnoF1wRz0bpPK91Hs1hAOfYMW6rFOHVqE
9yQV2QQDAiscTrxiwrkC8e5I571f/FVUJqV7WddrnR/VWkpS/RTjiQ9c4oZlI4YD
zVMlAwdmrZYYgFuQDAbfu9KoM/WGKuHXow6EUtx1eCg1aLdBLXvJUkeNwvhzggZq
S+0MKG9I/NvdK3O9lMJZ+sF8PIWUTPvbMtKzvgWXgxULvjtB5sdO4JraFF4dt1QN
Des4AYDwRb/HPIQJw5Cg/TzkP1/Zk+pbohK3mgA8C6G7fyYkieVAtWWeOJb3vHFJ
DikyxCeXdq/gRLSrlTIX8QbO2NJHXQn9bM0/YjPRkKKLg14aarvVtAhLQsMub2ky
J/JshJXG+gPMhYV80hFsFgshAU9Fi/UTX5ZPY/gzEEoNl/W8hcj+g5jvrPPTx7q9
6WLIqXED1RTwu94SwzgTwP2z3RVtAVVW2/SHCxu3qZt1e5IkAcBSEBwQh3+tAOsI
X+ykeyHX1oiI6lSeDageGU099GzGN5ZOaTdV/TCXOD2P8iLIi1SrwJnIjc7pEb21
5uSEf3w5o5BBLyTWo4ybdeFE7ji1H9CJFPFh78W6UjljXQ/4hi7LbHOjtelSnlPO
iDQ+7eqo0bJv5bJt0V9/vf7kHPmKezWDHMFAmAY28lZnQCRDRFQCWKNoKb1BlqS1
Mavbf7gUD0GY9VqXVTloGb5fUbSQWtTXtW3a+Q7giBi2s+enTOpv3JOBMaRc+VH/
hzV2ganmThX9o7F+0cKVXFic+mwRMp3z4azCXfn5tctY/ltTvn7cfJirkZoGl+yy
9DOMJO4wRoeJdlfCAMnMvsqh/s7lbT18gnCJqff/bd19/EEDTmSWLeFSY8dhzZL+
+s8BR7hJdh5F5UKLBYVD2BXrNk5fmXr2qx0BiVV67hLfT8T2CSyBCIWex8r4Ufmu
77IUBOQ7ewqulIcg0BnV2A8LuPg5Jwjy1TqwRKaQR/5I2+ga9TPyueDnQIWCXYaQ
P9rHgxEvlP/CJ0tGEsTInqk4ZSmT2DQpcrqblWhcJo2OzFVFM5+9QocUtNQPIZWI
97JwNTFmD/vq362Nthmm7+wzQ95l2dCiGGj3Bm3ARNy/Zgu9oQQsQvp/l6q0xpmw
kiXY5scUfj13mHl+mb5GMTaqEo5IntZH0Ylq9E478fosFf95YIYEoOwZJRa9kEyN
nApWgKbGGwIq1nQHz3Gp78WjN7rvgddoTBRLkoQzO1I8qpb4tiFHYRdvLJvodHC6
PS4XO4JU7qDX9kUnyH1buH4SNyxMJU2bNoUy0a+517x+tQluEmb9KlGoq4fF6yb9
tQRg2+i90OGhr+ReAx6TxqlfxiWxxj1fUmoKm2L9SreSHsB7tGPnl4iZ8xI3BwWy
A8uC0Orzkv5JMjLZTFqZiYhNOenDN3BJvtFnIqXzSv4qRB3hoaRcUPbmGrdtmtMX
1PKxTVo0sI4JdGeB1XaYuMiM7k4vENLNfVF6LY/bEhkvv8S90CPWvURWP7rsq5wT
oXJQWBljMGsbtO7uFd1xbz0AdLTjWqZtW+dypNnVKExAWsB10mpxL1Yrkh/gftoi
n9jCNqrAPtz81J5cZHBRqSwELwevaFJiT6df8CmLw0u2HBkQnn+eElZviGC09pir
bzDfeZ3iVmPEUFn75z3eNq32nD24UbTas3rbT3kNegFh2j6OzxgMCeLZ/798foFE
fcujn6XGnz9bqe1hWgF8wOZAIvlHUnZKMm8IHGaZJwrEq1e4iB+PnGMCkdsEP+dM
SJVhu+PEGCAVhi/sxKCVKjKF4hxNdDC4wLNysTmbTSDKIBDD3B86X+GBA6EW9o47
rCxHqQrYPADLI5vOAVdMbrXi6wEPJpXjviv28nCcu6zvdJC8yZtWNs7Xm4BtmH50
ox6kGjheAmT49LHe+Txq3aLqSavxPwpyovSnznxxmSxKkZf1p7rPtrM+ZfYMpAEL
7Izx/gAR//QOarCwHVIQL68VXmnqiO0BIjfKbo6P6l9Ny2+mwnaYsvWQgLmxADU7
5fykN+Vgazd5SZzLAjXtWQ4LcFdhzl/HnzFKmKaYkUqkFIWk20jPCAnLwyVzP9fI
h/RoWLGGCQvtUKOimew7UXSBYYF9lKd59tbhOe8KQdmI63z+7t2Zm5Dw8v3ik2bw
ui/F0FmExmT4YGodHc3zb+foH2OgKW/cjPwUJP0UqusxkaVt0N2CCr0nOs+4mvxh
wvU9+8qhbJneNgDa1yLBkXLybHqtdfRC+jmn6EVIutSnPPob1hTjIJ6ScVVgRQmE
txqXXp8DW+f01gOIquw8Fq2h7QC+NAw8eKH+CBLvQuQP3Bu6vOS5m6uCn1SIp6YQ
vOhO2E0VgANBfFjc6x7RiS6KHkdTAS6DPd8nP4jxpU4ngHRQKKFVNAAUDYyDFZVL
Tbp/NkY2jZyWtW9DDf7sq5OjT0gwOLppISFFSuSLcpUpuYzyx9trL9pvYoASowlo
vL4Q7aKrNUcerA7vqWgEOL8PTYBTp95uSz6VFnn7+hyeMBrsqE/1MykCWqA+zJBt
i0Buqva5MqS0kd+cACsr7BtNvLLEPBhHlUpoviU8pixiXLP49dpKjs+K4Jyc669J
VslRG8297JyNJGLelfc4247yHviWsJFBuJ29fhzTUfOiKilZ+zQYBncwA7rSMevE
lnm4dQQxt+BGaq7gHrEtnX/wGnLKHEvXYe3xJd0YGEcvSav/qI6aO2x7b0lWjabV
VLqNLspy3h5QRmy5ZBn6n3OJGzyFzFTDxLHjXZrR85HGlds1fEdeV9FVdMMLeerB
4optpzqeszUVJWbRR9Pt4lu84qHN83G/e5JDqFx9NJuHRpoPmvaSveo7nbSWOC5v
lwcrcFIhOGways2A+97qww+KMBzMKXu/h4d8ZPujvJqeTQr8UpSk97Os7YO4jRDG
BiUVMZWqoPumbjzLm2qA7TQ/U8mKr8gS5DcoeNYc7neo+s5wOqj7tf1D8PG4fP/J
in5/KGJUrYr9J8AHOLvk0KuYnyJA1Vp/+y3TNV657ybEpX2Ut3QvJ3/dyuKAirRI
aE6kQnO+bOxXXZqhtsRI5OFPjvpG+OzJ/MyQDGUPBM6B227cuSXF55XP60cbFGrm
7yxk16TBYeckuuuLDw0/Jy+5JPD2UlPRM382JKlREyYLmI4BEQ0cvgZmGixgDRKq
dScc/1IAtPhbiMSM1XfOsawLmUSkx4gs6Ncap4VoOFxlwunEMoX+zLMuAVOhkJlm
cJ8sj7DC918DzFvXHTJ2pWIHC4xG1BCncFS/IT5cFJ4NajX6NlnmYBbrH3QEZTkp
PGy7ZiDLddwLXtNZgeTcFlVG6i/4cLb53goPiRS28s3NjNiV8+qAhGby379cGe8r
es58z45kmj4UjE05oEgFW6DN8tg5JxROocUrLNbGWta+auzgSe8f2j3EFWzkXn3z
wXR0+yvnN1WwgiHkIyPuncwS97f/CwLU/0ezm+zVDpAFyvEW5hmxfUIdloml8W8F
u+TB46AlXzwPMHK3Nce9w8lOgIutP2R7yybk+8/TqsST5ntS4dfk4W36/zpOqNe8
K3G2q2nsL2c2ovTIk9j0rIqsnpB0H3vWlmS7j9V2T2iOPD5NF3KuoTglfOyk3Z5e
bhf/rB/Ls1LZC0TuqUshlPDczS9TI9TvPBtMlLL1y6sczCS6buE+D2i2+4oW2eIe
zJTKvH9XKAimCyqjsCBW7ZvyHH79hRFBDUj9ED9A0fyN8Y8F+rcY2rrKrlW1NLQf
JFUblCZTYo0QuSutMoJJxwefvSntczFOqyNjl0mVyVxNuyIContMwpd8mjMo31a9
oQZdG6Gog2nd1SatkN5m2KjP1RpCQQu71rAB7IROeaeyo6ap70zgMxBZZooy0z3u
ypSvf+3FN2aM1hzeMCrWorqywzlDsZmKqVQjlH46F5/Y8k5mxQHRVUJdMwRnhC03
paJUV+g1DCqWWxFbfMBSF2vUGgS3fX5y2X/x7/VEbboWx+9vkcj6kvO/xKbbUYJh
zTHYZV2WsN5cMkIAJ+NfI3Rp6SZT/2B0pxtju8Dkf0dl0hGsfijyeFusH40vpfXk
MNWM4FwqEf4qoxl0s7pqYMtEJk5d3efwzRiJmD023MxLlFEQk3KiItkYza+I3uHu
19iZ9Q80kkUN8tek4Xlh4bw2pl2e+TFMhFC9rwP3cZED4EuUHlI9kGzJUiBYFLLD
RED6v0nXhGGv+HPEMTDPNI0GAm9hyUpOGOznbs4hoVy8bTb09deXB4EJnvgo8B5H
ZI/gyqYVys/zQQD1gOYljZoBXU0pqhrqiLLVA1GEjJkQHyBOTBH3fshaKTbhf1pI
Eo7gPwWNhfayIHJIufT7xfyRyYlc3IZh2K1Xu99foYM271hB8BjElBc+zBrSS5E1
JeAxO2OuAW48MpLYcLzpQOWQJcizkTYIRfAhGE7yel1g43oX0cq9tnW0wcmUMFzH
jGQWgJGydiN3g1i9KvHygkD9h7RBvfjdwdD2gQWYPXY+5USwRYjjeiAhIBHNTGG9
7DIlWMwkLA3ODGEauldxvm9mlmXU4yew33Rvm9eotiLPJsTFI4QJqmzg8aQEacHx
CycpYiEx1Ek8jKZO65kMNpEiHKbOnO4Sb1KCkaxo+bfYL2aZ2u/lGYQExVxUWnpV
FHddlhysiHGQg9iI436iR3I/1LRwqn7PdgcYkbOLf2iW6qbmBqyB36OlxGHgHW8P
STSEk+bn06DQpHjieuUqVldYYMlMKEu+WWEM2XLkNqYgV+97bOP2vCS5dB7+H0TB
MbcmATfzBB6L6jkmpjMwOvXTn1NrVilfXCnPwLZYJ3U1pfup/OotyVzPuiVvfTgB
kkJQlhQosjE9Tz/sL7ngQ9NNdwkd5L5r0n38pP9Kj8/xFXECqsu3OAz1MVptTH7Z
4LlrSkHX5xcbxmFYwmkFICQogJ0Ghr0UUvnf9lRc6iMO7Q1JOGEky9bl1KnIqu7T
83Ac7WdRXq9mCRhznrZakaUM3pGNnBimWWBnqcC6B9GlNA7ffJk2b6u18aqL7jc/
C5HJrNkM78SsO5Th/xkkE8Fi4gdtnkqUa/0COv9Q3LDoKTFD8DSL7r4zGvu/M8bM
XIEFhUdgOLeiVH3yIxcLg8wh6JthQXWj67LPlUhR8/YAPYyONTe0VA7Tcgcyzxk0
y1FUSOxTQYQZtFBPHQMJuRd11N3WUPHlmfBRI1R3bN5mWt1kEp68vQPKqJo7s+wz
iwGSpbAw6TxDuCobSVIBQUoAmdJgGv15Evr6S3U4bHv42sx/fWcxf18yIgWQMG8E
srjbudSsUkwtTzmxGkxawdaYwjzMFlO6bNTo4Ev+lnmbLdWvDWuGNtNeC/lsPtzM
lh9CxyC4fdhuSIaBmNzz+OfpxflRbn04uMy5Ywqv/VKaCdl7QiQa36QYNN6W5Oh1
tOghM7i9oraugVVBRobu8D3+RJp7NEERPaBxvZZSumkGF/r4wR4YfLGeDkHj+57y
6zor6JF5mKsZJfVGmy4ljjednSwQypBxlxj1sU/+crJtATvpEcB1p9m1+gyGSAQC
1vMbJwk9AhAimCoMHGrjsYqE5oxj1CbKGEolCxEtqE4RbUTmEUoL/4wq4f+5fpOT
6d07ZGhjCOFKJDMqs2+7qqOJ4k2IDhb3G3554gKxhMOPcKzZMUuca1a4svY+WZhA
nF7d6zqP3qBoSMeVeLpDdjjyotdkIkJAmW22RGoUALcPBO5qqOQI7OjqG9zTi63J
u4Rn2RFm0scOyP66EoXNx9SJs+ShRhiQVEXWpMZXvXuxylLjbzj8tJPMp3RXbFtR
vKQJ0uJgs5FEYJy6dzIP/Y0nb3sZ1xNMWr0UraGGIcg7E6sq3A3kgD3ZNTb0b961
h7E9+5NeRYyXFcz1g9uQt5hXN/l/T2F1cAj32qG22sb0Y9f8YXLki8wydcmnredc
mCGcsA2MybWClAkmR1vo0oG4s7JI5T0dcm8P0kQ/wcTzwBRQSFOgciJRLaEqZlsk
6dMK+hJ4Weoztev1i0oXz84daPCjj0FEsNkvw4y0uvPJtaTjEfiNB8297Jj4UQLi
oi1Gtl0ylmKp1dSHnssQ8SMt6wgKlaA/nsuKsUlwqGtX6OUGHkcy4p1TukUUAMiE
UtEppcQPxqF6n/D3DVBY18BIhFZSv5cP1PYh7VK8g+DTo04dgBUXfzX5Zgeyg+nE
6TMkfP9d3L9HsjWqMp9Um14LG1KcLTmK7l4UdXpDBN9QFoCnNl+yZK9GfZbe4Eob
cymfro81HkZMZnFtdLt2QDrfnaO5REcSo+YxnWo7QS5TXqLUJnQkDHYyuXf5hUT1
Ud1UA0yqfyntM0XLXe5HZqS66gKwkTxUf/NGk5EjpDwcPeYjemLTXp22KOjS2+8m
0FOYEP5GOEDyRSkZgkYuISnNsJfOJsH5CQbZP7OI9Qb7A44xoUPXpMb6kidkZV24
x3MJRaQaVdw82H89YHalxUGo85iKYe0d0uCqlAONTNRa9kjZcuELIMN8nA3p6SIW
imBJdEpr/qOOe2YsflYcyZs77oZeoSbvE+akYd9AOUkaGwoGoxv1D9ClfPU9sfYr
dAGVjf2iaGTA18C1JxSk3oXgUwsr8exRv7NWj0Qz1KLdnUxrtouqB/mWGsuY9l76
tnaHJb6pBJQKzneDbVVdXTAamiohMef2GV2ZusXA/7p6WXiAbeKC/uEa8atLfbp1
Z2HX0060dSYACwdQcx/otsj3qyD5ZP5BFjgOMV2TxfhONHFtROZHGGpuC0fzpHwX
BMfFDq/X4yBTk2SPw9sEGsi7EM8nJU61QUb/X36ku7Uqjjg1tH4xEtH7pAm+uw7o
AfgwmMloWPiJWmRbl5NNHNfzxHqxUpne1rhFFAAFDCWrWUPz7CBcz1v4PuAeIpU2
sPsq5tQY9zFlGsVcUM8jC02nJP7z3pf5P50eRPasX6/c2TUo8UjtWG5DNljyE+9A
TzXny1AXqKt25CJmSZAj7msB80sepzoCSb3mkZUIHWg3aHZT86n4qIlbhGhx0v3q
cI/GbMxrfzaCRLInJiAooui/6W7Zg+RHxCIbw7/BJikPI0erLmJJyrvG4Qcv6OcO
UCNslzgCP9niq9UlJEIo990A152g6tZjArerYky4xMVARyuH17OzpXmogb1WlOsB
Aoboa9c2D8nIMrPsIlIRt2GEWaE0DKpkK7GEDp3ctMBp46yS3FFeZmWy/MF/bBkV
Ohpif4zSL+6Xjgye+IdHelkvlIEmOuAfOIelKk2kZyPYNvsChsUufa5wm2nOY6wk
8koOKVZrscfVL9V80AVjLFs67Cp17apdaqoDVphZNvCEi8EFvnTnIZcBrdgSsHEo
YtU9DDg4XuyEbuCbT0szEYVMoEhM2G/naRKA+9Uucxhp0q2whjeCKgsGxSW6TArk
zrvDtLlCYZ7rtdk7LgNpIfDXZLPSmbLOd+T/vJiGHuBSjL+STESRnapg46Tiz7su
Zr82uZdm20sbu3bk5HH+e7H40WFRjsYDLgjV6VADig0voTMougUUGPoMMy2plIwb
kTte7ld/ppUvJhjYNTAMhMEPygQ5xOPHDx2o+QD7gaZC3By4+vrzfDmMzba1KnTA
EL9KM4Y9JJC/uqmFvhcSXFf+Prtd6GZw4Vo/GhpZXG3ViAtI3Dgf+iHOP39e/wwl
csfpvWt/UN6aPXGATO3BRBozWp6o8ED5uOun2W0dzEKiQQgGTojDtTJ4l+c0K3RK
FsD6l7Q+boQ+F8J+sdMfVd3m5of4lRVOPA3aaWSG3MgaHvN2xge2ZkOTpJ8uKIRa
JUmwSGxRWbWHn8KDsoXzju7SZn3VDUjhzGHwLotmtnzHDjd/fKpuURMNI3QNpdJs
xViYPiYUYb+fQfGHSsqmmZu/kEW5cJfDuC2s2UnDxjMEieUxe1ESnThMGdRdzVba
8y/YaULwiyOphqWG0p7Km/PI27DDZUA4FPCbLE//7l4En1FCkGhpMvlz1PHDBCCb
aFrR3Q5Ehpp9m1tGQ2XJWhOxgFAjzb0K9q2rMBV79/lRXctW7AoHRHN6E+Uc7Ma4
W+WFFXGMT85caNQ+KWlW3T48BH3bdEGvMtFFBN9P0rekME9lK7nCqdzy8N4EKDuA
8Dv5Ir674l6jFANcRu+M2K4tjSKlfcq2bwN/Wnhf71bFTW/mh8g8d0hh9/8c2AUu
HC719sp0DypoeWWDpb5QiMwjROL68pugppUSRtCB/pyE6MZbBkzYE/FCD0aE+1pG
LdBVQllEhAd50TodeR0yrTVldA2Bok77fNLkqRNk4xrcw12B97aYz70FP8PnYCbW
905iaATFoieyE7BfjSpLfdLFDcEMmpVG16o3JAbsRdk+HVCX8f5ParghcpykoqCf
iqoCvc4dVwvL8L/1qVhrI9mH0uTgMnygXPFsEPKmXRS2+j5MtJ7ACee020W0I/NW
d1svsSDt8ZoM1oB/qryQRw0iYva+A2Nh8CNQ/nCh5/tOpKWP95Qszy9ztArdZrTl
Ixm8lUE975WHipHXSMcizZqZ3TfNAkwAR/UZcI3oVCNa8BJtNbdBioQ5rUUpipnw
YZhLioq6/+g9tEcwWw7cdOtJhUrFughJHzLUZOlrZ0otdaq76EVUBoGNSbNM2yim
W+qA4Dwm4gjl7dOLjBHQnAXo1qZxX+ODc76HOhIJMRgHqCOMdqUQUaLBz7lNM9i3
Esq9Zwgx9wBSzUZ1f3ikm1y7cwRAD96iO5nNQLYRMYhCJS6R7YY8dsOuaw0Rjpfn
CEGgjAK+9GYgkw6mavAmJ7cjiNdaOp+208co1s8BjmNBwqynw5+wjiTxlh+ken8T
ANX8SSXRWH2FjRDlB78jvzx+103Ctl/Ps0bzSJUQfjyTb72byHpPk4YDVYLetiBT
KFhDfQC2+0/y2SyJK5YmWkC610rymqiWNPh8qgjojkv7pdVjPWs2xA+iGU5a9aPv
sSs6KD/M+bv6Dv5diPzc/rzaGGa/z3ss7Isr9Z1qebqgizhioJ2MPcIbjJD/QKJX
uTFUGEkAsQhHhj30nYsWMzrr+aEZlhm7EAQuFAuxj79nVrlpimeClZe3O9lgqn25
Wo6rquFlpVXh/6Y5YL+dHDuEMgG7GPP1W0cUwfq0JShthkai/pXt2J+wofl3SlU5
0MlvB+13ikdIX2d0xQUvZAv3BxKmn87hl827I7R2Zx+DJjD8ZSygrknXTNvRADGE
O53L1el5c/fu++reHexGyMKf57nJsoTtfA9ekjMtpz4gT/ZJUp0d/r1CM0bCnuCm
k0dVi9+l+MwAZ0CUHBarBZlNn+F+0SgnlcurS+KidaaDLKkhKhn67R+AcuSl0mrb
XRObatrDyjBOtVn/qHr7uXQja0nEOnS+8H0m9AlKHtCUvoBhcWpceTHRWcY41MTh
M8v1ovK+44Yl7vMNcUWjXXxoQHQ4kOEe9bXfT9XwrOgFiCuI2QKHVn+Q2I5Wxsmv
Sn2kXizKWZyBHjUgUHHG0MjrYDeuUtLUP/V6ZjdKXnNbHGpKs+/4QiOgM4y8ozD/
aBuMY7CO6SpKywXPlO34UistZ8jqyh+AxCyXO1LEGBnR/5WxyKtBcAbMB8WRnF1X
SZRINYowC+krinNA0FmdHKwBaYFmLELGBwo/b2fIRcCFVeKObwSI0Qgs4pjHMMea
nSS4bySXjN+ZwiL0HNuhT6mgCDRy3fWFEQpUlu4ERPE/ZdQnZLoOhPRGEZPXi2Jl
p6/XBLCkuVid2hITxhtkbtxD4WAt6HFPYdiz042Giaz0wdmGxfpsgQ5DFhk/xskn
mm62fWPG9uu52kaIrsb7ugM0lIwmAKHk3xPEpIzEd2PLdKN5yHcMTfvT1L68jB7d
Sl6gpj3Rh1rEIC0EhnWe1mdhWyDdcZBuyqejFLaeoe8iVOvZSUDQf7Dytpj84Yrm
xVghhJi6KxmI8tyPSKyqVW2Cy3Kgmh3stvD7w6z/1WJ3l6H7izMuy+DxNtx0OGB+
hGa5CdseC7pI8s/57/y16JjijgqkT38t87TBB5OUjzaHd49R7iDNgJoygHEBco7H
fy1gNv1TrLFgfH3PNvoSQgViwBpMl2e+8DaQmgji0gJw1ogfV5Th5rx+cCHCgFHT
dwAYAsGinEcNHOVtQWwtD13vJRWXn+fCpAhdq3tGq2tlIXZ6cbOhybf8HMH+20h5
hD/ILSy4VofSccRscnH0CVIF9Mck1FPYjrvzpoT7OifgiB6W4zrB98Dyw3dRGQKY
nCxB4Min/eMepCKE1VIm22Sg+rjj6/Q2cy1TD9L1lmAGVmIR6LBlrMIs72YKJFBt
6mTRy465auVY/jUkinC8o5E4BH+Hx0Gr7hvyW0HeHdvrBNX28ZvBhRbQYJ6aQFbM
gofmYcdQ+nICzlLN5V8wbCLxkSsUUz8rabbncXOKVnpC2uX7UDIYP5HJQbwj2maP
4ma7x9awYSQV4J0GGuNsAYHCXpTpWvydWISvl/AR9eYxGZJHRuMuFdU1gicvntS4
l7j6Zmn0Xpf+buhbm4A7gXfrnlhhBdcYpcqyfcmJ3c7Re5axBHdUON17uv3Ed+Sk
M1FWn/UPgg1EYhNS3/jKxPv3Vw/nrolzxfmKPFeXcTEjxzqRzYVvv7u32YsMuh4E
sywCUyy+4x2WQDwK6OYp538s3J2xvGy2jxlvTeXFgDMYCrG9PP5PPEVpD6Bmsgsd
Jt5a+UOBCiDqBHDRirDx9sghuzFxeGkCcwCeAOHxtX5gx+YLhHevJ+mudvOJNzXO
AloOCP9+/c0zxawVKh19UifOmL3xzg5aUyTQtjYPFhupE8PY51f5gmE2XS9CpPUz
Be7fKaaGuH7PeKH9e5lLdsWZDd7+vN/7RELS9qgaTrq9EN5YUNS9Ybhg+dxeziX8
g/H5qH4oNpAtEM+qoZDTMv/V0QCpUW3nC4pTbjj+JmuSTfsHLGShwd5xbGDDVQgp
gkEmTLHathlu5vzdaWJybteAgsZz7fn7YOWrKjGxHWGS3AWgtMPq0mSp5q82JP9/
T79TDSMFWirEyK2z5VjMXiV2RZXm1pm5nQ+ztF9/adtmXiG+CYpoQgVP3DYXaw/P
T9FurGdFIcz5J/I+U/xYqCx6LKjTIb1KHWlXOI79Ird7UWobpRoHK4iQ9nSzrPul
I6nbayZ8wynxRR8G+4yU2wLAnZu9QXL7GFYcedgPTCsHhy7cgcSDRBKtXacmZ+Td
8E7l+XyUKaV0Rg5nJf4h7JZN8KSyBgQeP0xsdWKdoZ35E7XN1zhomiqApw0IRIhS
3PrtOlKLr2R6dGhuPCED+0QRUGSJq7oqS7rR4NQt2H5riIeIBGjBfCt8X/wkJvPT
CXxSfF17b4oyYWyussfyszN1+5Zceb1+QwXkEBfX/FINJ8JMO6ah/EAa8it0AB/0
TjgRj7mIJyR2R08y5uClm93Dl8cE5UqcqrUEILEggf5T+XrJ5JDkNN1RO3ua4ang
afXxPSYSYT+tuLAY92fAkvn/NZl6OX8Eic0xK5Mmx0tvpfUGPG5rJcBJfhLi9xoG
8UvSiQavRhOjQz/62kXK3gUEfyejE8bDPoxOkTdiYTdYtJrHhJiJeK3qiaP7Tyfd
ufFqySJzGNYK8qBfo1E+I66Ov4nwBDyT/ZTnbZovqlAWHkhm163minemYchZK+58
G8igXrUZU7ZknzgIG1Xf/iOTDDasHkHamZqsbE23PZYdDEXU4ulCsOIZZLCzFbC1
I06+bgjF0F8nlJ7/UojRKWWGu71GSILO6bgU8n4g+Gkz/Rv3ZUmSvfPBYrI+2QGT
lsNNY2xM4duht6zEunoWpWjt4BPqGsbj37mi00PSbkkSSCHkxoNADqpoXSK5oOyC
btvy+sAmez7KSIw+iBsmZrZJs14UYA4y72dvnGtK9+nPYtyjLC/vLa4Gy08XiOJ4
EevHf/PFvlX0Cqdwe5h5BEdcL7Omrh5YytfX+K6VG6MBV0sOszMxxB7t9PYRC50I
Gws58MRVrV3Aso+dDTus1tuFTeHnqJouo+sKbKCehXJxekn16NaYzSodTwefRrJI
5nHwDDNlLdgXZCBGnpVmPDWTjwkOLXbLVf7hJPogUgYwTTqABc1SVSHlb/JRKAQx
bX0lonuNt8nllfGJChD1EjV6AnLI6xESIumz+rXYucDmtLZrach95/BtE4fbmGxo
FD99Lvx/H9ti8Os51DCMOccST214mtH4cdj2fuRXGFBK8SruYLxY5aASpXRUkxVl
1/f5XHozgn+9kNpAujwgNg0W4aeEADNH2IZtxoY8jWyivZtrS5hbceJLGx+vE92W
V2pNmAeCaLSH4WAU0jEOiDBNHnHNDc6zQ9PMFhulUIpeVfexxpmw2UCjunYfglAI
sqMooPUX6fBMRZoM8DJ5P4pNLfWNodomE6uTkfjpuORjlmbqA+nuqQSfC3QsAbdH
TESyhBAoPnpJEUAu2iD+1SdHMI6TlWkoV+3lzK4aAxOVGn0UThbxP5FBaT2ZmtTA
vJRQu/FbxLUIAYuthqnyxiE2kG5M6YBkboybqr9r0QkJMxch5D2uhLjkaceXAWOY
bQrDubDlR1m56hNKt703T5CPXdsjaNYjUAj2BZffvK/kTSmELC8NbtBqZotIqFSS
ZIn8QPICo5R/5b1sVCsYCKYSj5ewLeedVuWfHqdQN8iI+a9J1LUG0aU0o6ZTJmTY
oONaMOsveQTa7guk1Fy89WHUqA1y8ehDCzUO48eVU/Wq9bsZbpa+40GO5hTDwFBr
6FROsM8h3yfI9Bpnf2QfH/ASj4OnCfSQsUsLrOSsnzMqtcgxjUrxYu0AaxAX4zYB
t+RbsBrSv/+YHZSst+49l7wFeNPrt3znyo/5OWwuUJRTxnFtqee+gzIJdA87Ihme
9G3FachHa3ddTuTQbwaml7Ix95NDSEjbZJujpi07MIC7FhgB/qm8Dmdt6K9gFKvb
SgY/4N3SI2sCav7o0pqRYWgNie4oWIcMBQiJqxSDEi5V/49nf22YDfctDu8huy+E
+x9sMLt/SVz9kNH0L+PwmkqK0XmjlhI6KBePTOx8kaIHJMdX2u4pKDcGkNXivWuW
jixBlmAyJtb0jfSpSEV4NH2ZXMw8O+4M8gay8ilKuUYJYJV3IoAmlDQMGHEaZyC5
SUaXHgkWhCqx3LXiuwc7k2PB2bJKYqtkK+FFfdE7VxOTE1SukSY4waETOS6/kaxd
wZbENDGBXB1LIc0d54F9+ZazvlMQ2PvEMkKHCvv9xLXqF+tSFJTgpacybdiZmGrz
cWO6Y5b0v7aM2E78DF+VbWaJqSxRyTVtieickdpQQGk35XDMcF90C0Toyg1HgveP
62okUpgJQa543TePQNViaLT2rHSmmM5w75j4rX9ux0W2X258JEW0UyLixkcAwndX
lypgDWBwr+/cwLmpcj0ZvBHUIaEWWeGZh6ZJskEpU/kKoQxfCDOPvjVNalqYY7VA
lI7/sunicvHt4CEVdOiEt9y1dYGN7ydLJsQzeZSZnAcVqiD2JP8/oTLaubcDAmnW
vjm6Is1Zbx9Iuyob4rwh592AtqesfyPt9E/c+Ozm99qzDUFoK7elOL5Gw5s2DM70
wFjE4Es+o0PswFH8PUmL+QPTuGkatY0zPx5zBHZSbE2NpqH9Hy2Oh/gxoJrj6hJ6
PMjegflkrFFCCb//dve5+LMw5r1jYHgm0NHrmvrbLZF+PfPPnrIgqhXJM5hsSCoD
SeB2/WCSKHtOxV8L4jX5CwJaWQiTJwc8Onz8loX5xzygFziMByCpkpFmS5PO1Hao
d7/irGebshFBS4U8BWXc2rvYnCNYem5Y0P9lYNo0A/XC+qMpgPoiEotGj9fRHlMk
3gpNokbGLUJQeDlOgA/SCJjulBDUP+1dYhKv3m3dpAtVCru664HaVdJTshCTAIUf
eA7x1ogLfd4E+0f6+aRcP4sEojc/CLvty97wTDJkHZCZMU1EgZHu+TZP1mL+x2bo
+aLPkb/K7WvTPjrr/sHiA8xifG0lkY8w4of2rx5JCXsh1Rcx+W6QfIYCWuaeF49S
nibIibR2rsGxryBLgU0fQR6AAGCwxkU2fQ+tFjJq5AXtEm0zTlkMRQ42pmvZZoic
nxs7Q8SUWwGymI096oFIWIu/k9Pf9yfgpq9n1cfZvXs0CV8Q7a5yS4rzf6typMjg
UN4KpzsqqDFVklN0vXxHnvfST0Bg+cPr48Lh0DcYU4mxqwYLlsQc9JRJIRKa7Kup
Q9oFkZ178CZRCyF7cMTxmJekSvAtqt8hfzffBd0xmeyIy7zkCaQYeQBS2yFlvRyO
q8F9ngKqxezp7tpw2qyQ3A32+BjFL9S3uyYC5QahCpVRkiwGs8hhR4IGxGk2EnxI
9OfI7lBHr2TaEvH4jbM3stdxi7yd2h8KFlcrQR75BwIvtWVPQ260tZR5Tv401+o1
hqP/pvwH75vbsEZwJqK1UhAf6efD0qoDP5bcars18Ufdo+j3v+t67exeZfqNmg6/
p06I2A5svJ6iz2ll3b40lQQ/4L2e1zyVyFrwY0klT14F15/kvqby1QnokpPp6dQ+
QECaENF2yYtiHRW2pQZmv7wryTQe1dx+9xJFtbubjvY9jAn4zctRG1+UBWLd2gSt
ax2pvxQJbql522ogPZvmSRPwAoSx+LSDnGVGq9ig4px4YUSVblcfYHc99tDZrk7B
BK7Geus7uL0sfHLemCVSRCjXQ/fkJ4wgA9rIctzGwNK7aMqiiX2YEisDLEp9oXNh
WA8ctfWX0NMDs7kx8ZmzJbpjZzV8iusIGWPGOlcXa26e3FdmY7l3awggdyAoRomf
RDs3FRtwXkvqNmXaQulr5MVCDKeqfZYR3k3lCmuxmM/IXLF7dtASSVKIcrvT87SS
wAjVdILtZaVxRFrOaRD2WKY90Fka1I2NLy7aO7Oiblv66lyv373C/1zjC2S1I/2Q
7Qnt1UhKhSncuBmSClE3cCX5qSpJk4IBFYfqreCFjKjAQt5ad9nj0rdsug1kq7aS
HW01iDV2u0hVFDdez+pessiplL3+kOSN4VRbLIWPe0jjOQQPxPTK9UftXst/hFYk
uGN4BLeJtGoexR/HjtepzXhOUlODQnlBIoZhUQOghd8FTlRR/tci4oiH9YUrhyXq
FrMuN62826PnHFDxoUfOp9zew2rCGycm27c71yXjKi1K0FzvzpGRAL1lVyFEC9tA
YQRrBgpkGbjXfmg01rBW4HlIh5fuRmajyyB2nIi3eDfzw/FxzcMI9x4iEupEJa25
FjxZs9viC/G92iNuW0qv82kEEjMdc10ntIr/ZEvAjiaADkdF+fsdxWnt7V74su2b
vQSqasHasb0dOdrVlPYT+Dc9ULYDhfmhBEsA7AOf0y8U/0QRqXDZ2SiZkQeIfJGC
Rw0L1Nr1/42ebXAp9DtLH0zmTilB2f8+D7/FHKHu6XIaU61WBHMxKQBb2enh6fGD
iOEC06uTqSCqN3+k0coGDiP+OsanBOdBFJhswPG5M5PcObL0/031GnSLJazFplUn
CMNdx8OthICekgTr2wUEyguyllSiMU5ZisGznikdu3Rb12AQbrMNixvmC8HYHBCn
ajENK7W1x+rWn0mB9NUeVffmgldXiBCo8HTDns/aCJErYJycXteaom9A/V6ZOOQq
Ku0/zrRJ2KkJu66wtrhxRkwI0193X3etjKnPTTLu3x1ynx8/xrA7f5K7Uw/2xAW0
+XyBuINR5BFccmc/b5+VPecR69hi1Z4czu/FC6wYIsmTn6fTI9z1h6JrtzXiv3Bf
Wsw08Z1jiS51LKAf6I/Kb8Cs5DnGUhGgHezMgFEUtDrLaSGywTp/qakCBcFy+tf7
hdsADJprzvXWKMNUVbSh7hR3szpsik+kU6RvNiSXgY1krEvZkTKGHrRiG1jNhN3l
rjTLyxW/J+YxG8G2+EJrrZ3/OHDr0LV2wDzc/z6yI54PV7CMBKXcR+60FwVixHwU
e8cUSpcNehLASzcMDk9Sa/wTFqr5GASDVnu14oTZsjUgrU/SRfxqP9qJ6dRjCfp+
hbPJ9fr6rcE17JiFl01nfrOYbJZ1Abws71we42FluyTPxHaxqnqvpPGpEbSLaWLt
rsgQSXOAqxzXhGb1kGlSv3A6GxO9mIvX65DAunagdKpKISxbOAS9z097CHT/EleZ
viqk4NDcqoE9FhY0mx37cxEakFPlXRDtgbpjlcNao5RxmMKT3pcAv57felujcZiN
lVO3vbw8Yfbj6Gih5bwJIdnNp84kwf7++3F0EURB5OgwQ+EKXmsWOf8DGk9VGCly
pJPG+1S24i65B9eqqN4/nIVjKKsktKJekL73eV1eN2K71fdt4zqC1vkIaZN3Gsh2
CYiatWiaOvAV10M7GOiSceSnEIFlfrDBCCbaUyxB/b7tUxhGoQim6CMASat9s/37
05UxxJtQ9CtJPeCpuQyzBf/Hzl35y2Rf1vepXwBVG6t5aHXH6atxNLdAeEIHOgcI
mtTxwLYMK7M1BAOgnGVHApnGuAF8zX8cPgfr3VAgq0ZQ4qScwGmQPXfIuBFxuVc7
iCm9EVCwgfXx7D8bSzI+SJUmN13PQPiRi4tV/EiwNep+TEYHV26adaLhzOTPn9FZ
HpWOc2D6epwxYhuFjZlpZp3PT4Pve11RMW9QqD2xiyEfcbdXp8yoycbk3rWcTBTR
il4QgzELpeVa1cx/8x7PUtl6LaGMwRuBz8Wy3aSOg7yx1Qh0ENq0PIuBZNTnTUfD
NQxqiPk2I/qHb3ESF1RoOA12CtS2tQ6XOPqRItLMcvUHDQOOxZp2KbsE+AWm4pCv
D5QaiK0VioHt2Q89L+HCWfPicbXR4zd7DgXAFo7cxCQ4SsdbfH5w4C4XLoyqDeWt
L53veDWpZejA5IyEehBAl6CSDdehWJUrK682qKsvwGi3lkEttM9FR8xid17QNP1x
89VDflncpJ67sqwVpieBWmEGcSpaddcyCfbq6Q+Cb+pQXhorvH1b9R6AIdltw8h0
iIELbj7oL8SURtX83gIs/fGRHf6/aZXUgzl0BKuNZYkDMjAn0wyNwDukbDwcTkg2
DzwK0UCYrSrtzOrgkf5r1IKO16Kr9qz7vszSgcX+uX2rQc4ISQmwiXGQW8xnzg8d
Pb/0q1U37qdL/LufyQioNENvNEhzGu3x+/saxSDqocQfvc+yuO2L71Fzcx2m1Y64
QkZgMfGjfktXEb/R0OOSSy5uLnoFfT6asByTCVdM9ehADkm0uYdSQo72q3/WTvkq
ckMElFz17yI5rbkRR6yzNUPeULUZrGeBT/v2Uc0FjlA8BcxelJ/ZthbQaXrlwglf
JDxwYkeH/PtLYez4dRMvuaOA20rVAr5NelrZu9YJVWMmBZtn2YFbsPgtZR8i/SF7
b7lbktSizn1s7VdqWfwfRXRS1PY131LVdI0dlg6J2U6EVeuNeDEZQvmxZs46kQbg
7H8EUOhCtx4+hOxSkjlc8pI3tcwbe0zJYXTna7niEd67EzmR+l1WV91FLsEoXWBh
FpKzWkaLCXIjGFg49LZm5/dU/JzuiNpMQGkj0auLrCeehXZt4OTfVLmOPiSEZMLK
3IyaVM6j+goGeG1qSyGZU7WXD8PPdKQ8wHp2+u4x9pbNhbRbQKb4HkPO9+CbYSv5
aZgt+Z40V3Ti1iBWkoFgs/R1apcAXEpEUyMA0U4aZ2+HGxq16rs/GtwYyVImQgGx
JW5Yy7m1yc2JqH5h6Pa17ROXfzFv7DkBPMS5hDQkPunMF7YfdrDA6IzcL++25rWq
x+KU58EQQSG1VGTxrYILQP5dM4aHBAw5EP+f3nkuTn3lM+6sbxo+iR78q0e9NEVa
eIMoOdb1XG4/o5GGK3bSlvdkJd+YPEPKsJkNA7JTDt30E4toR5zoDJS/lWGszPUI
eUexameWUumfxesPa9EfV4PPbenHASR4VbzzjFL8EU5s5ds7PANYh5E5IDotR6Vt
rU6XJAposKGBfQyscag95s64ROkoHaOWG8iHQNszQzZVbBGGEEOdX1rx+Ag78zrS
1xg6EWdLFHZfP6utn1lPSUinfzQpfzUec3l7XoA6SxV2eVSr6kiFZNBs1t3sAwqf
hqdGtCIa+o6XH1JHvbkg5fXHmdPpeGsRSdlTSWT31LdpMuDmY1Dc0E0/CTTTDZPf
KUB6mobo0HRBQADeN7sl8QyWTHgu+cS2lC3BPjL1/lVBXjhf5a4YAkl5HRz/uaP5
aAs8O/+wfUmC5BTaZ8lg6MRN6zwMi6gf4xr3MUESw2woUdfovR4umtACZ4KM22n8
/D2Fmp56DOKSuPBUpKyQ5gtkdJKclJG26fsrEPok2+oaVGG1y4qTPIMEf1DHgtiI
dfIKeFepDzmvM9+ma7H8wP8pGyEy+Qs/uLcjYJpoyaw6t7eJSPnLmMdLcLGL5xye
VU1igIjqxAZT782FHe+2HzfvLq8A9RwqyjCq1FZ5xT2IX0Zp1eY6dtrVoxoKh37C
dMqDIUjaQjL+WVe8sdsQ+JrJGO2sGqLUFmXgLNn0BP2XtLuOqK21cMRCq1dU9gug
ljGTNBoUt5Gez4/QK+WsEonA9+Bm8aNEfbFFdc7GgAXTncZH/dMz6SrUBZMq5YbQ
BJBgwIrGBbmw1EWSVcKRqGoo9GfJnjhWIM9G0OXfSfp4AQyQeok7ql/U3laNtEeS
BnE8Y9+lWc55jgJYyaG87KEAEtn65Bh/lQLTNR3BEXJ2jZi82bi71FpIsC/Dw7j9
/Vu7Hx+2UYdYACPnwgjHT9J9zSVryPQmZeN47AWVcom44yG99KR2c8oDHCvT5wza
ET5w1UetuULD7IevL7j6oGU758cidgJBAPy/tzLNLPsqdLT40mmN1ABjnqyC/tFp
Edzi/ZBZ8yitJFu0pqCW0QfT+HPOf76tysACbeC5vRtItD7sdjoSTI2SiJ11QGj9
ki+UVNQI+pEP7/KCgLE7LNdIthg/H4bj/Fq7l45Tt3HGU0qjUfTwCSSguFaR+SHr
0tajmxLOmN2R1t2+5J7TeprubPq+A846VQsqvtqhPm//gXSGOVJIol/aq/Lztc6K
nlTtVYALgDGI2UC+c2hxM2hNC626QdItDdTTJ5TfH7oV7gJBL+rw71KpTQlVOAC2
iBVAL/ODTZQhXdE5tAgJbV7FaR/uGbrgfpaDqr//yPAU5590+03jQELswD+GbkN2
MWqSDHxRtJd6aEe2Mgf0y5lzlH5xnvYMVB85lGVd1cYEqXJe9NfAwLjaGCMREqOv
cmbMbTciWNpJp44WmQb6gMQe9vm0Uh13YP6djiMT4arb4rARL50HOMN8Zjtkg3xm
5EC8Ui4UIDS8CIDsfVctWBiLGn8SFgPwF/6PVouTY4ugHPDKcTNGawiz5BNeENRY
LdHubgsFdQk1QYbI5awAiJsOQdP6UBf2t/cOyBT9jD5Fk4J7Gfnk235BRbA105be
dTDH5xfDXKwxXJeHRaq2fTaqPQGXsY6spqWXDLkCezAnJLSxcXydQG3kCZU7ZO9q
zLEJuFZJ15M3/65iMle1+l8E0qu80qOw0hoRCsQ4ETuz1q4/lPW/8ZIWqSDG1dCI
skgCrmMIUaVHjR2ul6/E+5aHz3HtuIXRQaKSWjye6iZAeMTG0oYXTKqF+NbYnU4G
qQP1AZn+h2zFp5N+bAx467unIYYDQDXUV8RkUXvWNV2/E+wpSKWKL62a315mU9iZ
L4b+HXAuK5ZBYwc0bWzI9nrRk+T7dbsi5kN2dqIV+dgG7GsqHk1/A1UsVO6IEQrz
TUZVYbvRF23POMHYKGszcQPeGz/hYoxm9EHXqN/63qsiVW64ngQouTN/kklVRkRe
VyrhqYxTOrbUEO8tVcgxLK+Z5HhovCe4X4d27f9Au0aoR4eFRuFWrmhZSkR5IGC/
0kFuwwbDBLaRq59ub8x8d6gIKFYy0Qk8Qo1AcVxmYmSSShVwzorbQdLYc+Zj/oWS
MIxLK0rSZYitiZHgI713z0SbpWfVOnkZfOUV6FPB+wfvFmHpdF3yOkS3jfeqK7Tu
zcXlRPPH8uJddndPPuMVBx/RSlV/GV0C6FRAKky3gyijLN9VBeEPNcsnciPoyPYM
XFSKllDYdDnaEnYr2FabT+nUn4dF1JX7ZdHiiJhu06id7m8MHFfHKvMLcJe1drCg
ZeRabvX2glpnJ/GZhfTiaCfN8aEQCJSs8IlGeYtI6X3edtcB4L31a+Thc6rz01Jw
37h3jNzJ84eV+eE8bJpeI6GBmnv/Y+mJHM2T30KnsbVB/H1DjbpY/MiV+Jq5U3fS
T1MLxz4dBT5dQNQdmdR85i9hhquvdFvOETYR2IyBybHG7iIH9SE4keQ22Ano7irl
iIuis5j/2BygQuw4WVZP5eXPI+CK9gVlZO/nopMRalRSTvgaAC++KJi4161QOWma
528VJi5MyLPmROAR/flK5j9g92Dx41gauh7C07R/V/Uvmst/2e6/lK1RVzrvWcOP
YGAUnJm8LcP+009zq0y7qEXxhZyzyqVFUigCBTOTdxtc5Nb40BvB90oyWhzLUg4e
S5iCAX6laCR1RhvQzNULwYuFlexF73okcdRiTLO6IRHH6wPiox2pVVrcaVDK2N0L
RSPfQqe2qe38KLX0JVHwBpF3TBDESHjrxWbz7MY0vRPZH1bJ/KPJKnBOlMizVY/D
0N4LIOJ2S2n0b0/gm4CZJXrMyxki3IO9UdAjPSK3/blRPDcm+poUGWwLRGAF5pyV
yazmcXM++H3RY854tllRjnphCScE/uzrFryy7YkiKL5DSlPQ/A2yFcVJrC6WyBbi
Hl4o2cKnE03RTfOAgCDmj5fnteDLE/m+mHYFX4i3ab511m9va/EhEvdrFf0gcoTG
/iqjN5yt4x/wOE/lSqd6lqqriqWv2ebU2E1T06xdBavdmgCim87rpmQN5ZhPC6Rl
xZEfYI8OyYRjZ+6oFv2xZw3EMi13lqr57bTIkT2EsIFRNC1Dmz7DH0b0mFQV27bs
+8a++tSoaYVdvC0eGUU7T4h+Q3CxMWj4zB/8FECzaufdy+4rgyerUQKiHrMbpzN6
aqU0d7YhKpZ0v3/zo0Xzz96AMiojuQCBQI7oOoQUHiYb2kVA8ws2xEc4w+E752qC
W4wObfy5waPsZ0ZhqUub62WKEIiZxp+O0/82bG9f5uoGth9xgi2Ogssyu4j373uu
23RKE91Y7S8wlzJMam6z9ksrUxCdR5vd+m49xxzB4cPSpOq/9fROAnN8pg/xWJbs
AyCfYgUXVyXkMaZrV68J7plYEJiA9K6rkm8TCpA3hq1XURoyPRVsmbtSDXYwSbcD
N7X7yD2izyEWm9uV8sEX17cUTgLmGSoMaJnlxynLJo0sC6ExnlynI+aEDMOK9brG
qYBs8ltaLDouVRsNa30Ri1iOPzwa/pi7rYHQrNY1bPcIKxFF2QyodIQu5U/XDJ5n
z7H+VX8MEb8D+T3nRfX6oMJTMlpy3WUUqOhxIjTHqrED9k1GUrTwDyipMsN/JPrq
pn8GtVprfVRPoOEaQw6g9UrWK9bbRkJeqFcBtdsm6036aWDCP9bSnRUrVxIeMwX4
t4yjIZcJv4rLhUkKyS+wuG3wc0KsY9p7NWVC+9Qgm9d44F4A/51ACOBCI2abUbCQ
w/jAwlH3CWf/ozpH0jJCEqXHQisAjM6phvAvJ0MWDLgdoXURyf7L85QnPYFpnstM
xGpI9MgQXlTwdZiuuwGGX6rRRMqfSEAitxxPQLUr06J87yHOaLy/ZQqKhPnEqmp8
e+MXk4LOJE8FfHdWkxw74IpwsaVVC7e1mAcPSmZ055WR5Xf5kjy2Y0wA4ZSKodZg
1bZPMufdZ7vGBDiUiJvi/95cC+G+xRlRiBUTeyJbI5zCcyhLMoggb3x2ZBszYzEc
UIIM68/PwSYHJ9FhN4AzvgOGF1WI5VALU4vmawbCaXecdMa32+jlj+eaxNNujht1
EER5FxpQqk7nDXITgavg5VIe2FzOn6WWwens85vK9I0nSqtVVn4F7w/LqrY6uDAr
kAcu8W5RVMTm497IM5G7c4G9oX/MTh01tUwBOs5X15C6efE/d5fG3eIHtPjlhWxv
09Bxpl21INYgexgHK92V0ESKJXO7IOu7X2gYiJcD5nefWDaU3J12vR3vvhgTeBMy
MxwzL9ahOTnPVNGm0odYQB2GyJTxNXb0xTv1CQkOrC52rydbwV6Y6C2hodC+TZ19
TpyCx5sGAva5f50L7Jmb76x8ZhVOmQXLc7JqvxhnIhTfgUloKJwOPC1YZjc0to1A
8AfpxIQkx6cK4ZrXQ567q21Y89KRxWBY/pWW4hRGLaEdD4k6Xbnh2AR2vKgKOopu
RZPE9bg2Tkv++Tx4mxrR5+2jjIG/N9xLU2n6UZggTgyCNrLWfASkceBWD+gE4xgv
egT6UpCCrYG8lm9EmVRB87yEds0f7BfSAcgdThUBfapL7iUNqYtf8yD73B7lFeng
HIGO0it71wVqlbsLzSLgoE8wEU5myFWkAinAvcrc+YQq5A/ob68GveipZnbb8hZj
n1dyeZ6q4zJSR2UErmLpIytJhHogRYAMYgC06JCJdlO5DCF1+jdgu2KQ4BWZLyYR
FssL0WBEbMomduXGWi8R4njDQI0n3o/v/YspXqeMxOxmN2DLFiYLt+4h5kfQsUxG
2PJOxkJOpgrKg7NrGZ/ftDBICFqR40h4fybVfDl6MO+vwZnqtTT+ujN6NQWg/hw9
VLA5Izu0fqMmZMFdnjmgnqu4MxRwmiEbAUp80Ji4jfK45lI7vaBXmWARJN9oH7qH
QYCeJZH6tt08NLrq/44u61njdLszzjlm9++768zNJn/G9NJN2K13x5mXm29uVlFx
DtRj7QmKIJlPxkT4q37DPKc/GGrD8ZXjSLjTQsT303sDhVROnrExLlue3MGr2u1w
ZggWwVfwhxfEVyGloDUmEno3iXyF8d6CcH3PsKaMj7nojig0S0yzVVG6RNvwEgdC
RuVOOwu01JYf4eJIkRg8Ssk9KzTNT6SRFpwGOynD/9fEUXbWLHqEn+GGdUKS3AKp
stq79mm3MUSR7zEit54yRfDgQZJ9homO6f/AkYQQvYCAHv+gKnP8MLuqz4kTyKZs
RWML8Ll1PtwLXj6oUTHVhOpnW4aUe9iwvckypJNPONw2qqTZl15lLRqJRXcGiIQg
Q+kNQCu+0CMCTcwr5Gl7C+mMroBZlcef26nGDVqmJ8h5Yi+iV45VytZQ39geKSa1
Dfn7EsjMqYPV0mbHX5tm31tL0uV1L0C+vhyevzlzW1yDIGHEravexsYT8Q6zmD8B
3sU9B+/eFVfR0lK7KU6JREaXuRJV2v4//RhrrXybv7O9ftZObrtSr/qyBV/+4ZOq
0UnpisZJk3gNZqico1/CSec6xiT5p/DdUnMTqSPZBCx+ACP21h5RNltSyHf+NjJp
VprCO/bhgGDD93qFqi8t++EY6HyAPNzv1SRyXDhR9vLsk+3+05ZdRq4Icur4lsC8
zy7bwAgITCMn/qX6/gKi8hu12UpMAJnFOoXLs/iH/NyyCFnYCjc1ojaj/btNETKl
4NeYtT26flREKoEagyYPV9ePrxznXcC6HIf0vsVeyeRkHaFhYYdp7uYKa8sDqLei
rzyMD9T3ut6rvvtSwUCNTjFyXhnWCijH3lkMvJkekP1lGE+qkmV/oJIGf2gLvzvr
ktgP3CFgBKBrUyBvY4qk8HiMB3XXPz2/ZymHU+9gx2j9vIhFrC1tLBQslrvH1oH/
nIrcp8PBQvHxJnlw/I+Z4aEolMNy8mevYe/Agjz6KgtPpSi52P1xrudvS+9LnNvU
VdJp0tO9gVBTEGyftIts36ZqF3wV0CxEqfqVXzSgi4vA3FgGrY6AXowIZHGI48w0
h/NCaxnuYCDwj3SlfmSBRkpL59+hZ54LOJoZUPgnN3njr+yeQC3trI3SIA11KOUQ
vtq9cPcZOca2pUnWsCIBzT/rDWpJDq3XT55WEklSd7x9XlRp6wB6XYOCYY7rfMNo
4QbQQEZ11QHjLrV4ztpkiCmIo/yQ01iww9/ovv9AjImKUQumTfnvPOaCN4EDtLjz
p1nNbDntm3cVgvpueJUyE6hdsoJa5UpdEPsGJllQCI322nc99FpqOpt+/jHnCAq6
rV3TuKV7ly8XkZ8eflg0yv2+BldkRGgSEnzl/XMQJ5XRbXJjMvfkgLy17bUOdg3h
CKjObOjE2YW/oWsSJe+Goo7w1/L6GPnvZs3mfIJ7Q+fcfJTCF7Kv5aidWQ4NK8zO
tmwxNhQr0sInerZ7Qk5MFVMgs0WGSjVxlit0MFudKZlaYme0GsdGjCKoK0Lu1ZOh
UqbsXjVlM13VDTPrVQ/L7AjUyMdC99depLRC+32+XZVroRQrPNxa7sOrAWo3PX/h
TOArcz6I42D3ewfAyt9uGbPqCJOB6NYSj+Jyb/sGjtH1SfvDoAsG3Za+qKgV56nL
Ybrj3O+RxQxe46H4rHvYlzLKJxaoAeRvKjOkx5q3UlimWOWsRlsDgOPD3Hj9lmMG
g9MYojQgMNeFBu/ibHPGlsXkB/xlMONelvcdinZxc+t16pkDvVFgwOpZqbywmYbP
S9dJmnv0VvYWkO50vJ6TH+QCoKMcKvlb+x8zupANDzB0fGDLBY9YzfkGyjkVEKCc
QeBbdqEbKbKHNsKc79OifX5HhTEELJJJZH3ieWYL26Qf/XPgCdvqY+EeKkTAfRD2
bjq8e0C9QS8sZRnRORPEn0Jkw1nXfysvgLEDaxWy+tSbkEztRaidqain8paEN6tX
vTKnKh9gupT4O6NmxhOOiLspKSZhZQOZG7oR9uvAZYll5ErsoUY2d657+QbaS51E
DGsN07A+9xutAnqgI2m/2vvgJ25hpCwFltzVHRvEGW7eMo2dz70Rks3hwy6o7fcl
xyt33DUL75DpOkrfqzXr0Ye48u4M9CJ+F1MJKAUBmigJJvQgGDWWjhYUJAwshZhT
vLdr1NtRqhfPoh0VdpkDmPnf/bK8kra6xgJnsMBQDAOHiltMf5evNQWF7KoEkK39
bCgntz0mZF3qd55PThsI+lkNb2SLn+V575/tlEqAAjN3/pw2nO4aSotEde9nUKsw
jx34Erduts8Ecmt9tmp42mPzAJHqoY8qoAgIpYA47nPHtNh1IVBrhnDt+47m7F9b
e6vNCsZKVAVE22dmnO3lc01gts6/EolxANdW/U55WKSV/FiQ+fFbPV/iBXM9QYsr
by0eK+Ekv36x0Ysh+nsrSHTYKEXTjKe0u0K7SW3Ok131W4qKqOSjrBB5sshHRHe+
Tv5k11u8p15yU1M9XDIcJ29510J+18Ls5rvL8/bkPGy11R+bjE2flS0gqeV31fc5
uulTOHitVJOEsRc6Qqr7BUnm9A8Twdol0gwjEmSlZbzTILrbPL94lxGvXCInNCWf
vLnk22xmzZl64WXr4YOpDqLSp/wA/zQRtBjGA6H8P9Fvdw+Nz69Eh1aCutAx0SiU
1YR6r/8c/6HUUwjkn3FW5hY856fcfeGunFj2xPsf8pzruxwKBVGQ+9TuUAa5UsT4
mA6oYS3/WPpGxiwF6fzRNMVPMjkl39pi9sC+gk7Wm8VmwzhXfOuhts47RD6nozza
8DVPFzLKl6OCFL5Zw4V/siMHFnaT/fueFZtFdcuRysTnUSXa9k/A3beDhVeRIW5d
LaUXZltQ/x5L7vinY4dXvf7F90ZdGwcaXBrNfV2uW3clGPSRzcyFMj1Egg3J3EUY
1V0SdZxBtOXL1Z2InviI01mirQBmh4ylU+QQ4xvuFx9zzLMm6P4+ih6nQ95M6G6G
ii/csl/gpkxBCfqdUfzoIiIjZI76mwfeDIGAjI61C8V01xhzvcP3eggn1fbij2tZ
+cH4VZdidCjBLbsBs1XFh8XOVe5h+Vc4ZTX89Rr8T6mY8AklNQv7m15Ix+h+AH9U
kVX6bcALgrHpavBhgyqZFhuuUWAQ2kw1o6dSQgBKLz3W7IUTkHDt/1CMAdddCdqq
niOLx7qBG6AnyFFYgquYYvp+VdzACd8LmPitBa1khadc55nxWgo1fhVvPGwYEhwy
kYkgds5wDaJmL/OZxL7NcE9+1rZ0X71icrnyXQpBmkWfR0moO1M3ODoWN7ieyOQa
YMphugkW/to2YsbFR8s/QE0dBso15OcsSmPLnh2mUbW3JYzCqOKvJ0ay6vsWlW73
814qAXpj4AS9X/6x3/45LKovaUG5+o2qWM0dUQzc3AFUUXkHMhQwHPoR8Z8Ws8EC
o3guihs5ea3weDKZuGYmMOaIALFaGh9tWoSRW1zkrwvcsDHnqVluCJ2WIvoX2oy8
LcmzNu0WQTO7VsvWCVx5lHBxu+qwpulEwmqMBNDMv4rwd7gRhlT8LGFaNqU8x7Bg
NnODGVafezLltcr2Cp4N3grWrIuqZrh2d5r/9IkuZVZnRi2Bgw6PsDC+kIM6mQaH
74Aj+IGJjkYh2FfLkOb3gmxvWV/hLy7aXXAO0+XvwOfC6mkGcq8p1drlg+J/1zZ6
vdcYaNTZcV5vxYoWG86Llx0D0EdTcIaphNtYQrqMZ0Vs4qG9IsvmNow1NOJ9Tr7Q
WbMJpfmJHvRpK78+gnYIjLg8anD1SSE0E9IpvIo9ZzGLFmQC97b1LXCjhhwXlIn/
fEers88AnBHt71qV+/XbViviDzjsiJH4c2et30/I/CEsYGFMjeDGMzgBKQrqgbdL
H1NS8nKxm2wL38FODoxHBcDdoK8EXrmTARsYy6h3Q1ey7apyooFrecJgGwau/aaQ
YUrn7bb8zG+OtTT3DDPQVXzP0azJFSFfk73pSnIU+qe9HMd5aY4IvN0dXclFFIa6
GGO0X5RzEueBOxjlczDligSD/dsm3Wgf+M1Y1I833FRvUTowGFrWpDovrTJ8zfR2
hCA1fg9a+L3IocDT9r/+OPAHSbNrK8VVUitmfO+5sl9XZQVYjJrTY0Sp6TgkSQQn
H2wZAxUayd2+WJvj4UV1Nj+XiTBVdh1p5FpN72eFuooG1mIQCIZEoTwcjLoTYCf1
tMxPjxKIzzhaHovTbaQo8QpBNqm7Jn1zzGa8IHLqtnStB0CRzBuMLApOZ8AMEz3U
hRa/n3bL+v2JlbIG0vs0qQ4Uof/kSq27x1eRBkSuif49aVDpNCYypDTZRyn5TLn/
UdihlrJEnRYPyuHp6crm6lpe98zGIWGgREjGZCAgBB4HfDYhawMYuvw8ua4muH9B
u8orGoDHsgOlMYtbZN87DG8Zws1ZXhK85su/hBMNcejYH3Nv2X40Ih6WDgLLQ+iR
nL2Yam0x7qU7EEmP4YBGhWdV8T0c/kLGZ770tAYUap2AwRSW7xZXM8tfui0emam5
gfFIsqXIoZA0tYUQY25xPbFq8lAdhbGZNUmCITxdmY6plW2INIZoYb4GqdpwJ83W
X02zgKWsouJZbRXd5uEc5iZgWjFTZEGVIrRuywwgd7hne0Cqq2ukwLYRgYcAqRus
iRL267ieTnvGYQiminA5G7ULQro25gj9ioQd+RLsthXp8BXl9EUdluDuRFAgV6zQ
1Tn8DUmC0ML6f2gCQx22og+dq3OC9FmX6SbdXvhx2Y1OGNccOdoTpFglCkCXfQ80
GQlV+A/xadd/zn77KHrsdXDy2Tgf3f2xr8IBw+x1yz9USv15PenJdnAy+C9UPUnT
mw5MNotnEZexf6pQJcDL7xp7SuFxMHM4kvYih1K/1/xtHbPRQrjLfV4k6rUeM8qm
6OoWbC7ggjrtRO4eNEg4YEp5kh7Dt3sUJjlXfrBdqVvqQp7mo2S7A4YfRcpK64M6
9yrJebFdRJxbJCkgpL8xFyLKJua/mQ8Bic4JiNrNt2dVsYMzVDNDwmYaU46xJR3d
UKvOvAmxnRKUg538XglKfx5edH3XOa44o4Dv2FwL06An+599b5FG9JM3yvXZF6uT
R3T1Z49Kc1FoDqM7SHF1TdCW6wVqHmVLNVQYG6mANmAbgVYiXYxxna9BlBjbmzEc
r+2thNgKc9lH+TQ9yF3LDzS+JVLFLiEbmrSYyRA5SCsv6LnCq8sC5PW1JT8ZA99h
/ZvLH6bRandipJvqNq5vtWx2kdppcyRxEsO9Fi2TdVxCFKrePICKOz9ncYpy1bKW
o7DGM3K1mxM58WYbS35m5SfphCaOqkJOQYQLjvw2uY77HcFBLk09qvu/16vUeR2d
m2rVY4A0ghMYOXeAo8KyqHBkrDI78rGJzCSP3X+NwZXrhQwomifNulHwHVMqih16
UrS97xuVrc7JuIq8xRmktoqig6MVPxGOdawshtOqxpnJWGdEwGNREEDMF1Qsb3RR
DJTuBP/PKe9lqDTvUVZmood8aATmctTl03/YvPtg6loGTigkiiQAz6dFO6sxEQEr
qhtGoLzwc+XQahzlb6kv48BkopX6LXepeeErVYTYQ1ZyLEDQ1CbrSO0ITOOQWAZo
JadiUgw9LKbiqL3u5cwDYrCD/YF2cc/OODtPUQd6JCsgtP3fxifl5lKmlTKRdLKh
3HkdAGrDZLe2P128ESDda3uc9j6omtWt4FAb96K9hvrYYoN++JoJts6K0IkknHZm
YFLTxaFM8KZZzeAt4wxQZp+L8EhBQ1Nu7I8Eqz4Uo0QZEamTVJ3hHhKa2xWmCvda
Wmp5lE5Z2alFZsYPe9AxtmrzR0ooqZCm79zMDpHjH9SGmlRkwpJZLxDU8oEObQP8
Jv/ARlPK0rgg5Db9sO0wpwrqmJ6+NEbFueVera1VsVpZ16hU9o6rrhTibzea6R9N
5ge40sC4IpvyAE5P6s0LQoFqKSj5YPNQDH24SXGoIw/kdF17Ac/INW4uz+heM51/
b0EOW/a/RmLV9GLS/DKS6UfTXtGgntnNyE42c/WwX3d0OLOmPTg+hEVnntYTmSR5
+KMhmrODwPoEb/iB+wIlS8Ohsh+sh14cP65fwmS/mQKNDd93SJHKUZuI51Uw02KI
YrNoQFy5U3FCx8v4AQuQ9+UUhxyAvYt2K5mGvBQUopVz0Pud/V42Iv+8n2K1h+1B
6QJuqQGWtk0IbVkYafm8TeD1TJfrCJ+ry7hZwKPTpVe5U2kpQIRO/izWrLVR7Sj4
QKpbvEIdTXisOcVTqA5GHoccI9bHFrK/QiaFz12gTwFVmwfz6vvtnndMQZKF+YLn
tXt5AfelDNmXfedebf4RUpsOs3CsLHmcqD+IuI3vV57aTIpsKYPABGpUg9Rb6Ia8
d9EbTk8i4YM56zoe4VLJdY/dKSo41e6EigCnt6OLyG0h8jY7ASIqiY7M12UvndYw
YBc0+HKPrOvKy+J2Z3eW147rInpXqsajGb1mEOiXRhUQ5EaOs5GAJ7XmOB3hxAir
+dPaIWYfcarcQfoxh7NVl+Kg8VsD/tfO97wa/RwOc49tJ31J0Us6tN1+VfquFRjA
ZPQ9B9eI1s/DA6DRl100/OwnTiNpvp0khfdsmGz8SexVCDGJKgcc34vUr+eWo/Z6
xhO1x5R4Z+QvN2YpxwfLA5cFBbRJe64VraZlT8Zrpszuc4blJp1NuCfY9kq7pu89
AlQD8krY+wyY2W1+6tCu3GSibRzKEMP7KPq1WOSMZQePM8S4oIF63PSzz3Zqq5Sr
12WA5APRfiQamqpHsf1LcsmzHFYOmOc0LTx4KUXOg6rsM0Me8sq2I/jj4Z5wRxhz
afQqYg+Q5T2SO5ZpvFaAelKA9RaulNAPxxfXe7MVLdawOMb188Gf0KqtB1WWOHWE
TpcZ0ftiATc5sloOMQV2vr/lWsZmRzliEm6kvlxTRTRXzfjRRKBowkiXZQ33a63m
f48GfBkSap/JJk1OV2r2PoeDpTBMRiLLJwuWFtFlZTwQAchgs1rQXZsaZyF02upi
UE3A4YowMid7krBwIkyWN12eNgB6xWhHr9yQOvAaTY3Nw2j/Y93P8sl2E/toisTp
cVN8N/Tkjr4RLcJA1Eyb8rTcTJfExr42YobV7FdSnqsm5uilguonrQJm6m5ZIkt+
fTCkOI0xZZizZ2Q7DmxkUlJmBd054ymKGKnnpsuxtPdFVogBO+nyWasIRrbrroem
BfSjsinEy4tdNnSAe2le7ePMpMZC5cyVacyyVfq4/S9sISnReN4QEj6Y6Noll1h5
hlm2FyBYp3sJoPvHd60X80sR/NLQQ61ugdFNXbyWSMndUWFWmkLk6fnvPag1cCFr
WJdaKweGP8LBGSpuCcq3DkRrljRrTShhLYVTprpCdUNMGMCD4EseQD/wP3waeHtG
LizvfE1M4zgS89uTet9ksfXEOJt2Qku+DIF9x+DKUAM3EmEHlHNzWLL3aKrK8yyg
tqmgif+1OqOWCt6QbfPhHhkSNnO905aIwDo4vn3wnkpUs4Oc0h61gC6lCjzZGzQK
9cWOA7Zg+sui+mtLi2CcPkqBAKWxOE2/baUFuJ7vsjE1wNlu/Q0uxzNklgh4TnjU
azpjSA3gBSYMDfryqZ23hnm8mSTS4vMARo0AqxKTay8azcJlysYjyIfRbsSXS6gO
SAdY/n5MqRr9VPVXsrQl8kF8FFqS6naLeF2oOoBeifSaDqICekLKPDw4obOgJz8B
9IwsBtLXKkb20rbTDkxnvCke6kWFc93e6PViilX+nb5wPGRiotkPKVUF5C3zbL0Y
RGqS6PtTTDe9Bbo/qqBtBxRfVeeDt5ARGr1j2t6jYdgBBiOA5IslcFyBVR38llv5
ClIY3+cGGit70QnS5l+lwtyJqg8Ibq/r6BeXftWudqn/msEX1WIUE29+8YnCoWe3
4w3KQZ3xA7tBO9mgg4tBuBFgIN+aeZvgtSmK9/vikkbHz+JiySU8pkc9pO3WcNbm
RRDJJDt1TeBfwIeGyZRrPA4ubvf02lFwAHndXZeCsMLGWf3bzDE/OVKnMF79KM7f
z3dFKzXDxCO/Z48tB2O+VjoSYURydRBIYrQKU1rVp+4LTsOgDhzpWnwyxVcRTILx
xrKpJAItQMKN1EQ5YjLU/C4tio51iusuEaEHy2hGOvVbuy9GYQWqoF9VNBcy2qzq
1Fhd9CkSxfaMUjwGDrfF++qerqpaDAiWoHHwQ2/V0rpA1dn0mC33d2xsnObkhPyT
T2L6ggwTc58gGnxGYgHWZafG4uBj+7nSMIro5pTSErvDCzRaWXrzSZN2z7pGAKXQ
54fWHMFCdSIMxIQGMEDyomjRyjS+7fT5f1QcWyiIfSK2sUWr7xWABPsF0qIkgU6+
lVcOI0rCHNg0DRUhb6HQjs+8JPeVKds/mqDC0fsReMqr3qwjsbG6IiDqctuRML9I
9yiiyC4SdebfHWKT4jBmvzm3rUYmZ6aTAdWJZ7PknyQpY+2JMQlDbRuEEGlogekf
7o7jBHx2PLjC8NmZN6fOeiSUakryE9dhYogV3BmcpSvSsBvi9bjTlUtm6QMZD9Dj
w7y3rLsYMzZKwsnDdR+81V4JNzp/aEmyP/n97vxoe8HCQymHJJdghMSedNyjLCgx
tgIqzF61fZYg6I/O35c20Jm04RkHcXkARUToIWzTvMvXNFl7KzqS7c3jJazDUp7o
nCHpLvN9RD18YFgi5FoyZ3/FLlwRWMsMn9LhxCm+kT737e6nzl0JUULREMq6YUcI
c5tVKeTp6cI4Lq6WvuecmxGbcW8rDfmftAymOSCo11HR5KTYTNIRTFJjrHRv1dgH
sDrZzTaWLCHUkU9b1I4PIWw5uRDwzHJIktt1tGU6RDAX4RpJqB46EAsw2NGZQLfA
PpJdUqLPHQbZ/mVb5EZKLmn2nO1WS3aCWbHBkFU+XtcKw7JiGsYCSk+dO+pgLVnk
mMiWXWTXwDtGgIhn4IKQKz5a7DGJSwC1/fR2/EHIZJ3bFvGGTWP+Wab9jH5g694h
8P0UK8+Fwy3mXra3fGso3FdtaLVMiSyrHjHnhphAt0lzYrgTg7g5ovWDYGuoXaHU
eQorw6uUvEUE0MoeH676dm59qQJ1cFMSPJIfLA6a+6oW8r0l1dd6bOtb9SM2ysbj
NC1l1CBWPUbon3Em9KR7aSzAY16JFQfJLBU6VqMm2yMN+yg4nX7G/JcNU3sMhULY
KVxJiTfdzZl4lB7Md7R0gi+7V4k6cvmQh3t3lVDQR8PVcIv11ojGJVlpojboZi/6
kb5J33+DE71s3PjXQSt8UTx4TOnKRK+Riur4eXhQ9uKJFbBKv3eDYLFWZWeOa4u2
jKhGIc0XAn2qgiELQT4rxRHfNboqnKv6B2pI2VuBWjul088phW2hKM8RYS8MwpzT
83DDiDG9QFL0bl0lhjkSenHkKyQ4LHeFiBDO+FOMAdT06z/94jw/q4gPc/EVYAxT
/8cvgkTDMrRBuJYyeCCcE01XY33909fEVy2MTSQdMJtb8CORSFYjzQEjbKWD5qX1
zlgvrcQ9HZhZpcv7HPdHpQltZlS61lULqgl8EXkXQH6IyY4aM+4KLXHOsOeR2rKJ
pVkVVDFsGHQCM/Rum3w1/Z6qkYN2MGkdXsuZ2FN4kAInj0/sKMYG2W6xzoU9VsL4
yABug1dVC7i5/rshhOIPPCTGsRQOADxWxd8gOt78oEkXH/HB0cKZy/fld3RCBpT7
esu65OmYVrkjYzVYkw7cZmIvAw8/luqZeo18XDjpikqFLhrOCiJhtySsiNkMFWft
/rCIHqyvwWf3AoZYME0beAi7kg0UF8JyOdfRhWBAoJERmsqNEpxxDHI66sHHr61e
oZukda43Bu9EHQVZaXRG12rBuvCcEX4QtQVaXI3MhLq0XkyZDG0BX9vp8iFN82nP
ZDP965mN9IGUkr1e8FHWV3xJ9Zz1uCgRLs5G7pGNhFKbZUI/PsywX8sjstDbZVjd
rNco37K6dd+uddYTj9BrLQj30qAeJJtATwOv91vfDk01E8irJr/3+omAXpDKGYDn
RMmHqn/Uk7ZNohQc1DcEfPfgiM8hfUUInz7BTTVHY//17+KvFqpBe1ukrVhK6ec/
Zyzy+SibQvGhwHrcvCmfGTMJCBzX6rMGZJTKb2P+Rww9WKfQ9JgnXf/JhoEYoKcZ
pibWF5klW9aVomPYWooX4AMEnhsDSIkxgdKL3LIbrqieFiJ5qnEgamuPdB1/VHTU
fnuCvJIUHRMIhxDUBBhQTBq6FGrdbUq4PUnymN1Ju4yd+qETAoUYRE89KrRv6iAT
FbGi6nUhAd30mDaE8Oc/jG+i1q2aUsE0O9UJcxVhzVoqKJbqQNfZsxHuliGwG7Nl
Vp8yt1VZebAtcUQYoyL9qkxaJNf820BjvgN2X60+XKj7exnAhzk7PRKbSP+Jkz+g
TEy0y6xCfI28lsEyDpW5/adYXWklHWO1L5dKzFnSl+MAtN1c2nEv6E4PR8Yuv+Y3
V/Bx+w3xBWXl3+PEsKCNLot0o1qhcc4HAxqWX+yaKnYSgCz9fcJxo8VFDsXwtoAj
op01P0tysXOf0UFsFG5Lb1rIp2ZrjjpqeB0uw3dGAo/7dSjfNGoFuxTHCXnrDjzA
95TBcwFClsGKlFkU/be24L8JyqB3WKk43HcoRAL8J1CZuWhu95diUN8Qsk1iBp+a
31gF1EKgN+1hTWeLlJyAMHmkFC5134Aw3YLlntuGjb9gJkIskqeZmzcLvVXUs4rv
25ZEsuUFO/dwesdUb9MdhHW7wsf9KLQTlU3L/vN5W0sojOA1LPK7XX6V1Y61GoXF
IH/6pFk0pym1YbwXZUcvxLH9cT42hKMZzpqvaEa9ehgfWtVv9ydVX9h1/P0IJ8gy
kqOF7mtAN/ewPNJgc9UyPTvPiyaGUtRcptYEFH+n4OctZ2AJK1ISgmscZwMa7qwd
Zq2gmYCdekWToL02MV+MISRXcZmBc0gNaJavdZ6LUF8g1z5BEeprclENxRVC3Dkl
u+eP0D/WFdSlKoLFHbMVg7croMY2UyMUnIitf31q+/x3h3mtAUzCaWRBNUB0oMr+
c+mR+d/Zom0V7LqXuPmeiNxZzLDSN7uAVHbdu0EMiUZorAJ9nvxCK1LawcCqhyR5
cyCY59Z8OReIt0OUc9nPn4D6qgrrhAEMJHY4NgF+jaL90fOAfujkP4jBO8NDvUOy
YpOfD0UCSjKJZwdsdtxRW6zP3mgtkNl2Sye5z//OYxtcxc+CK4vnMhw9XKrmPHfA
qqFNLHGRVY+hErTegnoI93DZT6bVHLYdgtmxU2mPVXnyxwMu7mr4IyF8ayKvqmw6
7nd9mDZJPAPKu5e3QDW9Yyow4FjTijB7NedyYkrVsPXLCAc7dE/954U6cosxND7g
WlTpSyuoXS2sNU3Z7qo7arueAv/i1IfUxQAut7oap/lw7x9vQc34/7vh3Zg4EGQq
PLzbpLwW+BH+qnn0gSSeqnrBa7iC533SQG0yOhZF9AmBKChpUUfeWnsK5ACTf7Qu
/Uopu5zRKoEznidVYjdmcWi4EF14ZS0tWL0MwCn1rxQkvYs3WHfVXJldrkVumdgi
OyUi8LKOBSV+9RKk7SaYoqU9u4VnSM1Fiy8TEuZDXUFQZYE21fhLRO+bo1YuxByc
pV0Od3Xq8ElMpObfg3sFxaWdNtMjSRSPOlX33BLdZ2PY8sOBcyPUKlXj4eNIQ1vp
m5NW9M9fq5FfZwE1AG7mDZxfasTcv6Nkx4z+RV06SZ0ThsYAiJ9sxUr903TUijIg
f+zs6YF5O3hVToBavoMz4mtKRsSSIkNCcaXIxuFrrQzGhbO9VaPrKW1I5KxODruq
turvgJtMyV92t+z+D8WJWCUBC/G5HfU5ZhNqi7afR/zEIBf86cHWZ6GqldVLKlVo
sUJBi8/4b7N0yA8neXgAD/xzbO0JwpoA6XJ//SiydNSseR+1Pc7DJJ58lzxvmmaC
Ee35YQVJAvH0puKcKX3fHuwWevAyoWJreA1EiZi7Bdyf5464lFOZ2OuKqe6HaYVf
tlQxgPKqZ+7mgRpHZ10nxwJ0xrfgh7IKDUiDQiqBQ6LiSsgip51hawdwCxSDnWsn
Wbh9bqjjUVKkCBtL+fgADq7e49zz7FYQcIS9S7/ZIKVKxNBqtE3mpyPtAStJzA3T
ZJCPij0Iz5CiWgyFrD1JcOwhuSOxW9y0KYICtQ4ck7wgSPWZi9sVQiHw3YgVN3FA
EJF6cPRJLuPRSROrCKyYel5duqSZn7ry5wJZP3rvakXFJ/HyF38NYFBAKaaQr1yi
RR+uGm+SHJScWH5vcWZZVve68pbrHqcK6LRGZ6SQQvvPGpb+60eNnG7xZVw3qBk4
9xHEgL3LOlBkSlkECzbVMuYwIrUWUriJBPE3RFerLNXV5I2uyQgA9bI8pgOguCnb
SOuFJ+KjD3ExL1ShyKdTOEHuYc7rKUXAs7zrfoue2NB6eDAm+L/x2QouA+R2DTw7
Ju5+xc/x6jdls3KGIjd3VDWgqAi3yhHS34nIDNGzPqrsuO3oaopXFvJ6/FrGEHJX
uqzgfXtb+ZaGtU8aopULuS5fOwwUPHkYi9+4AL2952RZCNmMuntLn7DYUsHLziQO
r91ufCTy4Nsf0zP1OCGXp0zzn3qP3+i283JPVEb/+nK+/kDDdmjrBN8VGzgKwsSg
D0nT09696HMGYky5MvPcvGL1Zk7Z8tpFYeWAON3+FfiOosHkcMj5PQkgrX2b3zAb
Tdq6y+nITulFj/FQOj6/EZ3/6HCXlJNSqpY3adAkWm1sMT0lWJaaH4R94mJnEw3N
kPRDhvSCf2PG/QN3voYqnuZV5rEgP/3a8CXAEXFROH52XOKdBAMrJWi4tsGR59xk
XBa6c8FhgZyYp5BJzptJ7p0D3AN0Dv+UuNKJMg8KLchTZbVvQxsNn0WjrIGpQhJZ
KaKfv4zTlLyQUP1x9myQj5ZZusYeAj9MRiMyb/3ORys8/wDLkMQCopC7gOPWt40n
v9V8LKaSUJzF/qZSwi/qYqtFgNNvM1ThxNEybSKMSZAxcwNNipp6nEQhyv6ZsupD
waCF5iu2YADMc/6vxPf61RQhhzzZ07sggF+8wwETZgsg36nKPEq+C14yorv8lPqa
wAog1ahQYvI28R7Je+DTETGHhijFXMpBqoIR849J5fa646HmnD39CC3BW4vULAUV
27fHsB54RSBcE0ZOpEZzcN7LI+SHvogm78XNPGKouDR3ywbYI6ucnbgwWUyVDB9b
CA6yXG35NpxR/Q4VXhv4xUvLUdBkgHmJKJJiwBGB2QJ6RzVIl7z4qEzJA9TAqYNz
oM25XMtr6ciHnb1yc8P+Vvy4Zgr+4RNjYaxNZiRBlNEKhZc4o+nyYPtQKNq332I0
jvGP+tRUyyIm0yjFNbqNeCDWYfoIjfH39RxqF/GqZTz/l7d/h3RPnIj01OQCJMY4
gt95TqRyqRvTyTnB/Mi7ZKEmWQ/PgQqfvaGm7CI7aeWwJIBCRNwfizOsFPL2jVsG
MkOprnwqb1u+x9Gkgt7Z8XDODsy0SYMCx9ppar9WiJApKAigGNqHAGf4f1obI5pr
28Oalj6qTJmdwGT4LBHM/fI9upspULYlD9c0LM5EY6g3tBeV88XZnAe7hqQvdEEU
2ASyAGBA6y34s0xwM2vXCyP37ikNjxgeQFyOhWnejM+ub5cIIkVAIiuzDUllicIv
41J1EyD8i6Cx3LTPO9y4oWMJC2dOL717OlJZo15U6tCj1MZcF02mfqV80AWjDM64
0olyaSfsV3i9o/rqlAy2AHJ0ivQJ5tOdakjpvOutX7nezXTBkWeef7KGRxI/KJdZ
m/4kJKAZz2TR7+1ulSqQqHi8tA0/c0FFb6p0HZnlagGaIncZVHfev4ifQKzKM66A
+rvl0mPaNDr2dS0hhJVAstUsqusrodQ7HTnxKfNF0ayBtBlN69mcVzn46bB97EjP
j9QmoSKcSg0Wdxn14xqbOPg+S4jiQxw1eTBS9EvGNdstbHONb9C5OJ4R8rPFHOc/
J1fb94d7BdmTOiRDnbiI8JuJfqW+BMtenPYU6J/OoY8xCQ/ZH52JB+HTvDRkCqsm
dSQx/oMmaBhEXpUr4dGTh0wQ1AGuSyEUXl4dfnM8zkRqAZJtK7lTDtg5fKjILIwy
ZlHOEoVwc6rN5gRFZnwcWIAlguQej0CgAjPcM+Tg24vV48nfhCjbUUNcbsB4xOvX
lyFlxOpgW7EcD9pOK4FLicesW9dzSzWrH5AORXytzvSYQCbgE1EUVenOvUeW8X1z
5By7W6Pj8xaabIdtr2EVYHi4fPupDnJX/pQyOxk7fmC2KgrbqUkIRZdD+ak4iCb6
ANLEAtxWX0+hiEZDwtBeX7yBoatvZzWJUEpJZChYC4puMfQQmmfEu9kiZiwP+CZD
LGVy81W5lorwS+z28D1LEL9XXetRsmfrMI89WPVn6jtZv9lh4wrfwWmPpbTeHzTZ
AXvliMqPQTDHal6/Ho0ozWUUqXvZJJqHKqv9vTdlZ+Y0SyVu9RX/xQTguCFNpJRB
zQPxIuY3/4OJbfuRplllVVmiSFFcCjYlLoA5CYpHasPu8qzK/CmtvrIsJEMJJ6TE
7WfctEtcUz+UmPj7dDL7V90MDzWQ0+xHu/MzvZiEXwSS7wCn1FeV2j8Twtq5ZpIp
NzKh7z3M86CY7n99B2+jx5i0aA1WvYZU+Epqz8b+CwmMphqJ7zw+wNKfVVp/ZWPH
UQnMTf0MRy+aVLIeipSJoYhNLAt+fqk4cItNm2tGeUjjzNafR2OIRqSGkbr7RXlJ
539xhJCoToveu6TiZtDfCKr4QCpaBzDcsTD7s3EG7XIf7AZKIGgtZD7klFtK1r4f
Fnx/F2/H1YTGQ0+B3QWVFoYwRDN2Z77T8oTByojh2L7WY6sIVRunLWodN+YOro51
GEs+MsWfJR2o0Zy8hjlNZNBNX0N+DRYot5QdBcryp3uUu+elx4NR1h3qZQS2r4Ja
apbs+5hBkJjDN1DelPFJuBOlwc9S/zaLuGHjGajsCiZ/PpY0hbpmyOXhdrO9d+py
oXeGyYwyQY1MPlOmb/rrV/Zmfchv7wx47kk/z2O4KKNymEEIk0GJ5pmEDZjaEOH+
P1feQg0zYuEYsTNVIcuStpHfMVna+0SqkOy52gDn58jgypRwwmBU4zRby5JdOqQC
xO9KABii89vbjhhgjbMQ0NH8NiIYZ6eo0A56xssVt+K/szzu0oAUWXRCWUmyy+/B
Q2MbcuT02aw9NXKlTUwqP9d1X+jOzYD5Th20fi24bP9nmSETv7lRwzdoyRnwu2L3
EeKwoFEWXQTlXurCthK9rVkgJaG/BFpAlv+sc4RHy0TlbXXk6SA7DSUU4NSciUiS
Cbr/ciDVEE3MgnxuKYj5K8Ke6R4+MyHopFbAX7vo9OSuXLwZvmAIKx8yI4+h4ly2
pJ1jptlfAeCYqeJI2OstHSKFifFR9fA8e+K4GCP/wV43r5dyo3K3VAW6u1RCSRTG
+2Qp3gho4t+HdbgABx1bqONYuHLCEOTZPJ4LdnJ8bQW+zCtu0pnuRd+8BqxzjmPj
BYbdf4g0q7Q/Ag35g6RQw6KeWTnIQ7+yFPRl5S/ITvTllnAYt6q8EK1iGG35jzr7
v/YEciPwdjiFBsmkyxNLApkDeDXqxxF3LwqXNVYx8u5Z09mjGhvPBKNiqeTrRSYw
Dj1SIwNA6HypmCCI2baFnLUJkGvLWIlT++YL9h2mGW+LMtm5DW4To6oiitRTNR+g
LZpoJWA3F4qQ+pV7l4mCvNkRaxWCb3eJ2JRrNMboJrMN/+oixvtW6upFdVwfz3Ol
zwMYkBeDJBXQuCyYEi3gIJ2udcJc5W56IqOcPc7oTfeaZbqnCNhY09D7n9w7fWcG
415Zc3YnddroMmwWb76niPxMcFao5yTLMR4xefYjiLMS83ZrMXEGZ9jJIyzD+uFy
U71sJNK956RV3IQ104TcSq7K2b1BpFQOPwjfdhpG6Q+GkwYKHbM1Uzspthmec1i3
ChmcN2toL78TitACWJ8reNy55P74f1zeIb3WMKtD4iWDC+hn9Aj1gGAr1u1VoDcC
OR3pWYJ1YHlAFQ90UuZ8kSGzKg20OJfJ8Tv0jjcXsXPbpHpOW8JRdwU1ELsdHqBQ
5BEzokvSEDlijy7rASxU8uUjmGVq2h++gm+AlBmC1mtdAtYeCjVpV5VGWEssN5oQ
nPUj6O3CJNiMVS7UPB0paICr3+GF2RTkUTy2fRfuG5zZeBEfN+80BbksK9M1zpZc
aQF/+Uw5v+uZKe5pEYusB8IEjAs5dk734HZFmVerOD6JXTxhEh3OAu4ogaWq3Ouv
IPAhCrcfeA47/v8pNFDmP0YDxHKnWnHxw/nwHcCqaix7d4u7FJPkk4JgttZCRQuE
+wSG9f44bnxNhew9nFZCg1L6RTQNCOR28dk5H8kD7Fwi2gHs8OACJQxTrAHuQDUd
RFhZyKslMeU1qSBAMmwUZoWy0hYVT3tl0oSodhiy5MUaTkzEi1cL8JoNevSEO2tV
1QAQj70VBZs3HI/EK3yRBeaFeZEY+9HSzwirEAdhmwF2hQ/hTXlZYnDuAxrRBRPv
JRCAm8GI5p4ZokLyVkGneWPonL7AdF2+ruVlpeJkp/apOCnf8r5LBm8bN7+Ip7UY
ZTRnFW2zLOlKawne115tsTEkdWjPKY0a2qaExEbxDHRtG70oTaAF48hBqSITy5Q7
/k+0WBHshpDRkzLsrvGxKScHzvoHC7A9uynkunLCfPyJxjiQcumGxYXE3ng7n5gd
LdONuYBciGwz2hvXFCaws2N4dXcA48NZv9ggOm036g5URNHqEckit00qUbsH/ozD
Twd/W5U1oxDQhOqOdoVmlbj8lRo0sp2kIKun7pZ6qpDqwsZiKka0nAqkJ5qcLwRu
uYMi8RGCYMSvfafJIanXG2Jr/ZsE3HW9/t5xm8ci64VpI8F6T6/5cHpKwQ/Hv/1s
oUpiDu32f9IchB0GlDbmfBDpmOAfI1M/XvvJD4nyPnMZs2RyImTF0K92m1nufZAU
xvipzjmS0mm3QQfDEctPti28ckwdpRu9pJxDe8iil9ngnnd4IQVlQ7id54we5yDX
NyE6Za7BMrHpbvtX5VB7kwexHReVxgQyegYD8/fK+qS4uElXgag6DPqNWFlcZsW4
N4KkrxmFbiLb3KjsxuG3oH++D8biZ0DKoFB4zPrM/NCfnz++ajWkVN4GO+CKZ2Sb
3cvmxgN2g0SfgkEjXKn+wroZ/eH3w86DaIXP+yI3QYUGp8VlW1mQtKtpDqtu5vgA
gF7nTM4QSnZjifXBa7t2ap0DSRiGs4lGwfKgRZ/9y5xU2ZMytkaRhFQd+UwI7Tee
nqSrR9280iQOvOYc4DrURYDUTumYQJJey+c/l7kkn5cMMvkOMi+NfrL4d8BGyltq
m754N7H/NGTMq8venxJ4RqDTjF+TKY5iOzuR4T8Vx6Vsogy8ChtTkA3a+qx/6XPe
Mevl2j4B45WIy7Pk1k7YctQopWMbKBUDERHae9nyk1Ze0pMRLjM/GMbtqwaXwKiH
FXOfrmiTE2adLP3epWwHFxWV7oMrcMmmX8EQT437QDJ2ZxoLekQf59b6xIQGcrSH
vBdzsoYCqWM0g1izgSkkzmcg6ngGT0W0q4WjJHXJ2yD6uBQyzxR+XZF9QVMKwTdP
ysOPeLRVgOtocz2NGcX1WhCj/o00q8MRPyFNa7pLZLCgEDMwf3GGxyn8domeB3sN
h4hIZhWut5qZ6A9nQn9O131h4quF4OOm6qn7KP6M7oRVSrY4E/a8hvYaub7zdojJ
52VpP7lWsITcj5WZsC1sf3cNLRN+YkaNb3Q/tEEM/u+LanEpiEl3z+hLyCZ3CXL9
XeEeVdVFBlg/r9gmiR6kG27054Z9njDGIQKsrUq3MJEM8fReg0BE8v6tkz1fI/Ux
9PNkcJaE5rIIMUt1O7D2vCooug8GlEk7QYG7Yf4zVIf1hNm/DTr+gy1wLEaRf+Oi
OUen4yj7vtGbNMj8QKvnk2/Edo/RZ5paS5bfax76hxxxR8Z+qCbWUx1zUBX3PUHf
n+XpMjK6D/7bCyeMv6AA7LhPILguF8Vxa0l/N8s1MSzKN7hVfnw2CqpIW/siYoXw
vCIHgm0yMRKod356p+pEbHZY0CfMlw8WqIrW6b9o6Ey4CtcC+n5UxkcA05n2i+bf
7reGaS5rmW5r7F67f6NdhTN7yIGLOagWDsDipGxUn/w6c/M/Slvoa0vmvH8umv+p
aDUS/hxKhlkTHlehEa4lxFIlLqPz1nguSFLbZriCVUk4/upqfNXkyZCO2+3zUpfS
3UZD0i5SIMjFvKlXcNw/nwFLerWfULp+7QIijoAHNqDt1GCy7tJb4OKgZ2DBCPTA
3mRUYm/1IVichjbo/evHPp0XqKSPC3nda+4X0htjjPHvd4024D/lRTXQ2J4ZtP2t
+Xu6m9ZEYd2qXW13U8gYaanbhPNqzYN4RQlsMDavRrG5jVJbYt2EGTLey5BXPWBI
ccaOLrCukSQjEkaX3CGLnYBaY1SbXL0G+l9L2ECDbMqmvllR9pqN/h230XMNcAMG
PyAlc6pWQ4j9e2ZLPAl1k/kjN9GMhixKxyYslj8rU2NfHHoy5HHEdAtpm+Mm2W9H
J4xOd6wQozYhKbYEsQDq+tO0XFJX1okzuw/gdNNwpMjbC6T7WoiFQhqGyKUf5jdY
dfyydaF7LM0IYznKec3ELxCPil1OER/vnmWBGXL/h4U6aH5M7lWsqBV4+oU7ZGoU
Sh/yyyjI4e7XZVPQA7xIe38vvWwTGyURT7Ocf0mmf99NQIs8sv2Em559u8JWx+s+
fOdB5hND0f5dSqW/Zv4sFDnxRAAa9jC9QPkHlA9uTtH9k9D0vXutUl5jDM5uVuRy
OtYaxrX6Yo3GKndYQreGkonYopzo061XKtMlp+FDqvJnKAhKIZoiVXBgLfFp4HWT
j+qCMAvZGQzQg4Z3qTsIj+LapKA+Ds9HXDlGSkrYwbjF81+1jHw0NIBp1Ijzzfzh
nIKo2rl+tzndBiBJG8U4UEjD9sHzUMyCKTuSapYlEldUvBR3ukdE9zV8kS7Aczmq
f625tuXBoHlyFiijEN/OMMXmvl6Aq7U9vmcKCrmGwCRHUJ8e604nvYPLhec2rLnX
Mfc4hMOxydEq1eHXy80mTorlGg54463Wn4BdlHjSFKADSF+9uhkubG3QoooqaRCr
2D9+UUesPLI9PV0/3EA4W0GIwH4SUT12KF0MD+6RkBTeh/FIx4aEbDmJJMNadbTP
HtGn9BuT/OwzCFBmMq0ewEToWlr6ZVpGNRiyHDnp4DijYZ0bZErzfjAnMl18EFB3
H5R9fxTO300Utt3OxSrLSUEn9QsvRh+J2qG5bodFENeWckNtcYzGEAnsdXN59PJ3
Ej+B4J+HiaF3YPmmzEm7wJm2TVc3pe0kze0ajL6IIeS/hHMpbXRbnNYXoqHSekKI
i6DMGw5zNUf/xao5eB3LZh1I4p/bcs70fjszyrus9ld3iXw3a1f2QB3cGwL0HiyV
isNJPGUO9RzAzZGTzBN/Y4O2njLXljCJBMn7OiQn5X8VCJgRMmQL2mzsY0fYiTOv
Ux4H6oHKv5X6cAhPULsZY6kr5fEhWhANhfZs1E0sgXl8QJHDLdd2rAdhcKOOPfO4
c0qoBjsl4oGKSRLivqGD4YkEGc3m9REB90cFgITrZ7J1AEi+9W9BW724hTFbmb54
jNqk/s/E3ODF9bewmZe50JhPSZGSKRmobePPZ7sPKcUPEaH0ftOMSOoVYe8CSw3B
18Cquhtv8jYwa9A2mWlOl7YNwBjBT0dA1MvEBBfF8nVLVfFyuxEHwrgHcm6Jv6rf
nCBKblBqGvtyV88/exH3SenDD9WyzIk43C0BDIMA+ZfwWOc63dueus351Cna+6Ox
8Jwwv3krQZP6OKjSBPfCRDwkgrCS4qafgCh0pnJuc9ntoP19AkSVnfmogsZWvNyr
/GFNLGImdVwnhSPV9VblxSK2p9BXwvU58f8s9JebDspIhJ338yZbg3LDES9AdL/Z
vEHEob+QdgDmczKtbo/DsfDRAe4daxP/UySkH/NVUvc+mwHEOdIPTcDYbu6x8dqb
2QldV9jSnEqgDjdiiDXMxB5cbyhBzkVnGk23BUHWQkoSVeaEMJ5q9C/L2q0hd6mr
y4ni9vmXO/AdjSHEkn5uLZUoxjH0Sp+ixvUh+CR0MPasHlAKheJn8XdvgdewEPmB
FSstPB4s6X5FEARAV2JkIEc7b64y0kuhypr3f6SLWId2eb0JEKSX2s74B57DG9c0
c5IDWCDNskZfXcL6g+Rcp4D8H+7u/IK3nlCydPhnNXGtTxHWZ2f0XpjuEHI5tuQ3
6NI5IAmIaHAQW6Wuwpvi/1uYovWKrPaM1Nj15WS2KD3nU6Be9ldMVvAWsOUFgqlO
gAL9VN/D1NznIwhju0Btl4RlzGDC9+eCzKScXTxSiffCOchfMerMzh9nKpuUBw4Q
l+fC6jKJJHJD7K0R9Yd81tYDwrFY6llaaGpNxygl4OzHERnTPVp8q9MvKB7pI7TR
NguN6qH6HYzZKZubvl49VMr7iMU2Z5uLsKUXkyx7pGOSQINJsiDSVB2h5Qh4f5lp
8pFMAC1CoolXFUz2SrmH9ZxgZJb8pMpKBI6o84D66JsfiO1S3JF5BGdY2z2KMcPr
J6ldtAjv12Tgp2u7CWeUIabb1m1PwHktP7q6mKWVK6xbMleZdOkZcWZyxkF/z+v5
H/m1FNDWjk0XjwZiPbYCXvHQf1l1uD8eP5HFw7Ux5edKDWtliO/q0lFTXox0OJoz
XMTLnGNe1rIc/ZwADMQvE++RM2jREJHxOPi5qmoUTlw/eF7I61MKSApBP/EUuq/u
Mu5czxid5nwIfFYaV5XuYXNUnidqBhutFtCppn3BY9ENcC/L+72nxtg61o1jIDku
/U64KO1sVjnv6sRhaUuIH3iCCRq6W5Rdt59nka9wq5rVZ8EHFpMltIjzEF6rFqpr
I9pnQ7agSHtFuFRnQys2eRlXYGY0inc1/APJpTMUwroyFu8Heg2Sx2MM8qsaF6Cw
/7BekUCvBQOvFI5B2WSYgQy16x6Ebv+shLN60TMVAe8J+RaZzjNarkgTDIflafpR
PTmTxgPxqIpk1lAEJpL7FcnBJ8Dnw4fKq5AyaO8IfHYpS5wWKT4GRJi1x3w+35Jz
BFIRnBwWi2PRAzKxvHj6Y7PMmW8Je8pCsflLI8W4AXasUAfjoTHd7afphyulDEHX
RSo2C4sBV14sJ30/42pbifMcOwum13+OVqo3G6l5lgdr0MVaddr15fNLN4LhuDwC
OojqBSZ9bXfIySv0q2CxC7anaaJwwBYzszkzOa0OaOUoXApHrmbUOJlntujbEkDM
i/hTGBGBwOwuKiKoL8BdGC/OE2RTcGJAb4RA52UsAY850nUMuZyjSVnJBblnV3Uf
jqGGmgPeOYYjtslXio2wg3TCLtVVSyFYT1G9EyW6h2aOjEyLu7ZKt3uE5jRVDW54
lUcPLZlyf+rT2CahRfm5T76H+MoEB/4bhugGWZ7LgzW7RK5uCLsJksSoRDeadK2J
8HMwocQsMg0yOwMwP7Q7UEg4EPsDmbXf+mdK2huuxDguSPw7iV1WVvhGhmDd1zF/
LR4rhGnN5W4UTwUjdwjbMc3E027mpOd3CRD556RrEjYKkUBXPd3AvXN5V2zrLOiK
2ab7SDoX4rhPSaZxHIfRHLt2G7rK5lygvduOz2shyIbxy5q3DH1ixe5wy/KwlHw6
OSvXo35AGwFGMy6d/h9gfow39kU0/GR1GW5eeQNYE1LKNnmkEBFge0VrNvP+T9Oo
qPTGpa32bU4bowaV8sMV66/u+AGRZbA86v1UVzNavNCG2hDnfCwNED45809goyVa
G684ZXHMYRoYVtbNh10EgK4G4aQVRARkMjz70oZPBmeirE2FgLgOqvuHnHdIazeU
UMQ30IZZ2UCL1wcOsqxjqbe6FLGhkItQrKKiiKYpHrpTYhkHYpjkS7ARd8CRi+i8
0UqX6NiNKVkYdwUfALQ2Ygd4hWkIxRwrIHD8kDLYyYpTtLRjWw8yr2MqHJFC+xjs
QA0me68P1NC55M+O8E1PkJUBdpN056FA1bgS4Ci031LXW3CDCBSgEsJRfysegXyg
j7asYzyRjLfB3Rah0b8XsybtwI8N+/P7ZRxtiK3sFbXSs6/usLHfeG0vqaBVhSwQ
wZw4b+dBbtrjtIZDqeU5jpwGBR74tI5riWRCZI2SQsQzdrwumAaSHC21RO9LCb8Y
o9b8+ysfMTo5npEFKnhd50oItuvHe4XSIrtTi+687261BiEmlcGFI1rZqaiZZywf
a6LS3aA5KEIpY5XSDPV85T1JKvMWAG1ULCmKZcvtGRdGNLaDoTXtlZOQghPIrMXm
fNzDdiUdkSYgDRcS7y/n7c+P/CxgUR/I+VfD+Rz0lX949mG565CnqmlQMDqAMLzu
f6JbkGNSTXdXeyKoluzROQTdFRK62RQiNi6kHeXY9zgGvo8b0ziyFjr73aHuKmhn
Iojxf6LLSXptFTMU+SyERuP5XvFMR/A4XdTnSwLhTcKHLnDCDt6TesGPcyN5YBky
0ljrGWsTgyMEL/fmdp9mBY/tJ/oqMFOq7Ab7FsjAlfLPVo3DYuF2qhS9Fo09BtZL
KW8EHx9W9NogVrS+fAnx4Lxbxh00MuuhxPc4gJD66EXGClYjF41J+Mf1nyTNRoST
BRF2xKDChHkgyRVMP2iItFm48RnYk+CSyO95ol4NWFvujEDVE9v/ffJBp+YnVRuz
ywTyFX8Ap2Jl79jILqFsoDQcW/5nVreIJFx7PCDvxutqp/+ZfHnoW3s5XsgGFPYo
bdpxDQOjJ4BlsyYYrLmtBhbTy7xm6QW6KCEwQ5C89/I3rqAh5Nz43JFc/57ye2gR
2dbWfr5KFee3Vx6GpHDTOHZZNLegnrLaWUbQ/Kln2aie5B+l9ZZ1OzFeMfWWC3wl
MZwTfgTZR+5n4nEsEo1ViDDxVC3l24h72QHIlSeYYnKfCrK9ZySPrJRtoFzzuKhQ
FJYOO29I9XoTg0rvcK1titJYQysxvi75zstlSxd8jzr/x5RqBUyre+ZYBmfESrzb
n4L4juRlw1oHiwGkv3OXv5JJKrAyUU99vRm4vibl5o+NG7xrLFf5riqLfiPcnsgC
rX8gcvPgIw6SbvgQVDWgdHyRPVXEbeFQZfXlnrCw5yr1LFXujhBw6i7gD2aPlYod
ZLC9BZix6XIldesYrHmoX3HpEQVyvmoUtZXhNWZF1IlcAZMZCpNO6oczimBTpvOU
l+VgGSrRg+tP4Z1g6UMe7A3vKQapPoc7mEvuHQ+ZZw/1k7G1Enw+9N/Zv2tehqwL
2vZ+bDbRDywI8btRBgJbXtZyQwKpuwPPU3EmZGp8rvpLwbiW6uLhvoTMqz4YX4x6
2oiXk6ROzh4XXAyJG6F7gLaoft3NKr/uikH6sQ+z9i4MOATQAuhjKXYAw221ataM
2J8m3UNZlTO1gvCkcW1xzFWBoxM317ol43SUR6siuj2o+m/7eINLtF3ilI6/VJz+
SO6ZJ+FbkSIH54Frji+Jzu4wY8WvozHKjCzsdjDDqgrfJAIFOVdjhQ+2V+9mWyoL
2INmgdVF0oQJno7WlUwH50P3sF+zssbpHkl64Sh+5YDb6EdSV3AXo1IuwGMXrNCT
Z0LyZK4FZ+lhKlFEGjT+S2IUMtZIatr/KQS99Q0cxwE1oBwvUw/UIYDBmSGWURSe
ZcDzfZG4VR+uggJp6AL4KoPB2O8qWz8jN9GQe93e0l7jbv2ksXURBnpPJWg5HGuC
Qoika+DfIYOR6KgoE5KobSgmyB5uxuPKZ1DPoiQZI8k2P4loWQkmpaNoHsqjahHl
B/wruczW6Dg0zXopowJaMAb+DQcTtcxmbvN9b/Wa3f9kjJiw2oHMze2O2EQ53i88
g0AAMwN1UnBgYV0X5MdEyN55Qx8egB6pPk6nNdwdR2uKtrSizZ1qTdK7o++HTs4D
Mk1WC0+KEsDvFJ1eocKW7ktk4VX7jSoKgZSBUuWTNyzL8yaravOJ8otH3Z0zkJWO
JjSnzlPmSa2iJ99G15eNc9PLa995K1Mg41KsGTWcJOX+wUq/ys0p0I9QJlloChah
g1Gui3yelv0Odvf6k8T5Li+Fge1wAns8ZuD4/jq3Cco6xv25wVD+GjLlIRkjGry9
Brsmw+8fhQPIJBqyUHvBjYUfbTsc6Y1k1yEPngMr4yshLE2WXRHqL7/Ja3yI8/G/
zVWAXGNp8qqINXa51IXXa/RzFSwNuHlvLW3FAPtReUZ2JHv8j06ByzmZdzKRFoD8
+G8nKBjwFQROzhyVI/Q1Z0faDkezSQphgXWlLQV9PwRYr/oDlvzAr4uNW0x4VxD4
YEJHzaMa9DiVYUmlURmQiUiRNRsN8FCR4KQRrb+HbvnPlxI/235HKa1nuGsJy+Xm
h7loBVA50MP+fcsWD2/ZHS7tDoIwxD7goVfutBP1AAeK5VzJkS4YVCGT3WoPLBdB
QT0kSzNwfVwx4nFdnGQQHyCL6gi8oaiWy/t1cog75KFy7EFUCcQHbdXn/c5MvdqR
mVeXxfJ5J6rZ/x4Mlek0M+zZpF9K+nZZuz+H8IUIHrOcXeOAXuQ7aiF2ZXKt9EF5
gqNdbCKvRnIWQDdyW15UcbqKCRtLf6DTEDID4/l/QF4P8Z0MgvzVQEuBI/OOZe75
gevCMEih6+IJnrQTdEndfZRnX2VRaySTp73IOarGVpXjmAdUEwQvO22J1I7+kYE9
bYHPOVUJJg3XvXpWK5DWKwMziJuh9w4hRujvBnxjyOeX4B5NlXqm9mEguymU5vm7
kEpfi8NYC7EfRTGE74Ww3BF+P3NA6cRrDrqJ1inuXfDKG/Mew1rvQ0FjF2VO1yHz
5yhuo8W8hB3P//c9M0rJnr+yeujj2Ya9Lb0CIyrrlb4CafjYlNirOZgFxl3d70bm
zG1Zf1FUyyIvL602aUHCET1SsDGJnS0LZRLCWe2GDtveyXUFCJpirF+8IvRws6nY
ijr5BFG1OoawVQ2n3BsQdKLcv267cR0e8LE1rJA16g2ou1QKYrXJTeqvxq9mxQxV
Kg6HXLKr6hqbu8QESLs9bMuuEPTG24P2CzTn1JEK9vppwmL7Gak6AAxWeJGL4lGT
TIJ9BnexMicOPzWMzftIuaZnZ47+GZNLa6vnj8kVfNkMPDb8QClKBRXbZ899Lc5z
BuEAG16TrJlGv0coChbx/wWY6fI17ZsntezYurJsZnahUKdO/jgh/WG6qpBDRlxS
wDGC6YOjCIFyprx2oU56w4/60C4lk2Una4GI6qUzPMLG5tL28TJJOkPgMcZpKy/h
hluUrWDQvB/W6WXs+W3d62FvGAaBUUerT3GSgpDWf0iKKegtttAsaPwpBkDdU/Xw
iP59zamy3Vr071RSTuhQ8YjZEV6JLGPUkGWVVhLnU++ielGD9sRFrIbApUIUHlnZ
day+sGRGmmKP2ly3n+vnfxMVCcvT247G0ry27mLZNPrnjCoaMO0qPbqNvpP860o+
nkkq0WfYw/SfsawK/pXthn6s8zq2uYXJ+IMOEMxxgj1FYVUBbNwFDCNid+rIbVsd
ozOep/qNbtbT6778J1uzOkhUfHt/P08OhZbOrJ2SnJfLxBtQdzGWWEpm13wsWNbU
BNOnfKGoALX84Qg7352SA0VKwUtdV2IQx8MgTU0GSYuDXonbnczzALccR+fMrCMO
GetB+RjT0+iAmKDYLrUtEhjUHOr7FxSrzN1MK11Semd58SPGq2mz/V/ADJ6CihCH
U+Ev/KdfCkR9EM+NN/4EcBg4XXIzfOwWEjvUHv/TVlLS8WFI1pzl0q7DB+LdQ7tN
59yTyJKZXbypqjjmstSnpf2ihMa6xJNgohtkML/jxHR105uZ/qATUY99uTy6bwFT
p5W+t/gzzV4TbXpN20wP9pqjJ5xZWoKe4YX83UcIxcXKoGNdQ7dQK1D/WSghM4je
ZgJIo+OOLbn6MBXYsyFTk+I0rh1rWtg9qxQbvS9tj1uqbIN6+s0SVKf32gravlTr
aXAPlJNy9Gz/0pIa7StOaY15alpi8gYu0QsnePmQDYtjdw2nRNMrmnYpWmvu1bd2
uKzK3FRaqrKxLR3zV1LLzxs/KnqRHVmlFtaNeBIVA6JiJn6zNJEFkLWz9iFagMZG
FFZ8eqj80URS+oVAyZNJBC2kLJB+r5sEoATL/dKiqY+VlvRPhXUgn2rZc75Njpwp
65oeSlEwuKxxz3NeXwxtvLsOv4o9UZ0la0DnhTMimCfQgN/xG4BCWfvlFhTnghPD
3z8cW12E1mWeawCIcWhNDbsbs0uYXlDY6Kxmj2svfB7xDWh2XfYt29nmMHoPLIjG
0u+D8OD4DgLaglwl9jOjpntHH9n9iJLichtKuYoWoRW1vU2FZAeISAMfyQzmj9Kj
b60hFTxVVNiKKhDgwAA6lW1OTZFXws2ufBZYufs9K+khvGiS8ExzdFG8xI615U3z
LwRorNDBUkWxeNjSc2HCsda43u0f5qYVOlWk+BTGv8mvqYTSkNLgSb+c7VSXH53j
a6XFKBB1tbZyCztpGo+RsLqfdtwAIgCWNZmMANHfMNETQ0QfsQ7/oGyLQn479SZ3
liJfR9kyW9YLdSbRrai1VAgvrbCCE8GcpoMQ9orzh9zUw2z3jTcquf8bWwSfp1oN
KKpJ+9vNTZKHKduttYAtQW2CkDHusPTHOTPMO00lczqA0Z/SACkSn8xuQZ8BHqet
igzIu1InlmNUfQzztzlXDBXRLuLBEbQA0dVd+0egt10UrLj4LF16BnJ6DMGsVUKL
uM0HhXyQra2zcAZbWAEmIpN8QGLV75NOWQ8/4LyNyTgmkIJIDeiu4YeNTiGbWfHC
vhb4LgBcUemW06god+8pXljy4Vb3tB5vkldtuHCYZEmQuSav4iKtI4FsXJ8/GLsW
La0NtpZHkiwGE027BU2+3wC4Y4qBicHN7kqhoZuU5KbbzR8ttWjUustqsU+b/Ibe
qhKUHaid3Qs5b49zMlubZmWh1GWBeEWSe9nCfwg3mf5K5Vol/G8f7CylihTjL6ut
Y+9QIe5THM5NRK3ag+dHcH+jgezRDWI9/sbVOxJUJot5MdZL7z0NZQ7OajsmaB6b
OxaSh3xnbMtyBeLv25NoyrTQWjcNVMJCduBcahMfDDCUuH/LC9BE3/mU8RRocBGL
6IqUPWmXJZUB5V+gngzJ32PaNMMVsUzsKmg+J6fvTAcne2gLRuTQ6P/HEY6kdYRI
+sVynmra19ZmcBujq6InEjIAd+VYPMvbaYRNno0KZblPjb3J6nPrV7s+gnvJvEF3
Bxc0ddr0yHqARPQo13UpQk07wjMt6PKNgUyhUMOfQc5v9+gbe4FO1+zQuAoWnbQ9
1F0Q0QR1dYtrEP4RQNoRo8llLEMdCa4fI/aI02z7T5PM0xbr73eWld1I9Dkmg1yF
JhVfO+FL67jPFTlQsHIZKO33nTq26DgFMKQAZqCND1+D2SP901AGNrcQqAAQBgKW
2NHaHEOO3AvjmuWZzkYOmsa6sU7T1F3YM0eZsf5NgD0xo7Ksi1AebCGviSFBFi3j
yUhCgJ3518EnGa+2QlRp4vNNoNWQs2KaQyrE1Z1+6aboCMEljytnXc0dwE5BX600
lk9PwYz3yYvfaVLjQp0ye94Sg7pYs/SBsFcpIRDiNU9nNgZRN14BhRsuMcD8P/Qs
fMlNkkfhnh2YntBI6+jDfI1xAFlQL0Ab+oyd92W62/KZev9WvW8MTSYwH1O16vIt
MtQM3AJNbvthp4IoEwdhUqMkVn+QpqVnUKxMnvinRLeZRX70y4dNeb/1yuO8aDS8
afWQxHlKQb/jiD+ReZT01GDpHrRhjh8kXrGZl/4RBiCtAX7jDtnGXjfKoaehtqV4
rSIPOs2OD/7Ok1NmY7Qc/sJ+uULAvzmIVX9aINt8ZKsCxy/v5rQiYxzyW0VcOYnC
zTk+fioqah/IVqAxSZFJQ+Tnkn5CJ4Dw2hjeFylQ34fN6cXvJqxIc6a90dM2mB3y
SV3FEdl+DDnGMshcJSo0dZWldHeXOQueOQUiOA9SvJ27x5hatbpQy9rmgTB5jLif
NSOyNdhZjYoVb3Q2WM+J5uGx7zGloFhgb+fSlbzBKiKH1OTcKEEWAHdt4PyHrt/+
0VeBShrPXIzLSMT7tglOeGzRz81KICntxHQisKSglqVebtCVJq3uHKSIfB91MhsO
XopXe4dRz7oq/vbO5Q3bTnluHXFrnoc75lZ2CA6T0je4PPFUlrBCr0pm5u0xRlZE
IIMdrHIhzWsgS0pX/cjGsFlFmBOgsSbXgze3wuioDhYbGFUASUF6O46xDyDlLOx5
Y9f+qz6IfoXp9HGXOKCKcscIrT7mYbjvX5OdiaH9jc3s0bdU5hD2WV8QdcNltIvk
9hliN2MsQt6UJuj4S3LuYtws6/S8Fp7nTRuUcIdiGIVB/sFpIAgXYpKSQ8voRX1i
G4D/GmFbwkZA4oLIsPVnt9OdEnn6jM8yVuKpia5xo67JZweQjQu4dxD//XlZLZ/C
I+4/axA0tJqAaxT2Q4G+FihxQWsYmUmE818UmW6SWNiZo78Xk+Te86ZF+D6AaLas
GKlEhBnIaR9u+2pqXA+hlnz20epx8JLa/NXMtmSGTjn2NzyGYaPXkKKUEEBW83mO
9/8i+sU+yw29Ll84CXYeKiOquhqIAQ55b3cl2dbFDoVALixsjewmzCQPZ0wnglPY
xPFHNv2OXba/Ui+/M24t6I8oaKTgfJ1Z8A0slMj/wiAemGyFbQB0du9Y4c1AW+hG
fnS8beyWQorz8yW5u5/CZgnHNZhtzKqyNmFKtiIO0TLdeErYGoVnS77vMDzquEZZ
KeJOdYZyl1Ujh2JIsk17J0HsuXrqgNst0frsaZsQgnTAIyjvjNbQ5hQ+10fHLgzE
cMh5+a22HNfOXCn96qoJgYEo6H3kzVtFzWjZAYO/6AEdbOCF7QLhTdTjaYQsmuSm
QOtjwyhz/C2JKqjgUi1TONmXNBB5zi0PYrsvHZW7xi2+CEZOb2AMQJWSZUMJxt6b
qbbr78e4tKnyrpGSyLFN6F1hrapRI3I5BidyqsUZESgF3EuE5qveJIUcEbmA4KmR
va53drQw0K74O3YC+OAY6ZpHVNpr8IMw1jTdb4FiKZPzrl35DopO40yJrQu0DDYn
gVn0CzjL8OL/QMqjKlpltFRJbVm2M7N70IbUUZbzveL1r0tgH3DGeqggsOi6d+Ee
poCmgAs/lPIidKmo4KX0pEZb9DeCEYoj5CXSLZWSlvpRx5iosddYRDe+4KzYv2U8
ZFtj7+hj+/z4y/h+RdtXrJO6zuX6NpnrYSaLlsj/umjg1bXVCXgDD+T/8+AvcYu6
EcNFkWPT7qNdTD1bRo1Ib+HS8EMFYbDnC0AH0vLruwh/7BO6GgpIa8gYUJ+/8rvI
qSYsYectYhojIWkhKFqZOUnA4iYHodNHITwYh2wyjizMhhKGmzWQL4Xh8zoG50fy
zNK7LkrZ9T3vNJDcCha2+lRdleqoGx9C1O556VowWBiHC98atJZDvVhwVaBWpd1n
/lNalejFXFjCQncbBTyTd7Q2n4nk5EYVUj9SQPTUxXjqx93Nh89Nhej/Xoyrudei
DUptrY2LeE/QCZ6N+aDDHwT2QLNouTWdZuOy0ZTGnKOuyIcFIjXfYlohh1eDSZV/
RDx1tUtQcglCb4td8Qdx5t5fWVkeZY2hPghIkX2ecte0cOJ7U7LNQbvtMiHrJL7G
5Qt8Ga0ooKK32SD3UgF0BhbkEbHN1uozetMM5ZI6XlecTi9jcU/4JL+BdfdxIZAG
naR0sxQLhUiAhPZOuFlOElcjXiw2dOw9A26M/pW66lANK7imOoKsot/YMWXys7Wn
HykzW5QuJmx9KlTD7NDXJZVogIPJJV+vCJoQZ+YMbot+oPgH6q3hDROBW+Do40tG
lyAkp9ljPEum5jQklDq1y8kM/MwuLV3asXuJW6hKxGLt7uI7ERHx5jUhFjHIr27/
GnNI10zpkCakQe5/g3jClOsOpohUA3NUsJMWYkysfhkrtACxHD8INHTkbvI8+Umu
RKaWCSf0HyMgoC2g73b2m/CN1fqh3PkygeLLq0pRLkx178ohwnB3hbPK0j+BxJsy
Q99txvi+6zGTLKrbATgNy5ucNnCe0Bmeq2HjG8/zckUq5XZNymz+DcQJr8+k4YCy
ZU97h+2xyT6+k5umee/qWMritzjq148bkpI1aIBjXYlMHyetgfXXrLWrnoOKk8A5
PY5ztmnKv3mSiB7Sb6smlPLHWixfO8j+D7e2odoB+KWIgRcGU8XuXAPR6Qsv+kYQ
xzRwgRVODt1tCbgI3wsTmBKSnFjD7pt9AggUg7b7+8RfCuS7UpS4RnB03rxhD09l
ZlzgOTbDB8ym2hPFAnfyi1yqaSa6ds9Mtn+wztLAm+xBaKdvIFkRvgBaDxYC5tr7
cWtY+rOfR85ngQ5QCnI2Seuv7DiP0+mzb9Kde7wp8R+tyKkDLPoSQU4J1Rd4DGK8
QQUmUYappHJulMBFcFSSXeK8t1NgL9uqo7511+XsLBGrEhLQyRbC79ncVYNN2oT3
/PcPMddpkK3e4cdl0EkeKuRi6eSqR7+A/it9b7y8Pm49QbKhDJgURPCnvcpNNGJA
LAnqK4rAgYd7r07gdYZnbKVDz5Im/Ss1kgp+VbECf9hN/ffurD4i3pLdvdKZIzW1
gXQq4C4eKZkRo9JFO/7ZapBP5kZPWAtaskh8jnbSJhCod6wZjp7KrMh7EYlpRIB2
25ala4qcb4W03K875fGIW9yL23uGufzZ5bn8qrghKb0X3sRQvmj4SiJZTD1E+coG
2Pg6Fy8aPUvOGxGgcCv916fL5GeV8n3zfodA8px5YXO3kX+2q2mU0aLBROMOI12c
hTl+sWVwC+yx3Uo7FF9f9X1QMTNnd62VQNlwUdnhbs+65s/pTPAhlRaSLTr66P55
QSItcjbHhY1R3jziMWM2zWLtp2YyTByapvPX9WJU+wUmOMdZ1b1W+RrVZSSRDISW
PvpZ1z91l1d/dlHXORaASn3cBnZLcs6N+Z6BdvIx1o+iAkQzQWmaA//u5zwYtU3E
SMqEgFWjFvcyNB7hntV/qJ4wYCv4omC2Tb8vGzmy2WAAMSMSo5XB2CgKfJ4IfdK+
LQmFFa9MNd36xsAJrYkWRRjBwF5IkyURosN0dfSg3kgN3OvGm21KDYbt1TS7MhNw
lMAAW9wmSO6fecwqBzxfFHgWxBqpzbwvnALwFZ1btEVbTEhBN9aVeObkMLfUD3i/
OVYGIG2dKJ15Sg7KfwFx/qruW7cfEJlzEjYHLeZSnn/tangZ5hwSy9mJSgXLj+NP
gQ7wlMJwzxbTCSMg+cbYSb/yTq803ef+/SttOK2lGXEqwUWRnjD2zn0Gu+wwM5XT
yZdaoE2/KrTHRrWmYx8yxblRfzW9qJ+6l1o9l+WfHSFrO3DNv9wMb67eio9/InJO
t7vo8VnHWQ8NkGq4RCupCpNcr/P5XQqFeh8mIVsCvNxNCIBREANdicGBtp2OtzxP
YwBh8AbTnO0krySkLxJ+Eqj2ghVxIZf1KMTpew2X/vZEPey0Ug+5z1qYR/Fs0pyN
1I86z2Eorv3P7YSaGWZb25Dpta4/OKM7efAABYKTnQw34ulUtsrB0LPfmzCtS8Gv
SwjpzhGAvdpM5D3xGmTa93xQF7zIysPafd6exb0fXflqSOFh2EZu1TNwmbTrsp1P
P03lv0VMVa18H527JGm5tc3TyvOKOFVo+Xzwoj6yYWMvP4D7j+1wyL6HIVAAgcDK
h8uUrR6mrVk8hbXIht65UdMkEjBklp5T6lj4hZSljcw1QuegIW3QQj9itVRg9Vyx
uVh956RfATDJLCn2rgZaFNNpZHDwLrKApyayBFOPJpUaVrplgoEJDEjNBWooxsGb
2MlVBZ36QHDlhfQTUrfq2asL4gVXsFH+qwem+m/n/ZiqMpYbrXv0E0yD+SPM76CQ
/PUSR0yaDc0wZ9NpnBIUiQEqvqQqJstxIwHEUoo9BwunQ/cOwmlCvKL+DCaWSwIA
F+v08FZh8gp5LsmSYDfxX62FCMRkd0oHzcYyVNsobn4pTWQPiJgoPA4tcrFA5XWm
pqaUdAJw+VlAyTnzN63Iw19b4frxbjnmtkV5uOHTe6NCRaAcJexl33TA0jEFPi1w
OZS2aoynvJoblA71fVIPOd0ISG76R4doQjeK3CL22poGnSGqQMzAFYTdkTQuBbYq
HHOrCioGJiqR0vpW6/0VBetFlR/PYXwl4/7IBZvR9kFbMDoS75PBEHYmMg2mFsdA
NUZYlsKwJLih7AX9rP+o9XUQqGKUdszoJ0kAJ42Bkr/kLmcBsSlEM17qHkbP6Beg
MwLH8s0RnB3eYLLbMMk87NCsnpmg/qwXWj6yH6DzdhwTCVPVQwqFDspnk+LE5C2B
NhUxgrwj9ppgidhN3ovC0FZmcxWJmYm2JUpAg3VmO2tX8v86bydB7csLCw/Qs10N
N2ivk+scqMF9GVKN6Ap9lOHVRFBRKupNkaBM436tyTakPMCkA/16BX1zGxUdWo5e
NHsQio/X5UMvM/a05fyltAPcL8GqmP8UTe/hnsmaCfvyIgwKrW1YcoDBFrLcGTVI
H84g0ZF1WQxAL/dIUpjHL2/thlcXnL2Zy7jHhQuUzwSqHLS39d38tduRKJSYsphp
QkLquEHUfIpOMzDeVTHt1R7ZSR5NnwjPHnieDZoOMRfFXtzjpEqFnVmslvtjohnf
CvOCqaB2xEGhF4iwlItbYE7dHHJxp8lldyn+GFJAiBbzLmzmrSZ6CaBJ8GWSeZtk
QIDFeIP/A/c1yEpi0G5awBqvJNTKC+SdKxCWPuF64bjpEEKsAi66potjc2IMbyrh
3auYHOcfJ4FF6Wn7SN0n832ag3fbP4CmupGqySoF6joqr+eED1dP7L2M22s/lRQb
SkT8vBCMC23SHowPDDdmZbCrq4wAJPhC3aRmfi8Co4omwKNr78By/w/2J3IqwhUQ
K19fjv4ODMVm27MnclgioXZgTO1oUyX8D2d+oZb/guqj47gP8s3SBDEVvxyUzrgw
1wMPNHU5KwDWTeGSy5mOH9h5oWpPNPXhQiidTyioEtQ2Oc6hQh0oEOcVeP+jIuCa
5QKb01gEYXcTAeR8zyUKKYlSXbBBqPDxNuiqqLC9e4CllYHYn3EM2pxB564uCZ3h
HCIjnbrVLFdGTwc4cjhbFdEdrxpH3nRmOOQ1wBwF4Jh2Hm4V5UMLshc3D50TNxoM
ieidVDjea8VUvQ5RTuX5H2VZHJw+BX/LGYdLoUny3g70Ww7ftbx1C1uWFDBZt1cz
t6KUJ50nkq/jYRaY0muE/T3hkxMbrQzkbXNUT1BQAYXx/8R4CGqIiOg+M2jYaEBY
OC7CebXUm64qFD+2aHsFvxuyopyqTNx+FuESLyqqCc8d2Yj+OIVCIu6+Sslgm4P/
yWDdmlTKWLTglaWjWKvoY6C6FYYXYhlMVpjnS3ek8iC62bod1mcmI6SEzXiuWkLJ
ljnYPJqZf/7IBHLLNOs69pReXbuvhmemHYRZVz5xumCLugEJNBoZIkJkEdq6s6a9
wLw+vl+X9QuJ1I10AievQe31MWwJ7o+uUA4GxF/wqpB4nSjAhGWP8iCPQ6GI4bam
FDivi8oxrWh2LOu07gasXHz1lEIlpn+vPmptqR7HA+echqkal/lumGFwXKW5wIjs
WhBpZWgfzedh3EPncnM19MjuhPOUz+9fKW0o0h+MemDVkHTiL+Ez7+hUePIKvGx7
gESccenAEU+v3mMAyUeuMZT1Cj7cJctZrYtgfI3LiQ1ml4wcDtkSNGGNaidxBl/t
kUu5hHbTqBxicBFK0NWLdyEChxzmXrIXaSduncPmrjpGAOzcYvMAEZgtkzzPq9mk
OJkNeqce4r+v1Xigp19zWMurtuJ7ZkGEYeSOysmGObP9DszydTWKlFwq/ypUlotB
uwVSZNm09dEhCapKGSXNTuO2LDW8XBgHsXpG4sbrESAEsLeOGL5E0Tddf5bytBw2
k466xpBBaAO213vsST/LFw0JK/A5cYn4647+F9iZiuUt7bKXJkb99gOxdA/WNKxt
R1fcBqrlXjMsaSLrXj5+mlSdJTq9odwv14W88sohhG9/FU0z3ndb0RndUo8vQl6m
PbLksUZOJmvlTCvKJHIzgBnQSBqUeSFbMKy8Gke5ojNhCWzuXjF5AZ777KkYmF9X
EFmf7kwXzoJm+YdBhDfdON5HwW4k1W32z6PSb37oH3slA7NUEl8Qs2C6NX4hD/Ui
NbNFJmwmVbskJb7BGrThb0wgRGp2XvpyA4s10Pql++MC9j3TEbZ1RGEZtQFX5utJ
spRWS8YMPURXwoF3MY/gsQGgrvGwyTZp/AUaD662wwo8BR9zfql/Gmt5fbTsxJu8
hNLKz8wGA4YUgx4rwtUpVWi4KU+joWnFkhf86Sfvpj4F5J4gvNolkqvlvhlLHjsx
3iaTpyisG/m4BaYbfnMKZdN9dfn013svqZAS0e8pghYcVQu8mAKtNISEvdi8Gq+s
hS5XOu7/tieK7xYPpTgZlr5wZveYs/8OtE+9jyIFPux56FmPfCi6HUzo7LHXXJKA
k/7+KI6c9kZcIkJk1R1n6E5Lgzxdz+EROSRk62lAF/faBK6eAJ4fwYH3sB5i0FxF
SGKJBFFBmdX0+5+eoWXVD1luaUp4xIjckedzbpTeMW433Fy6GJXU1dTNdDRQrflD
BVkL/qZysZW7iAARnHUISs9uuVuYgp7VxdqJUeROvaUA4vjmaEgXCdd645cCiwCC
Fh2FyFExrK/BNmhifnx9bsVQgq3BaqjbQIaJHMwNgVxBoT2hXsRxf1uJAWcA4wDe
tEXYYOD2sEF1M9CsEzz+IVHDD5EhylipHsrL6JTbq4TNodNSttunvaQTcWlmadqw
jBe1sIGZp+4u5gw22oz/eu9eYQOET5+Dijqz8JZ39SPJWiu6IMb0ANu+LE/ujBCD
vSPAnFlxJZnhTe1fdRDFt4pcvNIJER1GVfm/ZjuuPQO2GgWQm2eLQeCTiMO0ujp0
5pMpYQsVbXW0l/tlkH4Cy0WM2AKrZigipZfBCd5EpXTBgmQiiKoDl1qDEVQPBkcS
LOU65I2rc1pa3ScNFbkTtaSGdCqcRJTsLem5mJ8i4vsP/dkXRgnovXJvtdUuFAVF
pU8MfPI6vIRzJPC3EQONe/KCs/6QtvMXpr2IUEgUmwNv2nCrrVMMm7aU5I5XVPle
cTOvZT9R5iFVNFW7pLtTCLGWpxGWTFIztHQK49CgSMi/20memTHEayAth8P8gJvq
faCh0HnVul+0zsvW4sNTfYkJY/VSOJdeO30jMPpNQ/7A9VEL3YJk0BaTP/Z/VmEF
Y7NLo0kZHWLvkFCuGnc7F4HInxaIBJ27U3LpgH1kmfiunOxWtkcx1Bae/17tyJ+E
20m6HfBh09fW03on3Qx/p4uVbkyD42LRK2Pk7xLaiih6pRSEa6i6D7IKvbZzFBpQ
lCKGnUsC3SRwe9asQbFhhZjGlQ+We3E7Kz3ZjMMDQFNopxLetKuTEh0Nq3/P0den
hGDiKuiEdJHmP5YdK7IxKj5hcxogJ6239WKs3dl4NI3cssLugUGLKK2ewY2B7LsP
8q7Tn1/Q0J5F2KFkr29rbd3Bb8h//FebPMp3F2JXMBT3rC0YUEx/jjQAcmfPKzTu
vcF+gVwiKFb+vBgRTRS30PouvmPmk1OepizsG90OZwIkMMbpVCaxApuRkNl6EWSN
WRnIjgrGX7aYVhdQ4L684BRa6pMR7ahH8zYBlJy7ZAYYNrpAji6NoV2GfXsYiiQk
uC7Lrie7RE3xrNtgcEq0Js105RNB45RCqpHWYVSSl1jsxkl4ynTTuVw4AdRO1d3/
/gD1eN1zyB+Khyx89gYGpu4tz5L1/Dfsn2tBMz4nPvmtGplgpd9VwtN5hq7DCF7w
8I1YavjU+E+SJykdRF3zbdh81WAse9Emgyy7ksd29dAo2mt+YdpMrjlW9IRUj4aq
XvuvnKebJ3uyLh5w6ZUGnFax7jHEmTPfqUZRiJJbzG2WhYnFs6SdJGRaKEV4zCAK
tVsnq8Gh12OOmMrgKJQ31s8VGpb4PgGnpxc5HJiepiyJjLhRvQLY65WhZcB/5aH5
m/p+fdEG9wib2nONfOCpDiNW7rK7J2deRlr1qZRyeRDwe1P23D2V0W4+hkr7mR1a
VxHe5dbnigEj4HLgbQQap244exujfeoG7aEAt5QMCzMPqdA03VWfj0P7JOTcw1j0
5DQIetkDqBG/z7Is8VuZ8+kvVF8TfcR6x0LoXChVE7HBuWzdT9e2w27KS5qvuwkd
Gr1xfL63dMj0p5SwKB7m1VQpAUX+UyjbyB2NdMO5OPz61rJf9UGiUaFdcdRNThkU
Cizl6r753ApD4byZCjt+fyobIrZX5aBtmI/T+JsUd5qk3y3l+wdac53mVpDlLVKT
+y/Y+kmBTHDpIMJmiPYE8JseYzNqC0tR2goy3w5vZSyUEGoif9dXQLIgjddCzBZM
K16QJqpd5mKEZxd1fJztqylGP+5A66HEifPzqP+4wnqJac9BaDBlrMwxCBlYzWpP
B/62buGs4lXREwX6TcYOuoZp+7/T7BJyrgjK2yM3ZZViC+6TINSgqov1pfuutEDR
AXQlkEDx/0rsPPX5nJtSEEXCGiFOIcUaXQvn6RaeOthiERwSuFo08bCPCV2mImBc
r81qrCfUdx8Nbj+KudHwqr/oneCdNi1dE/2RVNctf/xwTdm3sPf6BMaOKtTj1M03
g6CDhsScrWl8/HSmXHMdwuabYZ7FJuh0iesQBw6JscwcAeBqJcGHOb2GHGG8DGpT
I0m80j1g7AWQe6jey5oKJXdMnsV8zNRcrfME/c2UKP2oikTTA1lrColAExZgn/HC
UZUU4aeQu4HaCd7PBQCIqR2wQ2XoCJgxdiO7uILUr+ebBXqB03Fc7o1F6eBzD+W5
vLa+VOO0HdrKW1syC1cJbXShyRdfNuD2kh/AJcvxAd//nYbZDMZF2yb4osJxpMdb
e+fs8wu+3h6mFYoUviffFMBjndkJfcGz3kNVqp7ieRqZl8wliIOJR87y6Mp6OeQR
cZtXcbc8gigHTAQHt9IjzWe9J5LP5Gn15l7GUfGASk9IA/44U0q8oAPKeK5Vpb1E
Ho9+DHqfqidWBJmP/h0bQ+E9RjRoJfg2cvPWgNCLum+xWSVIcvDHxo4tzXx3dALe
jaC7GmRUmKH3mTpzq1rK+GDEHEgOeGMmfgKLlC+4liI6XDcINldOBaavpbzggrIn
1YIhglua/wlb1dr/zdFXXxtSs9oVB0ImWeXYsKQVJ9QCpYa4wNN03vS+JcXJj3ZF
7Epl3iiALVWZavGialGH0i3rh8Q9dyvqAkT25+uMRgZy4dzHezU58TFktDDKOsLo
auEV26e2udBshJ4dT0Y2oYLZP1lATX4HdeFRT0sPGKUIxstsUTqHdaf2AzioUP/6
Bn7+oh5ueq+v6IRaCQh8Apk8t8dSGzeQB/PJGjKSzW2qksiZK3t16Ybvk2L6lXQS
jFxz/KVqmX75gqD6cNBE7Hn/A1BP/xDlyvSthutCU9jnJRqxPL3GKvzHSo+WDqlZ
IBWw3OD4aIvnZZnDAgx6jGnrsQgUWNy+nGOH7mU9PuJnrA3CG4HtjZuMfDtc3GSl
DshxLwtqrITidSXWNfSkK+PfFx3BNzotVfem989laL++4iZX5iZpwQ5E0ARvWLeD
rDZWEFz+G3OVLEoFAJMd8+NjabGPokpm/uVRshHt7Z9zIyg891ab6+0lYmqtxunm
rIlPCRCRN6j7hz2/01hfELo+aN2HY4424Omx7iOOjtt5OBOLTGQ2QyCNYsApvjb1
dvCn3L6mKdheudUT8G40ZidmoD4PaYLKnZ9WRzBnX1Hn7KtVbMZ+ogv+jBthhZRd
o7tWseuzANZeKuslBHCP7XPLT8xYkX7P+4YIT0c4T4C2v2K1S74lAg+SZExYVtJa
ESyxTjPDxxWHYeoDlllnmALUT49aFhA0QDJwQzaPoElc5WfXem7VYdlBYwiZJVfN
A5xBo0inpupcOis/MJMUpOVo4hr7H+IFSH/A1dfogAho0cjbt3viONGQ0Fsfybug
DXaTjeFLhgsNJuH5wWHkp03jeqfO4Zb2ZTN+tBRGqL2Yl2UgMTnZ4ecC2hGnjYRS
tOPjxgxZ7+m6x6XXbtLUAAS2qu+eA4/L8rd9YVs9JZ+Z9vmZsqxDy6ueNrXj0BM+
uILoaShGOdgbMedUi/R5eP+uRrIQx7uo1PBD+EnWImUL38Q9QhlVp4c9xTakiaH9
nwmsj0cBaKyVBudnGfMYcKwXeX+JH89V0rskD6rE31ZQnd0jTOM8SQ2b+dsfhgTr
BwMROm/+D60CiFr99iEqgq1KLoG3gCMkjU7ji6eWACEIrxirF0bK9ujgxqx69WqQ
Swd7FTXX4xMG1OFvaIp/6ZjChwjr8lsDRMbU06Pq8yAfn4kUPMLXOsvxGazPWZq7
f81OGLTtb/XCCq5Oqn6Hs81KgNwE+UA+AMGfeuzOOEP/qSjVAy/dj/2bvMET9iQR
2cGhVj0aL5FymuKmC0pL+8+3Zy51OiXLdNmrho3LkdVL3FBQiFhtEJeXGfmFHxCL
joPaLeUqeoZg5t/Jc7AKgW5+RyWTb8q6NZdTXxLzkLAFL9A2SlKQfhpNyPVcJ66T
JYZokV3BhQ4yp0Qiug6nqBw9JOB6JtiNEXNTLNn4TsR2lfdYGS61TLJpotpFSyhR
esRp65l19fdC/gYSJgwzXVnXzAZFYz4ivI8o+6iGtJe3l53/AF3n6YtlA+dCLb7a
J5jiIcl5EwKMNWdQv4chDMsuLDhR4Mt3jdlvWCzd7H8PnnaDgXfjF7cKEC3YmUtV
sIg9StopvVetTBV+u6ROqifXQL+EG5HxTYP6YRQgKxJE2xC4SgmZySR235hs8tV1
JDDtHlZ+FgXFeiJ4xr6IERLN20WbfG56BlE1OUAymP7JP67h1B5h3fpBfZ0ClUY5
UpsSrmsDJKoYAcn0mchdjAOWgb+0WkjCMSWIS7VwE5uoe8sspUsQsATAOzB2sMa8
9KeGoC21nLHMHD6YN0hk4VwNfXFhHeQp/erEGi2Q1WUWiEBvVNvsBWmEmXvanfKv
vhFX8p8JE6Q3ZYf62KzuF+c/yDbh/tsu3uCbLccaumU6323oNfTOTQXuWXNrtgia
Qc+BILWkTLFLhHdq6redZwFMvhECNGoPZpd4FGKEY2tpn2erjRYdmOvtoG4qttvM
utksKmJczHuUbbLRbB5cwym87Yy53Moc5dQ0Y65umwj5YUcUXE/1UHh22wXjMeGV
QxfrLbyAiieP7HbJKy8jOtwreXPY9WZMlfnekTfAUV51VUiTiYd2U/4d5tgIOjc5
eZDZyDpqjF83b495VEZoMapbyFAW2g0yz8OGd50feNueKBsobg1qAsRt5hGGdVH+
L8boHXS3EvFFyWm7WXoT7FyKkS8XUOSVDekHfEDuyUzYu7Pzv1oUAPSA2cyeogo0
XjcJnk9GvxUKcmdak2aq7lyxwvyI8w+dDPbGKyO0r5JoCHOHzCRn3VzxuNWdulyB
dvZFLM2AW1kyjz9jF9N1bgDclnGTKhdaLTcmwPWjeXIV0n5aiWLjgwojIGcV0jkV
mxsHP6taAzLWZmq70idza25VSkxLyETtEjwzeN2oAn1lu7FJh7Cg4Dx5Ylvw98hN
Addl5hprq42nCyl2dX3lOQ5Xas+Az/DhP/MG25Sc92ca1PGQZ/tNbrvUl96Ebmbg
5pUaS8o0N9/rLhQ9Vp+vACmHicEvYl52X+F9Un17uBYb+Xf3f/N0MzXMrrvL4LC6
+mvgCCKVumpxCjuzvjElDbV+B5ZK2uCacu1sYYpFh3oWOSLrK7FxMfqtDUPe2iXS
HhD2hbG+cuTFRE8YFLEPjH2zcXHCGZLpd5WAMt1qIrgs7W33VjYP3lxliEx3IrRz
0YROWv5Q2+pxrHdnv5o8EMHy4MbJ8BKUF3AEVsU1A7w2aeLVIaroslO7fi1WF5Zx
AH/VeSSimQ+yVd7cWKRk3+FkIm3MCCyXIdAF9cR889RsWx2aF5HLKhDWDt8IEI6t
RKI5XoQp3lyI/W7MoPHVlQ+Z6CfbAl9IeJ+AxKVmoIMijAesIwdxmAbMLvXCZH0l
+WHD5aDzTMcLdoVe/mJnvzo0VsOjO2RR987LxcTs3N6UTOJJlEHD6NIKfaWLo0LV
MXVquN2Ha5s+i/Fiz7ZgOfEtSp5V9kr7FX5xD+sPEPw/s4QBQogkLnGjsSC2smfW
CoxdNFteml2/lZooNg7Lw7Oqesz0wI4IUKcItvFj02VAxAv/Pc5+5RPxvh1Lawy8
sGm2Yhu/R4/m/NmZt9l7SPr64zikI9FU/s5YBTnUZ91Z7fKyeAVlNgM9jhNsKWY5
XFndvpO4J9rfgDRikXVglNB0ps/DiU03x5X31aSIemFrjFZT7rOrXYAfhvFyncTQ
oj43NjBxNVF+tDN+LYE8QPWeTrtau2aDSXNrjonqFo0wkgFceu93v6h0CsQpAsrr
l9qNhPcZS1V8IF0nISX5Ql8hNkEH5OTFII1sA+QlWA2z+LMnGhmNpul2wYOFOsEs
4ONHF//A/hosjxO/ghYr+DXE69JaU6glR2ZRe7KhJ4XJrdPU6ot8tQn5xXIAphWz
srIkHe59EcAbapOzCF6cIaxWD5Uf0uGl/6RR4m5jkXjJZeVyiekme5vOcm8q4lBa
aHGE0F7Nty+X/gnW4ZRM+swyBCw4qHZYYQtb/KMyvH87Ec4kTpY26f8MIY1R4smw
/+h27sEo6m99gsJQimYVNVKZP+OS5rQX6Kk+9IWPV0D8uIUMXxa4fVfIEgd2ZYP0
iev+LgTec9vFbLhSgOVm13wqD/36JTtcQ885WWiu4jEcnDZ0/nAXqrumqywO3h3A
TfqghEX077RzuPoCHnIYfyQl5uXPlctB0/86jVguMFIjJAAB2EtMYXonxE/ZtzTo
a+zh52XaqudpXBmIG4mBRRlrny2/JYU62XjL1VoJ/Ee25Z8PJpbomjtpplSxB7YZ
Covbvy9iK3rrLgw1MkyDNIiEoemnrCPhBXgyu3UOGyUA4pGkgaMT4c5viFl4BkG+
W/jIG0LeYOq9vrVhpj6aT/NBNScODSG8+ZBDXSi8P2zxsGrs0nRLw9NFz4a5mv6r
dt8aeb+c1UEH3UQtqvhBIkfXNDOZ5w8oyNKke7/UfrW5Uzs+lZAMJDLIygL3+Lpv
2+2LgJi71BreRkwCbgkDLEPeXehpFmlPrSc9eXhZfClmXqjzjLsmewnsN3+KX2tf
Em64+cHCT/htBMKsY8RtoSa0lm9uqBLmZaSyXM06hJ1hxPtzbAfmvqQTYYFcXSPg
vEEpyqRzwgZitU2bl6cruuxNHyRroVlEhwZP1tBGdpu9DkGh55JYK+Ox1k5qxhyW
3GZQgtFn58CrUQhevrKan7iNuYOU6SuF3kXK3ylRIUTzVLrYkignc4wokctHr6YB
FUT87/iS6Qg+K7Azw7XWOiie0vp0uVvjJpTuC9fHNyPJUbfc8oy0Ae0nNDES7nWk
JFJS3niRM3Sty1yVnIgwtQYUPUZZKOLY5ac6pQFXfJxuiqbFgZLEW/mTRHyAOjQ6
prtY1QN68ERxrD0tZpLbFyXU3uCbIx1eWE8FzQUhZBEs3+2vcs+EO2YSkFyo5bQ/
BjEV7oMx9EclxpBO6pbswE5/dr+lL7oTMREEveDcMFLqENDimAL7mqRACnbS9XaR
nIaFrxDebXZ4Q4D2jPEGhchp97Skdv8HoT2MBFkqInKLB0T8pLm9/mtCd9poXvF9
4bFYNf904khWtAHSKEv3Nc5pLPzkJG85bFsARP4FmC+FZjPKRCgl82Dhs/KFlImA
kt1e/RTXwF/NCUIWlVIAhUPAZ/CCqmQ/MboWO5y5ZWv+j+Q2hbg9clDi1mstkfnt
S6lH88b0qOVfu/yk5egiaUqKVpLJCh3XQ0sXuUenbS7HQcARdUIKAknygaUOPOpM
qx1bUBz6l+YbolLJhVLkFgr/ZJioUkU770g5xuf9cKN+IKKyq2E6MGS5oARk8jtI
B+oo6joWSFm/ljV9E0CzeERxXL9VLojQZFWDTIx9QKCAvE190tDJV80qje8WnLdl
yoFJHZ7LWmOsbLg3EEB8iqufBlHx0Rau3n0WlIKH6WXw+yj/wXpNFhOnMSuVdVuh
DhqdmmUChYlyyAbNOh7do2StM/fHuWzNOMyWcLC55nL0BvaeTbYbqnp7KvQVGs46
UkTaqobDDUzE0LzfISfmHRFrNk6LgsvJYfS2rHFUwzd4Y71MPLNtzWJ00qc9rXoM
JyTlbV8BQ7/zWWzZfDRR6mHz4CGO8QwuGHtrIFIgqwJubW7WsK1fFG+JTgdCl/Kn
WxNF4Pjmpjo7vOlUYf9d5NB4gW0XwFB7RNtZ3wWAeWcctOT2krvV4lMP7bNIEc1V
Ald05PvdhxFx/zS2K7ZH9i4jbkn0sFsfdUNNMP+NuM/ATmD58gY5VPbR/w99qhWC
Pa7TCvqC+UmmBvEmkdqdjEbNr+3xMtF4IkVXp0+12yI7v89z/n3ClMMnNc2A5J4h
B5pyeCLqBR0v3loCkb1A5j6bngMFC0M0byNYs9RI4yJ4/ELpubpvMlzNmR1oxViu
YD4NWICs7ESM55k4F0wJyHXVWUnvqwRKrMG4HF9o2o0yY1axVpQS5Esa2/MoKBWy
4XXfNsuVHgq9v5sbbW5ZyuWRbgQsYE+Rjau66/LRbQ5EdoFRNQfdahH6ETfL9asI
FQVHA8FH5D32+IjXFWzBWYqZ0tBjwptky3kPQcacEKdu9yTDJXQLqCM/zAFvRUGL
VUZHBhMRz1oBdVUPJqGEzbDNYK07NhAI3lJn7UJu89Z8kfFBQuwR29cgvLNdbTJf
1o6OmbSbEZ4wy+QUCd8Het4ccwZJFyvBgikD/Hj+YIWcIthjPU5bKh6DCrbKQK4k
BEtM3wx83w3+E3CmW2RT/ShIu/wDqpWMgQSfgwrkvTdDU+/AawKUt0qhWREcUoV/
SI4xlm+XkWy/d0wwk+C9v8v4dZbCgXJC3lRqJ8VQhD6WiuNgcmMFcUFsU46w1leN
YGzivB30uqGYAJDxtngbQzcmL/N0NykcPm6GQR1mjiP/pmvwaEN5ofWR6suxKrRN
2UpfL5ux48SbGjHGbIrm4N+pgl3bCM2dE7bwgNBG64fsNnAWseq0EVT3w7kgHRck
zqj7gm/xAIvmNHkOGR5B0McTCGKNCjGxiyzn0FiKJeki0037a5rd3OrhIWSzTZKq
YiTSTTtIy1reHLL10HCszJNuB66h3a38cTwASBJeeqz+mXZz2mLMnzndXIoEnuSl
Bsxl9HzzkBnKCBIJBDA3Rprw9KDaAiiozdoyIsgFl0o88Kckt4p0oumtQDkhxOpU
/LI32oRosOuJvUu8MzCNvxIv0KL4ycabdP2fMQweHr9Huw60KSg1k/c927Dl0R6C
isHIHoQMKbft0X3dzqo79J2uMlYYj/LrmqquQrBE9NT5OiVBntb4t/aKP6kA7au5
XlpOFg2j2WtHwgkPDpLNYnXtIy1inmx7+lJhZHGq/jNc544VtQHEXpbIPOadj1wD
jtTBZGPEOsliZlciH/M/aw5/0pwN6YgFJ0heMWB6j2NkvlHzLnpXMNfhwNzPg+Wj
9fVjipW00QNUPLeMOBwUv3zmfxVZ2RB72sBDOrFRS9cEaBsyJYBIFWGt0wsx+pLm
oXS4GeIXqsM01zxxYABBcQkj/7PM8idLh4lA2DLo3+TqPmFScVC4wKXMOIthMsop
32wiHx14Gg3Va8zqCrfLB6fcFAoZV1O9pr9N81BuEODv7s+JRWoD+ZfYeAVlNPlu
4BeFtYOQfJOnQs8Xkfe19n8esO4U2y7juM5PE/Kh01+g2PY50hQsVSQxuesIcs9m
TO2HONug7EJxt1+clhrQHZr+7LaWRQSxGrmp+k0ehkBURQbfmbzzi4UK+5kGYQud
htxOxpb2D43PhqyfU5f1DmpWnkHOXlqdLvW0I2mQZEy0tJaGkqmfpOPBkvnTFQa3
YZ84fWxq7SQ4Q20Tw4gxtfmqwum28Q1XIBw5mA7hD0SwrqxGIkaN2ZecjIqpogN4
NsZHdJ0USfSe915vwZkJsXRHwlAdwaA+oMKecd9TcrN6sm5DSDaGW0Hr3tGFWPWJ
kV/+kJFaruBikxfr1vPvzsXXwu+jkmlVI5MX5xplAS2GmTJSHHgoTnqncDhjPKYV
etrL5kxElwOY3hRbVIXWVQOnJRMG4qnvnCDqu4K4RTbBbRkyJYbfQylQV3uC84wI
eutdLgBV9/PnE3KYECRlyJwzkUYDinjeF2hLTstUwHEv2EIfSSMm5Pi4cKwn+W2c
g0OYF0/2IbGThomB+LDVtgbE8wyQaA3G5ZBBeCR6JDz8CaZ2RSqRWMXibUkf+tWr
3SdouPT1nuM2cJNLTDU6VBmZMQoHkqKr3J0baApu6o0v5eZWL8ACT+ItIQnRf3j0
GkiKZVctnbHnqg7P5xDSoaTMSqBPYnvB/qzO/IBG+K0x4IkBGk6uh9JPMbbbQYxe
t91Ltn6kUFoEFZrUQMoEFvUJdZB1EezWsAiyf6GwbMLaXrG7lNY9ZN8fYSB9y+iM
1jpl45YYs0Rt3RYTqqYS0TfsmFJ0GEzJGDHXajJ1xBpmXy+Qs53viFdhpRLz1n3X
/aim4p6UfBweR11psyzpOdFX2mJwaL49nqvUfGmNLK46YF70qUlKoq8kZ5FYWY4Z
F4U+jBtX8WUAxmAQGN/BwnWFLbn33orhVndeqBmxLtSS15kg66jq3GZ+IMPBVPrr
vJLJRUiIfcMVxRM7RGCGoOtJZad/WGKONCZpB7/9QFhyYejLe7khOZaXaNHIWjrd
qPGIzvLSMuGItW7895OIdb/Um8qMbfqJDdT7THD0OeNFtwziv8c4X9qWVW9UWbx2
a/1EizkA9FWCFtcvkzSZbO9iInh1SZVoLPzaZqZcdL7yALTpHMVDeDAZip4zQnFw
EVKBYKaWxWIUfdvNuOpJiDkXpRBzOvUmxDrlDWduwRL/NUhyHwXVAU3icawooU8n
Bhw0GZsCz8Yz7fL7Szp4w4EesDCKK3Vtq3LH3KXi59RWpWqoCDbOUIWBewQ6tRQZ
1rfDGoUc6+nIbAFfKk3gqVeoQg1yEqT1bQn8cctLll67/OEsXlf3818FXLmnACqF
m8jktEMrkoqcfAZkPUPZwFtIaELWo4Aw6l9YdnHVrdzJ21OsyV+8C35j3MDcGpNW
faxDkoUkwENRohtzREEHNOYosEA6HutoAQMDOQoZItq87MAMzydb+Z/bsoAHMLkU
GxVDQ6vfsX4VY3vMelwqJhNzrsUvxHTF97HKhSZ/JZi+p+WCVJ1WAWwNI7jrV4Ii
46WptfuwMdKJEUV8hCf6iFqSpB6WXskxW3Z8lqxKGuuUUXRQu6ZzxR6bpaHfyQ+0
L55LQrUsO8MvSHtMbj//aEJINXKcfoc2N3UUHzKMdizwtCXWRg/f9k6gpvnID6gd
dGsEsj4SbCfW/REV8tNDV1AitbjEiF8IAkrwPL0IANeeMZDTEHE0x4lgrM6yA6TQ
xsSl/crUSLW785hSwxYl07ytSI7jDjEgeV3R1pUmklVm/DeVV9GbID7swMmH7sgr
LP6egsZnc7lRQ8OIWhUQmg+OnYEfTZFaO5oare+m0X4hBAdpBtdSFdVydw7Tvs1o
LXyWNYOXXtPeTb1wC1wOJ0T5SP3D21jceb1XKLJCNprumbpDR4DA+6T5XW+qHEd9
6U73i/XCUAKQXZ7Njfc0AKsIxHAO2SERJf38ZIX/OvBeWT/s+aON8d5/HXxihGR8
TBskH/xfC+ZJqEiC2uTf5pTlIJomiedvPhU+LXOx6rHZnLSc12VnlXgGkWL2XEAP
V4/rt3I4eXK9Gr/bBDrguZdhq9mgcerEg7BnatAP1TFctBdtlWDAHJBeFft5+e53
hxuaA+AZkBWTcQZ+5Oaa2tX8KNw3cAmj79i5xYVxG6Jxzx663ktl3Udq7JUDu15J
zfQvtIcsrykM8qqIj/gFXU7Gpr0qKhyM9y9KdytRNRg/CKDwty2o8sx8GzLywb0m
JHhB8Jn57I7JzjEr37Lh9gODre39Zd5FGBTGDY7MB9j7vooecdCk4rFz+xS0TuxX
nz1d/1wyc+Zq2RUgi1KPaojtQzNLyXJ6dPPudm+/4mc3SKeQbr+dVLP+fHqALOnn
Q7YnB09dJ9XLfZ3ilxIcpCcdAruRqEU8JG7ZRnoY1bGGYhnCW9Tdmb+QknOxz80l
f89o40fMhjizyiEp55WyWNv9LLBQNPUzxoej3Yq8hpu6P5Hu1iMYBG23nENJEYVO
n6OQCAoBTFGIBw5MD0lLnqgBCym9Iv3/tNGVAJBEzRIt/04JXig3bO6nDCklrbKB
NIdLYtxUhCPAGx31AMjdhxkFTdeNCPjunXMX/CGn7BlIuwl2m8nokdDZ2cKwvRiw
/0I2PAAthX4o/Hbc86r7okx5klA4zA5ua01sz3BgRm/XXzTkyGuD1AZLajKBy/7G
4IHJZJCff+slkZizKcMddCHcY9f3/0OAAEWIuFwidmKc6Yw/xH5qLPGrAhF1XCs5
65DuhAQzTl93Gf5b3zpZHg0LNwr9w8+ih1i6VhyrFpEC42C8ByxSYMFXLxQy3TkG
RqBfLWYkYMV4R+jMBXwfZuprW5w2FSKRng5PGQuJ+hHTmcDTZugpn1ZaUdMwK+2u
hB6QZaUnfkCJrekZno7AKDF9RQuBkJEe6kavYKgOFes9QmKmcIBiMoGhgoQoU4p4
K5eS7Fvq3oOHIXNXcTQQOoN/00YFM2szo29514Ks9HSMO+tJ7BZW1/NwCh4wr7tm
4U1AHdI4btvVaDhu0CPHxVZG3fqNdfMHCMW0OJLPdGq1JLTMODAvF3fzD7erf4pq
JI9N2T1usJWQvySv6E5A/r15rpHwn2T2H1E3pytvPtLu7qZppoiTsfWOGOFPspyS
xp2roCOpuxA2D2saPVlYej2mr+m2RaPqqQGXl0aYC1th8CcIKS10lbyGF6NWEzne
LPNdJpq1qnGeMs7VCkcD8Ez9zenYBjee/fN54DthvBSg0fQhOyffw2cgVNCdbGYP
vJ1TQue3xc+0sYcLlqRvXMSHvqrD+6wQln5LJjLtdSN3VFq9WzJ7Q/4H+v2qmajv
L7LgzjWPSAO25KVRPCxt8IC/7PV3qjP+Xn4KzG+UK+L7vHqv4OYkGHAhx5pHMIDt
MpqGWIXks1yToWkoxN+dmNkEcbj80uSQ46RfvqEj6Zi1I/VX4/drO+rLMHnDKsSf
1xk5X9Jwig/f5BZOyjJ+8naU1S2ausrAvbiLPCNtoAKsOi3QrRuUtDBf6eUySnTa
4k8TGgsYX0cn/98hfjkwP/+7j1/V5FZ5BAByyrp9Y7DlGJ5Ejy2JrGzYSYEd76+S
9YoshciHC2P1+IgMOEqQXz+H71efARypZe1oABH9jUtkMLU0mZXn1iY1QQiQkVJH
BcppEjWvVZx2edaMxKX/zSIbA/AdGpVnWTaJbw5QYyckIgOcO2J+Z5DgOQpyPW0G
4wl6BlUF+J9wmGLWu38p9+Nq0lqT06z4/QQ+fmRe665xqQk3Nz1TDqMD9wsO4BiF
Vsztamp17BUinSqnDcl5pkcR3+rUPHCcBE4SjnYLihZHVEeMOaPvoPJQGQ+ZkKb5
6pGftcXx6G7rBExZe8LDAMFr8u9vaZ1x4ooSYmgGwaykxwvKVGDU5dclneT0pUZf
2mz8J0TlDL/ajfX3vd4eCFZgiHEs41+i6sRLSdHaVMLY4uAU37mYcbmGXTEFbVY6
qmasFyM6SO7t69e39rSbCUOl8Zj7cQDbERyLlB+7eERcL4Y6R3cMkxREQXurn68O
oSh+KnmnPJtya0cizzZMU10MYX4WV+MK/PD6APi+95UJwY7KACJLsZWsuj30GONN
m6wnZMwoYIlZAr5UIWw4Nv+PsLfySxBYTIWtspZ7TttwUNwpePXq6a7D2eK88hYd
PK1dylCbFjS7OKZep1foluFJctNbmTrriSkWe6YZpyXB3Sg77AXG+LxO3leKB0hK
dDfH43Yv64L/QMlP7oKPm42N3mI0K6dBM8zKn14aeWblcnizMTPINhsEsTFHM5BB
VtB8Yji/KjmYlRYc8la71bTUslxXKfRN+Zofvhs4IArGW10BHNTIqkofaLzlM7QM
ASc6z1wbKhZdpcTpUbf3gaPhZM04xGQCPFKsWsvMeK7vLoAXXdhO+ERIBDVf2+yY
MpJOLC6RgXI7cJuy9F3mOgo6dNp/O1U4bS3qg8w3D833/zLtYiklMkBRiWX0CZ5L
ioB7pFYoJYksstCDfMZrcvxN8HHSadBRLm71vAEE0ErEIO+D2PdmsydT2rZgXgpI
uAORG8jFyH2TVMrNE7mTc+MjoWrIJ6klI/SIMmg5RNfXPGH/cvLa++9mhQXj1iqM
5Gwx1O+thswSQG2ESCh6bshm1CGC8A51Niu7i1q2pyuhxmC6MUs+mvl4xUX+LPZV
s2EtVrcCMQOBZq9xpohW86Ws796BwNsXDJ+mbF89LfVvj3N1VuhcoQOXIzE9j6WM
m94W4j4sihGn6uQZfH01qkRrjC9s2F+LPu8kqejZFZZE81FmfcUYFLxuxZiBHAI9
Gh2+AHHZmQB1WbaoMVR1f3Rp6H/tZ+KOmYsvKiMom+8eMJdquDRkNVGCYg0Vi95F
PjhWXPIju2bTEz7s7JVzTG+KAjHZRlEi66OUxxaqiCR61FGAdmrFKngwTNqZATdh
h7SyWPyBnSgmHeSkE97Pmgd4DwzReuLSW+3aQOwTvzfWMg47lhpCKq4thBy01CCq
dBRzLwa/46VA9SlzcP8egpe+P/HZSyOBcnKQ8p4JajBSKkoKtq6KBi0djEBY0W+C
ud2pEstFsAvkhgG8U7xVnxqGFB2TFfZ4eb5Bxae9GCUVHqN8XAPUthyATcyO7+4C
lgRbhIbP8x61RHQUgVOT3IvbNyyEFJPEX/evFSIjxVbBbffxCMUwlCxND/m29cdk
IVFpnk+0LYAwPT4/7DY0F6rRMS5lNTVDqCsw5z4NmkUwkUfyA3OmomD5kDIMLrl5
VL1VPrrxQsOIvL4u5PNxa86ah9RxZo+cuVISX6Qh85PHJS9xvVncHt/URh39klE1
FdZk6U4x1sA/SPlKTgjgo91YqB1WTpyZJM9v+oaG92tM0KVm+/ZpbJYNaU0Ev5+J
XzPR8WR0Btwb7Cb3DumnD+rnHXjQ9uxUFco8RMZpjFivNYUbfYPWSWXBaiPKSpIo
AxDcsnhzneXVb6MEeGvgb1irWsHLFcR3wVYBUVFbmumJ+qCR0UNSlyVHJ47eJrGY
7BsYxgCidGp8oTEV7tMuq3AFSdIAUgDcyNSTTN/4IufCTV3AvXz3wg24QftxBDv/
pz9hQLsQJYmiFIJ5APNseD8fiAlQSrCGpYGWRQc0jzqoY2PC7vjp6LEvv+IftLOx
2gbssBlbqWDkqqs1aMAD+4rIUMvWZD+arFTp2FIkKjnTtkcInbKJo4Tr2se32Efr
RVoUE3SbFWxfn3Fzm514GrhuYDeYogltGY4QbTahH+hNi4G8jTVKMy00Sv0JUVJg
9b8VQE+0Eqp2C9SAQZgu5kPFJ2qk8Wp5NSJMpaXtEdlqXTAaPJLR9UKgQ5AHib5P
+oRJqiTQN1MUEJR3y+lDJuG4acczOEpzQN/Tbay6egZxRYgEv1NMTIFgSVHv4l2d
BkRE3mMymTeYHbjpaZJc75kWwKhK6dOyfuzJjo4HCsP6EeC5iSkFj8zgPi1u/1Tx
uEM9tfZUwgdAUylMHeayxpJPYrnlh2SlW8DUxnyxzzXKdO8n++sqp2wIMiANVsYS
qrYFvrN483RXdDNU3Xl5sw0l31UWl1TmqhTtt5UmfCmdas1JibKIJIkFuQLqJ6TH
CLiZL5eEjuHOf6koxhIQHpmv4Wd/2q4ntGA7NPYwOJNh538Rji0KYteqJckb0pd0
f6PrC1aF6wmFGnr5VO3SYCEureizaBPH3HutIdKdPYAB6X7/v8LfxNy8d0p4+SiE
TjcQ1zi1IIvhuYuA9JARYGzirNp9WRve2NnSbTpoukCfqUd3B0vupiHI52tt2BjA
J8rg00LuWHkuaCibde/U+B0iHRiLVvPswWRgJfFJRpJ1hr8NQq2HfT+pwWGbPT8F
ZDWuxWGBc4JMBriNDKgHJJMWsS5d/oqnRj4ng3ONp6dajD13vNXT75WYBBrMlrHB
rOl111WBOGeXWm1kbr06ZPsYMqKUGlLrXs0jKfUXHWvo1xkwvNNgQk18amHFeClu
8J1TsTsNTig6TzV9oYuEB760L0Vb1YfChT8FoZl1Z614IyCGyTF1YB7rShstbOXr
WGOhhpSj0mt/1p3bGcb2OtWa3FOcY41cnd7iVQaint+DexArDqJmPSfTsDMS0pZv
C3dbDeGqh07V5bkpVH/3GNHeB2sEQInXYr2bcUFEhzgElKzJU85jkDUgPpA7CJkK
ocyjgWruJIDYjdJHM7kzz00BLRlNhK4ZlYjRGyKm8WjVl81vfnZsF4PxfrCUh6o8
v1A+LhB/aKuNUCFnuqHjQKQ5DLhZ/cytdMWrafNf41/7BVkDep/bQbu8AY1iaqF4
fuYWiYWk6aNADZwC5z9vogX/VMo+2lCAKzhnHgt3Ygrrt5mFED/pHPyCZ4KPCdJy
7OMfahYd1KXn3KzunLLNMs8HsFOCo/GqQCJB7gGmeGcqEdSBT65PrpoWj2X91YdJ
smYFBSmabezVVjswBkslar8suQfnd4fLS0NmKt0EAnKgUvhenKwNMK94QMqiKEww
y0F6AS18qr3QItOaDXAVnDJiLMBwSo43b11ezEpk1kbitw/Ga9bmjUP5i8MjVVSP
1o0lm9lKI3Og+Z/6KVmtRyful+W7XE0Ess3PKY+mkJaYXJonUYhtWrk7SRToSqBJ
2Wfajc1QJb/Gfk04aNXWJZIHYcGfl+nDIGIkySFHq8AX0jtAaNhZYAbgmz4WKik2
HVgV52SLLm367T7izcf5Xy7ctjSN86BjF61IYkZklmBS+sXof8VhX56Wfg3NzREp
NvaiH18a8ut2Sr4/SXsReYDsIb1uwNF4Qd5gva5jlsOW5a7UhMZlyn2s/WDeUlH9
JBUDQZpv6yHeX49Bg1GFVNKnH+Oc8bNmFQauxGv9MqtBZTGuLXC0Az6XhQ+zO0sE
bQK6Y3Q7ff0OA9T5VaZ4kiGnECr8aNBN3seX5ft9rzRdNV1Nppu+sio0DNIKocqw
OengIzslt4Z71aqw8uMr86oH263tTwA3WxGU5OFO+9xo1jOi5CVWIL+O796LerRM
hF2XpTL9xGv/0WTqt3N1VPwy8hAYv5QMTfo+800fEhqADxa/wzsUTggTbELCo2HK
4ay9ApaA77nV8yUvX7iUQ7Nx5w6LElieM9PSnv2GybLMldImYs3pRO4horAKElH4
b9xH5//aPyMXkbp99IHoi2YujUh1eCRP2IBZo65+oFdsXe2bkUQ117Px1GvXTXQD
1c+6oNgKgzeE0GN+NZQnyImgcKgIFQcS6tVRywJJtiHaIjdnZBV+BM8zvW1ZzS+C
7G/d9/X6Sa32LqirEhuJsYS6BQnkqKbacruVRdgNDlQbpa3Tt1VfLq/44hW+718f
s1rdJak69tgNOPUndkQn+XXXTs61jTrT73d6iz/V663eFpyp+9CUMBok6NZyHuQH
tU0gRb2DqTqMneAeHoymTOUq2rIyikmSkVicPUIJCkLNTZLVZR6QpO0sxJJQ9OVW
gUl+UJ0uRB2zDafS3Qt3qX6f11ax9+IDhdiBUq8An5MMj4Oasl7qk1xLXccB4+s1
YX0tKzBe8DkS4uPn94yrkmopVPFFypGdXgYPLnoPBHhvnClWVqc0SGPhqk+TDB9t
Q42QqcSSpgV9rmjYNMC0lBCjc9tl92mqjpsc/ACTpGdYndRVo/QrtBgL+uIrMeIh
T4MFGlLaDw/Ct6e4WLV9xd42ZWsvAELrh+nHUCglpdh0XqDOkx18FohqDCXEX2vI
fdZenD6qZK6uph+1EEYotcoFSUM591o9mLok7ZszX/AWvrZpE02XdbIdPcSfWnCz
1vqZOiEUx8UuS1F0UIwpTa11QooBSNm5He+i4UuyV07REIXD2T5B9TdZTy3AFHwu
XzVLj8HO91qNYaGzPJ8x3GADqm8Yt0+iEpelYkBraIIn0tf0kxgb9OEG9/7MOhlE
x+5/w7GJ/ccSabzgDzG6EdewrculPSn7BrWxQna/u3wioMEPQHZKK+dZw1uJqNYq
s/f1ZlfOWmUJa6Cv5cb7OaikInLPd9nDJaBPLIu2oKP2XTaWMMrEbK967gdOGLE7
tgC1+Y6Rd1uFxzoqYxlO7FFH28MOtRNw0K1KfaTmvfyKjcCU+ZqklH2+Ok7l2rBc
3Sc9qw+kwczvVm980kDQTUcOqyrxNX6nBjnKt0o/P3yD61M0y7cnuV8BkK5/sgu8
HfS9LJO/+vv1LEcIJCRDjXwx6dVbVt9bL8KBsHcC7N1apzuczqmYtZlLZHShCYly
gdPB32ADbUbotHZXR2PSl7RUFP18GUn3EzEfKmUrW0KLr+5HSe0pA1gHd5Oo616e
yZTwKYiooyZodDvBlWgzsT2J1Uosue2MI4a9NLa4wy+/7j555DNdj8e5/7QDZJfc
IVA/8yiulDrssOOadfWWoMSJWEauseFcdx0H2AIxJW6bkv2qSlzpXKuypWaKrcd4
Q2GHidxm5lcmmoc/GxsXj6ky0eSu9Rr6MFs/kCxFbrY+S09L0dJAhU+57seVxvOW
ckJDL/mmsW1vyvzhgfs+HGe21Cq6PouLhZ0QRuW0sfLMirr/o/JsvwRQ4FEBsRU6
LHfO2d4X8Q9q0PMovlliGLQvAsLQHWe/1P5n8U7qazcIVflk6yZufTUoAyzeUIBN
k89tWphqT8GzPf/BA/mClv5Rnr/2rf6Kk/b+mP/GKNa/xo0ULEv1iXU2WeHKuJjp
xCtPxW37mADPWj5yqQEmiY4pRXpkzHZZATFdza+OynTbUJdv9X3fO1sgytcEBInO
7EAyFo+8EVlDxZjkkjvoLMx1DZUhyjXB7qN1fLLQ0F6tSR8IgXQviCkpGFxBcHeX
tvREw6OJUoDvRh2i8QlfPlSlz4aPMuGtw/abWsR0aqgggTF5d1KQ1YgobfKzASSU
fb1YBTTjgyG9XFiuxzTE3btBQY+OneaOwKZcrPCfEhj54Z1LQGnlL+Ly76RddzXd
8es7E8IV5K14T+Tmy9JDTLc6lncjg7P1poWDfGJXAfyBneFSZxEJF/SiZYcdqDG1
rCVXPMFcY/j7dqOZSjHCNv7YgKUMAv/qjV77mz4C8lPNHPaZpKq3+vomCQ4nItD3
wn75AjBEm/oI98zBgPrWNfJ5kvzd1CoA0+mjOSXMRy9ZmziXChilF8rLsAJdDEId
EpsCD+jQZ7U5fiCrvCQ02O/MsZogBqf+BSuW2CRN92D8ri3UfJ8gre9ufzoxvsbl
Sawr4a40Oll7ugDeGtLZ4QX5brCA0CyBHIfKTXmjG4IRYbBiBpoitFFqYuOcXa/p
Gk6KYm9GaSCMSh2eGnCrEKbD/BN9fuJOrxrBIufvIdcVD/+XPcVhbKlbc0CF3f2I
MqN/QOtYT+EjXP2u766amRcNBWzkOOilH3px7GLObqN9VgPFUFtPHqGenzDhPltk
jQtclVgt7aX6uIIN10XjkvvocWoaEFQLyrBc05hPEmSTSQvgvM3c3vhiis+g94Lx
kGTTB0gLuiyhGhnp/ipF03NOUJ6yXbazvOF5dtA0ZHfYoURsEOnDIGDQEaa7JDLR
dtncTuEseQVvS6ol7EpVLzdXfUM4Sd2f8GNfuWWIY+9lpI+ZNkh9R/YW16laPe8k
bfvFOXBXkXXXLCBsFhml0CbFAoqdviCu5nEVn87zC+a7kuqt6/zRfSvojH6Hli+S
g3kpum+59ODpMBjKKjuMgFhK8WgfIKgqi2XfVaUzPXPwvaZUD1Rp51w+7KLBGhx0
jJS3kuhNy9WrFy5GO8RZrQ9v32uqs2H8pCtCh3PysLZK6m09Dp3fEm+cCnC9mtx0
rx2sZjp3J2+Wr4jhXEk55CnN2+604Y1CFJmyTusUFOAImc0X8Ia3PCno8mTfQJVv
JW7L9fb+s95FEKy0qGmwyZoINVztP5/pQpGEeEg08IC0vfLC3PvU8xnDmUEvD0VM
eIf5ES+3PuRfzdE08WGUd5SXipeuf68896xIfkJY4Aw9EX0ypbw1NI06PkT29I8A
caI8C+4lQ1EkGb6jDpYNRikeSbzH0lZHCIEPn2c9Rpx2k9IqAxPcbOvp67iBh7a1
TpRH/SkCcm3tJeYpMVgAuOpAU5vhKx2DIiycylzxX/udxPfJHakZf3TE9Jq+MPgT
7cx9v75a6ukB59c066cCBxiX4CGbj7S7lohasYJEl/60UHWYl+2GRPvmb2hPVlha
pCbxQCuz+OyhTdcAmxVLiZtuhgiAENLbk3lRYrCRHtpUsMo1IqXH19ELjnATbPfM
Wyj3QLfQjtrSK8Cw+bWkaXWvfWPzY96sD39Rtr35wvZqLXcv7whP2dGEWMqzGyRd
yHpm/VW7Pd/e8nPFxNaLWTvD/bLIG9Is5f9ekHXdo+TPPwrYfOFpWjeBujE6VoWN
0zyVzeANZdaFWmmOOHaFJMl6CXgGOme0GsKARUPvH2X83nFNjAn+X2hz4ZM4QyDX
n2RXgxgRHZ3RZvQBPwRPG06wK44M67kR2NLbHvqqK9beJQbBzP/Ui1dnDtbh9auG
Vc2wTYA2PZZMEnlLv0/6PqR8xWlB980wxGf967BMZ+ciVdTH//kuJGf7JpYRxtgM
bqwHy3SsMCiz5KprRyQiHmaRKKL/Edma0wfon9/TkJuZm4M9nVjilsl2XsE4tt7Y
LdiRj+A0hEXjGOv4Pk7pF6e0pBB9Qrka71qIrPXYP+yaAGo53zvFOFN2OmpNNoPY
yxfN9MFEINyE8vQ6jpKefYSLWCqh846u1fshHYtwD22IyRfoUYJUkOTD8qla4nYw
AwEcv1Na+TaUyuWH51lMn5PiBm6zd5JYSb34pPLFj+DXJCS7Ha6fuTmqHN7Qtkjj
RiwNWDWjcow8R6jXiEdSMaYm/GtKmC3MF+RdqP7etCVqBxPfldNxrg/KYtioeITm
EIR1yaWpoC6ar2UTRUdbi1I38Mgv5sGaU9TUKczh4fEPlEDjD8DZtbxoxQAoPonL
0wg7QRALKl9IQKEJkclqd1y/62StO8W8vkPxZCcDzZHNAu036mG1OYk+PDgmLE6X
JiDMCluCj2z3NyWZ+M4HB9Rc5/IkLr8IuxZFHefXDI/bCHWFirrySr7I9H7RySlx
ZZcvE+1oaBpbSimGjzXhq2qVMCnjBqma3gtbbGrKCmsTaypk8Ak37P+axZ1GuH50
yIWzMHa/vMGfQL5zj69HXPLmuy2+uYkcySBRV6J299akxQAAlMhGvr0KvZKrga0A
uyagaaapPNwds22hTvlsyhab4n9BcjjLEu8G2JAryWAWmDhJsnO2WcbM9J6sATw/
YzcaeO35mYUviMTF6HJ3qNDwAxgK5KaPX3yJlnY+pxjFKfDE2/sLSd7UGileuEKK
f+bhViz3NavnE2dQzH5RlEcpPwbYPv48C4Akc1WKSW2RsqJmCm5bBfu0KWauNjBB
U/xFjf85eXtDJAmQfJCimbWj3ZT6Iehjg3tWIuo+PR8j5t2hq3n3rbgeGqczK/ko
eC2HPxAPi1EJut6s6Ca5jsiG0DQYvhOR7Uk2eUPofuKmWbsukqEzoKxZKkzg0YnX
Ui57ooa/rnAoZPq7xx6jwJNyTv/pd/7yQI/BnqzQtEP92GU0kay+KjXl+YndnIpU
visckjAouVKkQpPZ8haG/rUy0lPEAKgALok3inpOhFTNCLmf9pmnx5Fpmy+XdAXx
m4Sj7QO+j/zMLCCusXDfLQIsRiBbbd9L/W/9OePZsmDsKYuAe8Nl6+k2sx1r55Ss
difl7vlezjmy4uo5WI8Ngh43SGCXsE1JLuvoaTUmf/goFBxemDkxpcAu3EaUmTkX
TRmWRcY3SMxCTzvWUJ0ieCWe9Sy4xCq4sCQbr2fD1p7299jWy8k+/JBg7RA/XbEM
xeOtxEDuuKRjOXa3gy4esmDg8mJ2Xj86sMn6CwcDe4s1IU/PsRbCXV/JAbebOmG5
xlf+xE8oCgAjzpBJ5aGu8yhHlnmWYN2t8qtE8L7IsqsrJ71vCsck2BTwMOwQ60UL
bfPMABsz83OU2k3Q7RxdG31BPflDgox5XBpL02+SRrtD4yIAq+ODBejxL1U0juVa
YKCUw6PjgEVeW9bWzQfyVG47VUwrHnT3xPczWtdG1HytladLZbJfhy9zeb851IAd
TmykmXdqAnP0p5Lyb0gb+ulBapNJ/KSeqVAE0B/pZMa2DHkE54ft78VnY6je67bY
p9o9GwFafVmcl5zjHdWwnMb8VTKO1cvGIKJWelEYjlmJ3dIj8ISsXQ8F8aAm5akC
6YiIzS+1Gb4BlSbC+VlV0Ej9mXmoDiwGwwQFgalBeJB2xx9xU9IvCOrd9TyRHkb1
ut4KtmRO15uIowILSBJUzd3JjuKxRe6lJAAASDxYDSoVcF97PqbPIC6LAxo7urEI
zBrSnn3dGUG2yjpNmYFer111pXh9YVCUJ+FEiyegoE/lXIDW6M4aHCixAMS5X6YX
bjlFSi4ZTbGpKcgHtj/6Jhsk9ISvBHxL51iv2jdLblKVUMQHKsGPyWeDpwrzeZih
q3k842aIw9EbY8RpEZVYvcKD/1nnSEahqRocpUSzpD/m5uxGROkLAMckObt2UYqS
ZVmhmZcEZvS5WrFxbtruT09cQTTaUELZygXjcwZloNehKUZKsWmumy9c+F5yEU00
DBYNEcb78ELvMOrvCXn7+1y8P344eX0Htvp3U/SUtUcJ71Uxl86wtB1Z22DpGxss
vH+jv5WUxvDdRvPftBfsRx+T6lJ7BcIAkVRPtzsSH+3L6e1VZHlIcCnHmoh33JEt
R6FpgbNsaaRvmPYzyRUHyL562sYbau9dWHWrkugCiSP28FOARo1sMpti/ZMWVuUT
act9MqEaajsBfeN9SbuVoR5tnDn/xd0Tvx7JxTFiU1R5VcPDgDl1NtInzl5ji3Kz
93e8BrBg8RK54xtEQYB5bE7NESOy/SqnrJQJYUhb+d62aPC8AJvawlk10pADgmUr
u/Ys2mskFgB3fm9/LHyIO/WehEq7pOzoFocLZpg1tmc+zL1hLcss/QRYTXRsyEJo
5CiSDORjjJgTEhgSzam6b3h7rgiC9hzUHTpLpx9g8sLj2EtR4aHX2/TqkPgp+JCv
pKPGWeVifKzdvPaE2sVgJIbvUxE382fEbe7OpccvnaUUkwMLnLntEVcEQvsALhqV
NJY/jgsOYOC3jMlkPgUgcrjnUa4Y/7iJ3gJXborH+yTX1yUvWGA86Auo2LGjNpeU
sV8ac/YjUeQIvjg9b++iiDyw7Jr5zSMqbZP25aQB86+iF4k9TMpRW9dEL6WsmtVn
fys1leMelysKrzZ68/JPwzoZkYWhgU0LfI9KdcQq4RQMwU0ozgkB0hzmIJPMGadQ
rQl79ZOAB5KOjDokL3mn9aHk3KYI7Urg61ssfNDAw3Gz960bVtDezT1SBL13DZ4c
4twZn9wieCLCuwoIPjuIt0RPEwKHekogq3zYiJiZucGaJ0n2G0oAis0h0yOeTjjt
gQFOW+370mCAtAGj4XHS5oxgqLsZRbn7H2eeC+DXb23VfCGi4h1xd4c6jzlZMC2r
rXXM8paZAryf+3B4StBCuIKRbfZr/94TUwjyQuZlcsOTRrGCZRNgZicBr2gA4jZV
Kq+iMMJQC932kjQIIgx/spgdm4/jzfx5vh0zRV5OF7Fe2kuy2E8W8+yuMO8dN6Dj
0YyrbRsTFTzSbJilePZx1mRgALGEuFFiN5e1vkbR8q7cbPFBzVZyNnzhv8w8ZElG
6H3fFz0QsaZkjrnbsAw4vdVOc0IzHuEK12YqRe1d+X85ohipvm4pQICoPZnwIfA0
IlPfXAIu8mOnrhc+zsewDiSekz4s4x3g/nMwh89JQh2VNB+8BrLIHmDmV6UMuRDO
vn0msEZs7YB22YaKgkmcgmq4WKZNJUP4b+1yeCYehtcfFXG2S7oyixbMI6pTchOu
F1KfPqrtUlM6moGqYwi9sc5wLFEaMvJiZoLsFB1torvAoX/cKX5R1l0C2DuGA/wU
v13pO/yypj17hnVBBBwu1D00UGD2bER+WkcO86w3GK6KL/dQ97CLGHMCt5VfdmbF
kEsisLDz7o4k6xo5EQrNErGnFD35nkIqSMVNswGPEsItvPWkWqNMkm6sSqFa07j4
J25gF6RgcDFsbKhpYu8HBTmCgqwARPq3CD5v4CbUhxReXIFpbWyhBhA8tdJ3/zF4
lVLPJCW10ymVwVu7HNdBgTggxJ1H6kUJUDJrgvdVk5pxWEYoKamOmrPBASE7beNn
dTiZBvYzKxykYW7lME8UhHI9wSEUgxQ1s/u64JPVJL2DDTLuX0yPdrDIn4drmCRw
shlVDJPbZvv/58e1txdIxo1ahfGfd8ldwfrls+DhcOL8mQHVsSA1Lo+L3MH6isn1
ib7pbrjA+0l9MeG8f40NmQEa7J/UyupaFm+vZUZ3m6A131UBIARmyn9re11kgBAK
jksZTiL0ODF3R+YZcCoyUCzJodudZi2syeq/Qs2FcLiONplmtM+hY+nyzFQ0XINm
WMInR9XYhZp1Lpq8sPTJgpd/kfLpnW4+hmOWatdWMN0/c0Ys0XgnQfVwNFlNaFPi
cj+xfaP0cMbKT3cyJVWpowP+hrIIV5urmBIV9I8dpdvmSVs3XMO2zmyAMXh5uYyB
AdBNVfaJubr4ul49c42j7z9Ry4+5dTYHvHi60npIUc7hCKlUHdyM00G8uVXa7E6Z
iNu1uk0pfs37677CjL4SIAMYtTvDDUt/Ac/NCUxPlkNwmwbjRnPsDHMON6RuxX2Y
r528etIXeQ3mFkfgX5GyuvbvDQ5laMThLEYzfBhvJi0TLN2nKBwiAXF25bO/zzNF
GtSN0uaXmc0nj8i/Q9QrA8umg9M/rY7Otgqd2CSQpfr92QOXtHrrHYMzeSjceaCB
DFlCAwYp2cOtDwW1d9ZLPJTfLXmzp3wJ1XOaZ9U2t+O22r5vVVCkQfcI7VOdfCzL
TzdeN9GhQfE/6lh6trOjh0AEOtUW8Ku1cgfOGxTbkaC2mNBE+cKplq/IHyOk7fOS
0+XIQlJ9rH4pb/gX2n/SZvQRh/5ZODiZVMb96P1w8wIOTGXVEoI/icHHehWVIYiV
ChF5k0ruWSgOwgQYYJb3ma3XT6EY3iTV7LlMit/UyBpZOMhSXX+rjDVyRxMr5dHY
P1ot9/XFa0yvhUHfqtMhsuTyZ/ZOfN1goV/AUJ+IqOGPoL+w0mg21pe3ZJ94yKWy
xUMauxDgmgbmlEP30X3GImfFjQiXsnng+3hi1HjqksjNNfDnZYPuPzB5hf2BbWyg
+GwkX3ADjUFCsWZ83F5K5DHINt45M4P7lbmHgHYlPiRzSGMoJQMTQjTwTJ+GWmYu
LSvOwAjKMC0xKgfMri9B+RAGdwnZDEy5fSpkdWZussblUAC7O3qSwgf3+c7/36O8
MuLDzmJx7wi65g82Q9fH/9Gp/SMeXE5c+ZImudGw6MXBuuj1HPIz9CuCrcQd64I7
z7ux1xj0fdTXxpVWWBp1CZu80AWC0Z+JjIxRyw1kNoMR6ryEr562yOuFpHws+mt2
Tv+UgUJgRQrYx40icQtabfACYdovfO/qIwWipy58GXzIbDaorwFxQTJvSe9twc9+
G6qYA5WqLG6HWbsKIOk/RY0g5bqZaRU83EWoKv+b86u1hivhR7MD36II0XLltGEN
4aD9sc6+GHHyc2kHf+GY1+g6VjyShqQ2EVZMtvknScBsusQ+Ud62JQURWmTiV0RB
yso7OsWWNFtayoKfja5LsT/d3PnzYwQ/X6WkXZ4E7G7CQfL69Kv3+y+C/u8v0zRR
cBaBaUNYA+d7jyj5sIo6iw/eqwfYxeeL+SX9OVE6Bk0O1+7SvamtLoO2cf1psiwB
15HS4mRK0exAcOeS+tohIJFYpCh2JjMWCLtZxVKjDTL7JdNg3pwrGjH2HY9r6xH/
RC10zQEw8uxNZNSQceDUnMXw9B7awY/pNihIYLaPBcM9U28YDYhRbyeIIxLCVVAD
LRPTsjowagDzLAh2q3+7HFSou9BaLD9kJ8zT/7Sa+A1BY+pAaq0+Y6fsfaPWvqMb
Xw15CfOaLpbGH0HymOIf0TeuqLeiScq3BOwB/4HSMhVawL5E+TA8AuN838Qr865r
Nl10i7peTxba9Eg1+HRJEZ8jh//L7CNnSGI2Xgxoyzz/qo7mpAZ7BzVauYVnbgOY
ogGBnW8g2MmY+QE4kgZ2in/u2jUNoLRSrOQyHMauO1daQQjxVBLee5waBRew9wcJ
mlfRo2PROcvEB3HzrfBZah/hDBQ37Wtvi9FGqmetG3AFL4k/PgUvcPL01HqfxU0A
nbWvBMzL4Ki6TOKlUE3M18daKhFOCMAXNSs4NtZBYpr7LaATIZIZ7gE2htrdwDD6
mDKY8V4aaOWveottDj91qWG3cxpjwNWzotAikbQi4CVX+boRTTZ41OGPNskVIQNp
Y3tRE3ZZVQtphaN30UnXKkJvc4c3eL6kEsyXSJP86T0aOhtX8X69AYEsh0nhDYDn
Zhowe1p3RtkkZuiGgy1yalxKrVhHK5q56OpWRMaabssvYskuv3pm0TQ4EpjrI2iG
UAoimQY4qZaQw1X8EOhMH0q7d5XjYuGGJF3itbdz3jDTDGbLcfFUpcxcouWHfi7H
L8Qzk4mR7T5mL/vFEjtyfCcv8c3acCMyywvBGk888F7iNbZRv2GGdd+5pEzoOvPc
Hp95De1zbaELwYzPj8d3kq9TyzS4F6BvrU7MQonGhm0pTWuSdwp3mo00ZR9AErZ8
qLe5+l/Vk4ODRw6Ajxeh27f8ZjbvTB5aDTlGK8VJ6Zjao2/5meXMjMrHtd9RZ7c2
1skZv3v+TniAM7K6MVzri1PgjYAozk40UaTVtkxj250xQ3NuhlH+FmwosxvHKUzj
m63Dwcwro/8NNo8E6zrQwGEm6EjfaCBXhMMoR/MlqKeqfKKH+S4epmBOX8EWjLOK
YT7qI3rvcfbwufhpPo9mmLZBtYpNMeTZ4dfPnSaE6xaNCFU2JIzYAiGpaqUKLAvg
/NIRFPKUJ2sMFc5SIG8TKGD35rVSdi47Bmu2TDcCYIRmY1kCy59LS0xQIxfbmUL/
/3XmpR1Q6DGWkK2aUxzgJ35RcNTFNR1ptkhKxwAskHQcPXwKTMkIrrevN6cppOKk
DWed4MrxwT1zYCuHiZbjztFkqFTLvtApCSCJG9KwP3LQuQtUl1TmbkFAiUq60Fz9
Jc6tkan95rGpNS1fsDiVvLfX0WZJ98O3YHCUR7FzJPISbcKaXxpGl4veqTI+6Wlr
2oO368I6pEPW8psHcpAZVPLPF3iDRotob49wweXent8kuExqhe28hbdkVgayD+Vq
RD3ShgO30Gsf5c3ucUMNIi2pDV/1P7DpToA8zL0AAp/KVojGP2KJuoZV72WAZIPa
c7DaGVa3wgGqy/a+csc22OPMhOWfYTWe8qaiEpaaBmByy1HvMnmng7MyQdQYORCP
G6RJ2xAtZvQ4r5HIr+U7SnynNlBEJ8s0SXQFuQVPPZnI0OQGLwU6i/GovqAg6ku1
fFR/2sx+Jq4kDV+qenC3oOrHlbvUkCmRAZWe3RDkbskUxxwcTSTqD8jK/GVmccoH
tr5ubbu/bkgUzMLYDir1Q4GbA0TqUMbCxQUt/UfENfn9RwBUJX0Ib2YUjZSPTuDl
UWavPAUkpJg6eo84pn3MaKZCo67KHGBosrYOfjPtziFI82f1ph3sPQ09c1iFCNpg
yH0nOX8ZIYyH9p7EXZLCizcljgtj+70zHB9+yWQd72614aaJ+0nwjT3swFPB7QZS
XcU/mwuZdx55R+CuEgdVMi3Fwm2hBwQ2oRTaXM1Xcz8Ml/0KnXgeC2Yy/eJsD3Py
Fs/d2xz+xAdo4msCJvQ1mqzlW0EbUxkKpT9SFiKSSiUufTLp7EIqruK3pqsexVcP
kc/pGR93FZaZi414OY9ptqlYxDeggfhfNi/kvU4PWHIEswijTqoREiTV1M9FRQVw
mXEh34Im6SPUzciZoae1LXpoklwRODsVVn3NaVWaKSmRPsVeeOqdIZJby198/Gpi
EXd1DvxnPiOAgEGWKLpUcBkxAIdhJ6OHbKyssLlpa6NlmqIeLcqR5bUDUdnWa/iE
T1XEMTho7Fv5OAwTqomIiq18OxFmUS1tbTdqeMw7s5v3UH7M3mIZecgVjOTZ/7Kk
sZK8hu7UlR2YaYeFEHJBlMSmLQc44EI9Dijn5eLuvywNpV3f9eclKyebhajbPZyi
jaTcVarc7sr09nO+4QoYSbihnJLv7oPM5uw2Kx/yKfYBhWJIevVmhpTWposNnvLU
9VZFqy7NwQzXM0C+aLtIvLVRmk2C7FURmqCkn8yW2I6TQ2oQgslfaSoqLt4QJbH9
m+JZ4HifOzNZtaWosv3oaMuOoo7gGS1tIGjlOwzUrMYA66g6Crg0N2xP5wit4oH1
+6doh4qx3B+Vf8CpdweaWu+fwBENuEg541PJCQkKHmeJ8qJFk32+XoRJxxY9+Rib
EN+xMXGsfIuE8sKkHEgeYJ5mOeNxo+Ldy6sIKOYL+xT8Z5qpCaCZXLVAR8NvxCwa
DxOw0FhlktFSAMS70gbVmkRjKK5iGVD9JJqpcjLTeqDSiB0uzEaiNDd+mr+sRUR8
7CCjyd1B8EPijEhEeilnEfsS9/DJezSpXc+1w6hlkTErkuNhxxtEs3EnHmNfN+MU
MkLeak1B9i+A8UfQI4H4Yl+pCMdzGehevQDPYWM54JEOHWGnqop4xxd7JwtfnW7S
DZ0g2Pn8XpUSfEmUaDIbsJC5pbewoL2B/gVI2f0o3ERKOslHeZssOmaSjCyd9hk8
8VItW1nvdXgiYmqK7nQVVcyqsRPFwU4+T7Al4pqtMOfcgot7m12zXwI2iG0G5XVh
J02sE5xlT6AfYgnBYwnrSEDUUPbVwxMt5tmiOml5PPtfl3P570KvOlhi6XiZXNKe
+x6USpAqX1Qit06hN61yyToCWSmbBzly/fnHkgOe+QQl2eOkylYe78Vt0+SVFyvR
7Ni+cUesM3LxQFFaBULbPlqd6LLrOIyUt6dBsOYyD9sjp9iTOaIMmFgn7br3IjiR
WF0o8RI2Or27d+3EB2AHYV1UTZ5/CpRCgzlRd5FD0EQ9RRqezmGt6/1UYF0Fzbs4
dZcwgY4uJe8Zu+e1bWxuqNt8wULA0mEp7fWwaoCSgHSkVZOLgsWJPTa2I3TAzU6Q
fFOh2ERy/2yVYnlF96lu8XZZPhhk0B1uBOHz3amatkoQIjq+FJ+tbS/FZaL7rCXf
wYNxs9Le3mv+ignq/NDzS2S+AFO0mPUQ29DWTYmCIWssAP7OVAkYucN8JEDqIg1C
tgfenBA9oFQVD1XGjCl+7AjhPQ3P4HkaRYxOgNSZPTmNO6bFxQ8VZ6JVCTyPFI0k
wMo6EjUFBPabfUMzalVHJ1P+RweYoXCQ7tptylFN97OndIQLdQlkH79Oa/HFyxU0
6laUom/dRpukNRg2SGa+bF41KNqw7AjKqXLFsDSmLSiOO850IU6lbP8iSjJQRW4U
Mfm9J0iDHqz7K9JLV+fbewcvpow8CYUT4bSg4Y0EHWiLZGakQgU5Gisix4v6jo/8
297h1KzkHURKEyqX/hpNvvGlUWWPM0Nr+U9mB93ctDQSppHJXy9xtJrBjWvCd2k7
eb42PA5k15yfZ5Xqpzo8RPFv/bQyan0VMx3pqdzjpf1aZCzHcTOYFQHPw1EcDSSX
Z0sXJc18ebsxbS13nr3M7IvNlcxT3rz13P3F5N+ZTN8MR0c+R+9bEE+vyUgGMSfa
bPGC2MfgqwPrE9ThfzHKRwC9qHPyhXatS6s9HBuHa05vrcTB2TlBwZIcpY0n7r00
Y55O+BXrYRhqXkB/Ttr2QzzmQBQIZ5knXRIGDrgKDYI2YTeZK98fYkeYWuWdDmBb
zy/M2VDMMA+6O1VnWQogWfZ23G8H5J2qGF8lXFs/GkOJlA4IhTGNiscOB15AWpP9
bbZCePAmVWJH/HPL/nycYVvn+/NX9PObp968ZBSeZ7Z3y0RkBz6P9yQJBqyzGMmy
HicHzvsv3m8vvUoYPkLWHmmAmYdDfh8RUDoyWkdLB+nBNGAxkVN3TP7at7CyPKan
ECxaDdkft0BIj6TW04omxiN30z5GLcsBGyG/xxUlbIgluWZrSwZI10iBBGZteYBp
tIaJ54moC4F6guMjzJKEKqy+ceMTpgh10SF4WZU4neHLIzlG/YQPnDRm6kGPzn0l
yEruYAgmphOA1/ivFEN2mF33+RAi42nDQclUGNiUIdBLiiB2oICdZT3pNOdXXF5m
9uVidw+Mx8hSYDgClOMGkRdgoUa/bkhLvSsY4F9UsllyiVHspW+FwSyYCCM/NHP3
SMQRaVuNsCR9LHHmS0NWZcYiq8zcQm2z4yVqgantLMGQ08f8HjATRbrN8RhH8dXY
1FOFHy6qx6bCHG2asW8AzJpfgw8lQlfpdi6aXI5S1X9qn964WHVG+0x6CXLshvj8
MOl4SWYeTXNvYdRZ+3w6ohEQGijWjcPUwiC5FkOFXKi5VPIO41PQorNsY7xWEZmu
WB9Yx5j0HNVnBbjQGsk6d3lwfYvf+fW1R4qc5BKV/OXUGcs70JIgVjNwoJ0b+dGA
QnlrQ2fCDDjcVoF4MI0ChKr2bz+5hLT4YhKpgyyuCiHN3sH03uy91vSnLUMACxLw
9h0HTvu61X8f1I8PR7Sg6+fm7BHIyehIsqfw56GjvfkG1u9xPyYMobPygxi8YXPy
gSCZdNyQ1uzrtM8E61oFWjh6PLeYgMlbKB6O0HpFHt15Cp5skC5lM95hiSJCiSFo
KzYebY8SNO8Df6ZTOyJtin+2RTWIhp3IgcJZMr6Sk1O29VAJRst1bhlWdBuw3k/g
gZNIAN1ozxLPaskck9iUJgzqg5GeJuXlUzguBZZ6ZDJHecPQ1vhlrycxaFL7jjob
89x0Zea9y0ESezvPA1sGocnnUFuIwPStXTQazIj9YFXSYxqT2JZbVrf1PnEB9Usf
9oi7blpS9lxaQkbikvG+R2s0hg3lIql671Kv5kOcip5RR1mrBj8igH5dpnWvijhB
CFEW25H7MvMOTn7idGEpspoOgHZ6rig5GYhK07IT/BEGlHj3NpE2Fy5H+9Ua2fM1
mP6zHqhTQTcNSFNBwEFrKO7lAbxF/cKNbQUiF5nzhVMeWoe7iVrNkv8hejuTDi9g
tWVuZZedUB3p2o1OF8FRErH8/nNBk2FtlHnJvJFG7RZm/lfHWI78fJ+IOM1rR5QK
8knRMfFf2PJybfBFsW0iBYL8uwwNASYmPERnuTtgDlBmaLL5wb336gcOL4r+Dhbs
uYVk2K0hyW9CRXJ2u7/8wDTTS9CnmzQIrhhwMPDCZcvToMePVFzvFVbpaclAZw6K
Ya/Xv3kg+p9hJzL0I0sBQ2BdeBuioca1X2Ek+Z2lmweMD5+xxuOaZwR0HFcY9kll
Gms3VL5lkDs3US9Dds18HQiesIQGnBx7PvS+IrA2f6Xk7KJZyFvSsLqe5iZJaPvK
9m7qP7iKYys7e2d8xNuE07FOBi9cgGQkDduNP9NG0794TdJt8IJSlDLwgVsgn8pb
BebvVBN3vy0Q+hCzNcrgSKVexEX3rxGEppIYiLt6Vv+Pdfu/F5SUcvrnrHsPuFnf
LelPvTCSj9iiObF7qmJTxdHOKKM7W/4HEoleD96MOyWHZry13oCORHfuP47T3Xg/
w6frgc3mfeAlAQw87xrtKr48HabUWZt7lRRUb797xnUvqV7SGm/CD70dRY+aPsLr
JZ1YpnO+YdXh/kkSwQ6UdtJfd0REmnws4RBnkoPjbd4A+JCBAriziIerX67M2+YB
R+gzbIN5PFVwishS9SHB2D/yprJc7h7k3tZw3t0lN5SwcscMs4WdN59HYeWkCnil
RygFx59gqi4IUAZ+isN5os5ulyYkj5sodeDxpuXNxKU1sJdeUPyqUhC80XzJECjA
qGhux74c1kNwA/x4D/5+ufeQAs4eDb3K+UjhP7kBA67wILkD/2b8jA7ZW6v//5k6
Qg7rtwYSv/RZb5nLY45Kz2B2rbMpavQcW5vFYO7MDWa6O+Q3ulnOZZFa3kpMHVYJ
yaZXI3t7RxR1agBemo5MSfWR1Ep7DFVeHcs67lVpivdSI8qP1loF4n4uhtkR5cqO
sU2bbMIfU3VcmVQLW2l7IGijBO4fFq7V/PppJbcj8hE9qxRBOIXwDyZl1pTzJ7rO
52NPevu2Xr1sFqVTXIkFy2kn/0iOZIiCFGZ0dV8Fbp1+SiMdZ4+Z7udrgedQV7WN
9vjdphkjwcRSuFr4J/jyyoUT7LBcWsbw7ZM7NUqOBz8SZiirh6oLrcVb0rgGF9ez
iuVknkzXh81aCYEP1U5kY/cck5CYNelQM143lVsoaaFI/j5NChMUBxYXUaa5L94a
6bKbsZSRizi0PkPyknDXjQS4Vcq4rfqyUv78LjyhgDaBHj7m2p2J2U/98/Q5YxeH
K9VMM/QIcxWCkPrRUPe75F3hQ2E+uC+CRGSlCPqeQx3YaqjGTu7doJrwU6nKPIgR
heLD5JGvd6J7vR9V+g0PUgHt43MdvQ33OdF6PWW4FUAqdCt1IoRxE/pkvB3XGiSE
5c8IiHnuhWRuAVgFdVMq3hXz8bOnB6HDnhmGSm5z1Y3nlSLfq88NP2fIDm6gQWT+
ta24f9Pen1N+KSBiskJtJOC8yOdG3KLVHazQjPeERzkgde7PxvMHhos/kkoc+yTt
xBFQbmSsyFYq8jr7JJBEKYCuoNLV+kVAVIyvYxHjytEMg3R5EDhZbnT7hXUJzVDi
jxOAFcaRoKK8QKDJXN0bA0zxbQOL3LqMLBkPGNj5CeSP6nG1leFqjBicTzJwbJYq
zJmToBT3yyV1Ogw4bcijdgJP0DJMCsGzZDDJavZi81J3m3UeF2h5aVMuZ/uxgBKG
aGKMRejSUYqe20SCju4hrmoHpnbiq8x6MMGI3sfmGDJHORyheO35o5T/fxDDuFza
ReIYDMO43CqG9NiYBjQmD0CL/2AMv9+7QYDY7TfSwwaEaNEs38tdNFxjKotIdFJ+
ycY6d832rvGS4Ecf5Sl0+FOjFGKfxpkaH0OfRaH8dqHrFQHv+8Z+faxClcyenNZ1
031YPCsXGAR+SUh4PbBkLtaHZfrPevBSe2L0UPsUeEvga/7qKSFb42fRJfrCHpO+
kdu1p6h3c/vT+P8+CoX7c//EleYpk5TVnSNl5w8pWEZvJvj8V6cTw8thnuJgyYwo
cTnW+a825LSgOVyQZQCfV2NeavE5EUhu8dLpNZQgO4hlhStVk7U7qLsWwbZYFL5j
+jB1xxxY0M3rsTzgu/hdh6WHEzOXzgSteDYSc7ZmSEXvMLxh3PHrC4A0FZbaclZD
On9PokmAr2glQ36z1skmZsvB/Zp0aoGNl11Z5/1qsEB3RLTQKWPdt3pZaEDvuGSm
+vhiEaQAUjUO2suxFqnqoD1ajFpMIKntCwoFmzQ31Ih8tFcgYLMM0onqZD1W8GmX
ZcKY1jIs3fpM00AikbzQ14DZbjkGU9Zl7Ndsc4HEJEiuCNqHKCxnDmrGP5s4TB4K
hHxGwEchaj9wu0TghKSllhH+KzeJqkrfh594L9fEa26PUHWwyYtOP47ireqHpAs2
pfSOW55+OCxADeQVLIQekkAbp5wl/ZqFn4S5jSSBUIqdxBo3JR8uTPbqFvAmnN/c
f/BAGZ73HJ5UQQYM7iwiUIwVHNY3idZDbA8PGmna7VuZ5qMJAs+63lPXcHjKmy4B
NyRiY/xAbXWSAtERmmNJPmpuvSlhD0097Z9r/Q2IksgYbU0iwMPIKSjs2MUL7ykk
uNQMHsZIWPSxJo5z4w3G/A5N1is7ngP2xD1WodliyGxTKYz6QGMC42DYR2vUUydM
C0qdlAennlboNaJCSBkuW2HNLS5qcrHgHGHuj+yZEE9BH0YVlle1qKFf5rHSeFK5
4UWstG7sArLGiIMlGkam1982uLF3JlOpBIFWBqboZ0EBYuntyqThsNj4Rvqi7v6D
34y4EqW1lL2Ufg2X4llYOfH9pDLkcFGp2+ZIAu4XXF+A2w7lPgsKdxu7wEZf6F+T
vtF9cFP/BZRKNR63vMBuHKBu1QjMToKrFkx15lczgr6k84ScGYTedPr1N2XF+t7a
yQwUTQLo77vdhugQJmpvppHjTC7aAzJUXUB7535KUYH0JOh05+MvyRslT+MyrldO
fAz7eLPCgLKcniiwfl+nJWGTe7Ah0/6zaZk8dtjkPYGzpYZJqlbZOJ0quhG++bK1
X+mYVUNk+26SsQJwIZXCg1G7x+vw54pdFcWbraAwoDxHL59QxL3oaONE9RQJDOxf
gJBCdvUJXtGpVLUZqXdHBk9GYkZqwmDNfBJMmOho1emGU0wHq6PHpxeEksZWegY4
pbJ+9BMaSHDZXkmRt/SKe5t9yoe/31h0Dt4+XgbuW8askDAXEuhjuF68oPZgl5NW
971bQZX0YE3sEOAAmJ4TFSA3GhGWzLC/8l8z3ZrdS5FvSp7COqxeGEUT0ozZJPww
ZuKyug7MHoLMT2VuM5U9wrwcePj56Dzn2bHbB+uJmn93fPrwG23knAIxC0XGq1UM
8kcxYyWtk6B+Yjm9SGMNdY8fEndHepbbh7x6WA4eBNSNA0SD/hWLBr1SAj8ScIcS
2Z41L0y0CY7t02BenyX0rkqwVMgOVJGsQ50ImqYFfQXt70NScVFc8pYNHX96ialX
ZZnrkpfronFFzhlEmGRqSfbDyKB2sczMwwUCWgTYjI00+vPwfNVpy0ntn7hxUDDY
PsJnjuCHOAVTGL7LoTZB1Gc1a8oTNVu/jJdsM9sy5vePBd6rl/fg+Gvo5mXt1GAo
h9azMnnVQnJiyg0yG7JHmzAYhGMGJxXBotaGwbNHz9T2sCqxXKwu+OaAlgHpckog
9iYbE7fXjuNzq5SFb2uodGB746UliQdPqeu7/6iN//hGdCjHKtdHu9OkK33rJ2L4
cj3zVgcOY5NL0jMFXWHgCJu7e5Vgi+x+7QUJiJV+PrzW55+jGAKwWAVckRL/16k2
a+5IXfW2gsWQfRYlEDxsHPa9f8xjqJ0BNwzPulZIQ2Q7ApT9CBo+nzc+3mvzXFTs
IVvG6wJhAD8BiHRCsRWBsd59nkMott83gIgSKM0v3tsV/ft4yJsZw4aiM3OxEfnY
tQWfMDt5hWkEBwcI2ZfVqONSpgnqIOglGjKQqnoAga5xUSBwIOY0hePxOJFTPVQE
XjLHWvlQRJw9cg12Kqj4Fyl0KmlqxBt4aL9p1dnfSH7bLOoRcJzIpGGvjzr4ZDam
UoHVF/kxO9PDsJm3RRzMglBnoISDyM0hnswO2BdbLxO8tkLteJaONYgx2LFz4pY6
IEGtHZLUl/X3wRFZ0IMmUtSdDQ8AyXauQjWjy4iImJCGwu1ShEk0oCw+ofe1uBrJ
dTlQ9lr9mhiUQccs1iOnTw+WCsRCEj0JUs4ppsbd+tQU/mBeJAKJlCGK8hToL5sv
TyUgNmwMwmFjRY6VdHS47ebZZ0mpQ9INoxDLIkekfUTQeFq2FT0KTtcRdJ4w0OGR
9oO9vkUhNaCzvql6oKiarWCXCwHB3Drt9moRhzhDpxyjqiZRf42QH9HaLDW/Z8eA
ZZb5XyoNyajoN+8caQRdQRxCwxDuxNQv7DrEoCbmvODRcqisQqBppWtZtTdIe9MK
uIL20mxMpAHjl0ygFA32jLu1d6kFpjWtQfwbYB8oT+IZkb3MfdUKVOBy6HteHnfl
fCqC2IP6OLFK7+JEpMJ9SVcGJKBumMcNWzo15zVvkUsMBLiPdiXWyHXiSTXhoy+j
xnlIlRgkDFGNGGA1VOAbnKqjEeEjhAZZ4LQJodrKugcFLIWFi9qfMprys6s1Kv4C
vMhdvxwCZ15FCJTrg2LnpeSkiIs6AA5G50KbXIdslkUcLxbRQzGffdzO7sYggAcJ
O83a/8bpI0L6cygCHMIwGXuhL4QywHbhT14r+uWfKQnWQVMs0ub//G9p8Yrdq+Mk
1hr0vytoZVEAu9WHgzgtbL+Rhq+4aCPH3VlCBKwRHq14bZozcdo+rBA5e9t16OUx
NNGBNqYPOFlarQZly6SRf0yVQ2/WjJTNqdclpzRG0PUmtznLwSjEj/b2v8QatUnu
8yQdWkowMpEmPk7gAKDP/ZQnVb5tKFvUP2UtunTrLQlcWgByPcDybKaHxfJ1seha
UiX2qeJPiZTcYbrG68A1i+DMBwyJXmbEkufAnhrUjzo5jn1ACpL8rg2xdiyqbhAt
DAuaNDES1dRDLMui5pO2rB2Kwep37k/WMJopDQSSOtYF8Ly22cbMdOU5lWibNmmP
mx8BoidypUescr20Ipnvm5pxdUhXlyJ2vZHwiEu83EYp8n3gACOTW7JroDslO/L9
Tw4Q9sSPFOU6UiEh4yXtd/ui3v4BONXdqwwz6A4p9Xt0X4QfheePBUckQD0fzbDz
GdGPoKJISTklKKXQw2FqgQswLv6Cw6DGMKbHsS6sTW5Wq3u4+KRMzH4cGkhTa2oD
BeRXsB//l54kpLQhFuvpqxnyVPN8ymtb8S0nxUuMDf1r4TZaa9pJg8XivDctQRA4
EmZp9teb+kF1d4n6S9bCp7gnNJrmeczadSU7nxKuYYWdwreSdUcL4NGcul0Sq+Qn
rCetEusiT0yoSg3fp0USzhkEBcaQns1P/x7ELIHbUxnge05bYebA1y/u82gRU2Va
qsMRw1qjzO2AgvqfCCXihR2j+o9tEj1UD+q4hdl5038TxQhVzFdtMWYrvBfJjOMe
Avx4PkYsD6Bn3EHxCdH+sVJwxuj9dF1PGFEVulj2/ZZH9jpWaVPeFm18QbUQnltp
4q+ZUTVrVJD306MUAab+3jMUlJAyn4IfBFd0Fg9/dbWmQZR1ZbVyrAYqVAPg2CKm
/pSwKS0ceAn4pXRZvcX5e55O00wS/s39jbX5AVWsyt1W/JXr9vHJ2PeJHCCKermq
TLHh588LcfyJGPP/dghC4uUPx9p838gXMYa0MdVsOkoI+kmeov2JohLuq2qZ65XN
ESKknTjLGsXv/uHFfkGeVB7dseQvty9mFk+TCZu+NsT9v9ri02vSnXKJW3vXPkeF
sRcePMC3SrWYYwsvF0hkiUd7axNLJ9knMWhqYVUcbQxPV9vRc4W4rHbpZjUAqnO3
rTzLMwpUoA8Jgk6rRaZUL4W3vETGGyO0rY34dcQJatdkQ6eVre8OqO2CciG9Fn2b
gzGRO4Q1LmLK9RR4K9rL3z/glMM+kv4S8EJdFXzi+Gq9CM8zz8FPry5FgENJnL8F
HXBcvPcGyS/fhE6UQwXwGygxpiVVSoih/ndc310wqwURIQoRt351TruOu3068zVo
iTMxGju6Qbk5fy5NVsQZUCYZq4fBOPRswps/EcxSfMq73olYafMKRGeGCuX+aDbU
ar8itlEIWwXcsv6J66tSIjk6XDNs3XYDr4w9UHMyFaD5/0ZcqjsgQgMWXn1ovGKe
bFGnOZkx6o0JB+uPHWi7tzipUoOhzOW6Zote17jd/kRePH1ClEVoy0l3xF2OV97T
KAHgukiI40Jec3Yc//VTwTLXk9EX8W0s4zf5Li3D67lIyJjvnXSxROusjm9oViFl
x8Q37RClGcgs2See//uxT2wpzZ4dQSRqUJYVd+H3Df2WwdsY/VCLE03Zixsazxxy
y9qEnqWPPW4I910rL0CmIfQspK9Ifjqi+OrMM8PvEP2ZXkt25UCUdRbI65W2MsBh
LqHvMoNYdj9HiVaDzfx1Tn0A+q246JtKF9evMlKbTxc+XEtJAAk6siU25RszltNN
If7bKRpN5RTf2VaNL/kgUXlBVZwO9f2CfVxAiQ0eDxUZXpuT4P0IvKbrHMbDttDR
MQdMjyONm8yXlq6ZN6n22Xm0P9db3h7bxirMNEkbaY9DGknXAD/Ax64poJa8kxh+
1V4R9uKxEBe+rknkpgAfSJ18P3kAU2NoQBVcJzIq0YrTKFmoni9dKdSW4XF0KkJD
6KuM8vci1XKxSLMez0xT8+6Y3y2OhffJFfqi8PyFEtPRd7i9nsFDxwp5+uN3d0vF
SjskaE1iEPMKwvOYT2WOxcjexB1TK0sMEfOXt0QgacLNsX0s1jdvSwbcu3SxkYvx
RKbiXDrk/3y4p79wKkcckDLQUhK1sU0DrdxJHUcvRtZVl1sbrXg+NowOeeW1wvgp
tN/+fNRUNSHlF73pTvHc3MynByx4QI0wxW8BOEXKlk/7bY+8UD5Hc+m1GC+fUgfC
IpL63h97kD2z3iAgegVSEigVhNUZb6zLCan/agP5Xst+31jA2Ubn4zy2+2SNCVml
vmfB2mMHggT3mFstFmoOwCNl7wDalhgJIQLH2u71k1MQ6ISJmj7iWxn1coHRR+K6
4u11SCKw2CXfkkwJ7bboW7gJ3+gPIDk0v0hdcEa8Ek79JDj7sg5/Mj2M93zEET13
aKBy00YizbhbpjiW939e9s18FdcPNwO1BphCEzWP3XP1Is+zGn036ZGVCXFCqsoC
qfMsHZ4uYIX9ltwE36GUIzG7cpAmyAkH4xaF+u0FqNYYYTE3iziK83C5/MB39cu8
vrypElfpZmzQz7h6I6boGk4y0ARwWhpqwFEfJD+aEpEaHElGm+WTKZJM8JIyycnp
qXeqllHqsFiLtIVnnL90H7o1yYBhFvdLwI8XR3M72IkeyKOK7LAbN7q6j1aQgqIS
5ksD4Tcbushr/Ez4DyG70RAZGPf1TLGWoYW1BWcSIeYf+FYsn38kzvXN6NWx+dhi
7rT7WKZo6+1euWG0nHzEx0wjbCBOmEDWy9hWHTDj4vDUYpKC5dR4pG1JS3zPm36L
T/1e98Fov8YBkiebUgT/b7QhjJgs99IqD8B2xl/+rrLTkpbZJQu/eJGECiq2v0xy
/ifry+NvsI789yfL+YJs9SSh3qXOdVMIacnFBSOMdbLDbvje1tvAUmUA9yBVtuAe
xCmMwwmeZVuURITsiq2+u+kzPTk6wVg8WcfsuD9/bc8DAcK1hcefbBjBzYRvItb4
wt7T1jHg8c5YuQZHnwtmny17N2TINn6qMR33FP6YZvfYwQWBxnazYvL/R83S/Fre
EsRNcbexV1PF+9Wofa23iOFw9NBzt7RXlFuerr6tAkHECVl2Q5mTXg9rcAyQ9Vn8
kQiUs64kILLuBWPunfn0+a0KZvn0RyNbD/7Hmbr9S6WzKxIsDS1o78pNlz+5R06I
0CnI32fJaY3xYb7LF4XFz6BxJEfhYEMG6V7E5uzK0YlT6Li66V9m3gVtXY/3gGbO
4pMxZGZDMbm5vE3IvdkSDZAWZSn3ipzREsfV7ahdTZyP75DhYkR97t6Ai8jnKDQA
kPvtmsX4o6cIrt/kjjFxZMIPKZ5YrfkeGDpjNckQc0nA86quKP23mgvtlWXPuAB6
I2WfFdTBhJWMDCAveML8C6ZY68UpDIM4YTHMLzVJFWLKmQOigUu0CyiJfEg26ip4
QlJAO+1uES1crVXyl42QKmxScuBeDhmEb0avnAOgPdzZO2iV+oB2cEPC/DLfxAU2
0dwuPO0gtVpP0A0mz17lnvOOIpMNurTLiXTUCEbJ4UnzP4MHbRzwWmcgkFh90xtw
5CNcrWxJvSZhck8oa53OoZoIYA5zGEfBmOoBfZRlAe9E+xKy5l6aGIx4ypug7Sa9
rlJeHX4n18O3MzRPlH53P7QWdps2rPovSyh2cwt7WbEeMAa9sfO7DAUVlh3Kkj3Q
XiddkhZTznN1xctMNlzhO9DGiT7Jj877HmrgbPyYsGgd6zbmQQ7CBtoMbvrai/y1
qmyWB2t8X4fKG4ViijcqBUpM8ZEd9B14fXCC8DrH/mAvUBAQkOAgc1qba1cs1Ypd
4Vv1z7QEA5z8PLhlyFCFMG5IyB0dutEdFdo9E2ThDbHdBbfKt4H1w0lAejpo1peo
s9aytLGkW2d8xtymbUPqb5LoC74GOmh3MTKJ1uTrxs+mtSkLau2DmotiFISTXxmu
u3m+R5576lcHWRf9HE5+85h/cXiWg2ev8I6NNrA8wR/ykTXRwAKq7PHcRu5VX5e3
yc1L/Wc2xXjJMmGxiE8tF7Nefm7hX79s1zfTQGKZUN3DY1T76koDxVi8/tWJPZMe
In5mXLYToOmITWUBQ/TTYecmqhUgrOHDCkjCA6ylixcL3l14/InnsuW+/hLfGXqX
Lw5UdsiyEL4QrpUf7RGDvYgiagT4zclCLrYOAbIwZxHI8hXY7T0gVP31DBmLzP/q
23tiqArUUjTZZqx6XoIYFZydVub+Mhy3gs9NTHIkgzq60vWMUF82u6kCCNiw8OyJ
wxP5QiC9xd66U+U9d4aGWUtKGFVfNMHyWSUhEBTA9C17T1L2nPZZTOigWtr7XsNE
BzGxD7AXYH2nbotfY+fIxgKnwgsUspXqNKWtRMliaOE6DnIbrmv5bQnXKq3Y285z
qqZg8E/jmU0cKm2UfFD5fYwfvceeuXYNjP2okWupNTa5CZoQxHyJh1SFaaCIlbx5
3JRypDjeCwz2ECx4BL1tbWP2YNhv1vvHD28ZZdo3a2XXKQVkJGjAYdbivTAqlrDy
XKFbHDvrJf7ZqISIzcoanggbviFEPxhAnu3nyvmfsoOGvzHyIUoCIUnG/J5JXQOF
Z6VCaT9NLgIXOBr7Xu0Sq7gdN9ozHyt3iGXJ8FerxRCeeT5nrRuWJiGsk3FaX62a
3u9zS/r5vYgGd8MqIuQ8X88G3YTUdqMvAwxiWr8Nr6wg0pmkRYfkX7yBeUGZJbl6
G3E0tMbIqC/ATRwM3riBiCQB+v1UtAP4z1OxrSxdnlcLpNLw5Tym2u8f1dS9+fHx
nNv9Bl68Zg/d2AsfMPwyDAOBM9i1iAGDaKoLCSNKHPgyN8Ftzv9A4RjKaKEfrWzE
wPsrqLvNKFCo11hYINUA1piWQNB7syLMllys2Utt4IRnE79Z/+78bdV9fxXm6Wzc
LY4beX0V0tsaRX3E13oXOsBj5gPm+UX1dXRcJGDlEYoHsTDhcr3v8ekk1mVbbvl2
6mJKHwSsUG/7IchFAWWQg1xDUlI0jYmCMxjU+mricQ23aTyS4W72q4vlt99VwfCx
npwsIBKNT4kc47bgT9Uwt3mSbVoo3WZL2/XRPckc7OqLRNG6X8naZDlmzq2kj1lg
uMNEPasiHJ8BCIO/RHk2YHj4Y3cobsqhVVFvNOsxXB85IJ5D2FLuzjDJE7rL3g9i
KXTjS88ywfAR5XcbCSasYO1ScLVM0q8tx+b2IrQ+KGuRxtRWVmBay/Cwep1Um7Ir
dbkOvPsFtmFNsGZek20lmZ4/B794PFvM7JFdr03Qe/0IkchXwGcMFV7y/FnS08L3
+DuBaA62yDOB1GosX6iacM1XNHs1lnxnFtTcCxwpOndVzze5m97TkHb/kGpULfzq
Hai9jRWtZb+WD8ci+VTaFzKVP5qGiLPxrR1xaPXnefZVccFSf+JAA84dKgt+II8P
EOOfd5cFd0ncPaNd6L+WCwXfjWP72peKkGykBJ1o1hP8Oa/niFibZ56kY9D7ibcL
c1gprHu0K2a12d2SDv4m1N4LKlod0Nt2pdVi3F92wV53VC7ckREin0ocQ/PBLVVI
b8XIFW1VLoeCynPX1v4SgJfQzs/AzPg/Z8Y4yELTF3bpL/BKJfx6Mn3dOf23qv/E
EoO6mqE9zD0dfyxTQmHwYO++/TtiN/mYAZA5my97GAEqCIF+HUiE9GhzJqOBtG/t
c18LZACDRknDkKf4V7Fn8Q5dnHoCAcYYfY8hTjH6k11beNsYGHeaQ+fzc5hOtdUF
aZsr9BY3PqAkeTkRLth9sOSlOakXRvw2jocLgDZBQ56qRLcnOVNDyx2MjPTDrWev
YgUJCyd1je3G9QoTMXb4WiBbEqBxrd0y5qAjNOyWQFvNl7qPl4+RKhLc0WFw/8AO
VD/OczCMc04SJ3KN5PkxbyT1PB+q5vXIeoohLN9UWG3isRCT3bzzWKdbP58x5UD+
hMktJVhIBkvVx4kDsQQ4CHwECAo4l/C5ikk8QTy7aSTRNbiS8azrVo6IX/bOo/Wj
SkPWR4xk2SaO7hacOYTNI7hU2v8gfswlLjR5aqZ2V6guoGNMvEtqhFHWg4lw3ENP
Ck1MM7CQHjvqEpSLRI/IDgsVex0cE3WpUMWIvwdDSU/eDggUtlKrPygHlsBEDjR4
cpbvkZfG1reeFfpXALXsZC3yeoeRL26HKzVQlcnJ7JrdpJJw1YLO81nH64t0QmS2
2yQXgsI9htkjmtIN4eNK/FjEj0D3qtR61jlTm11Or+XNYSJ9GOurznbiCu2Jwf5f
OtT1Qkh2k0+HMSEUKAVVUws58ZPGw4hYnkkalBSQJboBJQygszIhKwYs7J+0NMHi
yrE2PG7xThEzZuFpilzbb4wF3SjfUkYgG5YOQIBmMqfZWWHVb1VDcZoaOttnJFdP
cLup2md8dxYFby1/FFHZwAuBf2cSzu8lUEH/80lONJ/KuL6U1/AGYcS/HIlnx2pN
Ht8z0UVHq/VTA93P0pS/Sx+v+Wip8cImTtZvwd1uFrPtUXB0gnpHKltDABIadeu8
/2xdCtPDz0aJhiqTUcediFgsPxUfm6afCOLyCRCSHoqKeWLapbIYgzoU/d6da6yu
y6hykmBGpmdHE0ZHDab8TFaGEgYwygXrRnFlJEgUtVlmLiAdsrp9uQyzPsht43Cr
HpmJ66fBpiL88rjqislhslBU8EugdkPRP/5vg52bgd3sezzLahbGGM8jEeBBBeB/
NJfPzCS60MeVeHlkRVY7/Crg3MmvXqjTOBD0fQDwNwxb8O6VtJ6J67JGl1siTzbg
S1U0JT76lGwOQqHpw94/7eCf0MNVLpgQANTL/LM22BtAk3fnCCtv+c9hcCXC1468
UFsnCwkl0ZdWAfQS1rESZt5T2WAEN1O0UsZeEt4PYAQbhB1WMtnaX68C/Aq4NnZ2
DBcA5SCF8iK7/icnFA3XeBzk9sFzJ6PALjwrC7xjY8VirkJW1527Y9k2cal0SX52
H0xA3zOJdaKkl+cKsKtrxsxNsBAfrrFWovO1DFJqdCJKuP4nQv/N/OOA2ZTrNE+H
X2HALcz7aMf4COfx6bR/9S7+dzCqY6/84WPGLwv1D8iE/utVRYLVyPJ45FcBzklT
nPX1sBnmdm4q2PyYTjsPgelvPV3F3NVrW6tAcFLIYY5i9fgwKMAxXPV5+StMOEET
52IzcORtFplJwY2a200Hm+cUvQzOOxtHCx2FNgKOsbhIsS3STmen4ujD9152j/uW
O93hbiWPngoh2io8XEU037szaOw0pPeEJkS/QHSLHMuxbfn1cO+Vl0NrjbhU5qES
e/QhINuY5zAgIE6QOJ/ZFXiG6EnF7KBFgxtUhMMNeA2mxjsk75KX6i8gvX80ky+h
SUNaBXDKtMHMXAZUHt7ew5cT9HDH38s7KDYi70s3r5pgkUp1Ob6nO/dYSsGXwSev
0KsLTI+lLaqCCM6TyFFCCmT9wLOKff4PYVqngScDc/Rju9Q30zAecScKaViNtN0f
CYurWUlaTsWhpuY/KwY8l/E9bXbejlV5p7Vf5hMPlfN4gXQ0+IZK55vOlGhOu6tk
KlneA69LAD3wQ9Ay4epedeBtkxqPhcPNHZqRsUNNO9MZ6Pl9KYwPBKsQaKOdu7I7
KUVOY9HzRSGGJMr8tc+RH72Tuh+MFEsz9p8JRTIQhXOLXMUmebGpfCSDJL8PQZ+p
FNsKxqJGzfIoVFBtBrGNmspvGJb06aT8lF2V4vUX/QBxRUvIAR8hMADgaV6dbWdu
arpZ5qETtF+QNAGZZE+YGYzvRCaCnjW/bIJDMKN1wKMIlxYvYXTdPBiuIHrr/IKn
alPiq5LnprnDJ9iD5GDt6/pPa4rHwmfXnw5M5v7q1Y5DQAEcspReisFjhIgiZucx
+gzMB9vM7MomONK48D+2F+Z+YNOIcZPQjeJbFcSQiSz380kd49zfSXQ6J9wDn3PH
MKIQYzWO2TN7qJ9CqpmSHVTpjOU5eyancO68jmeT2bNribIX+oRWELIV9MQIU//C
/PZNTwuVRqtafu5whvrLvpLDufs1BxIM+BCKyHmDF/ezU/++165CHc1taBroiEMw
rnIESDLv6JewClfybFl1YOC19QYjpGog5uX30lhK0Mr3tG0801Gz1lvqVMsqjZG5
SFT7h/EU21kcJl7IbWoRZE+o9x3MaCzGOY4t6PE5QGMwysVwaQKK8u7z/ZQYa0jm
pEbweirOO/oIMG48Fz2dXrtUtVJ8XKyCCMeU1Vmpf6LE9K7an5nOYu/BBPkDsVFl
gnhcabMYh+M+V/GJ5stoN6l9ps6TzQDfduFt1mRoGTxAbTzZ+9Ci4p7wMorjqq+K
zi9ZGjILJarNFzf3503ViOEQY8cGG4rLFNCEosQUmYamTbbqpHX9V1XcuHpl6UO4
QOikrjwirW0DDDz0QX0BfCzvUR/0yhL/R3hEfQySo9SEKMeRCgKABsnhxabJy6XV
Fv78STqt3t7FrtH7orGGEGRxQ4CLN0sNQrKDpewU4hUWAj4hwcWJoVAJ6ccYDoE4
PXL+obVj/pqCaaeVTm4YValLJDk092bkeCnIhXV/DZfoKsGFw1I7QWTpyrnOkzFs
Fme7ugzxEoWwwFKHWc5KP2gO8vWzf1Ge/QyjbAPsiSU0L0cWyFL9Q0MJgf7RqBTV
PDmdgQH6RByTbmSrVFW2SVcfoHPWLxsAiL054PS4BjPh7EXn9vrtL3m4bO/gHjnw
x+TxOCHVxdy2NFWEVyBcKvAPJp6NEP3z7bMZhtUptKxw2dl5nqVnatydh0AnkgXh
jnzoEakMfopgzMeHqjeqFzo06rCFsNeXKzMusiGDrZ07EHk2YGNN7jI326mdNidc
EKjNcH5JTGtC+FmNi2tSw4RgFG2DwzUbsgY7YjhJ/qXvKaeSGHGDjCO7337nlr3W
jtK1/pJVyUwblN7tcUfDVNjGSlOVOF0OHBXWp4qZTMZJjH1qiCFbTttTFi1wVTAn
PSiNzBbh0rBZ5LVdzrOIFi86bbgVy38c7mMZOwuJaxIwP3qAGdfDAoJN5YIvGZ/1
c0mml6E++tCzMKxDsXrLfiz75FT5s4ZAHhscHRrbgLbM5XNpX+knkYreQlpxQwAO
PHehZFeD1Qb0jldPxRAqKRxHrvcu4wJCTohO/SUHJpPmFV+x5NjnxZPdV9XXy7tt
beOubSkPZNJK8fu7+jBI4WfzKNTp47oZQidiU/mAk4sEMmKGaA/nuDdFyW37R6gk
hPw+ebMmWcc4hwPvyXvRPcK49CC9q0ioQX7lvCE55wZPJeOOeknwlP9/D117mt25
UjwhRLsvn/M3lZMF4WhPcqsLRiqHgS0K55xhCu5MMtYPr1hUiRvoLQRn+rzpStl+
ELPnOloMNptU3+Cby0JZwv+nShyDZHJ3NekTTsxpEb6enQ9Y/jTDfhFU1t3FWZV/
sUVXkpydwhSQUWOFV0aR4tGjt8FUwIHo6TaeL9aOyEewI7K1JQd3LjRd1NlFUBvm
2w2LWvQ22eAezy5edwiBqn4hIjydIuacNUeVlKIxgMrhyISUKOVIXppKCYK6dZtn
FPUA+UemVl2koBIqSZIMgA2AZIFxn+kftmfLJhLHm4irq5NPID+5g90tAbcFxPpH
d2exN4GMfL77IL0o3FT8KeCMuGDB4UoxryQUrC9I0a8/m44k9iyHI29RevssqX6N
q6F0KrU5C24MyrW51nk0VG3wgx1Su0N0cmd40Jnl/Jj4UyILz2kzw4aNqM5luDW7
9r+7BBRFXQyoCfR2+ghIh74zbsia8GJUfNnETZOx2/wsG+fVc2aSsEaPL7+Sce8I
3ri7otGJZ2lZgR3ylCpkK1qR6nEwKDAsAcR7QaTe0qX46+OlhybOPR0rDOGK3vu0
hGrAGZNjsYi+HkIDb5gtUOp3ljP3HvLpZi4XE4dqYy8noV2UZV8yF3oEqm6c+jxd
tbhCg/QwiPFGk+f7z9xMs2L4M/aX5SS8hDJlc5cpZZTflOiheHH2U6sIjjlyUiM8
PDKUk6EwP7OfgEXgbXRMON0YqNtH5WHcVsF0dqYM8aatMgBmB8eRAJQpPlq2yBkH
mKtO2gHYy4ZyhNk5ckIJadg5/+sktSVnNwI4hJhWO3P54KkRpmlWFZ5qqB4uGBtK
81mZgJDLc8Gei9L8LIOCfaV7n//vd2Xx/AA3bqg7HQcn7TjCn93G1/AsUxuyYj7c
QrOK09XOGGIJ/X3IUHHVGx1R4jFEg6H3Clz3pyocFibUT8A4TBdF2FrgASh/eaPK
Pwyb2iJKBKE5XvCX7Ci1bVQVDBjDPKu+bi73SbVjlPwaMerTTWRg+Ffjlo1cNtb9
RIDAAN8ntL20efxqPPE0WlmK5Na263pUZc5k5tUztKk1fyyv5yQIeTzeglqMIlEF
anRxDX+ed4TXr2WChzXUfEjhVVIhU1VbFcnFdHHT/KpnCumwEVOTOqPX38tqTKMJ
nq76cyiFKTTET0kieFxix14FQCEhssmMR5S9+hEKX4NqKBuFaLFUyLgFYQq4NKtJ
+mZ2BKjCKz0ra2aaRVTXc2OyQCzv0U8Ll0XeGkOK+nzpbwnLHkbE3gnkp6o/dXF6
gO0khIXS8pBWHn3DReZQvtLEN3zsK2icPp8MyFJEpSbTmmPCHDwnDeS9DKLBlTJ0
jTXoAwZ6Ls875l0esWIMph3H3as0FsPuGLH06lGAs/plewCbs3Wkmw2744y2NL8M
3tXBnz55H6VBwgneGR7A1KC2nW2akZOmlSLOdAN3bzaGH9ex1kwNHGL1e4MC8Twh
hepfAvtB5mnok4xAn4wODluTQeFbFnnbWxu4xvb7D84GIxldO/ux3xJWIK16DmZF
DnUhikkCus4O/h/ciLc6sijQmgcERLJNMJNrnPMqEKdGp4rdGtIrE+rzAN+NYCvN
PPshgLAYSKR5BKDqRM6tHGYDm0YtKh2CDP5jxh3c/SjKGUuJkBLsXZJGWJHfWykr
tgcs4EaQOJHJg8WGQ0tqi63PD6cwcRxLybUhfXkjEVhEjjKUqigSvHvyAVhlLD4a
Sn0ORiRve/HYXYMxjgF0jc84PN4Jb0NSl++R4gqSiUVNuX2cf7tC4CASLrSrHqLh
J6DwL22PPDM0O6QsL7n03ROaoATeALKA0fuTLASA6nxSRQakVj3XrS/W63ICAYgd
vVhsg4l8hqgJFtYxhplXTwOjQSsD+4u2El2femw1wo2gUdjnqFLsCf6qHBL0nV/L
wrmxnTkCiiUVnstezVgNUKOto9bdV2pdbK7/Zzy29K2EAAeBeeyCyaWboLA+vlKG
b8HGdvb502VbYiIlfn6LrmcHzDkWlZFuWENyAk0LVjwcSp7UIpNsTwW9ufqLBuaJ
rgDIJq9OCZbHfPewIQwDXwqiL57IOTv5it5eEIcNpSY4Uv10X9MoiF2HShjz/u4V
oF6VzOJ5krOt+Yl4/b8g5eMwyBfFIxLU/3pCfMZDHVRMoPyxqwpj+N7qWhD4gUb4
9cv3zMUg9aNatzld3dfUQ1HE4XTb1H5dt8SgWneqEh3b+pcm2I/qjPkNIQeqXAsl
UC1gRkrDOvURiBagsqK/iKP7LTaFQCyZtEov8RMT59V28EaNemZ2CnNM9+MwNqwD
TnTVEx0pS7qp2KNaBXqRMCbC6fghp9razsABAo/938oZJ7apsTdG2xW2Ao5q1eA3
JB5xAX373h+4ojGHIbHlLN3LsNnNDqG5n9p3Hr7OZkFPUvSBqH1cWuydoQLI4MZT
OHBfK4xDU1THr2hHQZwYENVetCY8MYrYBAZU8iWkqCe1stpXSaPmNw3J9kqMhQae
pZL0v2ZKenShBLTaMNKYkC9eY1ZuhhsD+vefNrF2flR4y4yFXEHAupjeVaNZbae+
xYoNkD4BkrG+W0k6D9jlE0WBfqoDrJESmqc6d2kykGsCKiNZrYfRCV6GDjXWnvA0
GgPzjIHa4dSJus4kQithC2k+7BTIUO4PDIEJ21mKNAUQw9Ekk7ZNy5Pz3E8eH53J
StdQq4VmpZz7qHJc9P1LrtbzuueMHTzkL1b57qFsGqe3O43LygevecP7n9eA3dKY
4rp5HtT7nJ6Dn+NO4icZ7qAGXopjz3v7MF3GigxtHezaqfJvQJeOGZRsNZgN8cet
8+l1xNIzc6lSms2nHj3Ga775IYcKzzFHm2DMMQOoR4bjQZw641gvm5spZu4ZIjMy
/gz5wFuO9mloccmU7iRpRebvQrz49kI8o16nbGl7Sa4IysvTIXOgACYBYrhQywYk
NGq43Z37kxw++ruVXFwBioutix5rLfZ82gzPFnVsf2Yja685mORjCZok94bixlzd
zLu5VJq3VAPWZt0Ie0NIMEkF/OVm0cqYYiSmQqzJSTRGA3M/daNQwb1roQmsnckl
Of2bbDGpEgxrtuAB+Nr/JdR54vvWtlIfvVkuFXdHGk88lwVbJWAL/XcZEd1NrCk+
/v3/uoHVMj12rXWsNUgUgvybAWqj6guiH4Pm/ZS7rBU/tgniyyyCCs5Z8QGMlRZw
9jSwY8PEhxU3rPXN+/e0HcHVWo/zohXaA6v9fDr0C3PIzi9JNEARc370rguyH3wB
Y+VMlgTPpauEozab7WitFRc6s1zRnvnxPoTXFy1zfgmTGDsywemlsy7ewz64gQL5
G0EcVSWPXwxpwU8EbgUdw4bbzW83i4IQBVjUTeXzP19WeVmr5gAh8+oOXqXMiQMI
eCkJzO2niDPtRbR+TGyxHax9eF6L7IMq9DMGUzublOk7TkOJEvLaS6pKAdMgMjCN
OhrUHPtxIe6prZj6Sc1BJEuF3LTEWJLgCU1q/JThVjkAHJ+xybjXKZ0YOeKA4SFY
RbexHuxvU44ua/5V5hCVFkjzBMwipSBtVC4zZ4qhhLR71Lh2lX7EFMwZ4ZvwiJQY
Nf/9OuU0sJvy2VdPkeVH5Z40eZcOW2IRA67N5wTurxiwO1SI2vQNsi1nfI0Fc4cY
fCa7mNT6E1kNvWfq2/P7LkWD6VX0cy2o0o24FM7GUgxtY5mhJoIYsvrIPiQrOAs5
F2DECEWpDrDmJtctlxSqHuVBIpQQHMUNsU5+zVqdlbOF0Ig48Ppb0GzrfTtBxtlK
Db3MMQq4FKPYWsQP58TXN+V+N6yYtTepCmLUZ2NyQaK/QyfCam52Ttl5zmgBXNiD
OjhQgrtnSDrBJIMFgaREWliDehn1cn0jjO7TYPwi60BTW2NJIAVJt9cZ03WdKWzy
EbUUxe2vPKYwDZno4SeO6qClCk5DKagIMd+5XarsavfBByemCLQGZuzEzifRRyr3
pSlCoZruZh9PT8VvzardkBZPDLUv4QSRqALff8bVHxXm/ZBV7hoHko//f5uLrrSi
dSNBXfropVVJ/Ca9sfSY/jY7hi2pfqcMqBgK3B3jb3dbKmIFeQ0lBhxkgTx5xP1w
L2SuuKKqhQUFOJ3fvSOO9ZgYOUZUYnJYd0wwm83RmpmZJnY6Tv3y5yqb/L9qrH5S
Hz/dBgPeRaeq9O/8fsRspX33z5t/MWu1ZXPaHdldh220Ai4ydsXBB9lUOSp11chA
cihi/jrQ4VPv6Skz4tcEmwPJeylAjbkzVI/LIr6xT9NJe1umih89W48YgxAuwSx6
aAmnCqkuAwkatIi1b4IZ0vmId3kTarqjRhBoDlvdva5tB60dkrZYIaM+ifgb1f3H
xwp4lWeZindcvWwWk6Vy+60hoJn6PLMU/cSDnVzpSbdYK2DURLxIgxNu27Q22PNS
y5o5uRp9BqgYwer1gPPymEPATT2hp+d0dRqLNu4eukCWOw3IXGc4yu33NcOgZH4z
Xnl9SifF2nF1jWwYEtb6xgrPxfY4I1nz2EkdRc8bip/MmE8DyjVODVpMEg1fSDYZ
a1Ogwxbb2JchtdrtyYR+b92nCzCEQbqfh2dAmJ3xXBLD0f8iXqi2YM+bqSP6OB87
A/YtEMDpCVcMe3E+A1bGHG9PU9DMcL+o+3epzM1kW1EyDJ4/VVKqctl/7Btl/R5W
0oC7Mpd9noZY3zB+MfCY0Y1BTX0VASatNGG3PpKrV+65S3YhhDJRcWRFgWssaDwL
wkxjjg9DbsYVoXRUEfEOAB/R/AdpzqTC18+aiRrSn5TxxOqRz4NzGahT2rNJN4Iz
TE9QNnKRuyOWRZXs7OSjyYFM2O8S9BfpVW7/ip7U5x3tpDoe67Bzsy5wjP0Tivlu
4s1lIKTCK8GqAjWvVhu3Sv80H6PE04d5YoCuP7VCTQzzBLswzKZCgY1pzx3uK1VE
r4lzYHSkuFC+Zu0h+RcCIxlP5D6nElLhBq5XSs/vNlUOiaq/MST2PJWQgV27kigb
JHE+0MO7vvax8C1Xdi72NbgAE5bP1jF8Y852T8Yc2tB7cdyNE1b8ZLLLLqOOXsgI
eMEWPgvc/khbWecB2KL6VmTWwf6m0h4Cxp4qrALvU2YVu/MR7cUdM69mJq91iUdQ
PkzdPUG4PRKGxlH9qQZNba8yqFGrruMTxDgkW29HZeTTQ28MeBUEukxt102SMCdC
SdFxvoUgbULd7fAzSL7Pzgv6+NfduVxGfKbCnnr1xcw/GNaN4jNZipa+K5iWhCrB
bDotvkQg/zY8RPtjkjnPqEJPVeYTj2bc3j/P/CJ5qrfFRSPNngOEIuHV3JTNmFhD
xfEPauwpB5C/MDT7SM8fpe2QHrIZffxpjp8Zvmka9bVOIZdNQc/17cw9Sb9SO2lP
mXuL18d4Bb98r6FmHbwjFmFZXGIVb8S7rW9PQD9YUFX+7FxHTUzjF3BWaKNq1NU4
N7Wsrt7GeWIjeFv/jo3B6Bk5EdLV7Z1YI6KWmsTTufcbcCJLbGdPBxAK/4nKGrt1
wOtIbvSLFWnfbzdstxWIM8nsADfW2bkmOEnZadTThY09OHMZ+8COQP8UNQarYYfG
+T3JmnETFfpHw/E+zVXthMpqwgiKTupPaK4J05j3wfif5DIh+OKu0b8S22iJtvwW
wmWrOemXfQD2kPk7Ju2E+84EiUiTAF9yfbPhodURb7rdOWflHX/t1ZpiHaQCPVCp
tR/YyewU4h1w3mGe7lIjW6Xj6cZ1hf2rpc5s7tkklZOqNc5FkAv8sorkxRqm6M+6
AQ7/sAKrNPb2YTBMAQsJ2JMfX8zJC/8yOOc4C4sVKQ+piHPlvQjHp/Nfn59EFTn6
sX/d2Zprr0XBERMTF1Ii6XymvDwiIp0jgOdOt+oNb4b7qk0lcZR8HxTpzgDH5V/8
X8N3Y1JRRJsiGAJHJIs3t1rw6zMkcaLBC0Fxv8ZLKt2J6giADgd0R6P2T8wLlqZE
2uz60XX7MG0SZHkGlAyJJo0Y43U0HxdobnnwjUYZBSqV0aVgjLgMsb/kb1qxdfX/
LAEHb3OBa4JC2/GgxJeMnP2WF2OZwSELrBRymrfm1ohoebQMSYCmKV+PsHz+xhtS
0gAGP6aLSTXtCEsOYdgGtxvjV7z6P4CEKMuhQ7d7nxKzjmIExTV+Gepw1PQDsm1D
QRipfRIm0VLeQGaqfkr+3NzCL4/b7etNSnRqc9KaG/J0P+qYJc8nyTds4uuHFlN9
k3UMrMq0l6utW9CDFZoTzA/WjibrzL34W3wgEFw770sCsGJltLy6Otjp1+0SZWO7
J/mTubZbPtHx46Y6uHhQB0YZMYcX14ydzHIWyJ26tZb5YiUvOlJIW+ShLO0ZGYnu
Kz52D6++qjnJrvDq5jkBA8wcQgOLd/2y078KDBS2IzV7gSummQ3481PXafVvZapq
Jamnwpy4j4gewizN5qkIdKrYeWicQdLFLaoIgGan13PmR9Ec5fa4/LorlLkgPmY2
L4GKZh/yHxVxMXF/WTLBfx6dy+KE1v2p3r8HqKDe739UzOIXEEZbn9K/k3nMB1bG
Dxuy6+UVMdjUQXBmDo5klXFZogvUGlf1HSFeEc3w3j345id//Bf9Qkp0H4jjd/9G
Oh0faPMqP9yuqoYN/QA4Lkt+o5VUyQuPK+eP5UDddRAR10HvO56RgRTmOEXOfjQM
NCuW6YfdB7hzyHpkYYGHjRs8u9651Yq2N2hdgB2oQ1o9oplQz/FThdxx/2xi+Tng
MbVqOe70VSFDTrwqzjYs1alEfvreMsOcu4WCAiCxw4NhNHuYHAOnFNnbHr9EoOzq
F8pbOLdv/AmUAjrEdccypcJgkpmG9Eq/PtgTu7Mn3lkojLug4lV5+oPYXikpD/94
Y5/7D94/s+5ZA2tCqFlJTdeBcmRkvd6rWZRwzYTiuPuHzIGd0UehpXuIZ3/G/Ulg
qKZHDqquqBVQjNBYjlrNUCXo2Hp0vIt/qb7Uf03AtMHE6OgNEUPCXDnplNZtRFTM
oL8/iYCZxnsmIkE28Hxnq+XGhxwPmyg1AIC9WG7H96Tcp+1kOZIAAm0TGBOmMacy
27mDnoMmRrq5WnVy9Z6WV4EWb/sbm2X3ef67YABnOEyZxj6ATzEzyCNwLmgNbte1
kbJ8mba6/p5nDjvVYRBdQsGCt609J96i8UTMFFGiq4UBxedcepBb6IYGm1amyBqx
TeD9c37VFJsGI9dmZxeCEBwknV0y92Y3w3x1YJgXQw4aGhnI4r8IGtQjN5id895G
eSVN3z/uGFQQa9hwNtWAUkfgINosjXZQ6ME4vqgJlvi/d6336OjloGdmWcW/Suur
IXry/iZ6mbNXKTODvMk0/zcA1+BxniRGTORxi90ZO6WF7iAJ2AhHtBNp9i5cBtnG
PPbJaVzuGXkrTwARqBMQx0NM1LiINOVUrFTINsix/vcbiC9U18eJWcs6Lx3P7YrO
Y6JXMYZe4uP2w/ZGF5hZxxFl9EFW5W8uvvizIt/uSfZs7WYZorP64RyeCMhKWNzd
pT8xbvZ3ffFSRhOSNrrjaXk3XUdp2g2MZbXpCEnXE5460jEH+UYTloTVCSPkXkaz
rf4LkSLgEuUuVU/8Zmt/xSuIJOAOlXSxX1FQhXA9p+zUFHAq5+6vHtX3RlMJWNwF
e6/WSwacBv/U3NnOERzwyavKvhkhAYfbjhfoOy9AVJvg6H50kpmeskG4qATBPCaE
WtpXIE1X599ebaiLlun/YIe6/PcvoT20mwch93t4mpwfAiTLUY6K2q4GTYzdUXTI
gCCWIfOJvaHbqtwDKoqIzNwzoEItL1q3IquLVgKjoMCTRZoPHwqy9VtIljqK5wBq
MCNK4e54y+nDsNahynLElBvWDA78gS+1q5yQ1Q+0awecZYSZ4WBDMeTYzBX+G//c
Li/DY1qe4Vb2Dlf63RRvL0hwQbgRkxOwxCz6+m6q/fM9oxRBXo3GINA1loH6ZWLj
iXTht3sQBYu+f8Sqy/F2rF6lqD6h+CnYIm9b4yi/OlJgeBkAiyJ3XRtfvjUQk05n
mHm+Fe0jTUY4kPcXfAOeoH1ilNDoyk/POjS06lafH3x5UKN4cNo/PmxAh8PvSZi8
Pmy7Tg3tVl1qBDrm7OOHEE0wVlltdvi8VQc7QXOX9qbrcdv2Q3tUbSmplsQqJbv1
A8BFnyVe2izBqjrb8fblQ3QLC/nqk9DfW8NM7miH6uisKP3RkTSjrLpW9NRFxscY
sthOLDkJn3BJHhWhqpKWYcI85KhAWUbscQeQ9KqRE2/NRku3+iIohVXstZfISZvU
RnDpqzDQ5P7kB4cDss39FvBXkxRmqMMtS2W1H8Y/pXuzK2QPQAvizh2BJAlwR0Bp
tvgUNPcfeEYOkNJnFzBSq7z+1MlOqbuJizjScDuW+dasZDQaWnTbeUC7T2eZTL83
XOoks5nH2SNxVqhEtSTkQtL/Q+V8n3CPrNg79ir9drpvLR3YemmfCjlMwPpArZ1b
Wyrs2nFaYiKlMOCAxeZy7XQJSN5fML/1/0s/vR/MeOyBLuDWqcvEYCcZr3VvshiX
1pjfhplv9ri5QROPsl6e2fe68ou6KlOqiHssxUblW3nfz7NmBQK/AtYg0m++Jioq
qpI1pfGmwq/wzu5ClQ57pjdOfQ53qQaQtJjXbm1UjnfUEvVhrMWsDhO+Fn3bL5UX
AiTzYfarKbAwUxkAnRsZCJ5AP7Uo2MR2PygWHk8r46GfvCr8uev6WYEX4Pqj7yjD
inmeK9LfF7qdMioRH7zHzaMhbQkOZe+N2DTZWZGI6sTG8EnTrbiv3jzGP85CjdSq
dSYlfNkdtZtp6Ce2jtsXlUcjym59VI67sZxtSbfDZoFiB6xr4w/SSrFeOTz350Ya
zPxLaVABNaH2AwxzHBHdCLcYqiLxtUzt9ws3nLdERLHiqFrO49fgWKVBAXyUdstx
A95N/3S5k+2LllmHdh2PF6kIPVfT+V9l9ZtsgxvTH8vmEs4tqsUlDpTQoqcnZtLM
7R0Nr8hojI3628zKDZ5c/6qbvrQTU1C/6jv6VO8wsMthFBL8jXCQOdKCIVAm0oY3
xnLPbMqwWFaaPC9/aN4evkyANAu5nSffQkyn02BB6o+I1nO+3bAZ3cW5PfniTzvl
bD8U1YiSdcXnFexvaCDe8BYFFdUJ4um5oIgN7SimuZ3nKM9OtMo/OyJaPm7jm9kB
DPOlsC8aXaK7GA1bqboh7blV/63Kz1Uii/H7Lho9WroVmApTXgoL4tkekwu46fuI
Ohg/3paxCxvQRYE6mN9uaG1qvMr8jH/bHNvDu7+0sEwICUtMMcAsl6YRyoTnFi+u
0LaMOSdTylIUJXQqYfJ4/eJn+6XMLW4fSy88VbtWNwbiHlfPJTnGS5Lw1Zm1FiMa
ypU6k/yOSXJkY5JOvMu0QCw/AiCoRWJ/mJ0kDqosaz7w1Gzk5KRo4xMTmroEJ+Sz
C+XEZKuz8NcaP00j1WxcfMh+e2IhOTzvrM9hiyYKicIL+uGfdvh1CkxqbIT2HUqw
HLNhmpl3GG0voodaWxU7MxR+kc5OpDYQIIvck1OgTLOuxMVFejLcybbtVQK4JnQQ
kqlsF8bbqPM4dCa9M9aMmq7WW069BZAGO4CwgpevP2ZIr1JGMchFgFu5gPznbhB5
8+spEm6nwR7+/V2KvbXx47+XAqTGBChSJufGxu5MpOm8YWv+ZpANB/mRbnPn5mY9
/szCqRmp9Ml5vxZacICoDfwXwEuuvI2fF8PvWwQx5Z59MxOieTZmLHxBnSxFbogD
qRhG/ZcaNFtejXKzFvrE8+nSZSel+E4hcHlO+b2/6CKQWlBMLIcOWpBCdtmqDFMv
VkGrKJca2rSgMGBOOk7T1NIrC66RbmIsSSvR6JK/LFuh1gxXRqBhKgpIY1kCrUt+
8ImrN1dX/yZI1w+KWayQXu6EfbvONaj6igutBsJnq10m8oi8/TRaPEw0hD7SBaB9
qsHM5K8gm2W3m7Q+MHK9I0HUJy/gzyHjPjVAA/lqxsKQ03XaReLBw4icZ74xB66l
968BludEHd46wtaTxpcXIM/iy4OlowMrghzQylxly81UZ0nbr1sGlkCziFpHFxTS
2dox0u9z/T/EGrK5vHKUUjkt92GehEzMWdFKwsnP+4UbkCnUy6RrRuVlnQxGdNmG
3p3exTF6EQmO85HmRO+SdMv/yafDcyU4FEezrehUPyp/OrFoTe5RdG1JpfPOlfN8
YytwIT/KNoyimr/kn9tKMCU6+WKeiYL/2MIs/gUXAHluB2AcAK9UtYQ4MODG9ZYN
5OuJZuWnpygVMUcL1cExD4Jc1eZmEVOQZkDjvgu47hvKjVXYS/WOSH80CgnjXBVn
JCm40TkMTDZJsiX+CcP+fqG2mIVA5wrMEcR6RI2CdvMrif8Y8qgR5VtaatiVlvH+
kkvg9kuVekFhELPfTk5UTlHntaexyO+2OCq1mOT3dN6San0sVXsAAwC2QHYs7rwW
PZBCuhf3EhShFeZXCettynAsZK4x3SHrNqZNXW74K1qHVQR9fdKcGDvuhcLU0fdy
ASTdo577PAiA0Dw+LlfBjqqvblBc4u2lWUQIqPd4P0VlFfyVK4BFRXEJpeki3S/9
GFmZthBxMBHMchizqHoF1vUweYNSEpZBE6DhSQ1b4nkD0RqOxW/DYpAYiuU8BGAV
quGrtoJBy8szX3OBjkcIwmrFC6ga43DZhaj+OMmghiBE1lyO/Ou5uOkiXktIXNng
QvS6ajrjK9036zy6TTPZc3Ji17/UB74rVWG0iI46hjlqrSwmgoe7SCFZmBoEcHRp
Z9/DD8KZtMdQl+/iIF4SAHT9o7V4/pKaOtIGHWwI4n0raqKWbU0Mx14wFcxgrmzp
FleagtHcBD7puCyauwVilqHJAm/gBJ/aqvRnAKXBrCYupDp6DzbO3yVgRYItMezH
Xf3U/gricibk/uNfGQKQdEpO64SKjnMOeXjZ/PyrNwa8JmFW5JvEv3ocYhnlZPqI
y69yCmCArgLxDFyR10NanaFCCPtsHEBRVgA09RDjB66IUTbmOxwDwqgKhetcesNx
s9UJDJQS9w30txpP9OHg90Zwssvy6DPFT2k/3T6WNuMkkImhcuqZNMGEcUq+DlUc
tDSRrJbLdHS8sr0EPb1vsSTsbaXbIFaZXe35bXPdNiT+Uw8Pc4pU8H9uj1T0iNYR
/qLVHy9QL4bUj4PAvG20YxmLF/y6Ag7/S423M7KTnQaZKC6S45zoUQLm58396SBQ
qvoIwhrFUbhH3I6f63ZkRJhmU9AAvIYUTrHGkZZWTnzTg1QMMWRB5OMHdH+fsiDO
YwRdz1i1TNU7sgkwUhuEHB1EkzZw950qEzHwxfhgwMkIewIw54VHuPnfbGBUMLOE
BblKCnF5BDqJoLf5n6ztb6K6gOPmem1Rcml42uYx/7PNYrbZMoxRzbzRFLRdv/tQ
QfDtYYl9LqPWs1QhgP7fsETxGvuM8yibzvVXMZKivSZ6vdjqBDIdwd86JJg3jEZA
etqGmfou5SqiIE16MH/Y5r9tS9Yd3UNK2LGoOkWQ5DW894Q0G4VoThGedAkqSDMY
TOBpkdhtvdUYurTLuSqWCON7AA7lBLLuiB6LLCvmxM25Tt0iTFVZpNgMdi8niowl
jQWEClYXe03anJL+qiKAMR3gcLGcehQzmFQD38fai/Ix845hqbp4E9ime0WnLc1r
k1ioCzj5ZAeZtKfwpD0RHS41lmbw9yDTcPKE9evcnMV3JR2BKoG1nOgVIYABN2F1
ISF3s7pmJLmhddvI1yVkseSTc56S9pN4TsNN6IG2LDs4fojy9FOuvE1grx9EcRK7
Y4TVl6oqWLhBhYGYwVCCbMA7ZZOdka9IMM2MjjEbLCeFFrJ6Si4EF2nWuUWWv9XL
g8RVkY4RPAjMksDDY+uNOFBOQZfEAw38zyewqlW+aOmzE+AUwJyberFGz22Z9Y2H
CaoR/V0w/xMEr7etkETtmQogSGTNKHXZIVmFxGUH1O3zm4tdASmOxNBmZGCPTCye
vkp9mvo33qSIwyIPd+ylCVpnKhnCdjvDUriNbHOpxzAzSxa0ovAsaZEEE+FJnHab
fhr/t3kaYOUzxbnhtIQ5Lsf7XPkF5Lb6Wd1iY+t2jBle4jz9XS+TxuplkT8YoYGV
MxaEMzoSDJz7A0IwZfO9zzPZyBb6gZY2ZHrq1N4I2HrJJG9N7bxxOWsuYKuWMYhx
ejxViAzTvVnNA1xuKBkemoDfmIs0NQAuEZ/6fbQ4fuQkjLMUXJqJrSQfm9mUtH2N
hGiWypDvxbDUdAvukRhcl2MI31ZuiPN06NrmFXPLJBdLhQmfB7TiCbl3T5KBkBIc
ruklc7bDMh19FtTQx4idhFdrwNjsRkw9xb/8/x/rWPkF8B0imNNtrzMOM82riAy0
zBxbY9+2yYJy6BDaEQs+DnCVDEihJWOnc9LBEhuoJZsoO/B7VKx0U3R+DHf/qqiB
bXb9lQVWP8r6bmmEzjV9ZJBoefsv1F6XB16QC9RH5cas6MK8g75fCADC+J9UnSfB
Fvps89FUxHoD+nDV51ZUtCwbL7UEEqHQNWk4b/eRpevYOpSh8rxSu40cNizWlMcC
tB2e69w9Knbg8uroOAHVgkfErXV8dfFRAQ4uI28Ef76+juihZy0s0NIvBD3xvwEk
3p74qh/nyPjj1A5Z0PrXYsVESBLF4Xtt5GAQDKFQpzZFPX6zoqqtl0Nb85IMeJqi
ll9/pb4l1tGubY4OBMAMTXtizQ+asy70WpKycxHM8uPxIPK9t7UIW60m5G5r1tKR
jd6sAb7mL5C0tUHw8rkMd8OSoJwMjV1x6aIH+of9AdK0BUudkETA+aYmk1p8PYJh
pThk0q/CaAKxvaavWtta/vjle3960T0Gc2ECGvcOQgEtYsAsmf+wHUTa/bhXfyTb
1UpgbalMeEidUgHKDxbobGNKs87GIQodfRGn6toq5WgpERjDo59Abgowpk/2SlPq
dxlTMCzY3Y0bTfRzMFg1qKQpo6z8XcdT0Ab4s7w7PkG3IBYFvs8WwfzDjQsJHZR2
6pLLxSj8CmOx0/M4Yyn/MTG2lla23fXK0jY4JuIDOvIb5JsUetmWA/2B3ynqlNY/
vtX3BJ6fxT4/XHHri33hWwiAOlNfu/juwimCj6U+qCEA1qWcFDRSw3uPg2URyr5H
ajwWR6vUDG/ygoJnnsEfvMbuFb2tcpwH6KqWP6rM19xg7I6nD4gNzr03tW+VQfsu
MUpRNBVwyT0bEtI4I0ooBiIar4at230EIbtbkwk/cpKgSJzw5zZ2dJ10DtjN5Xb6
aKQDtwwnXWLCDM4igu0liejBE2d95DZpA4icFskpMO8AZ3uG/nFaW1tblEbmWEGg
H3jnuWLLXiC9Tit6MhYCl5XcwD1RPtPd/MkyD8PcM8aT3cOwOIuGWyjHBaYFPSRN
kZ9tSUMDfKKxpAys3hanL/UBav7dONGJHu3pJlHQQhX5fR8UMSgGgSS5PdiR5wy1
G7KS7CIkVRdyqnG4Z7LlZwviW+RtlL+q+uomhr7HSfn8n19Z+hxVIs6w8hx1NTkZ
xwgzPYLP2g9AtwC4620ldXxIfjYShpPeBCqM3YpN0+piMwnujEzIISY106sk/yqk
TgGPt6lGXTy75Xr+TYziKPOBpjQnq7u8Q4t+/RAvttc9iy1Qs59++BJ1+gRQonKc
rXeb0V2Vl/0Q1GNWrxVIG54ysTg3rCaKkGdaE+zI4xAFMOP/QH/1wA5A6X0Knat3
KK9M/bOonAduug4zlF3qNgi9JdSy1ubQrUNO8eCAbRXXXBqJGpMBrybyoRmgoHdq
ew0wnAIDopuit9UNz94TKkCRoYkVAWQdf5fbBF57PwJcc6Ih6oTR5LzY5xuNkokz
ueYd67yfIrGtbgpUdM7LzL5ODWCaVcvNP/CTqqy3ZIW3Cqo02DcZMUbmsWFBWtfj
DXhG3aCzfIxwgYXZXWGWYXqzlSl22bd2fGH6EU7QAREOKSCeh5YBV+Cu1+z3UTCz
Bkh97K1k0CvWoywsW8O2cmhZp5EwK4o95hyqr7wHv0yR05JuZHuxmGmh6n/pWjEn
s3jzhPG1ehrDpB/ex2sggxz/ifKGfiZ4nnk2W5P4KmV0vsEgnFgBbzzIhZUqWDz3
CQN+GsgMkOtj+RQ9e1sMCc8Izg5A5xlU2HtOatoPX9kvWHz/Ig04lYbpMe0a+bvr
cwxGBP9xXWRIA6CGHJSJVOYOFE6yQ4QDicvfeEaIODX1v9P28lL9x0fNFB+iEdiL
Un8BI3LQr+tszaH+VK6ycQpEmlbjTglyQAw2dQv0azz6oMwePM57eg7mtOHnq0NE
Kx88+itlvxXMqeM5D66jUtKEsRu9IdNAdGLtQZ4/svYyTcy+6UPhSDmx1XAR7/yr
3Cozz+67ujzgg7+alWt5uIygqwLGn6STlzFtH4O+6DmYVV5tOEAxUe8+gVSHOvec
UjPM5wTTigmk/3HBj/N6OALsA7crdJ+fz9JxMASDVqgCiTLLI6+ur0hiOBvw/wCX
kLcPVc1Y4pwyPTd+9dsKDxi2Zj5A9nLR9iFUhhBXB2uFlQWzCmiV+hoHv8nQRo/0
fYapeG4Wljp440QQ5UwcSa27ffAFaPMqXuJYe7ARRx/wnSBmCHY9rmlh727gbcyc
M6TRy4zuUC1VCQDwso9Dx41BhYm8pG+PSn6SBHUF8h7MMWHjpUfqtyMgQ2z4ACYO
wX0e0QPme2bwzQEAr9Q4N0myZoPJjClClc8Jj6ZqoCRvwdd+0fDW0hJa0uvtbLeB
WRDfxPLIN/5sHpX09sRVJ6JK6+ah1fvLv1AI9X5uOQkA27rd84P3Y9XKHdLfs4k9
IIl0d/hpmOfvahZQ6vyJ0OI5s5TDnsKLyJ2XpMCZkty7xLU6wnI5VfBmj4tiILY3
xDNjxbcPxrpucMWmD+DGaKyQF9S9LYCW2tnxyN5gOoLrCoBYzCEcUIiUrLI04pR7
7lYFtni+Yd2eAGE0mcokkffYQzFspOGd59AMUycC5z0qyPeTb3wnQMnwnGzHHxyH
7+r6NQD2G4ENWf2pkgY3e2ii9TKsZjqu6/FvXSi4s0cnNRC6NMIb3XQmzRBAimlY
w50YHEjfUCOXIfVUdA8dNwNL62ZDkVSbgmnZbhxbn6qiMt6ENIaFSE3Pofjr5w2L
au5t8FY41HcOZ+jWXOoa2I3ROb5Fu3emejd6AXmgnkteibohwFyOSq/5qBKYeMD/
yzIotA7s6Uix9oeM5pcaKaQynLe0GwqRsSmqfxgQWlvGSWRGMvbv4B5AUVigQGBt
7WwffGLkfLHbCGqDPcQ177zS7iWMnCUUySJdU6++Jit/2JD91RkeC7xhbTfMQmB2
Joeqx1PtJ/YjfxsH38SOtn2dVDkQs6a4oy4vgFyqUP3Mx+OueOfuGWdfvDPVUVyt
eUo/sneMiurRLSrAF5AzEQazztfvMzNH3CPS0nwmcc2yS7YQTR8hffhX9ay1eI2G
1NraqxC9jCqGQooEjdypX0VB5nio141naVq5pXpc5sjnMmIjqsPCNn+iEA2jmh1p
+dOcnczqgc57jV6ntoH1lWIOw/CHMUGLMu36CobBRg7+U3/uMfkytfI6WogkTg1Q
gl0Fh82XE5aNNrBPAUBCb7Bbcs/Pe6zA8FWy9B1a+GNoc1ZLc0vcrQ68FniWCUMM
E9NjiUFvpNcTcmmJRfSqMorA5lZrLeg+XI2wywIAhvBmtmVamLQUgAu6l9xnAYrQ
yiOgQxu0u99/B0puHg5dCFzs/13ugsgZ23f9jIXahMBdDHR3agS4Xgh8LODBtRIF
t2wlGDW8vM4GWyWJZQjuafUahVukKCMFgEOlIjn1CLeUkYoBbXyQD94e5R/fuLM0
GGgw3as8nWwdygLVgcC++DQhZ7ELSC7nv2bkbUqTomobW4mFuo6JAQfYPoOnnvFb
fzxu0zlbmI3Qz3ig6UvzgPuCbqNqBI6ikpFzieZy2967rhYQSFgeO7dwGmkYrgTP
/6TkNGdK+cpKUifvgwQgWSQcpuAR1kQKIi/hr8E8wEikIk1Dmk0EnKLwOuY8nSY2
7uFHJh+4/xmjBivoyVe0pmvUUtxaY/FKmS2j9FJBixMNTEbp8PXMUdRuLxngx/77
LOW2QEeqm+PjeqRqdc2h6YdZi1cckRc4xloyGx1hjC4g2kGVKNc8C/aY+0OGbW88
4uq1GZEbjTLKdhw2RhGK4IuAqljJx9veNotD8mwkPcp5D3F7NGCC0MM9SX8IRPCc
qPvXSFGGmsM6DXmmvU4Gu/C2sYm0X0Rx+N+364zk6gnLJ1IKaQsAcbJ2vdr5f2y+
owZnMJu0kCQ3n907q453TH8ULvYFSP2aUZk84u/ptpNOUmQnVHH1doChU6qnlddP
cVE2R3Lf3IC7GYBSMQv9363ONWfGB5ApqNFSfFc5lTsN9uhX3qMhEoyus20gNtIE
zQUW8VUpACDHz0mT1Oeu5HhTJ3zuZOPMrq017fBDL1dOyHOHgXgwFre6C8oBXUkN
oYpx+iY01sLyR1GjJnv/uP4uzjfOoTKN3bNj2tW0ZUSE0znGIqxWIDtlMFDaJQk9
pF5KuUo94e7Nd1ipRejL0qqqyHLi2BSMPnXuOu2irYkuUN+PxFUQTiiSQhZptgGT
oz6Oksw3yJ58xUaDTz0r7mcCMB1nM6LRSknljbKn8RRl3F18Ezwj56bwawfQKj17
Lljc8EXu2/IkXdzuAn0NNc8ca8+9DUwCIh4FJg0OIZLCy5ssUDQYcnfjTq3oWyRz
F/6MkSvyFCEJBerb/9NWoACPdakDqdU5+j4wKNdDxn/0Nq9NK/KG4rGCSTT/mVvX
5wUppJoGeh5nrH6EA3oNBYAJcJtFHAEN3+11epGYLP43qO9R0Nli3fETBxI7q3yY
FzdHDtm/n0OS/waDiyLib4giXuEavmZkOmPMIBRiE54066/nRDjtudtzHsMCTqiQ
ZgMHCGfoUFLg6y0ZIAU7ufMGICeOrvifsOag/xF+/Vo7q3zkZTdA7G7XdS2l9zJy
NM9QoBKZ+uORVmxkYedn9IFcL8xvBVBYYR5xv9W97b7w7eLpo7k56CHi1rfJy70d
EBN6JYNBPgg3UmmdYlwHyNrBv1Nx6vINtrMcFgL1+CCRCKe4G01JKb/KYjUP/qwO
a7luvvRa+GhW8QPPFdviYK5l1jvSNl4jSGm7OnwfSqDNRbE5BVd8R/YEcgE5xATI
UGfXMuKY171Z2qC5vNlc7j2RNGFxinlsEPuS1WcOK9yZRSUuPxsOk3QNf2HcZwBB
CkMfNPSE2OGu0mCvQ3D0CxSzjqETe3OXQcb313uvvuoVbXeRhCj+18Sr08OhWK6D
6h0lIGmqlJmiQOughn1K0AFZj6yGzOuHbdgRvHXyLzTP0Xho0ymuHZs+kBufL3FU
zZDd8zEh1kmNZbxcSHuZvSDIYD6gb5a9po2SZ5ZsFi4931gARzWgnkx5nAlq8Oxg
a+TfpCnGLt0Q5KbfxpbiHsNnt8Yog4fcSCQGFuaXhHE3bGzYWzjXUrT2WYl4RZpu
Czt1I3MSKcorK7BHiSUQgYCNA1EjMjYGHmO6Bj5uTN95CsUk+wIQvtJ8m0naalkn
+VQ8KmStUJR2QRwLySWtUPbXFjIgn/dijweqPPC1wgQEatLo6dQtMCIG73IQwpSt
1jW35vBuYd/9yFBs/DvCygNvd/kMsYRIVciJX7IumQu+R0tBefkziHmGMvfxG6vm
4+mh7uZaRj9qQcDFkLwPgS6FyO95obA+VTryj8jc9qxZta9YieMqPZgetYBdTcei
xQ4PlhvrnewfqQjKsXP5AebI1WsEQdEc75qqJed7pShPawGPEWNY1P4kOmsMR89V
s0PnQ67IaZjDXPEaFH342zHmiYa1MAr9Hd0wpn63X8bGQCtjNbA2s/QIpRQmCB/t
6/Qv2aLXFrMSdH6i/JtUwGeAIS4ufViSi9c4AZ1wsdn/7iYgU4795zcNRnfczJFk
obwpLG5m3ptELnx+5SwnLFJpTiSWIinXo2Xw8eTYZSTxdVfJKLefY7Fbp5yafMw6
Zi8WzTHNMtlC3rqTnDf6nSWrZGrcSRw3Z6xRuqLXQbS6+xBeQYEtbj7buSCzGjbV
dl7kStSjzaHIDLrXw2weEq4Jkkzuy6T+LKJnGU8CngHbdrlDNhnZku0esVfFnfN3
VkAkM+mJ7NcGvIx4mKVUDFx4Uxc6quDFU2hbbqxsJihF7iqBwpqq1C6QmJBKwx95
Kqgv2EoNr20fEICPgG5/J9TckWO/PuuI8rfGF2YwOpcqKPThJbqcXRdxsVYgjQgM
8OtHaEZHItuZJbBjIzEcHt7k0RYVczUhyYYU7WqyFD0NaTYTIb2i8YQasxf2LZFc
BEqdjBAVdaMB2IdI2hg+vh7WruZbChmVlBGurBQr9Qr8Ys6WBKcaiWIyFj+bY+LR
qN4AIpNCMDPM0pjdRZgw0rQSsXJXymrzC1pzQKxOD+Yj0+nxreTWnJ/ukN0Gq6Fw
b9YYYPhnbrKFzcodFHaJ27Q9Mvff1EJ4wZ1L0z+91llK+Cdn+re0m77JnOOiKRVX
nYXtVQuUYxOzrpoYmHb/eMFCI9MLno+JQVsoWm3WacAohZLRdvWe50pCPGWajpYx
9UhKCtrd1HacZ2m8tcpOStyF1jJfxdFx0thJTXa1znJX2T6XPOT2B2BpjC5DvkC7
2t6CADAclm2eDkEoV+Z8t7Vn0m/uHVNr9MS+kgYsA1J0gV8wKxBePTWQc5zAqYRE
RoufKUA0jUsD93RGDZhNb26+yY5ufUzQnMJ9KenZJ6YDOSc1b2SEQpBwvo6+w+uq
e6HCthy8VMMlbujKfyFnl2g/UEZ73MIWvJZJFg7+YWFQGMXTGgHbocUHanVZ/10i
+STrBFRTJDkCPEmG+AXv034eDPx3RB9OYZjlwF49ST2AMd62MGOtamMWv2Nul4qM
/ytyL3xPLTgA/n828SUsIVX3cOyrD1kTBq1UuVAdhElB1+35QT8PEJSB10/BM2V/
h6n/KBwP2eYYyYvE1mIgbi/JjOD94gNgynYibprZz/yWlOdsEEpJ/iWJiPN8KYw8
bnfWElLyr2w4sCa0E/CL3BJD5AvTEMXd2dQOLkLKzx9a66fSC9Ni8ej+JJwyFQHz
BRj3d6UJOsVcjqtAlfxGrGQ/wURj4+zbfcpSmDDfTro6fECgVvmEqi74vNJRrtu2
1Mbsirs0TtWBYfOS1gqFKuvOgIhCftcZXrcQWNELXDI2aHy4n+dCVRksphPIKA47
KLbF6a50h9vfixIpdEe40G6O2+QFCHQK5yng9pvnImQMp1DLLrCLIWk0zdjWMCRm
c5wfGZ8XdwC9xSdQCN9Mf2vUX1VO7cuG53JX7e5Z5VjlaKVTQtBqUIihtmiKo6LP
m3z3MRsfnGYsjGKkT0o5oOGexHNzMeKwixfYye32mhGeIyDvn4L/gjgFVy4QLcJ0
dMtIdWMfHpajec42GK1z5FMN4RAAhQclbKkVQQIi8UKNqRELkpUJPx3QExnTfoFN
Qv5wuxXfSJJ/FbzuFyc2s1TE5PDl/5unPOEI1rSpglBA7gOs+gm1VHIjv6zdWcIZ
DI4hjbWytzmHmW5FTOuchIIcAjZE652/d2UT4KK29AXt+9J46HUJQFHAQi9j2VGq
0h38or3ZBZgclfiOe98L+NDDf8rb3kXmmQrDgichltH17IbqUqcgLaydi2n8LH4j
MmdWS053sc5RsK1gg3W0gwikBWBWzRCo/5cUxeDGD8eZr8OL0AlWddXdX6+lV/u4
0uKgRyF/xW5pyAeE5T+a3WrOJ+xCnjJWCdG00WhWU6Sk7dHKkf476EXJkEcUqdDA
/tEZeY57yjEVZdGLRpiB2Qxv1yIcpzyo4g6W/5nEG2dBbKk1aHWZVGMK34619uFi
QRd2zllcxhQYKMYXaLm1iAcnL4NrtLAdWkOoF6rtHnbd6YR/uCO9v5yT0oT7gjdX
/C985PgEupzoSyPjI99QUHrkOWRiGkLKwMnksdMrpqA8gJPwrUpr6t9WMx+r+tIp
JfltM1XzkGyqa3k2gjRTU7Afvfl6jnv9RszV4bsuF9fhQ7/vRrVK2xn36wUcuw5q
zI5jhT28fLoEKpiOHgWj5SOCLlQ/f+Oj/2vmm9pLcRCqZoieMdCzeGrBiYnEKtLX
QsJNSh23dJ6OW/CGHaJkJcoH4T51Lzr5ZqXM0Z+afKjAsa3fLlBHvvp4Iund5jhr
BlQF2zYrLUrNjzqGQNtQHfVFF+9tFbPEGwb/PKpulXyY3VRSMiL4wsbCm46dp2Et
EAQA/vUSVqQQbEGgHjlKNuDRSA+hYaVDxfHjE6i99cYx+SZ1m5d6mGetRB6ZmPBq
vapSxWLbIb2mRNZ3+qOVFWVgN29v54JoKx0ng4flEfNk9bF7TuHVbwM86kh0dP8G
1v2SRHL2Djbf7P4pY93VJ9oxiiBenKyrZUeMARdg99mSCZvA1KO252QaqH7AuDJm
PySm2tgpYgY6uYZaLBOQv6UnpQU6Cd6lPdl89h84ZK0y5pfHK3xwVaTqSd3jJ5J6
W296EKeSoP9W7bsY85BSchmJLPSJkZd5uYI4AUz3n5a5ZB/JpIuoipt6E0+FS4AV
3Q1xzBjyRKYXRUxCgmEvGa57wRnbMyas2caWQlpqA8wtXD35JM9AlKQ+N9348en1
cfYMy709478bZYsT9rJrm/emen75RxQNDt4ILT/L+fynVAOaZSKWGL6Ih30U9Lfd
tZPg3mBeIJwpt+L/mJZVhxehknWIGO7Lnqgr8Ki1p6E9HlvDZA9vBj5rtIq4VmuN
P/TjJUg1e6wQ9yZGNRgn2Buu7dmHIbeZXGh6zR6cwz5ynrDHWBefmZskk3A7KG/l
di/zT7kAD8LcK6e2Ms+sHm5BfE4qa1tB77tbnDv484Tl/ur8lK6PdvThhX98Yc6e
eus1WQDcSki6JNOk5UgDp7STFn+6ReVkMXStuC7f/DSW31+pUpQssUg9mGfYTLuq
TsNGkhN21ANnZZ8JYPhW//Fz1zKyU4OSsJgtK1/umbgDxBXU+episWnZQIRNFPjQ
dAvNOTZVW1cuNX9QE2gjuBC4L6qmRdEANDi8hSsOHvDO9xTUAGBgpSXY0NLdV1Sw
LCzi8C6X3hMiGrgcjpF/Z9o7Rlm82SFmLEUi3hHKJQYm9R6bwXqd+IfbtDynFXbD
WCPRjseNZ0+ibRqVGz+4pNioA4AZrdFq2WhYVIvkOI0GbXXORlJSuyJHNIMvp4Ik
TtmSyIY1kIHowjsCQuEkV+S1oyZb9M3U37gZwJ2KSq18vk3nGwnOSSCjfrf6Lq1R
lxoXi/Ea0vr2nAfxIZrsGygb+D4fTF6SI2VYkb5SaRZBHYHPh/QP9Y1rDa6E79hu
2+vpd2vLHjRNVnvNxMyM6/nuDcirkg/YWMnT9B7H2AbCwzEaOw2FcBVRs5HfOTTr
Euop2sc5owKcEnvWGGckkJ/4+EociOCBRU/DQI6fzqgUG9hSoackIe/47Sle9V08
8tpUcF8mZTx8982keXg0OxLlUVq6RdBMAoUJsEKrRl82sTYiTL7suDuCYEqMXhVZ
WLxf+mbAQrIjtFXfGrozJHkaWBgJoy1Sik7LANuBy+G7F/NyLIplVa6eVTjqpXBv
etJiaOc2ctORuA6LjU5aaMAAunK8vjXnBiX9H+44dBQsypesPUdOW1aO7Wyf0t/R
mHsVVmKqUT79X5WwGdE62ZMkeyvxmtaX1ZlFI3jU9xYvdwvG5BK4WIU2J0EjqmFJ
EzC1c67L7jTud8VnBa0cJ1LNoZsUiSqw3RfBPzSyhrVNIotDmBsjLcEXw4SFdmqh
3j1/8InUKEbXAqQme7XDvKDCeu81TNBVQdQSKlorVtCmmGTL5xhVUL0QExIF5aMv
fkNr/dS+Dnzt3ITUW6NVHZJWETLSMTlovpUtyjvE0jmEtH2GTQLV+0o0aK1evAxt
blL0vQAAN1LHZIeQfrFskxeU+NpV00vLK0GENAjPJJrXmEZyu2io6sCnZVALRGBk
CRV36PRhqgO/aFSM84njLTrp5vchtCaB4uUBM+1FMS9hdSZRlKEbNt/OP6rA2nbZ
yE9vjbwqpIKrMDnm3a402073vOq0sEOBILnT2xFnB4pkbHHsxbKOWmbe9wLQTMd+
7y+PK44Ne1b9JR6o0Z/26dYvXXkl53IiJXiNy7rt5WaYMbOLfhdYXhKTUwu890hl
EAXfQzUipb2DAbTTcP3y7E9r5GYuRu3FeW7OOxm7LK6p/aZVXtPjRfEIkP2U/QiR
eGtBPj5YegKBhhCipafaZwaOTeMt9U3kK1taJFOxWT64d1+pjWhi3vNhJvbQXt9Y
GG4eDQzR5/MhTIoH0sNsIuuk9uLOHWDSJRXGmaqlDI8KWf+6MZ/T5x/wfoYgHWaO
UEkg4wVCvRLQ7aGosHTzDlRDt4K0w2i113nWM+lm66knLXYLiwB5WjhY8iMnH1/L
rwn7V1PLkKLkObp3lPgY2OYcbLPRyGYiRhgkEczKh6NDzXYL1uw/T7qlv5uHk6kS
0Bfj/7oUKfhAQiAflUfNLBtn86ycRqIVIqjb3JceYw2qKQLLRSjPkpeSy/6xQWHA
edPnJh2cMUATeurL00Rza6W3T9ldjwUJxJrItEDJG+LwIRYS79mZ7Ml25S6A/9+K
wuI7aJBvmng9pILWiwnCUxhdWb/I0vFIxwwgmIACbR2Evgak2B1XOPrdhBCEYLdl
TmORu1q+v2YYX/VicPaa1OtuUx452fuHfz2eVwdUnYJPmcupR4WcP6I0flmkyOBG
TcYn/Bs+AGPcZBDRdjHdIvtbTNc3p2dwGfMyLadmOv5C6ppal9Z68nNgo/EAqzr4
RIQh1fWfFm2A0+cn1IRsJ/Uqhsl9K5nuY6BF7ae84O5cJbpZ0ThtKWGRvIWYGl48
GYYoDAfdTcVPA0XbQe/vg6ugFwCbC6yAsHmU6ufXDIoUuGTJvK2yQY59P+AImv/g
TjGu5Tx6U2VDNtFVpFeBhEYwRFNYEhxycyEI3sadfd/1FA78VLnsTSX1iC6s6QUh
Ao1Ufc2y7TT0NMdgEejIkr2B6KR7sCe8o8/zpgwyJuj0YUuoJ7sc/QUinYN5m3U7
GWYg4r7OMaDbfC602njfR51hGKKTYvTp/oZd2UItSsKyEoj13IekuEVADbfeAY2a
m1XWuGzCHd48B4qD7d3lEFMh76upfb4uIKxez5ALN1E/Vyg+a+CgsXMgoZoSkugO
cyJ5hdDVe0jdym4vZh5+FUAyVXOEKTo5jUzHxTsknNSqgZGcXiriQjMzd6mmr07I
o6r8/PLONqhaMOhz9+C2XBQLHq0dhyuV/zPbtN6lFqi48mca/OJJKb7NzFjm5Xln
Zb9dFlpuJI+QyCKsKsROrc3UDVY6BASPFisL80OuIXWs0H8iFj1oImrxoYxJXRPC
uoB2cVFdLs8+zKJBRssD1BnzKBOjlvA5Y5a+QidhwU60iINNgHE4ZXOMNGdr+jhS
NhNsSCfAar4im32Zp+7kbItxGKMjx1WhMf5pTGPQHmj3MvXpLVWbd2muP5ML5390
gKDrU84NJEruRFjApDNio/R0RE+LBTQLpGlgs7Jl98Ws2f2jofDmp9QSRpW3Pr2t
+7DlZN45EhmQlGl8U7moibSZIn2Z5z9ULl7dKyE4auZ1c1D2x4Cmr6F3HpJIjif4
u/KMgIyl2flxpxEZC5ZtpAbWiDPODwNQwaSWct9ldqm9W+3YNv6aEuTPIhH0NoSA
Xj6TTES9Vtyji5EqTLHkt3+6YjmOjBrDaJAxHD6iOxKr24VBrNOb/e6/U+BOXh30
ig69BCGhKB8vYfwEFnxHNpD+SZGzicNMpJOVAu+GSXZviTvKbrf1gpJsaGpKX7jp
hDaPT5EKbMgcHW/Pcldd0HCbqsA6a/JZLeKY4GKdAa+35nR8arBSf8lO/YVrjV9S
J5aQxi4kNZtItDb23J46VuX8Ln5XdIgRW0CvNxkRgTQguwlRRWNS5viN7lBABejK
bjf2KHSE6KrVwT33jKVR0bfMLkL/ExowEnWKbM6vHSl7Px960kLRQn0I5MNw2Vm6
ELnMd8xpWBbgn5aNYVfdzTttpsst/ex8Zm/VQnwKIkv+sptjcQhUVoAJ/KkaV5yI
8BCzlIlAJSXu7AUfbmybUAcBrOb6MNlBQ7Qa1jVR62U2XybElwPEnRYulPTaqi24
UPpe7Gq90D3vWyQ3nzz16wTp++as2FwEc/4t1/Q2TwlV1P/u9ntoMEIUZOzVOCmD
ITZ4OLRnyF+NbsYYo3G6dQE7gaO3TnzIxTEWgTLvwxe04hB6XJFEg5K5o0u/igdB
9nI1Ob7k8hNJ4xztk22UZDOHeEUq3auUHO5kdYXegGhB7lpq/JOp/zh6z1RIF6Ek
yIyyeaDa1uN3RKdAXZ8UYxwPOevZJjnIE3QeCTClSnCNZ5zSs6OsI1zBtXxWvmCM
FKti+qZA8fPVrLVJCtpXRn1pwFRs+xYRMzf19kumCIlxwn7VwURCx+eNMQEte5Ex
2dlSTiIEzzJCUw3Yty72JkXzmv7bB/bGHhUi16I+y2udJOdACUkKK15GfZPdN435
rVmwP5LQEn7gRvTXj1Xb7cRmHmi3sgzsY70ywQKSbOXWEJEWgVxJtAuu+40v6kyb
rLcZ4XguZ7+K7bbyBytDDkrHWnTQE+dMyOTi1YynGc/6QdI/c9cQdE0VfspBe3S/
mTx3AvIgJ6KCxCtesZuSEWM5TAD+P71oPXnbiE2Mdj8pcJe9U91C1We189z2vkzn
H2ICLTXtq3PYO2a9VjwgInXXGdr3OsvYth3nbVR/lIrCmdk9HtSatCBZvb8VK2Ap
oRoI24UXh03+fVfDNA+QHYHVM2GtF5JjAOq92KOCOaBsraxW9sXExEj2uNZrPXxy
nchvGfxMIV6/FTsXsHlt4V97Kle7PYwHFiCBFM8vwvfW9gFbeK7htiGGhqIfoDMA
UisyV4cqv272A9SGlt8dPYISl6KhhIVgFQ2E0x5rt91sOLW28gejgSB7dE8b4tYR
2E9IzuID17iQTwc7rIqOaI5cYzDPgY+BlTuhenfyOJFIqJJKdlT6zfN/4JmAoxWK
sRV2eZ56fOCxdIT4N8PnTGpZIkCUCuOhJwCEd/dyAW4DThdHDwyK21FyVr4VKxM5
J4h7F5Xgr1gi1lkwTbUtiWwEnv9mTu2R3GaFfCF/aCUtUJXY2Lk3xk2jmla2CAWe
1m6YzfukNk93Xh0lYiy7UJJDp/KPUHpsP6il3+eFovmQ47jWjzXuEQ0jkfv0jD0j
arht9sAaTUmCFsyjDMNOCrYKO/hZWeF3XYU/moYO/zog1eYZjEhXUa3IbHEXVcDB
iJfywp5PL6z88Qu9gKUL/AH8cYnzlCbRc3DkOobmBSXDcJPxHUTKfoJxO/5ZSwT0
ruLfBIenfP7vmF4OgcjqWeDCPz0i7VSguULsRwxC6zBeBAtOK1b6pCUTBgOzEigK
Y7n+duFplm7Aw3axb3/BHu9JREjJgWd9cMrvroU+ArSYCOBxrqJGbkvu5JBlXPpY
wDjoKdhabfBrlU16PM4eYs5tk6E8BzFSzAGe156UW1P2kkYgFS/Q5sAbfjtvYIWg
YcbQ79j89cW8l3avMw/6uwG2+nZm1dtUhq1u9Y2Hg5vUKGW4TRAmIfzQO5BxDaTK
wgpBxj+kHfcoyUl1YtGw5VaAvosugDiqOa1MOv+TStbeX+8i4XAnQRt66yN60Txs
YPsg1vfmpJs6gfPSyNIlznGXZDP5j1ONI7pqfyrTDL7KfCXvH7adPJm/zNTpYSmm
BxVcBkgVRUZJO7ryznE4lOJD036IFn0MVM82Gc/5pMGMxOS7yemfB4d8Y/Cl2B7n
c+iskYE9ZWSQNP/hIXw7YMZFOBWaCENE7tRxflmHwgExH5ge0rpTnHAxLdYsBqW8
6LfvdE4Up4cbxPTdedd2MCGL93Mw8ixP6LrsiIq2L3znIRvLgdAuS6BPrj7lrPRq
POLRbBJfPk2EsjARuCRNB35lVIfvlTXpuZJ+wJ6fzVVslNxbakfBI9AMTP1nPnPz
Sx/UNw3oJ4fcMJiI/kqm2U8N2sq3YmPk2qVi5QDVoMqkHcT+ZR5hztsqA8eXOVrj
Aw6rmrAj+2rB1Oyu+u79xx6i2sclQquVSWzkN/MwlI5vXOwub28kWcrqY9OsU6L6
0cNVhkZnbR8ph+g3KHYaTqaeXX1F6Q4O87XgoR5dpnIbcMs3ooownFQXruueJIFe
abnuFnlg7qhsg8PWzJnuuiRd3ota9QHPlpk7zT20/QrPOmGS8/SgS2Dv0oWraImP
ISuQWL3uVH4DIC5U+JJR6pClcpUqRNMJvYe8luMT1t2z7FTBTclBKOZEEPGNiLFE
i4zGpodQ7CZSVQYFSicJH9XgGtQW9H85vOhXTPJ1YzYC/MCSg3PqXWK+RefoLe1y
N9oCOAAIxaIsQ2uzYUu3sZDeZUo2Qn1ArGrFDZ5uq5sAI5rFYsF5u4kR6unbvwOb
jZv67r8fOfCWRAt4X9nTi4ioSu7VdZ7qg7+zkNqksbpaoxf7b9enycsyce8MhyIp
LquJK6sy4k5Uy8pSfVSXlbJH/JNDG48iynTcgyPLwAZWILjQys8kwQycXD8LNpO1
1FVT+2B8ccGbaVeripFeLBCkB6OiIBnd5h6llOTPsMKRj2IDCTMHgvbi/IPvPlhC
dZpQyOTkjRzEUw4Ll8nDdr6bHuTl7osHMhlwYKUhgM7v/W+ezTGObqO8/D/1Raq+
1EV8V/i38HzdKSjwN8fqFAPC09mK9fifex221PISs1rg5V6pMtPIWS7GxdtfaN2U
IlD3N90kiKh3hFLczFi0kcF2pRtdSkHWG7ugbMmgUJOh6uTRHI04z53frgpNQcmt
uhrEHsj3scfEkJCgDOvQsua+v74QFN/Wpvyc7GE5Zz/n40xBNgCSmysoNxnfxSgv
hn0yd27j5KXgEVaR0Sgx0ChxpJjRr9Cmi/DarzUEgE6knDC9QJ3jf1CegCbfMW1u
j0RBiF4vkhJOXKx5FZy6sGhBvaAPKOwIcNgglPIPb/MRB8lLY0zuItU6rD0Sn3vN
CIcQ9QnAK5dsKmD0kqLrzChy19lzdzPGUZFTbXaKA+sSCixkR5QOo1JA+B9jomTz
zeoMjncUdxqUqxQIzQLqXj6rAiJIkLRad3avTyYYVGvFClSgJAYDJ96CVIeGqx6j
pygUan+GTpVHPP+OXquLknYPRm8AQUHkQYR2mIGWUh57jB9j4bVhotr8f+SfyDYi
HbRhJKqBy1begew3G535CoH/4sBqC5a/lPnZZb5zYJyZiLvZM/Csm2UiGQKm40Sq
6pKme8+PZAGxn+pAVXITGehjPq7TGNhJbk7GrvqRMeKgVCVeygnOWfA1u1yk/Ug1
EFX8d3C/CQnkTuLwj3BJmsWmgnKV1cd/8PliJKDjQO9AmuvMtc40Pi2q/ht5RJby
uygfGvyGFKPUDMy8+TwZBraRQd7JyUwmVod3GI5FX1cqatjga12X7eBwGLfq0R58
rimzOUh9L/wU3eSVgN2TXSETMndR07gjQD6Gw/hfyLYppw1yPh7RfD9i56c+gTHX
GA+a6hCORaCemCmbGcz7Blljd/D7N5FFY2Hgskm6rj30i6eZGP8uvzgGQa7zY4hY
JN3YYHTFdt8/ydbAgqTnxRnYxVVcH5GcBtVc/ns71MRLqQEZ2VfNF0iaYcaDhiNI
fbsJovrZenhbIzXdtUYigLixfFjnGgJD12s6c5i+In+M1GbROi5a3Zr5kXmkfGIr
p01uaxWXeNVQsqN+4FoUYOquJ7LtKaZAks2P9QbCMyYi8WF+20gBeAQYMCPhPbRz
xYctKGXZczIdejdF5UdHGIhyJDV7CFtSmObUP2MAnC03CBiXi8sDGDzwD2IjcgHQ
SaVjsfZEnE09uRixL5YTNFW/ZHT17zmoNcoYySJ4oGM3sQkbdotw7hx6kOvV2aJS
8+gayhRBrxiVpIdtIF7ma1eIaJIbBKn3/e3BxZaDAZvwxxi2Zj8SMh04bN0tuNXI
aOqxcNcWyy9q0QnwJBV7+T3PDCOvNlhPN5PUgARI0WjYj8Y2YDDc1KGwi70K8BPo
Bxvboyt+k1tJga4w5oXWFaynqVDfVBZfCpJvxzP/ModC8lGJIIKs2bu8gzSUwGVz
/bcI4Hfv2PkT0ioZjkArFwMh/DHhF1s4m428M30mO1E9HVijtwgnRVosTc1ffZCG
B6w6Al97PbFtriendED1Rf7JJ+lSy04zGjR8+TkoQiE0shtn0ji6pvlP/QLmkLvj
XQAM/pku5QLJY+qAtMca+nc5rmbOjS9QoVF8Kp9Kctt+UnfEDREfrH7E/dLkws5j
qOeHezAs7mIU5yvfjsv1ftWx3k9UyhvbQEvLAEMO5hvlYb1kdDENZXJj4ZczAu7g
GY8jiwLj67TVfijzXMrZ4lgvEdDJTZ83nxCPvU2wurj76SN6UU4bAb39Tze/AkKM
DL/3mJOTSIGsmvcqEefU5H2qxYj5o0RTMiIPXliDPbAiHLNj9H69dqrDoNtqT4W/
TnmzfR8e48ie3EYdX/daB5c1WcocxmBsjQjxXWvOo4pojwMfGky3vjU5fb5VmPak
JmxDB/ZdnyaNHfZsgxpWMhAtgAu2/wvaoevfFWFeaCbvJI1Kx2FJsWHxmZfXvrXL
Ze3rZqtMVBrrCRDjkJdlWjSsHIiEsqFpMZAXpNwxUj/rBCLjA9gEjuXdoMHNQphE
QCdAK8HsJmyaMZm5d4DdhXo80VPjCjls2L0AjC1+LXSdxNSUN/RvgqM3857uaIxd
+ycTCcz2CCkLUuugctR3ZTCJdKIrwDHYEraW0y/mSu8FM8kflzfb8QeY+UBsyVj4
hGiMLeJV94USv/OWuv95Q1WkrzNisDb0UpOwP7zcoSyiqRKN8Gm1dBnTkrk3OSsD
OAXJ/MWv4jkk0jtrC2HjlgbqbMtDQLw0ItmuDOt29BSra4wJtN0OLfm2TIjYqLQk
kjCoaFWPWqFSiXd1ddwFxDDdPDjrKn/TUAWtR/7yoTI+1gt8X04GOrJiO7YbM+I9
+M7aN5T6wCIubown8Iry+jllqH5O+12SVTKj2gZs/OOd27mYJHPtRH2WNe1C46tL
BnpoafekWBmhDmTV4+VsX8OVyLBn5UPcx7Nhs4MuMUVzd/sI5eFvp8XYgTNqafuz
ODYsRRBvceBLoqRRInM91LvAouGZgrXay+S4HGtjOxAimc/gtSrWjIqaz1SEAOhC
YL1NnT48kbwDrjkIf8zc8AZvGJAkDjRu1+rzqzP4nVvjfpxebdWgMbRS80nA7qNX
63zs/SyCyC2Q5SJQE0dOlaWkdnPtA3/Y5eFF/AV3Dxf1QeRFEY3q0SNst10kiu2u
WPugTjDTRQNPR7qvbQ/jXsu7DSKy4sZ5oqBS2kYe/ex+BkZA10UmFzjEw0Wg95ej
hGTOj1epybHoZh2Cflbs8abnEQZeUWanTy3cTwD9hQzUVbeLNLw0buboI/Sp0+rz
rnLPAoJATDFtO0SXMYBgbb52x68ZzWpwWCtHTOwW07qS3QlIiA4GGaeYqGh0QBdt
SyDtJp98U9UVdmAHhnHUyCo0Tas7pxu0ryV/n95PjnkUJfsxlXU62UaGsi2//xKG
eG/q8E8ReBFPrMLOTlghaMdUTCRMY921yEQWqIhM6zUCpq/SOA3C802AIJpQy/p1
EiwPg9hOW2ZYrA8Iwk4n2gX7YGHSrMgQ7DBGiXOTvvcJrY7Vowd27JFzB/A2AC+6
K4s0rb1kznjh20/5yAJ+YBRdaQveaTfnCjO9+hdZ01IDe9YhinHqBIoR/XG84kc3
HsaxKVw8AOMXZzkC0d91GqZKlyqBq3M5S6QuZ9SRfCOfKtTacL5NE+qJgNyWw9w1
fCIXkF1vSBA3XPhYh4BwwOEDx+Dxvw8yXrTMu+89QA0n5ZrKU3hX6Awu+vgARHA5
hdElZ/IzOJopGo9IPoA43zaZqIqLlhYeus40+YIdJWanIdIVo3nqpLNdDa6atO1+
H8GsIEICfgB6jCZVU64PT+EQdI5OQX+EfALy5FfVVDWdMU5F9OcrDgT0R6Uv0ELB
ecPZATkaWpbJY+agNwJrn+SzhNo1ZatH4+k522NU3X545xb/muA3WPHm1sk4ph4P
GZPzWNqzb+ih0MByUvCqwcO83VeWwl0RiCB3QXbryA1rOiv/uYz7FGfggM68RKty
SMHk6iMHQlrAA+/fhSVGKVxnnLhprEOUqFjD0ph+RHQtxvGvWJfyVsS0HXS8m/Vb
T+QWXhKtTRvymeLxB2Soe8OIFfy5G6R1Z83V/D6b/WQOipJ2IR1B7lqUCEX5vs+Y
LQ8qy4z/C7oTM3trXpAeyRZ121y20WpELyi4oNXRx1ZYR0jVCdW5uHRVr2WfAvv0
LDlLl9faWdZg6zLwSIYnsj6A08WpEIvGX10mNioxUDtu2g99okDx0S7WNedXpizA
OUKGnA80lSGp+iHaR7tu2F45vuY/UFLbqQ97SuWr99bKGc/Sw0mosB1LUShB6QJC
q/iVyr/RAj+bxzvc17YTncKjJF4jAcRdM2hA0BHiv/4G0zg4eleigwlYCmsQb8Ir
sW5xhMwJbs5/Gc/sLBtbkRaUKQSZkGq6JWPYZEP+xL8cqk5SEIWEMDWbUWL0yVuM
cEW1zbJPT/DSgVMhcmkLhed7mqKZvy+QrccfwvKw9nzl11tDlze/T9ITiZ3KpYDL
QY3M5Ob9CzzQJW/nOyBdoeV/qDJme8oyF0S/FcoTEI9C6M8j5jNAKIu0odpPtGJj
RULK9pclInzfuDdm8/XSq+wMjOmM1Eb6dWf8lGW1sGIfKgqGr9MoBeuLebC6YsLl
Yh+Nhv6T7uLnK5/aCWLCEimZm8YKkdcZE2S2XD2nK+feVuiqLbXR32FQJBZRDTqR
9JMiDm4B/ULbFD1vA4OSo93F3SgflC92o+8dnPDRR2gexeUiryv9WZ6gqCLEayDS
A1mYl+hJ7C2wrC+LKEPD8+mW6fFllnBZV/QoMoZv5GGmxAslyRTaDTYmdG5dDr/e
cXSNMD3qZduJHaLH1ZJfl3UfrIzFHFQwbTxkxbo+5pT1laNp25YZ3XFtCh+4jArk
bn3CiNT3NY5/ax4VZRnOYtIimuhiA2JbR7YzGMKcq0o/fhvHhPD5UffJQBQmI6sT
DJfPewDASQMS+kxhE67cf0rKCKXWG/LNN8MLRNur6R1p8KEbuZX1zfkoV7P3FhTr
IfNjTkWNJoIepPam8Hzc2KAGEHfr81gWaGnbJMhSrlja1Up1hEDNgDPlr+ueIi4c
bxKNcaDNQk3O+sPnoMxIrCJ/3GNS+Npz/Vq/CNli0kZXxOjq2O5VZ4akR+F8ZXFA
8NnDGJbW6hDEID3WCHE9/RFzlgFMeKY2tbArJUtLwE413uIifyet/Y8Fi4MHx3vY
ez3lTGBSU3NyAqTQr+EnIS/Ow8SUD5J2HX6E03k2qpTazc45U8zQA5EMB+brMLVl
VKKmSdGknowOThxnTm5oAct27LFiDMpWU2vMwgrXR07sWs35md6nSoBfQkIKC1TT
awRnpBWF32rUWfCrLJOQLntt5QhJGIwtADSpyF8NjNNWpGyMBqO0ekHDNrMy5iV/
ovhvT9i1qQHlxwi8tbFgGgyQi1Zip+Wfzzlscx2BSjNUSBkTUC+vRWf2AS0hx5bc
vWQ69KmTfhe0CmzFuQ63/nb1P3Hv0SfLHWiOPpGl4KCErKZ+0IaC/cB+fO67Mgio
HlW8ZOu7vPAlzpQR3P7hQnExwd2idfwkS0bL5OtVPgO7ZMHGhPfaGYLNiId3H4g+
aSeOY3x7KdIVe9+FIp24OeWH/lXeVjDKjQJ+ESndGO7ZegwBBpZFkyQ3Rl7boto+
bSnMIIdROFQHyF+inDvbwQqAasOnMDOqlN7xcNy/L9TliTQNsgxMRydyvFptvdAA
SVfAEoy/rQCXX3C3YYdQxskyboyiyKce8SYWtMZKHTRcUXGKiZkic3akiBVN0zka
JchwzlGz8sKuVzu92CD/oIw5q9mfZV1wAr2gL28EpJoe0ceXNucZKIMHU3m/Yv2F
yvJ3YgTU906MOLvs21NosPe5aOEpCXbkgMe3ebuZsM6raLmn65hGgqLuv31xIZEV
cTR12K5KXPRT0Zqzm79wpngldgW5IRnMD4oEMHFOAbJ/VRKy94TA9TKyNqxD8+F7
xugvsO8aARKLLcYzFYiY9X3ZMqFekYeR5ld9GDiPp+YcdrazhtLcNU7jbMu+lpv9
uzXIjtrb+Oat1GNifgNLLYoknBQhuT6QzfFmbpwvN9mrWvPlUds4oer5Q6p6/1r8
RW7zdiOPVc82/UL4bTewkK7XTbBh91eELzV7eC2wcRj4RS1ZneBy/iMbr7qQFcSd
0nOtyutX8jWEtkPtdmrPk2yXIrAoCzxuwjBvQSdA8nKqkK0JW8Z2+5MM1iUsQ/Ia
31K6/Kkwz4uTYC8SaJQMiULz9i02jBJ0a5mZtAizuRMz9x/U5Vas6NqOt+qd5oTv
c7ZA9MuW0ZTZQi4hR2YE7PAOMjbBwOy6Fc2m0frn8YwYPipE4oUvmi+FcjpiS/RI
wDLd29wSPq+RPQx/AIOSsfU5Md4FSSjLbDF7sQzNCUat26co99VW3nx7nw3XAgf/
j5I9E8qoedONtq+HJfcD+WywgP+Jc/XYLiJbgng5VrlV9F7L2zCWoFsd9vlHD88v
If24Cyzdk9spebz9d3qxnE/bTYdUJ9QkE/mC7LjRZlKLdzsVo7TABWGiTJtTsaWx
/XqYCnvjbBavXXoZ9KauY8PhDym8bUpn+nlsvqImoNVZm9hwXnmsKVETzZJqYwVa
3VEEulh5SzMKCoy2nHpknsZPjymPLAxHJbgCJfFuS1pZ4OjMeb3QdUZ9Pc9QQ3h2
MClA+xeFrefU/9EJsIFXDbsHbX9tEurOnCfWr05Bdp1tET1wwLPlKiCvUtPKxxlB
pa+ku1Vql8g/oRZ52goGafBeEJPZ1fI3UqG8abKO8BqJ3tTdzY5EIz/1/vNuBT5V
rp4FW9xwnVrFAhUNxPCOLlTkRHdzQmarOq7k8Zs2YmJGV8JtLWbsmFQNgcPcHCo4
xVHPt4JCgq0LkgHUmt6KjwJp3m9lSJxZi73A3xsdxwv+MhdgLDkoump5rW3J6HtY
03+ybQl64I2kdeaL3FqaTaMzrL19bIoB2vRgjypLSOo59fHaeR0x1f0Vc45ufcJ7
zBookK5FslKmxcFoylyD233of8rhrpjISEg5Y0PQAhA5oiUXHP+xfF9SQEvmXXTf
a70FOttzL/Pu59hC66OoMCmU4/1WAq1trCa8AM1l0ldudtK/sp9focoxnWn8anP0
XP266F9xWANcLKpvLK6ijUgOj0kvgRHRc6YIyja7J2vQDVDCsB5LXV62IuLTelKC
7dFllR1/GFi8UL2POGqHmp4JWjMJ1FKpe2RtTizOWoTnD5wA3s7n1G+4VubAYUZc
hDFsLBI3+mcMap2AmTtOqbQ1BYPkrFLhOWe8slhm8ltNywTPHTqDweRmDZNZSiN0
q+qsA+g1HuvPB/EgAS0lCg6ZSEDyeC/AP9dxNRXcEa/YffpOjAtTGcztrOHW7zum
j/+VoZB6X9G9Yr7shtAWALTD1mY7+lSLUhsfQo+jrpFH1jMOQ4oAx/TmwY+5006J
mDlMt7ke6kT9PJrLYjNK+VeYGmC5PTQrTtL4dptPzMz2XFEntPyf3H4K7gbhsV8w
JI8hfMdIq+OSWK6hDmeleeGH5a0sObsd3jex7IVkWMtInUd2/DySt9Nu6QdTB9aV
RyExw6UN1pE9w8a2A/QXD61yP40n+ktt9FQT8hZl3tb4WnjGN5MLBcHNprBJY6LW
2PHfyY/hl4F/WEiiYte6Axu/oluBVXaxxDNL7QjWAYz7dtoVa7ZuhPYVkbDqqdTu
zn1YS+79ox87bTdSqci149jG6koxXYVfcZo/2Mh5JbW4zDcl8zBASuZeiXBJYvLY
qwSHD8/pr4G/dbx6iMGt/GNECIWVCKLuv6y64Pn3NkNuJAT8Kk6UnrbfUV8nmWt5
ihEmBhZVYnN+A4Z3vw07xtSRgWVjvnXdyAVxAJHJjUOTRsW1GnvceF62cCFxXhxy
QIFOkYrgacuEMOPH9od/yhI9H/rVq5sZ/k+PhF1eMlzV4B+0Ke5L0KFM4MhBjIjr
0PbnykpxJshNc4Wrn0v8EJ42mmuvtRbFJs39LCKtu6zg6PJwXdcBKK7nr91qKbmH
cQOoEdEK7+QzCajllujq8L7VwxUaLQEF48+r7VhNCAy74A1ZIzjDcJ22J8QkdCA1
YgzzUYVHlk72zZZnAJAZAIgTi3x+AlYDhlXIR0yJ/+4wZqt/un6FAhEnHbe+hUWT
qvqSi5UOHS/Rhj4hubCjq/4Vb+D/JaYHi6fD4HOVelcWG08HWnOMZBM75eHD5XjR
YLCDb+3f3kQzfty8fj5JByhKAgVM5ynqhoH48sVDZArjmkPCFNfrYNQrteiTAcs4
W5HL2/VOh3in2U/RZNcYRzc5RCUcIwaWLjuXCkQq1CZw78RVjSW+wx7J0Do6bd8u
NBr3TmaTzfNwr1AshsYK/dSW+DQbQOIwnU0UT5Rz2bDl59BatlqWqgeH5/0aPiqo
YmyCnbaW5lS21DH93Dc3EPxuUtQYGj3z3yJln/u1HkpZwGo/PEfPYL9YaPVXBJ1G
H2H4A0hjLa8lbeVD+r+jE7ffzPM44cE4QnR/PcrAmEdfcW0bkv/9yHE+bCujyMro
bOErbLYyu6MAaOgQz42QciveciFrJebpptAFogk1M93n+WI8Rlv1TJwDzJQbwgQS
Cvar6BCq9r00/zp/dAjPnzQVbW0Qh55atQur2iWpOSqTC3ZR7yiZJmN+LERVZqCt
NDooM/SciI7auQy4cI82MkioK2deT2ffnW97YKi/6K+1YxpYGuVhk1RcivsufqOB
9q6U3+S3lFJjFxoHKY9S2m0Jh2a+GB3K2In6Z4mIjRgE0nmJsFSQP4oUaV5Hfmbb
tAf07Wy1i9vVFyttzvw8yNOBjsCeBciNL9BqlJl0fgLQ2lzxcM9zpfqdBDvZV+HB
D0BUR/1xty3BOCr17OHjBN/CENb4hyFDyEDvDlEj5Iw9tKFNOWyWISso6TIcCPep
akfMBKRvpfkW5gzqIgrrExRiewCEFZ3s+D770nmydP5vKfnQdVVMcPB+DO4cM3F3
orR35Uyrdcdk5LK2svEVpqROhkRZpzoiZdy3O0b/SmtOI4iL0rwiiH1saY9gK6PF
jr7PNCgtPr5ghweJ1Y5w6/plhU3PUoGrrEoTCErMWi45vYZR4adW1GM9uRS2d1cY
q/6LvsXJ4UNQvJNTxVbydpTM3fx0LWa+iuVNKIjj5/fydOdK2M5LqFVktyhWYvqe
pIF14I83T1ds6mdlVNpmhekxwE8XqA613DTdz06WMsNlHwH4qYOwjXaRcbgDXoZJ
GfNelEPBzQQ8eg6DkUG8/dZUhePSYIS00AERLhQUD5UGoqwpJ6j4R+ztZwtUlW59
F29cyG5YDQ0olCoyOMoWQRXIE+tnMyBo1crpfPO2/oZSMUGC9Dc2I2qOIYqzRDJz
M+8Hzr8wBBs3esfbf/XYwLJAIldEPDFPm7879iTOi0/Vt3Kay/vUav+rx0I0nwzt
VjMLL6t8fWGAckjKO+2yI4MxrkD7AeIkK4WrT5EJADVXZMejw6A/yt4bxxYcu2ZX
aGzHTPqxA86lInxLyGYqCdFLCP/b/Xy1p9WK/PFrrYqKt0+NW3xYdpgaW7Mg4+nw
KpBJ4W2EqtBEtmELGOoZTdGaOgme1tV2dMHsj4dRYQkfR2QhMmjTGykz9wdkt57b
TOubRcwZdxLAg9jYX9wscD/uD2LQBA/Dufvi5qNy4T+IeG1HMlYQEigFv117pKLC
nVZE6XyRgsBCxQTeZY3oh+l//NswzFHhCWoO5KGaiUQvmx6TuUhJ57QMTWMUDZSw
mdb8YEjN/uSdNxwHo7ZUQfDE0e2sKbfsUBLecNfWEVnlT8Tidrl4fpakZRWNnHl7
9ASzjaYi2/rW1yYofDMT5csG6HZ+rnZxyGbwTPOnSlVlfOvru8PDp18cr0FhhKFL
/d6D/puOol0dMI7nZwFwpRkdZx93c4QWMpfKVsf2FRe5CU8jFW6+3Eu03+1hPTVg
rwFjwKRX10ain5ZFTm9f35Omo9Q24z0rU1W7cXkTdobN5yKlNZhCsBzY+zxz3uu3
VAVsh05GS5g7bwsFkUjKKi6BJx2zJTMet5VIr0mJDLfmKs9KrLryxDpPEx52TwHY
TtobkoMFHVVhJmfwGu8EJHQxu6qykIVMCPeSB00VwWfPg4zUJozIfqq1d5A2S4a+
yqVEYPuGnweXVHmLFeNx/HPQC0guzbVkZQl3IYHXJi6tnB5ddGZhFGMHC0AqUWJ7
Bq7SVWClMC21VEN57+cZqa8RAjtwC4iUnMza6sDflaDPePoCNp6eAEluVo9Wa1Te
WbeT1mhS2cTmBxzaG5aSvfQ2FJeotc9ajrPPMuzcQyiNrgOcxmTRycF8ExtvNZv4
G9IEsIjTtj8kzhhgxBvN086amKKs9Q9JWatjRVoLz9ycOFey4BQIkW9Zlg4VSjXG
nRKFP7xrJQIG/FH9Q7jr3rtAU4FQ6EGQkwnGpLvtFAlR0Dcryg8NNMV/D2B3fhxd
yqRoFvytm92iS1qjECM/aeqhNO3AfqeU0QmWvUterpBQJYqNc6fqEZ6hwYsp9YpW
9y4KHtqnUHRJJQyuvXBAP8R6lvgan2A74fiw99+M4UawbqXLMcEpz46493gN1PxQ
xmlMYxrbaFMwjGnmuuOvUHWBMcWFjVJbGYAMz+43TzmLzk0qqWnQmVh3sLsTO7n/
1XfGi40ptNafLylQUamHS+Lcym/R3gUov86VtsknoI2f6zPpR+6u1pBzQyD6rtoB
RQBL19U2uAfsM/idEtscVw6/OVk4jEXQKr0TfMuLVAZ0eYuOH7mJzTm8pKKHM3n3
kc4nx0AczLkFbnd+Vxm83G5KTkplUk5i1vGpTJN7nDDl+d/kEhGHBneSYiXTLaaf
YevzKU8HyP5cyfnRzUuKXNwmzYyg+ZuDuNpGQ8qwR3XCFlHKLASjFSNtxdNhx46W
B2XHhaQfZUVE+thuHPLOQDZFOs90A8NpZYIR0QXCp3UIaPVoWSjeB8KPsqV4aNhM
lka1Xe4Hvy1nOvQMSH9SJhUgvmJ9IXnHK8zAQQ7eaPwjK/MToFaJxXLz0SweJTs0
K6NCD/psmE/Si244u3Dy9DgXxElsW3DgcLkVNwsUqaYmE306Gs+MoFIAtvqMgSiW
rJuw+ABLvDk2t1ShzGdNVnBDbRqWKhZB9VWpUCX+q2St3uexzPVA5gZhXDEheYnF
B/fGnE3y73Yd2I6lcn/8L/iWXPTBKI0ZfB9FKhmYgC3ra1RI86Q8xksdWGoJvtRP
odGir36uigvhmDdBjkQ7ZG50mquE9ujqQvAMHTWG2ES98ANGv0Fno9Na4xhlx7po
nCZuY+vx/DAPwVMNBTH12sd4WY9zW1XE20dIkXPxK/Hp1Eg6yFDmzWSzQhN6ZcBn
4bHD4dryMzk8nDkcFbL1UOFugzrYDhQd7e5CyjJ8H3Hsv8cvlsOHKJK9fX4JEkp1
RoSh6cLOffmRx1VUT3YhvoBLngKwVQ2VXvBoF39XdScrh9ks5+gWxSCQm41egwBr
zu3lMzUSmtlj0cTwDQGNe5byqyeUwlo1YTVbvj661SwlW2EL/gcYK0VLU/iq5TDQ
hHao6dkVyS0zmyLT2nLiA/w2Z5hytmac9q2J1Pr/1TpnWshddiQKM2XrxO6e6H/a
aAYmBkFSEeJc37Yfh5snWeq5ZmoAz/V7jr83qi7/JOBNQwG+NAOlBf0YALTyNdmP
6ibJ4V1L1R81VHIoa3FVwvgboKgVrjXnC6WxNymCdFNqKnpe2O/ee7LaYMBLW1CL
UGgNT2dD+1a7Z8xqjP0/j2+EcL4EZNx+8ofsMlk4AbdDstZrJkCfmvll/qtMSZd4
4Cf6hM6U5dR2VyVxJrXSAhGqOKI0oPXlQO0ONucnYHM5RavrHHiF6IhFd7Pep/r3
UjAgrNkHc2zCRKCNn9qRIqCCSF1NI2pTsRVnLhI1yS49LulfGW7aSoWL8M+S4GlE
C0aqG7OmLksA3mWIhTi0pIh7aI3gV73J7VaIybGU8LP0Ft4sTZqmiob1W5fj0+DJ
FJ2CMfrypaeDPOe0hre7tJOAvDKURQosELYKGaYeNoJnY67EAm54uMkTax380O6r
Mivkc3MPhEomeLh6uFRzqfWLGRrAJPN6AB4UqQjASGGgjQMr3/MizWdBES+4PWQ6
M992Ep+9ra9f9ilgkJ321qtgyoHxpjqWJ4LiRG+eNgKlxvlYpLyuP7E38XwbRO89
ccj4YUvBHvZMamIggsYh1RREuJC2JvyvHQh5U5NTQxvenN2jr2YHbPoLG6R8kLLt
i1efhZogwcrGkkP7hJfo0FRQJvT4ObMKsYfNBzz6Sw+5+tDKEZt1Zi+4cqrqII8E
AHUKs/d7vula8vEsMXSOOB1m/5HKQ9BGxxOY1UABItn03PKIeNfHgk4tiaIaUcur
rpp1JdFZNCvEsQcZPaSCzOI+Ws+f6EXTWdJCfnb/MzVacbYy75U56wBmqTXvUIe8
xSGxw4MGHoZW/t1tb1P7K5vMXokkQy3I2JCjxqe5naynyudW1ZjCcPo5LXIkGHkR
D828X4ADcnBXotyLz1d7WhKR+XQpIyyOMBGB+ibDMsNfwkrTBy6HbRqKL1UI6Sw9
fQQfnZtT+ETQmfcMpdRbe7yeZnbUDyKtFP6xxmhusFRWfK8uEzUpmgosbqJju82n
A7A0qx9vZvsrNeMiofOZztOeHe4iAVdsctCVT2kgbaMuhEhqst1Ji68JJChrneXg
2p3x+Y/rSnhjujCQ5LfEdyuxm5xioFMoMjFhOdBg4kg4RjWry0c0PdvNpGCiSVtQ
fWFC6Tqn1NIxbhn6D1QDPavNotZDKhk/fO82EbPIXhP+Fggj5x7GrdPAy53hLold
coye4LExhpxd5ZdGgCO2c/GSWkz+PNipCzt18ZKFFk+RtxD5+oaVsHH3mfrNGd/N
ONJWb4tbcPmvJZ70SS9fcOqrMlLPEM8/JOZ3nV6C8m+iOUhloTDAzYbp8e3KwMjH
vLLDGvjyJe/V0MtFhmVJgKkI1XvrIa0OqOd1Mp5dOyUfg+fmKGU9pnovPhjew1dN
XRh3iz7rx9CqaUSftqsH90m1SyNjrATeXKqQ/jruly4EmwBqwGPnmw0tVNYxETOd
/+qq9YupgH82uzpFYnYw10Ictu6uwSFg8o0t/qnMPVoX3c1Uim1ePZRyG/d1EUKn
al3jVFjkQA3vAQJnqIwGCtkIGyDRTH3GHkoo6B9Oy+JVmf95OM9l234dTFEgajfI
BdaVu8l7T9Ullr6wwC7imL6aM1iqw/JWWrzXyDz7kA3wfeDil86Zzgo4jht7onGT
RdLzyltou7o5q0HLpGZqTA8evZwJp1n8pUxFdZgIfxX3caXD9BSVbzmH/2nWaacZ
paWy4CSdZiODHe+bN6Bk07TKq5IpWIxbM4mpeeKYe4CxxNAe33pnNGZQ4a7iSKQp
Jc7GzmoEpjH8Ku+v7ePI4/sk3FCMxoDRiU4oWiWw3tjU6G+gcxYtSpwMneMnIaXb
hRVOkzqinPd1gebZN4ZeTGOhFLe5BYJWiyHi2mlCIfifIUfR18JPNQizGYmhX55K
mDmeQq3Uk4cBSY7tjPTVf9KqjPHLvY3hSgbtr6EeuB05BrrWyMHEyNOvZjGBiM9A
UT1h4JWcfoaKXdk7aAZsZZEdz9glNeoK7rJrpmWnyFKbygKMSIZo2jzJz+EMcI93
PLj+Uh4hpX0YvHj0+SwLXdBVSC+G2F3hBiUShQDJ3N2/RiPqjewHXilkIqE9P8Gu
XoyC+Ckn0zLWdy5GGUfHrsAVB85Aj6LbofuiDDQqYjHVjzzrtrc3oSbHI3JieUDw
bWZhGSQWCNth6icqSXLEipdqn65d5Pqar71YIiO6YhyoD+52qwWgyVBtRe1fshFi
1VRv6J2y8oz0cXtj6f73C+ITWgbZst0Cxw9W3/nYdMva6XwnYhv0FO2Y6WswNJD1
xAjC+KBcjEuny5yOqEUoA0Y7TIVPEYG5oSCZKTjLOdqQUvAWnpwZqQNxlWpT36GO
qmpZevNfBDSyAmqKYiMbNSeTVUG04zeM6nr0tKhT/sgmBfDDPh3Zw6KggVlLLQoW
zAPLpQrG/6sKHnESgGtuQEeChNNel78vTu4pd901hTKKXJMvtiIJmL5IZ8WxLmTg
FqXwxv28OvETyNgLhfZOM+fzX2k7FNDB0Fs0mMWcAjM5hT0Ye48EtkdpmsjKgdyo
WYoc3cqNgFJVrOnP+JFCsHBgsVjZ7zboYnOt11yvIGw3SAljHkffXBcFppsT7H8E
ROBo6cO7+Lz3phig8hlbedtnjvagUgDd7ekcJPuAB/U2FSggDuJt7IyVUwDtJyNM
/LWBsDCvPMRCrMgn7Qc/AMvExXCNPhbqzLhQQqX8PIeWKUgDyzGpTX3K2tk3UNBb
uPK59/Q0eWhQ3cCtbIzN1yXfdyWa8F7kqOSJ1GJtEh4a43WOE1/z5nqQ664t/ue6
jSUSbRWqcXVlitwhavvC6grHO9wDBfes1aBcoeq3Lh7pfvFki8FHFAUtk3AWiRg+
IA9jidmx81y/YM8+MyXpRMpZJwliKlV7vewveureBcnM2AldZF7eEXEkeMtwtPNI
wG32W4tpmbCcQSIILVyeal3kTSZgOMk7mfqJFScUHzow0iU3n8lrvMh2HnGJoT6X
aS0TL2fK+pfHp+NrRZV8mNpuOac48CqvrbfTvg7IyuIYWXWxV4AnlYmoFeTm6FaK
kd4NG8aP3OwOF1E/u8uEQBd7aGFKs7UAS/RCSJw9SVBT6Q775meoG/liwudGvb7G
h+1tU9k4XsBmzkqrfiUcUUjU1/8hKsgHnxTMkxRZ8WVOvS/dkVtT3uK7CcZyBuTJ
JsrlzFur7l1bjQENzovmI+QK+5UB47FzpT5zreegsa4cnbMnDNMalUhQEFFpyeD4
u7Zl8QS83+8USZupASTAIbY4kpRlxLEiiDNaw9jFf7sGn7DsDdvkr42ZNE6txnW0
M8ekbYPOYi6Ek3X+YKDDGTBEFNkUyJe2OxlWIdShRZJgliTLERJ0J9zXxT3X4nWo
FloDQQ2dQDF2pJEMmvWGs+Q2dik7KU3kOkOyaKNlQDT2UHNs0vMWz0UK+k2rgVSr
09So8WL1jkgFCgKkgrHVojLyUetoir0cWHbs2uG1J+FrPQ7xJ9bXr3a4xnksZNAe
kyyS6s2RgvAsCKwgPhUQx2h2xSRDV6xKvIeIERab6mg7jh1afPwkVtici+XOvxrU
aULbow0AyD1N6FM0dwUbrHYk1yRY+lD9/di6PWly9zQTBGDogLsGCIMVdH/EQ9Ha
xVkvEIGNMGcSL0dseozRNdRell4ev5Ne58Od9+EeJTpgzU1l6TaXdHBODoOPYOfh
eMcngj6ddlMUNiPuuAB/heyJyWvfQm88gNCtKQxJeFAV0HUSwu0VeRFhzQojQms4
xGGObbYNKnTAuaH9hNgKH/3shkxli/DrDQZoV9Xt+iS5O2tjRmmR9dIt3CVQhgGW
lWOs/uQJsp/+DAT4xqtkmK7eySubxwRFly0J2AkCeiqUUnPAXNXEpsVw2XM1PhFK
Y1GEsJYOIWzoGGK8HElHLjKArOy/X3BcEaAwRyR/TJwz5UWcQUSHxyEqCxJvMQun
8DPWQH4lQjQO4IpVHEEcfT3UdYGKYgiOObsI7d/JIMrkntiZ4t5HLsFHEc+uHP5j
6+dtGw3RDwHdNg8my7eM7OuYahJC9H4R6LFZSpzc5E5QSlWXwPoCAOfwys17i7/0
cPFRYtcw6mJnKZtkgsokR8yNzY8hVLznwTBtu3UGJQwF2vuu0sW8ZRgobxgE9NTn
KFiKB6Z18xhwu7VpT24hweNdNTBKLaMQPqoAaarV0BQWe7b7JlJZeYsXgX3OIQ0x
hyrQ/kE2xIH+/w25duDjMNF08lEZ1uC3+U/5OSeP9UDf9+ELoxTe65gVb+XLPAh1
SlI7yWjV7DV1Ep5UKOj3czt+EoV0KOwUS4z9CBbEjWUl4U1UCbqvTS1x+y7jjHPR
wZS/pi3AgcHVf7STwhlDcfvgX8CCxnV8WEF1nH9vU/v5BIKHSDEHVMzV8nV3+Jtn
xAtmpJZQETWj4KL1JRZA8VQLb1G8e1JdLzWFQNUvwmLW2ybh7cPUVRunChZOm2le
yTBLUPXxuEk/Zw40DVh0bhsO6qDXLON3F/XCyc+7AG33maTS9vonePc4IWepyu6Y
+MmoNvplStivLkmVJqHyYz64e1+8inDV0yEgJ7e7N9qb1TvoMrgHCWJ2UqqUyifZ
OgZYik0quEdYaeXd3hQYQNeEIKBwC9y1BByuhR5jdQV3vr0pXkn3k8bEl1R9eNsH
AqlDZZcQdMgyaGEm8lFaID7JeM2ORo+HYGNohZc8uAHG07dtohRace6tflmgDfl8
/vK3qs7SmvU1zUxBq69h+xjPR47MyHPyhKtU7lqQ6XZ/3GPcLmaXXMj2v5oV1n6t
9S7s2CAGIkBMiEhTWQzPR3x31YJKS8r9ihXUptWJY7stkCHfcMqsY+ma3NNQhmJw
58j26Mk3at7ioiMO1p4NpY5OVYu0pp7TYDdlo/jIeAu6kdQVHC3ZrsNPbJwZmsL0
o2ztPGtggLP/p83pwKG35+xBHQ6r/VPou6vofXtgW4vPkcO8xQRRkMlJfYeT7RXf
zeAQLwE1HiwQX8aRENcsH7fcTInzDl+1LkaCqyHaZ23+24+cFgjLaZvP1UtITCcc
dpXvq5Osq8MqtdfdvZlPahgntAlZ1082js3q3qYvir/BRMIxsHwGepdNi1twxcQB
OwZt+LKcA9uOPb2TYAZ7AAp0bnaGCsnWcgZtqk7EZwN4wxOgoRYgSBOoW+VI0a4n
JMbjkOLAovKkmqAnel0EPHCFjg3CuT+VjEJ5mi1WbFGdzVB+o5UiOt5mWXXTrq+Q
aTu4H9nn2KJiqr7XT1FczfLKmDWDWzEMxy6RtA318izUQoQuQ1VZ0vop0Sr+N20r
/DQIMSNTNuoSdizcOEvCZ+age4gPlXSN/sGWGwWYOr6Lg6ICOlsvbfHcnoDrqQaI
tLbq1L9u0SvzjMI4eve1mEwtMzn+4yFosKq217Xs7TSpduvVygDfrUEdpIncZGX6
T8WOqUnLYILG/a3jTEMTxd9EJoLTVtuX1cedjUBE1prjdEZGCoJop8pb6f3EoqJg
/whviKmUK4tJ28mkOcOeaMVqJ7S2iRRvjA91j1TRngSYWYXVMX4pVAQq5deSp8+2
ESuyW7L5Z4FlUOsTl9gRn9tD3t4RdOPOXbDhyv16TZhT4uJigHY8bQfSpoeEmVdL
BtqjdEkcvDFCGmO2hSHzv8avPzIwCLeRP/qa+s+RR9+M0L/E5B/tV5+nGryjp8GN
GGtTsD1vlhqD5ao9FuaXPMepXkENZZhVrT2wvkcgz4kxiLQ9OvHua77lnyPTvK/T
txZWCPSVOiE3hsa1l7zAEgmIoa6ObY36HE9qACZuAl4lmAXZx3b6t12DMevMe/MW
OxS9t4VZmgu0vtL8uOZGV/VWKOvZC800hXIU6H60azSAIGas/+ShECQm7Xw2GLOe
UJ1qHgKzW9NBkmFneNZafNdCK7Z4i6x+jAEKCLT6dl7BuD/4aClmymy8FKG2E8Ni
iCtMAvB8YzRc5JsRuvgXM2UMHoovNU4WOUmLROx8EInx/ZqaHq3AJFKYzMSIX24i
UK64bHIEzGcPE23/QvzoW+ZDN9Wi9Ip2DD3DshfOdZAXbADKBMy4CPRODMCjTxXI
OH3Hfg6eVaLhpErkvgUUyb7WHqzBFs9WmbWpORnnycBLC3KS4viiiC7Ji7g4QR1F
CCieHkPzzTlYcY8pzW4IVFnUelKArp2mEVnYBs6FmZhqPsl7s0kIJFrX92T+Lsag
nJxOZf1mS03wUE+K+C3LTEvZsj8dzzlLzLf2EGUwQgaBYe/JFW/ikTLFXpBfzrDF
6atTM4GKZl6WfRt7GDyP91OEvHHo8Shu86yPzWSjQjpxS8mrwkt/0rxxv7AGSkTK
MkTcJGDwMHI+aZJPQfvPOB3yWYzPWki3U5A2vNJf3jmXmhoGtRMZyEX+tW8uCslP
tJXuy04aELlLn7Sq3gjlDhooTdGA/05Ak8NmC6FbwPu7ifNIxwd2s/aeC/6ZweVu
kiWm4mqfmuhfsuIHNcfx8CcwASEBqLGpB6+tLILnWyVtl4gMsnJ1k9/CoNqueBGz
T8c2b9ju+9F0XX7EtpBeegYtb6vrQCraTun2vRVN/K5eQ8K1+2kW+4tJgWFJCG3X
QB0+m2C3eIpRg8b+Tgnw1CUoVI1KLG0UfPMjNvHPLEiOcEJLr4fdlEjv7ehIvanm
In2Sau/waUBO+so9e4upfHMHMmJjVfSxVowo0KwoGRQfOmLu0tgWUGoplry0HNbW
sWfygjDVKbYfxG17+yaXFI72MtFQXylXQ9VnXA689WFHX83++0fWhh+s3Zek2PjG
hUr0tsVcvwIN7MInlM/gCXHy6a2aLwLZvNyuwkUHrfukrjqC2LADNsQsJs1TttOF
+8LTIxVDE9WQWxU4nK+UhmGmLYd7h8+D8DaQrWor+MxLTFR1WlUYgBVAAIR/RdPb
E0/j9VhayT60a0e0P9tbgYuMVqFAS0As6MYbSC6pKMDL0x1UC7CPJZGCI8OEycD5
nBmHGWFF2BxZRa6ZL52LfvvjQh8KkGjOW295ph801jPbH5qG2vGIA1sg0KFA0Ns/
ggLrJ70rzWaqbASDJGoZVQv2L88VtNI68sl7dpUDVKicvIOTaD3bhPG3Rd4ZCGw2
PZh5Q1Y4Nj5TFdcl8yQxUAwOuz6zXUCz5S80MssIr4F+VZZxxTN28KwCR9JcWmU9
GgKHIDjpsqvkA7Sq1zv2bSq8YUBsYSk44OlFJwBn+JGIbomJFoH8obyzaYlMrTj/
Em3MoDnff/mzfxfPQPVOS0ankZ9vjfw9+gnhKtr8CC94TcLtPN+iwf1RKkyLFABC
BCb6GfSwZRPOEgGKPgS335femAnFEGODSH27MzeTdDz9zT2Y8VifWs0DsyYY4NnR
1o/S6PXoYEyEFObGH1A+58Fuo/TwP4FJ/9QAqdTUybDJ/XR428inatRyibW/L6TN
iw0szE7GJLUjT+fpmwsWnFyFsM+j5fUnQZ941MNAvFjsMW4qOESBVb6i1llW7RQe
wydg/d01Vmjz8Be+WTkHeegJIusr93Q0xd3mygdiWzKyvbFcCCJmk9WORXB/q4Tp
ANDUfJAFWWLy5WPY3qaYjyGrwdOxxKeiLPNjKyOdbE42g3DgBLD4RCILosIo5fpW
LcLNQJy+nsjTRwnsNi9G+UsbblikxsTaw1iekcdsi7dUW3lUEP1B5Z7Hc/Mq0IR1
A7SGNviRdFnTkg6sBQB8KJ4qMVJJ8JwFJKSYhs99LG/e8NRVvB44SNAIn9QkJW5A
o74CA/xefFMIFxO5Nj3NLOZVOD3IfZ5cPjW57PyHGso8W0gD6qHrPn2F5I+UJKI/
fnd8Ncli9rJzNU2kHa2DcQSGGBuL2hllKOpp4QxKU+6LN9MyawN3ZRsRDfFkNEMm
bAGCa9rUD2y89SixC2GJzu0Fc0yCgaMNaQ2dQbGW4GnrUc63pWty85gqPxH2wmZR
j7jW9nLGBIxrsVLzL5gAbDPuMawvR+eUEIPfdpahf9k8p7r+Duz3d6r0SGBV0sOj
zOSzLiP0AqYwcBR5l49WOaEH+74R5lsg9LQvOD6nZJOON5agjpEpTcOx5zxxqXj4
1tSMt7DlX8/ga3pWKDuJZFLWiH9tn8qHtZXVBUebtEfhPxIpwK21BccWZQZvO0xO
rWcfYQAaZAPCeP51SqSroo+9z636+JV2PXPxUD+sTBT+YXCg1W2S4cf0l6sJgXvM
IxXkIDqR1NkjXzPdnHfxe0A+WpLSb0WvvqADst924dFb46y4Pz1jrEIvQ4Y1EMR7
ASKZBGF7K2Twz9BXSTJfG/1aQnahLjIIVReleazeBJDJn7XmnVvQT80soZvSlRSk
L5c51/vyRF4kT1rjLIdzeYZJpTUCWDdnz5yFMFEDhlphrFxF1qptnmLcAZvCeezQ
RoJYtoNKXi7LPvMegNTJ1bcMoxztapNFC7LpQzY5/sHmry9rlGSW9BlvZkhiBHqh
g4oo6BzlKv+twu8xZwkzgYrH/ascc3WlS55/8uEiyjyea0x0PPN+6dMOm25YFl/b
1cTCkp26E9sOCSgVuhESRsJPXgRV3//UWblCrZ/DLBCvgML7lG+Ot7HbSS5DLvOP
dwTFB8pS7BHY70HRxBz0Hq3ndXGsi6FuBmyaMWqqQ15z3jMFPTBHAbSmE5hhIbTJ
mroxrb83BrZzd/mHEPAfOow4be4n4Q0QhreGtzdJ7TXZIezvua5fRUl8WFpavXVl
Qu/rJ63xwaSpOXL5EKCA/qi1AXLb3hLbI6gj+wKN0EOcwGgH/dgmcblDK9ICB9mW
NM8j870OAqmV4Q+/jw+NBeXO4c1AePd//C66cfMABTAGVXRnZ1mZ3Rt5j2Vt58Nc
H+qiNOjtivdQBDM1d6uUNDrYBUwnxdaRJWwuuOdT10+fkpHxk9HMnEW6/jq9Zm+t
fTxWe4VIuVMt6NmWT3S1jQqBDIFElVAoh7r7LIuQ3P/OT9SUfY+berjcLTtmnZy9
4rqG5cBrJm9o38IKVArJF3WFZmEFPyEkFLo/SaPIoeb8zKHEAfCGKeXLRBBDg2L/
vVf/Fe+8tVBRG0Z+tPXtBCIFAqBcq5uRrnxmuNMalBfb8Fwi0MODJxbpyeTj740h
3SbYIVdw5eBjLXqgmMFgjaO8A5SaTK7omDkHMXHSt3oBCUpcxr4PHfZMUCZJzxl8
LjOZieDcNbJoHGGnaDoVSUxR2Pm3Tq+D/mSmnbMhD+2OPz8uC2GsPrjmNog5pWzB
iDnpxTX+ofsAlCZdrG7KKJT0NBGv1xqyacf+0NAxALgJSWg3wzmIOC+1FhYViS6F
0Ef5mvxv8WwjKFToOzIyxIrBRDqI/ePtTlL4SK1c/V1NSO4UGEsiuSae4xyWtQHO
J/2IANQMM+QHmyPWDeFLjiLrEUxV6ZzR8fzwahak+pU2fD/Q9iqXBUfpuSnDfBLn
5Ib6Sg8yNSWtvw8Hu4cdC8axCSmaaNRsFkRYzK/y2kk/rigt+2uMjUY4u6yXT0xo
XdoaJ3DdqAGFaSCKc9FgtJV9d7zclVQpkx8DYKxTsPLh491Etoob0ekHy0ixGoP5
u3izlWZ/sTVSVAq7NbD2/ChN65JEM98vBxI28ICW4AQGKgmomqo2a7lmoT0LIuDE
WDQ+w8rQEpTW+dpn3dXxfEfHS5JD6j5T9xGwHB1YH9pTPWWSR9fNvWTee6TQLZhx
YW99q7Tsp1qebLz0RkCEHmkHrw3Hv5RZA07WRQNnB0FGY2J9WZICv4bT1sUs9V6e
8G+VjUGSc248Elxc6SErrH17ufwUuTf944i6sEw9Ej1c7mdb5TQ3iqcjZ7rXHIUS
qlGhz3BIFTnGA7XlMI6jk+zfaHHDdej1hCqow4CFjy4BO9Z2Wn4eKrpkDwbSXVmg
XOvIi9V2s35ItTT97q4ODkzSnTIH+xBPCAjEjRHceIxBfhmObna9PwglQTwYnGYx
8s4GsBnjeP/9VQ9QHzddFw9YWvL2Bj6FthQVaiRZzUccAn3XYLulX52M23x/iUUQ
gLGNGR5H2p2mh78lkZW3sEofM5kfzYIgTOYF+gBvOLVJ3WfIYpiBvO4qOUc3frY5
Tkk13/uBZfFCgmQuxzzp/xgAoSN3jf2RQeXwmZiKilmd3O43mR8lyCRz+DHIhCn8
lgkZNAV2aBGjiHhhPxbYm1XBtX8C7/75H8Z4UVyMO2ET4AAvye3X3U97MII8V25n
VM5RoZ0yanWlPVYt306GysRG+3YhXTdN8kre+GEcM2lfJLvRudwEWTekrVHWAvFU
5xkg6q6CacXyx/7Fc7Dym9z7e7NwBQGcI4YeX1MwWR3P2waGWIAZSra5K8i8S8oq
1+PKApmZx2hPbwNEZu8ylElA9FxCpQTUXtVHz6A69ktyG+Y0+yZPjHxfCPhAm+KE
UVWzFIjDI3H+vdJ2FXpR7q0jLkhlQrVxSu6Q//wfdPgYuVcw+6TXJtPcKO1RWZI7
j+JjUoHKZBJLqTiADmrX5dtOue+zxMlCERYtXUH5Oz4txzP5TG8i5guPiXg9ldVs
TrRmIshQtEfRplsAEHaqyuqnPi/fShyquvPGee0VSSzW6U2a7pM7YgUcHhZJRprO
tJF1dOISDV7eXQEE5QrKpZJjeGMnBVDcRR3/4Hc5yLK6qxyA21sbLp9g07aJuLnM
vFBlPIftBddMlx8gi0Bj1yK4c2GI2GVqTXzZmjEvlS29JJRkIdHO8SHlMIUS6krN
+sJepDaT2LrHNtzl//AcGsZX7h0Z4LEv6PiMwby6UzYc2+YPvOuT00NyezqZhusN
PiSgC+Z9+eHbl/yPXgsBHYHXBwjm7SWAiX96L5j/PwBifMVzGKui4K+ZxCfvUrqg
RhXfgvW/pybF4yzUpb1+eg1S7un4WWV644G2yK3S6AMYDFb9j5nVVXKjN3+m+kX4
bXRnkUiFK/1cpjyy1KM0Hdt7vZ4qVYa4SPT9DOx8KqGIaCDatZNb115N+e7S2NMu
bip2QbIkewIlXTEIciDsChBBwD7tu/QfxFb9qsoaBElNeqQRmL4Mt/lREHxS912O
u4tPFX5ogL+cwJmehtjcL5TegmqBGqS1Kk+tLQswnk7f+w83KYvX1ANx8nCkipMo
h7m2pCFdeX0mDvRGg8fBTK5gK9ppOiPB1arwQn51AQIeB4KTQU2NPnn0JJvDLA7d
4SWYA71jhs456Z8ZFunFoup4dKbE0jzIOHVbKCVWs8mdREbdz3RrBlnFnoyXYKrF
EW9ROPydmiucoCwC6COZB162Gz8UkV2hza+SJC0qWPI9Igad3bFt7ibOEsljIL14
tZCQy6zt398Aios5lPt4Xmd0319VkuSypQMPy0ATrU3D0mqbuOyewbzCLhJCL5B7
VFDileuiGnc9d8QEaY7+7VqXaoYeQQRvEppSeW195b2mXA+QbpNfN+WMrf5x0LJW
ukVc9DLincNH1ug6L/JuOhnhyIo6NMeHCNkbezCmDchOLhrYk4w4GMbzXlGPIiJU
wOXu3sPdSnX5ZAxILuGKHOFuAsWqy+w98haHp92a0bkqowwyUt4Y2Xn799OAla37
0npdlwuDgP411FTFmHw/Ja6f2MaVTG7U3jPM9rAKUY2e78/2ykJdu+qjvt2ZacAY
l8OgMKrRUojumRj25QiE6Gj2oX7+lM50H6eY67kk4O2zCJ9LmGZ/bTZsbep/zoFy
KdrrLYqjRyUHiV2cgNWlmuy2YAqqJeOdd2ksJGIwE2gxL+c9aVYR+2zPkpXsDdTi
1CTCGBlVRLORXATG1wEpVOM1jPi6pDv0x/KWMKVJka8Dk53TONs7azD5OjwEnsdz
dG/Rp8kJ2hdF5morUtWql5ZWM6sahQgbGC2sFBXcNEZdZtyi484n5WjIRKsaLx0j
CfAHvftiq7krasOK08+OUatpl3sHeA0rpHXduttzDp5F8o3QFn8O6kThcnj9ShSt
/4AXhw7CKuBO5Du4bn8gi+o34xaUXeiYzOe0Jn+occ6wsuu2xkjFpqqiTW4SsHmH
GOY3MYSCMzLAMIwzt9hX06uCsT9vBglRH30MwI6RfO99Ye/UU/xo0OAYDHaXMrdm
fF3UXr8SnihZsJdB2iXPqXI8X/vPnTw5ACTsSvRSdm9nApZvdPEQogmG4D5UZjCJ
RgLLPnZRN46XNqeQWXOg+i1MMiHUfnRLX7UeupQwjE7lWIGrSEVQBDMVT24aOMMR
85eU1HGKd08s5H6N9Bfu7iD1v312Nq4tGnVt907KC2Fo2FdcFEVvmaxXU5AaduaD
MCqlq7eRiW+Gs7Ho5BM8ooEDt4ICaPjjJEOPbnzTg+FspAjrjFYCtXl7WwerykhN
JYkBRMpWhWZZQZSZ8tup2dmcFq9khGg5t+Oheie0jxTbS0KCS8pnBUvcDTh62xk9
4tm5bPM5e9+wo28cQTI4YlulQDzJRadAqBFy4fEBKk1TNJL3cuer5DemtENQYH7w
CIhjQj3EXpXtHngm0KmthLLXF9gZvQKw4sKm8Bc6p4sfRzYgNHkUsFpAa3uHnzTT
8PKKpL17FVDO8be9yDQcCDQh2YaTzUnVlLeqVsmvNXwpQv8fc/sWHxnOqxWf2oHu
I/JOxH6w0AJgRT2ok2J5eZXKe7pBE7zXuRHWcRd20jB5YZd9GdSo8DDQ5Ik0Eit8
x3j/vq1PNIQ/ic69/KYH4wuviJx0983J1U03Vo9y0kQaThU/ARqAc0d+gLnqOX7J
nW5uTtExSKqW2ouygJFKilsJ69GI7FXdbYQABqVDwmt4QBSP8WpsPjhsZe0DiV3t
kUtzw6JvB20i1S2xQQxiRKtrvnpEFgxm3Zp0g/VKGcWbs6H4HcY1MpPDjLdIrNh1
Ss7TjlJEKLL9/OiMmSUmW+9ZNRciI4y2Gvrotn5cAs+a8uRmNiReD5dmyi2kEi7r
YdK2NDIX9rO5BErfh/dXcRuV2Z1Y9g+OGZysees5nWA11OkKNo9Moswwe3mNaH20
30Ix7m8ToFpR/WvtppjteqZHZbhog/28rFG/2aF9gJzUj6E1dhGN4uXFJIoiR+QT
wrIMzGycMDAn09LpAH3toAX33/LP6aoX8/qXy6Y+CgeoKVs1/VUkLjDzwCd96jFP
zhawyDpCQoqNyZGZZA4QHxSK/JbXuI7luIb81F7vNgin8pPV86CKJf/d3n3fkgsw
Kl6dYR2TKITeybHgRO9NP4EQMkIFT60Uo+qRba+z+hUoAn8KMF1g1os3PxmyUYfX
cbjecLpPlwVGTs9fcKa8HP6vSpd2CTqU50KWOwAPBNneUpRsCMHvn5r4RBkqhILP
Ohco6OcUOutlj71hO9HNQbTYySA7q4kF94OG5WYsFGaDM9C3u36p8DxMXF9klTm2
zxDquRbJWKb28bc+thXunqfp4UrVutwwTQ2eYb0x5dK49dwMWXU/o6Q3bf8FrCwp
cBj3zbmv25xr49YbhFP5gqHawPw/8q619AdG6uQkzEWZK5zM1eBYWhu7yHX/zfNm
SwyU612o4UQ5oT2FgkR4K5ixJhzhl16ehsM9D3WUT3haAE6bBzgGIXUrTZcaqLuV
2+aOmgV5WOGjT/iwVOUdK4as0xRvQ5gm09tCWfeuFEVfYfidQZeYDoAS/0np2M4w
JsxHoGSiK/obhBgX9L54Tf/EhMZ2X0M5FYFBSv1t2h652OYIGJ8RSqc189lthpkp
uxYFIofuDA7vgABnRI1WkI0+wyqIw39fh0T6VhCfnKklyW/Qfpja3cni/BUjQ+Yw
BZxeA4ciL0RgL2ZjmcwZGFIDZ6HU/2fqTCL6NgWuBukDdol6MTHV4J3faEB+Nh7j
D0DOHx53oOzGL6m5ZrU/UNELM6jQBBzLlkPIH3FG7evS0B0rdm+TwrZzL2y6m4kV
h0Y8a7pWG/tdTH/yGbAE67gopLHk7bXpNqUSpwpeOHgvqhjIPzRSp8gVyjgRiKYP
DD+fRMuYH2e8DnXJFfH9J2uKiu/UfV3rOBMus1cuxpadzUdeQ414j8AHvoeZraqG
tKqpGDzM97z8CabmKjIciLii2X1pUGDjUgmfKz8/1kG5VhtelC07v9Vs71EAMGH8
BiduHsx9xnBFrFLenTcyFFpvxzr4yEOPW013MarKTr5uN5KTvpjsE1p1a8NRFx+a
8tQm59xnOG5xjus1MIfU1IaMYR1KKzt86IiteWFYbh0eZgoIFmE6tpIYGgu8JnDw
8wzVNBi2Kid2PjQryzftKBihdpUpW44Hh4xOtsc/MH3NW2dd9mPmHaYvujEFE5bp
IOT96FmPBouDxzIYJr5YsyMPVnAJi+e9xTSFjtflsF1sn3XHX6noyk6g2lBuGNlo
vs6HplYwkFXR+uOhus487AjpQCf34miCO+mDmpWyvxhA+81Dx4GWslWxl96FU65n
vW3CD0OewaQZmTAz+Tz4t6C2JRx4Ydrtfk7PheFGp3Sv2EKyYmDeb6MaG8B0yODG
Yf4CJlK4RsHPLtKnN1YZU0eKKpcC5EdxZyd/0l/lttu1/iNo3hOxOQrubC21Dndo
/UCaanrS/xiIxrAveFoU1/KaWq0c7ltrDeewgaWBAnhe28TFQoLY7HjYIikot+Ho
46b4g+Y8o9Eth/NcFEt/Ssx6S67gfRYPg9g6uciZK3co0f4ysvJkcRDVJm3P9jja
NGHXvFdY+vkQHYOZodDjVtg4UrhSVoE6w+wMXK46Dy16F3ntnGD0wz/zURfPwYsW
qPyIlchLIpnq+31JjEmvRimS7iQlRptucnEawrHTYw4FRBUk9WeqO9XOFkRGKPxS
U5R+BgSFwx4Q5PnD5H7K9NZSkmDSA2iA4fpZO9T3K8NIq/hfJ3iDJ8wx9ZUxxgFk
rrjxXuOTrtr5/w6At8y7LLFnohNDlyHia00SlCoVL3gfh5Vs0GEzXcY0s3Ya6PS4
r1zS6+W4+XpPavgw/OWOqEZQaqr1tbx7KU30fGznty/pa3rmshyY8cv8wG5Tl2It
EO9cBn9vYz0bv6UttcIDnESdOhkZeOlKATBfDtqkOmchy3Pyj2xl/0q0MsCQA5KD
bzqcTZpiSLMUND87RWV9RGB+97NB66NZCaNtwgyN/ls7Gw3ZmK4Af/RnNqxZjdgV
6NA9cXpaWiyxQW1w9RriJ2om+MD/atkdAkfkBleLroMcXai6jJsPPuouRuwmi2cX
2+ur4QPDFj3Qmiw0yl7jvwYHswwsi5zuNiCUV3GyGoFpGezwuMmKfeTy9q2V3NCi
D+4AdDhhDEpclF8pO/CwGWJyXfcDcV9+mLfe+wuiyyzyYqkI8lN29etetKccCVeN
xxym9j7LcjSrRQ+PnVy1VMYFN+o3wGFqcMysz8sYGkVGgicOX4sIRpyuFXdOqXyz
ygtk//zNI6RkI4+o2ShhZXsa9uaf1gOBUIpnipT2vJiSYBvhpjHBoE/Cymp6H+7E
5JGoDHXr1E1MIt37Hd9MRL74JDFtKeCl2DChFWXfRnThF/nYooqIGG7jVRV6wxRX
j3jxpkApMk/NtsXjwLeBxyzgErv4+T/eA7ITJPBwiNq4kE1DemOxmHsevJeLTk1p
0YDyTXf0EtdXnDqn/eZzHC3dJbUUEA8Bx3rMukO/ttwt5sJJg9ofAjhkNbaNpSkz
wH3RuW+Gu2//S7ShguMryjMBobWKtNj/mM3bGKdLW1K4idRq2y7EvFfi1MDglRP2
zeF8bE5Uxwvyniv4TFLNhDvADO5rZe7+vdHxcErWcguZygMO30JbjFq1z4+VnbDb
4W34noKAH5tAGpGSZOmYIx2XETx3PeMFRJa2r1LKSvjKEgA2EmBkz+fGKt4ItP8m
7Xpov6TjCswtWziKuBBKe/jjTYUY1sEvFJ09/7EWyOqtRmNWRGG9eaKMT4eX40KU
Lem42zx0eg4hxn9AHDr9RmNwt4YabxAK2++SYcAjgMmhAlnSeANT2CRnUq/42AQN
hhGw7h05T0qtRScF+hXvyw7+FPXwFA0zuM3mpjNaTZHSSUhNZ9opmQaGRe7jNEez
2VBdqQ5u9lWnOHlE4zoB4V8Br+pn5ZudxZInLuRmGxUqJBwUuDsJnbQ+HTO5bSHp
4nHdGM4rLcFr55xaNqeMAJZcfNE+HYe/AYTZXoYcLvgQnsyFUSbirc2udYfStnZD
fHGjVtBngAgvBY6gX0G3rN3Ii+XkJJOwYztPPwfDkxioJ7/34McAMWEvzfMIPCez
vnqgq8BuoZDAS9qfzf6fSYQhZ0lsHwxiMBirpGUVn1Yton3jf1VuQ1WhDdiunolJ
wN6C5xwQj9/6Ogox6Lq2Mb2vj9VFI+K1G+nvEVupCcLJlIeltoBx3dhrt3/R3c3A
FHBvw5quEqOaqLZCqml5cKhUDCjMDH470QGFCGTu0uUGaCxaOJURdINztD/Q5d/L
nHGnei07WLmE2TpdSQLs8YVhCtzF/TeIv0q4BULeHZJExnoHS4KxtGQDKUfPB/ok
GFItzrjgihwV5QbTTIUu50GozW5AZGzJYbFS/xCdwYUk/o0zfxYXyDMVCAmNYnei
jcEuWubijo4POFNASRcVkeVhyooxnr9OsT5pAY3wcIAdZvApgZi3UyDBoYqLKmi3
T71M4sKL1Moccv7iUcE0/BPBJTnrkJ7YkKQOETShsVUs0P/7Fjha7yWGWUYwZle7
4Xr/XPyBfSeQ41OKlEuPjjGKI0W6r5QmaEz8TKeZl0WZ8hjSTNC04o1cHU04IwC2
/Ux+MIemwlrmuVjJj+kdRsXIBIcP0lzRjCwy0tdWpB19eTUA92aD4zG7bbiNOOGq
9SlpYCyE8R+sEd21d1x1xRVNQgMjFSQceMAsb0V7nG/KS1Kfhjd2xtu6y3+ZRK+4
nM59J7sJ/iMUVpE94aM2+5tm9zDpEh6lEYP+bfT6B0LunxBfc10prIbVGZwy5dN9
1yAzK0MoHIAMjItyYdu4h11RlFADENSXQmg29CyFNc59qH9pfCiV8vwTAvJQvuAn
F2O4O+YHYDgw2rgfnTFzGDtyJ3QQVlBogZHzEkVgz5lcCF3SyhIhrqWK2XannUt7
FeItUZ7VzeUnm+UDiTz8z8FQJBFSvtL2OZIZoVSJRfI5OYvw51tDEt3Il82T6JVN
NlBVo4I0g7APqvfCDrPkZG3hQbywC6SXHKglfuTwB3+W6gNUEktzp1yKZeDSJ2Rb
efrx+Uv07lgakxqfzzHPwtwTphmSEWQPSPn9toElSJFBJsPHjdV0YdsIl+iLSdX0
dPDc2JN26JwKPUPOlaTmgT56sRspcaFNdii/gjE+a0PWE+4Q1LGEhZMQ1p/Xr0rB
fYZfPGM9iO2gx534bzZJcpG9zZcQmc52iO40Bk1SNA16SVic62DZp6F6LbUaRxbx
+6HEEGfVs8p8h9zphGi1JeAiWTIvBPzadax73SXeHrrd6XlO4QXdpYtsx8CE1xnn
OKxpoVllY/0SubvDoVKOkRSFLO2vMq6WusGld06IjGY68NoDcmfMvi9/jwK9R+F/
hE3sWbP26Qe9SnVWF6tFpdpcnBUqpCrw/I7Q4XpH1RLorHPKPfCmDPb1b1X77rvL
h8W0kiHjwl8z4Gya+5CP+ZpwsPrcrF2pwuIoSgmzMPj4YyKPjVoZrzEKhKQt2r9D
AB/hBe9RjzHiWe94GVRDOW27cfxGxB6eXsG25nMg1oMRUnvLhnfxBQvOxlFzLavC
eb8CLdfzQ4Xvu+XkmBFZUPRPjYpQGfY8gaxZmMK8hlzMkV74bMy66ButNEwVZGuU
/dr8YrZ1//zfb93yNOAFSbR+yP9kn9fBpoAr+T/4OcOAkwQpAT2deqqG8LTAA21x
2t3l8ar0XbQ0cAbv4FH7QCJMparRLm2dUHJraqEuQ3zUgvMJXS4XRrFMtTGJSMa3
QqVt4wfRHhP3t8bhQKCoEuaVR6i27LV/on0NGaDd3Fw10IqhZuaix7Mdwf/6/50f
IlNB30HQlrWXMidqshtQS3ECE9L7fmAk4cbmomCC5qqGOQmOS0+BxptE3+WJ62Ar
jqbnEUrEDqpqlnvdSYs6RLz+gBkKwwaq/AtaW3mOrW/YXaSE/wwkikD5ApCi8Qyj
bQDqlxMv0KYA2NmFnoEj8rxhoXaok/wZXhiuvsns1kSkuvxF4JGBm5ApR4tZZatB
RQIDLE9zxZKr3blhNwPHzGmqaVDJhsrdzpXnMPp/0l8rHXCzOkTkfhApZw3BOw8O
Dr2u5CZrgcLd2/QikFLlqwRkgeCO+aoYeSGoOd/Pn1as6fBfZPwaB0uPYXrT18oc
sgnaI+AcdS9/w38EIZipZWQIaIw3ckr4cTTdadcbfh7voLyVaHcHclQEmqYAsv8C
RgTfpm9iqLi1RH487xdVzSubWL+8o/wlogydGDpnSbDE1QR6c8LLazbYkhcACaO1
/Wif+Uu5rIp17ps2kmOkqrJjRLJRNMNYUTywnHAjHUp0tOYHJf/HNYNfkkf7ocbo
/oUHQT3mJXbc46081S3fWrH/T6v72Qe2/1q5PoXNLcs50KCY0eA1EGiTcnH3+tf2
oQc1xOnZv9JJLatcSAEsb74iLJ3SAsEdmbdm5G73uZJdi0v5OnHHHM56kuBFWUoH
MkVlSnobjo8Gefr5yaPVB4aNJVp7kRC4lwyY0VqAV1W0HC0KAICeEqjd9576RnkJ
RSGh/mhe5u/BCD8XSPGUjXrnB3gdy7po9IPWpqPQrAV3emAfL1P/bXx+seRxAF5L
Of1pEu8pq1D+ODb3iWqvC88rGrr7Hz5azqHKg7Afz/uN7h0CfTW8SVzPzhl05dMG
PVC18ngAQ5Ag4n40pqoBprFk6XPRqGTRLFm98P3UJNXYfI7c+sF7AxBeZToPDBhq
uKuwQanzNa/Ka47SKENtJfGBS2Fcgz57ceeNl7HouULT+TeoqScLi0BtsCz3mhWl
3BatHjBGQ92OjHAuakVyXx5bLuhcvUAdV1KYXkXmExAijSjEQoAU4Wu7oOe7LBam
g6BAUvbeM+wjpGNzVeytXtrwyEXlZBkYeKImzJ1vXltgOSioM9cA2/Mk759JpRTR
FQbZJ+COdWKEmsa0h134RUuOxbCKjCAJ8xDfXoqDmfje4vpMf+LHz+przhptN388
kbRN/HBCMehNwSKuS/OOVmyYRzmqlVgkrwmHU1CcLjhYPOqXbnji02ctob0/EWK+
/SrDGRvJwLaivxBbX6lUHFrhxomjARbVJ1Je9T+5rqmlghS6YaqM8RQ+I9lmRrHu
PHRglZwlPdxtAv9ZYOesOBisMZZ9NsNvAbGmXcWM+O4zygd6Q44kMbVBNzm9HpUV
EFbMeMRPQZI1ntn84o6pGnGpO9rNUMusRFnxf1fGx3k58y2K/xV9qvCxCOK9YgoU
kHxMnKkQEs0zwfEQXp+vqN0VZRQFF7+uwGWW0/vLrtPuszq7c6Azp6TZK6JQfTWM
O2c47dq7w6Q1TUXLXPp9V43b09cGwL4DKaFi1eAqZJI+AyDY4EfPSP7WhGANryea
TyJGJSGzS9Cd3yoIXH6q18WWc+MEYInSFqaUPdaiIj8G3QjWdTWsQ0posoQiEv9s
2auD9y5vmnYb21CjR+tjCvcTZBQuCuuV+UVDAMqYe/RgS8DtmVIFfgO9VaTsTDFm
aVEaAIc/VKYEIDtaMm/jpCxdxM6yuT3Eau8feYerf7V1XXxw60zVxRFnbZoOBYR0
pdjqgXni62EATwyUn9Ym8GG9s7Ml+PSGl4BgjTZE4VPV2i3mJopNIrvqQwZiiFwK
5ShtwVoYySqyLaWaN7TiEyKy4EiiET5kHnf0MAJ7HApAkHZSCsmcMn8sqQxH3TJC
AyAe/e94hvX9ZtTeqChatwAQLVgLg8ChSu6EC4tp36DRpkpCI4u4o6yJyOy1c9K3
vmDW9pOHX4J9q+2oz5hdBGJBPFvAWyWUHoxoaSakNGGlIAxsUDwr/hHzRzDzwfXr
SVA13ZUqtHZn+Q2uP662eznM+Vv4ym+4cCsSZguxFeT5CzuQemvSQaY/0ZZtvmV9
t2wf500OGEEk2Bwre7iPwmcy53b1volfZz6X6Z7bb0ksVw74Jj2rjP+5doUnoWHd
RDDA9VV6Z8Zqv7pbsyt/5BW5G/K/hK4QzFy3PZbUTz9hMoP/cdj4ZoNvO/KkWCPM
TAAdS/qRhV9/hQ8cwhc8zNr1sKuy4EAcGsKaHKQP9cW/UA3gxiEh3r9NedH5/gqX
3HLpZjLWh3AdXv3BKDnUllaqKInRigtrznazPD54an3htwtIWPgilMzJWHLRKRqb
BH4aca13hVI20h1Ce5NWmg9zBsT6/ojIgz9iz3pJ0SQ9ClA4t9H35hVEeJGHHp/1
hMVuyVUd3gUxZ3lGlLceh/C7UCjp28s8M/HqEKjwWOk0TSUqrTTFW+qBZ/tXzA+F
gsj9wRkjW80sUOQyrMEQssUK/fAS4g0n1dqJ5lh3Ptw865/Ly3OnFfPStqLM8mP0
42O9fpNNsDL+TilK2/5Eb73QWT19NzQHBSCt0NMIMsjtheTBTDAYCO7Ef1qn0bC0
MDZAZuImFdDKAjXFl9RT4P/l2uCfSEUDymsGrGi2TsLtzJR3ZoOJbnklqsyvxFBI
V5WCGrZb/DxiwU1U1KmSlIeXZztwjtbnowJ1V+pUQwGmnPHjWKS37QQROIa6zSs6
Ytc9xzcrErEIz2JA+vY46piBI5CULtdRILEYcpLBfR8ABR7q6cXVwjiVigP6F5/Z
RgtdvdmXoro8rCNgD3E4+ZS/dg1tPTCrEciG4F96NWarim7igmSOKme1axHoZuvo
Y838dgdobMghY9S3sDnYzlFHp9/rADMURK3/0QE7vt5jHvHiL1C7rlUWvnMkyVJj
kJhc1ZqlF3/y0mWXOvaWw97G/Vs03oIn3STr5fJdwEGGLwRVYtzgrfB2qhK3NWJ0
2qoZCL0GRoLdQyAaDMlUFOJVJ/v/W2IQaDzG9uD5YGBtBCeRvc6lvmWaJzLvlGzH
oWCxZa+AtUaKytau5R0UtdX5N5WHGQubgTtXQx3y0uAcW+2JTv/xqqbjuiaTnhBi
chLBFPLLtu0f5EKJoISlfCG0tzVgyt91RV14wHezHxqC5g3YKYI46XYs0XwN/8Uo
IX4dyVYNBBGCPN8MFoJFjnESLoF4QXggS0/na36Hs4T8pVuQbk33kHsqYaK0wD43
cE5Rs0jnzlQ60d7keGAYuI6h8gP00BmiN4IEO1+sb8HyVxhLSB4Kk3CW8bWksU2F
SBlZfzQO1V/AVdg0INcI6ubwDUYCl9XrIqCJK8JvmZxUrOc5IvhFU0XM1xM1wLKj
qJ4bJz+hr0LzMpyRSH03eiEOpqoQyCqOB+FWEN3lQzCLqcTNvPkPevNByKp/ibTB
aEbLtLiSQLE3XMza/cK+OoAFnmGlH2SV0M+kDm22v4TlA88VIMf7SQUY3z/VkEiv
aqvA53QtrACn8gOcTI2l9V9g/1YpQuNEz7RfHWIH8M9yqULRbViZ42DODOoKP/Cy
lk6QrqCPu9PS2g7SW7eWRJTxwRvmZTk8JYuv0DOD9MtzQHCqAKKrL6e/4YXtTg6h
/nAcM7wzyGsgMxPo/X6zgCIKJ0ukX3e4cDRhCxBbXnvIJMgqM1sPKnu0OvHqaxkW
IR4kBzuvuURnvtWqrRstBFFIH5lgLZo4HYRUBk5/oDOl+TI0TeUPIpNkpoMBmB5E
0pYM8u0NOoHoHILX4xLOphC+8QH4YQSYgsM3dm7hWfddyk2mFBGmx86wSyje+Aja
8A+/IjRL41izC5AF5ci78f829z+ZhrY/Lt2UI1TWZgxm0Z1i/gLJ73dNSOm4FZGV
Lvtb+sPBAb7+EekQOgG09jSTEw+tneB67dqotMBqI5U5G50LbSslVcfpxGbgBKDV
IFCK9IUsPNa6kTUEoMZj5db9sglLV+fMtZRjyrbAwmo05/jtZWuc/J/GKkhwoxS0
l5h74bOhdbtBGzmyw5M5lehzj0XifG4owtFpWcdQ1Cn1Ed+K3hR4sq2dWHLdARRn
Hmi39ccje0T//lVxz262FS3Bqwd33oXsmm6skx/nvu7/jGwmloHniMPt7QOkDeVt
xdmu87nMMK805CGIhVRAP4CDM0oMG9Obn1lujOnqiG1t3t9uB3tWHHo8b/JaKGVk
UCCsiCyLpTr1OSqJAjg/Yo0u0P1fKjUYk4gdF+C4Q8/x0IZG9G+MmZNDy3Z+mlbl
IJ55Zwn2syCvevZEEYqB5QB5f4+CMm/B5fd//s0dFLZuFFB72FR6PAVv/m1EZKMg
S37cO1+tmkrwYODoPF3wqdKSJiXrt9UNfhSBPngtOhW92SRFpJYzi44b1nlEmqWG
Sv4IWdt9AMwrE08K+Rjvu3WtUGFi4lBc1sxnTF8uAjeeRXiwVzt7ylYu2qi6QF/x
flk4ps2N1f1C0z5sdYCbGUrBzUGqT5atkL68lLxprgl8qwKRZgNUu7hIv/lxZ5Zu
Qgni8nFPZEUTZVQXURKQ/PsoP5QlgjT9GNz3Fcop258TcFY6zXUV6B2sXkfqIw7N
cWKsvZlKGs0084lY/K6s7gHdiW+xettDA6F0xyGc1nwZe7ushowiVjmNntpUobsn
IYHUMU0SF3qy9EGAMZR2anxPvX66Hbtt/LkDOZt1MSE9Fb+3XrRHBBkFIW0XdkrK
/IVDU4eLzYhnSnoxYRFkic/8isCRcAVOpfzXEgWJRChWhR+NQERqkR/qm0S+KXr1
p/4WOnXGyokqInaJNp7X6PcDK9VwWBLHygLQBNTDuBILEOrkZB82xjb3t01pOTWB
Hhkz8iGQ8G8cjz0usw+7MKQR+ucAoH9jpiXqykJE9MugEeUVCerISZwR2/A9RUMn
ztFtPChSMHga7J41wTDxHBMZtErDU1QJB6tAlAeEhRys5UwV+9ZyMnwMgfRf5ucq
LUebFVPSDZ0KLo0hykVhpt7opCXGk/aMHlUTLPilL0EfwnsHN9bZYk1jM4Gkc8TH
i4Gj0z76MvV8uMbBz4qcNJxWmxCwZXu1p9t1pm2OkfY87M/EOhAN4MgVN26FxxJn
onJYHrEoY7a81TXGyxRMbYFZGywbTqrjt7ijhh7qZ9DG7o1qFNYfXtJ8ftuvAXQS
le2y2hy2a0RW7hxOs2d7cIhZqkDD6jiMASt9tC+P6varI4cZHMqRCD+oZprnKut5
NdY5gdL/QpLE+uP+BAid8x19TW4fDWLo9eqVFn+Lo4nQKHs8cYVEJAbh3pPqIB4E
bQndxnDD6QwDGvgp071/f0Cs4iyHezlLakzcJVAr4RnWDXJiXOPJ2gWeRM3/LDmE
pxjs7j2N1HxXH8wHDKYF597qkastfqcuDrJxONELPlUsa1pTRpgkENy3zrlmPjIR
tHk4SfEXyAeHTv02dD0EZWIPwengOhnuW16Sw8mGppvH8gm7IHRZLWuxui3Wsfrz
vOA4i8qFu4IHHtImdJK3SiiMTvZ7DjlFqYhPmGq/Rbwz9/ep7cvzqh7E8UrkUWtg
siyX59mKOpaLnceBAw+f+Q2+H+W6nMmYoBdUv4KSt/K0QeTy5mWAuwo7VEJeWEhg
puq9hl/Qpq/0asuUNX34KohTUL0sXkO8qhQbz8ZuuInYtDIkmgirv3EOf+DPkmTf
V/U79Hri1VECO0Kl9eQKFvKwrLvDlUhG8X20rNYGyB+dCLemLhvJ+elKoGtMDJnA
oaArEEm3ex8vuxNwvoa409XUcbgtYCZKznas6CKQWv1INfwe+kxa905koAQtyT1l
x4vE8j4K16it//xhugqr0jrxENPhSpRYnrXmsN0SGIfLHb00qWZg2w5YlK0gX3dT
kOr2jIvl97rag5XIJb6v/4VxGnOR2kOmFCcMFu8E4pCpV+7XyEUxGcVupYiLHUt6
Pia/vvsr7bla8Z0ObH6L+NoR3ls0CV91lOC1/8J94XiQwnBQIrPBmd8QKMVTMcg3
l3bnEpKPjdcm4p50MqHruoPQCnU7M+YSEzpCndq5ekGeULJbvJsQFQImJHsIvJph
IVlG9EjIwOxBpvEEPUL0+UEvadVUjI8WHxSmZznwKU0j0znQ6ETHCpghg/kSEQlN
Gk5K+6EcPWQ4xdyDD6iSo40v6RwfLPD0WrLrTglC82NsIxQhKXv0l3WEKkbme6J2
1cHAm5Tj1E4jwGy/1ZTjfIiUeOt2irpCE5ZZZH6BNmYzcRgr+P8nCPm9CV5isoBO
7EKm2CX8ixT3AJBOo0IUmYV4dBm+rEFakx7Gh4EGEk/ORp3aVMxS+5dGQxflB+lP
0pGV7vjlSZ7ozDl3Ydl+Dl3OhgXN0DDiJXDGjHQxDbgZX6bXibKkyEJHVYAE5x8w
YEjgopikw6ETz4WGm3qAycsz1rU65lowJnMINUqIlFzjUPqZqYCXk9fOBkmZ9jAj
HJ0QkVA8+07wPttyNvmhIFL8dbp2gWlh1T3BttLkxoHkIKtrgcANA4Dym/perhJn
6CnWaNTcUFYrQRMuvs/SDBHEehkx1KCUp2aCXtVBo6EggwX/XwGp6Ucc18sFMuVk
GPamCKo9pVy/iXzv24e5EHrel1oiclC1zBasqEoECPOawVbBck2g6nMbh9x7ec2N
KfylV9oQ3V1zrRGQjoHLJVnGW1Kc2rXIT76JodFVvq0gUL//v1t1IP1wrvh/fSnM
H/fCKzEOLgOWbk5fEHMIanxQwLttG/t8Gpm6b8LbvyGofZ7fGUBNe3DBA0neetRR
lGvO9j8y3CIwccYD1qIJw0jmrjvG+fCHbupt7mX8hWtKNaNg1O1WesB/s2xh1wfb
YXVgH+vn/fOn8GrUjbkKlpNjuS0Zk0Y2XIeUln63D+vs76QAduaBnlCXc4kJMY0h
vFAAScws6f0xZSEoVBMkRat1sz3MOT7EhBpNLg1n0vea7255hE2AhrqPFjvOnf4R
H9zUcy6O4uimdkT5c1NZSx9BhfXLbpLGWyNAb0caBMXf+4vFoG/Nj9OekW4VgAgb
QwxSnYHgBeTnvyqm5JDhdEhtcDSZfXjWY7T2XDl84zJhZrhKjjSgvc6ziOzIhmS1
BjHZDCBwq49ogHKcrqlJF/OeUJ09+CIQ1LB8e2svuOB3s4VOiEj/jZgRPzdNNZr3
P+ydCe7cepFlT7FETVJs2OR0SIRhZmoD6FR45PJMITWWmTvp+J6CmA0hiBDHA5aL
G+ZvV2IxD3d1cwDIe+bfPqHItBxryDDRhLtSH/taIGqDwS8d0UcCpgmZ5dISRtQ6
m33n68DGp2D6Zjf/4vO6xIjc3pTGVlzRY2sTH5ehqkJi/U9GMIWP070ORfIRCy0y
2R2hK+J9RKZaZKG7oX8hjBgKVI0cgrtodsiVirJEQnttUpm5WbXvQzZfLgBoJKjQ
3mfjLofelJF1W0XX1fJT0+5sN1CbTJfjQwBD9ROgiYBkpZ3SGW5sb4ZUfekTgVrU
CEWkHjCcbJuhq5H4YKbY2FvITQok1uNJH51L6Ca4bxvDxPkTazl2/ReVEAUdu0FI
kmJBUakBehJqjpNDLNmLt6/TG/Dd5Op3D4Gi76ph6psHOY4UgjRvH3U63UQrwlb2
MgEsPcKPguCn6vpnfF1ri+yaruncE+bXHL/kmdU/7DB87CvdDKex/ZtL488Mmv/G
06dgwSRktKCffA7ysVBu8jxglyQCa8CF5QXsO88R3NunB64yMo6dN4d6x31bUT3Z
ENhJJtsNAOauPxLnAk4hYZ8LmMBhVPObFrNr0WUH7WEoJOWWcLMZ+aSA6leyyHfw
jlMZ1C4d20mqyoL8grvCrueBlPOCbdTKVsw8/eotLryAtUxge6oUBS2e9sWc9fE8
Tlx1puOMyxT1y34ly5124KBujf+7+pvZ1YCY+z858sD891WnyXZZHwiIbDRJHlXV
guDcritVoETnhz7/jYZpvNDsaMExJvRlUNxqfYDmcxkD0bHjswVZILqF45x8DuWk
jLfNU1+1jlNK8E4kSTfIuWb/xNOqET4Q0tGHeDvs72+DZ9/kqb+oD9a1WNBnU68k
KTu51Sv0+Dwxuoz0kDh6jvninTysu3ZQaDxApRrkiRNQd4O8shMzo4s/IyxF0hWH
Cjwa3uDZ22gp4vcJH4ZD78aITgM6JXgf9GqoFfD246nw0MMoOr8RKSv76R99Qu/X
0YogVmJTnsjrO/M1jvQgS2bA4plKsp9tPyycWWfusrx1bLH3VE57PB5oWEayOazF
SkDqy65z1/Dqz2p/qLfqwXnFm38dnk8NVtb94JZA4/nWcYK7aIywdsQdumT5T4Op
kfYkOTWII/cDUs1An8lt3EZh1a860Rl3OHCoIzdzxk3vs7T6/s3b7BlyUbaLJIyb
WFuPlb3QrD7rdpbWh05oC8veCvle2/oLrIiid2P3k17nh9aMmZGO0/E0fI05EB20
+cv9LWXQfs+v0NYeQiTcKPUHvlV34D6/vRgu7uu10IGu2D92KZXSBiSq3ilQwdZ1
kWC7MwpXxoj8WWw2Q/bZCuPkohwikzUJEc20dyYqoXNZ2Z+xOUpFbq3sxaRIp3eu
3zP5bUBfkMpj8jNFDZW0TkkihgxxEKjeHf36QiHlyJ3tH7qVXV6ATDghveZLj0Yf
fzTC0I2EwE4EPmsFa1WkA64FTcXJmdIV7oAbGQNcdq8fBiCY59ymxWF812X1UX8U
m9UpBCIM6/YEsaOmq59BugCU1KRzau0iW/ogL9vuWEuh/QRwI5Y/7B/yfVac6XCK
uN/PEy8yJI32En179rQuOgwUbxWvexC8JKEa6JOwZ5QMDQZjzeMyJLkaN6lokAth
aop2FO4R/8vpGPRvse/dFH1uUncu8PEFe7TeBcWBMjv5v8dOkqENcG0GckaFKxd3
Ub+bGb1Rdvzi0HvKPqhx0lnsOemnYwBoHl3x/H/LoRjSdnnqk7LSDspUVwTseP/Z
jmUCOzc3SOud2IwtQZSJR8+nVmRqLyaSWV56yJlnJR+K2OSDaBeIVcYjObmS1cAF
vC05Wd+so7SLYJfBBtC9kl2OL2FlgPG3M7aS0PmpYiB3qjym66reibI3BSZ2WzwD
UMhfoiAVOj/09kTgzkmEr++aLhze9/5QUfnbG8m4130mx3xCDC5D+obgBJWnJvrv
3SZqQcy8BR9lAHfBbm4NxvrU/T+MbGG4kdeJueuRLmsL2AD5PPwJLsBp1tKSm7yM
ia+GPUL9x6Nj4HCegpvVnek98cKBwKbbEY+CpV1PwrbM2SoGcds5odN/gqja+WUb
76sEM4crXVrUM/V8ULPwgBCO2FXaNs8M8PIZlfokfAQNVrfS2TsL/CDlZ96Hu+3h
q2e9nJ+7qh5gjAah+VUvFpdb98iR8RpVFtZ0ows6djpkopJjYRZHIILZcw48QjSq
u/0I8F8wWtsa+2WV1D3ZAom4wfhDKMGQgsrEDF3vjSnqWsoFySgjd3NAbuK+Wqfb
pwrRA83JUZ21m73q9OASHXJMekjvJZAyl9wSkhdxGO8DHNYc1Ug+9+feEQSMV6zE
bEM/HgAsUB9dLQL4hs/vxlxIxav5As7i078GwZuNP93005FyqhWM/1iIYw9lFXjD
OPCBPt9SptM2lyv7ERdyJu6qIemr8bRWvRxS9lwPPp9J2cO7KEZ5/way41UeDbe4
I7kExpFhJ43qMjyXC9AmLPflhuMcRzod8UVdH2cVmWAiTYTNp9cL9P2Q5yneIQ4s
xOlVYevnA0phGE0sPsD+bc6E7/o21Vw+TXcDZf9WM9ZJPJlYsB2l+jq0HU2M7ALf
BzlIOmHHFLcB4DsqYNsUgR/iYMLt4MMAG17r+CCG0b0FaEmSBuk18T7NOsJH7kba
5Y6q7TWjhPdQxQEkF4wljpF5lT3p4SXAtwLikYJ6xNINbztjiEmBKFT5kN1O7c5T
06PUhv6dWzGm3tjjrbV8xJ/M3lJuHnAQJY/whBFL5BisIc4zSTRdl7FCuNG9ZHys
o1AMub5Bjk4mmUJEZeFpwrK8CysrqZVH7LHTrHuhx9R97JXVkR0UipRMq5q24q+L
QfVhJ9vHTlnhYRWY5/KLro/+arMcKKPjf6kKATJJ8xv4UJlupq3b+/3UMo2RqBEn
49irfXNt3Y9IpC3gqVeV0eHk3NE7pl1SE09xEDWKs+sjw4V+yx45+tlrlqm6J0FQ
1mMHKkkj7pIoMa/oczY2S8jVgkSOlk//hl+rc89dUIwZHL7+JkPA8V4IHy3pt4Wb
B7fV7kueHylChV64My7JFzRHCQAj11ol4jMz1W1CTCtoZ3HlDrplE2L8CKAXDkQr
h8kKADZFf8OTPEdDgB2d7fq7j/XkZp/TM7rtUODvNLV+pOcnqo/z4wK0aBJ0L/H4
sDM5El6H3cZ8zQCEcwjaZoMhZH2biGllIyolWM4TWGuumvm/OxXFO/WddoOu82KO
tqsu83uWuovPu1wuQ+FmrQvQOv1wEE9JThhANixNDegx38E43oyvrCqTmYt2xkF9
9vrBKQ0Br5my5EoxbxGxOX2BYaeRY8xI4kAZpUodyeGGjijyQ4oqFu64EBREGpOz
dZyspsEQ+ECSnhtT/dG6GzuSduwjj2B2mJo77aGWiZCa/LpZQ4dHEg2+GBUPeydT
qI2kLKTj0y53CZvu7KHDZmRqpLZQvZp9enPg+s0/5lVWiMEp8qWCQiNcPt/0F1nR
i/Wo8EXs3yoH76oUKzSKHkiLh6tjEfBRz2PVJNkVPVO8w7UE6kLzwd/L39GNn9Fb
dfpEtNSpFDcnjLiVAHLbwEe2JhEdAEM5hr0gNgyTId7jsxHKOhbW5KP/FY0q28Zz
b/wZRZjBY1ezrKGqNAhmg7eP9IQLjSAg/4pWSLLJjqUqiypH31wpjavwTNq4Oikb
LGzxpWp1Rs6kHZF3IqPjV2Yjfw1d2JCLl3Ynakb+AGshM3cgukIwhmZd0GtirImP
y576Fla1aR0agxwiBzg7HS6sH0uTQV6zMXRCO0eZAeiGQWdmP+fHCKe0ITqDx5pM
lGZTYC1gEYW/mqjbGhTd5WTCUgpsJWkW8ruGvkwfhy0AWkTVvUB8L6moafUfFRe1
r0NJ/usBxsnUv29676PEB0R6CzCKP5APXDdmbdXUbaxrRvUUMYkqXM9aCkXHnvux
F687dTjqWvDGpM22qhJikc9qBnb/iqgEMfk4xSI/APTdGcEpnH+f1CU+efybqA5q
7ahQ2I6K2oPGjNmKDxhX14dCklGZORdVmgaNpGvm753cN3UO3axfMEF9d60hp+ts
NOX0QMgMmC9s0ZmG5dEzU5qU+5xosGPITMVS0qCtw5oMgNBH78InsTFzMFAe0hax
emTWFt91cgymAr7rdW2BA4fIP+Q8A7ba3uC0o85qMmO7jBwOTDAveTo9ow/h3Awj
GLf0wAr8ItbRob3VIdAv25YTnnnUNStaQeKgtYKv3E62EC6JCJ/JzfZh7bcPqHip
L6VgjqfDXavvFDTTYGcUNk9kuj5Df+u/u8sEevApXuuM7n1jWhin1+qGX40bsrnP
Xsdg+7INTx4Rf457G+IQAxCOMZKVgqlDEIoOCJlOFauIAeMgTZE2xpCyGiLsl+Hb
YQrXMFX5tL70R7qla4beUq0zEs2tEyCmBdZHGA5AQ9uyZWoMN7qP4deKbl/hwTIh
4HWXbohtseL3vixADwcxevk3cn8DGDc6djm+0pVL8XFHkdoNKwaOnKcYiLsufVt3
TPgJxDKxFIc9sPJfFeHDX/hqj85G+/BCZFbyTNU3npSO6bS1lm2p49IAW7D7Jqe4
iQUuOJM2u46AdgVurNz8h/J+1+Bwyp14jHf0PkyzAu6JEcxrDoBIKH8R1itmLhbq
ymhLp5AlyWXg1sclhcFMpaPB+M6HnK3DWo63PxMtXL3C3kaLFevmu5pON/C7JFX0
/yqG0z871gr1w2pNS2TQvDYvhpSflxwOihPSJHR8u6K0YmslBE3IEih/1yME09OS
/Pr3XODZjfGp/mTHftmcQYk6wKS5z3u24Hs8GV5w9j8XZgHWmk+wCWCrheT8FGMk
eVEOm0Vdikq6YQfRFcH27CcRK7ofIF/ciDjOup1r1RVvgFdryaIQ2Q//IRZ9ZWxI
cz0ZrnjTNMC2zv+aQZuAEpIiecO4araOfeLXdWlQukSKMj9mOP7+koFw/ALCEI02
eG2J9mefkyq38UjdHOp6baMoAdbQkGFbV2f3R8ULSt4adn0sgmgJKizAtKdPGxQX
Wu9N2qOWCAiWULGLdB1/3OmaiI5judsXgYp2K5R6dsYHJcobPohARNJiboKGi1ZA
DQfybFnDxrQsQ6U8M+UVDFEFP4BGmpFKeYlFjRoZbpO1rZ1Oj2Mod7Vod8FuS73B
DO6bOir1qb8YWBqaazaxBfa96U48J3I2oAkRZGC9o2VpG7ztJdM+IZtYmPBGUIXr
ELjKB9l56+NeXZ9x1ZNr7WytQ6+4d4IzXLKyx3MH71/8LN+/+bCGyySBaRK80vQV
X4+VVNPdculMUvuVA1mGw0tDmrcU82xhJ8WIlx4BujYW8rUbR4DyyomN5P9Fxsjx
rrGbbtaefZv5DGc8ZbBEsl9biGFZD6Y+aXVBEq8IoyqBudMD/XPoHY+eSXVrJ+qC
zI+i7Ieo4hwtoCc0dVA/xFmb5GB6mrHb21j2/ueurdVHx+TBji+YJTq6PGnPYwDe
PtP7Y+g/BWsU+El95y7YC3w+1X/6G4ztBm2FS4efHrOSXWyRnoui2Y1YYH+0jDm6
7718NV9OqhHEkY86HMcZnD5T8dutfmXSAO+k8w1NJ+FZlvy1Hh0JQRiX5jZrtwwb
A7Irpq861jW11hk6JElrN7naNW30jc4hvb/SwSF51YJxO8ah6RjTOddzSRyjMD7w
Z2P4Hx5G2aL993KoTNiiemTtJBM2OQ3iI2098RlAiekKT0kjm9fTRZV+1nkx6lzN
fS2NXX7AYY5nUOujjXjBX/tsfMqjKeciFP3nu4rvCV9em/ye+eTPObuGBSn6K9Un
70JhvN0UhFEZVRaK8y6ELeeLzIUpg8kL+zXWJNcwyFTVBFKzPyxEqFnMaxtnykFj
M9RrLSBlqJisik9W25MVDrXKhzoR6h5gJZUvCUKxSWEqCl39SB7rYPduYJrJKuAa
ucP9Qi5bBBVoP1VBQDZJOIJ2IOfoCQtGLMEJwnSTc8hjxGWDpNo2SwhEDj8zWM+W
KF6n4WbFI7Q0NJOomXc+scChMDcNKDJ6jhPihlFQJNBEBxT72guZ9fltUcvV1EPU
vqyOQGFQ5W1xKFt2xFvU/MqUwO2CuAslkvFnfEohFLZ0pJRPvROTpNSrUJURo1eq
xK48iPsFcA0Zy5t54MO7AgpwS+44qg5Gsyk06rQa0gM7FEBC9mtHnLOmy3/0mDGa
xYhiSLSLx/ERPlTy+K3VctpCmttKnDo47nv/oJRP2jMprLuzLaZMtKVlf0xeY/1W
fUYPmBI05uWI/KYWqCZSU1iPrEQgZ4Fa2ZdyFtymbWXyl+1joh2EH3kLPOSxuIcu
Ry9zW6uAp1Tzj3AzNlfAwXndUugjuxAzyLrqmRzTMy3KbXycdGaHPtjMAUVCbn+L
xexNrbDRPygKSS9YR6j4DfXlV+UXXwKtQF8Dt5R2+U6GfzpF8MbSxiej5yPqoC8h
WvPRZ984tUhDqEQUCOKPkkPw3jI5uj9ShyLJwbhtvJL4PJCIgZcuMkMc6ScBnpN3
Wzi+yFTNSlFOnRTF438yiwKA88GCmFXgO1PXO85fthOFcAYI4qe4xhcxyyBjfBVh
zxKMuXjra1Zd1fre90nX9+bJMq/Qt+GSD4ykei9G60b/lrQioWKFeytP7wgncI3O
nIx3dbhK/0ejK9R3HwZfmT+h5nLjPZ74UzqATmspHjAz6frDJ7V9p6D/aOebBDip
60vgJiWeA2AfJb4jqQ/c6LegeCbj1z8W8OqYcEdc4gip/cjzcGf5u0FsigBrCN1W
mdzkYw2PmB/PmQvIzKeMG1uZg9v3BR62qEvOeoTdTwLF37nmGFJ67E+LOaTfav63
HeTcuo1XiRFrUtxMX2qbEeOZfJqFOgUCflgoJjlrTB6lZWnnnrWTHQNiQJ0Hu6pi
9I7PO/QUHwBMsP7pXYzNX7nUFTdNaD28ExffavIvUTz9f18Az9G4i08GAiu+IEN+
swprJt72sI/NSCN+1npQL4YlTITOR6ijqbBAt8CjA5H2jcmTFhFtUZngUciZQpwd
k39dIrNXUwpnyTjudDOdYVM+C20AtDss7GWZJTr7qAfh7ZBpiAk8gBtmzCBEJS7/
5q/qdD14XAMeePq8SrRYTVcPWeGt0tQ/rETo3A7Qp9GZaePg62r30EKws8W5tuto
QlvnC66i2ZbsOTcNFk9pXj+hJZmLYRp3CmpEYwfjiQmCommk6h23IY0XoIEHnAwL
GEFTjx9j06Mq0Fi7ZyB19klSNq5qsFpnd73TtCs7lgJNBLPc0vMFH3s3kJJjUoIC
wb6h22fCm0eZIokRSP58gr81KNZtCIsXJaKuwmeaDZv+uXwOGi96SlB1TC4VZxq4
Ts6o85kElpwB414GP+zuLGF7n/YCsAKpW8uAWRpPoyhD/AhpWxAHbr5TjRSw8ZXN
fMkNRTYI7ypTkSEhGuo3u6svgbV7lO0U3WYyyPWaNGoQCyq+QHjRH745yvBH00yo
un/31cpw+e5Z2NLc0dAdgHJ8+s8ZMIUVHcxMRpTcLtUaMCYYAoLOB7SKwzhR/Rs7
DuxPPIUM835lfaYgoam5kkMz3ycgEEAxlGnfT9EgPrWjmFyYO6rRcZAuvcZcp2oR
vyhQUjWPYBKyh3osc50KUedoycVe4GH4LqV2zpOeJLXVJmU3ARBFN8w+PpVNvNrW
9Q/PnYeo27A04gnrdKe54+zLQeYITUe2031wBvLv10q8qcrc32G3Szj/RyUgGNv+
K1OIY2FZ4Jj5UMdTc83yGXPqA5GL/YQ3+kYEGw6Xha65INn16/LAoiR+jDhQSyJy
Ge9GLzzSrGh73h3KuFeZPThnRyeCc4UsQEkxPmlBKopTimPvtKVxXjJ3fOjx/BS6
maTCJF0yO+GBaGZZyceSYtZh8EE0xsJ53Agr7ddv/3l21dpyaJJ5V1RTR+zOyr+2
yq2nsoOozwFOg+weRjB63anHNrNHDrLgite1NOOMaVy9mloWk5dBsI2EMlQDF2AU
Y+bRpP/WeT9jaLpy1ibNbGkKPoCgHjPUkHnKIM1B0QgXNhT8cm941l6nzFZr6UJJ
oFkWc2CEoXx3h62TQQ+N8B4fnj/jHHLmkP+p+eRPgvsHTwxIaoY8J//zNnONC4kd
iHvYUEnMHeH0zgT0/CQUaoO+8PMSNl6iF6WGL8U9oq3w3nRt9V5V9iiardEjDZ/A
6YW5sNHq/Vx6G1YjvAHVjCHRl5RC9xDtoxKPylWm75Qhpg/DzmAcBSfl7g7qLW/d
tLlkl2HFB/c6alp26QOXK8dFFtw7Bu8cDBy1guBJT3eIOiEZWtSoWIFFfAWFVQZu
fv24TsvJP0PrA/KOgDbRZMcf5pcamS9a+Y8TvV+lFN3NchZFC5R60etdY6Gh0Oem
A8KY9DWeCVfqh5hLI67hwDzvvX5LSwSVkdSw+WrP5dmfOtkmfS58wLW4lzrST5WU
aKSXE+1Lwys3zsHIUTyXJ70u+rQkOWjq5o0NCVf7yQzJXtEDtPmvRhgO2+1m3HVQ
CMaYDqAK0guNsVbS5u+domRJDbdiBRy8NuRoUtq8oBZb9ECVmwN4glQsw7pHmTNk
3tGRSLM3VfttRtga6Z9ugR/564un9++YY0V4sDPPWaxurtyWoCWB4KnkwJARvdsJ
v8vW8KqJWS85nMATZ2mUD8E7Lf1DQQpCD0/GBnNw4GprlwxZBcxObzzAuYV1/LNq
uWc3LtPXfaWIURerETDJ0JNKtoRCWDo1xs2fwnT2tEXYeWjiFpgD7NyEnFm80PQP
mkahUopuKYBbxj9n0NdewRgNFGBDhSMLUQ7I5gk+tAgOVhwnZhokJsr1RA4M36hG
ZoyLUnRjBkZfeZ3WWR8RPjNP4+woyjvK0CKQO5kCeIq8Wn4NrQjmNLS+cR2iL1PR
KSoT9cRd4n/Ym1tKgnzlg5nxudcal6Vd/g51ZUoFiWabPHhmowYAS9coZUAX13yq
ZdrI8rOIg4ihxWowtNfR+1X+aavlEJYcgWuvB38LxulDTI+f1U0Xg/rn2ohnDAkX
LMtv0iA57WnajXF1jrJETvs5EymFS/PygyWJZuoD/hWM3COO8Wn6A5N+wciPxpi4
TXXp6iNOHFhIBi8X4q326Iztkha+No8yCn9asn9EAhNGvjwSllmk+EhL0/4lHwyp
ONpYWTdCNDn6PKoUNoipyk3fhPeWhwrwCqHAa/nC6Rpu2HY35GdK/uurVnwjwMEc
o12oB4XPmNDLbgwlox9QinNzPS7ZkG0r0Fy34VS7/AC7K5xiwInwjoM2LurWg4xM
ai2QmSWl4RXOGeAEnpRxc77ALJK11upD4SYbcsTkJ4V6Kz7gW2NJ5WkvPLm5lhkR
Al7s+3oG9Nv8zYxIWKp9UeWxsKvwPU2GNDzF+il9fp233gK1jwPLx8e7V8MUfv7n
Ti7N6V1+kXgTvtDL9JAXH3B8A3epwW5VUl2/rD7Wjb5MhVnVhV9Cr6sQctmn6lZq
l9li/Tr6WFBQoR+YNXQik4kAb154L82JLQMfep+HTf/6nedh+4Z2STtXt6uJdGRz
UnYvwoRsFFLpF+4mi83AtmQh8/F7wvgVmb6mu0au19adVsehK4QZ4JaBsrXFbjUE
E0J8eSZIO+vHOn/eBbKQfQ+yKn7REyHyQy1pAcVFf9RevrgcFCXw/fbntSLGshMz
KLNxzEPYqbtPSVZRlxa86dHJRyxROXYFQqgLEv8+pg9AAqnjAZPtjvLUc8MOahll
kY7g0me05w+2J+dnu8WdStRVsh9Ko6MJXyuOwoXj0OTep4TKUFWQQh6KqwxTpoIK
fxmv5Z/UYT+VVmQ/MvCiKgoOGXg4QT9+LExL7pVbkKDEl9dqX8LvUPUvU1z2hFRQ
XxrNsBSAHlvFRm1hFLN9Ep+tKPjT7p2rFTb4SaG3jxQLIbJcMhgNHblIgi1c/jhv
zNgBpFLYd3nxzWEv/zRbtB0Ccd9SbPzOEnxG0cVjRMHEmEC0+ZZ4T1383kncnJ/1
iXp37J/voAdj/b9dNAJbb7TbLQaGdD48L2MDeuwTwKs8SBFUxAPaeCzcJGfsZvHq
Zfu0kB3qCUDMnxWrTC5IFE9ZVWGMB1U8AYEulnInz/hJ20A/9w7Sc2rda5PmaK5l
MIq19/aX+cb7mpntyXD6CE/xTKFO1GE2xNFLuGnfIlN5BmmiOWhT30ws0I8l0zcQ
W1bSG3UzXchHCGlJUchagG+VFiluehCqMhKwxLlTAS05ZrmMw+EJHDRvppW/GKC6
cYo2wu9h8L8VTENu6XJXD9+z1fkHWBiqKk88DN10P0qWIXVaHpkqUPw9xD5F4yuE
LLpF35+n5d8q/TVf6rIbRb/xb7cIi/YVLIfJf4IXApDjsA4vb1NtbmSU9mN+liiy
hzHu3/RLbydT2vxS5bdQcMT+1I7HzO1V1nRWBPR87xuyI04HPsZzzwMrg+rN8phP
rF2ooAiRImuP216lNTHQN10kbgfNXzxq0n7hbnvoIsB2fuzsFH5YeuCoXqsHPFgn
WUm1ps2vju+iD7TqMBOlCdQSUFv4hC7YVglC6WBpo1hnaR8hAaKdbLCDWWGN+w5+
+dLTP9XGnxS2Vmegt6XU/1P3kWhDT8TBDjNUYpY9gc9pjxrOsTLK02SbC1XiMTgq
N8f6OJ4Pav1wmN7vR8EDLv+ydxbljYQVl2T6O/U8G1kfzs3kxNc4u3XjB94d3NeA
6t/QxqdihHNXca0M1fR7fXFPzVUcmT6fUkHDnBOHzgsitlviSipawTlkEp5y0St/
qV6H8BugqOuFDZp3o6wdP4yuyOe2xd6bP+DH5NE/ql1mJSbjR1dkSXfeR5bMQF8e
NFvRL1CkbI2/BbgsV7fJqnX+XES4rrNprXzWRiONzl4IQrteGu7Y2kUHIChTiCbH
SvAJ+eDv8OyZhtTFzjMqEsAkdogVe3XfIJnpNQVgOvnHy1QOmSTQrlZjIa0k1C5x
CMLaqReuLtkOJOYq3A3yAjtM3defQj9RIsdd/IH4GCK/lv0cDqLQ+Pcgdinb5YSA
AzSFxMtEyab5sJOiv22nUYvxDF2y5Ol8eT9JEgV/tgiO9PDkoMxK0/GierJrPFcE
9Rzf93D/ZJg3wG84r7pggPmTn0UVixlsum1LhPaUe+fMHapvjUDRYpCxkW9BfvcE
dwLs2JS77yJGxepknwjbd/Odyqo6l59nKx4NSCqWC5pTo6gfqwIrnarzNtsi/uxD
Z51MIAtXbQPl7UtoIFM/Dtzx2sCqstvRypBLALPtQI3X1i7E3gK9xXIZo7hVnNdc
BVh3f0asI95bk8vx0hLEG4LKscKXYw+MYAFkOLJtVuiU66bwDdk0VV3eW9d/53b7
IZcGBk7rO+WiFiHnoLM5yaocNdHf3niaaLSRvLK1/1Nk5grl+yi3W7XKQCbrVneb
EKkwTd7Qc5+FZkR6kHfToNwL9Mylc7S9ObBgMV050CvIcdJ8eIS5HIMEoRdYNnyr
hBp2YH29FHtFWT4ug/N0CDAdlUrSTZ+Ftet41c5ZndXG2IKWoVIcX8Q5hv71/xZb
+aJ+0fOeAw+j1TqR4yBdGZ1WS6InLUPOJvX5XoFsia/j7Ba+MmlXQcgj0RCt9KR3
79OLnbcJN2WrQ13xnHk5+PSnp8nA8BOUF1pc7AXPtzh430Zyj4REufJV8yY+YaCg
E/YIrIWYNyUJ+78emOjO7m6oZEd5uW2zsQLm02KDYoLRtyKXBhbcHKcWSbeElRzT
LVtt7xUdpo4ly+j0GQSlLiqIJhL+Znpg7chie7IWnA/1xl9YeIzUQjq0bPnk3DJk
0k4kZtKxlk9e57crROwR7jybhVWyeOBvm5Xl3myKqDmk2w+PLjT7bv69HCr6i0KE
uFT/0V3jFy+M63TMu3Y58BuehYhi3AAEGltLyb52fr0CL1PCcu8Fkr6ytXedy8p4
gyoAFxCT9bj/O+VGfr9aKbi33/e/3xWukHn9YyW1ntCBL3G7M/WzKJhyLx+ApR5P
tG/jRzpYm5rqxWZlqkrhx5CRFxBer7aNpfvtmbOPrAq88RLtFiCTQYT8NbOqg41D
fUGJcAu2EfjBWHZLa2jBj37ve07PWa0y9MvPlmOBv/LAWep9dDQpoozdJcp7s4hZ
XLEcMAkC55F85uk1RAsF1+U9vqr3nMQyWyGlx0bdCg+Sq0142/1agl1d77lAPE4/
NVy5z9L5HzJwq6eEYLH7oOTVBHTefsvt/JWmFsA1/75VPvz7v/rWEe4FxnOXGFSY
ZRIB/hvxDAJSZkL5XFbCZNXQ/qh6KoSiB/xbIluScd8K9x76vQmIVOSEF82X2mh1
y/n5zSOUYpaSzTKSkKuDCGLXGkPK0hUor+MB19CKXJNZuO71iyB7/Ia5zsUhw+9w
vhPLExAy3XiYVnYmLQ2K4KV7h95gQ5Z86T7mBBRP2zzLRS+jswb+/zwd52uuR2/2
sD0uojnxe3WmEYpGy4/DBHQt6tkvSekbhvTTNSqEjYXJN+avs212eGVdtlPr2PlJ
PkLlHo9er5/GwN9WMdZZkaSpnA3577ThwuT3sGmnyUxIqPKbIpbBGGK5bhq+pO+q
whgjc7x7F0Zm4BtQh0IbFUxCZJuetMrUWi/RN9MKUSOHmtVhZJtjXJjOdN+0FsvV
AzRjKrUB96VZMZPz0z6Mzu7DAyCZ63og/AB/H57xYr2UxTKS/NP8lsDXlmzftsMM
lLhFqGfrUpk/xyqtPc/qQe/RqeaQq2bGzovEO06Et7alTjgVme+0CMmQpypJDwmW
7WYUXubOXqfRdRJyFEZK4ilxx7efkf67+sno7JwbKEKuixOeJZcYp/wOUXp9we6w
z3xt35RePsSTDJzeLsSPm32t7WJLI1I9k3R4AyoJY+L8GjAFdxprg7jkYbk83Je9
vBxkRsjJbrqxQNqDq70XyUzo7rUReblmnoq2fRItBoIVkYhfOEKyEprw0F4e8yDZ
88ImQhBOXbeIq6i2kPjflT9giDRs97965/ANNaMIAzAD3ljKJdPdgO4yBi7o+oER
93VlFLxN1LS5bs8Ee92x6gsJ5+ktVHcGgUq4Efi5NCKHZxcL6Yz66Z8MeLGPZv5/
QQzgaBbONLnVtOxenf9nGkO9wJnYIvpzYWmt+NvS0JRPrGQmu+T5XbxDgxhiG1S5
vRKiO/5JwkdAFpT199Ei16/IxOyD9B23jMKiAuF2M7OzGUfmX4BJtdTNHELoud2E
3x/d++UFhBoUGIxRJ++Dxz75++UwEyY8Qjr7InRIGZN182kKhgLlqEimZnYLdAmq
YJL9BCYuqnecXkOPP/aNQrsjDGGtiAJjg77CJQKFHcMTvaV+koKFm1Atn58kiZTq
SBJh6M1KXGAuJHzFS29Ece16Qv7m/8Z9Oqgdx8TIEEzlG095D4VVi5KlDqKtxuF3
A+VuZTd7hwsc64BYHUkFW+IC4/OwhNiXmnsSrRahwUtXcK1DEy0IzuDAuaUgu5pX
52bRs+1PsRS4N4ymEV+vhIBiemSrOrAcTvu1Qu5h8PSSvcLLoY2IEZVfqsV7fRSf
/l4gh2C4BQECfIg/T8advQDIQzmvNqjAtFD4PpP73AlOMcJuPlRwFKEY/Sp5KJcq
fvyb/gauBAJFn35ZztT1V3E/ZNmwlgwrihZEetIbPuZjr5m+J8ykOHFVN2CUj7Fd
o7nHiNFQZVKs6TXzZ7moOeTldJHM/J2L8feMPG66S2MQX3cXXkyRLMolx21pfZJn
KX6P2aTVuBHvysskxkQuQrZGG11xJaSmjMtJH6KyE+z4w0QeQSIcnPTdQGOWNW5w
7wY5lQpXiUJ5yAIFhpdwhGhPXXnHYa5digRt1BoUfsPOG9NNmZ7nRaewlhmJMU/g
TCht59nytsMxW9qsJZEV3op1oAXSoc/douuPieKWghfN/AtVhc/7i6TQcZsZ5qhn
JzAmJoeD8KRGAxAQagtVmvKoHGWwgjsrsxwmTDHVn9vrP3bOJGyC7C/ojDzgxKzJ
PFNKFxasZUw0hzwyABlCBPJbox9Iqcs82NDoxurPEdCCR3pqkHSYQl4/53wShTu0
m2NpzZtJxKXq1eNobCoaxkDo72aAGkW6iiAV2Ul9uT3qRmUthKml3ClN9ANhcy2r
NXq7tc3TdMACPQKpyKYV11JseJ4PVExcIEcaUpNr/yX1Q0FeG2QQY6xQG6JNKSk1
wNvCNPO/NkfU16Rlb6ZhJZJq+Wt/1dcptpbhIb/nrFGJf6Q9C8RvbuE96Am1yJhM
wKZH6gFytO071u716Jk8uQA6DXchJlVymeBg8BXclYC5CB1QvOErw+rs06xxFfuW
l4lnOUAp1vD+bTZc4evuvmhLBx904ZoMXdkGoCVZaKR5Z4sSnrmcESK1UbPWwR5H
jZ+zZOE5mzVqoW3poyFl6ZYxkdqzDNBfVeUvjuKUj6cpNL7zCSaN95X3lzDJ4TXZ
mvjrP+tuqmaQn6rLJSFPq+lSpG1ls2fKybMns0qpscSHhLfbDm2cxUKRD/cRmiK+
Rmg4jWZcfaePPGbQigymmD/0s+zOUPi19XtuEZrx7jll5C4I0Dq+vS4tJWfMBMqC
MYzD00HlbwT+yNJeeFzInw0I/2DLmwoS5CGPARL8uiWKEeuy2JYkcYLIo7j9PnJt
yIvmoUewXHePocjlzPsGgirQzCHzHNntguGXPkFaauBKY3rPZPBUOJzGh0/1wSJK
d+2WPmdwx+Rn8GEVzUnktf89jW2krCS+oEh5VFhagD2IizQAWpUZGWvELARcoknB
Wc0J7U+ZEpZAn8swNLC8jv0sldtqNSU1O0bb5BBu9tWbxdQe9E5UUxGwVfmfC4sw
RTFxnCnbwy+yBAgYGFX9y5HB1c5WfkPdvUiGdRudrVk1mZqMmWhpAwIRFCyBZMs8
EFkwoTXZZnooHjfTYMG1bTiHbLUYyISUsyNuqIcQmhGaThO3g8564fStxQ9u0SkB
YbhMMM5jWUYcvxZpIA2pEAxOqlcGQElCmevq6zKZY+LDt0CvAKoAULLBdRUsD5ES
A3b1Wqw/3Q3hTMWT0GyW2S+eGxYDDPSGmCK0/wwcav8g8vinw73fLC9v1vCVgdy8
Va7msPG85cwPfDQ+1maDXR8l0rHEWuc15qCeJrHM4FvDNwpmMr/bS5DXPDg8tWhv
2cHpvkv3S7EcYDobLbp5uhXWK/GRbdvtnQbpFrG22ua+vi8IR/L+hRzVIIUCXS3r
8mr2i/zhdWG1cSEisDWP+FuQXVMCqyow21EeVU2jGctmmMdhi7vs5q+56DnMFc4H
VflRK7ycZvXio3YIZJMZ8oyqfevl1U/AcOczl63yl8NWesjtkcKQ0yfEeB/fYtbd
ymJjtwNwyKnDF3HEJ4WYyWigcQz1w/f2fUIN2OAHYXysIo/GdhcTPKm3jIPK9KYR
+QzAoL8rgsSKsZjfEkFx/CeuFl49ucwPPcQcQRA8Fn2vBFGFd1S4FmL7sOQKr5dv
GG7DTq0+kbIUNHRTLizEg4TS3uaaIL6LcnDERRF5FZXoVrdqFPAZ6vir5OIXKPMI
LM+sH7xt5BPddqKCoPRd//ktVY+Pkf7o4WYwQiHaM+vZcAjOT0RoQSKnaM4toYGG
054GhSFcEpGv4zqpVjSCLeoXcExa65wEP26j3n4vJy/jGXmIa+DrdbFE/IgfhKkJ
J0ri37D5HffQsDCy1y/I4Jd4jnylcsn/LkhdDyeu+byfQX771u7vc2iDx0xu18RD
QYT+nbR+DRDoBOtM1m1JQxKM+4OH0W3UfyOKI1FmtSYvlix8lBS9j8TAwn5ra56f
F5zYFTWCRjAXGSHAevuGkTfeDPwiEkREwRc8gWjitVjMd/Cd78EGQvsfyeiIh3+Y
SVnU4tSQUiL5av5cV9EzQm5m7f9jMP4O3ohYYNoAX4RpTFyKLceEo1d9ekTJb31/
wOaSFl3F7+qIEZ+2AhxKRmmXiuBaXnZoVlNAhyzi71M7OCb6aSIPSOGfq2mysyew
/H7Grm0JzwiUczgOdM3RkSdfRcgLkWHWKtDOu0Nwlg9aZrqf45r5AMnnFTvXSmsV
TcX4GGNqD9/2BnPmJVR/rUPKT+4jjzzvswxxw90Ao//PxVc4x4vTC4Fvu/kN071s
Neh58q5KL2dUUCueg+6h/9I2Mspbh00JmT9cPzc9noEYWPdJTlMl7VH7LqSX48+W
puADqlJzM3+ymkILngMRBuQcLmjcPPB6q5u24PxY6Z3GvkdhfxhtNGZZTBKq4Y8M
3xuzj+tlEElQhOLqVwSw9OSjiv+1rsMeYurdMZp3ZSa8jLuLzwpPIRejVQSaK6T0
LswhPGofNY2xGPNsEPLQznACODmzRAJMKAGfbdhkwWm6mVY3zX6X7GKxzJbSH0HJ
y9biImpygsb7K37eSHgX6tj9JOgtJhpZ2jiWaCv0gIEXSvE+OL4ZM5OpW2Jlzlq3
MLtsKTDDNHF4sxfn9cvUTOdIa9f1z7a7pR11V9BRXNUpiAVOS657jrA3RaeiToi3
vxpWLBsAghAxgBQNKebWJrA0biuTKEhMkhLYxFvsJTYVC8nRCzhxPR6Vsjm8ODeu
RHTotV2JruAUoL/d5k+vLP6JuBd8wLd9vPAVhC61SQY4utOA4POpi+mWqNewpUJR
t24IPafen3actsYUbVnnboRJdBuDCCYBpBiJONfbkXlCM+Poz3mIUUnp+JlRxPUx
6GICdtwo4p34uig3HTrXiy0E+ALP52fsprkZkh7tPR+Ici5OZp9GcCqHZlx6KLhu
hPUOAiGpDrsQFRQTi3wsHLL08yyfdPeeIyOBVjpP9kwJ6+eRqx4cXGG/QDYpDtME
PUrnrTd4bThtD3cA4ikfJa/alqe7n1SpxtyMYoUD5fJVgzwj/Dh0wXe22lsyGNhR
aC7QtwRuwiMztR8YOCx/cMKugMWr1p91FhN8YL8lSRurjfV24rHrcY6PYK/E3qP/
tsPcimI98cU7Rbs4KQyJZ71JtxZvyDjYFS2yWf9H7oh0S8c6AWpFWc48rVZ/fQwJ
FtjeFaZVdJmXRcBFQovk/iuKJQdHW6BEo3pQ6S4P1yHG0q4OSxVaZCP8HMF0sQX/
fnsypP9Yzb2cfa8bU6ucj1lk82M37Zd2+CJGoU/cvekPDniDw3+jPDZ6QHzwHEe1
y4zyrOvyZQwPZJm/wkSXaBjeU9rlhar4aMUQDi2ul6GSDgoNhVFYHukdFuVxnDKA
Ppexqh5whLyQHfd1hWY7Geenbs1a5xrMRjSef+jLEvvDcHO6VWBC2BoVWawa1ehz
QL1BLq8EnG1w9O9qGsIwcGPgQV0sOnqRyghlbxJbgNcwu8I3S0roq6XvAxuqSf0V
7nnu/wnkDVF5FlreIc6T9FKkiRAUB+Zoyj2QAGtvjV6Ne7Pj+Cr+9l4Fy/tVQ1Gx
aEvNHJRxMsUX9oCo3+toyHeA8F5d3oVpoAaAidBpfGn+olHQqdbv59cQnggg0dVF
ObTm3BonRWRS1d7fOzqOaVseae7WQ1QJc/0x07XbAYED71mDRAxcgYR1/WD4+v5o
QZPqI2d0UzsBrZxhAXCM9q9oy8aXN/lC9dTmaBaxj3eaB8sHnTnqLWR304PKEN51
5iYbLBPSVO5xH2tVo3VLZ4bIG1Og68F8xHHSGXWWhYzUGQXdXHyV7csJ3u7lBdwF
2ypCngj38x+GQK3DZL31nh5VYnNjSwUdkpEzAHmbnVDOnJHYqcsRxO6iGJz3jcgS
vX8p5l/OuADofU7djO8ixTaWaTkTWIRimwOdr6q6TneA75KRA3gcT0Wtcr1HddI2
UrqFQqWTP6eVzv5EEPgwoyT4oN3zex94oedl0sOBITKFzhHwJo/4143xeQuN8R3W
IifjeINk4fpnIvc1btRMA2sDRFhpAaVcrCtmvL4EGlRgwXdybInTqyA2IFNDT3DB
bOfEBtAQwgmif+riUqrF0FeBsd3en0bl0puZdBgJIJ/eUr627lvt48jKRMIZmj6h
jVbXW0d8Oqt8Yi82CSfhLzzgAJ40eVdEI0v9E8mjAgNIQKbpJvlQ3cu+o8SMJ9/P
DDzEUiRsb10/TQE0exBWs+qshCzOYkTZHrR2WFygBTnxmmqLu/TwuxInv96LfHcV
moe4qSw5veBomPgLKeQaQ2P3XVrxI7P+bfbtU17TpSvIl7/q0wVRZgU2UNyAkpdY
TGB2swWFL+velGf+nadY+O1EIOum3BBSlyXz7AaVBvjctjQSoLenUPTAo5EznDw1
5C0iNCp4Ax+871dW4txcMkOp8W135IF5+XoCBl9pFrxF6U00PmZAurh2ZBV+cWg9
ZAR3NXFBtGCt1VbvrU2jEGo8SjJby8JTEUtTlVCz57neSzGRRj5xT1lDNaet8PJg
6Ng+s2e9U2oVUIolxgQIP4z+Wd4kfBhEZW18BE0OgcvM3l9NL5DV0DHaByi6Bslq
vHD1h9qIjX0zQ/h8+7UGADe6s43/EkVFoKfVU7ic4BodH6ZvY/m9l9N3ObymN6Sk
KqJxziCLRAK375dhVrfuIh9G2hbe7UOi5F+booniXGCjrH6Mdz9Vt9kTWTRwSaPO
UOn8Ua3UL8Tl/7jecgt83AjWmhdFQyHxc4JGn4isPA8SZvBLP1wmPUGtE3o/839C
4jRTUlhgzsdVVGD7gN+nO9t2cFoYkxmhIvabAVgSA3keSzY9py5VQcokheQst8xJ
/U+1huYdka0gaTfIbC8ecPz4lBdoFWO36BJ1dmfZPqe+wHbnPePFsqgA8gQwvcr/
2NRDpW2i5cXC+AYMokMJ/fo8LwF7GdjV8mnnA7IYlNe4dNZjzl19K7tANlEHKKjq
8T2ObjPeB4PFZAIBe8gUEXGaxEza8+ZXAzt3/WQS5enMSOEWTt2p3bOcl+d2igC/
Rt0xyqYPUVSFnfivKrRNIIrICMUSmhdYQF005lJA14840pm0x2W2ym1H3wwoodJ1
peOtbNr88cG+ahwM3b1wB5LJcBUSjk916DrYzwwqyu0u9ewyR74I1kf4XOON8EEh
0v2ub0q6UcRZYAJwIDHBLci3D1GBmRbQCiV6tyOOv+pElOVYiyX15JJgoqOANPtx
JFO2MDdp8FLkAmCUk6pHcnrsluTxh4CdLShVUuU+T9IoNYVvuzdSLmSwSwmDAjY3
myMp0XMyYdIbgJMfzvmUGyCxSAZhnEqi9mF2rJOesw/SHpuYvxoZ9rYYiwj36Wbd
URQ05QEfpDELFmmXyCvp0hUBJ+Uf/aZY1iePsh5bPfgs0d3BWwinmQwSmxkDA6T5
kti7Vksn/iTjfScK2A8BVFD34UQeLz5Dor6ILtEG1vI4UJVtVN90IUt8xLsVqnqy
v8oExxhAWm9zTYXyYGTXfAS9llvN7gTY1yjAqbX9S8hSG6LeHof1mZ6FAuwZDX/D
hTYzcNcJjBKnU7Dkym8Ky25VD/jFPxelqtKe1/bCWUPHN9IbjZWIiShk3mq1lppv
K8ny0Qp4ZaUkieadEuFfFCb5afXq1tvli91w/LCi0FWvbA1Qn5hDDuf2N2I+IL6K
j7iOks663v/WC9sCZVphtfWZt7fGIn62gy1tcoy07yDKoLA7huT8vHkjO4iBYGzB
K9pldrMdS9fbUB05bywZfuZGYA6Il0QWU3bOW8hY4b7SA6BfdCJvLjDOpdZprtaE
LUQls0LXuI7o9s9yY5LwPPSY+spbWor1NXqfsgd/m2vrMzuNLOZ4inyf481Kd/KN
94rX3JyeT9VlTOd4rZ2pkwdXiHbO3g9tfmAyAfZjK/2Kf4tGrZwvA6vIRgI4+zVr
2bLejvrnL9AsdFvadcOIl1nPcMf3qM0TroQcP0Ru+YzpyKBIbW/3GGlJ8WHnx8cK
4B164uPlYdu0oMyhdKjkw9ju+41eLjbZPrX2TAn9g3JiP/N+1el0lkWoWgmeBH87
w52VS50fG2h3yRMC1dLxlFv50VhtIDdMq+rln7YbpujVD4VUaXor+VP/yhe0FOb9
wnG0R/XzbhqrmbX5ZYNdI1vUchidWJrvQXGNHWcKj8BfbUMht8ujFci0OkL1SJZl
mE30iZD9MwMF+zGVpExDgQ0k/v7r4PISHDX9nmPTgsOGJJAstOueoW3jqaVvXgTO
7e/z4w0umG2e2Eitp8KxUlqb6g7lRwqY0m7OfrxtXEIldEAyEewlR5tHAH4fTvw8
4CFmySkUoHgF4IVasFl5fmtaBp+3LIy4gkuGkQ1A+ysH8jKE9F2aVHzrHddVclmD
pds4YseBlXp6T7QxEpXv9RteuIOvpNxhEA1V9F+qFF/1h5bK+PnIJqKq3FcrauAA
URnwcOENlT7qkmuYHASQ6DCwZCxjZDm6t5iX+HtDETS2OSOuqPYPTG1Ges6KQFnZ
4FpRk/5343bevmMuvgZqmSQE8x8oVeAjelIJw4ZhExWCUPTTwdDFrE1/YAjK6OLv
c4w8/TkkbTlu9YvoTcFhX2sBbB2qp796KB4ASpEj9ou2ZCbO83iiLgg0vU7Y5G2Q
eNlONYzHHQy3gaS4d3X12yTcUQixjKs0EKJBQ9O2GoULCGWK3raIxVxAKMuvwpRN
Q7JI2Va9pTOMPIb8WDrYo9p8Emx1+yDe6Rul7gxPRqVpyMwK4hJrhi1PL913EvKv
th2ZkkZbA/uUrrLgSTSB/vVub1DTYHWW0bzbiMejrCMwzDl5LwbguyxKgFT9vNht
q/s+PivyPQtSmBOb+l44C5YgtvXGwDWMbZ1BKqftwQJlAIdDUA0abA+WTThPoxLj
2nsmrlO+pHBwxdd0rzXRcHpuupO553WC4lswEtyjjcqX0kXgsyRNEz5t6xpYTrv7
aYNYxOilTDrz/lNzGIsJMl2iQY+Db01/rLS19pLMFqmxXuCGNxdSK3KnK/nEiK0i
uoxs0MsSxoQjqQ88RZEgfdSWzJxhmeVgeFtHNKNa5560p4k362Ul+yogiRkJC2bI
EXRdJh+NwYeVRysdYbSqSLRKLsUC6t9deqeUqKCBtot4ik+7EVh+29eeyObxAZyY
zlbOhW2DvKDGEZYiKY5JNbVddRn0dKqsZ62H3Te/IhpP1fhLLP6BwQfSNaLngIYB
a7CoXarP0vQ1RsYp3gfNdyVRzDiDKsfURyKwE+Iu36dhwdrZQpYDWjLdQGThkjUc
tkiSxpMb18yrNnq0DsOJuya80fs/NsgdVbqOCRc3imymoDV02Rs7l+G4HaoTkywJ
AFPM8MXAsWORSLG3WEU5I91NOHR1fnDxBF/RG525MyqPQxXW5KD3KEzPwVhs2rAm
wbDRjC0nbpB/rajJeEQ2txUgKSgwxlDkq2YMZxDnKtX5ZHQ7ThW8Yku8NfWhJMFE
KUnKDmiCU1gAtvMGf/eyptS3ENTWauF5Lg+DZraW6vgb3NlZ4POwH01s1BEWXvpb
0t+sy0z1XCMZx327NdppB/IzniLNzLOl+bY9cCqmwbSIDXn7QJ/nI97LcPw6DS7O
kZNkefVHCSEQsc6FhozOROJDGVWwPFah0+7+95KIavGENhci2PfdiOyDm7/ZQYt/
MQbTOGGGvtTSObbYWpE2njbIXhPd5cyEOZafDYtveWfy8k67SK8WHWhjcChAAVN2
ieqUDpa7zfr8Xmb9bBYPnXwNzY2uLXhPZ7TAONs+FCvdX76u8+1uI0VajPHwafPl
fNGPMHM2Bk4V6DnCE4STvlNsGlxz3C3knh37zOn0ZVe4BgtulsRT5Pr4RWisvxX2
bu1meQXrgxe4ID2AeHd9kyk2Nt+3TrvzdO2xXbS11dk6jcj9vIIhZCT5QGzpE0kd
AlBQyc0GAAcQc7NN3FNk2xgm8bSsLG1DqJBdYdRRwdL9Ppm4IsRSKmo046BnH7gF
M9uejX01qBZsUKtLhGabY8b+HyFbJ4dET031H//jeedoDSrD05eWOoF4FTxNTGCE
39wvNvCEmfuLKFqevWi2lALxSe5G2sMJMQpEYH1tVsqneD32G/l8KxiHzMtXFBJa
nZtBpfZ2LBYBATAQjVmqKdOXA71k7MTecwqk7xW8H2epHzyKyshu1j0Ph2k8y+kf
u9fqNVafs7NskhgzIqkiLQ46b/tkAm3MBr5PtEUjJxO+ywM6p+r4pWZXc48e/qTw
Vvjqa8xlJO4exuTlaKI11Zw3uPuQu9zsZlrRtvWmrqtctbKsfKG7QCa9Nb6ZsxlE
3LXb9i88iyO46qmq6zToymKpG7OJgmS2/7Mc7cWGYEGvSD8QFEuj8OnLfdWmhzNx
vadnWPMs8em2Ej8DOVscHF5E3Xd3vJwXP2FIJ5T6AKxsuoWr/7aYM8tIUemY3Hg6
XHhG96ac6OvMNZDIBqy3bhY03YUlBSec4qjzRUZmhhOt3CaSa1OeTTiosrb76cl+
ikGd3ayDnuo5FARKGqA1x+VwfFZ5PjCnYrbnQi9J8Zd0k5Ftgpha8eP8SCFJY4Z2
xtjZ7sBoHJOejqsISCmfG18+yOlIcRwUQl1LwnYIEtJNfxWNzFGkJxnpMzNwarI0
R1L/baBm75AY12drMA5RgFO1Q1tq0FQH194GYNy1AlahPdktrq4CoSOu3xupK52+
AAqxys1TALNDG741hMlMrAbXSxmdmmPGv/qtKE8lsEWmNrcZtHjJYeGNI795t7p0
RUxHcPvicX8AaMQiaPygIvDUksSWS423enxGd4TE/PwzZdMa4CXTm/fhI3WtlaoV
GMbp4Uep8RNkwv0bZ6/i97AIdua+gQ9FyGDpT6KabQXibJ2DzPSKfxbUPLeoaCzs
yQNBi4Mnp9tJFF9SGjPz2oSz9JgoMGSWgS30yKcSCnK9bXQca1dn9RZOatepVsge
TwdQ4SFRMsieQ+QKesFrxKSxpAWdS/6N+tHVEDd8a46y51tPv9tmVHTwgtz9A9to
i09a81MNbP48aPOX47xOTtgnLHJ2oNn7kq5wqv8ySjlLucmV2IqsFFDMdnUjQT0q
DTw2CXdNt7QOemYUtWTlp+MH28UwMCtWXvj1Nj3WuUAdMzl6f9c/Q4WGOjxO/Ehw
QmDh1uxo2hdJw6ZpMDUFjwkFwiOZveIutyJAJfjk80fTG5Hiab7NTXUD0PpAAe+5
u+e7VEBp/tinjkfOBfjp5ZkV6L32ZHZNNFKJAaZWuPidU0mboiXUeHgEalEKh+ET
8tVH0XXVlR8Xes+E8nCFAelqW/06d1FFO1dPwsbaicCNfImX911IPClgWrpGHYwL
Dcks2bmgyzMJtcu9dYDVbVuindNdcRcMEcfpLJ6QU7QYkFmY+Eies2fkxntCdB/P
eIG02pc1HCap1uBOL4lTc7t/qmypmY0zdeetQfNVd7Mv4q2sTC99CUyNc2cNn7sO
OW8IRG6h8FO2Z6HEKPkhYnR5r6j3T+rWrgf9WiVdH1RP8PxH+ytqKaa9rQ8T/Tiw
OtWtOMrVm6poDv668K8FAJFQ9e/RUs2zchEyA0RW1WzeAXVbT0t6VkUDgtD7F76C
j0LsQitLwY8xoPRaOPuBixy3M8cUJ9rkhMIzpHTlkTMor1zTqcklot2f9BBCxlNH
ppklDQrRMrzJVTkj0MAFprg6xh9loXWkSUyKuUEQqCCX6dI2i00VZvx0mBhG5oTZ
1Bu1D5fenDgQYFox7XkZLetGEsEO5TBKf87wfOYvTTYmXLq/Fbt+5C0Q3kFoo8gJ
jeEut2kZJhGXrgD7WAPQrIkvHSi2gWwBN7KwV/SaViNT+s19gysAS7WkLpXFqdoi
7Sy/BUJB7Uma/q/ABmdIa4z2OSeXvvL7Qk3t8eQj/bSy2dTCOinANZnWDzMDZJgF
HKPr62LZsORy0UrTWDkErhIiVFJkB9+G4tGcTYURh5lvRoWq8s/yhwocS8oZ81MO
NsJJLGto7/rOa45TJ1UEIKcXM6ttiyRocwtj7aNaYmTIZ5P2GntSrR7tT9nY8jZV
q2qx5gx9b2SJM8AVEMd3cpn6EZgBwoF7qMd0M5Fik0GHnUJolOMl76k879eHYHm/
VlnEjMPv8hQW+XxlhjykbjQVyYFKlsDJcxFLdzYekdu0bMnHqy8sjvCPDtFGoWHx
UJuCfZJFVoYYm0wilg7jJjY5Ny7AOMSerJevwBGyD5P0yQZmTrogCT7l1xcpsPCW
p4MELx8Or9xT+1pBg3bCDIywOYYMloUTG+QkXc0EP60pEHYy2mnAPS9CbjrVW5YF
fBl0OAi37f08OZ/kZ+Pmx5LgD1GJyRDQA13uuhfl9DQt44gcALlSQP5W12PXUMgT
e1jkSR0h6O+DcVchxwCB9q4i7GdfHwdf3MknAAI1J78Tq97zu+efyECr138SCf5j
ok39UuAxRay8DpFPvd4Qc4amO2adj36wUZzc7jAzxG6scOQdQMUHkmA3YvaiQ6IH
ytuzKvwdzyWncWERfCF2/V/ci5bXRUR4bE20y/6Zjzz5w+TCkIBhgmTmgEk1u8W6
9abMOW1uvvRq98tz+d+JQaMDjespAgDNcLIzgYBjk9d+8pvW28uxLNkibFr2uC0f
Wa9R+0aJfDzf+IAaSzaSFduQanbX0B+sg7voOR7/mi586LPQdrJT3DwdqYtzNikJ
HTpgqd17WSCiMhuwFRkpeM5fLUa9JJQPxJclTKVUFVnzKSPpr+M3B75BGGwcSqw5
WvCvlQEaJCOUudKDWJzEzlYFw/AkJMphbOP7cU+NM/IWXlZ/LYzsyTU3eqyog+Qu
++q1GFQJj5EV9ej6CLAWhRkz5IBiOT+TXu2mJaPpeyRpNe5rTS9jMyXlWpqdKo6l
3D3ZI/qDg3Kb8vNTlKY6UMn4bfm5doPLePJLIJ47UW4gMIPWELjC2TNvwfZECE16
8OuICy4FGYWFfmMyGBGsfKTNjqLJlJY2pFWqeEU7AOJ9VSOGWwhg9Xx4cPH/g+9M
KK44Ko02OiIsdYU+SbBJPi3PLufo7HypJIcrnj1+a/kiTvQBrkTwfBVDIoftgovh
dM6IXEo0Idot3o8WKeZq9FFFtChlreiFzczpYP/EsL7Oivj6JH1ORSxeekCMJsHw
5eKjfJMAOHf80XB93lEcq5vFy46RoqqZCaZyp5l+kRY5zH/G3VRAJ6qRCUk3/d7v
oXV4qaZUk+FtYNQyaQcNePHUYpDW+48hJRXw3lHN4+L4WYst8hSsnO/mHcLbBhHy
NNU9+xosHrHuPEq71UlMqZLEKi/kvWlnYbqeHYcVKEFrNLXeGToz5CB8nH/x51xo
/NbdxfBTeh+pqkUfSwbiCIAV0NsT2PoTDnIIS5k8vRRHOYEEp9zVE27it/S4SezQ
VeDPKSXV1E0UuTbTwJtVFnIPHAqSl87T8mTc9Yrz1ErjaOkpRl+P3GNC5T5DwZGg
dwEF/kLPG0KBlcG0C88h6gp/7T+e/AcNTL5j35TXln2dtuOWh+HjOgNlnUZHcq6B
noojBtpZVPohNz94ijVykejSQbC0yBB4ZoRm6vBiLHIVfWwvornAhXIBTvxnFjTR
0RBn7+nR1VYyqZ5jLfj90f64crJvlRBF996pb6m1TrSDBu1NoxkTFQm8ISEtF6vL
9ZGUgamgtePZTpFs7aR29awnmjcGWdG+Frlxy5MHCvRmL88kMZbkJLBwa82b4pTl
vVmA4tp9uDseATS8or5HxFNpf1KlXXI2A0xwOPy8aPMAIQkMMWcmu5LGrbYia2/Q
mwh6ugO4JzySFvNom6gEQ+ln18YGrUvgbYAgSA4ZBkJ3lk9cldV5thAlSrDD2vFk
japwB/sM5UddQ0NPNrv//jYR8zvpFzAFF1kmMY9uVKBg7Rd+uPm+ab4jdEZllSMU
sfjaYz4cTSChzQ+GWjeE1nAMiPg1CcDButcKHOdPO0r16w31XmaQCiDg3CbjhcNb
wFkJ1OWniN1qvNgzjXoSnb6i6TeUXUgRo1ZBUWW0HvX5DrH7q4Mhn1F7jQ7WdPOi
AJuBY0DlKscp+4igPEGn4fEd5bJYUm6g94i4GUK+TWEES9l4/NmsO02o8DTXY+mj
0Iejg5RuWbhh/rPnXVAdWJ1w/J69QzHhBDbaaeQWKCL3a9uNc/OSQs5Ww3KR/p9X
AWbizLFDhB9inMlJ6r8ut39/acxODK2sOUhKl/8vdhSAMonAggQgZXb8LDYNMZuI
EdjIQwDYUPeppvrwkRh2cn9wE1H/GwTofUJco3ekslGOP0vCBFi1BmN32SaA8WH9
kZotPtH/3ffaEH5eQTy2OOIj+LuQ6ivxj5MmJaS3Bgpyi2888FZj3s5aZieavx+A
s+ZF3bqO9Xf5+nlQgKWLP/8+UNgp03cxkILw2N9yNXus+9z0QXyCO7KMeZnHzxgu
xZiwjCFbEzoEhQtYPfqDUAezHzjwEtmUIybqC7se1NJB2sZCMeYATU5JDLppq9nE
ft5gwMLSwtpc1VOWW3QPgLShLkpr1tWXTwFwwoC7Rd+Np9Rjh1+A2BFBWPn6bVxa
M68NYg+Ub3sTeiwXt2SAHkB9nx3muLkcn06fo7sJrIt4lvk3fawcCnJ+1GGVKr9m
SQUeGJ/Lbe3p5Prpm+7TPLJXRVheyMfIhzEEk5Ym1gjgTg3Ntqf1UO3sTmDQswHn
ovQcziSMae1QlIC6CLNhKi6XUlDmnyprinbBxNexei4+y1RmI90l9vH4rPIARUcz
QoaJD09FVMK+3TgN0iRdhcckZMpkjoo+tk9lsAdbsS0EEhJzXKZwkLJqo0HNMsys
/wAl2O8wBRqemy5tiIc1fe++UBiT+8id+RnYsiScmwVjBHrRNJ2u56TKlELzmIoA
F2nzniiFP4yprezvHUQP5GzisgAj7dLSkQATeiwNvp9wKB1w4+kQGR6a24prfNzt
1qjAs8he0G8mACMFoEzRXhcMHctkWZdCebXRMCFbtlx37dBBnqUMm32wdCEVvvkj
9j+9aTPMVr+1GITFNlKXbZ1I7ZthzPcKDCTzxYTpB0bjE57e6fiNZcC7tzvaCqA3
ify1I4WN9IKrHZRXxDSkEXdM4UaNfJUSX6GAnnlv0TMWyyOuVFieY2nBhkqY8OAQ
OW8RjmTjt6rd0ssSEdsctOwnalnf4OIzI2iu1F8ctCDgTTor+pBs7MUr/v62TI/q
NPBy018yALVQSu+tfank+VGZCoqeFVSe9anUQwF59ltS4+lTnTuoJWU08V/SvmmI
o5LPZb72mm5l771yUvb0cDvZRKg2oHwKg3OHy5uRYKnumeO0PA7Y9V4XtjAZbgwS
ISQTXv5B1kKMJaEfZPBckOMVnm3VI8K0Q4fLrJ7MQVhlKOmf/v1J9jI+jPqNDEA+
lWW7wQ6OU1Fe1N6hc699FjnAg41dUz8lU47dhZdyGhkaDdFsIW5+hLP6D5jKK3zr
TeFUaeUM35wGTzB8EvoT9JigTnaahvksIPgOJxcehNN5CrXc3ROJMqt1sesiZI60
c5n8nwX9wo5tRUQBd/OpbGg+kYZsUfbKnhK2nVhp52sEn1RIB7bWpOkVQIkRJMii
kAZiMTr11Kwa6RRTnzkTbILRqjuxdWlUxYA4df94hUIL2IfnlWsn5WiPmxGcZ/VA
ocV8SsuIlFvcKb0K4K0GQNskqlB7cR5QCWe7oojfyjtlOtv2LOUWZwdrPISEcGFb
73CJ45mkiT6fmCEh2iscTGAYUU62AQiJN8tdFWznIw+b/1CfxmGLKgr7A32zSSPz
iHLtxxu3X2/PP1s0VxDrV+YS6AXVKXkoSRVd2hEygb4WioNYSQx/e8GhzULEH5L3
cIaEcKoZUwmR4EDpjb/2+YoCbFqZY9rvCjZc3wU+bW+nq4C0eT+i1mNT1bxpYDmI
p3N4puTpF15iQjsot9gblvNibzZT2n3QLjlEPGk76BTa3rOu9df+bzzUvHvDiYpN
OLLeqbSsxQWsorUPWZOAYnS9LkWv9q40ExHYw3DcI6OYGgZNVcwijHgAz3jugzRT
udyXyFIXpBXGjKQZhqz6noI+fRzw1DuumtO/dfuJDRCXVskaR0xBo7IaaLzeL94i
icg+u+LrbJeu5lVOqwQwFXnYeN7KZ90JFdEGpx4oGTD4NTou2Oum+xBzeqedeko8
TBRufStIvb7RlGQf/P1S3t/olZISQ5fxv5w/YQSPeCajmwqiHxGT3U4aMzk82fCU
XTYk3vb1Uyc/Z3sA8ncPBJq75ksc521SH47fnJ10DnKL7k0doW6y6MjJvEkJJVyM
EhsMuCx4vQIFSvsWDAo3Gq5nOXmeUrTPl8G+ZT/xpFeWfVzqYj0hK9XCQXbbYe/n
ntDFXUnRK+Z+8eLVwn/by0EmI1pFb9OvrHzPdwF+n6vdA2F1p/fcbO/+Z00LK43c
+qkdcb1SFC33WZmxyPt3SZiAcvjJt+sZCV+3U66jDW8JjxBbK8iUmdW2dgzSZ4xD
rL3nwGA7AhdyAMSJeutxTH8tS+nQsWvBE7VesQshfRYxCIb3ybWa5p5loUJDd7Mz
NKdulzTBv7WBDHOwLwLA95qOUZGEzxYtqdNFcMqrbwSkSn1nPb+EBboPVcl94hhQ
5DTAcJQ5+BOONHETN5wKApr4rii3SqagKV25P9JnzNsScvgA0GQYevlkerV4YAEl
1BLasKDEx2rigLV9whLJeZDJh+aWs9Glvq/A8VysyngITT8IW/iaHnt9WpbG7G22
EQb4TOIyeP4pdtDpT/6/65qM22CuducXIyPuzUOa0CcfblTLD9FXTRkxj4PJjjf1
l4fL1ssMLG3R47cVPeNiHLUKfvRSmKWTNkiE5TX9lbVf3CHLTqKgmAPDDy/ECkSs
ODeGCd3PH5AjrYGJQ7KSDALMw86WL/78IIfzLf527wXUzcyt28DEDp5lT9tMpIEl
LDS6GaKLocDSp73UZtobEaflESiEhbAYVOuDKk6mzQY1TLgq947nzd9kQl7In37x
KW165h+SKcf1CStcYTIBXDoo3eTV56zdiswWutJW0hTNc1HoWhjQzAWdXOINs2Ts
RBQZnL/2c5ezE4j2sM7ZptFEjntSDOYpYzOt/JBp/2uaT9wJweXGZ0e010ItXdDt
bkEpr/qyTmhCPLLDXwENA9g7B3IYvFD/04+9WMbSVvvAlNy1glQYzmFlF/aC9Q66
ty5YSZUYxqIZ3Dc1T+6LrGg9n4q5d/3NtlZlmJOE2L8ycN/CVB2idtPfBv+JmYH8
1hddfr8hPN+6kUXqYvyzA7IKVzi4k+F2riYZmeAsbSaZX47dweBLeolGKncaOomi
MDlyJO/110WJ01v2CxJ+ggBhYiZ21Lx1RxVhyp1xiLT3pHT3O21Ti8jK6VX3+V9r
hi5CMV8UGUVnRge5hT/0r1JQKR17E8ePjWOD8WDS7klfsbN8Z5fRBCDLA0SG0gji
Zs8v7t3QTrYwh7FV5hcqSsmrYdDPXbZ61cbn9VRVvL8C4gXzR3Dv1ooMnX95txjJ
IVQbBX1c3uSLT/sX6LF0JUN/gvlo+IvRJ/dGYxxIBu8+x0ITx9IHAwNN0b6RoNKL
klqq8JD4QmZEk4ODorutLMvLpMkF9HJxAlx4Wm3nJv4r73ch6sevcuPZO+IW28CZ
2wjxvq1byy7AOusk9iNQv1D5cvvgVvSJMtTAufQXB+B9RbQhEEqtB0nP9Tkvungp
V5hHVwfg16MGeBu0+1ympbTfo+Y+QN2IYtOdMIhODGLD3SorkULDyyxGjN8M3rvy
61CRsBt8Auwmu/LjqV/QqC7NXvOIGTl1Jl27j1ZIMwRUSzFilXCzhQDgyUvZshha
2NWID2Fl4gobURfSgtUBdjlk49etTixp+j2Zn0ub+SfElGGeEU6q2VrQx7H8RMi3
SiNXP2p17kUKc4qSqWE1vHuqIclbqCOTuq/nyA/SHLzaeAoLnm6G88abLvM5HCVE
bqlm6NQsJigya3z/CDH8tD0iGjwdWZEWiH8ycT6n9q0kLh4xyPAq7ExCGZ+nqJoD
Vw4Cvgg7PrSvUoyIbiWaWkrCQGU32SvcP2Y2iF0DImy8BuOgKopoa8A38VJeWjC6
1n+cFfluC1QzMay7MlpM4atekeCGVYNTyJHkapqhi3hf7IIJnpw5HYI6689L2HS5
KVkeFgLPn5Ii8wMGHKXzc8XoCfbGbgIPwQiRHggOXTdH21Cvz08Ggf618rAB6w3T
tT5WtzTRBga4jz5ttDBivJR8ie5eoYBMIaAGne5zzEj7QEu53ZkxlwQOSmzzmbSm
Ro63NwsSfyLwkqX9jM0qhEPR2b4mmpivcN1lY3PFcBzwuYPX1dogGyEQq+3+WFRt
MmgrAoxjzbMjYQYRdXp4mnBu0gvuJkermCHzXPBVNHeoYCOLXLXI1c8PetCOHpeG
3BTQYKhRN+yAwylmh1FBqi2SPaS0JrzshzKlGAm/jwbgN2LDlIi6JmRlpkpyv4l1
zB30DlcRx47jt54uhIqKjyFHuuK31g/bcShb91qyfVP3pe45VM9oABfQvBxsLLOw
Y+j2hUKZo1i9jCqMrSew1wExT7SQjiRX1Cm4hSq6bCMGNEZwuNzoM7kgXxXUPxW3
ZDBGgYv2OL93Fii3nMx6XgbxameOrU6o61mjntZUAYLpHwTcc/npQOA86uZYGntq
PiALkZySoOwyQBSTlmLXZ/gfcCQCJsq9bQXwQb9Tgk2X/yzI7UlEmjAg7LPyA9ay
uuJ4A5AMrOtUphT+aJE4dSdkQABVSSCcwGHC/WZaYzQB7wawh64nx4tCfuovsgDJ
8w3m2p/hqdzAIbfSpJJabXp79THmBDOgJFahyfqsxXOX3PRBJ1jcqfz3XAF9Kf6e
nPomx7S3IiFaqr/3YKpshQPQBS5155pgp0q5EEbZevdn1+pdPEfbVkVqCnYpGF+S
beVk/ZdjEKTJUfHf++baAIsDzE7NqLoXBn2BHo9psK6yamXjrsiJTzUaLxPz3Xw5
8jmCsOD10H6EpzhuxbL8F5ONK/SDa06qioLsyP+cKTlEd+IByBNu6iO/E+8JtTEO
qfx0V9mMG5q0fDNSZPhx0ZSjM2vOzPSfjuvHJkVZZ+iCiyzSdYr0zGwd/feE1tUu
XoGV7WBIDQZyDsxGIGa6XmxmFJnwquJyInBa4UX0dnajhJgE36qGOI9ju/wg8azH
xusp0moLBca26DKFBA3HrC9SHM85GCpUTg/TCJ7jBk7d7BEB6HyoFtRz+ONKwOOJ
9NRqcSyYOuLw6ZDwJWEytUedaUlDQU2ozPy75Fyz8AD/meInRlsjF9oMS9pn7c8v
PtjWVyJ8XKfGV9hM4LtOz2jFs6hyNTzZt8VJ33cjHefOsIyOjp2S3PkEny4BXjvG
gmLk26ORvCvTrtMMDaP7hWJxdYaQn7vHwbYJd54+SN3w0+6MHlhaHrd6/qO7wc1o
ywB1ocX3q+G4UIk7mmvdcZisHf9o9XcQwfMgerqJ1uKCjF5jRYNxounUsqTXCcnp
X2YNwsJaw4FUYaPx6v8SjTN4vaW5rhBICD4AeHDUl3M/8YI5MTHvTMPAF7M4HIGK
aH0H/szJKnJWSFzaxBQna12rZKaAhkINLV7U5n1cIPG+cbgBCgpUSVP/wZXJ8IrN
IFEc6uTnhPvezUZ7IlSWzmaZjy4/5j6Ud+5jWiK1h1PTA3vTxu26Q8XyB5cCuhuy
y3b2TVnX5uQy8+MA+xsBj6T80PB/J+PuumVPfLB2ZsySaPdG1EsHPy4OgGJqhXpf
esunCs9JEuctYM9CYWFsEQ9KyUmQyWuv3nWWa5szZBqkUZoITzAohQ9kolQjzqjy
Ryz54FxyQ1LwQ9IorN/8LuEAMq79TWTeeK2WxqQZuJWJSE213XF45/hMYQJTlsNa
+ukg5LkX602joq0Cy+uKy/R4JZecoLoXVQlh0MsU1gNVlq048jC3nViASOX3wGSo
Ybe75SU4BHeBlF6lnZGKrGLQqdeN+u1eCMYWH+cYcIBX/d0MgoV2HziWUAOcY7UU
Jw+cn43CVuCW9WHwOuRsHr85A9MlwyE/yjXaVc0MT+rUxNLKrKCtW/JshnsgKftI
+mdw1/1oFqh8XpfnN+B9EgusLUjINWksOxA60QgZNBunptQBu4ezR+D6wFCz4402
rRFavzMXp9vvf3jv9Ftw6dCmghYnsfK1STPrro4jIzKCHOwy/cSVzCv0MaqBbx+Y
XJXrp2B1sKWCi1IpoJewvxIRKbTgRsuTxrbw2Kj9QbBk8NEudjY/cRMcQVtEo8nd
XiKmJTzKd+QhVB9Ssh8ZcpxBbI4yq1ZyfHAclAMzGqcGD73CHVQmR40+cWw6MyQ8
HyHnv7RvxM+A9PGpHgLZENFbQ/tiOxVu1F8JP2VBf1ywyMkcrQX7L7zgWQ4ezVAr
EZYHX6SNN5LxsrPZbuhywoK91U9y5Wt6E/JGOy38MOk0pq4WM5FMi1fErPXtIMaU
bOaeMA4TstNMapsQSLLwXzHJ19hKRzpn7SUjBnClJWGnsL5tTqo1a4tFR3/GSxwu
TsfwUdZY4D1l4+hKphEXROBqyxlVkxgeXCMA8YLB3MAKDiq1os9+1W6mgEOBYIJ+
F9z+DQlFIh0kc9eAjBuw03IYUU4w5+V3puCglGMLISCPIyyZMSDX0sc4+iUaWZuT
6YlVguU2+fEVtao8qlz4YGe4i7LNAZdYqj+Wcg/7rnwjoM9SaZD3AWa/ENE8LVXS
1uHy5oszm7tXhdjVH73sM6+ViQaX/iJQH+g6jUc73LwIOsdS7IWSOEK3k/hFm/44
P0mE9qqMM5m/ZjUaLKQ1OXeHTHBh7nOysNsE+/v0/Iz1FAFK23kZoLUYEoMRxiuL
vb/XW7WbthHg0Pdj63z+Sa5eb6LGBEqfu9Rm6AZ3wDGeKzpesNuLZO3PxdnmfqET
+khFhmfjsPhkUzRIzXkEyFmLay9YHm0Qf9hUb9fYo7Km9KRujjNt5eM3p3zkh3og
898+qLevD/6bKdNVX65uXBSC6Vv0zxz2jT8IS2/eHM5OWILcbxbRil8DZ0+G8Pgi
TrFcDxcDBRMvKgfH2fsd0A88qbxEokcy8VqX6oYn7V2dwNZFq2EAtCgEsstAmXge
nVq2H6FD3ka64N+zhKSctstP4/0fLLCc55T64+NaAG0rAtmvQGU5rbxKLtJlOGi/
SYzeFxOVGnUAq9nUnbOxYgrQeBm44zslQHCjBddzpnKiI5cp4JuFiuryrg93Mj3+
gmKOSeYaQgIikiwXWNJr0hwy3UaiusmhZDNjCWXyj1+eh+BqUS9IlGh4lhNHh1V6
VssETV+j6McBE4lTqvQli1g9AxkyFdTUhgUp1veXgyFSgqd5o8C0EkzuvGnHNhXX
JidnWur+dQjf93cx/n0bsKyd6H14oT1iHbH48VWM2zyxHRhdikK2DpgsbPoZa66K
4LXtCqAZW1PGXiDAYSuS9mxYJ4dkNiWKFLw/Z5KP9iF3nWkq3quOX44oG5RtY230
XhkHVckHuuE5TbpouMltVMLfklWQrnjKSXlkMpzNUnjwyFCgxmKH5uw/EcTnDYCu
Yfe20QsXX1JHEgARr1Y+fvbGi/ixbNU76Uly2GsW1eRhbdNcyIK3cJHOBZ4bNC7W
4XM8JaQhgs45Ez41Zm9HigHFz6Wko+tJAN2l8QZ3Yw1L9SkX8x+Pw+QKpTYtFRP1
rAylPQExDHf31dHVfv4HL5/daeXw+rguWm7r9OpZXTf/ucF6H90sXYvgSlBS4HhG
FXXnpuXgHm8wuSVj/bbM+ClzDTMCZERIWe/mMMmdhE+jproGqe3S9+naxAb0gIiN
lKCLO6lKbVlhhuzPGFmSwz/SysJwSkeRleYRqysgTBdP/C+Euk26IKMCjS8LAAEj
XesUIsqr+/gJ0sBLCmIaHsDGDgxt+F9gWC0bUq/d+6BGWqT/+ZbvLz7lsWDpBIya
1NpvfviydE9u96dj/Nsd+3T6vDgSMVfkSBwn1iE21FJ4mb+fZOrd51DwMVjC90oW
+0565lidlvcr+Gb0DjzeSj5mbNdUz0rHZyybDOGZ89nh8c2+GZ4FbbOWxAwmmDAD
3hXdto6zvxe6sloOOqAagwkLfhnmnYu2/VRaRN6wu9m3TTaO6aBik4xO7wpVvomK
lHLbUuiO3s+6ZKwgkZZ8/qnCCFwSlty0deMFtulJLi3nq3vz3VF9BTKSnDXuCXyP
x1GCu+7KtBhDzMBuT2PGJJLEt/EVg4GQ+UsQdasG+bvLWKoYnXftjhIh1vqC4Efb
Rfj7PsjUmGtRMK9/Lsc9iB5/zdjK+/X1YR9kFIckJTKu4RltvJufBwFVdm7jEnGY
IRx+WF3x0k6vtMY3VGu6i6AAS/kIfcBECDTNfhUdjTXcqGX5d2q09X1LUtR6tpxs
XBPCIEHF+F7RUHoDtxTac1ROBqBvbo7Y/5YfWIfnerzBCp2SXGej4qLdfX/Gs0/i
LfRxClw0AH6NDcAtzn30Qx36bz4SMtNdJjL9IZVhNrbyeTpGZzgW/p0jQgUGUjy1
usSZVLAb5bdJz5+kdn93FBVJgnIpunzLZwNsigxea7VGkKygpopnro23kyihG83I
YK6GIPx2yaA4rrOBJPS6sSN+13eEguHTSEefuv67nKfUpfk3z3qN8S2sEuFOUIDI
RKijL+BXS85fdXe9bZnwc7C7pRiFVqR5lxT/rswYCsEvN2VlljkL033Zyn3tLeAt
0Wqssu3gJCONskE2AbCrxdG4SuhMxAGKrP/wgfvFD5yzIZPZDIYAQBdsyJRSRpZs
ks6/buCt/0xPiwKRtO/6l/cTNy0Wdcw02oMK53UbvPkZ5PNCFwm9dIcO4/6Oiduj
gwSjt7/3jAHmFIsWrFA2BWRwNvxgzI/FW2N1DjdwusW5qsGl3eAH+jDrPuLIgm5N
Xwd9Nau1fmvZEWu5b7I2KUCPK0YOi4JKePhi9k6RYKoZDL+z6J+ZneBw9t5YGf2J
Tia16yMbcRCrqoOCOSDY/QYRkF/gJI4201r6IwVoaDTfE1KNijG0FlMcFI6NYxSO
nhQqp6/VhsH+UrXjq16O1oFJlcQVJFWcuW0PXBlNqqC3bp8ip7wCVrUvMjVWxXi4
wpnHACZGJtHI35DmpM0cV+MOVZc3j2FK92XvXb5NTjuB0fMBMT6zq6EIpoN4HbiX
SOyABESr4nnw7vYDVW9qi9gGww6J722u2cLjDc8jQVBLRGEjOuePmRqCN7ywwb9b
hCRtze3bwm6Bfk8Ct5wTCkO9GfbDy+tmwzgXv24ueNrC8u+Q5tVDg0Is9aAQKP7j
Kq9dN2FEDplbcQYe8q3Wc0BFRr2KspN22xCKToHCSkBViEHIlz0PAFtMq1r0xmfq
Y0dl0p5ok1Iylwz6Irnsdr+OPWD+N8Dk/AjLXnnmviVv8y7mz0sXnNcO8bCAgf3O
9hB4pA3r+5psf5vPkgurX57KkQ0iSHORl0fBYljwGeLs/lvANj3eKcc9NuHqVzND
i4JLaBBdJI8OKKAlVEM7xV4tgsYThjzacNcenBWIITTy1h08zVTaZMFXmS4/lzW2
dIbANZ5ZR3YvH2vf6lAHtQ5NKcO4eLRK0iMcNuKwUhEIqA5XwFsxE/oeTLghgLm6
KtRUERK63fR50AlVhNFEc/Axwgf5xuzVZayJaMKQ3Unktb0jaRIbFegHUNkrpEBi
Y+URxrmzMBCKaqxZad/tJTp2/QHFHHd6MM6VHqaZ/C+vVwaAzZzenrGL4LVotjrb
ORgk2KZ8Ud5lzhqFp9l8tR5/frJXnL8RKxLn2uEA2Yi4dZpxRIy+VLiW0VFhaxCD
iKC2YYJoBuChjvGkA3y4iKZERr2YvdAhSnRRfZEUCEN60squrM22CMcz2DU26Vpj
pv1xyRhieDikWXiTvpsODWyapIRkaQ0haMnxaOS2fkbFnD2m0ONGK9G5vISRXLwU
IWOPz7nK8OU/ikgekB5RjqAhwvfHRYcOudEmTm+wtSU71l5Tc+jIg5N8NyXfPLHF
/kqfX2WykzXZfxFBiPt6b1kl3utkZkZufxcVclBm/Mv1D49I1zMOhGstWZno2N3b
Dtg+XHgxBlfM9JtSSwIdCV8oGZ7O3ZQsFSU2tkmpZytXdeSX0aafDfUH7JY9C2Ik
Aomz5e7nN/CX2b9c3vEUMybtREaUaSE88EvVEJZoFalsB6xPJxMBeRMLZcX85o/g
MGLq6HzA7DxPLhH5uvI5rhIbrsiqcxTt+3ko8ArmouLJMmY8Jt/i4i/dRRVF77dB
fweVCrxTlFHgBpC8UlQAhXoH2KVeTCeaj0OcSiLimsLNNrQxoYK8uggnQAH87bSh
mR+ZVvG5nCm5mU+DJIItYerkU/4lspKAuUHiIcZ6N/o9QssaYgbIbxOJHRbDHrXn
kB1Lq16pmLH5ReWHs87UakPocdE0d0cb+OcatsISVf0iqA+4H/0pve29eFqMA3QE
HRMKc7tS6CwVcNio3Ryh1/30eHIx/OLSHL9du3XRPorSub77VZFURRBuCbwZsBdT
Sw5rmmx9Hdw5s0QFc4SvZeGIRc6voyPC0R901/zeZiqcTxSTqVCYvbwlmHWF7zrk
agggnG+iT6Ovct7hhXQJTXrbGdqDd0044l8qDnlOEr2OJZs/9dyi17sDqmqsVa8X
K/R6TdryBXoEioBfg5H+NqGHMJORdrVdfFiuOp2ciEKK5iaSshHyy2BN+XxiLEwk
gysdFjFCykSCmznyBjVWANbMLAdiMxp/XdM2/fkwcI/qTQIrI71pS+079xX9GMqD
6oLBQ1+bHUAFt1hpIXdkqBf1a+SjZsumbnqKdSEs7ofXzBsr+BmrcWCxPmaFZA0n
OTZm69VsCVcnJLnI2xyZCSkjcpn9rR+wKukSgTb8P01H03uLF3M4A9Hf6kXZd/OI
QpVY8DPekmuuUk4V0IOyeacniz8T0WwiWPohed0XvBEB5SAAJpsXwgSQyoXG0Mld
rcrc5000HsCN4dMsPSiDJQ+O41huX1OR3c3K4DGo2wXY6yioSe8oppXiO31y9G3U
ZbJPgMwK8X4E8sBMauEeh7cha1g/mnQHE2sK5D32SRVWJ0P3NjMR8/bsOnwYEWkw
Iw99PLi4VlC6Tb3V5xkLndvQ96iwzO2ljB8YyPB8or/JvKB+vJI8QOh49hO5UE4A
YTC5nkDAzAuNeza+aD6a99FYy3fTDpRLFQutXd3bNAC8knE7nUlGiYyPRLVj1rMC
vnbEqiOLabnSZNOBN5NGf1GYHzrRGO88UuW6jGVuUpsEJgjZxNKegfWVPSjnaMQr
qjqhBtujwdlVvlRsnoJqFilRKPg1ntpdO40Y/aYzy2H46QYTp3qXnQPOeQVCZspd
4dG4hUM6YW7vOH3Wu+Ha3DtrG2NsI0/oRAfGFyXlnFru8HYforKOUvV9KB8KLaqI
c+1U23TO1UjoHIzBjLLCeaVFupTiWO7mSzGvXWfyZpL9yd+FUsEqb6pspQN3xWWI
Xkbv8sH64hGXxZFU4Hif+oFLCLsVBdeVPvduKlQhL8TxQ+YQPUh3DWcGZjKSGy4u
uEc6kFlcQ4x/8brUJJ3QBkel1iAiEXoptRVW2p9hHvoCOB0r4oSkGOowK7Ynch/3
6h14t/Zd9KVElx6acFpPnuvj3eY2NR7pJ9dEfoU9gApKf3Z33jlGGqUb+63yH2fn
hbeWlNhG7NQzIu0HaC7RBQAL0aH43xqyodhUzI9f/Di9q7VVOYHC1VCbQJGZALDq
FD3XiKbju4LCCUjVpslf+3jHqnrEjXQnXwIfR/Q9zVJi0hGihNyxMRInrFnG9SOd
CPD9cUnChAA/RrH8OS61Qfb7sAO2nREE1vXX+wBmxoXHeeVGOaKU4U8AMdvfA+Nh
tznesSODKwgx26VVxP3Ew82m+GOqQ5aY6PoIAPGItga0cnpNa4GhzpHgww62X/Lb
fzsDsM4NfKFuxwGzGqi1iFOY5vuQJIuAac+MXd/zMLiTO6jjsWwK5qCG9Qp1I37S
5bu/7XtBGfGcjh8Cdsfzp+ER2kOz72cq91v6jeBzBEZg3dmPs25x1eLNSvmVvABA
SYu7GGL+EgKbQCUoq2ShnNPq+UC7X99oLvHMzDfKKiSKTmPN+a/Q54bj+9sz5pZY
NCVaFbwV3agS61mtN3PDktWdYv+BfWh2cgNpeT4osJaDinLSEze61v8VTpeswhvX
MYZCKYmLhBHgSc7WtizMcVXXBAX0iBPH14GM2Uyv4ig5nZfKgI4hP7gooVH0r/ZG
y+hyly7AoWO/Ru0f5VJFlvUrSb+I7ir/F4Y4U+6A7YAeeKuRQ6GEAdl+kzacsrrS
DD4i3aRzk/YfyjEoMCKsy3zphLzuE9lGelGmlprk9xQFEDosAxZ19nL11HCwh98u
hlQT0ke6vGdid6s3cY7Cz3Gci2q4nTWl4P3OcsJp9a9WYOpHpBCTj3V7bie1TUgK
yiN3vx53P9e1sPXR67TzyBeqsaQsM2nwfK9XL82Q6zBblJVrEkq+fs8gG8/QtILl
N1ppbNpSjmd9UNzYJE+pncDRJq61YhY/ssQBQkdWf2uCOucWg/+k7EBJv2zu4NPJ
esqgSnPcUHdETZOBEsFKvYfDhzNK9ehlrvnlvO62w0EQV4YM0EUjL8MQE74HTx8y
PvKLGUb67ilUFPlPtfj/NfgqlxKq1SIDJqn+JP1iCMYtwBmyvQKz3/zckSKuoJBE
NYJyeWQRcTzqnbXN/dBDoLnFH4ILQF/8ogGQvqRMeeOqxiFK/EIcQ1abJkQQMXNV
+ikRX2AWKgnTEy02FGbvkEN94cdMX8P44/hiPbEKq+92sqE67GUYJwpvh5lGVeHM
zuBcCD4uWPBSBoc2TIN4W/TbihB5Ytts0IExKyjNCjW23nAuBhX0YUJfssqovmfc
zzx3CnZ2mgfwarL0TutUoT1Nd3LuFyshJiZXg61uptbTFyGoU4JR9Hi2VIkf2UPF
QyNQiQ+L45bgxE0Sv0lkrTHqp0vqFVcJrP19xUxrc3vzl+WJ1H/uuzvUxlp3dDkR
y0aLTyjwHu/mJ+b0U1IfXWeaQabL0n7x00AZstqkvgnA9LLbbaU/Hnh/LCHb+zmm
JtQEkajG7tW5glYBSqWteSPqnGPlQZwMGInwasQbqJhI3ESbzgp3RtvG90dBn9zx
8ci+ZuDSZDlYcAaPIjdWFIK/tVCyPb3R6S1/TTCMws1pam9f4GYt/bcazbRzkf1f
vwUQ6MSnxpE6MP6xIWwZqyJ4e9PmEuR87xyvLWbD6anqhUcmIub6E8f40cFSXssN
geOKYPVCuEu9X0mmzs50kGnM2C7I7WPiylexY8LVAbENi4LRsdhgOQnabz1SXp3e
GAHGAaB+DjMcTzrWg7IUiViEuWltWmkn9MxAwDlLkYCEFC6iVgm/39EqUZyUkERs
WLglE7mojqthCavy5Z/0ncMEGCHyJke59VbmXCa8wWCZv3nwRR1TXMZY7wl9O01e
sCOFjSbcZZxRQyud3B+2yc/emWn/mbsYAeAgm/5WY4pV4hjSFYtbQ67WLI8eYz5f
sh+cdQ8JKxHhnV8lV9pSzZPZmdjl9WBF5I6DFaW7IYCaPmmGzmlK52UQCVpOqOdd
oCX6T6DTGaFF32aUdO0eMvdAnVMlOcm3seMBTcEYGdEVEE0AMzelxsiTSaTOyJu4
BAIqRC9p+Z06PtBPTtJW4Nq/YdDKYVqyM8pcrftFqCw3OVXqUKA5AAAk5WPiOuhT
/a6xj309jPZeSVHRkZPO39yLhUxSgdXAzwSTFNGniaHBzjPCucaAasf5cBwI2DaU
VedspWVVCxKGCeVZOV5R9PHG67pYc/IfBGquo8L1jq3R/bGhAinNvsJG1F7Hgp5w
dwz8QBcw3O9KU/2AZ6hL/uh/e4Y4W5zmUPz3mFwMdTWX8Kq+Ee2+fTJvyb6IgIml
31r3wqtkXx7wwv72XTA4brEOWkA1dcW88S8KA36EM3OJGB9Qo+DidNhvu+AqxJWR
QeBVkl/bCRvF7yBl5c0gvWplliT47XNqoS0wGULUhQUP0JWo9afNJaeIcdpM7VLB
I6dTHYmfOVydTa/04Ra4RKMrElwfXyY9Fg9spFg65pInbiy/aRo7oo3iLrkg64bN
8x2jUYc5H3ZTUY0TrT9KkEwbnO8dYbwiY4ro2gAnWgrVRUo187iwcEmVJslMMFeJ
z/9U05hPh+lrUtVIo7Nw3/xk8oMNDXoEtn61kZ8C9aNtwA9ulUvUPin1DfOStrd4
Hi0+H9fqYEyXBQoZoBe2hI0bfoy+Qwr/RuKBWU49/eHov8psmi/Zo+EralMhpa0h
tU372kKvHhvyFYFt9RK99Bljq64ODt1tdx/soydbi0RLbeyPg1gH/8JvYqnZO+cm
gUdiezRQfbZSLOwsYD5WJA1pJQKiwAqsGVrwbXPEE9ge5rUhgMlcDl04yvyckbJ7
pmdvhDedmJmnz9XI/QdSBkGkyt4Hi4OSFEIVq1b7E0btOa7WeODUrc3x+ANmxN5R
JGpwRZEHbj/4kcnUNhLt4SYyGuyh6iHzfpdcG1NJ4a18uCwNgo1MDAhKe0g8i1PG
iYWRAdzq/DUAiXRrfTO8hllAX9pOz/Xjqzw/i8BDdb3Wly7nFOKPE6JpgGNv2qo1
vlSeQ5pZqe73cz4xTFUgABWIzOCi4e+CpquvI64a3bTc9P6zlp4RuT4R++2D6JzV
HG4OUkp6QGLGeHIdMWSRYOfIdhN5I0B+HWxQnvC3Sv0q5Mfc1li5tZQ4Fd10EIfE
UGEcq1G+vV5pWoaTffVG07tr8U1khDJhc1Hb3Lu5135QTFwdfY3uQ0zapXcarz0c
zFv2HU3BoTJqx60Gt8uvz0yvZy7JO652H68x/VGHg8yYQfOZhQhMh4JptVe489b1
/hUSoeXQXqM+pT3e06SKXg0l9+ogfi8toHxjQcGRhh+o484AZI2Kl5dpaTpZIYy6
y9FrnwHSEcnbID9ffWp9SoAo9Gne2xAvdYDuYE/ehOGBpP8jyYoE+w5TLWbcbb5d
iiufQySh9BhNj7z5k/YOwUejraCMZmIXeQYFIgrRiG78LHws+0LbyYzcrBWR3Pkj
Psi/0EJEHwnaGf+Pq5B48afPe9XasKiNYMi42vvnBKmg+7xgeN5xUTGaGuWT3sJC
zesjeDcGSao9m32eMw7Al9qMAVd7ePtGeAsUh4QP9tL0FQCucceKI6pS5eG65Hfr
OojehArfl0oWua0bQIn4LcCwRppJly9JnzO1/YZvKboLZaRVwT3tNHx6VQTyE7Vi
LR+83a5EKtaSePiIFf0+mVAPLJjch/Izk+IrG2SrSkMtAMKFMXsvzaQ6slmYhVzq
/cgl8G7u0/8RBwQ2tv7lEauKtqZaLH8rg+y/FCYM2uhgEbeup3VhHG0IW//eJsHg
YG7q/6G+ICARRW5YEgmXbXkivt+GkAlFt+XJoek3DdQDemc69Q02y+TG4XxhH6L5
Ys0UCE1j0lsBgPUlLKDkcTl90VOI5bzkjaBg2qRO3FJUON87g1dq9UwEYL0wQznq
kcforFdYw0QRL8XUMQxEC6dfAnz57QMF81KARNyxkRSdJsqUNcNcnsnW35Mo8r9b
X5BkqstSb2GK4vREBrzFxVs/JApcIQelIu47hEgEEy0VRRfmxBG89YdYqDTBfYft
ySjB9Mje7FWOBcllviRdeufYwFbyazVay4JtCfGSssS8VHic3xVoiru2jCePdY84
L/zOQEIzBkRXHDAZP6N3YkGLMFPk5M6KSPhpJhqf6grLKYxh71lzPfGE05F1uAVq
PMetVH+ttMvGN0Dn90kAUG25txr1LrDyhI5h7xvd8A5gxD7Ichd25lBR/5N7El48
ihE+aCX5GEDIT7ifxzNtfF5snVjtxXP2yeO6KQ/fWq6rbyNVwBDb/UxIbd4ft3oR
Rzyk7jnGzuZ1kP/AuEOzR6rXXzDoCq0+g5BjPu7CdsbMBhRizd44mEL+PqRsrpbe
hGT1dCu51pD49Sxkj8vQVbllVkfeYUlZIg5mhPbgj48LCVFhg4hZjXKfsdvB+LUo
a9XHUPzPjTrg7U5Oj/513zoPjyv9eiSSUzm7aS3iLa61zGPwz7CChkmY3CqSBYTf
Fzv4J1IQGbY1x1nj7nEJqgSuGGSaBhky2CdSzICZ1LQIAnxdw7N36/Yc0CpSU8Zb
Hc0QgkvtViSC5cHs3rxFvtz/CzRk28LhnCgaSJTkhZ0/vIV2pRpS8bPIDJLf+5Hy
/DVyqddNRru2oXbib4jTZNI9ds9YMxqgeBgkrQJrAxEOTZSxSPFUniKX19b8ejhB
TO/Jyuf4qUPqI4CEbpFDN/8dE8VsgDqAdrsGUQaLA4gEgJyDLN54Yi0WncI8TS6l
QbCwd8iSaczrBp5tSy8IZaQYeQamUPX0XcCYe+dLT+4HN8z4iroRcJIkYS38sJWp
ctsrLPKa98RhxuElTDCCFgIBj5/eWwnQOzES+RgEbcAR3KtyGNBgOEDeKcWDmFUN
V2N6N1fIZs7ERFClHmbYH4EAcmuqKG/wGqTcKfqnrmbkfOhcjrAuRCaIa8Mp2SEM
l7QECL5+lU5iWmUX3b9YXf9wSZeHq9sgMQIOaF0ABi6k691K/GjkkMkncpANq5fR
OCxdbRJYXoNES32Umjfb4kkbzW6gezoTUAG++JAh2xs0nO+qCdZz+slAfYqKRpUm
ltk4Ao6kPoJ36uNeSAeN9oC5SfkwPwKaKKvB0MPiicn0Dm0JzflgtkOPJTqIcqB3
MZLTaws4ffZO9W2N+zjnkEMJV5plH4iUZBTh/Q3UHAx5NqyrngneI6T3Q3neKDae
ys0RJkUuOs8AGJC8VEv6StiE0b4EdzPK7p6I9EVqEnNFy8NS+6kDQRIDdAqMC+SE
M/ceXoBnNciDdfVLsEhrD8YGLXZSD+nIbSP4bN2MqGxY+nv9HIRASEjpTKLccB7+
wsltXP+eSB81yb0KVCi1CCKV6mxw9btSR+TYVHDZT5zi/+0nIzWOeLB7cSW7hZ4v
83eJg0s0zwtx9Xi0FcZI/xpbCCFp5R41aFlGU12r44QCvm10qlIFbq/KWvAPmtSl
cwUDt0nb243d3TTL88X6imzq99UtwlQmptUXIP+S3DuDwApzLDBSt6rvBXftxJeE
g8HV/IUqfYHsmAqS9+e5crNQ8n6G06EOjT3lf8vInsRbfeN8LyicsvZGrVG2VM6t
FDZ18/ia1OrOjWcASHNbg+pJlGJZGBDUoY1mw4ZQMAudG43OvI+fIiiTnvyZ7U0A
aEXbMnmwiWnwjDSz3u82j89RAK2cPUXATTKzdywXNZFFdaiZh3x7yjLM2vK3/5IX
+ELInAapsD8fkmvdmTgqgoEilygGTnEZZc8JViGgQYoUGM/zVCwKthy+mgvwnvC0
6af+3GUvdfJyYggf6yT+PGH8m26NbmHS9Lhv/X0HsKsixGayKhIHJ/nLdfCjCDXu
dUxi+gL/jjpOX4xfOdHvNqYFtkm9/FmhaVGq/KqW2O9W7BYP8tENke9k0cZcxls0
VfrDjFTMxTmC7PY6vvje9C0JQUEaL1csGcjfCDPdmQiDLVuWmy08IZpT0tDSCmF9
6JoIAxCid2hgL89PaLqrr5pO/TSBQrVAuM81DslbkALe4MbjocHBb2rPirKmrKRo
8Btys0fR9S8Gyxc/OhoV8dDDtDoMQXIG8VnX129Ytz/F3hx14pm82GFXEtp1DM9O
3SE4RBT11tx/sHBLVrgp2ZEb6s0IkehBsK4s724scDgrudz4Crxmgt3I5IdkM/J9
NYkoyhf7U6KVz52O16kWM3E1On8tza0SSRWsDeTIan2h7enN9lWvaIA0Lrpc+6e4
J0EZmybot+EXiDohRlxiTAVl3vVsQtCaGnsZfQU2i7DH6m/v1euFiW5ABMh8ZnDy
9JZojDbF4kZuKuRIDC0y+jcSirL3xRA3yjTTSjghmnP5Z3eq6rKQHVkdy43/Xlr5
8l/R426qk9DmspcK/9jTb1aXIygqZQ4xgN1c+3mZ2kMS0sheXJwYiguJtfdnusdJ
3jQkxjX59/jJaYzQD/kc44JdLEUt1IijzUCcHBtoD+dsW4bxW9ShLWxKB/TvoLVf
Y8l8Vj+XON80J3jlEMgVYrUROzQfpe2xYgp7X7ENlssSZ4Z3VTy+SGVPjumkd1x5
3/+2DFbgcAZYZnyshLN8a5BllCYOsvrpYtJlqzwN1W/ylCECTlSac3P22kJ3JApv
4PKgJFndS05TBK0boBhSGl6zA80+04drTzuDHUkxmrzF3Lr0RWA/ZN2Wzh7dTqV8
n67zZfvwyA6iy86JfmejXrPj5b6PFhNOv8fz5a0+cWUxmeDhunJgnky+3RbenmvX
dHs8TobaSB16rSGS1XhAugYYs4iUr08O+uAfhAsmvL5dBO7iqrdjWu02DCMjg585
fqAIQ0T1XHJD/iw4kzayQ4HcMY141uKZft0tZ/+71rKvj8YB7XjqiFsQvwUKS9kw
yWVP4j4LzQk6cDk2IJMouN2uOT4u0hSH8WGAZuNgMxehmcoyHQYe/9zW/A7IE7PD
8tOVdFBWmrdGg/kY5PRkbGbGMdREeFdI9JcmPaqnrHenEgtFImuaXs+/nacoQIGx
uaeknTowodjqnjJfw3mZidWv7tZbGtjs+0lVQ8VbguFyu5sVETy5IlvCgYjTDA5Y
a+wPxiiUvCa0PNXMJNGdQhx4N0MICxc+vgwSS+d51Er6UyV45IYpVXWiHWpp7EMz
xiXhh/2kIRpg/c4QuhjOHEwlgvULOmawSIiT2dvdYELIQbRnYZ+sULmq2N7HD1jw
OmRRaPQFTCf8ngq5YsXBQuuKoGkKi5HfnwaX24HCdaDOcnav91GNOE1YpSZOFrIW
n3ikVorgU4cTG8j17c5guzU1lqmgkoL/9lRSt1s/Z+Kf/unPjdGqx7MbYil/jKie
/TmC+1H38SUCfZCt2MfEWFSoUinX7CtiuPX4DkspG63AAs9kFmvD7MF6m3aZAD7j
26JWTL6a1v0+Odg4OuM5hsUzdH659lihf0OYOn1Q5vD1Om7lJkF2OP8XVJWUP6UK
GIhGztxAINXTnYNC9KU1jip2mZnXtJ/9deYmelZeBKTevN29wCJCR2AREqslujnv
NxJVBshx43TzHz06O1BjeZYb6MIAWotutBjam3NjyaOfJpzXbao3QSj9UjuC+N0q
eYKDeywHCsROUIyLORStDHVGGsEib8466mPgnj9OouYXIeDE2hjtcdDY2b2ekQJx
KH9TE5Y1DunC+MxGa0NyhPd0/+G9TVnZSO++519OH2DoAqu9MluvXmc9ZFSerDGa
MumxK79knNMFrMorNVbKo8DrvKeTSkRwdALhB57RciHHymeZdC6Ssqn08cGhrXJx
bqfY7KnLPlgIPVgWHz4Wp81W4JtQQTDOak8elw5QOBLz0CzYUrHzaDNSvBl6DGfs
SVe8w9Z5I0mSRyLXR/guEwqQsU/vo2gB17N0O+hqDb9YhzCsUB5Cuv+xvdUZeONE
IxwwmbTLMLeHNUq6anibR4ek5Zs7p+X9QR1EdnLV/VhAbli1THC8bYdXVy3sWzQQ
pNneKEg1Z1927c2mp7mqvYzPTjYCWMpxY3LELVp0WGVA6TlpjFmf3RY+IlQv1IAX
qvU5B20bz67Jz+KI9QAd/alXHCShrtI9S+K9vohs0r/5eobfs6IDO8YcA6dy8bUP
jdTxzUZoGD5IeBhbo94psJCg+p70FGu30jRjFcqUWzH63BD3vYC065cyeJu3QwhK
QUEuZkEu1xHoeKG5O0XA0tbra3aTKFiebl0HmyVgkeYxAnE5xvwE6AWdj/EzQgAD
cgCn80Ri74VXlSrnvpjtlYTHUTNhmec+nVUZv5iiuzabYFXS/nUeprYBdDvy5MK/
krMp3NZTm7hoPFfM3sqh+gwGVsObW/8QHcq914pehedX1fyWCPb5atrxuve5tNmv
qIOWG6n+PCQXtjcliTsN+9rlItOC6RL4Gb5zoFpUdB6GyEhG68ZKuWdCJZkDR6IS
suAY8wkiyRX6JqVpx4PjTU7uHpy7gwF841ycd8qAgzqsMuOLUe3bU/ONbSwD6TJf
P9KDdX+u1hIo7OM7ij+xlkhgWFwZ7xFUUgm2vRzmo5QvxRXvgjzYPEteejFcwXZw
9W1VHqCu66FQBYh0MoMXnLSucCoJzvjGo8Jckfuz7N6fzAV7lasywPj0Ybr6JPyu
/uXXimUNKSVoPyliq7DMC9+xe1VxSuUku6vqHE8TwEk6fGylw31R2zOGH3vWq9z0
Ehp0tvZwTcPZMgbgcbakSEqUSlzuZ1BBKfUj9flfJPAn46OzC3QrWtfif7+1paNo
S9b+ouTV7ZMNqmvsItu1s/BOM0iWmio9eVV0absNvzW4xZyc1Z15TZMNH3Py8YKG
eJN69yHbddJ76PnI+qdtPnsp91v4IYl9E3ArEX5PbkrMvnu5pKbn//8UXAxacO4n
LOIivln26KDZs53B2RzBmJClN5MnHN6nXFgjBQCr5ulj0K+Zuy7KpnTkZfuVyGc1
8GnGY9ad6V3nrmN2DBQwPxRyi5t8/WyzpHuhv481c1oDuJDcpPNwV6D8VPQ2Z+FJ
FcSxowsXdy9eKz4swDMTDYVYSmO98upwunICWei/k7N77PW/VjwzwX6CQdTZHGKV
+d9xvXaks5QtClXy4QAczByNYdFv0HGLDGvDM/Y4NK4O+2TxcvWqkYDchver5Rmb
uvNhXIFNIDI9vPhdFgE8CDGtuU3WoEy1+kXO2ZGWpq8oOiWRNvNA9L66yA04RgoX
zfLgezsbqEgN8d/uXWEdtXNcIy/9JPl1pjGjPs+XV8wPhMVubY+84Jbb1JtM9B9Z
lyJp9gv91Q6lDkqfSnNAtaLj8QYaavwb8d2AqAtp5T1nVNLt9Aig8HhZkiMHidhA
/RaKErtG3CQH/dQBOhYOBkUHSsN6ye7HeVFsnYBVHYgAH/fpxh7j6cEPNQu6kuXc
6osjoQPoEsoeixM8ETu58NmLgviwt+3YbfPfvLsaDaRShVzAyXpI35/DL0Tnl224
z8nVNgkX0PGMxatmejcoO39j40ugLc0ihUfSYsaiTAabi44KfzdskRZJBHWk9XdC
lRncU0Okc7qvCamy/eieAVUYMnTDk+HpwsJxGHBwrquNp2/0g5SuX3jZjwDZ4OVM
DzIYmKz9iDzc3GpnahmtI03kr08tlurPlJQq7UNdYuZ7JMnjgBRCPDJHcSWWYn8c
QXWmIJZ7MAcNKtxXtmHDXycigoH6W2RN0of2yvU00kNKiZtfrP2bI3rA0cf+1xcq
exwaQHNtrl9U9H6lZwDS10byW7aC77vTwq6wQNIOi7dwRJgU25TjiURNMzcgFzNq
kQT63TQuVpCBNcYh6RJVfnxpCA1O9TW4/due3c4QskbTuQe4N090hx+g2zKKBoQj
WsPKIEukBJL/bvyhS4fTMAqmGUGsZxWpUc5hDHt0B6kGCY1T+QFJchMDbOEkkdKS
Kc2UwRweMlV/ARUhPlmx+rRvWYyOHpWkc9lhz5dAAbfHHPAl5ttubG+6DyGnQ0OH
0aN9qmpDAem6nI0V6y9c3rtOEeQivBkGMegjPR7Gr2prPWs3DK/ez/gmpcTx4ysC
h2lue+016YuP8+CBLQkZbtiVy/zRoh1YMY2Yd1jxvMS/MJFXEp2osDD6IttDYAAr
YL9ts70ZHN/IO1O1kt1oWKZtXwuDdwjiuHq6gy1XU5zHb3nyLkRwLomRVI82343T
xFbXIZyZ6k/XsQpBC2038Gky3QUD6s6oG7yv3pAgOz6Z+zcSrAdi4lRaDuURTRir
/0Xh93Ts8ipCvJdeEOp2vimQGLYuXkSem2kPWIEMbmE9Bzus6ycS4aKKb6VcmNqX
jwgs2rxcochaOadkEcTLNxs0S3+FkaMuSOox3O2K2gNh6TKdzn2DXrNdH5+5zAAm
WSRa/v796siTBUIDAwkXwRhYmy+l0cAhK4hcrkDKiwWPt4IWkh3XIz/0ANU9Q2oC
4nx1Wk9kstRN47ZwSfb93z57jVVpWzgp+c+8gIgzYwcqFNnAdt/MbsuezsZCFZxF
SnnqroNV9bylhuCh7dxbMKhMoy3Y2RW1MBlTfMPHdebKgtDcqG+2nsEe5+Jdrypv
06xE58wt+KKXcNKQG82QvRNf49xRr/g6q8WziVMqBX7K5yx8jQ3H6kdquRob0EtQ
80FqlP14/KOKIivQ4/8NlVvmYLezX2VfLd6sgPC81SqB85/I7vMfr5pcnSR5iLqB
MbLxy7wEA4JYhhqBnoT6HLFEiihZFyUt6Cg7BVeMwE/wlHm9QhtztsQ9PrMRSHoy
rP+32+Dji93ua0VAiAYJnfYMmcKYGv2b79sqEGrUOeZM4C8uQ3/6KkntoYZ1T5nd
YFv/cHElI4gH8Oam0vXghtSf/ecP9ylOiyE5BIwbw73JO6BJRMeUToNkGUM3Fq0m
MVPYeeaZ7LW2263UPFRmJ32lDS0FvVVXvATlm9/cJQZkp/fnwOxLZUS6vlHYgyyL
1jJ1055k8jpRd3GsrpLUSUCfLvx79n7NMDr39UsNA5+600oUQjGMGcQcdwEHV1RN
wNhbjpk+octOq/O80J6YUBmJLBH8Dq9j4V/f2t7/dZ43mQ/PwKHBBx3Y/Ru1cEM8
H0+0wS8s9rP+EeC4ViKBfc5MDgWcPSf5YCrg1+LrNlq+6DPKr495M3kuDMXCecy3
X+D7wSaBukFoo2vDVdeeKad54PUVYVC6hkMS8E4wvSa5hDJ2tvSOPIjhzAReO8+B
M0CG+/XF2vIbty7tkxd3QmJZjZb0p6SIGTy7L3W+1CvtBzcLrbQcRUYGtbo+OJK3
SV6mI8JGZUqr7MkvSGDUNXo7rIl6YdTlW99bsuZHxpOAU41BVeZfFGuGjYB29tpt
O3l4xHGu+ptm64GCkxwSKnswktcFiURYk7aoCm9lqXQomDa3AxPTO0tiH8yJhlbw
zgvxecziZvaFFsqGaJ0Nvv+kN0ZnavMZZsQ/iujW37a5X3WBuPItfiK2y53NbiiK
UaRUvoifPge7WN8Sfv+Qc7c5nEJdP9xhMGpl4oUU1oEI3uG0hNX03knR/VbRJdYt
WiBS549z68yq7AnpiBbKZygBKOdZhwdSK6kD8j47VIKPhTA0HVYqz5oTzUSWHLvw
r1MMMVoiWnMUh0JVrv49jAEnSpyq2DDGTNPf4bsqMrDkDDjRHvg1G5JUU9XpsFA+
GB4sQyeG9QZBJiPpJPCoj2XyM1n7lg/m0mFLl4yZ33rZQSphkhMUgxFmzSBHTK5+
cWeFqo6ZgOyQoGSEk1/gtfvYhhO8I35z6DeeHxw/effcneBsmF8Q5EHFSyv7nyhk
8PU/I+dqjwlXPRTcPoUw5hNJeB53wH/9d4TS90IYYlpFa2929mUPFF2TGC5ZfjEm
hG0m85syKJkl7PB2XTbysZmUJ6TXLTcJg914Ulqohy78G6ieE9loUbf0KAMIUcWM
LKoBDUxmv/iWJU/fRC/sFyIXEBAbiuVHWSFgrkVLlksb1/bdXdR5GnSmPopC3s0/
uRpY2MP2LwyrIyyHT0fm53Yg9RsAIRS4+k5AIenpjZs1aPz/WwXoCgrFtnESFyOm
zeVjKkMmfpLlw6ytrIEGom3rZXOzRiV7LwUdlmnLmuiw/v/pzK2MVGZpna4lr4R4
S/OPhKEu8a43JnEjPh/0GYtkqpYOo/nZUhVMgHWpGqa/L/9ZsyI1uGCp/xSIqWj9
Ez5Bwi2xOWZlKH5qcqZh8MKwVvyum83LBCo1jZNqRKcc+Pz/2jy+cm/gm73IALXP
OadBMqqwdunzjqI4ggxCCvqagljbrVaIYIK8mptiuVujmAYmcURQfrkhSr4S2L58
UR21U+jFnkEDsGgdnYr+EkhDJF6gdPdNITbH4C+q47Y3e8h8mXzK6s1aBrTZfUto
kubRcsk0NqJsSqb1Gyop0ULe65Uob5vB6GZqpu/EF0AtcgiVpEBT8H3sxQTAbYL+
K7X974WgWdeiO/WHW+X01wQHzcSV8LeatIfFj065h+yJtBKgZFjI+UIPr3ngg1Sy
Omsux81NFR5Yb4fbwTuPnnhKMznXSVQsHT0zcO7Vmz66eT1gyVjNK5Qj6TlluNaj
tdgHzDYXXeiwFOEZgGbl3qaCA/3on2ACW3uXZge3IKvU2lJoJ/6qRFVKYSTEs4oc
fhT4P81LAL8IjjVta8yBApinWZlre1D++eGpSBkoIEaLj/Dhv+B+oVMZ78Nw3WLc
JXXofeY12R4EkHJgmVbUmNvUmow1gq65iBzbvrYAF+7m393dqGIYIQyz4Vegrlp9
uylsuCnwuVb1dK7frBAuodxb7/ra7qDc2y0KnwWT4guaYBUSOMOdAVXASAk9CzPt
2CXDa+S8ydlistOX849UsrXYSKUfL/js5yF9nsyOTFktawbRQeG5hGYq2PvCnb+9
ayeMUcgqOZYgjaZXYGRbIXLwENnQk1Q+fSLaEv1+9ICMX9GScCR12A+c1W0qltkM
9NPKeysoDHViLC0NZO5Ttx8iJBHI11c66jVuKm6ZhUH3mvD5ZvFoZjh/9Fx+kCm6
xNiW/1cQUuMT5FwfbBpSeFFftlnSD828ajAGeiCcRkaufvqRx+7KRutyrkrmnZvh
//o1cJxTNVVyh7ybw3g2HlmpnIEoWxmNP553yWV07b6Spsubm7ai637fNh/88a14
t6xN775GW4YLMtwvB1qYJPZti6xaRDTUUi7dSDln0yikcvL0rWjbQVdED1B8CYi2
qNsW14hQgWkU/MtQ8/jkKvesV539djrcBwCOZ/YlnY/eGc9AcHG7PuXEgqpLgDuc
CkreSqQalRtaNwKt0WGc5R5j5lS6aOQ/ztmc7UFlv71OnHRq3CJ/Yu96bkWvnsd2
H+aKu7P1qp6iE3471OfdhuQjrsAq/wT1hMxOTUUF7PhuNvTKlqpjvCew8ycowVuV
r66nFv+BKWa08ffIq8Ukx6DlZHyj5IJAE/bqIKt288pQtg+729Mb0u5gLgMIlqlc
4BlRXZHnrSUPjX1htZ5kSF7JmDTdFX5EBfmpBehimJ9yUvWebG46yQ1lOwcgGzgr
RWcxqe77P0Ylz1KOqOFovm8bOpdkhwzNKuqjKbtZQJFiTP0DrpMUC3V9BfcTBAMj
KdBbzbV/ST4+SjFONqmV/uC9BSJ5kVsd9EyB9C2EndM/E9CwCxcyl5v3fRjTQT9v
0Bg/wE3oOCyNHhiI7gOXipgCEU3p9BUZ0YGsFvGShknod9Pu6LQptwL7isIBXCng
Fjfc5cc5XtvzgB4MWyRls6J1AuCH4bH2cpkHYqEOMoaIz4tlNJirOkjYlWU8kLv/
1jFFOIyklQSo8AXZGIVaZUlbCvU5GAfGFQF6oux5KOxKJUY/gpEQc9pogG3ubFob
e9O0QzO7AX3LeS3P6OEXNdRt6NdLdYc+X3gK+NF0qRn9fj/K2u44tg7FPGZuhJQD
Tdl5yYVZutfFeb/BcbW1dHl0/IA5ej5Zn2OnpFUlegH3CPLIO5yTDvjn7isWDj4t
hUHpoUGsL9Cu3vDiTZQFI0BI41xQxTHJxu/fkSC6Z55v0g2xH7wI1CmvoiwBZ3We
CHc1A0sj14ttSWgOaNLpMfIRyrTgEeybk4fXmuBl544EdYgDo4coLRaTwkPNVUtJ
uQMr/aqS7th3yukrP8k/vH0CGbV3VLj+i0Hb4TEwbsDNDlzIGS/H0Lk0YAdwHKzJ
uGJoAv8KRliim2zLUOLGGc419JmFR8E07VHPnOtxPIr4rTjNC87pXvIRng+vcl/F
1CxxMVswzSRYKN299tECaLdhMZzVm/dFdbQOYrw124Uc4TYfuCTUEUC/miwlU+2J
8OioJC5ExTkLqqGC8kx+a1RS/UVh3R9RESceN0rF5N6COBvj0XBE7ZDRsOc1Ip3s
yW5MQSr2Z5ejR7bB/xdzRUK2p39CbS5EV0Revlqjp5U1Mi4b4mO37sgwpdrUjktY
muo31sD6vUZnFQdjl0Rd0dKAMSpsYnwnGeiaGUbeKIB9B7cPyBl1SdzXRml8fV9T
jWnWdVpPm/UhW+704XxbhaWxVewRViHvnfM4WcyeddQY+Af1iwTGIeLHv3bQQ6SK
CO5+y1Mnkj7VUYYqc5rU0OuYOwr30NlYAXLOGUe4/4LRN38HwXjK1sg5XhS9aORt
RmWcLPf92c6svuK1bi/yvD1Ynt9V2NlN7rZeIw5MaXJAKUgpEU5edWWFxgwEwstM
YsRE1Yolbz/ktJl7j4LeowTySPfqgCJ3148FfcPVYw3qqYckLAXiaYn12z/q/zDr
dHsKpUjjbvGLgS2KJc20PFPrpu6qe/ROs+oiyqPH7pUU4CHqheUIUL5C2H73vJhI
j2gYkWn/gFvTQkKq5LKbnjEjwEpF9ucOTGgSkGhM1Jb04rafrJiZjBibG2hnJ9Qj
5XNxc0mux12PXbCz26HEuUj5DislnvOaYA9HMwQSY9/55V1O9ZyNjitfQ72oiB/m
U0H4ljSVTkcYXmFGlfYJNEdCMk6rtKkNDBEBgRMg7zVu/WYIZbqUfpqyVm9fHAel
UFF01C3JOyMtAlF4uUcBN9PnYCDn2xD6GTFe3TCDqK7w4bwcXQsuVugKHb9J3Stc
m2YJ7REcIfKUe9y1SjU3yjPLLW/JvjkQtYx4sd7HWcRZncpaZNrQgxBrAS0pkOHT
+AA1pDUQzmvE4OBD74wM3zCkg0THdobci5R8+oKKBWAw3AMGZyGoJRKNoy6UTG2a
3rsapsrqWhJpx6Z2jE0n3TzZARdU/ZFuchBKmW7mDj7cwc/+uknHtqQaKBS/jKvy
w+Tankq1GrDt43jHvCKu1I8soQhO3k8kQK2DbbN4cGzqwz6mruPQ7wJQzMdyoMPs
3Pt51EWTGc4OT0pRUQKx7HUBhhb1wh2mVCsgD1YKG70LWgBggWhj8JWJezCnOX2C
4wIAgC8i8bVjlbtVjchlN+BHThj28jl5I/GeyaLlPyDtKh8SKlJxOjHlVJzRv4jy
TOZa2JQnAuq+SXiBTvB1v1ECCM9gcaIZ6Y7KJbhaiFyrSf76RohaH+uHeSliyyBZ
hqyz8mL9LFQhQVZiPiEXhHTPPnoX7CibK2quflTW4F6YkyxPNLoQy57RUtG+achH
7sQTvp0DObT6VYmFVKFubenJ+4S2krJwBn8GhLhX0DzMQFvh92oBf7gV4ndbOIGj
iV5QR4MjfJ4Nv4djlgjCAeWWVZcwmZc2xVSn1nHqZdPFqOj/6HtOXbOBc0q2ht00
VfH7YtT34i8MiLaRuH17pJYHTw/TkY/uVrJEPNnL1GcUffphBVf5C7T1rF0AJEWD
hwjubPDM7N0rFYlTmvqJ/HFjzonlalsAhY03i+hhjmivCowEhrat5PxbNNwQQI6z
c5WYhESzg4Lgo7CVNaCnQgcki+hPeUEdM4N0UGvPzzLMS+/ZaX9O90SrFOYn0yfS
UWjE3napt1YGea+kVj3klqdPSgBw5RO8ukTPXyCM0kJqgaip2pypNUB6vvFkjjJ9
d7uIzDKlQR+5UEtYMGZAXQP+HVEB9/w+8nKFAhfZFbjbUqUeaJm8ad0bEf6wbiJo
pUA5QdIN7tyTVhaBxqBtqq7+tsGkjNKEFRMt/0ldDXoe4StxMoYbBziDC/cBjytA
6SswRBlFIKjkZPZslK5v+YveCs2pEegFz5I79HZ4Be4rdtyMF9vLsfQnGta47vJd
kQ4sKbJ0sJ1dw1GjyMQ06V/UZdf7MX1brHTdGGM4zMJG86ClnCq8ZqQz8ycMWKuR
DzEK3LHI42qfAA4/ujOzgBku7l0geSS5jBKmvn+vb3S8Uf8vhE5j95+dgkA8ih26
XIk9xqHzzGAeT9sVI4mvRhGMyBymWPeui2e7hlsUgMCIW/J+lGbP1iuIhL/EvTuE
7TYftNBtvtdnqNa2sMG82wHLOd4vGSwS/1f2qYImMEtWozCcTuzKSERTmSG8/Yq5
p6uhiKgqx+x5rHiR7KDDrZz+2wgQmThOsYT1rR2nnL0DK2RFlYOn9s4Yv3RzIQm7
t8JfTK4aSrxQ4LjShPOxTk24HGVhTpW7feZ959Df9PHzvLd2C63SmeOefMM/OoMe
Qn2HDgEhwA0BMskNPITXwtst5B8yU1JluWWeU97rsqH2KmTZTzv0cqSqbZp425fb
b7ESZAO1EQIeaenU2NPwSddlKYYkPrx+/vSeTenNxLjc67Wioz+S7fedx9BogZzi
pjAeLgUva3qVClNOlahe2ODXcDxiehMsKbuZBqRpRqd7RbZnOGIX5Rk9SIGwSt8C
AUvyrmT3SnnhwUAuEFeJKwiCvUDx7+BHAI8NmMh9HPDtJLQKiDi5MebkTr/u2qB7
DQY7k1dtMnxNDmpRzBztEKNda7FqGumBKi9oTVCjthoOSCSPMp6zMX6ySyXYWSXn
NcbQAwO76HC4/cdN81rFqhtttBnRDk2r/TLqRhyKa0ImI9C4MsViDnhAazAo9E3l
0OLerwjIcFdenIZKkhFtuqvmbrKoLmJNMX0knfNuZtroxoRwznveiRXw6n5xhXGw
Ey+SFvby7gF8BD0sDe3LOBedTiCunG5U9xmrspOq2TktKCrNI9OIb/iO4BLJQTBZ
4e2YjQIPCAKltXk6C+nXwMVfkt3nfRSgCOwk/rL37HwpY/RF5K6yKb1awpcnEUji
VD7556dGDUR6mz15T3VeVWtHZ+u6/Mjz6J9HO0pq8zZG0N3Z8g91+XfztJoAZyEr
OjzJZhF0A0PdVhMkRXImjPjNlOP2888UrBc5ZvzMgab9b2uezL7jxRQNRCaLGXQc
2SChRNhEtkShjAj9d60FNBPawvEAXPSJZ99TQKikqe75PaKZQNuvoiVvPQUFTfhJ
Hr8BphTZfMKlboIvPHxBZeo7CqgKF0dinszjtx6rEr2xB7IncEVHe7j3kC1JDyJy
wigWHCNKyxsUL2OskpuSrQWR9KWZYRclOIAkm6BwszmR069UHkwijJnh29wiOqzH
jmWJJtW4m4yX+UiRjl8a4F7xQUC20LapdMvt7r8FkY12uf0bwJzQksbdIR1AwgZg
7xMwBNaXkDw6OaSIVVwfUjaplbUGlaMZY6m4mg54M4vYlFIIlwnZEnOFfYPj+abP
Kl5zcV8cSSQu9Y2kmgh1BmGG7SJpvxNZZ862RVwUgtYUUGvxwPKbmxd9R0aw8kaJ
nH1TmEVf9JgGpsFO00ZbX0l6DrYVod35mPy3OOGgjnCLlOVamH8qHEJFFg7FeViD
Q7t7Sai3UD23VyhLkdqhwoax7fLofB6l4Gnq5Tl74q7mLLgzo74DFgD2zZjuqBuP
+avsvB6XzGY3ZUaT5585qbDvZ/l/UoVLWIW48aB4H0BxEygP6xRi0FiuRo6I8jy2
qSEYBXGF5mAMqlpkB/gjHj3xwtc50i1sJ2c74VsVnmveE3FQZiroTdpDX/5DPQ7k
2CDxmvriYKuvB2UEd9S6St5HiOLbG1lBEuI2tM79EzB605VfctG2ysGmhOjubgkC
amCg61/92TJuTdQnV8zM7sOHpOL/5C/B5N884WkIulZCbuEjw7obAzkjES4jZge1
CD1UYf9wnjnvclbiCYS9N9hwjUW5H7x7EhK4WmFo62YGaGxRRjNSzmbS58Qwby07
2r5notC/Ct54tl1VE8IU5/SRAEgmoXnHCdjDCKXukU1G/DYIhWY1BRFjApHrRBT5
157dLJOFfWZGZxJErbNCCy/1wnZ6DdwRql1vAFZ6pjp0hz4FGu44znW6Msfthsij
FJpxfMfYy48kaoipGjwa0r9W8AX3d9HGIWTHfpHnHCWBazcmhVao6TisZWArWzwi
zy0Np75n8nzM6L/uRj3fFajEwGWG3RVk5KokPuKm91j1OPUMHePreLMYBOZSz7Vu
TSRJrfFppn6zf6SzxA5tU93ALcGAX8UtoPc1d3dP2/jEqx9VPbZA6qASAOw942Js
YRkkxGK+jKmbIvCISOZJKjM3X8rM4563IUvUIe5GPBEURcLnhuaNmLSOf98GkX7s
eYLZNejPMa/pdhPL7n/3XQWgpkfYzuzt5cVUwly14OcEYJS2MlXMmm81qSDcAdBx
o3uDr8iKHlZghKTyMVjcyHPHtY2mbsaGLRCkNhQqE2nvM2pCklgwahcVqMDJO5qT
rAZ7tbMnicWFpSMg2N4k4QJv/FD6hnOLnkv5e/8e/ROoC4prynn8UPByF+wGzmtt
F7E9iqZc2AAdLEb+TdCJiE0OX4p/oaz297SGztzJK4QS5MOMWL6VZeoai3idOqge
VRAHkg7B1RpYVtcMxd+NUSy3vNRSWYTx1CQm1dSakz9gM+MC/XZL1YyBLiVCdQH0
ZirURfF0Ry6nmc9PaXmyoa6M1DqExS+QExcPiGeVnyFe665FBXR+Wr8Mt4oj3Eu4
YUpH5VJyGuZsXU2/oV+wB0wyeS6sRdVf3ao5etyX/MbBpLPmx/gtzOO86hjocUPH
jF7ajvhvfuNKF8OMV1NcTdtcdolSxS+GCmAIGDGeiSE5ujEGlezFCuUGJuPV81IE
glQbssk+UiUcghC2SHUsnTsx7H+dThFWi76HFvlS+FMJK5i+Nk7lbSV1VrgKXyuO
5j5yfslcf1ELgCVHXrdUqInLKxKGazzJhvFujNGMFuRiO2SvVb4BPIghNxTapbw6
uGuuE4VsVexublbxCtgGP9PUH80XQP9qmcVh6jCcwbXY3CugwttpqZcf51Z2tIS3
CJFGB32W6C47aKPX0INHndNmFUT3XAl50SMICBWNXZj10/nwWaPCQZTFvDKv+cfj
vdMgY9kUXQfgmRubC5w29yg3NPU2xWS8SWAWuujmiovS8pBboo/DFLDmuiq2yjOZ
ZCo810g4OMeiKm2MCbgyuZZ8VC/KDdoX0GsBIlP9Jj9EXmLl48lUskXvXcYvUvNV
VAIK5V59ai0JfcMU/qEz5yx4jfqHWQNGsoJ151dAH1KsnfodRaCsh58M+XUu3VYv
9J1XUXACu9/TcSXXL7U7oFNs0G4Vb/HKLyui+uJ+9drzPs5GoRi1ovmG9jFyL5Z+
HEVATayruqYzEM2sn44SJV6hTQLWNdUnS9SWVM/AQxMYM8/OUBl0biUNnOrZjuRb
BSypk11giv3Gf1ttc2dEJPWXrkQt6lReWIaM8rgld/wTaRjvQr4T9Mlar7pV6wmd
+ZJW/MX98nytDR6j1hXobl+C27FzUsw15mBQ5rEd1mS8n7DC7+EJD1jySDCN7e0A
lprIWYIpTcg9B5S6w1QTujW/y6wVGYkILp9b2q7XIlgPsHm4QqW3ivXwGPTJnl+z
CROltsqB315wWC41eZBsDk/TYd7fQE3JkHHH61WFZi6Agk79zlJxSIuJzm6YuQxr
E3afcgMalHHIae0YQDmQYAhaeFlDOzOLy4Kbjn86c/+WPJcemIQkDY51SFgEVBcZ
q9orqQAF3EOSZT2N2lH0Ok1aU4raaOA/65GebcAeYt3Ewkf01XAduMoW60wthWxa
6RMr7bBBuJ7EOmLZ2e/dplxcPRzF1MbkDlJTkwmVNUgEEEn8OFkPUZyLwkxBL5wZ
+T61Yteu7R4N1i937Tj1QDDrRaF5UqgtMRnBrGO95e01cBWDM059ssMIXXiAMr+y
r00dzbxfFjHtzUmBzf1TdLBpwNfYM0i6W3+LnRn8NSYwCNwA+N1q2b1I6EfHN0V/
7ZstSLS73RPUWipBja+FliQEdKPsFTpz1z+Fv5e+UEdBQfb6PbA2TZqj7lepLl+X
zKMsRjeNMrvmLrn+9hoY1acn4Ybd/JQgpKq08Xx6MJgfWnnn4LJOk9bIcouglJjy
fJH60pUgb2EXEtXSWMf2mm8rfUm7Lrd0W+1I5EK0MDm8UzDmVXA8+8nUkUIzkNa5
DQ75X9AQxU3KaUOXVDmieQR+CRNpbivfX9pAW5gbIaaQ0aSU9s5ZiS3hcN4euOwj
hTx7DqsdKf5baUZB3ABSrJYtdXn9nFpe1ecUFI8qtxC9bJqlUC7FALdKlTZjwpGH
Lo/iaSXthhVxe1m7NsJHnHMbovuGtu1po4DLxbB9yFklOndJvDR6K63MiIGzEkXt
2tMiqzQVUCLAvTT1Tmj/3OVRE0qWPLAeKZV9fTLQ5mOyhYhS/sDBPGSIrtBmmnAu
qkCh/A9tmrdKp1epOESPHyFo7G8/RhVnBShbHTuWBsXw7O83GtVpNB6lnTyQYBs5
4skaiuZ4c9OpctM6xkTpxao22QTqwgsoOnuij9z/p72fL/cWL95NfVny1mamqZ03
wvkTx/qCIuJLXTEkksW0L4rZw6LmtUZsqFY2PeqdgGezoknuq0mMgfB3aK5kbvvu
A1kopQ10drr6eqN1cDNtfiIEnAJFZg+XQptLUMGeszV+r2vinozKLKZxh9Rnjg4s
4Hl5zz21LCJAwoG/+oLhfsbg42ZHTbznzSqMWDZ7vSGldK9M/6ye1jjIJtFEEXwL
LbgEz31IEv23gGKbA11t28Q+nwcvK5+nMtwy733kE3Zb89kvzFgYxFxxe0hO973E
fpERaoTuQY/mh98dA/nnE/TiU+hjvu9h2mKjTsOap2vh8N4wtQnWTY99hJD3YBs/
LueTLdnrbaFG6bVgqNysCMmoCq+e0WBiUM2njRDin6EFZdeIw1Wl5TBoCQavbk4f
qflSZjLJ43CphinE+EbAGwiQwCnb8gsAGb1LJogXxR+rPghzoS86f8knWuFF5orA
MpTWe4ZiG+cMBklenm9BAvqvRo+XkDzoDConSgto0kcrrrhRyvhavV4eoEC3kgiJ
Dn+dsI0FUYg1f3MEl+F/B9FlurJFqq0N1T8H6BqeIIIAhQ9LDMNksaM9gBtPjIvm
lZiMrwU74Lx2+adfPXLZmRsvxvJu/20fX4KXAvEcV3PIUlTziQFBh9f7AxSyisWR
QFQQbyml+7EzMWHi122lQ5aTtBlXtM7NO7UaN061RNLAlmwEqBB+0Ff2oxqVpzcp
ND8IahFuXRqzCYC86RCrlFdkwUA8JniO4HbnXPY3PI+10tgwE3v4rMBPAV+3Ys67
rv6BMvRanBlFtdRukU8yX7ptbeyPX1fPxC8PCJXyjgMtwCOgvzAQQYTwnSp9rvLQ
9Bh7s3QgvgU/K1xcceqqciw2SZmE8ju8YZDAxjYj2dRHVvPIiRFrzxkHBAY2Sy4Y
ONLQF4XZ3Kch1OTstX/EqFtp9aLY4p+LZ1UTjvl2j5/Q6+U4/eopysORek7AcHB+
KiJUAGFUeVBE0lR92GHeQHJulRQ/MG+tnCN0TM8V78+P7nHXnZU0FpQgzMszmHWw
W4cMYqqj6xE51MfPew1VjwlfRiiYZ/NmbnlsY1RZQzgBXUWLhm7J0TN4zB9Ez2eQ
ep36D3d3DctT7Z/spE8H64rY1H/Hmb5jtGWB6EipqvjTaRIZioAZQUGjx25dbpZ9
uGXMkiWQeURKxFR31r8+MtoD1QFVePmlXAobg8TCrThzOClQewgFtaM1sA0ag03+
FNh/jCg/xYttWGHQKEn2ePZF1RsCuW+oyta+gUpsT/PK9wb5e9XujyJSbx+mB55i
+9/orZXsCz2b+aD0647uX57EO3CeVAuUsMLj0KxDNisSA+JGxtY6zl6+Q/6S9mBc
bWH1TG+suVe91jrqYzTJKwC2sRm9tFktptr5k3DWLv4rrtnDhXTSSYmsAgHCKH96
bvnIII2c7DZ9nHjKas6eBc6e6i/3TYuGRfxIgWjn9zXupLkI8DZn1OKd1eYMB/hR
lQWfK0/LltufC7sr3XUcggJ1LUSKSS9cJ+EQsc3Iz+5FRlOsUcOqttV0H/x47igt
RNCYxhRGnYkKpNEcMjbzijCSfFY8/46xDX7Y5/dwU4rgYZ8grOoG+o+o3KtmraKd
pkn1gcQ0iSvUb/L70HmoAeqfW93x6vrT70d5rPq2XEoIJ1meCBRqDUmXI2x3z7+c
rk2htjrcF7+weFnGXthjHe14lkuN8ajyNGPwQ0lJ2j2N9lg/TZzCnbW9KUck6Mxq
G7rMn9BSWjb3o/+m8G6eCrwxvg0Wq9E5ClYRBBI5AearJOZLd3axP7hBwbg5I9/D
TuISV59I55VqHWsoMf9gIziVChYo/RloI1O/PGa5fi3NJ36fZ0JOKo5ErfKwIqUk
5X5jMsXwuklXdhH5B6fFEysIUPeIhasS2PMERtVZDkTAUdRmT8lkH3YSxWtw6M2S
AuDN9mmCvlXvBUJfjmqcoY10OuswL1UQoDV0Wt3yaGjlobvSQ4T0iLjAJeaIt05v
KhWSvUR261/5UfWtc7bXHXwAA0+bx2v0KDbhiirQTuBhZMYqAepRXwemnLcj3Ufc
hwuzfwjKYEyYroeCassYcM6iLh+YejTsvNz9OX+7f4EHdRlmw9nC8j5WD4Wo7MKw
r9i/2IUYS/iWrPRwytCPVMN6vVAbjKxwJp2I0jrTezwXp5AzMIzdzaXrd3UIwrUZ
qwAw8ObQRp6QACjNrWHAlOlBEvFVcjt2KEbJsUaq+AX4W5iPtWGMBF70hq0MyYTq
H6b9SkFHSz/Jm+RGCgSZ/KPTwlLLrJK7BsIQl6payWB7fL0ShPJfG18IDK0XlEPS
MVqq2r66nk930Fzgh9Mlr9SmHkL//KEsa90Z6GAf9sc/4hc9AWOkaAsRt/cRZZ34
pkvF9twoU8Qslc+QgRCJbvF1kDochqw8X5ygMzLj5Q73fTYQrZ6Ypa6ipk5UNqEe
IKXIOy02nDSbObxZ/xkuOM9G/7rpdtP9b+KdYp57/42fPuwnulS8t2KHS7JZpnyT
sNSxKvt8MZoikIdgohb1o4WmNUeybhI91Q1ZH4MNKhgSRAL1hvoHChcOxj9zc+2q
EUX4GY1UFq24Yck/tVu3D09+5Qs8ysUMtsHm0j3aLu48xjPAeK4t+GMvBhEdGas1
hI1cSNWOXDxPMpu0bTYNEV0UiHqOORDIcRDjXoInJMRfIkze6wmssM1xSmTVdJwn
UfCaIke4xREtntbPPUCTcB4yVRQ8QvFqu+uOSe4N6LvwtwSHxqD9mBi0Jaatt36d
VUPmgrS6IQ3xVozlu4RfO5GBHKGgeHzeCKR0bkjb0u6A37tmB0C9vHbW8zMaJSIv
fzxvgHRvX5u5JGIkgZcxlhG9ajLqJeOPe92q7NQrjAK4BRo/WcUk3s2NFT/7U3aG
8MAFKFbRKOgiy8pE828kKeXLaPHnyGEE+PyE31cerrJWM68ojZu4OKqVgaKqk+RI
QrBx9HqdSg9FxsBwgxziP0lALtjxUAYfjBYli8T5IFPBDKRmuKs8U4/5iZcY7YxG
w4YC+T5eih91RK8S43ZQFWuXLhB2tMzzKq+3/QpHKvk5DcTkrIjv+t1rCUFaykkp
oivfzSWSq5U+Pu+tclYq67W5jzgS5W+vl/M00HV5YSBseX/sgRXqQ08ZZmRj1NsO
5v46NyEI9iLer1r87Q+Lwm5vvxdqQhQJEiFTIU3uXiPC1XD3jj+LQ6bKB5J+zUw2
ScwUO4pbjSVrbOHBsthpgrqnRn+1h6pDg+jrpaXpzx+40LHTCsdfnT+MHHpzjiel
Pqxv/0bIaql97wnTd8N1f9UI4ONDycIYgCa0tUVQl92oYml4dH6R/7EeqoSUMi2x
Ew25KwHqte1GWABomvwvZiIefIEyNMPD0u2Nbtsi0Nm9iFMAX24wPJ/Cpaq2b2CH
VwLn3h7doAK6w+uQ9VGauoP1m1Ql2JG5KbY+w7wS7sVW6hAUBoIyerVI5jHCEgjU
wGTC3OKOwMa127EQf/a4u+utYZe0Fe0ZZIk7ErL0wa+eKTH0cFdceaIM5zVRJzwy
/MPVxW+/jTd1XrYv4mWXLT4fFtFjpxGgZdMOtaZpFash6mLZiUYW2o9qPAmVOdpD
drV85yyMGU4R/XfEyr4kpMUtRyyteUwijmOY1hVheePRrrDoS9W38/yflBjOglYD
ygFryBETs4mKS0RcwjIf83ybkURR+JB26fQ0syTYHMzJqbkS1puFtOidrglnOsSU
pKfWlEMKnh+ArzdMBFD50Sr00j1g+8zKj949MOpMf4Y32oUqApYAr5GJPaieYxEW
mvlLEYshaxIdQWEy74CA3y1dPUqZhjIuRvmbKYNXSutTvs+I7//A7wdVIb/TB0bk
sGyhvCZfnQCGwXuUzDTzwPZIi/TLg5wkji5fTjSTLlXkPSHdMc0+xtxIYrkGpd77
z0/dtTXct2H7ehtLEHDTArETfHCT/5QazjKWrHV/ZQjKktKJrc28zygrVH65pcRX
b3uPUkwUR+2wOavPX8e8xhu9Kz8ZlubPiUq79+KybYYX4ag2cTZdf3SHwLc5UhSm
8vH8suy383yF80SGTvXiH6ujYdgcagne58rqyrUxNGhyOioxzFTxWka0kdCix+Rj
7tr6Z9PW+zHzish0cxT0WfkZOutSVEpUzlsKCVdVGQp6en/yM1GLQRsi4cpkSMIi
je7lSkiBvzuXIQ8zMbY5nPeUfMqbAbN2llqfbHtDJkyNr1tqSHNJ+PusgC0mdSRL
FZDv+oI2frqXTikvM2AWahgflzT+VBj8hJxPjEEe/HclrDDT+y4kLTPEtHOz+HpN
7fL/T0EsNbv1hrIFNbg9s6JpyIyAcGBo0LAu/AdOXPI+8zsBcL5T41nm8U5zScH3
Zw3qtOcFz8AshjIzTmVmTYFitIjT0Jr1DW9+hg8VLUfaTGkKWJHqiPWD2bUXajq8
iQ+NPw8x5mhn0I9ymVLJYwRVLmPxFPuzslQ2c0Y9CoePthfFC5hNl5Ymjgee/k5E
tKAxTLGt8zQtybj/Ikh0Uysy7U51HWc69Jfoth4nC5uFjyq9tkraDCcSi6+HH3nr
nhlQLPBWFYEKE23WteTIQg2mj72+VsJB/gwd3DpriWpsgi83/yDxKrwuiShOk4f/
Tt5coYbVGNY3DLixYcNcED4FP2QBx2OOu1u6wt8KlW8N8qr4VKHCZU1Vipf2f7lv
K+ST+Ltr0WfdpHtknDtuL+l/faWkI/ptI720C9Y46YChA184p1MMt/acoRJ8fdRr
qB6TnRsavFT86ZjXGa2PcubXucPAkdcN4ArylbuEKcFRc4L3hl9YV9o+oxVMqiI6
gMaH3lLzYNYXv0En+d/XYgAgaMtyGP/XAAvyptQlYth5aEqYbkbsuPU5mgFNs7VH
pJgAb06EBZmBEz7P3jzTC+p9XgLrO4ni8KwMSpgcPbvYz4wLJpV2NtR+2zpRfqy2
KRuJpM5FPO1HNVRWTRhKK2lraxjI1pngawMkxoDQNFVNsOy1ytvRz7gPWWzmMM3B
5BBOAvzAQfH1G4AF37AAMc7EYXCTMGoiJIMRfMogVahNta8DFodvTdXSbGxKZs9e
c4XwkYdam01u/nPET6ySGgzovjvTOuPFmK09tPxQliRokmEAUp2uH117CHXKejaL
WWiOwVu83ZT2+aKokZ9Vi286cyvyMr3g5AUIB3CwgYrKi6GrRJ+2ZBXM5nBEKFJ+
99+GT3mrM5N56T6V2Z4yympotZbSBwocyPXER9bVga0kMdy2QZvX0db8LbzrbBQW
RJWj/ZTqBFkl+0nbvuUFhuQs9RL94svfP9pKwIQeg+7FN5NbPcTTXLCi8+44OWDL
IZfrsqnVxf2EX25n/qiEVawzVyZLA+1HpLaASDGui5xsWMCMuBRZ7HnAm9vOO/Kt
d0UlATvI3b0xpe1Yxq4YY1MlCaXryTfB/fnCsVtaNgkLCi6M5GImTWQmfQ7Fjf9P
GDZ3XqVKbvdv/pRDjOXE2W9tBexKscVuhj1DN1lnmBQc8MPoUnqky2LWiCcyiq6a
Qcx+dzWe3c7NKXWwitKyrnmMaQgoYhcpI/YVDMmiiinZesULbuUb80gM72K+u/vd
5tP1JiGwYjq62B/TYgha/Gh2BOF50VG+sl8uBQYcaUFxdSS4hZn1vSzDXkIjJYnn
aAuiUP093TwILw4FsL2BOM4TNn+sX1/MWmWVBrAzncZXaDItig4PNo2W3/jrONzw
FHIXW3nx3YJapJF1bJ3b+NjhWllPVTXHrs/X3C3NmJw19x7OCHyw4E8KQAxFWrk8
T9pGrTT/10pgR8s46BKUHm/qmOIbMhwPqP+h7AlRG4Zd5IW/ik/sZ2xJSLmnKDlV
mivtLL1iKLS628uBiHLn4/zoec/bn95lkCLCpP11L8cFZthH+7UaszeEgXaZ+lXp
KxxKqeMbW5biaUPB7b5VVfL/Dyigwonix9y/nOEsmJHvOtER1LWC2RMdGNHytpit
jSYjKT6rPxirJgKsIrzAXphgYa2bFHdBFDqlGxT6yIxH7MgZYiYiIbyQer1u1c9E
kn4Dr2pP9mIJj8hebi7GTwWHpszi00/bbU/fhRtw9jznRnyGfHiupqUNXaHN/RIC
jUifPet3t6MwxG90Mx45eTFu7pyTj1hbcd5vU7sWn3ag3AYiRC7hlHzY4R97THcz
013yqBas6hboazzW7yBdW0iGNFLnSxsBUGiOBPCAt9y6xYAPiNzuNRVKlk37u0UA
aNwOlfMqmBvL6hE5iUVo1/xGYGrd8w/1XMVJFwLwl6l0sFmJcjR2DHLHgw3mHeK2
ICDagY268jXOBV1NFqaGE08pSjxm3Pl1bP8lqXktNJPVV/vwNJdgKNOojtLv9fFF
a889oU7RZRe4jgpwnA/zcLP4ehaW9isT3BEmLgjS3tbhY7I3FYD9aBADaBPawQnY
/d+VENM41AEmjwubwE8Q8HQ1ZYkOKcfdYCw19jj4ex5H8YMv5WzxBzq34E/1+ioU
ImJZtEx31xvjWz74meE4kymX898LS82eUpEpI5DQXivcg56pO+9w7xEBz7qVWC2J
R4ADgASlQUMFHcyzAjSSodubs/szHqyUKr2sOE36nBDhtmsgHkQqyR9PHzEsjCxq
Qih/H7HZPGR0LhgsxRCdzt2R11CN0SPXe4GWLmFQDejLCY1dRA1O7zxPIU6POVxx
cUF810fjBi/3DUExzggHW+CyuIh4zfzOGxh5sNdQV6FLRYXXZlroSyeRxK6eEeOc
l72ldY3ZGhumZKUQYnvR76AGUwIvO2LPW31wAeiGK3sZbjEuHvqeCCszMw2eBGyB
0Lk9ub7PF62tx76E7Zyk3HET8xbQZctYZdJTuf1qepK45H5Cg6B7VwAd8KOz4EZk
NYaJ47gHzMs12iaao/63T8Dbgsz27pEEsPCndghyM77MKEc8q5NTPPW/wffj/Qmw
ybuOZqQNBRfBtzEG18ltAvHOCQcgVrTzhlj24FUHIsAFTVCfz7GW1A3vGDBE+9yv
01iGjSMMJIXYyo82skPCjJ/yZuFCeD+HIAh1+EkiGsnbpaJ6DFOM2FmNaZ1F4+F5
arjPDh9apwstSDT/rN6QEBCxdAd45SmkYz/KtDTeUrI1ZlkTBHuhvM2SmPPVi/kn
rU6W729kYhm5DfVdNIIfJQBjBn6F9jwA0+H/1iAfOh2e9jOewevqk/aXWtbmFmZM
eF7AaRHeoNYRqxg+T5l40Aw/edIwme1oVr0vvJmPH3UFK1poBtqD6RAojT73WNvC
HiVXrHOnusFUfwqRNNNz/O5ka0/W1rGlkMNIqDGLtfVW4DznuaA1ajrKWZ490BRi
fWziAswO9Ug30nG6BFK3X2KOng27zWuLbg5+VNaZ8cc4f93x2mKM5/ftbkG+5w7f
ze6oukEnAQRJPK10aQaa1Ns1B/tvWvngaU6JIOgifl5J8d5eqV4DmAmTiiFC3Q0E
XBZNVpswhItihopj6yDEtRrZHc0kMSiY9Fo2J+m+tUYFVi38pJ1J80Tr3cByybwR
p497lxHkoVrld0NI4G9XFpEFqT523XqAtWmA5XGeU7Q3xVEL7cWAAEa18mAzOHdu
ZFbj3x4E7X7TFjYFqn9XSWqmdwHxOUStSqGPMwxURXTtdFpnrHqaZzWLxVTRKXoc
ygW42OfodoZ4Jc4Ds4WwgGNUteCkoB6CGZqyrR85GnsTxsmN9h0qTnTl/WyNpijh
Won/HORi07Qj1lSJtFcRIwpMT5TsYeGvA++Us//voiYsEnS13PKkXhaoP+syxgIq
+s/mvBdbF0yFN/jyPkMbPHpHHB038tSYPCfi5yOBGrEsHbAOpN36cEDt50H1u2Tm
svpG7wa6cNBLFhat6bGeXrxDBUBmXrYMU7HBWuXoxkUNsyms+ZsAKdE1sfh2GaoJ
wBs56xEhxr0qAnMko20pNWSaG5CvWGrr3G6pE4BK/DGfe8cUb23WFCQOQEH6i2hX
3Dl19gqfl0iWY8iIotUtOKneXwtC6muNFQP8DPr+eCfVQ4Y16OsaIHauPlWwwuZi
8xjil/XKcxtt4nG93oEhpchIONO6gYcokqeFpB9eWkqIOk7keNL5F/ugz773D3n+
4KFM62UwtOs++F6oQrwlDyBUpd0VjvhXBC58KxaPEyT3ksec5zSc/KcwY4ysWBug
aENTjTXW5F3OKR0mIboQ29hFHtTRaQtXVqWHx8jI3msDbPuF9s+mlno+gv5oEXcC
jT9JND4pVFIhK/YtJlXGA51vBQ0ITQwNdcwlJCj4ap3c6knCSPRXB/2cqOsxG+38
AxMPApeyZuANP8e9FLpdyTsr8H/Q/OFCcsD3PUsG9liR6O8t1YrVX/b/f+rBunUJ
4Yta0I2rQptMdWzmS7SbGBPQRvZS5vg69NU6Zqt62fQEiou+ESJFV2DghrQQAZo/
apSARfyGByTM+tNGyEZmBW54YVk0eRKiWBcvgHlkdmKEHp5XF6ZcNOc1R80cpZ0O
PfV4c2MraPDFicklWZZI/voIesIrUEfuvfLGYHSVyx7T9U6n+DTm/m4yoIsYgc2c
m5iqycvHkoxK84Cy8k2mFegudOosFO8o9lldfBssekGgi2DDagkK7678oUsPy3Fp
+AZPQ485YhRMMLGUR01Zsrp4WdxX7sSMRHwua6ROWYWMu8Uif+A56VkId/6kexAI
6+IM8xx3ftUf9Zzbrkr52x/DVjI2BK71z9wvoprSE9ihaiS42euclc9nx2tOGZOE
0mm9neOCHIcmuYRxPqSzt+odheXVRadg2ZTINhsGALAoCebs6kCpO+UUIYpzCPwh
2CSG/fBfDm3zvIIzRr+6DIcoftwO3RgxrTwjg91kkCuP2cI451QeWPmZHQReYyIA
Jgf0xjvhOUOk1UU4HveEjahrEcTVOBIGIZldiFtsCPTSbIhjJrf4v0xQVnncgXE5
deYbnIk/P5nisV9eKvS5ku0ab4/R7oby74ynBnuFZfzDakyHqLn669qVc7J6QTwa
W8fIklgAJM0s31tkLFeqSk4OUoTl2Ku/4ra0GeNLL+X2mDWavhQtl/sqcpCDUTZL
AcF+c/LLODOhxlHHOh2EPq7mxRBXW6GM0HTRr9O1Ff4YcqKoQ8kC7wyWX+vAgBaR
SUZNBbkhlPZmQMEGaSQzZJ/2alDwmjzU0SCFlNDcn2bIdQU7/tKlZyXR7ogk1Nwg
L6XY0FqZgYlKYtK9GXPwirJb4n1MmPYULeTIgChDtxpwMb9QPUlSZWCwY3nsFeI6
8ZqgFzOrWGu8noc55tr7WUxAkEo9UnKNer6ftyMPsVzrhSqnp5W7i/0qNlsGxTJt
sAJoh5Are8Nj2mlSvXQobnuGzloBCT317wuFA+8t+KHSUF/VTnb4F+GmhnVcZfRl
SZ/a5iPQxFbRs3iwZK+MKqASdzUoKk4zFXnV8yIHgjuaUGuQndftZu1s3WXrs7PR
hLgwcCZGjYkHZpJs79OQzRpavoaG50XycDEkbbWDhKqpOpAn46EctzVzRlDobgJb
x9nddDyfadnm564LUHzmdaORRPH/Q7RKl2oBsRFRB/vuKGd2Ms7hcPONcsipOiUs
jId2Z0J5slQn/8IL0nRinaSt3Z6cST9dBu1y+urVhK2zOk4DZmR6Y+ne5OR42paK
96fblj4xaRXgDZgZtQVe9UIyZmGGPBdBnNQJU0X2XlDAyCpN/+61dWnv3gCOXWxx
jnT3slfD08NBE++QEcgqGh+/bh7ZuVJ7zSOV5YQKSbTsdk+Nxl5eaQDFtjiOUmir
b2GUYaKRS9g5pX2l9yy2IYx6pdb1thTOwDpfPfIT7F07A15XBeQsxqSQtHE1oOSE
kT3AYuowPROrIfamYz5NO3JCUIwltw6/mAPXyjEvwgzF10n1cbUgTtrz57eoxauC
rqhXp2mfGJ2w2ebvtXjscJ3gR20h1W95PykdBBlmBofm89uw9WGoucwazkiclbWJ
fMnUdegcATvPC3iCMBC1Tkd2h8jdHg0Uj9yMNP2rgK1Lt6AmsW8w1RLiVnFr5+bj
0KqQqMzvyGbdT67XT0chCZw3GK5AGjsODrT5KcErAKIhcofG0hCIa+m7aiHh4f4o
jLMHL0JXUa4SnWO6/Ik730bKx5T4lFN0d9hjBYMSoiQnnTUNfQB4i53nq/Qghw3n
NCs4GMb1OtZ+E3lF3QFxMqRHk2vdgr8KWd6lt+fZ2cadU9B3UYFop/9ej1HXz9IG
2wlefBfdMFAbEYEvr3MTBQ5AT/5WfyAch+9npmDW1H8dwnmR78QeJUmuRwPee90M
TkJxb7k5CFyBGEXjym/I9JMI2c5q6Cai9VwO6262410Qyq5FcmBLvJVUt6xYtkB0
xcT5ucs17vRRCjXGfiLMG4qAuABpthUw21uDGtyP7m+UAXq+0hKbzJHyX/hrBJN6
WVR3GYoNcsjeZFDHRg06P1904U76q09HkrWa2pyu7kf1pzKjS/3Db+xDkLH/XpIY
BbPdZW9sS+qkBjEn/x2hwkTlTnzbvXrur50gvvbMqPlFHOOtuuC22UrlNq6sB3at
+RNoMzmG88mZ5euKM0JlTueT6SIVxwBu6GrsKZjuee5olnsDYtjJMu5KE+K8yQOW
Dzcr4rZBaLrRhmLz+toHk4ipB4bDKzXTm8jAv53OdVNQJhcG+ANReSHZYnuLJc80
fktL2FuMi+S77xvn5q8upOJsrREUEfVdC0Vrbv35kPyC+SqCV1WrhOUWG1VAQQLF
rnn6paEs3buMrnFUZuBM4OxW+P3Cxmjp23I2IB6jHwhNd8/Mt0lI69nyGr4e/GMe
jxuC0OmFkb8vlDJV5yAYO/z/CMt4v7LMf1ZATWo427tRQAV4tXu1JoSHSs3Au5dp
YsrnRYm5NvAOZvoLPRL9rVliwftFETRLfic7V99V4Y59Em0uTmSTuUZqOSaZPPb+
NRRhJoDEy/F1cGarAuhKAcwupMFP1M37DfpJ7D0vHaH5b5TVQ9V+aVHitWYNixkj
oQyKOnXG3vzFaLZXd7rg2mTk6tIyxbpBAYGNcxgLs9I890YzZ/jvjLqG9Nwv+xXc
l6b5StuEp8CrrzRy2m/tYgU94A9IqYsphQpkZ/f3vYLDrBQ0dkXE/yxlHI9ZEMSq
e95o3T5mr8wEWAUvoXBNGQTtANSvT56KiJCwbBLYj4EIz0AF1H7/W2UrMgBcjLq6
f1k/D7tudS4ZKAiOBTbIDSdxIJgrNc4JW4kAzZ07QLsKX2ocmhjESPCUkIL+Et7O
nD+kpez/MuZ8g5kRy+iGUJMIpjlxZiHQVZtO3Yu4EK5gfFMwnI+AqkE+G0i49mcS
yL65FLSbZiliPGDjseTAFVq0hYk64jGlU0e9yT9AwlFv0sb4ywGDBeRQBAOw7Xn5
P0dD7OyIjDwuGcaQ8PZKevunLbHzjjWRw9vgqzZ82zv+zwras/ejrrT6NMRZKelY
L9VZt/lybSmG93i++85TNr1bDdFp5zxzu58f11xlX/C4Be2neTgL7aqBrkPvM8LS
iv5NN4XHub2rGiDNJlOzEhLw6AZPxHAgBEge3KAlSkL4MGv5DPeYOgsJuq0DGDAx
vYjCm89aGAx+uT161EYcPEtmJ9ike0sUaaUDAFLVm5HOg/CsY86POgu4gGhczm30
nXqUtNf3XPu/LhG9J4eotrDyEPskKPxh9ijSrSnSi7uSpZJFvW66OfHVLptrGn1P
1mWreazXg6X/AXhCu9L70FzttLqRpEdzdn28GNwYlWh6TPGWAmVh8KwiRiYDv2iy
CNne/l1CYvFscqeJDViaJmhR1txoEoV3ZwS/HaNdyx6lFr9dmOOHzHRNklQB8X1q
QCXbGDKkKP9CDqonZ5U6qSDznwFG1dg7qRsdaPgIt8VJ1tfpjAqf25pyMK+V/ddi
MSKHi2W65dErGAQqpRmvEQqJNL4mNlZh5ATNBAaMvy/MShrhAxwjOTT6PtpTCNKH
SWLStBmmGDLmAg84lZGehbYV3p4e4LFOAG1St8bhT0giHhi6++Ti/0ACYUDImo2V
fVSw1RnJYJ1H/Gwc/dPjpVU+ocYFlCK0jLqHYTxeVBYYTkpOkj5HUYGTeo0s86e5
4HOVLhwskCHxL8LhKSOIDuHmnUIiTHT9VnLcBApayiKoZlwjes1o8dPyDYWvH73/
aBl2YinIjfeML4WEltfAJmOFBY+k72WSAfHUos6qHjzbewfQDhkAAk/20MUc/Auk
4LvU8uGgJVY4FWKvwmerbPUmTtwwAFGzOMKUuJP1Zrnd/TX+3iuqdz7nD7sW+S/+
a+uFMJPybtUFOmqnf2M0QWYEiBehaKCHZMuq042+5KwWagcb7Q75Rx4OiiynJkQ0
SdouwM3HFJ6EPmciGNiUrcLP5oT8+Fnh/6ppObd/9DI2cieFwMdqI7CUFJfdwTxZ
B8mEkheSQvQ9dTl3+j2RfYZj2DI2SQ+JNr1ColXeYGX9UbrePrKs4SHOkeVlxTvS
A6nw7PVyGocK+h/pT+BmGRTeOsFRhnCtmFQTSnr29rpySwzFPK6gNMW2i2W06cwa
e7gOWCZmQzrK4GOMIdBI7b+FBEWYZ4Oia3PvVqoRaM6R2DNYoKfwDodLUTWHVJTJ
YVhIHZ1E48TOlPD7aaa7Tp9VGYqEe9JJeR5ZP7Ulj68T2cnd90EGJKweU+HphUr/
r3Bnzd5ePXYJlIadx55LboOAZJdPYYuUProoAiI/pDfA/6tQALEyxYLc/0tQ4CWT
T+/0g7vrW7/HbQ6XECJpEqZlWpy5Dt6bUN6pFX93mXdiTw+XydYAqNrFV/K/VPcm
/ViNpjZel6H/xBECEndp2pbLI89nZ6xFJG9msnWR8oBEMiQrHQuZdB20BId67KgO
847gztDzbj6wYlfcRDfuJeTcRz8qMbq8Z84epoq9KlNw7RhsNYUoldncZE1bKF2n
OtaRljwIA30tx8Xua9xl8Ulz+z+7jRA1onXUViCWCoUZhDXyDbc2VGuPx1iRvKBr
xIopU7sQOFEEkID3UnyGug/GFRoJSl8jxaOi/P4PCCCs4kY/L4HTUm71sj1qBYVm
HfCTwJZmlRiJkghKbAp5j9NHDTwB0mAmfkMkWGD257n4E2SSWUKlFzOS0sB96G03
4TYMc1HliO4yGnW1/h/BhN4nrJPsblsX1vmaVyqz4VkFp6uH57j2IiMIiP1z/RiT
Ubk3RFUiGmEMN+4z1Wu5vAD+LoiAFGVK9QqItDZA6C/RBs+hajV2abIVbkf/uVoe
Hgw2SAvVR1ZaWVCBSBV6oIfwwsOnp4cbfzLzV2R9GFoFXta+T/gJMWfqFBPFkgaB
W+uwyiNMRZTLtmAD5CpewPPYe/N/wK/OPsihval4FtZL4Aik8Oed7u9IE3T1k0/0
TlhL+VMc6VrrHX2mpwrjEVi2lHOz5XOsbIHb9mkXwJ0t4fCkgKn/E33rBtctmlsp
aeorVppsSNWgyO7yFB9ONf/6mRSIQF3myXW451+PfCXe+u/zWts06OnM7kWoWxmh
0xe16gJBaxrnzfqnLFS9I+5arScGDpz2Yp+6kMPhcRBFwGAmtUs4nYInuwasozRm
F5tCORFt869U9sRJG5vQwHRsN1gP4JFLogdSdNnUKLGQgu/arU3UcpW1em9TnZpW
6UtNHZVZ9bJoYTTRHFVs24kP0eY2PezMLSD5Ff5GvkbtJrHCcstbX+vJb4EmR/JH
CxjdEYmzVu71R5xMXm4FFGfV6htgBOWZLDlaJYFntSlK0OKAckFI8kjaIMfAnT4r
nFbVqWmjBticpSE9Mi57O0+FT+vCeCiLg1cZTFpQKQBaUX4r8T+u5/AJiS8W8BKx
+6hyw/U9MN/kmz9e3izB7s/skt736tBR0KKT56zMU3z/pcryVXcxBZdzQvSa1iUo
tZn7Me45NiaYAoDySWJ/SJlS2mPdlhXFbhUiKh4JujHNBnS/jTOUvRHu3v9fFQkT
TKog0V6CaDTLbGmGc9ESzN8Evm6wr4zvxnsPRuB368m0blS7FOAOCDmWFUwxhiin
UNpT5BONhy8YGqiMJrcRohXYKZCVrrB+lFVzRpyJ4WU0SKV4/3DAoKCp/0XAC9xz
p4K/DDfNdW5cnd8X9jrS2VWpv0ZeuAAwbd3HCq4tc3tSM9Hh4BnH0lGJye2VBDw/
+TZBX1CIR4s1/XIngv6ZVODbVzeP2AcBOuCyvYp2GfuT++KFC3t4KXQEWvCWZs5v
AdGSGcSG34Tj74GVAoRyOhnra1ywO9fhGA5Rgxhuj+4z/g3PWm/uZaTU5/xPIDQ4
IKOCYordUaFfb3yIUvJoyM8brdq7yXe6LN37nUNCtlGGj4Vz9jLObxo59s7JFq8U
qIwO+qK9OKuYBfIT/3fg1JSDMQ646Szj6KPYSOk/4Qnfj+UoOFwLUVXY6Xt1EyY9
FtvxMLrBTS2POzqGS0+8nIWawADHSwT0l0xVwgFR/OFiQ6rvvYwNEUorbI/oFvuy
fPWszWyZxehCeZANGA78/7VqUpQht3Me2nLIHVrt/Fsw5bUJiCd9az3X6R0CfNJG
JQQ1zTYjL1wu+L/JQNbWToXf2ZTjsJcNAvWm/G47J6NXI27MQn/wdgMf0CyFuDh1
vQs0P+mMVpBGvLVubnZabM4lgdKmr2YyxirW+UeABSvP8Fr2KobowTlIi/J9OYIu
iMUNg7c+2AMftMmMCg6S+wjC74EBN1ZxHsZN0EHlTkMK1aDCZ7z+dpxCqV5bvpiw
d+jz8qDAch7LeKJ5z4JPrRlYAQmIvZ+UJUbW3inR8bBM8Ltf1E1ScuElkb2yLLgW
b+eVXCNPVxKG2KKa4k+fV5CF/ytTsO0HSIRHTA7KgUP226z4Fattem4p9DWlgY3B
LNlIHIj8muiEc9cEJQSah3U7NBBq+0XxLJdcBfvYrmIwFO9BeCYbx4qLHYOLeTxh
rFkqbgGuaZFzOILkXBqNMovK6t7KqSYK/ktsO9TNyl8kDz95+tXpFHxASHaFN9S7
IGiPdsZ/aHV5DavlbdXLMeHg4FHZ3CahRgTBYMEHtzZ6aYVQ7e1K9bP+7OYnyttL
RDv7oqUaHJuxR5keNXyzjQ1eJrtsbbrTiHFLK3rT3QIUmHqvAh5b8rdSy4U6Z1ML
USJ+8FxOpyIESoCQWRkyWS9JjpN/mbogMjFhRKnCij/dzP52EaFEpbbCWbG/FaXW
WFxEBNp48lD6aF5jlv2NNqxxDURT8hILKHDs9+Uo+5W3e9G+1pCnsw4Vbd8mr+xA
jLCsOM0Gd1Sk00BgMYYy3LTX0OUQOAYzfD4AZB1NP2JvMJZLZ2vnHi15FmrkpoyS
PRUp2tbujwcK1xFDyy36yFV7jk6JjEbcNvTEpnUL3DeLZG1aNihu82nZh1TE07oj
HXv+X6Qs45LAcXgqU4E/vqW2Za7g/8Ivs605spFnnHYAal7Czkckg2xreS2FXO0w
+3TMnXX/ot428iZabdqbcunLeB7ojAkgegqj4uM/CwDYdgL47Lu7FMPT0TXXaiy3
ah0FyJiAT0Axz9v/gZjSDm56BXSlPJGrM2RX1To14Hp11/lzNny6G/0VD3o2jRS9
hegSFM6Yyx2mX9S+Ds6k+QwG1TPPHgoci3UsBhBt4ToPwRdlYeozxwynrAM7Kgmt
OV9ZWIMvY1zww7igMOANpk3StfiJVXhRVN0VFF47Lyf9zR+wa9JYSTy6Ol/CbaNA
DQgu4HnacvxaLfVIY6qn4wI2zcKY4DsmnaLP6i5krZaT+SMDR/MQxTM/itO8nDgb
fgpXVDG2XB4aRJYZ0Gy/gTKUXQXVB6GBdWNoNhX5B+OUePgGEvsGyTqy2cwqOHKR
55PQ+M+QUGW4w9zKfE0kWLLrzPQ+jHrguJyqtKeMLv/1JT1QuFuatCLd/AmqhUmP
hL5JICs9nboKRZcfwmVzNGJOwrri1Q/ykVbQ1qYS/gCFX74XGUzh7pO1Csg0L/sy
UCdtFZ9+jDjXuNyFg+vJkq0O2aok1ufxRL4Qw+++cVWP5KFVMkI+xl78MJq+Suwo
65VCJI0UsheQWz95ArFqyj/iIA1/lzOMd4uuzeGR0Z1grAqfkXeuHX8P3UEMD4Ke
RxbAxsLgrbfBYJ+mnbBZEkvelm5huIKrMxKSzZzIcj5kItfXYDGZsCWbCw99TfgT
7RUzoPy1/nFaNqGaVmo/G9Jew3wg9NFBW7LFYvPz6vlKALLVGtCz2Lw6ujfQRwF0
/2WgBWMqGZBBqcpePaDMfK0kjxsKuDFHAetiqbcYtHlekZ+awyU4RrROfLwlMSHq
HVdyJuOf54yJ9LxA2TN644GlLnYL2HZ0HpsFsswscXonzVX63FlGeejFjGZQ1F6V
eES84nmnD/1Pai0NaoeD6dwSu5WKnRIdBDB0KJ1IyFE+icxKLvLQwdqBs7xDG6rR
AEeYVjMgHjhV5MB58h5bVapXRZ4wXANSrGUlbdmiG5ooitxWr58cozKV8awuJV8S
rfuE/P5uqmU2pnc4OMuAGTeJWE2B1maZAxcfJKvLKogmY5oN8YubEqr6tkH6OfU0
Y/Vxi+4AhIIhluQijp0HGIyeeR0AIIVGla6QpGRge8B5wGtF+zaB8xWZHKtg4O+0
kE12SQQdJzyN9UKTRVonflQXahuAPl7CLlCjIXjJAr1zcyt18cAk3KIgHK5JZ4nF
IbSwanuN/vntWAaqtZJ8oihXEKRXCevBl5q9lZXycSyetJsGpCFjeqcNQ05VxQog
zh2rJp2NRIAa5h1wNBvxuTt10k9/xqWqilrpHecXjNTePVP/yWgiywcJ8gOPs8D+
bc7DfEnkFSg8U+CE4rPTNo1k5ZH5HXVXyDTmUsiL69hOj/EDyqrm0UUCwS26Mifu
oM8hMzsnU10yslE0wzhNcFhk8257xuj8YsQmKTDnya4GLzOcAxxk5E230Du7legn
5lWtLNVMvz19udGp9k+WJUFRlpFbt97GrkRmXZx31VmTzPix4scoCx3R0ThHQufZ
X4XRwQCwR3yyqBsE6FWbP5JFXIRjhPhPFro0pFYi94LmSvsd+cFza0cmouRNRT2x
7tx27+lyud1WOcH3DZL2Kob2xF8B406W36vXkjmYfPJ4tmJqg/fh9cIIQx+EfQ/I
T+bq5rSB9vnUJ05CLVawfQxSvBzLuIAg0Rx7oFx63l7ejjmtJbn96PZjyKMhgJTy
SlxXEEqBYLOfiXLDXqpdxTbgscTJ7/fDEXHvjFTAoXoEryYZtY+qBt0bRqWcspbc
B0t+GtGp3ve/jllojRSuqtrb2jdWr7mwjO9eMoJJr/v5nNGIxEXFb8t5uGvVTbT0
OxrbCdtoW/x3iA4HK8dFl64unJa3ojn3YJIVQ2+fUOTOWKmdp9BD1XLsi3qfpCcO
OrOMC3v//hu/jQa1g/StvQsGEQSphyqjOBW/5MpdpqZz1SBCLxjjgoCqJjgr4H3+
n3OIzRB7xbRDuFY1Koh56UlTnFubfxiiYBKjNPikiP8MbG+OEBuOcdXYzv/NyPc+
+Yd/0fPOMppfFncLDOEdznqh2Kj7jwg/wGdgKOdd5RzBlh+lixR6m3ydoxZm6JcK
QUb2DDvwvT1vwelOjrZeZ/Q8M5wjtSiQTaZLAw1+E3p4amKeHZLG4IvsIT8m7WSD
iNIHnYH2iOm8ypmW4YkEx9rAs31Ir46dzs+yoHzst/uNM/JmCrmAysvLieBc8sPd
qBIBglQldQqDQFC/QzNvxujHQ5clqkUqNsq5q1sD7wY5q/e9ELRtpOibGPrnidbo
S1S+8CJC++AIDOXJ1fHdZPVG2U86P1oXEP8XBmxL2E7MDyyrz1JQJgbQRi04h2zJ
anZihRXnt3maYeo+2EzusA+MAEMAUVidymjoOci1FTf/5CTJDBN9CJb/FldFYRAZ
HCACAaNI4Sur/q5jEeF1z0iC+N1ZsXTIi7UwB2rjaBrnFu/uAezbQe6wshbA7oZA
dizFnggFTf+HZ5vPlZ5Mv3RB2xNKCH6KkzDC1mJdw10yOT9sbgxQ5BmpjvidCF8o
JhQbi/ew8pxWqnEeVMBvkT/liwOstByC0iIFpZCOgyY59ANlksSCPcGJpbUf1aVe
4Q+D3Itekoqpx47Jv1MehrigzktJCJcU16bnUL0SVt4JXO6WwTTTc7+eXdUolpAY
1s3tOgOHCto2m3J4P6NOCgpZgaSXo8KDo/dXw6e4AZvpqm5P7h8Zldxf5Sls+Bup
dfZ44QpwtVbO4glYcsaHUVhnYrfzCAijktfuz8rPhTvkuHcgM1Xk8+55TW9+++BC
6WNL7xr5TmKlkhSzbNWUEclLXNZQLMgasxxqVm07BvtNAy9i5WgCMSHEu4MbyzpL
sqkkoKWplYzobrPjtwldI08BsFlV6K6zV0GiphEsAyB+Jv1dMkKScfttBjQDHcHA
dbbbUYWNhgAy+oUhICoYlQVAcnBKVEmun2LEXMa/Pb8s1vPaQOY/Z7fFNLkY36KI
3WSIwcM/enlfnQ+axtpXIIu0oaolE+1sJePEsin1J6yQf9jBms8lqJRq4euYslgg
TNY8lcOXuxFuyx7gXolxOMC1Qm37lke2DVUZbkbYsaRpRX4vfp+Y2jL55Ps6FwCY
hKqQXuytN5+sJ46mxTShnqnTOeno3P/x/JOJ36x+U4iDHxiWZXDc4B0lNC7Ewe2b
4kcHuFSpVlVTjAUZIjUBgmGfyh0CGjUGcNr8HTzrg8Ph8AIW1hgGosSdsGGxoph0
/N58kVBMco3cpb899HqTplLZqFzjPduu4lXGjVmGPg49dHvZ9/Sj1sO3czLIxar4
KtWEEslCnr3Rokf2hEK79ycwnWF51bpfNbndv4hJq/jRpcigVyvV/LntD6O9gn1M
hFkl9AxpFta2jzGDACP8QklsKrglu+pd6bqSbdzGfSvBJaAQN9EIJ9aHFKSC9Zl2
AY1oMomIpRBvLCWlXw/K4VyhGt9vDsQ9ryMEq/vFD7bGraDQro9g+g2yumaoVndw
2F6KzjQ7O112+ZbiTe2fsRdAcBaLdS5DpetyH+gEIrlzpxZYETudHsCFIicinh0X
PU+8vlbOIMIpb46WmFcWJ9DN6SVT7iDhnWRwd7FKphVMW4y4dVxycBMnin3OqrtT
p/KEJJAe2BJDpPlUPCxKwF+DeN3LQEjBrOuulUJxLWZ1oZj64+fkTdOUFkNPqWIw
MHpbTRYP9Nj3uqWBr1MydYjlUb9rl7bgQB3YzVrHGHNKlFNyXeMb2xik1d5uNX3b
f/R/XuEk+gdvyBoG/Y7WB07bm34alo+PRATFAoRMLG7zPIZ/wCZFasKkQnjYvygK
bKUSjI+9RdMsVbYfkjODNfa9AC3/PhFn7XaiiPG/3gE7Y08j7nOr7iMA5+7QsyEv
jAwJoBCKhU4jVUkQPVYaayp5mcsmfKcuF60O4wGvdjnpTjOeP+Es9C5RdgfyFHZF
ucSdlHa20Rh/1b4t5O7HS8JWwwuo7jjWFcMG5+V5Hi0DpUg43Ciz9qU8lk5eS+DR
6ChHpLuDsWPMwQRBEVc1bJfU7KOSD8D+ZR9PpAQKtAE+4ZlpmPifamjUQTUtuN96
fMTN7ZTRiiQqFESCOiO3gHVZ1wpyBz8gpENgjQkY+GE3CgSR3gaa9RL3FTSA/E/v
W1FGRG+Ytau+S5HTCiQKwgwFnQObwu1U9WY/nAtlJgURyZ5EQOWNKUS/NPHLcbrP
PIwZL6j88emIelzrv71kiCCqUJbPF7wLXEJANmh2pmVx8v0mbmghgQ7fjWHu2cCL
0t8eoP8uRTABc9SqpQkDL32Y8Q5PeoJr3YnafuZSqzAwzzNOaqmqk/GUjS8vIWM7
pJNi3FnOIryM5f6rV7I8dMFqMBipoVMHyYF5hmkungs0wZQ3i7R6dkDt4veFajdO
WDmV+Sm49BJn/emC5iEfYOYJqG50xgVnALP4XWv8K8H/yDH3SBCr1veV4AurFgMy
SswERRhwl0Qgjyp0i2jP2Tw5IKJKxAKvJhuxcNoJOOv1sX9Nh9MqmUVeju7pLiV8
801ZcJ8N4q1oGraD3sYVUr3Bs+aLaph9rhiv6AS+X7qG1Il6SSwFjdjc5Wtmdb0J
qyai1MdpkLSmkU/rbTouG/vdmeynyl41OdIfD1+j5ofowP6egE1uwJH5Cg0VPwdC
7OyYzho+QX1ceTmXy6IRw7EzCgFsavi0ZUnZmusp8pAy0duw09Nf3zoeIC3hcEX1
BXupFFpEcSoswBDqLmitCeKVvPz40IjdZzpHddjLotKca/foPFAEWwBivlsgzFIw
KuzLlQXzGS5eheW1LjiCKDOm06mPN5pAlsRbL6Za8ksiUon6zugcGR3NONNTEg+M
zRsdW0tJqksHrKGIMHtxpw6++Ma0xCBhy3eP3IAISbgCGTcrHIHCK23r+scTJmQc
RVLmFB+ObMKp3W5+zzDObcSMi8gRh8BEWfWNu3yHdV1dubnp1w30klhQ9VfOZZDE
W2T4DW1KFQgkeSUcQSDQa5EdfBkVGqsiOpqu7sm882kyjEjpSqqXPdTlHhbha5CJ
iuzlFBWpHbyDQ4p4Q2Wyk8ZXCdD38xIFHSztW/i9xRLODruTa78xyrOpJweGSph8
CX050xUxynJbhIJJQqHijSK6WL6P6J/lCuHiLrPoD0/R6i4ILwTokU0ksT9JyQ95
Dd8lLp9Y5Q83XGEA/yBx0vwFWnlBVep/DruIMIMZPbsILJJ4rY+i2ZGm1h/o+iZz
z1j/W0PMD1CgLErzUSMx/CiVSZ+jzT50fII1qeyFmvjtxIOX4i1KY3KuwJv4PvV3
BWsOPtn6HSr+E1KFdNRsWYNur2mHIlJ20E0binVGkurr3ZQwTULlGBjDvt0qc//G
TcrPtqej00MJg/+cxnlOS+FGmO8gs25OLth3YH7HcPPAEX99s6HP2UjEBjjCoDgW
3zMFljvgrkJeW7c1ItE2gOZrfohO56911is12S0DD6e7HQP/2gq5fu7OrkltqqDh
3hoTHUiAMYAxZ6k4kn7g9XOya/18QGuVPEd4uSgpPmBVqFCSHonbJd7US2Z39IC1
5yaQdGX3Vu+w3YmOaFeHMApbetxUcml+ZOawPR0JmyTQ6PCXsi5KYjr/kFy2XPPf
f+1ib2vbgQChxgMmfIb033akVYC4uYZ+yY4EJ4Egnu8EJeKknUuannGe3JGABH0T
e0IL40lhlmuPYddhClnfmCsczhzkzzSw/wrXyoabBE7DN/9h6R+JL8/GkKvwPB3O
wpWuLovE4lLVcW55VrWdh2xClkcQVimxQg0drr8uVYfVdY0G/kkrfbnCFv6t8bCK
AqaCdkuUN76xAV2aXPmzORJqbwufSZl3pPFlc36xDBmTKG78eVamPUeUmoZnnihg
HeuXRm8bpifK4Go5mudR4EyobilObFnWd4Vlz9tRKfXaMHX8SzftEqy/jIRYcMVW
qKLH9e7ArC/7MV20spF1yn11zB3W9sepLkWvuMkwnCYhFJkxs1WsONrM5aB5tMX5
sPy18GMizHQZndoXzVygk51E8p2NhO9yOdwUYTcXt+5BjOAxbh7eoxXDqUuemb59
9CRghjiIRZ+5y0mDDvUQV+TggjyXT/dLg3puaL4cKyCi2YZ+jq7FVsUSevUgB6hE
AdI2CtNz6KuoqSjyGeVqhU36v3CplPGpFePCLbDm5CGE+m5JD8hprcD0Fy4ozAWX
hDtBDMy8WLDa3OW8YIcbq7/R72uFoiV+rc1ty42EOI1Sjs51iwMt2EeO04Q6Wlpp
9wTzX/AJA9X3zCx4BX9qwSt9HRSy7kcVY1Q7wcm7/78Ri5POQc9EzXfyUJByn9Ur
M5Z5EGMkmb+nndEHiZjUa1DnMFaZYJxD51AlaaIFxvpN15eM3ND3/8Pab/606yXx
rGxDctfZVp8oUbC6P7wy0qW8zLfTjn1i5wMCM7boc0lR0Dm1VQAOhv3oAmwDI84v
4/nZH/Mwfxr4Ju1gDzud1E3muDZ28gPNkarmdXadxc9muJz7noiUXLxSnhsWP6YZ
ybQ10ReR/t71fwlJ0mqOivwuVmQVKTD1qREzczxu/uq5I0YkKrgxNJiibPqv98lQ
i057fajN1ryfjA3h/x35VCTfZeSFor8xrS55cIxAJE7Dw+YauaJvFSH1cqxX26vo
R+2ccPmckB5hAUC+DiYN6hlJxDxGQrbtYJ99yEtbKCXYbLx+XEBz25AFFGHdszoa
nocleX4aZ891XT/gotQ8HZDZpjyQZY95p8iGMLZdQ3o6GJ1jFl8BK+lNYAk32Sln
OqqWV05sI8VeQ2PkUCEYceV1D+V+d5FxGzo1tUd943yFOb+mqouE/j2j5GksIYaS
Hgot3FfasYAvdX3C3SEk3Ipst7WnGAImIG3Jo6w0jNbiUhCMXT2xqkRQqMEGe9hO
3msYKLwCK7vPycdno8jik0EKOSLIZDUnOfRsboYOWudhoyIGg8e1h53qHYmovlSV
V9O0C8sIumKQx8ZXE7q76QSy6fsjR1ohsQhNx9Ggk/3DmAj+1t0FEBs4OGJT44fc
sCreQDIGus2NukHsRJ3KZkm11EnOipjNgZSX/ZqGzPFQJ5969G47jsPLREd9JAdh
T3V7cM88AXe9pi4d1XETxqV5SHBaR0+tcVRka7Ur5hT0MFsFhXB+uqUHc9jV+r2r
1RKdVz3xerxXEMsrPkznQHM0t1WQgo8+GG97y9wiUZg/NZ17E6yL1/yWvBYHJpyT
FQ3WqTpPtP3HQ1wYfQnzO7KkBeoA1aDPzbZi9qWE13f87cGukCpFZAvHTYcNqF57
h2CMnku7fHqQS5RWR009mplSp07N6B6RqNzSwEGnvjzUCvhVV7TdHENaLbYuLvW6
Nl8xLP6JPOvWcT2XKq+Rd0lXP51MEGR0DVEVHDoZlaQR/EdnNx+NyTB0/cuU8HLC
76BWMJUdcYAR6ng2YN6LERO0b4T/Va/eoGXpmGo2C8iGM15rjLYW32Fu7VmJo0hq
CE++qr82QoZlbltHYZ9zKynVYz0hPXtSyJFnb1/xL8lZBteeOWfzzvoFWPuU18U8
XX9I7Eqso6aiPptlUQ6fUDb11RhMLdFLgVzvGlquVcDrMXmtJs1fhCPByBEZRpLB
a0dElLvbFynL14fe8e7YC21IJn6kWTfBRUqZE083l4S6vXHw4uodXfJUvVpyjyUJ
RfuRg4BuLAcS8YM0p+4AqfHY7TfD6QC89hngeVGGYesnHfTwGcQ/CdjS2kSnV7/0
+MdhW48LsJIa8x5yUWWXeFKXHgnJMW/3MyXXSy6cXmBNp/5y953ZjGnFQb5ChkOq
vLkGJ7nq3eYY4dOiis1c8ClC10zyeLwOyqERAC3OVsOWIykAwjDS6H4psvlx7UfQ
AbJAlGc30ElFZyxkmQ37mOr6MON6u1/Ur9nznoiwXnBsGVrqONE/Oy6N9w8CB7Xf
mGk3or/dBvaEKM+nL+cjcPTDAB3dlOMC2d1o0aggVMc9cu2bP6br6C3RLJMLt4rv
7SGE0jXuZOwxj6fqoIH4mvcRV31yrNIavnurpupqt7nPcvzlGRHP5sxARfIY5AAQ
k2wk6NOq/yXLlVDtmaighylRQxzHc3m8qvuVKF3ux9x5QbzTFl8D57rymin9ki7B
b/xlHM7c5zdazXpebwuliaOiVf+cET5SB8fMrQ5sbAtsHtoYkzZiD/bdsc6WoABd
2VYze1CGR6LXh+qSQMo245Js7Y53ttPaeECZgBHo3l/f08OoYyzNWnBhgzaHTc67
Dk8m1h7JUbJWhR1tMJRlUlhS3coYnsUWdmEBKkNuCu1kAhYMZzO8naBTYBml+JaX
5CnMYL5wg+M8UgQavtaG3Zyeq6c4JXrmUG9ZVGrSGLutqRo0ybDc7CKIJc51Al17
AOuQzlDRuUglTb/D/OlDTFiZcS9SUBdDb7IKWzVD5OislGEdjYV6kyaXLGHlT11S
ISx5B2TO0uWUO1WCvw+mZQwk6VpooHuNKXI2CbVMaphvjSjUhOmJTrqu0AX7AOiX
uj7koQtaKxCOJONOA485hDkpKB6uY/y9unjJoh84bvvIm0cbBLj+22czL9g71mVE
9Pk2REvbLzFzdY5VMFILZ0QlkuAt0A2yNUTi0HfRo+zS2Dc2rpCQlRB0mAiATfY1
gqV4Ib183Cv2+3e9XR9tJeX48nQjVfwtYuHcKEMlv8fPnHgq2aDUyzN9bltvcpxV
DPdkIJPDQ58KtqVkncIj3ePDVK08oBpFn0RLQvvCvabnV2eqmSkuUu/YsRUkvRE0
iicxG571wpB6QMCnGCqAi9AH1/+RS8ZBkliFKlIDnERuvOjo72togH13S4CzDs9O
j3jHXdoZOO1DYqhP0fI4xorkcCeNLvQmn1jDEyF9+sRaEbkBcQLzNIkkxMZB47tn
C/hjLTbjahSEUhc1Ar5AceY4IsdK9FVTIFcBxLpYshMv5wChbpaUMXJ2A07VJTiU
YDHUHE+ECsJ40tMWn1Va0CS8zXc1ErP1OfM41GVPWjvFtK4t4V9/GM1lQW14gsOf
TJYhSPu2LvYhM2lPKSwOze9bM2ToYv5c1bVXkBtwoplFVRkd0mHwsvIod+Z7JDIP
Ouv+RnrTitWNLetPSaDacJIQgtFIxPLUmU9Ci2FjkjFr2+KPtQz26d1ybgYdkUKv
bNFXu+HhwPKZL26vfmgAYXoN1cncAqBkAYsSsl9z33CrLwfp0pkEXQqlWN4764ss
ykrpzflmLzR+WJnXfYvGkand01M4vi5sXe/fjbum5q58sangfVcTWHXX+wPb8qRi
qdMxQPKyOpbNuIuBbUxh3boMCOPVDErLrwUk0VqxBEWaGpFEVNK0fhm7a/d50mQw
7EMP+gCWjzjTuagXqPYcC3Ao9XagecUehy8GIfh3b3YQQrUodSKMg2cQJpqjz2ma
TlajehwX9u0ckDeSlJ4/yuxq4YZMKr/ctrCbk/sPfwcMCW/N7OuR/Y5e7MFIhDrz
T0cvE/O6sGiWxiv56i4SdspuHG1OEiXOANT5dculDy8tJ1wFftFZD2WnJnHfQJWN
zO5zNVSKlStUVATlpPJuDtNaOyLY26BL4N7iXDJ+1zzp20eW8WvWEoXTVHgeVv/l
mIUC5AZPhrQEDgBXUMwuRvUe+hii0+hJb4ge9Di3ZxjAiGm3NGD6pvRC4OV96XOn
7byXEUssLoRHGUFEzmRm/3z41hU8RSewS5ARGNwO0r7boberZrJIaRUw+mlAtpQ2
bMOv16C5onTguh8Y5lurkq5GLr9m7dp+tKU4opvG8D+Wo3+McZAPtPMVyf1Gg9Ed
PINvp9TIxlH48ZiyjcHKzKkOrilWaUKEYXGDlYotWlJrPRJlU8zBXxGK6D1Ww4Cp
xZyP5pjv4hc8/aqB4/hlLi2LANdZn9yvtvS3Zuh5eTwFPlSZyb1gzsadaZc1mFWv
mvAg/azUgCWiNN1XRz3fZBv8pzb97PfeZd8WZt9tKD0OXa4Gb1ib1ERVPn2MEl+u
b5QVtFjwp/fzLZ06og15vTmDKuhYdUuv68xxGRLR0XTEGk+Y1l/axLK3BwmK6PP8
+Ynukkb6tDH7Fh46qyNjG2iTrf1qgZP0W+EsYwyzS3d6ocbznsBdTfkRWrvC++hO
IFivgdw24WC6tc7fur19ftfio2OMu3ehMfVkw3xNnSRXUvnnCpi/B0xbpM4dlES5
Jpc+891sGX85iFTRPDg1PVGOOzeIV1HBTjLM7flv0Q79y/5a2jc0/SXwPXH8XYS1
qYek3BWg4CV4+DYS7hmgMFkCr0/VMe2ojLxB4g5EuFpWnxV/3zN6F6JRDK8njNKd
pHwCeisgzdzzRg/7ALdx7b2J/qneTcfFIs0/2XpbvQwM/8QYeEwk+NpuyI/HfFG7
u4V/VtifXDnkLWcfdU9IAo2vxjI9wD1kQHaqHS/8MXiTRPZ9zYPszy+MY0+Jorfx
n3rqAbLUcsGlr4xq6V49p4S3wdS7M7jDUO+XyJCYoqyTMTK6NFVYCmm7P1zbCvzX
0BnU0/HaSmjbUdy4pvxLLn4o1vs57wwHXYeTtVrOnAJY7z6frN+AOGbGLif9CPGZ
LLbh5kCoJlmwbgOu80SqVZfqylVNqB1/M3WlQzyg0+zFmv3+ZaA6Nf/OWMtRqPwu
7JHUClD37bU6fpnQxz8C7qPYHI56CdSgxw+P9elendpp6bWO9idVsyrLXH1bb+oy
eTl83BPbrdUrhLx1YYOsKmU/UwDQAzO+9MC+UCBovmQELhgzoKSen0WFNGYnauO5
JDW6gq2dGOj/KeH82b8H594QPU4IjmAK2Tqn2rhu9KsbKnn9UFgd5t0NkspyRdWq
r7VHoEzMNK57fQFrfHhE8440pP36CJPV7vlsGrazI+T83pUfD/X9CSQI0YHYvhtM
EVGpuxvoK8SigYT2XH8X7ggpMUXP3rz1R47sm1j0hQxqnV8ZlwDltTr43s08ztBN
/uc/nDTu3/6bYz1kCkd+9ijNfyaGW/Xn/zaQQitjhjZikUjRBkfAY0V4AAQykjIz
WcIT25TgvCqb7iHK1bj3nr0FXkI1349bjfjQeQkbT06eak95xtS4mj6eIqaFlcej
/drW/cSqFbJhDcyuDdOkZ15pWehBr8JAbyuniM8f29/0/SHPdGT2FC7DYadqzIyP
PhScUDAtyndDzXihlcQlJ3hT3C2h961akkf4VZucpqwnrgTgBESy5S+FFO1QedBJ
K8W5bjRZQUnzXWldctuXuBJGaKON816cPCP+Jtp13CivH23Piplx0R+U3szSqQK7
H1qyJv06vm5Ta9WHIbYjZcKT/gZN5JGqumrA8Im6ZyqFdAzjg7rgMvx5GMKKxTdI
FeLjLJQ0ueST2P7Kxx11V4rrnzo9x42ScxN+Bp1c/k65ygfVSDfTHh1AtSbbJxeF
hlmHrJ7NMah8badj2R8yaTClg95C93JF6ks/LnrWWeau0g5tdTwCvAZ+C95dYiSC
4HdgmMHngvi3GLVTUyKPt19itkGdulTfVychlHn6mv7EMZql1YJ7MdAZWdiGK+cC
nUnFOTPj9vFMwZh0Ey5xxUu7OUzA97jJo7eBNtiD60k7GBxWFZdDcOyjXmXewAZ7
fVyPTCUSoppTOjpyVWuNvU2x3meH7nEYuxQepAbjsX3haTiKytbqXbL+jc8o+4FT
3UZeQjcDHid/dLYsR0NZy9NjTmHxqkhbhXmgjGWEQiPtri4nez26VOERkEjG0CP+
qJRmX/akY72OvSNAyqYj5pkiT14Ueh2cMv3c98mptTdOIP05BWpSmRfnmQ7y4PYX
1Wtpu5CjRbPhEmAbEgywRfQWSOfcv6OytZ3esj20+juc/2DpVKfbDOragXkAxxt0
2M6xaiRJhrwGHNLGpLxeMZHv+JswAqWUSMcmQdZ9aEloKJ0fiiFxA0YDAMtfNX7S
qNf272bgjlcSFfFlQfJIv3WzytP0GGHn5Z2jItnCzK9SQBHbKzHKtFFunhwzGnXo
e85zfRromV6skJdiUgDNqDaFs3AWTZZJ/Rk51GPx2QLY98NlG6MAACKrvPldKv7s
SRsi2KMO/Y+RRV0l/jaIfoLnWKp1wpIg49SRDUjb+iZK0HcR5K+NZ3FD/OOkN0wE
m33TqKZezhUOKFA2imQsDPyaHUMvCkRCj+h5BjawvOlxsL0r7gwneWDdloHcXWFN
4SdppadPYjjGaqrJq9S+vRuXopa9aZsJCvO5h4hOETsGMcJdIOpoie4977SMBKR3
/yRuphSPGhX754Q+o7/rBLyiEbgSVLpJHgVqywhzpiMgf0SHdhk4i2dLlp1qV3wr
OqQ6Foyhy8IGXzSIlKVExUhpf8P0aaqLFVI8xuNU74z+Sa0UMIWwMSnCBHitC4AF
Mxz1A9KYYk/QCc4U+vSF9a2FZrgZ2V18WiiyeDEkivSHPUqFqGE0BWTaZlMOA/kH
v9dSSOVnKrEJP2+DTERIy3mO4pTTglFkRk/3ZUo9l+GbToSIL/AuNwLE/B1gO660
s4A1gOjoKrXLCjSQG/neuk3KRXmOixQh1vzwd8g1ZF3jKJaPfPkYx/qASpsoHVg1
FmmGsE5xSFPhfix1dPvQWMNeAXN1qJOzgDOj3JgDSzM+Ym0euKrBwvvMng0BIJ7L
3qy7azbtyWt49CaNurEsAFXC7F2ouuZr7zzlGj1P/RFiFE0cVyOMCGA6Ah9ls7Cm
Zt1TUC9/tDu5Fxn4yuPsQ0XgeRtdPhpyTvCs2KD49Zg1G8wME/SPTOZOMSTbIbj6
/6errWwbGnBi9G29Vc/f1Rq9TKfqWhAaKpcrgaEo6/B03DRciRktbfrvmV3sNE5x
eyppg/5TR1yxiT/NGATcgFp5ZaMudkK7UyH7N7hhcq2TH8iT8r/Q2IIeSiGItz8/
v+UwEsHncPOcQrTIy2V1jpM861KKEn5HedB8mgYnb/FUcXhfxmZtOUQoOBgeMDFq
I3MPI8GOsNnvs4bUOU49VgePv2YKjS+QyQ0w5IkYt6OCQnUfudR2vCgnP8OQQIZC
naOKMFJZZd1yNnwn/KeDsZ5nBfHP8eNQYD31dyn+wsWlObseDiqYAU8iUPT5D2vE
64s5jHa4E88MTfz5ETVEylTbsbESGBUdHVEnsKmhz7zr6W5OjQ43/yNWfw9tDlMC
bp1KSDlk1gRgzH6sOOUCTO1ahTRg9ss2bSqaWeVC+VEot5qY/MyWOcm0c3QB7LUp
vOZlUS1cRWv0soKlGOab4Jzg4W0lxIocMHpuKaeFEs9OwpsZtArKllGcEFBIJ8er
ZVNL3edHHZKanK9Yv3YX177KwGRaCyyKWDuSz1SKdlL6NxwT5Av27UI0oB6BxJYK
mLtjKk8O8WUgKbfvLbxUWuq6hofmSR1k9GfOfCUkOrCh/bSO52A/4s91TaGwAd21
uNKUy8ES7S3WgPJ4vBaHTXylL/nDJzJ6u+NVvCpIBZvlreFvyNhx+2bOBWQsOjdX
MKy9NGfe1qPz4rY83kf+hbmqKO0cbhMl+fo8bdv7Y97YNffk1emtO2ZPbOiGgfbf
QlSZlBYzmZXPLE+JUgqXUwdHXqZ1MQjY6ySQZXZTqC1tHdhxBMHUTT+2AcvvKwc/
tpzBUa3lSqNWoyCE+tSQpUUFfKHtddEU5uwKQIDk2t55Hy0EhiIZZEXCsMYGpp1O
MqDSaZl9wP9QOkFoyzB61lxuFnpDyn/r4qpAJRryngdbqkBU0jECpH7yL7xHe26J
9xQY3PeqBchkKfDhFSEA7SaQDyfmLwPkmgVKb9pYrjKXNYdpU7b2bEDaZcFPD/Oi
VrR9rwew0vKTKa5ohX1gJyYONE899GJcybEjyK6lQL5gmM5I1ahoasLm9HmQg83H
bds6j6RLNGUhzwVcZpZspnETY7tKA2xhYXc3da86NwU6RVUsL0LqFpCgkc5DYbg3
2Pw0EI6aV7vjmev1MJkIa51yOBuR9E4ZPxDJb40VlrH4cGPKWcQplje9cMbnmjiU
E36ytMsxhAp9larMf8TrHOsRFZXURSreOG/WVHktv/sVuUCldEIR7qToOeqEFVgw
uJWCnlSnXxDoMSGNM0YyG8L+9yHBZbHaNPmHDJ+dic7fUrOTDOKgJaUjO9KqywWR
BiRHnbSzirp+UzgbV2M7iMItuBbrj/v3eJIve82aml5YHM4xaKU8PiyVZ3VrFCcY
dmmTcNi3CDi0J1RIFZJIiu1DfaabCZ5Y8ToGbgbeU1h97a3KLxozNkzye4LogF4a
iV0APqky9is7SFB4UiwWp3yE+o8zZrVNcaVtt5tu2q3Evyq4+OJyiFlQ1tc7E8CV
fTuuxZ5u7032R5dZNZJlqFCD4+zDe0L+vNbzF3TGtO9FcrjfY36K5LtJW/zm3nRd
bglMbtFWhdgpuhduMV0NFnpf1DWwbAQ792sF22RVIu+L+WPaYzlezOdiOy/2FRI2
dSjTnXbRsxCBstW9bskilZURzUjtzcLYYGrFilRItcz/lF5svH7i/ACB29rq+V3I
x2a/rScFHFx5Lt/7npNFz4eszhYhoYQMVUI6N1QVuxha3kG7efF/A1xQq3qQJdU7
H2S56UzbL4vjox4sH9EOd+DfBec4czW9SCJy/wdh3DRm5beNvWQtKQOzDRO9TCpf
vLDiioPLMXgf2YEliY9eXtJ0JQdEhxxPHP2hLzxKhFYVmtA8Ghgn8zfYLaULQdh4
1tPFD5E/sjR9c5s6eHqRvW15YVeQwA2jenDg8V++3W/sI3t/D9YKd+dm8/+NQq2N
ZfFRuwwL63bPoSShw4xgd6Jhm1850Ipx9Jgry5HfXHoSW1jqOWGDrq63quhH4jK2
MTfnEmAQxknqV+OGoQhfSAUNld9Z43lfLNn1eP0epBV3YtXkKnORlJlexji61iYt
7sPXemCQeQDAQFHM1wALUDaHaunDH+5W7wi1v+WAYh9gVjeMUrEXOp9qzOczz5sB
JUmHm719x09rda0BBtWpRgYI0z5x4vpO+fuOHMwzwgX/jjTfTyAHMT/53DYTOYj7
2hbvpiYB+3RdXGjQ+bh0f+drG19unEVRGS4bQ2EBWDOcFz1FFwQtqATfRXBi9OWg
wLixP9ECXw14QQiH+WGgCb/vJvQMxYvYhniuv0foh+Qm0mEsGJGJE3dViDcLt+cH
3de0oYhPFTJVVJlYsSDjNI4T5MeEAUvze8C1DuFItgOiv2CrHu94qSgqDOFkazf0
NWfR1kCaEDVI4ATxnwfxlOx82VI6+YYhvvCz97JFCSttwE/g32gd+yuH2S/gtf6m
gSY1PKJBQ+oLswQK12w5l7WF5YLgfF1LHVR7KKQx38bV81DFa8nIyOHTZ7gE/QfU
5pvzEKTZbC8bzUyktB161hXOd469oLs4TLbobyygtuwO6h0mLmBRwDr8y5l/tooe
TeKRv2xD5UhVFySC3wIgiVRjhbozyALr1sFP4RFLWjy99E8LHMqMbULP1ixwFDvl
PqFzejtYX40KdHGFwpOAUTKZn5AC2GRECztl79TJFF8NoOpPRyMAJjWpmvOymwCG
oYTHMUdhWDHxwu085Je5w+At9reJOsayECMX0w121TTRdZzv16zDl2GupNm0yZhV
iwu2Y6EpLp49AcMBccbIv1Hp/YZ+NTAICAwmmVpO1XW73lrC/vP26kc/P2jMrqd3
ccAZ7CCG49kgkvIu/x+4DH18P4m3iSYfb07QYNFCPVAy/v0R5JRFJXf6nFqamvJH
ng5d4Ir4afRa6K7cC1XyPZE8s+iJ49I3AptSMyDtyzY51Sj8H7L3bHepGWDm6ZAZ
y1TR0w2Au54gA+ulImZrXKT9FPoEP/4H9R18HjcrLginm03Eq0zGbWEH1y/pHQ0b
63FhNoanNEUeUvvjJjYu4xlV2Keq8nqxVKDG2ZlRPsEwjNsCfMV3mHiCvK+PmE0O
KnjxOtjXVNdWQKWm8IDRwY+p64fv0+YWVFfJJS/AbkgNpDNe5YJ30+IjYMahE6we
HP4WbxtraBhA3Yaj6pTZFoMyGAL2j3YH8yIdvC+iMkRWVl4+BN+uT7xGMnoBjCLF
LwN/Nq9wBRjlJnHSQ7iz8HR37bCobumQvSTdoNMWKjFIxzf7ZlVgtTbH25lN9Shn
a7rr9aOH6zLnXpbrQpmQ6SGYVQUULDNrSPDK0ed8n6r2F6VpxmDAnw3C8F37Gabr
NW6UlACLJKLyb81LPnIu7uOc7vf1Lgk16WWq+kiF4Zm5TBkh8GtqSu8D5KhD5Tzy
URLqFyePLIVW7i6kqOv7TNclNCzmgWDvw/rO9AfEL5HVgSxedzWYu4xjEOV3oxq4
F8PY5xMF43fZffDYi/KIsyQXAzzWnkyxRg4toGyTTZWyPyyX1gTmStiX4EPrarRm
5bezGi48tWmejF9tS9w705BHtaG5XRgFnwosiIGsh/3a9NWXrC133KaYJHF3RlWw
kCgNnpZiBBHOLYuRKVp+VXIk8qIhzcDX4JvCLa7aqxa0EotPR0iA3PnVfmAbl0o5
ErMlbfatZiaS/cOhWUcB8VVZYMFYVZi12sbsBshRsQpTuje8d98PErtPkFBNn3vC
qkvezGea97KywDQ/7GUVPS+HtPEROAxzbN6UqEViYMtiU3Msl7eGUFjg3E/0abwB
NnkiT/ORleRnHNYQqdSOP/KeBtb44UJMHwxiOdmqQ/HUtUj0wUbpTRsbpBpjMgDb
aObzGpMVHS2NPHPKspaUtF8W6DrlUXCUm6nR49+b7I434qJt/NC8X0Zet2ZKkPUb
XOxpCMdN0zDP7xiNd3JTYRLK5CapUxYt/EIDi7U9CcoPtgOwcSlRGEOQLm97Qrmr
IagPhW4VQ4idI3952OV/7bS5CJCsv6wctZFr8YSIPlUZORp4GfKTdVmDrTMKsaTK
E2qg3AdSyxMsOZzKDaldquKLRTBtiAaEyU+mwdh00GEch6lketIWwYVC0fT7jyBS
Q/PvmpsL4KQD4dgcVE1vLPxMDJKrSh/804Er7dKRlJKMy7PrERbTLbB7Dq5/6Hv8
/qp2SRGXOC3aD9hgj2GO9OYe2MhqaM6qJ1oLsNMkASwd7FbqS/eW8N3vmLejQYKf
aQBoDI7Jbejq/EwOG/iOHPuoGN0jcb+EGlh/cEgi1wJ1yl1YwdL/jeXpdMce3LcZ
wCCtW5Ughy2mLsHUYTfw9c9XvFZGKR0PJWyZVyhmcH6yraZe+TGRDdPBdft5cFJP
X6iINtiyPnclmafNLWKPpekjbLUEtyRemzSH3xnkfljmh3wahpUu1l/nqA7nybYa
N6+5XpE/bVkV63z730tNcM7Rhft0s3ljgLNp8Y/cf1xL6T1a9Nu+RFUixRnsuf3G
f1j4WqnrF/FxKRpcH3q5dwtdRNkE05Gwgop/3cr7eFWwYuxaNB3rUwA4gCWrQV0W
kJT9MF1EG809xjMH6I2gNc3EJwn82kGcZZ8WkaozBwYIhby6S/xZFPiVI4P9oWwV
TXlUOH3BB32zjnbwkfG0DzwjfoGaj+rx+MZb24tN58WPkhIX8OXhaaow9YpOm4gi
4rduujlEnZb3lCvsatOC1xdwdiIh7/9nZvhErKQS/w9lucSpCfhVs0OE/o5qzfmX
6tXp7jF8/aC22F7alTkbhbAmUUd+eFcSzf4OfTvBVQ1u1zg8gn1BX11A4lD8uSTD
cPuHcOx5Uc3U+l90hbDS/7igW5h+WOJ5VZZdVfgd5vo5PuAQRHYRuS504GWFMfXR
KGAE0kxQj2o8nLQKWvBw0ltnfLhnckBqrA4w1ztBWhAzGb5zn81v1T2QWu3SdHlf
Z0/O5cfMskH3hOVq0/YS8F2BlhOvvlMmwbHJfndIvLNoPG4++UZx7b/88f7O44BX
mvF956KryKnGzENZF0XDc5OPusm3xMEswSWAfcuM/IDVKvrlvcqSiVhWBAMmgLPX
4we2TO7zgPZxOGolznjqHCwupy+ah6N+kOyWtDowxZdWqRBOVzllRBMaYGnhe8sC
LY+RkNdeQlZinzHTvTh7kVGxgKB9qmUWZ9Iob+iVWO03q+RDY8A4ZM1rs6gnW2o1
LcTiyt6WK1+tZj7tVChXUn8Tg4KYmXBCRIL58wcA8Awz/ufPKgCrnw17b6G6hAmz
yC8cW6S/BB1k5CipEEPfVtMxsV6GcjYcCSNXkabxnPcpzMVSz2fyElWEaMvH1lCo
IgBZufB0LZ+ZNzkO6tcNJl5NrBr0jb/PL+uVemYJNjo9fIesw32mBQ4TBBh14vrZ
FCP6fP23pWo8y2JyBE5Cfq5r/oitbruSHdWElmi3LiyL/Obqpn+nKR4s/Rr60sp7
lu3NrlE2sj1jFiP4G4A/NTb6b7JLD0QfMSZrAnpTCQXytU8qFuvT0PT77NGPqz4h
pinvxDIYy2yPob8LY2EyV0ycgj2i5AXlD1HbOiNE5q27VTkpLsckI1qOZjod3g/A
ss+cpv8G7O+xET5IfyEt6QvJ7cCPl8/3d0wLGywhCKe0IK8gUYnbpXY9XzUNev+y
E+q0sZTLLSjqQDcms3+xpsSO/eo6eeBV5tvOOEw6kBv0mjtGmPlgoeLz8CG4LPBX
D86bedstjOWifAW6/+a2Mv0r4hDZBB/9ORIJ17tCrJhOmygZsjNAjIXTba73hsyY
0137uWGxoh1mi4uRtXB5TQ6HFhtKizhEVv53RH6dxjPs76JuP4zlh5pO9dpcb6T1
tpO14xYagFVjo7Lgc37DKkFbBGurNw6lePC/0TiOeOFUBLn2jT9sVqeIuwfOLfXI
bXw8jw7IR0i53SD6V8kvYxpYd2nQ/3eX5C53FHzbo9um4NzSwyaUm7KJo/R7JT5s
ruiXyKwjSTwYqFZl0i1NnTx8k73l0Vma6C9MTkIUAECPJ+K30Q3aPr9ZSxjrrtcF
RH7GPXSIkMwkF4+nvJNvsAWx9Pdd+ljTDzIM4WbF4t5BIPBVJjABgGFxt+I+SVMd
6EpOBTdlfMxhJyT1Qx/ls50yVcijDfYdH/mwd+OL5Hz4yero0BTg+vv/6DwS7S3K
BUmHKL2qcLUWRA3w0gnF0iYEO0qHMJVnIlpBcdvxUR6vPyug30aYBllJIjupG5Dr
QDlnzcrS6glhZVHojo55ffhMmaFeVrslWr66ZdPrg3A9lZez2IJANKlnWFullsPf
2lOmW33vDeXJmF3mwCScjhSZRX6vmhpkeBVJeWXPa0bToCiV1IR44z93xQemZfhg
GzbH3k8PWhViLk38i/U+AnmKwX0eDhsqtP8H98JXhFuuedSmzIlM/399KvEsCZsc
PUQKE/UT2NYlhRIDsjURJDyJkZy3dbhOfhdREwbN0BRDKAVKOVM4bqfuvxw2bvEd
RhERRoIINa0EPwQ97lMNar+33W9uZYQgfccob7w75N5OBfBHZYKhG1ahhAgN1NOA
i/EAx50kxXWm4kJqfCRAL8VH3eLOKZIIS3hJR73wYvtbit/BN7MxlVCpN53ErXts
gobY1kt6860IM91vdyDzCaIA3DCTMZAwtN6UHqWlopnkNbaPLeqgPZkt+hrrrAKs
1xU5jn/qrfCGvJM+plhm3D+uSWlVciKbLvuTIT4WropjXV+HhrDn3Uur/HkzVi1U
5PzLF7RCoxS+nARGbDvMkf1n+PCAJIEmR+XHyM/+OTC66qSpykXm+Am/mt6WVxBp
pW24sLnod61iTRPIR3u4q8sHiRbPi7nyf3Qy2ZgkuMQzsaPXFzdrx0WqMY+HM1r8
f8OnNwnkkB9Ra9/3pcgPA8fa9makxJ6i6Fi6gLmp4L2fvJ5mfZDsx0ngXTxZ2nO5
MmykBHhJAdQUd/65r1IozM57zHAFI4+9y313z8adyJ0HQToDJM2PS1WLorTR4GKw
78jfj0oI11cb1pfXX/EwwzKhzGH5uqacF7VbA+yPSWS6Cl4+xJE6F2JZ46ykPJSO
PdHCyPXzGoIO3fifKvzbMDxuoTzwlpp71ql+OH/aYy6thbG7kbtlxjFcBXYQ7LZq
6ReHxS0vk6qt473gLKPoh/qfJ9Fz6JthT+8sz78bAJD3L/hvHwO0fIX2xDiYiAbM
XdzCX1cth99c2Y+6T0zdI8vXxLdI3OYJK4W2Cdez7qd00mwxsrwW6bVctoiKEzjA
hL8PjirM9i3AiNKtjD9ysJijJ+visxjPyRe1z/lid9MBO4lfjO5zHqJLzM4G73Nw
uJ5Uz+SCs7lZO3qduFwN2GUtQkKd1tHb0SypWHDHKlKZ6w2XPlvclmF/lJKMnKUy
n4pT4+4VUyPL/r3Ta0kKyrD0dfO9zIorr78oQBtIxesLkWTpnLLLBpkiLtZQVPCL
NqdQF2slQ+LekKMUqA7FDinJ02LAT/OeSlOOsI7Op3eABBqgYkRzpAR3T4AY6N85
RrtPKyi+RW/aRoZLdS4XwLpPFY5bZ1ypCMkrHKa1LXQA5y81sm6eu6vDwOfhXn/2
kh3gIjy9qaPXQcieyNKlRID1DVKQfqN9u4tJTes5hGLPMMrPBpwo1s3wvk4rKP8J
LNkCtq0685Bsh6yozAq6foYpD+IT1X8d5lkqD7xlt5W9WF3opb3dHRgn79lxnD3t
er2z3kN9aYKs4qWoPHOY2P+ZPLETNNno0yW7QLn/E4b1kJ2IOiUXufm1mDeL01cA
TMBaAXtcripYKLBuwYf3D1rNdEm5VXeWoA+4zyEj8dOGV6xYJZe0ceL+HknL7XXk
jUtzdPCbmqNf+L5+IbksiX7BTtXvt+jn1HUECkEEvYKOlTluX3yJvwlkU6gwAtB+
jCtU5EvzYsVyyfrCWyhy7XT6dLaGcwrY7iz7RsDbxH2m7V9rc7pZgHq/mHKTMIjU
f5/xC7MXZDezsbRq0HZV2fdz6hSi/9FqgPrr8ZfKE2iEqlr3xz4ChHDAtwB3K+Ex
xDmZ5/OYHudB8JOcXaDWwwpSoP6yx6ovHXcYQprNgatVwF5TdMuDiA/HRR+Avz3x
uzeO05rObUCb/GhsHoAT2L53m3zJKUWtDl4MKtXfR/f9Hvq50GUEKqAJUPF3grSI
jbt635J6qpXAGWcgDes1wk1iEVcGWXlJJ73OTPnON0ydFbcimv0d2ua8FS/buUsS
xDvWY2i/+8siB4T2oK9b7YdKjpzvR0T7xO/rk1SEpKuvvnZF8wXqk264rbPrc9+N
VbI6WWMMWxT7TfijiLzjmW/lf4w26Mk7px2QI6eTRg+vvGgM+Yy6mctr4F5y0xDv
KqGqkuHADsc3VLEc9g8u3HP9/7ddQt7ACpw0IFxPSiunsHmp/N3BIfcywjIf7my7
kuOKtWrXk0pl5UD8Cuy0kdQHzEpxUFUHCrQyS0wUw5Cu2Qv0oUaC8tHQEnrG7B9V
aNVg99umW6ANnQOd/qmZDS1ylRdeFfOLWimkcUsLtIgDWZ3IFbLNJeWZ98u3bh7L
xriW/vNIi9EAo/mNk3xBOKfQsIMS4ayuG4c1q16na7Uk850q0/Jy5eWeWc11o2Ka
oZViJnmJIli14MZXIx8iR/4OZS5dZIuSGMRMulKNTNqsTMVjtPVbF5gldxx09/9Y
yEwgJ+k0dLyW9Uwte8ey7esg2NwV5r+5K+XQYKWC7tR824/48HG14RC2tF3TB4hv
SIzYMWINI/S1aK7zch5yB19RwL19+X+Cqr5NbEYRxgRQuzYuyAH2B/aSr9l968jy
ZUlWve8QcQf6F3XK+W5jf6LtPFS4s2Nn4MxfXP5cYPsaHGtUWm3Cfy2+SK5tlgqR
dYzbtIH4SvRc5hek+eYTm/p87Si1wRomYsjUz/lW72pJGu5m7SBLArRDiBQX5qCF
QDPXJ3e3Nsufh0cinD21kmB+WmoteIRqQE0uRBVZCPiJuLMD6+JwYQ4M4r9tqwB2
oQqMz4255miPKPUSFy3ApceJBQbgx/xi7Xjf0+OxAca4d+mXO+9jlyrvBaLgtc0y
fz2zvDkBcDpqrz4iJ89ChfDhE4Mv0qoBBmk0HRCGTnd0zSVfL42zMfSwDxVLIqXk
MEJVsy+rwFEt0xjreJIwpj5x7nYyD7xd99xbhFT6TOYo4WLZ68HdPjpiy9nGb2l4
aK1bNW953vEe1BQiTaIbnBicJY5yYRuLCql3XmB1/N+aWj8hx+uTTBnG7FxI1fwU
EppRzQi93Z0RbAMkDUb3jSKrovWnNbIElv4lVFOG5wZSReBjAbDqIDUBFwKex1oB
PFTwQeGb/eBvISuUHmNWpK0OAXfhcVnTAZqMr0GB22Yz+UO6efDVYuPpcHaEr8YZ
LRtI7Vjn2JB2hwKBNX/uCHsHC/iKI08wT8eqTDndULXALtKnhrk16d4lidV4WsVl
OzBQ6qZQ1ko0FHhVsSVe+QH/gSKTCp04rBCEErxSNJrCTX8R3uHcE7BbGAENHb3C
oceMqd0TjfaLX95XB6eVZx2DXBOZEJY5omEIsQIwrqdv68H/d02mTzbisC7FAoek
eulG6m+YesoJzdrV3Cedmz4QlKCxyk+wFDVi6rJqPH6cpEtCqCmhFs6T5Nsd57cV
l5kst7dfKeyYwJnXmYVXL4vwCHqT90yTRy5iTKhIrg5+I2B4iwAj6jF9l+eIWE3K
yWaHVcjGgRP3pPOCt1pv8jMKeD6YAWfVEMTa6s/9HF2pvJlGb5Ab3FSe4VUbz1Tp
hTg3pNDkKm84aWafb3C1e4A8NBQ2ZHWwLL0IOfiNQkHmNlnfuraM0Hrwuq04zC3r
/9LtQyGftQEjdgcRnFj1AkpqBq/UbhZPBvmyk6vUar0WMhNTP6SXvFovfj+D1TXy
LP6ayJ+JzTxsxesW+Yav4XWf0KanPivU5uTKDL1TmwNFvQYw8qGqZHsXk/ZysVhb
jOc3niLOUHuJHhRuAi74/esaEh0Cg084eMm0ORs+3YSNqIV8/1HIXbtuXAWmDZ/N
AShqptoENNBsi/vC808VfZvDcsg0OHMxzwQ8TRjaO5AzJSJ63yxYF7414sVJgAd5
m44Ftfrox2CGhhpclsK8KmDTpGuuGZi+fGf8k9tulDPWJ/hJ7psyddOh7zmIaR/E
7NraxX3d+mB3wsFTKH5Hahv20Xz5rzfTdo92x7otEotWSIWWhfrSOyTxud+Rj3j2
lLnoqAGiCzjDjUJphzyFjj3zeJGKkbT1Jm1/ts1IiMRUjzo2+mCRtyfAwCZZhVj3
zfHshU/rf9Wc2ooDsbAG/HZPu/1roEb65PEmqB+Q+Y6FwKmEFhfglBLaEqKOWOdE
+6+jVs/TIOth2gww38pvgo/a/T0uJ0QuJnu3+s1h1Oql9MOE4vZV2j4z2y3U3JUn
aF81vu3wdA3OBgEgOH1M67JUSPJlTX+66HVV2rXkhxMwpTRAEYueUE1+1ScqSHiQ
C6AH/uhmwqx/lAhrG4qeiq9VXpO8p10W2eSYhmzCZ688Z9Jhh07r31WZsq7/qAsw
kIz9I88ldzkqYTfUqy0ali8PSmFWTWt2EgGRZkD5Mhr/2UELc23/YsqUNO8CnPcQ
txqERurFckzKFrI6Hplb0fuZDryQEWeYJToMjg9LGQxYyjmxlZ0wNkaMN7gP65lG
iO+bYiHzv1RjW7XBznAullaI2O0RDdJv+DMRswbLpZ7/Z1vj9ijF0sAh5dvT0ArO
pxmC+E1Ps+lk7W9phuq4tB+0w+R5ItvZINq2xW5MoJxbBNfaEGCOx3QjhX25ojOF
OwsuqQkJLL3iAkiFXKWKaALlO3pTdt4CeqxqfAF2iSdQjKxc9EDdtCuv54kAqUdw
tr7pcGbVn/GcuTvcs5fGQkLxUOKysz3RFwah9dV9l4TmpNh4P3Uvwct/l9wuLfkx
d1pwN8g2FI2dej1VApbo25myyBS1eU3C6aaMFzjksW7R3nOU/nLXunBR2G00ADXe
leY/uBvrwAmoh1Q+FKCfo1kFfZu0WLN6Rb/9nkAH9dDUXqo/QSKCQBBkiNykIQlD
APDkBGAx5HQ7IrQHEV/N5Pp/ZTnjgPeTNZyVzidYA3C6rp80V09LbMfHj8XrMQe8
BsKVf5S/tTBBrRht/ErAiN50YLqR+NKztewdZMMoaiLb+f9/9MgjtzDWUlGIOWqX
bvQPHHwQUwMsezeAl7unfFEZTFwQxMppv6zMa1rDtsetOrrg1EijV2a98L70RpNM
jC0uZ0L6BgqpdzHKAvcmwVWCTIf66aAY3f6ZmIgl1To3TcIFiXecXWAn7yPYroSg
5XNUxXaqPAo6ceFESkM6NnS8583ta0DpwljP1XxycYfmqJpliH3mhRepkV4R4vw4
fZljbV1wo+X4usZajM6jEeE6BdVbWP4KDiJCE3/zBWBhCTRY3kzn0Cm+d5VTjVVN
UbagqTRBSb4hYMit7bTV7HsdO0W7j4UbN+ZBZ2aXL1ZXP43HVy7UroroSF6vTURQ
ZSHgGybCoOleYrxbFyVs3ClUtPIQsc7a9YCBWqku2jGiaK4hUuqyORnfDczUjhlD
cHrOivRXnGOGR+UIQEMiRI8f2L+jFFXVVu4MgrG/A5bjxtrqSufRvZtXZQni2DsR
y/wkpor9OkUcK69tQxCezy3mtGZ2ZOPWsi3ffjoWL+R+zbHC95mxqK5bVjpNFECt
I/YYu+GpRpKqKmQRX5R0UbpB8gSSBSmtWXIIH0pfjmNuC4uvuVL0DRwB9xWrKQFZ
SAc9k5XF17svl4e66qnVu9IfPfu6oU/f9iAft5KMJEaLspLJffxAbgERf26GBraa
DCykphoxT7vDVvzWHpq+gEQwoQlVPikNmk8Vv+CylUpj3hiGReKl00yYMN4YSpOD
CVrnp6ltAhOENMg1y707nKKyQhb57p18k01v+g7DEpq2G9FQnIYYvPW25WbJe6gi
1P1pDRWWgxffmKTIT0W8NzQXJmgFlihZoVY1e1jWqjOqFKDrVjkmpgJHjOx2Vp3C
xSF8+kyFAR/RJtZp1m8/qzdTtkjtR5DEF35R8z8cug0XLBxHMUn9CstA/9Dx9ud0
zSi7kVJZP0RhBoiDMakr7IHsO8gMzCUBNIqdO0SYfpYkZrIM+15Q/7FXKrLRQwYa
oXgRmAZNoOg1RgNh5GhEN+bfKCHeWCJuSs8ZNyq00YLWeOpq4joubn+c/SyYtFwJ
/xTtoYHYaCCiDD58FNqY2C7Jcz0fACeTlKpOHaoSkqBjPN8rDvULutl4rCqgkHM/
rBVFxX1zADE3qTzfYWVb1AWs8Y+PEhOtSOMPWRD5Fcxtwb3iKgGgqpjR7v4a9/bU
d+5ELnoiAHwYp6Ti8Azku9L6l8P9tYRgQGlFzIANZmfjrn8LGkttkeEi2KSSlFYp
a5KnDWtaHipTm5eDXP5jPINWXahORzJAX+9FnpKZkWto85JVWOACXLtXyOayXjkZ
jmwzSYrCo2RN2rOFX4OT/mXGhL0Clu/AT6RRP0kvdUO7OihG8uFNCCh26n333Y2D
xvkKYk/UpxNQxKRjjtf98dsJTX5yU+5EOlYomfGDpX8Gmc3RX/agA+ZFU3J3POUu
9C+ycE84rR6yp7mrpMiYKO13fQSrMMYnOaCIIEiSXHpEE251rMYD45GjgLx3KKGm
Uq6+afIxKMDwTqO7ypbog70+N9CYw7jvr2y214UFhtfnSGTwqXNN8nm0+dcRvzfW
pZW2UWUNrdLTXrDIL3/7Q6aGs8CjMXTr0EjoLZpsmHuY6lDXl2mq5Pz4MoYCQgio
8VfM9/Y3uC54d3kt8ibuqLR96X8X4LF1/iNpRMzqyTLMVF2OumIMxZMH9bZZwizr
YwJ3E5ywEJo/xfl077XvNRfNOH1KOx02UoYoz2aMBZjvVIlTMeGubmR22DCKfMUi
AReApEyXKb71j2gaePfIqEzepavBFgd6B+YWKYkKe8WKZB7mG6L0SOyepvpCToBP
r/P71hIMYUiNQBTXJC7g3Vy1etu1hEjtzIp8fi2XGATOMHxTKRCcLglmBO/ljeVv
9FnqawBkFvDw6ufGpbJjbN5V8I/lRSRaRE1O7bg854dWFFlyg24VVaREHgkJOaLQ
UF2hh10+n8kXlynDYJ/J3QwSxpnO+IkRunF1VQUtM21ZE7vVmMSmm0y3kkiaOnTN
vb16w6bMa8SxYsft6TiydQHjUhnF+0EvpUFewB/MFA003wOR3CbuiXZvQYSa4BwE
G5M9Rd2yp7uiu87xehrVI/xrh+rlT3BKOG0UVyCuLycybweO12TpRMUX+U6BxLck
u+qcCJDaoO8s2O0iSINV3xS+nnbQ1+Cs0/F3eeF4aFeQ81BWQs+8bGFhHX2W8Rvw
rdPsDesxbhaGUvm5eB86dJagABTezFYqM4zitNP3NQJAYa/KCSQHWyv4ytkkuWEV
4odvrBdlGbrRK1cFkOYGItYLyoF0TS2d+xfbH8fV/Ruke9kePBplDJ1/KqigOykc
aYfDIOt5bJAbskUgGP1SSVdZqzs/ZQqEEUfN60jvndDxrV8WpstSAy3mgBHYZmQu
ctlbRjCRG0o0O1skDx+sNwCutftTrhxHi65V98CBiUxQ6YJk33YyWBzwO5/fTCTQ
fYf3A+lLgeJLXWSNnAPltCIiPUXtvCHjC/Tgl/1E13WkzXKbBN4350xwyvfOOEk3
CymFXWc+v/AnFxpVl3mHBklMx8zttDDX5Sh7Rvv3JZ1rLYYJB38MRA4lKEVTmS91
w5uNgd3glmVYzs6pocJ0NoxZBgsumnGneh7DGPUc5YkIu2ipKVAYTY8X9P0Cwm++
8dTl32AYhtLgoRu+oDAnO0NtGgYSOUDzzF9OzeYJ+nF0N+6/kLmyp4OC0j953Kqq
pDLHfV9+PNuVW9G8RCKJ4yng+Jnw7EUY1899DH5B03RYyYmGEHpAKx/k1n1MXf2Z
8lyLkgGEXQC7337K/hK7eZAgs/PBWjUBGM8HJmgylTac0Yw1aU4KYeG7UmcBKFoT
06V5h4bf77fsVOug0zcK5lUyqAniQ7khwQggM3hf67+X+Qaeps7cGVZ977n7FHbN
XKASK7poMANIz3xEWoRd5B5XvNfC/jDRzpHdGBNoz9WnfUkrTaYzDHfiewOfWgVq
i6pk8Wmpy6xDMCzQvlIm1Rh2QgNaIL/y+ZwaGGQ4cMb58tsYn5HxVSygkzyQ9XP6
BzZOY62qdQikfLtQuWdB6tNFopb7vP49XvNCnGT4oYlbs/3gJVUYhGBSg65YJi86
160Sbe8mkhtTih7BNhuFmml7WHb9++Gr8KnLf+XoEjThk+Njcy/ZU/1zBXoo+JUF
6YCWk/YCZpmqxFompxVGw3ugGqp3jBdcMNAOVyt+sZjl6oyIlpnyvuIe3jHq/jkC
fyK4YbBvmhH1kmCKQwcE28hdoNu9z8xAmhN3FPfnqcGOdiT8RzDOYixzRqcIFvus
V0c8oDDDVXHBqPgFBvdaP24Uzf6Z0exj6HBEyjjvhNU+9yw3JOtuHIPG+HSXZpzE
m0Ni6eOLIW2UKmnCwgwjgA1y7Yms5K7IZcgEV7Eo7AgbXdYdaeb3kCb+fSZOm3E+
yKx5SdYWCWZ+jtyEls2NVlY40RSh0kW5nuIXyGRL87/jFymXprTHjhArhffVjrgG
2RPnMaE6b5M7/upR3hc+rQtCMpgDZPIoaR0DHmA0WLiG6CcIaeqGnC1Jt2VD8wn8
uikDoz+xy8JWGSkZscnOPRUhf86whm0nPijalPCo9tzHQTtcHSFEkaiBbcv3zlrU
aDvcZveoYWrOO9eZGqf8suvzti12KKOpwalotXgUr9eN9Y1aThDPMhqz1jGY099Y
i13nc5xELfjrAmvHxII1JovOLlRwEPxzMfveFh3SwTGCcn1Uq5OpCRratKxDRmXW
2S+2TXDCAWYLInGBoZjohnV43bVB5lhNmk32n2R6NHC0Fmaucv6tw/Aq0F+nlfox
4jwpMdVzfYS4OHTyy6QdvQqvnn9wPRzO5lt4XkNi3qNgCAcShEIoTLPUfEZbAu9R
YvjU9NNlwk6CoGNyxVreiM9Xpyzx7fDyt/pYrsw0ydGon8oI5Rf35eiO0HjDUM4K
AGVLFdTMNhf45wkehsTGHTMj2iK92WfKW1tAl7VCSkYBeA+aMQASUZkitRpvv0yu
pvK3Sd29Jpus2V9dWoArLulSRb1T/VUHoSkYz8r4QiTNuNlrZPpzvdoUGAeTlNIl
f5RPMBBQvPr9avS55rHD/kv+mT8bMivn9fEX32F/NicE9kix018Qfk6xTNR4zpvk
rBdoaEmfd6QGAE2+vYWDopQ9l08SMP4pnjXeT8eYdXSF9pI7xzU+LZwFk0d774s/
qazluZxHnWV0hRGJMsbIz3cS88T/Nr7lR+AT+4Gr5snfhhIkCB9KX+DLKMh382GQ
faFh0djNTyJHabmakKmb6x6Bfqe6UxDW340mN5YR/B2A8O8Hc+trBZXPxk/8honI
WpHHTYoSgMemctEZwJIXhauEG70vrxmEsFjjE20jIQz6o35VNXKYEy6teVg2Tk5p
/38+X9M2uJdLnSSrm1ookNIVzJwz4+ARS2E0GO/ZQ9Wf2gDpb988WSW0uIpPRtMB
GqvcxOL/zcEprBpJsF4ujEfdhLjbKyRYLzDgIRxYeCNqNpO6Vjm3fggwpjMw27gf
kNIVE+27LJPmwv6PkqrRvqhMbrylo9KmDnWroE/GaZDGBkllw3q0HHQR2BEMe0jL
ZHc9XManMRoj3dLSQJ6GgmWXwhXLmVoBWg8Fx3Lrj2sLa4IlncP4Nv5dW72gEyHj
CUn6wFwJAl2qAXHKkKyf7snN4l8ii2HyK0NrPpehfUGncMwHyoVRMBAHXThR8jzX
MHjUw/QNE4RkdVbbu8FIQlXCEUXAAX8SLcXqkok1sVNaCzwtHXch7YEYkJkZ2X1I
Bxjlfj/c0foR3G3xT7nLC0Do+DAVP5KXRyJ5N/M8x1s9/hb6xiByiVNCwi/Vn1Ha
9pCseDg7ZhI6mvbkN+hu9EWvV9MVfaE9N9VGYzXaKyarbuaVD9WURJWilhyy0cFq
Og4BnhljwzIFGKAqlobj4WDJHQtgnm91VETzbNiDK1cT8IW6bNBPQGCblQ8iawNo
jsCSm6R6cOPTSurt6CDBje4KwGhNgMHQCb/mX3GyD+bqCyjr3+df/npt93hJOzoy
hefT+rD3991bmV4i9gTAkihQMjtBbmwDsI92slC5Nc8pThKk5sJYSzXQlb1NeK0u
4pQttOPWmV1x+ZChdCnJLVb8CZo0z6dg21WrEW+ktzmYaPczchR4BKeZs+AexWP2
h75rOQFAEtAB+fqCaEB8vb6bl/RfAXDIdMU56Bm46gMLyRFgOS3IV8ZEiuGJsoi3
up/OjSQCTGuhisgNcVMikFG/bIwab6LPxznQeKq+JgRX75tG9kP9j2muTSBfLzAQ
cgNrV3C5KxJ6Z00A+mTnFGSm4yd2ZbZcRdNxkFj7BtyZH0FztaDzfCiiO0StjzEB
pAc2FSGxUwv1O8Ec2l2MR998kIeeNPqPXFfTUGskOKR0XRaFAS6K3Ht0umxCAcez
tzn+nLDyHWxT5uFp2cv/2xOJwX/HlCN2wCBfyHJ86xy0HkX+SPqyiUtcbMk4tCl9
7jivdVksQZL5M0GS6vQcucjF8IBQSu8+AldIs8/z7Mz3OkDXS91fIEOkf9QNtmRx
YFphvRpwx66FdaqVNHfNP6pWmYHhSIZcO3ge7LUFkTtikU/CScjmgUtPm43tEZQ8
u2jNVzK831S389kA8EpedcTFVRR28ZUydfZLtgI8+V5Op0JYcC1fspmBucIQa8Mi
CQ9zkdr5OgbjyXsMPCi6gXyTT7GQa3ODOCA5IWzAaTWi0bAEaeZw6QeT58Wr1h0W
zBNZgGhR4u/nmUVbVbgbFjLnpjSwpyuRwA3ob7M8Wmo7BDNecIjQNzaRxP/uwVnd
WWj9FqkYa/ZuT1sECOkX0H5AbIts1iP1u7BasQBKFU73s69QZmgx37FPIlH/A5uS
FhctOGL2d1wa9cHRVUJ7dJUtNd/IVEJxmlrqFouUMsNOiHqD3E61Wjni4B74iLkA
BFt/5yTBNtfYt+KwPRxBEDMhpF2yq4ovwTpsbd2VevFnNDLpVkRVxNC6snRoQlKg
Dh8AIWjJ0MhNK9negFqLqm0D7j27BlcjGKjkCv7TrNFpxAQpWrwI+GowO2IXbRcQ
isdBXLeo5D6aUzzJSjk+F8YBdomgfLIjnQQkhZMW0H7ar5OQXkG7KRtQcm1i+lud
FXxR4rNIc73+DqVfaTeInPWWHoalpYw8riabrm3ttplEj0OPCfhNGTaSvjcblsp1
zisBJxggCfwrx5X/5WSv6WRGspJOMQIV7YB+uChIdTcKF8d97GwBHQ7kXPmCFZWb
U1mJp5Wd3vfsKbe4i4p9M0T0jT3cytMl49Tq1VffOMpAkyBymXrmK+CkKGdDFH7v
ooG4gUxWwqQEMEMeqO+xMZnFyRSemPq0J4aZhdeV2qOTNPIUqVJZ4wk+FkWIFcNh
gFL/FF6+MHVwUcSBlVKYRE0ySx1wJnWAvPqWID7Aors7LYprvLnaDLZcOR3nTZEl
ZWvPZdt4J0ljWzX0zlXl6ayrrUQqj+CgV0El2RVPSwnPMTDRbwFrOaIrmbQcXcmK
om+z7dCaQnZqrStZq2kvEKJ79xAjrlBADGYutGC/jV7fpXPbwF6UNo3nsFmruxu3
0Ak1qsnOU1NbSSF8nxlHfR52xDEzzCSCxr8KJzs01k+DEVBsyMC1yl6GvuBKPXic
UYmyiCyjKZIm546NmoxgeBMzfkmR77qG8IXkcaV0k0o2uuG0mpC/K42pEHCZ67yU
Vuz5N6e+ycNevHF5smBdNO/OAnmZEtRe8ydtn7uzz2aBaMOOL7q2MgiFnpjebHj8
yw7fAGypyRZivcOnhdh9LOAZusFI6aSU3XGny5Sv0hGT4dY5/gEgLa5Opkkwz4HJ
rCXx25N5AiWgcAWXQgiyb1jK8wfZxGGji7jY0jsiKxaN0wrin2U2vCpljUSC5NN2
y0DEelDEzxhCNa+wSXn/czseQirir2oFxl2/NaiKqxbGbquV8JSSTmWIKGRi1s5U
5taab81u5/HScuNePsAmeI7tAb6/wKNsiJ4Ya+uz5ABc0xGWLnVrc7oymsdapnPa
z3sTmkRIjAE8qXxu+LTR6K5ZV9RBcMycMAyZSFMj1aeam3vUBNrqhUlrmSoS3AUz
CnfAPlljVEEfOxo5FtO1xhEN0dvmU+qvw9eNwxcd1JecItR9lBa27TVr1vdRilhF
0MBRI6pa/C/elRtoIlNsb4ja+IXAs9DuTmXB/AHihIWoBM2BeevEO8RoSJ/MPBSX
v73ubANeu7n+KWjSQiMNTywJFlkYT29vA5z7zIUu94N41qWx0YCPX16YVvgrL95l
3C7rBm59MVaZeUHaGbqOsfl2v+8fLF/EHoft2cYs7o8pBqAf+wEbIMjK/j9As3ds
yldbhajgzdwWPU4JdpF0t/Oj/NONq6p9XaxlzTGVEerf6T6ocrOTpVq8rPl4HRp4
Ln37tsEyyWTHL/RfzqCxEihgoprra7WhDM6XiDSlTpRNwfR4SfaPLyTzwN/gBNzk
ehtZfBJnhMrWBqyHCVt8f1pg/fkEix0J/NIwJyyNEioHiitiIRjAhDOcCdCP/Xmx
MM7DEpOXcX87+A7TSFyrnUihMOdVJK0kWMwxEL5J6DEG30+IaPthuWI6NuLtEDPf
kn1b4OGex2oNqSLNjsfbJt36KFFNfJGTjZRQut6anaxBxC9nwrsfFF25Do2xdviR
ka0wkyn3dN2VWbUApnqaosVyKBXMle8KD058eonCcbSSEAIKUWMMzc3rLZnUWAPf
iTnXHkQmp+HGmCxC1w9YeNhWJ73eF844ssD9fBIvuNKPWzdqBQR5MaJyVwTudNKy
D+9aupFJapQQKPC3inUwYZZ+FLyeLEh9lcBgjjshyLCYc9O/M31y6z3wIIgVo3U3
t4lzuuQtIJS+HmKImw++Fta8PDDSkHjd8C7kBrNCldb4u+ZXOxhhM906UyipPCoB
51dpa9jOFFWkHn7gdmeuGBnZIRzzjqtBqb5DpqeRSOTac+BdKlTZpJUIeVWVcDOk
hG1DQm3S1DC9WE4A0hpPGRQ1cJB/NJPhplQKgvvKczwMwSaCsOetrsLr8nZR2BXJ
BkIZR06zQRVIKWgKhF7JYA6hyTRJxNHgTvGSf6Cp6pwYhC928hxIgmmnmOb6sLCG
K0628F7WHYGuaefVJREob4qj/qKyeRWKpfmnKPw6MJlExjI/OiRKo62Wb6nvOapp
wPOrZ19uT04nw/tDTfwmjwGco7zWqvlNIb64S5jsqaPgBwHP/6IvU0bEdFZ/gD3W
4brjaZWn+qSnTFhVA2ao26sbVwWi2D4GUgHRn92jjEI46sVqwxKxXcg65KhdU2P3
KUelQRecIME2tUu5F6zMBODhrOLNxXh69BJUP1K72cOuLo7py4Eqy0CSCg9EBP4V
KTjn6emHLanFFzHecc+YgJbCgaDJnXCRvLo6irLHksw4YTp7zQk6XVGJc7uY5w/H
rJKrgmrvGlF9339cCb6wUXHRMaRGmIwyFw9tC+rIZqpXgytm+oc0FE71sGCs/26C
Fj6lu7ZTjFhuof77BNXC6sId8IrCB/JZDUjMwvZ9j3x8BS/m2Y5/Pn0tMZzB1jxx
AvqW/H3mgdE2ZF2gz+H/EX5yn6CmnTOkdwwBCqElf5bSqQLdDLyPpr89ZeV0/1Vj
5L/yBwZNGukY6VHkgT2HjIUCylLJGgeoFdKNW5blLZOhGuQ6khFdO60wa/QbGeU3
5ee8zQ+kRzn+qzbh9WN5l5xLND8TyEIaUCnd/jz5ix8G4jO+ZKiOMvLnft0wx/ss
BxkRJbb0xwUO1+KxyzC+87SanbVc0dcfyH9Up+AnL3QAUTMd1pEo86a8D613Hedh
cRuuaME6b7vO0dx7nlV32ssT+xOYVru4tqbS/Sm4P4C5SfHzAIFtyvyzJ3dwREYQ
B+O4FK71EWg5enNvXtFjB3LxeHh6Hf5NdNf6tkS6l96jlVew31QOYDdab5olgW5d
fzqqaUQRSHRzoLDDIaE/kkhdpjRNu12ZvphKF56vKWtWWFJSsGslGN7bbixqvWib
90HF/e2PBONTFcD7thYBeZ+zH/zfOax7OX+ZLjv0F5FXUxpiuMw83oV5+oxBYYlY
ruVLeQu28WFYGIffNBIgILqWTfSSCzkLhhRCWtMTAtsU6mpNLHA/4iqh6WazfWGa
UPiTBVUwgkCLL24drozGzdAK2vtmAToV/i0PAWNiXHHCIQbD+v/XBSHbTDg5RBuh
1+44JXnR8+Fy+VRvy+W9fJNG9cwRIRoqeZV21apTGAm1BLPNCunYFxixTRgc8EUt
OkfzxI32U6hBZbOKWzDFeUy2j4eHvUfU4/sk08FT2iIwtZ4PTlQmQG4kYRtdJWQZ
Tebz/CPmwUo4oTz1cjvQbAH6X8xG+DJrJPHpjKAvjyx4Kb50OxTQ4kSlJwL3P8LR
AtDGAk14UVynGpvwaOfAZwFusRBXVp+FiLU0qWV6ksJr4LNOELIkHszRgZrXkGPW
smSbrNyCYoNyyZjKZgR4ov4OAGspYlIP6HXnV2kg2aCVfuROMj3oSRbjah2gm0pG
LWvK49nZ1mXwhbvXud7x598zdIloUsG01ySwQGnNXQN1XDyCbdzbzUf2BA6+XbIk
84ACwSZUwlga8TmLi+4miKTGOTSPaXyApSUax4dhvgnD7/pt2quC++xnCCg5Y68O
FNpAwM5TUqlrZ5ZWjmjAQWsixXFK/jayeMZz22kwDzqw2xyJuJY4H5m3ekHfSYf9
FKbZbrZ4wrN2+6HGJQVduZwnUR4bFeKgzaLysaoMx2hyy7b77L2b1NYYhkvgt/0G
vCvDqMD2sj1c2MJIdjYZUF2uE3gVys3yEWarA4I5aEOvOi/a8Vpt/rjNo9Gbic/v
xJj95HalJoJoBjuzLRyDFaO1BW28Le6Fm6GcDDmi2gzY10BTqdIitKHeZ/EjW3Ba
yLxdXaHCoSld1VG/lVNHYRcdV43AhYMJES18i9xT4j9BWZjIm0MRGcTY7RRDdU4P
iHxhA2RSTQ0EHahagK1OzM07Z4dRsHKEGH6rauwAzPY4boNwJkAyu4zRynWbwjIO
YnwWW//H62E9W+0iYGWCHnn2ayKCejyuta9IW8ke6AIoA/cvIaSK2nI+b3dhbnsr
5Hi/iESZ2nmoxNp97A0xNF2JarWqT0PsjmL2xnt3uTbOfHBEaDn5Bp+e5Igi7Iwe
v/6lGKBeUnENeZgBgZtifPi1l3jFyQEXJJvL8oxCu7MkYDF63Psrr7RbBAp5fBJQ
1DcA7xt4+SEvtMQ6x4awRK3bnJIP7TqRiZcQE/fxKn9wk+ZaF9xpWjNljbtkrgpa
f++Yi6yskyD8dioNxQv3GUAIwU9qPMuiwuOdoxm9o8S4MQNaqZBaqkiFPTkZ3jsS
VKuotmT9GoegN7S5hrpLOcA4MXVub1ElEsFPdWYKhbt6laBg8kIHOSHFQyOYq+uk
0hdPu6zHpGKCsQLbRoVqq2NEgmmrZNsKXRs1S1PHwg6Dp9BmMDatRP6OYRKpQmKZ
XkfsLpxaDjJVqkxLg480omk4Bwd38niTUjpOzI7GZxTioQIUp8RK5iowz2CC0cI9
Tjr9bFCtFvoOCEaJvCHb9FMQuZVVEsPbFJpvjC4y7ylC5W0e7xzb9oj0iXoIDQnC
8QUiXDhKkEvRk+Xw1SaqTHl2xVCDXwEYL53pZkVNtw7mVaNtB4JhzsZmeH7u4io/
3G90dqDeEdhTsUvSlva80sRY7R0e6+SR9jTl1AOAhKdyYehfJBSX83n2E7oa7eiS
iOSDFsL6sD2fDlQA8fb1QNfhPPCBE7JqGxsGEFRvN6BBFet1Er9lEhJzfpj3PMdp
vffvNzFwO5sPb9rYq0jAvaqYZ443yMQz4gjgeTRJLB8hqw105+kN5G8gtkXJ1GAU
9kPxe3wW3itfb1ZLcuBFJ2sxL2SJphCMNI7eTB7ww2jdpC3C74EwV4Bw2dVv/m32
N1DRRoAT4x8lcmEQIXWcPPi1uDSS734nZWxljXf+VCxwHEJ3JD82rZsrow8ZDGjl
t3bIym8N8Yn3r2E4HNexQlzlu753LXJyG3QalgNDqr9d3CwL3YubhRE2JGBA7sPF
KZXNEJK/fWtAJN+EcVTgjsJ8UtnldrKy88ekcJbvw32zLJxwPeTZx7I7nqxwzTnX
022cK23lwDJJp8LWkX533D+BO77Ub7CwGJ//hj6qiKGhmMdvSSDHNYQNOfVdFlHQ
A5+yivIR4Z1EbSkhuiEMhZHUwg781+lE5AJcOMkoQTqb05KGYm6HFaOnSs8Af+4o
sO3K/TscXZHSJvsRa2jqPvzmr4BiCsNK11IkbEmvAcvn3K+ImAeoOzOGl6Esa45i
QOHnBkOP4p562fhFebQxIsdFHZryZSxqG5q6nSjEHrlpQ5V+MVjeQtFqeRClgcJE
oidv9aqVjv/eA07iAMydlL8k2gtH3yzg1h6bmwTp+eOeZKV7hQGobbuiRKWiXH7+
uP7nnVWZjMm76L0fF8zwclLRX6rGH08LhFIXJnq8DoCT0WKlTVYox0h9GeLlPi/o
pX6TMHlUrWb4HTiItPvMqqECneuuSOTYkm0jP6pUbNwDhA+tPoKrqwkkI+oR+BXh
vMh41hv6C+JYgHLGd+HRXGSP6F3ZgTm6PwFuDb/AsZYiPHS/potW/sWJXz5XNw5P
s11HrwPTxeU9+nYy26kt9bUfCXeaPSrN2RVaWeGFsPVE7lTbEAqbpe8e68Y4LIHN
GV+gGNRv9GGlHTmKlDWMq1qjkmgM4c2BkfgaMu3PurfnY0AxN15UtKHyNIENKSif
eFATbgEyoArdBjC3OgZIYNM/TTbRPAHsYCGAz8UosXvyOkvpRzUZhhONzKk1xVFK
Q8A6qZIQ1H4s7v4YLjpyy+p65ZTjg0bMG/JlHf4CSS/Sjkl+PEyrViFjqOWkwQYK
PIo6/gEodrZ3FWjfVj7MqSEdcoKzksXXc64JuCRKVcf1MI+rY743MsPjWNJORQks
a/Nz9QeQ8QvtOrJMRJVS/JHY7FC6Ll3ncqVOg2iceF/2FTHZDiHwuX1xBy6OfTur
3mtnV7Gahn3uH691Ouus51tWa4g3FtOm0mE+zz5PDPuBbxLVoWy9a+BAB8rJmuc2
c25+sQRqI1WckwVsxxke6un2PWGNJntBfNITvvRLmSHz+0gVGIt4/PMcjDQJ6a6w
9SVfFmKFr8I9o+JZ+OrTtduWH27NglLzq7MSEYVVbsCUzdpbBTq59p7JqW4m2xp0
+7ZetOm41a3I5hEuuRT6CMrFRM93g6BHad8HPJ8/w3I2PlVKRdISZ2mFD8vEEQ7T
kGvavRag27cWo/abZT/QIrqj/+cszsOZ48eEV/iuD9tjOlGgiABg53DcTm0A3h+C
CrRkzRzO86QiH/vwO1UnUIxSBHsn/QoIJLvDOg8PsssTdlcAUiu0dz5wVXA6d9dk
PteEMaFvh1ky6xOCcDnCeeRQ4TA4Wevx/EV/QQ04AxJ/NU3cm8usQR4Brv0tGWpl
F2k40lya/15oZUNJKCY47KLlOUhOu3TFe19ZpG6yQsOSZPBATeIAKZBTukVHnWGt
11DoC+/z4fAt6m3RHb3jinCvC3bVCBMiTKKhutqeem2+Ccoqqd1662be1ckzmdjR
hwRT8sppfFdsX0eqDE7hE9JDsB5gyhX8cOtFt+UWB2TVMfMMCw5iznsT8d3iFa0k
cDiy80VHo6aXfGgsQ+UCADEhHPeqvojXLlMWJlTBZaVIkpTKBkq6wM2wNoSB/Dse
z8cfClPRMtEx97OpW9UaPzIs4W7v3p/if81ANjPPZLBDuwzApFXqszFI2q3q8QbG
OIUFjAmY9Jdt9v+Y7zoxA4SuN5JdS3b4+PIG4a78fN2mA8gn05dkRpb7Hq5HNPjJ
5WvB5/yxOVVV7Lv7LiLQkLISQwwIaxvT53mNRhLqnkZA8CjYMAMoaOxK3ozAcQnc
rLU8v1+MEEgKg9dmnDKaDEJ0oNcA1Usxf4OJhQHb1Ga/Du2ppP05hx8JOcqJPR4f
A7Qm7rintbkZnQlOtYMR8fR0NBGLLshdJsGPrUXg8zJyFa+yRGW9sBbwuuTdEN4A
LQZ7r269QNHIVBrZBAQW6MUFkjaTUVqx+NSs6VsjBOi6NI0Sit+phmg8yhcy797T
z0QadAL5SRqA2Ys6gj2hl0N+Q9UN3KxqdIPuvADAZI7Sc277+Gv3SNVdAXjoiNeH
0oBFhQtCzH78vcohK4mMtopJKROWo8c8fqw3M9JPl/xxnbs5vltlhf5O7nhMjeMa
Y/Ls5MeVGYIDLs+l2g4oavqaNieD3XDczmaKwNKEOfjdEtrPhfmNbcquL1/flp2Y
mf+ub+DKaVRLK+/CV3a3c8F2/mxbZI7AZJvi0iGxj5MI9x+yMAZIW7fxmq4AENb4
l4VHyoHiFPik06yscwUObpB0v+AmuItS3FC3Nh70D5xXPk6Vfh9y1QwInPDnteS+
4WdrLJDxtANKieBQfTUkxsfBccQ5K7/BivenlLsV29k8Z0gSJBQQfUYe4TrSmUU2
YLH7UkTfnRoGtNUfN5micl//fcoaCLwlNlMgG7RUFQD+TIM+fah55/vNEtdOlevX
9Ae9q1Tvutk343An3BkxRnIBipGEC2e33eDB+RJoNZ0RegDHKNMJIkPjNN3OvxOh
AbSSX/pqMF0YNgjJTBsFLmI/K33+5vadu/3ceMQkxhPD44YIftkyuHd0NrJZVTS8
su743Knjad9hpWYv8PEfcNuPu68ESDkX8/dbTFDK1TgxeVPNclELKrspjD8cqVU+
EwrIG3ZcG1F1jEfXmVU1urK2Q9Bl0z0h4xtWl7J5zwlFDcTOhVYQHsx9UPH8BcwI
0hjn/D49B2P+bmjaT3AAKSdHtP1d8JDSd/2JSBsn/0AdYKOCenN60dbWLvomZCzt
7WzCiqAFih66LTQWijTeoyadZXJZq3KJXtUM/IsxVuPgVd+SpnjF+1vUznfOEuPQ
pH6BVku51DlShym2N3FRFJAmqk3QgCfhUEeLOo3IYCdylklkdAeSXsaAaW8s8Qgs
2HFxucoTWBjtZlEUbi68oAdzBX95rhpcCTs3uKSEcwHXXvYD3LLdGUAjBG6BI0DJ
+BFlBZPHfY7w5Yb/qjBYOylcAOaKPtqrc/LWNkXBGVqCqba+virqj9v70lBjbEKQ
S3x+UTzWhwmeuHUDMqIbZwYv5jjB3sUqriQJVYk7AJWup86+TLQN18lmgdQAhJnA
uPgMLc6G4oE7FvhCU3JcSaMFMeKX1blzCXh3NqxdGJN4mUabCHMr5oEY46aO35fq
a240pwoynCbPjTVQeT6tCvz+0WZOBV7CyX6noBcvsnZnrAqS5r00C8xR8ErNm751
wrNn9vQyZdak3O1AyAtluTrPF/hSr+zH5NRR5tG8KmtYOZwXXtuxcCqQV9ILUG8D
IOWWjcdKMtfThIUlGVgOnGC0sOzzS/VQ28RpEIaLxhDksGx13lpuP54MlgHkfZAg
WIi+RTtr0cuCYZFKGeVKWMH0NKyP43A7mbt++CDudMi8jltjysseYLIBh/FxQbAC
NtIg6IQ8Jw805mcA/JZ+75nnYw22gc6oy5MPu3UHxVFa/9KjCByNt+g1WxaCvOmY
p0PX1GJDkBYx5mVtdd0Wx2n9d9daZckXoZ8AL5OPpQhwG/3dcZhKh45v83uvT+WK
q++KX2M7PBPi/PoEEdg0wtRt8xtxbtwH89Zuo39DhAXItV3KwYXpcpm3gs4uHHDV
4c8WPLy7oZdwat8IGhu+K17zugpDn6ZtKBf9hCMrFbTOVUXgkPInxoHc0IJCnZJF
7YVY2o/ra4xYa6BMDxc54A+2S33sl1fdLw+G52C0yH7S7NCVb2ndYe6DvwOpd5Eu
zK34jsZOWVX9mgcBg68VkT5accwn561VK/dWZP0ybaMWivhTFZaGRFkJFV7Z2Lu+
y0qxIOuL3y6y+1mNSbcIChniuDpLNCJ8PlE+RXqmwyULYT3lTcJRcQwJp3ZsMslb
Rp4ndESZTDBojjpZwyUvom340L6iCkvNGA4GOHhl4IIyfQq/xJjFOIkbhkh+P8C8
HtKULqfe5Sf7ZnDOYKTDkArHo2YNCrccjsycwVKPhPU2RtG7ZgvGY+jjAK2iYlGR
tJn6Abb+MDoeIjJEOsz3ZJKjfpimDt7x9v0yiDSKTdpZGrn9Xn7Z8QevWJrTuGD4
8hvsfffGVybJnLTIYzg5DhpHz/jAYtIfBzut0tpAStNEVXyku9UouWThkGaL/vvn
Og+EMoa5LbulScafcNPNiQ8EnjjwOry64b3t6GE588+GsZ6l5Qj6rccMRTLEWr5X
kN+l97bv2wdbp9BGdGb/yj0CkQ6FVPXkv/NR3G4xJG2dFe4QeaR6w/XGMFQ9u4yB
YMYw1PIj8pa3B1JsChhbqsAYL24VRzC04vmDY5H/R/szxx0ibO61pE9IcPt1fziu
MdsPZXPtjJbNvJG13srW9R6VCv7+w1eNkHR4lGMvgVG8s84fOxP1IeUPImDUlchE
knImK6ldcIgUbYFCYuOgtuC7W5w1Os8zTWjB1A+ppkz1PBmFB4/qYvpKf+qAc1Do
FfQw5rHc9+PQ2inEnHMyTjJNCooTQbUfH5RhN7h+xm5iE2IKz289WonSGIaLqjlB
F5jOjm7pi6F5v5cMywB/9DNKQ3mM7+vthdhZq2jvxqQY5j3Os0uq8vegC9o4BJQl
+a1MssmBeeKWcl2/ofuxk1Oix07OLbVHFyNH8QQVR2b6qLJGCDYUZfW+wSxQVE7F
GPDQ+aHTih0TrZ9ScozaB3bP0iKVCGbaHaW/AmePq4CZ3WHBbC6HHvIPS+SPSryV
DbADcRIj4i7jEEwRz2b9ru0NmCYwacmUZ1f8MWS5XVMW3HArNvuOKBKVH5fQ7FqC
ugdj2lTQZvAYkqxhh4oj03GhsWCeG9A2TSTK05NHsJRK9BxT10HtOUJElRLWmVsC
WmOFwMBCW8LkaRSJdQEcQgBnfinc5otJ3RO88vNP00Yk9r18TCyDH6vdY25Nn/be
Rht4ajLPPdL8kJqkpmfPPHVw0+PECGvjomh/tWzir5w+X5oQuw/RtB0MsrcHXrBl
xeagi/QuhXPa46xzCOBKc5ksFFS02HrgXyT9d4VN/spDMEuLW8IPcH1xgdcaaAqD
yIzLtad+P8Wokr/mmtIvmIohBcOAi+QfBSBaysiPenJ74yHerZPEDqlzV5RkVISd
6xsDMGhrvyfKUQezeO4u3JEsYTvp3KW083zqwUO/2GLxecRMC29DB8PHEvLF7Pjw
bPSj9XhejyqCNq9/3SrQzWssI6Admsjz7WCxUcCGdciHR9xXaaC07WESyakQDw5n
1erO4nG0kfmKjZHyN/YXZZDAOYZCcfdciF+1SRi8htb0cW4tGN9TH9zCTXGV0VzU
1mO+dx46qcnwKoCx5hHNh7dMkfYobaOC2VxCoRps2Vfd7BhQdZYO7k6RjPP1gUA6
Rw9ingvUI1lJ+fj6OePLG+1VKPRrvCDXnT5qvUQ5Ofis4U2oKIkEaNqHzw92PjZF
y86vxYH7satfc0fbxntapwrJoPjNNJKUWqv7qF1c8uyujhrV6R4RRqQcOrALAlRf
1D+6LfQLz7OK3zp9fSGddtiRMnlOHVD958a+ak+VWr21S+pQ+ziaPwSPHiAAF0SV
E/bhtNw75gwrKcdPvszT6vUtPprUBxZC6VsgUw13p2AWS0MQt2kLeB60MnRljT0a
ghlyTmok7JGlD5Mj/OXZ2drUT4tfKsqeOqJRG4uOvAMyLgmbcWa5c92VFE0AQ0cN
fnoxBJPpJQXr0slQvxxNtSW1RUhzRvu5S1n2gyhDIT89KfS7UAmQlzHWi0GD0im0
JLgojrh7RPEjS4DAjY4oRz7iXcgnB8xfPox9SPs3qcup5YDLPxldv/PQK7KefZzQ
ESOtxMHODauDKrTQXDASuWJSasohXR1SCbvYYbbk+9KLoSfi0utecyFHFlt++SY9
ZjE73s+R7Cq6jUL8zBsuTQ2MqJrpzEwyPng1vdXVRWoHJTWR5Hp9Yn+gt9WBzBSs
gZEIPtNG7S93JYpjkVTCeXadtgXDwA0yLiToSvRBHVdeHkfZWcU3bP8kpwNu+dhJ
seIRv5hraT7f6er12jGWbIdk6TGWlLi0+/gb0TExfZjrHUR0mF6HcIWCD9KuVBxL
s+U2I/VJZwsv3Bqc1ZpyEw4GqfosXATk4JyjuZCLpSmhntgiQKkFfKTceQGbzNyK
c+8vYIf+mNIXuzt9MkYcOBEOL4hrIWeqrWGTbNxwsfs0AwaS9+L5EcBY0D4G14u3
HTuF2xZPWmzhnJudnS+PCTnWBTouGJdcZ7yS1b86m6xIUc5UgWHE38p7x7TfgDUk
aNeEG8jvB8MVjEm2NUvw3CQrEX5UpBRFgPgyTGzgM8p4FfyCEFcJfzu+TdhAOdBH
jv1+nI6BATUCFCtxh5LP4Pp47Z9wRYLlbKJSDkNaq6jDb+90eWhQalOR6MJWm4p/
BzAsfFEeIPM5yAiGxv6wqnHTuz7wF7WixbWXrq+7YU8NpXmv5WE4nhH1LFHs4lCe
ZQ5+/qYRJ8f0r/SvhBJzUanYe1leK/8jFZLmcx0dSuTa6dhvaNigTs3oXJaBWRrH
QAfdArRh2S4ktKsvzNaw+7XLOegwAojkwJ4Ddjhb5l58fbvYGLu8P9XPkPJs3zpS
qT4xKLZhnSXKl6q69d4zaPi7gGiScWmHN5w0gO1mvFonT1GvwDmlxeISN7a6V/2B
Tr7fQgD85omBbfTOO+x4FPDoVeL05gzBOY8Qi8N9EixMKlnGMuMoFZe0H+mbI07B
IPQOsTTIZ6pb1MnVYgKZmQVsUN//dcajv7bAlCvpHf00VC+5GYtFewhVFUJAxcwf
LXTzDblvMKAFFMy47lQz5qbSv0Nr4gDwd300RfWzAGfcl8ZfscqOo6pJAMa0Q3HJ
ENAK3nibCo7LoBca0Nz6l7ueyvgADuUI4srLiHFoXiw+ZKkNu0BjuNEduQ18cB/h
PdFLNyYhIzgcPgvhrTet9EgGcsZpfKY8s6DAYVd/KNnNrVMNxEg4C3SuLcQGZA/r
3c1h49AaED+6UbxfNXpZ2xdYjWoqNX9nHWjcs1XFurXQrkyHdKkiOB4L6yTHwtLT
la9+3/Dy5ybMcxTFX0ATR5Pe19Be7aOPEPwqvSJF7McMTk6PvJTpThhA+c+EZvh0
AGAi2i0AdJutFNHWuil/TK8pAWMSO9ne4qIiD5gHqFeMR1S5I42wpYFR/gD9UbXK
/z0kgdjl5cUz6c14FTPTk657Bt1Tqmyg186yzk6fBoKMTVYmjIrxTnJMT1XOyWlj
PTIfOHPKp09w9YqFcPuava1bMt66x5u1445qwWZLMI5j1y80jtmpaFeCIiPjvFnM
ekdpx2rMeAu7gdWgM6o+iCbgGsQ16G+SkRuILTKFMAp5UGWWA9WvdDuUb3qwJ5F0
r9trKMGHGmzl2lI6ZaQi/F9ODnRQgS4D6pKizB/r8klQtKu4bJeNlOEGRz3/1qmv
CzzgJPVxE528JVsa5O1RGSo+ivDWXGQMACIIyecumSJvgzLJMyvZahXpjkjCeySL
AafH6fwCTWNSwnF2VCzf8U6kaIO8sL8tKjVQmyl3mrnyBZS0HtffBUi7sv2Bb7uN
dwdhQk1r7bnh9KWyB0IDwtspvHV8Cifm9+F+KqxgG0HLwPWi9yOBaMUnJAgI38EM
FLTX8rGWWRJYXT9GG4tqj3wA3vlSaUFBmaGaSHgo9lexX+5UAMZ7gn/wU4TW9c2S
GWvsulljkyyo0YGEIbJ0KPYsrhVhOYVPog4Le0SmgoUOC2jfCcZoHiu3gvAd7HZB
DtI/yFso02GQ/aTJvxIMfaKxq0ohWk/4yon6OyzybxvrfX19polN2q4V71vvN/Nd
nrfNJNRQkhRL62z7ezLWvmkoMkUdLAnK71Freg8tFsExIOdjZNMt8gcg+bv78lQf
6MDtHBK7BT1jqB1G/R+I11QVHHctv2/7Dd2ZCscy01hbiMsKKBmwnU/L643xnf5i
JxbEce+fJxRruTCJq+Z68Dch0bahPI15yKZMzZbBQ/cZRV762TkHHIQxN2v8QBIU
1VG9ObrIt+hEs3bB++qcorVpcQGuGAuMvq6ObZKgGe0aEnL38yAFlAjzT0nV2b9Q
eMPDMKlAVH7ImrDZb/Z7OWKL+jbk3pw0WacoggREil59BNVOVtdHY+vMz9jgUD3e
n1Xdqrn12wqHShFfjkyIJjFtHb9/vsNyX9rNX03ETnwnwCd81JnmPZplNECO5XQe
mrUTgEywvDlt3136aXrhUdoQmm3EMiKybheMscMNneVjuk8LOKRU4G+Y+nmnmLLs
PQ6JiuIOcIKRVSktbs+QIBJwq6P4cBxU2jKLty0Tk4EJ88JhMNVLaREDvZqK+uzP
CXEdFXKe2CnCVFIFEm1eUqUxhoC0Jcab3srEdcKO4K4Fd0blPVLjozTmRA+sqr0L
xNDTnAfpPfAoOzVExjOZSAWnX4jjAbbZoeF0rlWMPcboT+PqS2HURUYmqpyv4Qbq
DFoTZgMiHpjJdS93gppUVYkFEdtOHGzlPBAMLFBeUSxL44t2g+4xhxSoyv0emnEe
soYF5Cca6k5KfOxmvrmuFl2mKPuDcLNR1+E010NdKQzHgWv1pmd+uBGM4x/LgfEy
5i9FU77REhsgkkPC6AxmkDFaw+qSb4H1IrXX0ny79gaFITrAjZmTGLdYO1vT2e1s
Vhzot+dJjPOQecBro7nlNjjecavEqrj63jTMj/Ro9H3xINpFEDWo2BR3ctfmQhV+
acAzA0Plf04h0ZVIuYzp0DttGV22yYy3eDcKtYMrdNNzPV0HzOhdxdCJUPiFFa6R
abfBRo7EWtSOqymY6um1+EZId8cXLKzlLfEJHvreoue4bGzN3JBXul69+gQV3gv6
n4QzE7JrYnug3BKOj4b6l0a+lXAfuMrJvlYh07A0tbrmYASKf50UpPtdfNX4fU+T
F6YfyfIA9i0Gp/pg3jtGgx45PHU8XBq3THft5Tp0rSjbEOEyKwEgtVRkL4uBWG2K
RW3OaUAjO4hLUNetXgvWWUQmgvQMfn1SDHLYkepvugD1QbFElI1DChWrezgxi8JP
IltwO+l2GwZ/ver8T0FuKa2an1XUkVQgM/RnRpYNUOglO6xpDwrkJvAiVy1CFjEv
LCaykdWC4iw0f56JyZbATaGJ6wRygaAGhWJcpaPArIXxZEqpSgeQUN0N74WSgCbZ
oAh/l+LEFosZxmuAB38bvCp/2prWSwkQGhfiHDitHYoasN7LFoS+ttoOyOCKmM5C
kdADVBXnPgmfBxXC0FgQqGPMWGMP5y7p9wvPGssXAK08EiX/TgEo5hgKBmPTrU71
z1kNtznWr4/nAVmJYP0x6UzhUIhBURMx/8r0C1P/+r50IdHWtliXXBGH+65czb9V
PbT1h9huL51NCHTmAVjt+3e+xgFhgXeDKBDPS8hZD03mJ8mCABZfsIGtxMSKXRux
+8+dEvIpcJb+S4/vxnE0WwRwI3a/gmG6Am8vzrMVjT8EJY2oSirtohgASWDQu989
HfpN87totvO76yHNMX8StVts+vV/te+VsurfwHHazXT2GengVmSdTF20xBeQStCs
6evef8kbgDZc6loNKGVeSSWBHEeoo5+zfcRJUkdd8JfRviYrv0tSfXdO2qfSOR5A
3YWrpRyA3g7imoC8s99IWqcv4rhX0aKte6ELUq0qDcn3p/ZuEKmBamxnFI6zGEsJ
aYv6qZAWtDRRn4u5eosN5u/VxIv/7FcD8zFK8fwYnvbmv2TGrMe2+X+OYpPxwCdo
uZKTDGBjpsqjdJhZrQ6GRco4ojGcOmqyO5QtQxceLOn86cJEfb60Wtxrx00VuZUo
bOaXZNe499Z/rKIrDWLT4dhw+nwy2hyu56nCMjv569IedACyVkazny0mn3nw51gf
y0WdxQR4JtWPQvzkc2cjMz737a4j+bgUKx3celvVEABv1Xq1uW+iszzYhzRpTNBM
SgTMZ4B+ScuPJCfeuPmUmwDW6Re7oULY5VxoRvpqRHAOEzS3O0CEzyFm+sWzNQSp
wdI22jVZTVk3X09H7xlSHsFvX43vCyX/Dqo6RAOVrxsdL6ITjNGH9OuQZIDw/BVv
/oqiRybLVswukvO4/Cxgj6qjed1jKOsepH+ztGlDfP/ZRbyRUxsWzlJIAjaCRcLR
dmZYPCMciPoBxr4zyz+IDa4+NWxZ8bsoCQsubJAnEBVrHju6YFmX0/yCD5jnKNx0
JaR2ZdwZ9XJkkFMDZULfybsclUTVJNsu/PJXl3UVPNsK1RiMrwbUMg5rRWkdOjuP
Js43IFH0PpLdMjZi8gXToUN8lvxnm84uKWhmwYp6fKwgpzy++z7kwN0xbcqo2e/a
RCY31kug4cgBh2WdyrhHD/tgVVwZzg7rxTOMoCQ7dKZJo+7Jx8JbxJcWsgzwpAdM
vdoEPHr6+okCPq7b8vUbuQYN1fBcLXEaCkbNXNmjd/0Ro/sYrlHbALIwO0kp8Frs
kQhopg94vCdBUbwdtQ4O05aek37oFxHBsrhMcs8qNDSMh2XbCk5LFOeZRawPj2yu
zZ3URc/HBQJ5nB9ALBdtiY60cj+ytZK5H5/Fx54Yoa8CPK7QBkIoEzFcfFmWZuCL
kUewwqpjajlfRjnfMWwiY6aJ+YUQ1j0Jv2Mn32vy+6LA0JoTPajV9fMRplAhyEBw
J8/ZKCjA1xpk0lC33r+4wAd5DJXu350wZVm3PgdX+4Z56R6glpGr8zci8feX9n54
cmzUorLtabFw+t73Qf3HTT1hBgpcJzEXSynMGZC8jCyGd8WUppwk3siGUF4bAQ49
LOSnO76RFkk7OMb2HQYIT1vaOj1KrX3Gb4S64hPZFWHhOorpg+qQzI3nJ8i4oJRY
YSrZruJpuPkByKm/Zv6Df7jaNpEycfsOcMYeTzgjtMH8RfRT20bXmFlnbUjeqqjV
clrqs60RWcaNVqhJFSJjfUmA5yo+etlyNrBIhNMbO2ma8peY+1imyN9fdDbBElVO
PTTQzAs8jfgc7niWIy4yB25rBI2Fe3X72VifSjPgeB0BwmkBZ9XQIXbIV18dONr9
fAu9x+RVQwF2jlnVEGNJs4qhyiCmCXluSS4QnPWguZzvEZru1xsj2qsmTyouaIol
Ol5geVRdWiliZ2rHBAGrkqW54Zo9PsSBYEK4kXxHVBd1kFvKMp+LTXcoeu/knvqm
5np1TwNhpvz6w91KP0xDWX+u5l//und5Mbon6IhWwYJukqm2sODy/0F4DxwMrnb1
ENZnBYpF3IGetzYK1lZdiBvCmgXW3JeXhTBR6e4brihK837c/STSY3jq1/M9xeD2
CIuYmpwkAjKfzwjTGpCNc49KiM58oy7LunGMaqrQS23mLPOopTH3K8bcv+dxiw3+
ZqE7Ux431fTbmR+DHuTBCSVjme4YtafzWpn25etVJ7IyXESKEIQa/06hMpfzz9V3
fSkJ7qGaxhxeaDkZSI/tB2BW3vRq4UpLWXBmGCjXSOJuZ+1bvA3OXwobpvG+Y1No
4dLMxaSYspc8yeBKr+opyKJ+T4mDI17yekWKZCEVqW0HnybRMdK5HbvfU5GkZiJU
HDqge9FvixkVVbrayPFX0A1IvmE//mFfXBphQDZZBCDWbSfadTqkzxPH/BMwyfSh
G6178G49m8zVlB/g+7wiAzGiP0zzgS0LY+4rwyPvOjkuHlFHsx9eq0yd5edkjVnd
j2iWwP7WD+54MWrcBkdr+xfj1oZts0FfFSr1ejW39kP+hdOuNx4tSUygBiwf5W3m
LBlINM6rHYF27hMIqrScz0RX8XSTmdTYj6xrJfTNvhUu/C0PeLGVYFvOGY3HXUbv
NOGkuxuKY/iT0GJYY9fbvrkvmp/6EreprSKJgcFOzcCWWL07vw6sjLA6Oe/tQXyw
4QWjOJMx8KpJcxFT+hNjwCJ9vNCIlCDGY1rUfN+OWz2FnBkPwkZ4gJb1cyVzGxji
QKu5sSfZePNqvJ2oP2Xs0rwS/0UL+KpG5Zj5R761kfJLeTlvJj9O6dg9OjjO8GHy
gyxEzAM0gRRxsVrFQZvhwTW/6LqRkJlU8GQrNhqnIH0bgTbtxqeVj/O3ls1BTbZW
yCr0uBRDoAzkVqmPzVaqYfeMV5/vBZ8/PWcaLudlzKxNMVk3sSqAiDqsY/MHqBs2
FeOpQR+ERCUMnPNKHhA2e5QGHKTjagcH25nW93tqGWpy9zhFMPgc0o76m4lCVezL
oL1214Hysm4STXSxmN2uSfpNNKlYM17F9KGa4BQ0UXkFR4b2Ad4uqx2gAZuCCkic
DpJsbIP9saKyMescKoeP4pPNWK9FsTZRqo/i/fOVh2Ai3GqzW81xK72tNChX3z25
vPn5+JEETlaAYkmlZWtbnHZj8Shxe9tkjmH5hTz73JXoOg9du77ehBcoXuFgs/QQ
GPPLldnFdQStHJJ0Kl5LZVElG0DGqu4wA7F6G4g093JojxMp9he4N05AX91M/5wY
E0fE0V6WI/CXpaS+2JbM/BEVPMFCzlEffQ6XyvOgFSqi1DCN/JUqACBIfnF3i4NN
39TsacQhk4vWLzRJLXzFkLn1WLBzmHt2zES+syACw0vTirMBmCUmTiD3SFJWyoEM
F4sTUu/AfkCggWTkRNXCZl0uM/oF91PvKwARpaqYucDuzrzgrTj7o6PwbqOtZc4e
+dB8Ykh10SkpJT0E+qKi7hdkqcrfOwoCQCvlAlaLFCSnmvl5m+ozmo+ev4TO76UI
8Y0Fdw+9tDutqtA143M2vCA1VYesdckY4Mk0tv2edVrUvidzMFCVRQHxwTiBwDTt
52ub4rYijfbHKKAN8PYatbZ9CjtQANZdYZOAA2xtTlgKTedXr4QXUz6/wNUV6KEw
5EZAR5sQzN7aBvi98nNg4pWGWX0wdfEjlxdmPGdUvx0s7hCB2S+jBpc4L6JWNLkl
At1tAkynJtlKcD2Jfw591QYmVRI0lUgmsPmdRbX3DfBgs19iiNwI8D3VpEOBs8x1
YyCBNLhZ4kbZo8dHHmG5WaVagPDrVc34o2QMo9z6V61n0EsqepkqsoLVwWbMCIT+
7pigW9YT0f1PWQtgfQsCdiQxIfgZmGZ1q1+PmXZY7e24mkTjky+uXZ0EIKkqAvO5
jgoAGRjMuP4qGK4+zo58pGpQ6ShEL3r+NXGXmC4TDhGV9v59XuvRFzbgwkiTTLaB
tWZaZvWq6oRQSPBsfsmASPv4PkSmIReTPI9V4QtuaZTKtbBNtWS0symYNW1wIj+1
xeATpEkVKgL2Jz7bbEXvZ9QTijFW048kb3Nop2hxMyNi3rtYrzP6ZoG34EE6QMlz
5pcBU75Y3fWxrIphXKNIoBeE7MY+2HrNvrOAVbvXXnqJWzU57prvAOqPPd1e9hfm
iD0oNsnbtxUpcebQlH7yCAlHOfZ1c45NDx0MiDlpRc9rHI6LkObOM9OUaq20Fxm7
g+0X2Wi6Se+LMGoIgLq63VlRN65Qd5tf0EKuRqYhmJqHQHG4kf4cUiIeIpSBJCLK
lf8WzO89NTzMpxAIGOjTaHhPrUc+7guFTEnHO1Mf5VVaUXH7+x0JZQfUotY583FY
hp+9vDMln6KQZv2vHYO1lzNvmLdARtUpEh+IpkDfUemcxz/tiyMLgnQctbT8DwHg
bsza30O621Eh2oxlXtDWYa5mZ+ieNvuS87IedA6ePI2AbodW1y6zOsgd1DrLPu2O
1xOdcINo+JwADy6k5iLqDZhtX0mL5sEilAi8eAI0Oj4sm9ZayI+bHBYzbqP5B7eb
eSvlxlc3O/HbSxQfmPC16q9zbMsW83nwGIZddiHvuuxIF/S6DtjGESk0HvWU9gza
K/y9pbNvF3vCjl7AlnNXXQoypGLOVzt7ZVM1KbSlqkuaH1lolE6ZMBm3sAqT+zsS
zrRb8g0TX5BYPDiXkCpU84i2RW1xbGRUPIP/KfTmDMzk+fHNlBzt3Yi2/EmPkuDe
8JA62D99Uql0QpsTLK+ljJqPQxwDjQbdubc2YxZtSez1GGNsYtvsSBYISK9bwzL9
ZFBHio7jFO81aIQWQBq2zuqVn9Y8CO+6R4iFqWGzUUnnR8AUW0XX9RSiOAC8+1bN
hMG5z3gcCCIHaI9TfXq9vfAyM1YTpIA4w3C5UGnEFfBv2FR/5KilbIbVVoirMYtE
+Zxhcdf5uzbjD0H1appbqmKicocfk/6NKAtsBBG/syGztwR33KsBRHltflCVvPNw
BOg+k2tKLChEdP2fjOx0IEnGT98dUG/hsMU0Y5pnf7GAHCGxkb0LnEJ8ZwmYx2tR
fx8IB2YhIWU7Aqd8LFfqvldC6l65xRpJQsa74fL0PW6X42a882Y93AZlO9RxkrCu
7bOfh09tTA3Fi5Dl+JpKpryZcyI6UF5/D12h2tlMQXINdZRaFj06X9/5iB+sFKPY
E7kFY7YHQRc1Do9RGUb8fUE3fNu5HSP6ekuq6gjIt8xND17LH6/tMBqii1UYzRuX
+AqSwU/UljvbQhHjQpJkyEEKAHEBA7hk6U+WIeZs8rJ4fDc7U50bsVxGS4Octj7g
q3Fnkm1didg7+0rVZc51X/9JH/SMdWqYFGy8/c77FW0zXh2UjZ0KtUl/7yJCfBJO
uRorjzAmsBPZj12ysgb1Oc551E15PpQdh51z1p87jcifktTc9uuOGf6QsUvrp82k
bxlCuYxyaroYT5VXlFBlFH6kQRjC/LWWzNpYbMHMBXfd8V8C2FDxrjoaKWRomkUN
obtoIdVhoF+UP9+pj18lMUuDo9JauiLIYmm6lCSVbg3DmLaS1Dk4gD0SW7HJH1EP
aCXcM2tApBj1fAHYQ8Dyl5vqQW/1Q3m7lz7povd1qqqJRjJcdv+fI04ZMVGAIF7E
+62Nucgb2rGltRLcoERWbplrCFecbPgwq+Me+70tyVTSPcZcPQ0lK3eERkLpzYxU
pNbZ7oh3vmcs4vwvzqQ6AK2bKuor4DLsdHUqT5RHR9PZ4NHss9yi1fYYURzqrPRD
7XGfIHt2dWi1MjNn0UWJiBWDtqaEcsdXNZJS0imxo/esSzYpbxxXt8vnK3dKNshG
lQiC2RZycEQWX+oPtyldSJ7KlwqXAWr3LrUjQVU55a3HzGd3UEZxHxYx/2raM87N
kDfnyzsXsqwd0eXQIKx17q3L4TC509W1Abfn7MeQY53Fg9Ofy3K9l8lVI0aT1UsR
C76OMF+phkLzavBqmcrGr+xwF5jJTF+YNQZf5ng3kHTnWmsaPB2WO+sePMA9Q82E
L48skLJn6v1rXTbSNCOGAKDLCwPBOtI77FSZGYOTWrBk8JLVpqoz9m8TDo3Qa2mH
w9cUtQ9Wt8HHkIapWCz6NApu+CmDPlEqFEjy9MO8QY9o9s+Xmyjr6bYX2heWvsAM
rjcM84r8yrkQWqEvgMqWA1Y5MM2WmO+OABTFqZ9+0U3jqXdZBs9sbPWyTU7k3xZ+
2HBpMvpSBMHN4aul/qfQYjHi1dZQg/70CTOrhrftxnstmBUZFeGE4t7DSpRuSEo+
XQHDjIAQoIaTp3RXU7eYrXKdiD2DJ/DRonltwNG5PJeuUUvccPorudr6mnN7v4V0
rMymKxd5NlxD5n4WuP6A063vGbySnIC1UOX7V/jUBmM7qEceaV7qCylXzKPCGHeg
JadjEEmGTBdrr2Stn87x0r3TGWO7a7f38MuxNnkAOsKdPFKUmXye3RaCH0pAn/sg
ikhroV9L/akx7khlEds5syB5Zayy/OTvN8BtEsRyXaapy8BYvWyBwWMsTrpMe5Ty
9Leu9l4YiKoFLZjr05369ZbudFyTvwJ6iIuGr6oXBq4h776bmSMSwdRabz2RpN3n
RMR0+7kMwWuRrjxO0QBMTtu1xuaJ7MrRhNyaYqHDxuxz/5Iv/KLKJFRoflSOjWEG
5qa2qWnE3Vuvk6ViOhmw16zhgGP6D+Nr3UjCb4uXUU0Gk3Wbdfj0VAe6XHdWcuB6
EGFEy070y627njA6Icij4iLY756T0ESNpHynoWZQU2ZSvcAKT0q3bRGDc+GCLxBN
dpCLHgIJp+id4O2E90mBwqEQVx9ENNPKBSi0bMK2tJqKdvZIqNMwSoIVrX+2e0zB
HFe4CAdpVsHtFjaIj/lPt3lEXo8bP6eYP8h/NS318XiW4WS6+DsRdxTG/H6DTQWf
kUmC99spsjaSo2YURtCp0RW1FiNOUZIG4NvQHyZD7ZwTkZD9dedr96eIJipuGVIn
vXxtuoDvlUkCON7i2mNLk7te1hJyfypjUEphDG5rtIG41GErwsYZVuzkzyU1xfzK
QCGDAWQhm7sIBqsVaSzk6IJ9rdH4dOUDMaRNx7idY1wmHQJAcXPAU+WzcV6wpKaH
2mYKoyPCfOGPTZBwW33+8LRjtH/X3495NYSrpn7Pf2xJWrS2lIidOniyv+ge0w2y
E0PASKoBRRCr1pZnj7BWOGbw6NYI+7jbv/yYLo2lmoz3w7fCVOgnnPZGT1K9ymr+
3ravsQDAkc36Y+T9FGW0pyU9G+FIoMDFvxuUXedXGT+g7atlFt7u5CTNTVG7N/xD
Me3b5OdwvxFuF/Kk0Ked7HRpUGs3Mvatsed+mrIwZAWvXfbgrMl8ElahHc7Adewq
X13ctMXf4IzUOCSEwO2ezxlt0I+0qXPo4OLlQw/LcN6yhlZ9irFg0L+ZaT3KMnx7
BZ2NsSlfsP/c2ajSuxJw+y45A03gXabE01lQ0O1/hPsHoPyua5yua2etX/LAaJIp
dEfdEY2VgwSDUz/JwUPml39B3PN1LFzcFvhQNOJBliyR8ezSIGiAZWo1UBMVmZtM
typK2hRK0AfWoXp6779Eh6yKAoaHBEIP94aWHZpocoSceL7htRz/HySboGr0SUOa
Ka8B9pHuByE6dtjzKSW4MJVAB61j0bS8m6b5LGh7J5MMOSoKwc6GAeYzuK91oJ5P
tsQ3gYtNQdWe4kBMbPoVnNHhUz2vwLFQqH+phG8y+ejeVBL37LLWcU9UbbeZ5GzS
ib/pDk3tLzrcIIUOPA78myxfF6ZyLN0dPdqSJDQSnhxWQj2FFWQiavKQorYvLMin
H2CkDuYctJRsBz3o/JWmxqI1hioJEWei/F67D0uAF2jfuX51pM49XcrDFTlCvow0
i1lr+UsTJ9fmD5YqYU15CSqxz/YlAMlcYWUpuYNB357KZ9hbkuWW2X0VZGL7IeJ3
XyTF50krk0Yt2Zh0mllJ7Mu2MpvJqee4vmk8DsyW/vJWuZIOB+Q4uagGE+9Cjc98
Rhlp7FvmX2ThxVb7k1WucaPh+7Z2Qsce2UPPjqO9O33LAiT13PCZuB20Xzn6+/RQ
Uh5Bq2DTlqVCtqgMpipiOeh4Puso/3lUhzIgfAstGk4C8qyDjZ2JkBVPUwOIHzZa
K3Tg3W62WQqc1Aq0s7/TnyTSxjHX9pYGzILIT072bQbFE4pSavKJ5KO8YZV8s0py
wAnRis4/AvvTtsRYbNhucKrwHV0S17WJiDTSdWuB3xI7EvIbuWR1Vg1+LSQO6TbV
QX8DslJiKoH8W8DrLWgTu+8rCyergt1a6v2aS6I0Asjjn5ZDhjzlyhmrq5xp8keG
G/RqLuPBKoedEbDma2U1Nd3kDvWIaaBz+sSVkTQUrHkBIKZKOL/IjLlSqGH0Svk4
4OUAMyUURWxkz2vRoQO6iTWsXeitieoJmDOyLlJh/Y/y2uy243yf9iTFfFgW486s
HA3aAXGs5guUdZgioJZgxgvuYTiGwIuU/ra9j/xUL+OoUQ5wxklviC14/kZkWdkw
090i/tBkrPLCM8TS/+HUCb/4w/8Ci+Ic/tCzttdf+rYRR2FO5ALYMdYt8BdA2MOm
yIksAwZXAsKDGCCMTXrolJSN0SKGOiAIWLRwO+Ydv7zMP9A4dzv5Y97s9f0UCJqX
t681kUrGmmQciLLvyqkP3n70c898VpFbJfhPnY0Wc3hUggBVpf1B7SHtl/QTBleu
I7DgtpIoFbj5KpoEa3jJ1BqboVESjIKkBAj3cKGlpZO+9QCEVri4ETvos0hxHkq0
7WfUo/F5py06OO2bTqgAZ4yudtjwP/Ofe3c4RKYzgKgCraJQnxs1CjyxVHAz7msG
v0ChyKFrCXX3lCPWKDhoK3Ad0aCbhmQgOSmqqsytRfga0muCGGsBYt5EIXtetVu7
dTpIuZalqx57r0PY7GXfe/6HtMrg9vCsphHDxY5tJheDNDp/+W5t8PmAHm9vdwss
hSMnb7QxNeeo+MLVDd7Lr7L+2hPQz576Q9w1D7f0lLvyum5sKMCU+D+B5FW6xqcJ
vvnc8rMPBbySzjL1XxkbNnNRjkybOzWHB+5nocAJBKJ80igpRFKM1+pyBLE+W8rC
YljcxJUqDVJbriWkCNBBJ4mEN/ROFq/rj0IkizDSl0u1TtMcJCItbcR+6UQLHX6w
Devn+H1jT0Ry4+eIIb1vgJslZSU0tlqUD+9aBw7GIIbxls68WWn15ePKYcZXIIEa
PKPBYULhdNQApnLecYmk645bg0uAMFhn+u6Y+fJvmt5a1yeOw69hevapR9h7pBJw
yGvY+2dpr7Qx+EOk/IdrVo128w8VZzywJ68HQWHVjtQw1Fd9Uxn/nIcczz3cM/Aj
fEHPyS2d5r6EooLzKD+cdJzycE715FYbow3Oh+Dm+QvX+kTC9dQVp8MDeF16Hpzr
50fiW3oc7Y5xB3s9IhPcJv+nsd3jEuYMMASYLFZI8cV6yYLPgN8eMHGADT9wlLiI
lTQ+avNfNlX0bdhmvpbjM5plLnJfmEP6mOGNDXV4rgS75I4rvijNf8CzoCGw6kq2
vNhSdBTE5pHlcEmVeaRp5xGlCcplWY/db+12EW9w6jJk3wOk3EdadIHU9ikDuovH
0lsUU8//ILI5bxZM8HIy0Lo3PJFqBsCYA+P2eJ826MTpkTZP3vzv+xIsChPdsy59
j61jHLVQJ6k4PyAcn5Ba05kWizVH9vdh5/wTAHT8xIJXmiN+IO/qr7fCguz/5eUg
oIJmOzfR+WIgLpWfHhFXR4yjw+EDO1LZ/AYTNSezBsoHXpxtgFpBE3igHWPmLjZZ
b3rKD0UIVAqNr2aHrT3yx4O2NyXYPnn3IATgiGNAIKXBllNMB2ZAGIG0rFWSE7Pq
YDxd4Owt3tUCwTLizE1ib58Jf423vXss3W+RceylUJ/AqJ7T4RtGxgmF0ylLzZZb
oLwiqaELHZ1kspRKG9SAnDHEG/mgBbMkJlszIqafl8PKvmisytLWTybQPUAlRqzR
lWz4dwcrrCZnoM2KL5EJ1xnoNJm89zxIhiMSHTWC5huBj35h3Zn3LAD7mlRgFJWr
4nqK/3aq/7vAMTsTFEUr4FEdz+XTU3Y9ugsKCtScfUrJ5lVPVKVz542kj9hZ5noj
37Kbahg36QCRqX8psIW5iNG7Vjn5nTpiXh+Yo0wFa83ZFP8Cjm70AKcHO06zvO0g
XPq6ZHWGKpowjIn4faKltqc0jHJcZPqyFoMJaECwI1AAns083EfBWs1KFdk43JYH
pJsTUU1oj617HhJxku1ZNzK54EokM4THLou3yl3rhQwduMegh9IzC0lLBub/1+d5
U0Rj8qca4zEKUARkbujn2ldu2ZwlACSHA2AcV5mvZbPBGYeep5adLPK8XVBiLwxF
2ep/Q3uvn76Gnl5fDKjEhOB8WWJOTo+fLyOz7T2fIH3cJMnfj0HuJEAdWuMaoDre
pz0di2H0e10MB0rTRlxOWD212eNYZFf9HL6G/SB0ZBu0QVsu7tgGpQ8QVZKCf/Al
wM54eYrME9sC9Be1QVwcojuYRhWT/b24f3wmmgtkDfyK2dVt5YUvPwPJVhxO57EJ
HoP7lSZn4TWtmzxxybaVRVX1tvYnBXBbKPUa9dWKl3+QdIIIQHOO5NvCb+xJSsPj
X4JWesGXYflBL1yHmw0YJhismUkOjzuyh02PKYbuNlHC5aLHtEbJLuUrJmQRU7cu
w3ksOgYRb/CzmwhGNpoafGzjhL6qQvqqX9zpvsRncj+dEc28Riv6nJSYmShLgRFr
90Uh6VFYM/gBOjc0GpWJMYEmsTtnue7QaeHFjQIVCYTCWqnch8OHc9FZQlZQ+Y70
1o8SyiAsVmcPMIg4h3ya+o4yVBxCZ6vVdflkaAG0SbJv4MMZgAJSO+QRlIGNR9mm
VBTA8grFBp1Ze0tsrobPH7sb+wlXUVAh5QWZexbE8yPpeQj20U8Mds7ZbCYDt08u
A2YzOi8iunvRSyxJyAcOaZ/oP5QpAwsmD5eB5rR4vO2Y3L7WIEUv2Uh/JJYUigS9
9fySCcb8GiWC0/Se58C/x3FZWEH9Uw5626/bY2ONH1wpQKne4sEXAT60B6TfL7N7
3/c7x0JHHqUDDDz4/VEERoct/yMntn4gIAHAlLalhzL7YM5/VNH0caiqosUMOfy7
SkcJBkDPrlg8oyHefOcXinZywLm20LTbFIQW5IvlV0ycj9M3j8h+2Z+E4nipyhR/
LQCnA0SnG+o3hJqDA3qBYwsZigRZXH4SRaAuZRxFKSK/hUjGn3xtdXUJUjvMoxKw
oMT4AJr55zC9rJxpU5EY33ZTl++T5pkUIx+JbR99j2MgHbEDbnjpZSxiFO4yGBe9
w3c7+WGXfSxUTE7/Exnrn7LqiFSO75lXJ5DKZQEAk6AuQVLPz23fNpUvb5oJugkM
zSg0OxnGfr8OXLj/WkEvpdfoX3OtCPBIYH3Dg/sbr1GVgBWz1p2Ieym4Dt7T3tSS
5TP3ZaThWWEXb4wvLMKR1FfvlUgdzXSBNHRJjanmgCe60HUMV9UVQHdsGP1h4VpK
EAMxAhw4Bqjoq5lpdTbXVDVSCz3YqJlkVe7Rk/5PDlLEPQ790CJ919Vo4aMRsnWe
sfmVanlCfpdt05zANmAGebtaMf8M4pplZ3eBmzlW1Xuk6uQ4Bc0ofqm76NkvUrWz
0v1McWVTK3nC6UdIrUEHEOGk5oL8eUPzeGNuKZrzdeyM5gP4xDulLatKZ1UV6Sw3
uDy1jDgOQj0efZxoBNtSRNR+lafBU04xU9cP57Z2bPerjVz85RLXARgLR6DqQCLA
7m8DvHKLh/a8Ga45Dm9VeE1lmbmVgvNEdEyJquWmCAj3TK22AYiY1jm3GxBFZOpy
5US5h5hiU5pCo3lGrCwWJDlLDUnDThrPiynoenDEE2HzJqbvNgeVC/zTMDzKWCcg
1oN53JwhINMWV440/5qILDuz0eboVL7GKcE8YCu5235cOuapOh1MemGSH5cRRty5
1LtqeitV0MxQNfyIiSWmWnOkFX3saAJbFgV3L9BBYR6uaYCTN5TGeuhS/g+na01e
xBdePpS5p1ivd21f3tOC8tUASlvqWUwYPZwgpz3hC4JD780BZf6zaS5d8Mz1j66m
xpolSRUeIxCznwYE1nO6keNjUeV9mTMzcoK2TF5WDQXsvoL6n3gROqL0/VOfP5o+
Xcvtx5Iw6Rr669YArLO0vnLtW/iFf3fAIMq5k7IRFMIhHFP6zfrmvp8IH2ILVKq9
ZSSvHc12gmWNstYsdw6omtKp3uYaqkKqBsHAC2ygdO7MbtvX1ztCRrFYOc28CVkY
1tuzTxJwOwip05YGF+gFJd6h8fQhlTei6Fdk3lkj1YdLLKaNdvIAUV8Gd55DzRdW
URj2lSskXwE1szS4GRJVAhgXxOeoCOLVXUrJiM9kqbF4KoEEt6XX4wPBMujPnB5E
7GbANj2qxAUErxCXfNcIanumrMi0ulgtgnblXpHweRnYmIOEk5BEgJBODZHxCDbS
8GSCuLHgcWvx9EXtgN8+r7LDsWX9zlCeavvAw/pgeY4pyhJTAWSYCcC6NGxbrkoF
KcwyfZa6Br0KN9njl81Iy2a8CK0zTDt6W5yIN8/swYXCmN8viIkWsSa9uLYdYS1A
3T3bQtUJxDb3HOqP44ksqxdR1SXRylDddVmhOWV4M4IrjDWiHUXL5i/KaAvPs4qz
LYstngJdngQP8T4A+m3v6CUhUiQ2bBkVT00QvfCL1zqRqDpI2JcRNkd6o16IMqHa
AX1dQKggvbLdnepLk75eEezx2z5R6nNrAOllN+HBiQFGcm0C/eKFDhxG8S6Kyjdl
C2k7prz85mvhYKYqkm7Zfk1RMG5moNVDZRrhgt2gR6YEf3l02X9Jc6vDVsTDBGFB
YHLQ83VJlNqmz04InYX9plWsUmyP3RZy8VlwZhkF9oF2jS/T/Nod3NYK3tTSbJyK
2XXQRMoBRjjVOq4HsS0JdTxuhGiynPUb+tRpfST1gk+kjmvZM1MsFdrKOa6W4n8x
j7EVUVxuVXsPPJ9UJa/wUFPfEK5qgOuymoJT9buPaKS7gjb3Hzg1137hOlHtc2kd
VdKYKswXRW0Ftec4GouW/q+B7NDl8PGAz0EiJf5g/eQC6sHwWhPZ00IbHb3CEm8d
KuRUlAJKwn693ZTekpK5CdlyuO8KDUpnS9JjzC5Uc/ayBKwfu7g4OYPX3QvGAz79
OJ13DQw7mLkn0d+j3+gQu5YFOOfaTb7ux0laI5urfAIHzBKF3OTM/kd9FqatyxzT
OILOHSxVUEHiRQqet2nyRJjeoF2vaMsIEE0ZFqCzft3xC43vx3Ff6DJdlY4mj1cy
z7xnvtnCl9JtqGXzgLP7nWoGh6toG5v42uLBdmsWvJ7HwTT8i6KDdgUu6GThXcd7
I1zubyiIiI5xe6dOVuN+dsXrMcUWIFYhGgg+6YHtmFnp6RUPpy+5pCfzroB1dVzR
I0BYD6hZN7u3Ob/siGBdjpcITYRGwoxPGPopRePkRnWQ+bjNwpwVu5/0FqfRnl9U
dNAsFI0T+uYU/mmYo9WMf91aSmoPxZ1ZmY8E1psG/92EJmuaTQVSL6JxDc+M+Sxk
Qho0/Cr5AHbihYwy3D+eAdBqZ9cFKl1uMELASV6bM+LfVhyCzC+mJA5WGCDWY983
OSfW5bLGzE/u+tiLQvNgAiHy/T/ZWPzDoowMdssgq6nvveQyJ1LCMhtUmVYFRvCr
3h24iF9uUGarBTCMS5IuO9vPs2YyL89A//pcom6UH6fQv43y5q7gUyCcfBcWe4Wf
0tFt8UWagPeWtv94xNh92Em1hv+AbPH3esBWy8ZF73d40AYZD8aVkoQFmV1Dt5Jn
mcf6/RQju4fKTj98mGaOyPYPt7alP+0mH9NOZ9bkocFiooZCVBjSKVkBtcPszEOQ
99gnnmAiWxdG7iBaRylHARR9z35d/j646Eg7A6LMjpiGP10UUELg9JlnI0aRUMxX
uwf84eJKezV+Sj+eOyai6xmPAf21mEEAECccdM2HeKdeB8wZP0x5mBIVXRwcBdN6
bsKq9Gjiq2AjqR7F2ZQOB5fgbFHEmGA57yAjpM4GtAloluvGz3tIbzmgQS9GVqlD
ZRUUOsZSAhDU8zHGBIA6QiFitoC6NvySGZsuzqOzwMmtTAey7yJSPoNV9pqr9Q5o
FzGt7ewsi1W3UcYD4wiKhJ7Oi5mFEGIMUGycBzQY7mkQ2m1gVhLwpeltsBwEHBvI
+narVYvwRaLcAmOP1VLCIOZKYNcru21/UW+Tm7gRxg5tjsfKywffHR1xtxugQ+6W
v+covOK2Z7yJ3Q85bs+q7VYCh3T5aK2JEj6YjZn9x/UfOqMcPMjlPKGw8mphZ7qj
qspFBNSlps5RUYzZ9MCCkPQu6qxza5NXMvq8HZ6NEDktfSOr2X/0JrscMPOwIiAa
tOB6eSSIX4CZYmevRrydoBPRPwBl965dRRVQnViEMJJXsMBmDVAdI8TC+Ege8z+P
/f+5FE3gmWCouvtPs8QDaM86vqCka0OVTIxjtqBXTbCnxv7ZJ76afCtBQBGqLg5q
fr+EvVVSBBl8vHrdN6sZn7A+tI5s6HsDOsRaPu4KN+WqdYg35ilKKQBOwuTfpKoI
yRjsmsGYDXlBJou4MwtRqE8OM+4H7u/GZjRxB3fFOUqkFnJi1YjFQFlh4NF+9PuK
Ph0IDl5J06FlTejqVCLE6oAXYqJbQU5Tvy8CILOalGaVKTunSgtokwvjd12ejD4y
9sOnPm1YmL+ZyA0C44xAqKVsQbQvmqkkQCtiHINrbrZDTnd0AaFS6ZnuSbkahTwh
B5T7zsH3oCIZ592jXnBYKH87zJ00j+AR0OTzaEY9W0Dtn44GHT3+dApri7tbgBhs
wO8UmvKe/qcMNVUVywCDgL5JFJZE80vTTzx34wVfjfJN5BLzwarGZnFQSxl2rQim
YFnSsrPtQKIxmDv0OEhuMawK313XVjeBYhEibpAxEImkk3JBELtsJXA0cwZ9hXzS
lHE+6wQlGFq0YzTstQqlxNF4tNmxdAaZQYSlaM20EMEHjFW7vh9vY1GjxwKI92X/
xfHuOnWRPcTHqpVNtLD+7PJnttY9upF8CFFhhWR8/oL2MIcE1d5jyEsn7nAyfWYO
6nlxt9QU5f7sR88rX0PcIQBBPIN29pmiEX01Q869EVVBI1xOj5S+Eq7yCCRRDSKl
UjVnXojp1kHWw2pJ4UCVGTjUKqfhpUGaspRtWMeCyCdno/LO9soPUMDx8mYz/cmt
M3Rz1dqgnK9vDaTatn4nEKoP+tDW3DeM5qQffZ3+IazmgfWi2znRZNwfiOTpJ2sD
NdU2LZX91bE6WTxifYA+gUaFm0CipSEbRnhw36g+BWoo8nZFejzlK2dIXH9FWdh6
NrDuSxf+X0hOSgupjKOlAJ2K9YPDxb1T441FUphrMQneEPmKYoT7RCZQagzsX5mK
ZID2JwqVT8yExenXjCJyMcBb8kox8zDBleg0woxIxCx0nCHAXkYejK/5YauXZnJb
uIR8FuAgJO5UlrbmVwWf1nuy0F7kWyOaNCpOoM8xGmM47wGL/0aWPqoO4GgxiJxT
XhTY1ADCHquo1qDKGFd1P7Ndoojx3nqpN6fHICDs7ip7BOK572Wt6QNF4R9FIiLb
WC3ejXmZB188SIcH5mA+Y0udDeyN50uXmhF7GXU7Mt/b8wfNPkr+3AU2CHLjf2Wc
PHCZ28tke7sLZ/SQx9WrhmMUFAYx3eppYosaGp9bzok7Rf8RFm/ZfD1WXIp/7hIo
03+Of0WX39ZmrH4jxTnn5MFPi4obSKYR4/cHfo4h2diDw2JjESCCxWYFSU3GDwnK
8Dwra6ITK5EtUttLixvyFTjgGKHsrDP35Gjeqh4wMizFeLHc+L6EqKzjkqlsUWwt
Z21F/KPeVYf7k5ZIq8Nd4Fg43Dcwa/KKwMvZtWSri4HCPrDEGN2MOUyjieQzfngY
DSFaZCmmJQDrgPAn05ML2VcZSiMvXN2gawclHrWkLS5yc5BgJvR0POkxMg1kMpyX
kmx7G1dGVLmmSOoVpeevl76iqPchKzJySwbCtFtEjFX0UvSc5mK+61vNteYIPoRA
GnJsfaqGVe1Ao9vDnYhZPz0Q80WB7FOyUzswwo3Rc38y1vcbPIZc/bkWRNu0aAXA
ju1CY7cFqlOrVJ8aRu4/r8tVTijHnYedoWUN9LbGtmulc5P+iYdZJzy0RctqJZhO
qa1+ikCoGVD4udeWxVsbmLmEFnoAv7p8mlF6/6BGBevLuiYf3bIqFzFx5QsgpKSf
SFwhM80WaNfVUqNNxa50hZeVAD5E7PmeMCgB/X18D5lDMXOObrGQ+a8Hwjr6ZJb/
KCXxMYyXQ+DoGdDQJmC/8frtxOO3VMH0NNpWQyvIQEyrwkgmhJQhppWlRCSTdX8h
TbQYFOrD0kLibTGs+ktX8mQO34/4eKY/VBuRJvD5R7kV3mnhIXD0mRwV/9BSzBst
83hNn0sD61yCyKbQzbby5G0VumxViyGoHy/LoyUFNA5QONa8sHNZ9HkWNizG4pz3
1lIq9iy3MI5QLQTE1gSLU4z91gWYLlSdSJg8/Sw3t2XhGNQlhWZQgCaFPAJx/WZ7
Xgmw+zlxaGB13S7B22YdavYRgRqzyL3plv9E7/6FfJ/0FN7s4bi3cDmKYfN/6uOY
K04dQF4qqfmEHz6SPun6JdtadOEA7Xj7Dt4Hu491j7fvKckgA4XcZDcQ5u/kQDoJ
cPbFlllEgHTBm30VXVSbffUMoftbIRBadbtyRQ0nobKCISqEjf39Vy2cvIUMOYQJ
ngMroPzQ9z8p8sG5+dMM1X18tdo3umIRpLH4CTvih3ySsyZJVII/fmBkRvfqQ/7/
PXX6L8H1r57tGrcVCU2i47PSgL5zvORMKArzM738nsxcA3NBpcl2Rk7uovKWgdQ3
Gt6kIE1kTfbcAXgLLj3/QmIdo2QWR2FDoLPofXgcrBu4xP+rG+XLG9PK6cX/39rZ
4Xhqy62aJJA3/WhXbQVsRPFPkpjbkpU/hk0I7K2Q9uVwPUhhD1IZsCubkJpojpxr
jfSpJV4bXSJAi4R5pzV8neF+lWI4krZnwa0X+RDeDvi0CoH4cbaVBhqwbjfAlNK7
vv02nt8HNSHXfarT/79z9qLAdjwUQtOtkAWJ0ULGCeXMacYHbG1DZRILec9mH/TD
odhYZXiBkbtXoOGZKJ1KHQNWCSeT1BJkLQ+OzsK3H+Yj/4legH6D9nANKE3rbicq
NGkT7k+hSdgKH1MbtemQg8jgW4ZUOtYRwWUINPbPyQLlRIR+EeRyrnIQqS9s89aF
ZQv0uUjxNdvAje6Hp/ohreobuUEB+3UwYJcERp1HBHIquzuvdAlLEXyHccSi+TjT
riTZjDtRdVVvjbjxZy87LT4X650tGBZyapZ/pCnlNpzuVZIugJUTrasW08V1dD9M
mhFIF16lAo8WIDwWnVWTVhXSl2k5G3KAccKntu/ALUsdJVc2+lGyJrJMhELtnCHA
3ogp5Znvq0eHct4VtcKnNbNilpX+fdUjBEnKZUjwPccklETJu6gyH+nob8MUKuCD
R7OcY4vbxxcH3S1hn77Z1wKYaulclsq70EcVpi0RLACC0vvmqfbebqVcROEyo00h
h/hlc+Z1moKBk//BB8wIB3KFpS0fNnQhYegH68PHa+9gJcLxQKIj1mqLP71o/6My
n7h+Qzm05JENSVCZDhuc6mWWr1fHzDG408XCBCq8Ky9zFVaS2wnbqmDuN8KRlt1T
cliZY6IE9GzwVEZC4qh0KT7selfWHGvuGGPqpsamuCImgyZ0A51NFHIHupBTFTT+
Y1rVpT2oWD5GmMT1hgIAB46j6HZ0YurP4rUod1g/RdFQP7bclDRCyBgsVZITUwtU
ZMXPVQbgiCsBUKJE6ysz/4evEZKs0kuGTehQK2mXs1TGt7oHJunaX2asJK5NQzuZ
3scpe9HmRq1WXsMiD7HNnpibKZOKEOTbwLvy0fXEntvL8bjGWBgVzBt/S4zdtJ2i
8AywPbXAelbQWTxNcVtLGjf/qWTT+Kaw9woWPDf2vyLMZT3EkTRTtGS7IyED7Xq0
geNoZabuL7Pv/0BZ8e+HW1ib7UTHdeAFJgVlYEgYx/1M2bGpGynLIYadGzRs5UzR
nj81uoSgg4RgYiHKs5jnPX/SFDyf8Rav5ugswwQzXbAQN+FuHdPDg4l5nRchTUKd
69lFJyBMQU8o93j8AiK6k2K8VGBOCBU1D23/kWtQwDNUrFDvhwkbRo/HK+3sLEZK
o3DHwWqz2ITjtQoCZnqC/d9W6Lp+DLzvTIgN2cDs1j32hklDKoESGUP8sANQuG2B
nU8WpHeMa0oWR0b2bW9e9s84CEGYhRAsGuqgZAcogkY26IG6L2TAkNAnvl6jYyCR
7lt7qazNBcHfF+AmRv4tBWC4f8xZSOkmxoZLqsah7oJ5sLxoN4LJKhC7/gOg8r8Z
8MOwPH8me3Le81lFB8fYaQ+w/Af53rEBJa7XJ5eakMgqL4UF3UUZ3iiqdXXOjZv3
mRr3veP41eluSwm0lwf+pHby/VNujMEKqFb+eYdS5JlBg9blicYEYRxU4bGU6ozE
HIkDgNsongNjESB7hblXssA2cjSzUGF1jT0+s8HDrnkMj+m6HhCwuiXGooxdhZWX
+29fJE+ro1MbYp5ByJ/TZaQGgY5I5VbytaAxnyroz+4UQceTzwTERTGQFqNFy06x
jGDG5wisHzDRaHRPteRHDgvONEcT4C1NA7u7B0sx0EEUPe9zl3kubXGYMY5d6X8L
rNhPORq3nwoe5dkPAhhSSCPgsmNik+b+iYU17mp/mwBhLBmSdtY1728eAQ/DxTiS
WSRh0LjRAaJxhOIBTtmd1boCEwfnyfU0hN4EeEX8fKxTNRfgNcM01+rd51DhFEMk
GSjukcLDLWbDPLNM0GdZTtdj3OOAf5+Guu8TPLa1WASsk9xBVsVE5IbVtsmlRv6J
PZJhV0Gj+AAhUdU1r5rYUBOtoLiYjDs4r5ZZNQwaYEbH8rEWLiN+gGZPvxp1B5Lg
J3PC+wceitnONWD1TcpJdHKva+XOVaufjRPdD2u6o6LruXO5oDmolkrgd3lA3sDN
Z1sQLsUFrQikFBcOrb8mO9hy9PG+KbH7Fz8RulkSSBluiUNt4YASmFrOV7wYEsE2
3ujP26icRqdSCmdT7mPLhAtejyk5Drj8owLePLpIposHlGjMSVpW29JGeUkgqRPX
dZeVfQ3YCXlLdr7nJYnbGoQ4R/dPdc9rfcTjsLOzApPH/ulQE47qVgEZNrfcdYyu
0jddTkNQovd4CQqhylQoE4z/yxcfWeHM4ycqeZEbQAxvFGFi9k3DQuAYd7frD0W1
RLlqqdEBoTtikOh3HGOh40pNWN28EwIhiry2SIId86QavIbp0pXxQR//OSRES0SI
LwZ6RQskhOMNQi+yc9mP9Lyyccwic1wIatHU20wH857YXHDrEsTDjeui9ZX/jZCj
hWnj5P6USoPcRh8p2R5NUisJfD1xk8yoSW/91jbQyCug2UIf99J6NpHDVCPT02Oe
FeWCKVrsDkDUS7Xs2bw9NmtUz5Lvo/RzAWH5tN5xzTJ6ue1vunPS/Ea1jFXHG+ds
wKkIHY1BRoJaMe0tRtte24hn7HRma0a/W9AH7HJeZa4vyUpyXMKLOFvRhwzueDZq
Zkkaae2wKBHRlXerVmMGogF7GIv7N9XubDQds83Q/yK3B0FmZEWevBf3XRzbThl4
g7x6JJAqOeYTGkORC+ovK3oqRV9jbII0P+sAge8q9Mynp6koKo0PHc2u2NxskAPF
u4fX0hJHX3ANyd8zmw4VuVlMAFnBbU+OZ3SNtlfL8dZVfDA0tH77uPgyaboEX8hd
HPnhJ9garHPkoKs9pDibhY734aNpZFxRjSTUlsYls7+VV3s/UjWue0pNbGyChjul
Zk/gD+E4hoEd88/IwvcTvjhUAHfYsntmFDlWzLIJCmpBJA4yknlhn3GA6XAj23+O
aByZeiz6B0kNnFWb1U9WnOMQE2WrZvDb6AR2Oq3mGV4PLZPiYdTCssxeHtv3/4LC
Jvw2xfh6nPIaxOe3/tY4ECrnNZ6GDvkvXcOS3d+U8xEh4eZyVKWIi2Kd9e7vPnmp
O2X8IqpYD8yVtgYUaHMZnYkp75Z7JpmCw2xsQ0A7FlOkR9RXqTEcMXLJqluKQ+Ai
9pdFT19Gnile4mApb1uGcHbiCWhfMjzKm4N8GLwdow0EPBi700xATxGmdw+Qv5e6
OYdwdFsW/MD0zB+yVH8iBD1XSlYiMtNmysrvbYheY2FfZTDtT9rrwmMtKbla28AZ
uG65ZBbVq1prE5lBIBbboSiuwD8S1Se9ALBav2Jb9KWkuvB1pv4McQc+nGjBilyR
q0q1TY/cyHG1MWtQUYv3vOpnq3uCBVPsMfIUqo2rUh/7mKttR7PjCvhu+OWtd8Vn
/v7F2HS6dpoc0kfiidTGxYEa05tjUJWwAhMUN9SkHsRW79x4+TwsOcQRPteFI3AK
ty183UV3cso8Qio/hE8cbmJtHOBLDC+7t6MMd9jQQCk649Er1k+WhxOJs/S8Xtzv
DmE1bHmX6ylrknZMfiCWWh+E2iQhX8cleCWKTjJyNvWN45UIxO29ddz+Sy1i32zv
CfLQUfiDH7WY92CMJKmZO9f7C+xG8WncXxFc+rUu8xn4mgxG02qcUOGxd2IxqYSF
R+RJT8ZttCzA4bowVVT0NbIG685WHrbxt7Z1/WD9ibk64uOBYrk+0+bAhPa6ASu9
La/N6oyCrZ91PLCCI3Hqrq/aWtBBYoqZvGuX3Sg0e7IPKne0clKQI3WQVt/anZIX
9lydvJo4WrLwuhwGckM6szCLp6jQLzfS1+S+Ib/P0ziXh3SqiOMBq2Kx+C8jJM1O
5hLxP5SaD8AEOk2eFe/iyIoTYwGBbFoMYm1QbXLxsICV92TDVU8+1LigEyvOBS6I
ppdSUL3HpmhZHboqB1k663lU6jjMC1w/EAOM0CLW2r417Vgl2AlvTbntFSy51DT2
unEySZW1AeuhYWPXx7R3sXP4QPXiVjzuTgiI1fxm+LqrIZgJp5lC/oKeSpKwJBNb
aInvE5PvQ4+KOENT9Sna8DG8f8D2TWTkpvsE/9xI6vfbq5zJmOuRv87cnbKsYEkI
o+qbmsOxrHNuYWNc1vOTn72wPYjB590sl/BPhfhqn+lAMeOkw29j97c4pmaP6J7a
mKDokkDkmXO4FkqFnilNK8wueanI7njmz+uDWyvja7K2yDOXyXf3h32Vn3Ny+2tc
M/gAQu9I1L6QebJtzAQxyQPrUOEwPjyGJfuHO/ZRE6YPUm3fOZfWGQtcIHhfmJdp
wf5GRswiL6+iYDIi1mnHOvZp7btnKi7cwQphaBDckaXZQqa4iRROp7Y2UqKsiAHI
T6EMXnjBz4r4irS3LZJg/JuIvtow266OZNroSgJrCVpbP1XmqtaHOPVDH9SvsBqn
/FFErPsbQAC7SjVyZccIoCLsT8T3NpGnBEvYCQwwXN+DUa1yKkVlck3GrL22v+MY
45Zb7QKhSiei3D0waW+EUGP1tc7w2biOu55MELE0JQmlBHFYYWbqcWWoUKVdtial
4+dvSc+tVWaqNCE3H+xAK0IQooLAE4bJjKd5P2SfbgI8o0AV/Z5+pIAe2nteC1bM
WfwVXkwuwHAjIeoJXQ9oAe6uUPtwue3mOuOIU1pr+jGkbnAUl3iq9H7YEaukHS4m
FfJ1QIMjMpoBRLxPYIjcPMDl/srwOBNc5zGVWRAbh94qlyPUudZWx4k/SkWISEWN
MfRXLEbJOvdlVV9cQ8hPQ1071BLUXqs6oM0ab7ViI9S1wsiZGhZnACUF2cPhPWNx
SC/ZoxYS5o26AG1yhLAtvsDZjiDv8sDB+1Tykm9hEUthb53oRPlfhcj1EYrNP8mf
gwbM6srm1IvgKmejp2riiHb+qAmJ/7qwZUpcfUHT3kypqGxODGOMGasrn+XxRrOy
5OdIK604V1/cN2eUxfn65JLkOv5HzQ+jQk0/dD6yT/Tr4hikvdAp1ujrJdANg5IE
po/iIVrFuqCk4Jlit14LIvwg4Gg6JwV5AOzdtlhmGY+bs1ZH7NTn8BWsZgVtE7B1
9nCGWgQbhc+rkdGki0vmpwgJbvRb8LHcnD80tYYZcqQvKMypRhPfcbMvQq4cqmCF
ujz9ybWa2MP4YrL9wa3qkBWc8uj6GBHUtbda5mzFDxolCB6ikd+3aJPo4B/i1uhC
Ft9oFHSFfLnBZJfWzIeS6q0avBUjMTgpVmz7BlQdtaO9mZL3RDXMhKByRDDYWSOC
RRX0i8retq9Z7oPYVFbOMUI9dg+KTfP6MS7BHbcQrcm6MOohUAMq5d9E96KkSjmk
Ys7dXFCBspB+ZZQdeZ+QSZ1MJM11OcaJFDrqyr83cSsJALmWm/GADudxNOpp00X7
1oa/KMxNOx9aislLniV/qcfT/OAukiPJzdHELxRP9Re6V/dMXiqaoRoXkQTHa4VQ
7sUguxrGuOHaOZliZZNxucJKX65K9EC1jwAM5zsoRA6a18e5+yrDflnKbehf+P0B
+63zNiKTfcIbKlK6yts87apzDue2BOJrTG65qNd3lpkehcD0hZ1/28ivOyYbDZRq
d7ODXpWrB3NxkkKGKcatFZCVbVP4Ag3bqvfGLJfK9QuhGIuoCf1Pk8y9ZGrZgRkA
T26cmBDRoquTMsjtfPufbl8S42zG2DlZg9YDPEZ3GvVxs80vt1epGeKm07ZHhrCy
suK7V2NN97EpoRuhMVH4GZnKYpeRnFQuhMRLMFEjwA7YxM+TNQcjlDsMkgXHuqnZ
EFtynnWbufBcclWjrrtC9FGkLXAZ2Ffj8dBmICr9/O8n4bMT4cI2cQB3GrNPCTRd
/em/5BSSrQlJuy4C7HMb5Vv5PU8Zf21F4UB+fS1akC80zMsI/sC+y9XeqVWWE6rd
8NPkgeeiNOm8lgrPcxqBv7nHeyf+PM1tscL/qzyYSKMBVAmPuQF+t6QUk701XRO4
hID5O23q32OEfBfCYeG7RlvRnifFt2BVIWqUS42onJ6FAtbxrDjZMJca37FS7Ot9
rZ1tE55ZE6AgJUN9Bl4JsrWOxpP/P08iix27hRX+0NAFkN4rmewuy+9YilKHfkxr
Z2k2kyW0pLkwP/Tph/HQczOeZZQrNr5XpNnvBeyv8GMrBgFgNdY3guuwh2dRYp8p
91p/I23836G33rIA9uC4xlhqgpYF4q8dhM4o8oJ9t4Ukbu8kTY20msJisiPqHzbI
z4dUCbU6+nA3QG0YOn+QWOYcidNvmejAfQYzaM65fKdpRG02BuRYA5WLnTzzoS60
/uJeiXlnLj5MvC4d5jeGwOE6jdHZvN0lRkrW+BJFLnQZAcn7lCGjpjVTq9HrScHX
UzSx/gnxiSsEnpG7yQ2upaocuGU2fMn73cwirddNDYK/g0eN6r3dKymiF56t7L9y
eV9P6cgamEiBt5KjjuarKfT9mmdOgGUEu39MOEu8zoWV+Hwk70tJhYNZwRHFhJUF
SVn1Si6DDjMlVJ4/eDtKs93E2ykmKafo4wZIuQuEctlHEtATGto1hPT2ndIxm2kl
cvSjeesu4YlhweuHgxzVDwzNxrIgJzFET+E22jSVVW4ZjxBG0JDcaVw8xs4nBRby
Orhfdlr4KAK3KDtmanuNsfWRvxCUp7DkCplD34UJVWB3FuoNUp00Vy3CB0DTT7gz
SWGovJCSz28epGPcj4fTdtHkCe6CteV2W9XnR0JMjuitK3KyKSCRPr9HroKjbWc1
Udtkx7I6sV7+wflB5tZLjNvvikoVOGSPzbJKT9nl5Ype0KycHkE18EA5pYM8DLGh
DxfssOhU8T8+aE3sQbOAfywQTU26g8LRhw2x1Acsryx+sP+af20AXcZ6p5YUqKbv
CJz0Xd5BAmLtyez4hwnHbW0mR2/85WXY2jZ4YHUZ1pD7R8fS512yBjMlyxqS98tY
W2Z5mafHIJ4A4QF1s35179rW1L47fYBC+veHf4pM5Sh5DO+QD9JfLMCXadxhOO5M
uMA7vV2zpTuIesn6pXEuqCTS2zKdO+s9EsK5qAl5kc0336fzCklTP5UpT0qXPCDK
Jq5V4TtZOuR0nzokmP6iBdy/v3H2UcuAOv5hhwaBbHxhWTFItbdqJVV3yFB4yrQQ
TtmOZTqwjHPqtkPN+/GvtMrAq5qvV5t0r/ErwCDv9TzA/khf3L5WVqpAe03pR23s
D15yj4u7uWq8wI1CBMOtsHjIMV/EdWMACeYlb+GS8r9B364kEN6+if1OiyxEpSPq
0fbGo073kMqs0cJgJH4v48+E0pGdNNDtmzjanUWUVONdXmM+WhbKX7vEVUvqv/7t
EUz33is1QCQJZpx/YlRvIDjw+75bNQ6Dl5CaY5fvYHamQlSBGs7M5UfkZBex76L/
OYeGvcs2S0OrTOCuSjrLxHLGqde7bjZyO7hXEmxzCykt29EJl7x5yLWq9omb0kUp
akC0ElJqVnbCxleK56+VqEIYIjYwZ+veKaByvOfWyg0F3lEyhiY5W2xfcfB1uipM
zItR/KBv9xMct7mSCv6ZpQpGSYz4QfRy/rgurw01GZqHTT0td+3mROkWYc9UbDR+
rZhDijyr8h5JWeDB/+NUJegYftW37zZdi5BheVFqjYSMh+Z5rQMnlDKNGv4wLOac
X/+FdkUE3F1ltEl/g01Q7v4zwu6oUKWJPsWeWgBVxi0LN+ivR9MIIkK0xM6/3K5R
FBUkedx7tI9STt+6f+3Tq/Aw64JWTJ0FezrX2vKQlApmJvncdzdDBsI0T0PdP7Vm
gONdVihQLTc9fvXhclLt7+BGpiw8WBTjl23t75JFl+ZvsHiaQDXcdkNuNyIT0vKt
shos1xb96iPFJb592Uaqe9JjiptjjgyB755SkeRegAI0+Rx7w1H1m9dH/1V4w3Ie
M4RC0sm3S41dpdLsFuiNSHBKvlTbpDxDtE8wSKNBPQZi1fNAH3v0CEIrDqPHUl8O
6LlEmSZcDu8NESEe2e/K46sE3CD0RCxecsEZJFUDWR/RVIgctbTJjDvyTjRAWsBS
dxmJwGQTph9vuU6yDQq9VY+EY2IW/UarFwdueeoQ7VsoorOwN7S6Bq4IrfzNGNZ2
eaGi0EB570bwYm6nhUIPNfg0/BSfOloxZOx5zGsSq66qRrM2WquDgbLSUog3sv/w
eNpsF/BtGEcLFs2qo/MjAiDkrL5QZlrNc+TBemyW1uRFUJzHPO+dIpW0ayIoisQI
nDPF/S/Zyure8JrzMwDdg98x1jmDf8UQNNUBXJIhP8JQmd2y6vmXagHSdtdzZgSo
3nIUCdwkiSjzcl/HKd+x76koCmCMktHYOzf8jMF6ZDMeQ91/nmywXhgO301KXC5V
TnvtUkXZrSij9qnRvewa0zl2jcPz5HqZ4RaXwDHdjKuda81pNr7hnqWgtYSANgY1
3bUkHiDo8qksA+6MXmwbRR0+EOYrMe1ZFwO5a5XNo7BslIOF1pQfOAt/Li+9xqUV
GzSI0HU//ytLBAMk4X++JLARXxZPMl9MHOBcreudMWZOELK3CByrZDuSp3KEbW8j
O0udxEdKxs4EGQYpCSk5YCDJXjOaHhRe9o5RGTC72thDc1ydNSyx2PH7/220Wf+K
m5YFs/pawbYJn2lNca4G3LcWwn+32qsV0O9AGt0nToHMwNg7L09QjqyQ6px0SZd3
pDeQ0VhN7JGODQun3cmO/eH5N2dO8AP++ja/V/hJVcty4TuqewRVa5XPmrqDKiQR
X6iBOtCVuAuTIBIbg0+2KA88+HKZ4ouys6oD53WRw/hmnQI7LqvfLMRTBZwdr5gy
QKek7Ls4mCqBpagnmjw8cruITQTV+gchLfASMHCSq7oKHo/Sq3mTlYc89EYXADiQ
A74zRYE8yknn3Ij4znCv5ivPoa4SXM3MVbqlyg3ok5DBN+RzVkWpzATwhL/ai+Iz
EsVx33gah5J/scYWaWRFckiTHD+Qe+9U2G0UMaCBsS2L0bw5qbzKM8f+rzgedHTr
qFeIJCkGMDonJeQkQQx2l2OiznnPUhdU3ilW7uhut5imSvYCnjQePIgoEy2qSzPr
k2M7qrqjeK1JeewsfDVNHt/sO9EOc5Tb+E7N0NAMfS/GJwf4ca5BdUsq3ECqBnQt
1+OMXVCUddE6uPBL7w87Zfhc+uDiN31xp9PMn+utWDAU79wbIUiKoWzwDCPpoxcA
1Lz6gFnF0CSwn+eT+N4kohYyJFYwntRPvnCuwIM/EHp1MuPlSJ4obxRriJQCghZ3
UwN3Ev6sBBQgFyDAcmize3qxw6cQt1bZaO5ZXV4wcO0rtGYNnubbHQiS7zMtDZfR
Fv855fgKPB/+Uogi973zFRU+sL+bW7O3CFnprd5QrZALVdu8SMIvD1bmjVHD7zE6
hqtqkmPbI5PwVrqGTh/X3hq1/641mS7uFA0/VN/R+LBbN4nhixIdCLkQ3Esqpnyb
5dRAyIsJHGcv+ZQNOa0XB1fDb5qJP7M+9lhuosdCkPZ+l3wwn3oy1CapiZv2LDQ+
NoEyyHnYX9jCrpYL9QTaxg1rGrJSGsAd413v/Vd3BnEjHRBdiltyrlbEvuR5mvYe
UIPiTcRrBVSqjhzYE9Xq5k9jbhF9DnKWhimx8z1qZ9fY88MYUm9jTAKYzFKFZKk7
o47ojt0c8yEv083qsqXz6hpp+S+RZiG+03qmJ2g7aascXb6kA45CcamCP9crxJEs
IdrHxviWXuHQBJMhjcUpvG38GtsjmdA8wqkTWai4nADpaxEjFZWxhLkYbR6hT4H6
YDGz7HVi767JidMMgGQOlAjQoS53SQpubcU4YGq8eOCQmJNRFIGZ+bsDnl+Yyqsl
fb5tU2EquZBpIJwndqIOIZ6v6heT+/5XM73b9+xl7JyvRJqfSM1ilizAnJj6kT/3
GbFpD9ZKQ/Z+v1jNysuKy6ZCQ54uSm5B2thAn1/5XXA2qjsLernIg4XGSqQZl2qM
eJaSVsmLe/I7lkaQICbPkns7yB9xzFGoMZ4vhNRpLowzojn9mMTwAgVabiZEEDEX
2LBnvaRJu+fPwj9qYfgqwwygImjXJy7KWjEP0LtjGdd39oOMzVwDgvYffw7P24dt
QbUPdJxwqmW5RNIorPfwcD4tmJtGcpUReSj31vgjWne9jLUuExGnY3SCjQglATNj
5U82dP+5xdjr1iKfainc6+ufLbV0GoV2xcJJo2NyEMZbJVpYDWZZSnbkrIkRB137
vupCANrNvq+kyjbyXgiHPtEzuFJaiA0euo9TsgyH7Cn1oKU9BPhEK6WvfHxIzqK2
Ya0InquCVXbGBaDKvvMauzrQLnBak9k4BYSkC+a9hbkhf+IFY5m3BALs2tWC7W+h
0QF7W+So1nONoF15FXSR4tf22cqJ53bu9BEpUtCwNy1hwQA3I//sMKBEllOEIDUB
tLCv+AEoQNtz68TrGWOcoW1K86Z1AJuLYzwIqdXCzbpQ6OfJgVJ31GSfAt0bllkh
KobFf2/h/TeFrCO0R+gah0HcbJ+5v59S8sda0RZdyRmh1/0CQ2siBsGeA3xuFswz
nS+5iYbhYmuPXtGqSKYNBcGDWReRgpcXx3hcG8Yuu+YO2gBLWegI5EcoX3HRT01u
X0hdPXTHc+z/Y578B8b/HUGQX834Fr/3UGuvrtvpin55RXqC2j7ZztSJhpvkYPM8
9kE/6tKFYnotBKcIXVPJWo5DWwRuf2vBEVbZgloJkrCcdlGOt25T9iVahYjNz4Yq
oOyGIwcRTlMH7TTWMNJ0lRjdsuv+d8ljZKMdHwAjJoMcDYjLsB7s5moHY4DnTRHy
wTR2pmi3SeKwqjLyI6IOWgvuwRbfL010UoOMrKnJIgGEMHOJuh9vOaIEO0FibYcC
yULdtvZxB706HZwf9lNMTt437JOOV1X4/LIUo9TnzPQyoKdEVp+GJs44z4WQ+PGL
rGRQl23hRpWKU7Q8O994cUmoOQlepZAdn0XnVtgjMDaEbpXhq2GTamuO+lzX67W8
wnZadWY+KnTxyeSysa6U6AGem9QclIISK2Y47WCZiRo92LJsFHNJcNLtDhbrIR47
k4wyTB4tNTBIxwsBVWJ7+7KdpC+MuPNwn1ttuJE1Pg3NYcjszZOxkSH7/oyRdM2t
42G55U5V2VvEtxNL6J66ZN5NtWWt+yaH8sFGLlApcDEFQDRIF/B9LK2C/DD1ESFz
X6/KpeNlQYTae6pNTAe+jLpaNpJZXOl1w1ffFjMruWZIsHBreANg5hcbgMMmAa2B
qxRVrn8IXGxo4e7Rse81gcb5NQXgg5tLH9Tk8KKrqZY6mgy3lDT6bRmHDbZQ80IQ
mIEpOUy6XtY1J+e5/DNUFRWCSstoGLixn0/ZzxEQHWPxKNZNuuwkZ3b61EmeY2GS
cxtZqPS3UDFufSkjlLa06H4wt7XGZpMMNutJUSVNW9zJaDj6Sej5QyDUrSese+lz
zxvkRA/0nWXojaGeZvKCDudlmQ1yEEq72P6FULDhEETCMaJQp4pwAgbbS3GLpr1p
9yyrBaOn/lRqC3lD8aX/IZTlWh4Lsj0aT2frHl6MbRaHttV3ICXgCJBUIknXYF50
UMiphmuEVL7FEOQVND+O2hKh8OAAIwbVPW7fiUsFG34Lqaixgyt0KPKAWi12+JAw
W8xLzy4NzgHK6+tJ+BdyahqChhwY/TcgOoUL4AY+D2w1klqUhtBLp+oOvCbxyHFN
cgoPxf42P2KMI3+/Q98rzwXQ6XHZNK8cUYnOSLA014xVWpv6W3sfYY6iRvFMxVDb
h2CAqj+/3TmhmU1KQJOwhu9mgbZi8dUeA6maZDwo7MTY4aJr+Mc+gOg6nXI5iZdF
NYSW457e1c4JkILrC2zIzZsR8wBD5XRpo4cj/uEpsg1OQ5/ypvI6VLBgzShpaSsc
9G6Hgv6/dLDDSpJVk/qY1zSFOdnpXMZ7Uy/lqACjvo41C++51ktH2HYXw/W5F1qL
i9WR47LH/zbKd5JFi2OPopupVP6jiOzvu4Y9ZmdaSgdrdZzCLzqSeCvr4lOBUr78
xfk9xmGWk3VC5IadblrZQK2vdepMtaBw8WCO8HsJmIaAc3CFWcGtEC7jevlncvJO
wXsrAHtYloIEqkhWjF/MkGvwC2Xzs/YUKEM59Bw42rMpjkEqOGnV+kugmQQDsYnY
D/prcJKJGEB4MT2Ry09CQyGv1KbvYAAWjdGbZPPSPsNe+0bm9RJ48wNqLnhTwc0c
QgISjNDRYCImWxB9M9Q8Ul0psd8MpWoZNGq8umyKwX2ERG7oHKU+R3ZWi1OV/2Ek
tM5e9EL9wm9yW74ClNCFrTcQgNVK115eWtRTD6Z692hLn+SUDhbvy8R242t6zP+X
62U7RrWwYyRKxWpf0iWHU/SEzykplEbbbqpqAZseeQTyoHkqL4NIZU/WgCCJy2d/
4gNirxWEzF6BovCtp6JHHoLvy7dkcx3LOWpd5xDfm0i2dtKIahoCXyH3kNtbPrjz
TNvXuROMSGQmVsbej3IEjmxLzmdQjdoKWP7501hX/Atx5i5ipbx31Xza93Unlvp6
VmexJtV4QpOCDA7OLDassI+fW/u6Ne+PTEkKj26Ce8wI9Noi8G7rK7u6zX+xgxyL
ljnGtjmBaGzohTmNKTIJLKId1dYocbP3TafhX2f4BqlzfAp+T1Wf3PYi37XAgNSy
PqpcewF8y9xlBJ/2XBT5OezCT0GpK2qEHmIP7FikZZUsm03xxdK8E4v2w9FWFRg1
Sb/pl6C6TPRhrt/SPa6jmpecpSaDC28PP0yYSUk2KSVR++ioLqQSU2LRHJrv/+Ws
Ns5XWjPHadDg0H/SvZpOpjLixh9AXbCsWGTQjExy3tWCLJozdvWInJawTtusIbsS
oTYh/TtJh9P9byvqIyR9i/wSDuhiMVXgTYtFcPK9hoso5TUG5EELNQaqvOtQ8/xt
v4uITSvKyUUt/9kkqwwEk8WCiS/1nwNNfFhkVqrwvQzXNfRswSIfQAY1VY/cmyPI
vKXR3dtNwXNizetnvTn4GgNDECYN21v+F/IoEMSnVcr8BDZ4XW0ryxn66VN/O8D0
LwEiC6pfzYcG/SAF556dHXdMlbB6/1cxE4QlR3nwPNq9x8LwcR/B49e/Wq36QFOC
z4ECfAIwwoWclvx4XTkN7UCxwd/0GIpDdTI2g9bSFS998BxXQPbsdfbp2vDHRSk2
9n1/21d8MbKbeAtpiIqTjBC3UdcLIDTziBGvrb20ZCc8bh0iBgWdUuW+Lp5nO5mu
bDrzsqtu13SLzaKzEDkAb3whj1vrQzzfbGYZ6JXiTNhKL4gPcS6TCZNmsq/zMfOa
vrehkwi5NQNviD/t2GA8ouktpWMyo1cvQBZaG96/VXWyOO4AOu6Wo+Ky+1OMlAuo
ylQJoqshYt8eWQ0aKe7xfkgCU3xswYQC/Vqld93NAl7SeHnWWqZUJGtYrKgsJT1l
vYoyk2s9S4/8LL8mk7ecwtY1xBP05C05jl9NGVEnDO5rUY2I+wikkqTXr2rQx69t
n9ZKP0kE4iOOKYoXNKOepp56+IjEV5p/c8nXxfpQZbHZvPFKjT2hYeXNDiUCLrgT
mD0JGkmKjVsvCIdIizbzkxUsYP9PMgAiaYVNxXjwSfj+3dUbNYaZsJHyaJOupbQu
s2wN10KYRXo6LMcbT7df7+3w0ij8PJFdC3p4BbuG1wCf3Cvcb5FUfncNABRQekF2
hJrAR8GWsxWBP/jvUgl3uvPzMEYFx5x8QOA9fmVS/jNvQY7kZ2BQyrbEoNMawQ2k
gHm6EhOmWQQmbMU6C3Ehl0yX22R4zxhGMYSZ5SXh9t8mc69HnPJUzecEdIS0craZ
03uLNkR+nlWA4mjHqJJEmTshvGn1oIHkdJSvNJYwZUf9D8dWYrIV1XPOGU3CKsXV
ArJDzT32+qN+UBZXqu1KdXP9gETrmV9kDJYjrsIY8L/zt+ju9QjKarlwCr2yAYeF
M3c7eyUn8kC4ytMYwaEa1xs3r7LLL/RktlABKZWbFAd8R70TXwEYeuYurUBfd71U
g1KmSDTVMrQVuhgJkpSXHar6d9E25DsAzHqRh8mQK6RZLqmbNzVgiDqgbOncAl6i
bbQf9NYge376XBnO2X80r587r7tRhJdqCC1NlfRTY/CZ9M+uBK6uUbnCjn671kdk
z6nACcBdY7o9vyYHU7IAmjAJxVajoDyRQ4brYL50zPcqWIpNmmiMsKwXkT/vwsMW
zcrwuAztpR23zLGQHFpea7ig+m88SLCUmhpIEXlSIm6x2VEkigIrTFTRBSvqTwTW
M2fcVZx97qApdbUviT4R+vHjfmgq8xNth+lnkV6vhn1+wCilWpZ5KEQLJM1tcEhK
50HsiueubiH+nXxRO4ZD/i0meLhi9YyP89LZzVoxpjjhi/k/ww/MEog1+hYmoS+I
x2WDelMLcLssTB6EKqQ63HilsKltYS2K8HYjuusbp4MdwayFBkQ6VfAAhNDvNxJy
82P+msiUy18pk3AhzkKt6gCBh0pNd82lRsNMXUHJjGFU+uBqYmKq5O+QgYbmPTG/
Xx0x9FMO7pZxWa39D4F9I8p7h4d8q6xhitWJcDse3YYnqxraY2m12uHrXJ2NzRD9
RWiblHmQpPtoo9yDqEvFoIUl7yLfmRQGtSzWhsNkQINsKQ+atEg+pWt8b9ZFA10U
77XQV8Yk6jrj6JBon2UsfdFtjMKuYHc7cMWJOvemojD1m8mWdSVpCWke2P+sMBS+
I4F9DuCmXtllcrDHA+IyrsBwOUdJG2IH3u2D3ptJewYiBf2Gm0BLeKmqAT1/L/2Y
4a682xeufMoEcNwUdAaxWyleSMbxaj8dKHF2VEYTMAWVFvO/W3kJZONE+zIKn5b9
x0NzpiTK52YT75AxVPBtnBaXqXimJOAaqbt06IHGg4Rg5U2mNdWWaxoCjqwoCRUz
jWFW/mKsbIH5SXyW5T+zoM8+FU9oQCTbsiHunXCQKkuhQrOD4bpd3mRCnohdQizQ
vTVdrY3Z7msopaie6XK3wFys6j6Ln/eeOO4Es6ThFJz2tD5alhYA0Lh0q87xTdxR
Y2Y3MF0TIC7MP/oQrVed6leOjNVwTXMXjLadnDzn/2NaF0ClZ1kkcAUJLaKYD0ve
uvIvVQUcy3DXgNCmaz+zn+Akbw0vDzLjf3CA1aSi+jTMZQWxzkvxtnadrd7fo9+v
LhuRwkm63ll+zHG+7uaCJU6hEL+3qrP7MbBK5LOfS4bmBWc0Jlay9+hE8DNcQ4Y2
WNj+eoVoJI2MuhvJW3itxntDqFlObVDcsRYzLPmab65u25wZYf9oaJRxdzjaAjnQ
/Hy/jwms+xeNC2LegTXpq2ZMY/MV5q78SwLyvJ0a+s3d/4mePtJTZ2w2+JM3ik3C
dDqyQlZID6PJDBZ6bO/1tm57Q9wK2XG3jcl0cxJHtQcRCShGbyA1j+n3FhnqsQ69
/GMaY7p+u1dc7n9tCiJz6NxT3+9N0muphCiC0ojm7p3wFU5grz1c24Ejl9FBiWPR
VcZgTSDeJe4nIY/6X9sxtFuqDqh7NSnycLQPhrlrZpbV2OIKX7WH+WHTcINCfSZa
197MnRsQAh6P80ZCdACEcBMJkf3c/TKPHvfo4kWZSt7t4wp7LjoEbnuIGsn/fY4k
zmu3MbZ6r5ztRf64mYwd3b7tRzxwypz7eVkYd+q6aWAPt+Uv5CjgkAKrjgz4X/iY
Aq4YgZ2LZ8TwUATQ9gwH/cQZrK3203K/MF4LqWBfaQZX9kTQv5inWONv2JoNH79+
fYnKMP0ctM9HK2fbWPOWzF5feddFgvg/oavXK3Mi99n7NVyUpwVvTShu/jryfFUn
LwKB9uKH1cqgbor8jNkG6T1vb2f2yCuI1lYgIQzwno0w03M1czQaNJQcTg91oPfo
NQyWQnkfo6FDmGnfZOUFnWx37icvZG1U9igwBesS9KDgf+XaQEAg2M6smxUCYebF
L+w/eiENx7uyX2d7ULg72k8a4s3+ziVf3cPxWgdjwqQLWFRE9tUVSN8i0cSP6EO/
Fq8/6olAoMKd9xmoW0hQ0m8ATU+ovMsQoD2nP6+ExdAa8LJFUSsFL2mgjY+s5db1
9S4/mRWcPEScsHl1H47Glez5A2yZyDtKNP4J2FKxesccFHWKOLu8f4YL4fWW3jFM
PiKRQNqudTOchC6k6l8OPRcW3hLrsBksc3p8eTx6l8cpvBrq2raARdCj+dhOgzGn
BZkIabAEah9rdzu4NIYNbJrS2tr+HzU2PyVJhUfw2KSD3CxdcG/9i1s8wYMt7k24
j0t6mUyjQFLJK+nWzbRzyPb4BeE5vPB0XU4HPRwMDeKap6UO4bVX0lalBwX/W/Ki
TW/v1/3jh1vUSIUpcCsVB54Rd5MiRBRdheL8twxYiITIwmhZrsSuXDQsc7S1kPNg
3dytL1N6/Ah6vVM4SE1B/SRP/Su9yZ8LqjYUb04iLr9sktC5olBqDS51SMXepO4r
d8gWL5qKgPwjGjius+p6BCfMlCgiLvzfayIgvgcT3Lo0bwFWHtM7UWPsOMbdu0eK
aU7inQUAr+Th6E9oBVTTcfwg7GdxQhz/WM6xillij0M/Rf8YG8pOusKOXmxXJsZH
lLhJtGqJcS4NlJXiaSE/rAWgkvo+MYmoDsyJHQir6yvnRnFT60z3FE+u3TXjKiei
d0wAmBPgHxaL0Wd0fSvJiVD5elfUOZ2xqOtRUPKwPaJ3grvPyP3eQAl7Br0dsL5w
CObqt01jb7UIwtEX55++enT2HBIo8ErLyP5c14mfvj2ufRspUsBH4K8EaY1+f+yB
QXp6n6h9pxQ++ivr76ILOYGpFgfLO5ZVCDviYAWAREbBhkxLaUnLp90ru9L1e9Xd
bRB9wjnWb4iwkaCemKypqCQft9CNsPmG1STn5rbV0wV7WHWmafbDTadpnEZ1QVOr
0jVTAgM0tlgRxWUDcxZb4RCM9BPdwKcxGUSEEyNzsPktADEDqDTA2c0lgf149hXr
MPfQDc0HtTWCdaW9HWeIRCbZ5upYREbR9JCAfxAASpYXNJy4eJNw9DVods98kJ4Z
Tf7/Zd5uIZlYaVEaiYBQQxErfY6KZ2boe8QpBLX9BtMemk3T68khH4kbf8gK9S4F
hHHRdBfu7JFqAeEmOe1QVSvdVYiASGscNw78iRoQSZ4zKWlcM5q4q5mw0/uZWMxh
ADt7uyLab6MRafdLQRKrWIFPbAxqPWwOplczhHm3CWmcrAw9tY95ES4LN2X6mmke
xGYtuMPpNZvKuHL69TkH970WQxs390DVBzjg28joieILt3Pwwz1tOJ+W6iL4XjV0
dUd2Bd8YZqbPbmPLG4nqy4b0KWwEx2be97JG9xvpY3kFD9EtHRaoIG+E9Mnz+UnC
AZ85JG9LLyV3Bno4vcI7OkPRnijdPj625ef8e583Fw6o7f67y69mA0fp8fguhAaX
QOT0p0VXlnzLGSaGj3/ZDEHFcUtqZGnb1riVQJbh2x+RWnHARo0A8Aa+Q+QrEP//
CWRaiLYxG977wXcFHYnRfktc35jmh0FSUaOp5IhubCU2RnbmHfLpPBNpbEM2sf51
TKtiPxVoK9fDoJiv4R8huM5fbHRgLIbx9IUcHcrMItrRjDEpktzR4siIVN64Z06G
0VHj0YVB5LMFw82xk5gYn69V6KvE/VgaUT/35ew9Tmc1EEpKOOlLPR2kELiOqvsr
bIghpPim7ErsutEtHB6WkwsRT6KLAxIckRTxpdM5clPOI649zZJ/Vhw5oS3OHR8I
Tl75vs68mWvROvUii5dM6j2NuQWP461sN5aU1GY23crGv7GuSoTJZxnwiqS218BF
nv4HxroDRfSYJs0R6g+iz6ohlbCbGcRzCy44MUqsZ9sg0Cu3Wybr2z5tGAPwQnsj
daWM0L+U+fJ9Tp8RNMBT+un9jbg9+5zn231vDtEddj+RY2sad9LzwBzOLiqBODwY
28Kw6ZSU7CpmZuRhofNgQqds78DqTpvug+vVf1/Hquj1DMP9nD46XNoTlb1nbtDt
/6yFvd+clSnqmXY7l6v6A721jJqmwix8HsFyNxRI/vVQvVsnKSLFkVDKHgaUO0Ik
4u5MV8cKTRYwejo64ETL2irUml03tTOWRkSfyMrxD2ZfcdtALJLvCvJu4WJvcUKt
vQZ50NdMFMot29unZmAfN5v6veOQSufH9VGQcq70/AymNoAlhNUcuZxPm/lRx08T
6YAJwzZ1SrALu+qUt1Y87+SRNjGG6QEkdFIFB2Pi0MNVl+6eqjzATy6PpleGaGw8
l68ZTFPcQhHXzcQP6OaNF+Aw4xHKkThui7RDtzvrEusiEUtL7+uKuG9HDEeiN4aV
KmbLE/xf3yd+1YjzFSRjdqPAGKMCQHP207SUQiG6mO/kIShay3kNdOTvr+Gt3N3P
ghCks4ClTS52sjd6EpyzVxuU/Wt371cSHPIllpWGveNCUwQ6U3Pja8Bw/zjouDuO
py7f2LOlD80dJ7Kyeh9NRmSMZtcsymWqVAx6DjPbkGXBDYyJ+SRUm6CfsC/gd5wy
OgIM+/NQqZS1KKSBoS7ORtx2lrmngncpCP9YyZFohrz0S11kNy7vy3nVllaaZLt6
orfMAbL6vnZ+u1TUfBFKV6gscM/gKXtre1OtvuX9d9H45WXP07L6EpWYZ5JbMgtA
7msqDUMHIfGsVB/IvnULNPkETveIeE3vRyCu+fyIFYXRpCh2dEUhkLnE3Dcc3dFS
Bm5STg0KJwe59uBf5lSuB7L9z1ApnHU9+xhy3sPaTcekQSdKv4Cia/p+kZlT7AKB
GlfDRJDB4v4GsxM28cey96vxaQbTG012+hnGtYi7SLun2MnGGiqdITAVFn4CkD1g
0WoocJ/55enMjxJ/XzScKXO6s7aP2LJc/UtQEfupgG7jNUR52mmDMHnE4m/9RsI9
0JpTuQTMFoenP+FkBNEBpkQOX06WioJUzLDcRNvZ0871+pozvdShmOEYSnC9KiSv
gm54uv+Xa0A/HnepMK9UGslYw7ZKhNsoBX4hKBZf7vFRiBvmx0aLqd0Df8h3K/fd
8GZXkwGWWIYuSNZOUjuusYEiQMFkmgAlku468ErKooQ8MqepVgIpQiFlhHd/F7CZ
B+cFWW5ooX3fl68/kohRizYJv+GjFpsb6h3C/I4gtMf2JnH8rnGDOqYW18KKxk13
Opq/I7549BzJZVO/+Dd+Uccu7YaLBYJXYM/3baO/Kg2M4gHjJxbGQ+HyNOJj8e2B
OAq6u0aG0iZrtmGG8KN9C7+zF4VtbbzF0dEewOSEqWVHknZ5vyKiHZHDsf98MTSD
nXPKFK71iezpwuws6nYTpWEjfiZkVOWG05YIqFIHEtF7bRKo+D8N+AWHgCq4F/Nt
k6Y9++8y3tUZEt6ySo1Pgcknz0pPyh1mqoGr3DGW7uPcFdtA8FlfXtBzIe5gvq4t
pwdZ6AEUsdh8sJkT3cRm7HysUFJxHHFSd8VM5uwUhqPZfBAIKmJq6HVQcOVBWK99
iRcZV8D6X2H42aZzf5OJF2TZZeLRB0P7UVo6YiLjdW77pWxnqi6lSz5Ix/K6pWgf
wFL28lmFydcl/TNgiznV7P4+KCFo+eVtlS9EHyPJpKK/J797dz5LNi3W8KDpgBqg
tkW4lgEDbJZ0m4EF9GdAYy0T0CIX8yck8LnZdW76ov4GoreStAXhdn9QLbdOR9cr
80Whtkh3eAlbyWeiDfI8XpM/AvC6qsQyT2tgdVHJMX5mR2XxGFYrhgIP8qE/Y+j8
oMx5l8sb5BIrEN/m0bv7ISxYb4lBOgQxLUZQw9utHWyoch7Z7JO7y3fQ1Do39IwP
aSzlkvVh3SJhQTzLPjTRgSFeRiDbXZjR8busagU5uUmFB2/U0EsvfdAXJr8Nsnhj
Xt4NebaJAS7Hcv4VfPUal1rvagADXDVH0IdmJuTcbXhj/6BMmWZDqM2ish1QEuks
vOd9Np/chcCVm8WnSS/NRWwAPt6YwDM5G8SEV9DiW0GyHHeYwB99ObtirmyDjYoA
tUCizyrifiW2Iv4ZNDwTed8QOZcG+6k9fGcoUYQTNlS1WyXYhchtxsDeUBys8VNE
lMhH6vb+LkWJhbqjcYVZKPg2trRD9HRTJDC3FcJKJNntarmd+ClAmtdhYLTD1dWc
QSYUevE8TNTB+kPHYEQy9p2q9U3h8kXGj+wRPHWoo86D8nIUGdLaArcr1mVE6V/W
m3m6+wFXM8KSlkRV9vS99ENy/zZW6renojn/OOdz3R5yUnc4Xm0X7nPO/6mVMuA8
40qaly0pFTXQdiyw77jhL+JIAnIERU1SL3VOzId7akpDVcn6DOdqsZD6JCJKjTqT
d+h6fPWH2SINL78cuDbx+fjOFlaIkH3bSLzMcrbV6psl3dIOc94rOv0vOSgmeqLP
53f1B68fkOTNjCP+5czYXgazLyiuPIVUtgV/6t/eGnb7g2iVdxMQDzCRNxcw2OYS
I8EAds0UcJsnS4nPLq+pHt4OrxfHCK+mTEf4RxRqEvBF6GC2NWXBSrYz6xbhlpDF
zDKkxSNdL6VgdlUg/cfMWS9GIRRd+K1KMeXW3SuSZuDLYDJwF+Xo50hdLeoIM5cA
mPv5Ct490tcDuBxaqPTtlG1kdewOEpx4YTLNg9jXXDXqL8EA83WIkytQ9eH5c4hE
lJFHlIsret6TMM0iDBYh/fYtYGmUn52QkIrzYWRPO+O7+bdddnKpOiajzMpxojLo
fEq+DZYaB47NL7ZIGr1J4rouqoFsT9R0uQ8iwJvye0irbWiu6Mk36Apq6cWfKY60
BoO24tBbbR4baIAEh0mcIr0WdvB9mhrHAZSMZXHCq3kpFs4yJUQuUblsjAuA5c/i
ojASj2L5+CpW6ZPC00ElgHn56F83yF+lY/vhv1x7Kc6Qwp371OGTes2YhaQ5HMqc
goDKMs2zmv946fAePBYYixKU2SOptu4ejSAbYFjH1r/YezXr86Q7+953FcRJ/CyZ
Yd8z0lMZPqWni1PUSCRhL/w0czWZFJyyF5zj8Q9jdtj7o5vnuEjyiGDn4TjKPcOw
ipT0jTHGmgeWIFYLsnh1K64I1fOh7JDwskR50PVyjrz7wXtx/eGcBrbbxxd0ttvm
AlmrIAhJJ85ICdLajlZmnXP6ZClHyuVfEqy9MUS2w0lIbXXyd/3leHfdQGuTR6K6
+FpXUnczGnmBPDqbtjGZ/Xfx9NUy+h1r6Opeq4/D/SIL9RQufNVM80TPI+OOetdh
8DaDOSjALOnx0+ZIc9tsBX3L/Hl6oPB0bXo30h2D8uZtLGdYMFgmNxLkGAYM1rnM
iZdYec4WGDYcwi1njIz1DrCXVtBOnarPqYUPYNHuECkPhu+wfG8BVw164YyrtMac
tHRMHfTzkQjFpQ3sfX3oHvjXrXq1oMzk+2uAkIKR/lk9AgqTpmjBuxxGv6UCIDvg
f+6wRzk0Lfdl02sFnP/HjbyNcENXLy68KYFoxZyFhqv2IijbYHuGOKhSiucusdg3
ajlyHEDInuWnItYtxJh8xTPPrTxgi6RQxJn8wnodG0qoC1Tzdyw1gfNm2W4kONQl
lVdpWR+aWORY99KbdTmIdUUjn4y8ueih+hMxw/QcySMd5jLbsiFi9AsQzzM28zJN
sIIlYGz9hF8qiNIZKuK24/xzxGf1UpDlP5lJvbudkC8pVIqO49d9lSouqlrjUKSI
wiH3xywLYt3klPiHt+RQAJ24q6V1G7qUGu1nSCGl6FedYQzOeJ8J+FNRW7p5ISRg
YKulV5Yv1j2oAnMZTPJd15Nqgwenf1XgpEt7bFcRZlIVsf3Cde4kg8Xrrag1aav+
P6Lwq4w5jFjjNLv3skgL2OBx11PSbiHnUbhKfipZkrLdRLkOaSFP6SrC2IOucFGS
B6jq8MCHswUdkwh3m3IwNKmKrzUdNVEqtkYPjsiFx+UnQ+VANpLpo9uyHoe/CE9N
IG326eQe9pHsm94X0iwbTERxGWkcqHpv1mfgDCKZrKYaEvyh7fEN761cY/2q6SOG
LWh/0iRqY6CrT3ySefkAC+IntMr4g5WNF9ssU5TPPWDriKnRAs/RdHVX0R73tHka
W5LxQVaw0C+672ZaOPvHKCVci0OdO7AUOmPbRTDTg/V9E5DI3PtgvLMfIfav7wT8
bPwFyp/oeIZqyFTPiWD9Xq2ehFWZKy/F+gvRMkfj2Q/E4S7fHG61OA/ZC2YJGCVi
o+z7WJB3OeTZIxdQlPfxUbiRT1wKoNft3E5Z9u0jZmP3037XCt0wVp2YYxvwbIC8
XmV/lCQTtQzjyIBzPPO7kjrL6zLhKpoQogM3vqa+wHb3jcO96UOX0zc6AFWOHDUc
iesp0ccCrN1/3sSZM1hcycXzdxyzf02bz+i0qpRZLDRKKIqO1AElYs2WTISWx5lR
izNDZ0PuVIRlvyqK7r4Qs+70bdyUfLFXJXc6yvbIae3Lvdkq6Tr4Zd8ZsTgx8XGv
r6qLxqpSLIsCZNezenJMvGryoRYu0LyNGK7GkkFQqyWZ04IRAnScSah0Jmz88EWj
nAIGUdeka/jXqM7pKhOdeb2Moxq8rr7PER1jov4K80F0TsyMt9ci7cLHMMIbKbqd
GbDwWM5CUfI4WQHAFJy2oh0lLIZUSQ4mHCox6TCgOHHtAzN4aeVQa9EI9HsxJos4
ppnm0gwdh5/mE5fXOu6v3dNioCpxus6A6YKB638nfMOJXDhoRG61ovvU2EYSMraI
qLYB0K91lpdltqpfqSVq9onb0jBzU5q7Y/mN3DTTq7k5GFsAreOGvMNW4k/U/eU5
/isI22dLcFoNZv+EGLODk6Lyl6lXN4YyHlGrg+08uFgrwm/6o3f7BWBM0GOME1a8
tF68KmRYlGuyKh/wmS+oesbkh/1lone0JskDQsi2j+fA5zHqIAC9Dk05fnq8n8Q6
Cpbl/k04XONp/DLtBygUDPQlY8zaVFHzEu2JBBhDQ0DzZJdW/WfBe6bf4vAZ6jbf
DcYen2vYK5a2N45hnj6XbLpkya67KAg4F3R8X4sg5OqTli5q5wpC7V/JTVzGmJfu
4DgZH6jLmrcrxLeltosp6ps6olhrOP41p5v+zYyk8SFTFy/p5wdHQ1GpSr8kEnbB
pOIPPtcz5jem0sEG9HGRob4dEJqngfZWN/C8lLUy9rqtMmXa7MfRWxCPSglSPpMQ
EqRsiQ6gVXGFeWL4ZT/a6YBGTw9iROpWsZiGw2EWZDUH1PllUieZkdtErsRKRYL2
GCzGdY4kBZRS3mXVNgMjm7Wc1X2imr3ES5jDyufH1DJqSYFjDHyTHmO5WIPWn6cW
tcVctUOgXuOnrf3t8tjkrunW71CIhAZ019WvaKwwluzSftNixgIXKRJP/OScr2GY
rdbDLSIwSVcRSoW4YR2JDBf7OhjyK2fNFTLuuCeGsZt+eiPVOwVoyRWULKCVzSnu
GaIMoHZ8NHalU9gBifMgS2eMxSaVD2OqbxiQekJEvcJODkbgNHJ+2TssMFZ9WXkU
YLC0Gz7R/6K+KRY+qoFeVUlCZESrf3hGI2mb0UDqAdwCJ7QLWFtrydnleDRLVPSX
KHZMJ2Vwd4tK0pxGUvbiUJ722fdirhr59VJZdz2zE53TPKvQ/YdtSW7Cj6ryAaEG
OCdkx1fNvIGj/mCvAQONMmo0l+bvvmcDjIVkpCroqdsLcVjw/z8H0KOuksvTmOPA
zLcRteyPB9pLPVHTgyQi7e5dx93sAmbt6jU/C4f1ISHSVtYEJkDKCUEgWPuD8do/
W/vMUGyeN+Dva2HgnVENH6cuUGKy00p4G1dyi3QfjgO/cx9r1ZewacxDPAM7+BZs
rmEdtJ/0n2T347Fc7r7ZymaPt6PIwUTaNY/GWP24Avm2FwX0M4D1eyZVmrNNk4Pv
zatHN1xeR83oUnxKtU15Md1rSDdo239GROGgvlD9oh7BELG9EyzEIBXiT3tbZP89
Aa3tX9gJQvjY6s+YFRHk1PHZ/W81ZgLtjd6v/kuzyi1SPT0A0J7S778OFksWGsFB
TSdKdpOONbMwfDYLlFcgATd1KV2Fcva8ZKlPHKK3bcuUqSrZIEWAUvH6Sw92pzJT
ZWI7uwKnf5/lopDLLZS+cAg4/41FIu/l5uL7oW5bE+d1TqXA9n0aU5dYzHE43mec
X2/HL1L0ddDLFARUO8Ea85HX+aUYLTRHOrrg5MV8iHXLWH+E1IQNE9TlV8LU2dnN
jD7i5foGgn/WjJYBzD5q/zenZ6MYk88kIjjmVQLF2QCSMFCjevoDiox/qMsNgHMF
SSVo/WzYmU+/noy1fBbEPqAu7Wr7CIVrS6JyAgAFc6FGlgMxo20CYMmP0oFOQC23
Gzc27FYMRPmu+13ia/BVaEfSaKZ0rDlCeYtJgsLMltJkI4btPxzOO/ThgRZG/vX8
/dD8phEjWEGFGVfgD0B8nXMcv9tpEVgreKwfmUSYlrzBdayTFLBVXSij+lBfjHG5
G4r3/DfiGiBALW16M8zTcI48LnZ0QnwPvo1HB9BANuycMoFVai7KafH1mph8yLLH
g4nWmI65e8JeMtoeTek12XAI9bYjHMzFRJxHQp1qhNilOjh2+omTnRUZeGqnR1xk
u9OdvyxXNjaX673NRFhhpAz9eMKsjygF/J3+eHXudqLqqbO2dQvPjvdOBGczjpc9
idHYM3Q3xpxKBSJ+n2z7IBAXaxHqI3GbHk7FKMEeMhP5qeu9czxaCOXKxU6obiRt
MlaUrMrFzGTp0X+MlcXcVyvCK+TorQof8wWXf8HxFTmMP5tONlEoxLjsvAywAOYO
22H5CRsUZ5BfQYhMztezFtEG0iRcp0/Xhft+U2oFaFU4UHKz5yzIpoGEdxFIcdB9
yjzVFZh1vzH1MYS3g5+pmrfGzpiet58w3cy47ti1iB64EC1df2iSU08DDKT+CCRh
kLWaHReAk3s2ujoQIuKmytcg8LoFQ5B1xcYfuwMCV9jivub6HUsTcgrOT9BR1wLw
HTlaNVR0mJJU1HfSTosNAI6NP+/+xhFXxUvX5wwC+Eq+ZDrBNZyAtt5toqUZNmvY
/b6Fcq/noaPB1EW1uK7fPff90BRYWG4AD+lsl85LUwUnCOYaSfZrG0vTM9lwO5oZ
OFnuVj3nmYOiGyg2xrfzDQA2grxpiJY7L97rLsRBEPhUfGTXJk6E8OgZdIqbesMO
OCEeAxxWIjNTb6wGb2VU3CkBv1LReENn/nJmVJVdqVVszrGFzjUKOyGXhjnvlY9J
0blf1rNZ4ufO5kXWWHcznh+Y4MiWcVCRIMWaylzA6+QsVjvldtg8eJU+T2VcNRi4
LH5BEcBWePaEXBwkCEsBaijY4/FwjXCJK6T4VbGNHL1lL8Dje65pOjz+0IdovcY1
nmx41wzVgT3eXBwu+6MtgDx5QEihe9N/IaKiBi9A09tRvaFZvc5ZQCv+TZVAYr8i
oqKon4Oxsp93BafRgm4PgzOI3AKQiFbI/mNOEN+aA8iigQ7BjWutWWtmVIeidd0G
2ksXZM+prE+3FuyWUQjad8ob7kncwoWv5h3bhjcNhKGYCmmWeZyqZAflZRVOiWjT
T6n0UR2yb9N95F/OFKZYsVmM0s/vsCzJV89Xqr1Jpf8Yy2LdHBpv0zcxes31bP6L
eeYo0gOd0HqICVKFleTTME1yFgHCFBeKjUz8BaQdO09LhssF5tOrAAKn5YTDV69z
uvgyZvo6RE9VK47L+SJSTSOGD3D8gjQltWszlKZXkQbISo0NGPJwWen3zP+05UMQ
GAndpR3E0zADVfgnI48ATQLPZjtvNNLjtqjdkcm66f4/ZZGGZqs4Wly7N5kbM7l2
6jAidovEjVWP0q8pfoNcifJJpK2DGwnlU19o+yKFY9Yg6IPJTkVpzgiUPx/fzj0j
qDz4gIzRuqYvE3gOQF8OfyZhIjpZHH24wgeKuIHtd5YNb/I3/0e5g0pEZNE9lZFA
32Nlshe7Tr3rExcRlAaFCqTUsOaiReYiutr8cO/HYg1R0QJ0h/YyWem5ixcf5aYX
Q+BplwDE+yIY7RdV/JmThAI48MZgvHiK+sYkXHmfmrQYqMI6OPdaGHMKMZ0z+O8A
oCN3Eq5bWYSILBsRswHouoxDEjQRtNnTH791fd3qfo+WEZNfyB+ERjpzu8gFr6NA
PI1V0BvzkbzJHt331o5Vp0uCngM6wOnoHSGpxJYJF5+ivZcakg3+oZgniCIVb9pM
cNZ0MXSkOsWfL0RBUTpjhU5dBH8qHJwclelWLkr8EapQJlrq3laqwPfvqM4vE4y9
1nbf2R/kp+HeY+a8b67aw+UpLnnXMjF1gboM82qdalVCVLeiIWF3tT9oqM/CtBG2
rOkpvq3bAg1du50WhEVOJtJu1vlQwgx/tE7qi9kNFyH618A1Qy4OkwA6lbnzsm+r
ioWBP+F4GFItcoiN7F0wrAB9pN9yfIsGT5W0SSZnryxInL/vz8EIbF/xk3TXL66v
MDZaHYPVHUIdv+MLZDoZut3w+Oewzen7tKJQ/pOT0DiKG4nmdHNX+IPboHNTI7I6
toSbF7KIfsQL8P24WQkGTJxc6Tf27DNBWPBKMWk3A3lnvjI/WzHqlX4sSC2rgTiI
VFvddHMrlRTuy/3n/2237dRn+hJQ+Y9e/YHC9DAZ1uiI18h9a6kd+IUf7KyMc02a
QROvRVnGwsnh1f/gfqyn2mrWCIYN5styxui6mjKTRIwjA+fxyMprw6oCfkc9J/uP
2lj5Zt91Fnd1qwZX/aK29JKM2GjUixTCMqtUSl/m0rhPgYdxJfaWq4/+B1h1QjBD
JuotKQFBRC+vH8iZoty3PF9WoH2k9ijuhFa6bbYf1pIllqfRgZ+50o6iZcMjaZog
ZKiYR94ZTPdQPiTjztd7AqxOad31YOpV+0syJm6o2i0cH0JUU+TbqSq7E+VF/UKD
uEjhtmk3PXDuZ93vkd9Fmwd8s+4b09aI5+0FHLiFBzih+1dSVshM0cieB27Ec3ju
g8XFb4LREJUlc+ckmk8y/s+1jazSmLT4rO5Gd5iXj6YuN56QxyAZKUq6g8ThgAyY
3YV6OuAJHJEo8sAxj+o10etcUAfFIiF4t7SINS9kUlQdtV1nOw4tlI/us9Zhwx5C
JuuVK//DcmiHyabTb+SqXOa+lEeYuP71LqdfrzNz4ejvjyBfp7hFjod2+9yLGATY
ZpAg62BwR0xNQJu+LJ6R2uUT3Kh0Lj3LCHuUsnMan1Ws6yTQ2HrhNNAtIJzGXjp3
CixkI9hR98QLwOEFGCRSRV7lBcqrjslaixsf+t9wUDNSkjwmd2Lci1BVeaqgosxO
Zs4OMKoppdbf4kZMnsSGP6/1vkKKMGLZvMKUiQ0huwXWSNoEArwQyhroAjGcEGbo
e3oHaqv4hyisC9iaXjMTJUQ/VlKcYplavBTf8QWwt/q1gFNoindnZK3xiwNfDBh/
yt9AIjFQfWK/FUaE48swzaFjwTxeAMWiL1m1FXiUbUrU04C8B2AFs238vW3hXCC9
Yo/7GbFdqiC05MMvjqjsw8plU7qy4qICeBEDfi8kcnhF54OMrLVTi07+Vq4A6MI9
ab7jC1WCrXadhpbE3A3dYmYI+f0GGxv0/r6h9YK9xd+Oc24W/KW06iofPFn7tntt
8v8a6jaWx0e6uFtKt+guh8p2RBRb/BcdbcM+PPpDzfxw0Hay2d3f7Wqp3/tKfk7E
2t3n6CaKDeJaGfBZXnX1HLfjXj2uxjMIFlHvkE+lUUsnRjMmkegoJPHygJCmbxTa
LB9f3VJIr7AMH0Oxpd+c1OImv2gZqH50kkRU/jgA3i7dLzukoWo+T5UImcxMqCpD
5enwKxTrHVJvW0oEWR4XmCcLWrlwkFiVG5T2+J7ukbNoSB47ynS2sDrY/Vh1VTpr
F293o4gHKmZUkWz1B9F/GkVcg1PmjL7ZdMauvqO1WPEQOnxmvGWAK6qr+fvJlvus
aES+y1qRP4ZJpI+S4Y25AjCasUFr8a0WJGw2vZ8hNnnRWyihnVEFjy8MYN5/NgLo
1V/bZEoxo41Y4KZvZKXuGFdGbcfgpAxYTMTewnmqrrM9HAzaOeNDkffHf5gn54t3
QBH5btFt7dnzjLucTVdFolsr6BUnAa4O0Hmc1fg2BbJXPxRqeW7reyzuCSU0Gdga
mw/CN5VYOnR+l1UkLHeGvkUqHXqZitIN6AXhVQaPz4ljJi779s892LYv34gjNZro
Z7aQxn/JBrU5cP6unTqpAK8+7nwJ3eER5pxy0ch2ZgyhNtvshwGlbNKNK4YrvoIM
e5FoslppSsM0jLyBCgB97UNp44tO0FSoWzVEABjOtcaE7i6IH0Mp7m/RernNth7p
cEfRg+BnuZ+f0JL0sBsQ13/qW1MZREEzl3OzNA4Nl3PVUAOJ4BGsp9ceF/3d1woF
rHxu2Zr/MQOzf4Hmn72x2lSMAasrtwi3dTjX95zgRr4U699WtvawyJznY3QBGTSv
muayMPw+eVKQFucBqOPPe4ojWx/qJzHrSgmO00EyjoXquglF/SpcZInEtfYXeSWp
JiVjtl+7ibXWqtlbnKA/Wihky4yKFgn7s/XKNkBcRFxJ6RhrB1ZkAr/CLj40etOX
NhQ6t6N4IhvnWut/eocYc/vjLulH5+izQNQNHMbtmMQQY/ceHuEuN1Ysq0PKk3FR
TTiJHwvJWTR74+kPAiY399rk7Cno4TaLJN4clEDGMgposksQcpZGp3OksV31CQBw
9NVvCCeL3TntXAz4J5Gu8G9wPjY6hFXXz3tHVM+kJeqE2bklVL7ScxABwkio1HMD
TEmFYyxv4Zya1H2aFxFS0PQ7w0aIOxFr3QoYc67rkFWJF5FlcTLSF+tY2mznHVst
3BcA4hVAIk15xsy/RJG+G65PTTh7oHiB2aIArwKazji2fPZzM1sDIv4gmcXD5P01
rY7OGoirAH2Ze52IASc5kZrSTij9mzgpKMVqlriW30fCm1ToVPM+LXXfv7k+7HA1
aGZ7pmKACWvUO2mrCxg6QURoLDdMa4wdIF0xXG0tKsEcUD4LtcwNyYdjvWlvuBuu
vj+cZYcyZMlDfJZ7Ll/m11MRGxbPM8AoNGwVgQdepXgnZa56StX1PnMNnU9QEU+5
0LNPU4PWaqPEypEAgu26L3PBJnBKCRc7zhCLastuGwUBewPwsghcOlMDwatEqzhx
FazBscJYvw7AgPfpZCI+PdLZAPG/05ib65D4d3t+aGxhLnEKQn4mISsgovGGCGZe
nnd0tyVhLKDzd6Mzxgc7912848X3w+Ih9E9frdlDBRoO0TgRnUVAKNfSbDc9LxWl
sXkGxdVSAvGxBbayhYg7Q4BuW/y6XB2mUYD12Q+x4cppIU9O1DRUL0OzhS+IKwos
JoN/WOzYXmZ3B8gb8rXgEC+hZY65dSX9G93tJtCwqdw0IMO8TaYk/lZkfzUqnzHg
CWi+yIZUBAg2tEwLrE3BdPuOWpW6jefgNp6wsoT9UoGj/qfCIDRUFD6AuS2jY3Jx
pG/rM2uQkUQeAOFO9SUzWgxnCUTsOD77c05iX1HivQKZc7cEASNRlMkrTOfhh7i6
4ItzrIPg357vBT6q67zQi8ec6cnwmKzBgG3NQnhRs7TkLAogdyAMRP51Qiq5Llrt
JC5M+tlohgfRZ6WlFVG3w9R3cDtNwQBdBibv7nL47twnCCC6UKeS5ZuiHiW2gDPS
t9rys3xT2OJhMA7pczNV/UKfbLNDlL0S7OOxYSOnjTktHnK8tsBOc7M6SPzrgx1r
yL6ykgx2ltflfFnmPzs2s6cQafX8gvrT7k9/TSg7lXiXYe8JexUTAY33GUzOPKeX
VsNCOtjynyLVyHf2Qg1LGIKal5FDoz9u150tyGiUmYKkI0f97rb2ikXTdji1+XW8
ypU78igNooQVB9Csey7jL0JTMcl+u+oTfcTEzHa0T+QnlW7D77I4aTx0lgD2gm91
5lEDlZwggucb9E5OhhDD/Q3gVBP/MSx+umIRjwDhtE7CO1h0VvdSvB8cqYbxk0j0
jk4rztOFe9pOFgsAOIRvUp6Xa9WSADMlA/wEHSF4PVR6UF+MW/nbCVg/F4rBuwV2
OVbjF2G2ZYv1E0DhEkFF/1ORaXQJhRbmMvc/zgo7HDJyxLjAiy+sJa1HxgbStPoS
chBZWbxDOXZCXkggE2cS7ls5BfZBUGk4logNpvAIlm1x8GAIm8FR/yjEH+JKry6J
cqB0UmbbJcSAYrOGzonHuloNSUcrEnRiAqtS8+NzqYKnos/r1X0h3Yc3EJowodx7
t92klJZjlTDxUAO2jOuO17nxiSyWU/R/rcS6K9USwVEa4ubK5VMIfy0dTQ+H6fq4
5la1IGroznUmTdgd51LCL69XpwSylwsmka1stcNVZ6+SZm8W08tJVORK/m764cYT
tavtFnDUqsJ2mqGvg8F1lxahY3fE2DRAfhkok/e1WnPKfAZw5l8UhS9HuYLE99+f
QJ9LggbhCdd/CE1BI3jEhXPoZbpkecGo94oBTIagrcE+eNcmjZc/Xt2a1FpujYQT
XtprTHj/vueBcCTRtmIdr+1ueUwiAv3JEEJ1DI3E9NWMba7wMfQzodZy3noPY3G3
tTlAhlb1lnZWkrSC/j0KxhMmsX9EC/1YljKMEO3yOg2C1rig1Fv5jmELgBZRmnum
eYiypbPCXY+hUzr7gUheAALUiyBYyL5/NGu0VmAdxuhXJGQcjypvbyZmevcwqt9x
LSxTpyg8jra88K6qAWfaKZgADOz7uWaPkg8VEBjnVcej77BLo/h01cb2fj6m0VYu
Wr9eB4dysukkibZTmPgefxlITNZqShZrksZP71IwBhV0nfLwq6D7tC7ID2PJ9oie
oWvwV4B3dlMm96gEGKZlogEtYXWqaE20CZFsScNQzdgbvF400zR6/pydtZGOyYWl
K4s3Fr5nkQg1Pd+ax9zXjGzsQRxIvQNekv1w1LeLalj2MsRMmd2C1Yxc/AJdk05H
nMwmIkw20ny5Z9ovdFpLPyFHpC9OjrIht8ztRYsX2Cs5NN/rbx2PSROSQ9tkkHn+
Fs22P0jSPqTsGGUB8yKnJIi6n5fkrKRV797KUdN/XhxFuauoCLm1uBKFP0MAwlv8
vFKKEu5wAzAvgPHttt36himojV6KQcnBHu7SO8XJJdAWviwoh1KDenBkL0UTfIT7
92MGOv+3KvozbpiTNgs8zeK+j1YkCoF+NoHv5BoYCLb/koulNqxhBVafnAdt/RFe
fC14Ww+OFuVWiO8tKvqW7wuLkA+LVfNzjQTmzXnL5jIHfCBwHq8oc22ZucPIDYEL
e64C+tFsMR1a0T3y2FMzsaXppA3Oi5fStK4WxNmT+GuixCAN/RV4OQ054Qck3cV+
Y05qAK6fSVNoBd5lPyD3ak+4pF/K0vtvca8NrK/5kBV+AuM2oCDSWLq4qHSjYIip
60zBrkSVQVDmpS6WJR8vjwpsTbm5lfJxxxrprLh3iBYBhDzgKBmmmJOUgBeAWAoV
H7tgPMK/qqZCKxbDUxWN67JPUGrvX7+z0JWddFMbFj+UhUjESBAvCvxUxcCnI9tt
p3jq9gyQgDj2xS7zvHVoEI2Hrl1E+luItromiDCav4edCYEmE6vCSLxWGzRmtx+5
Qs+IgP2YfJs6ZiJAWlTaqK1W4A2RtgVgIdE0GW2bOvIYjgHQg59vS9GeP5OMMOgA
4Xjka3In0dckLEpOoYxq5VyVmg8j1Bx6QZgiwt2wS1MKVSYogPqlpETYvso7RBkU
vWjCQROhfSBCRR6etd8mu7OgXS/+iJSh1nn6jqUQtz9hwQuCYS+VKA9G8ZitvGBR
VSBjg+u6JwupTReGnYPX/v71n4SsevRHkvlFfGaemZYhJYZMXhorEHnwXterwyO0
E1ABM/4Nvr9L+80h4Hl9d+xJbbzIImE9c1IgiG5w5f11fVva1bCqKLo6+iAdcSbi
72A5ziiaKWzjNB4mojIlc7ZcHtmbDN8mqEJXcSS2iLgO+GxUSAxxDHm6zrqdyO73
odnV9C9ZAcmwrehI9qtweQFR3eu7iLwS/pCGpedAlI3SLCJdOSBo+2IcnW9OJBfM
w/Y8r8xLMa4kN55PwtEF4x+lJByCacr0fzo/e3TX1KRxKRwTNjdgfqRViT+/rM1i
spG1yzLKo78BBn8DFlnDAnsLGIe522XoWIjZc2Pxl7t8Kh4WyJGR8UcfwxI1IOng
wR7LaObfpVqD8ufwv0ZVdCa2+yN0i+/CfZsl6UAO3MSCClDO6ukKBcyHQLEQHNJc
I0AkpLfqh6rLEWmB7gZAnVe3owHJSuxRCNcdeDPJY4FveMAFD8GrZKZ2U9/Olvqe
TruUWIxgQ5QoC5UdFNS3u/TuGmhuFjzrTotwqp3o+CFKCsTVDXPuus+Dvy4lQdFd
CyIEigKfmFwDmBNNtrQTp+RGinhs+38q1gTV4q3Cf8jDxifmcnr6Umq/HxUitfj0
MSRGCplm+Rai8itPLAuipdOFgK1w7l3XCmq2i1OSCcct3hq5G/tAv8GEeavv+JJO
L4N91Mz3OSGzdwSfk8wzIJMLqktDkKtijWnnc6nMe1zLt/UPBYKfrkSj6vhKu6tE
o2swBIB0m19XNc8OqbN5c4O1A6t61rWrM+7jBLaG6OH+wPKCKsyXDjtuLeQBsHeG
ujrVu8YEmQ8hQIn/ZJgv5huipj6hrouXzyN3ANQ11kNKRVjOC1/WabiIFIU+w3rB
sMbSANp+RwBveNbjaI3xGYt892W3O3Zq2FeUKq5quvcM3V9kmKWkoDscYxxpUfTT
869LxyXbqH3ZPNpc3iqFkTz07hdMV+bOrligoh34upwbbwSEC4KwRcSaTkbTT9Rg
GgA78yXKm+Pu8SPCFl8YE2P7rUbwL8mn5Qqet6WDZnpA4j8YySSou27WWhhll0iZ
eq902bNarvqiRObUAHozn2yQRArI4dHLkGOkyOvAZ4Bf9VK80Q86Q6ONEhH93+r0
D46EEkXAtE088BRdBFXTynAVhhmSLtpc1H+LGMt9nRXKVqYwGkLsh3tTjV3mbwg9
tBv3j/LwldbLA2o7EJSy5ArivwYmUbrEA27MmKvaZUegU/BySD4FHiCNJwbeLHGp
jx8zW3NGjNLSzRLpudtRnlz9NSA3pBpB29TjR5vlxAMPEP2N7G6BHxe1DftUFOaF
GFJnCMA7xePoKV0G/WNAOkKx07sa0gce8NmxOUrlBKj4pOTIO+wBrXtDYtmB6yQU
3u3MYCMPiC2fKZxJZGbRF+ktqNqL37y1RkrLsjsuojO4xha0WFk2JLpr2oGRNn6c
7HB2IV7PyUYRUPRLnwRkupp279Zs2JBBKNa/3cbBEQaoAe0xfiVYci5E29tZRFKD
PDl2rRgLnerXGVa0pyKCC9jAYgL7Aivv9DdRXnYK1P15HCYuuDyksE6gKD7YLAVu
KoEZv6AdAhnvIhTjDFtz1bj9Lwf6tM6qJua8gzF8zT1r0OlIWoBLx9EM9I5yjKQi
w6SzsYj7rSX8oyGfvml2LHrUfapcsIACQ1jKMuEE04S1Bl/rcYE1k2CvGV6J3JNP
BwqbXVa7yy9ulQrUbkPGyaVh0EpX0ec/CrYW56aZiM5x1638DozmJAWlS9B6fHra
UGhOAyWAOIJczdiIFKeTRuqTMwosc0z7hSCiAvefEQnLQrOb1kz2BN1JFVBpuXMa
L3faerH8zkjcbpsfcDM1saXL3dTrXLT+4kWbDTy7x0Bq0FlhB0xPUqGFdG/TOZ8k
SMaN0O2y9pi/eZyryhbHuo9CcuQWcMhoyaOzRFWW8KrDKGpATZeC3uAx2d1zHGQo
sf81f+3T9a6wXUPQHWhdtw+aWBQhkyozhWYf5hyBTtkWfl423MUT91Zi+xnqNcOv
26Qw+HiB1gcSdq1Bvopn7MmJ93a8VzQNeHo9I4v9MKwVcR9aCXlHvfPxk3Kv023D
rCTyqnNloi/ivB8yTpd7sEasDu38v9rTnpGSIj4hkxYp0y5QVyDLht2up13IKpUD
PbbZSE1SpXZbJgDOW02mTg8TmsLu8YLsmq1WsgGSiZhNVBiMnZL47mfRIB42U2nP
oCd9wqCYRfApW0g8JeHDWjlzG/onEBP+84u3lv6AfvPQckaPdeEzdYDXWB9Oto+1
xKjOKsG5ozgOoOBG3/glAmnFDXbh7iU0Povk4z6IMflJjEFiIJ5D5Mt7VJSd0c7a
NLd2+0gtDhWT5DdiMbBpoP72PcB+EUF2jXOmihl02xVX6asTwEzd2Xe6g8rrZEW4
Fd9KmcMcMu6fQ2UY4odzO6C8L6MxND8XmEXGH5DvyP3sqNLg3cA9CUsN+f0D5hpU
ONk1ovXRSRpvc2pku3rci4EUyHPIzUew6cafRs/8cnKtJ1L4xoQ6b6pEDpOLrVMc
2bI8Ubg6cvxXpmC9VwMtFoPzs3M5RKkGBhjN46fC0UgJ80ZSWJYBRshDg/0ccntR
QubZRJhkQy+PadDqM8u+vYG+zAQX5TgXOO8n4pj4mtlGCDRyOkwiouhiQcUpBocw
GA8kOuzRMTlBXqm27oRd93mA2cSVgKpJTkG1aagl5yVEZDPTIpMcBH3nFXYbBYg+
jO3tmcAw6tWWUPUNtOBSrLKWTIMyLyhFAU8HPDzR385PTa+WqmXTp0BGb5JFWE49
cPCilz3jJzFZ3eoikrhpXvVznrLztiaOGgrSvePsyd88gM4WSiWoKG6sD40JQQfp
XDWHxXxTDlxt50OMEfTj4SXI6jA9sOX+cg1/YrziutXoYTYJ8NBzGCanBCIQNnm3
ptFzJYAWDflGoz/Os343Kf/dhDueprnOA5rZOcAoI+aha+lT/slQVTpcl3eziyG6
lZC6TPbDjRjmrP1VpUxxkDXFbmQk5bCfGac01Y1Sblgu1+FP0ktJSncPxCvI9a2y
Daaxc63su/Hjg78IUMYWdlEC/jDV/9uDAO9iSXMxsORUCnU+vQ17U/rwUQXPyeLV
plLyykTFqHrZ1vTjWBvy0V0hpTd/LLUZvEz1/PitZl5//yDJG7aPrec3+a2I4ldf
2Lgmrug5zvEM3PUAWviNwSa7tTZsXxJcDoNlF9RqlCZxJQlZLQdMd08Wu8wr05P0
RJrr20uPc/SeujEGnyTc4TBHTRfgZfoC70K58oJRwzUjxue+jakQMLyL8Wmkuf6+
sEiqJNb8MC81qI6MS6fef4eW/zUHAqJpALURUR/aB1ZM55JAxJAGKW9W23jn1lGZ
k4NczAQI7gHKunAF2BKcGKUIfnzF25Jq795Ya3z50v3jOaDc1XzkdQIR4R8iECjs
OU2bfcGhrdxRbAdsTdTCqi0mMfbGXjbNmQbpqWYe8f3KzRvaqvVePsDXm+5jze/X
nmY6jn6YU6mm2WLjNUKoPOiPD9CUd3mad8GelOIO/uNJHT4BUURtKKbNpRNzzm7D
Y5gZK//5StQN3EyaqSwkznePOhICoV+3vEifoVLbGTOxvw7f0PRQYuJO/swr+f3q
ErLoG8ca4g1u76b3x+HddxuYcp0tTcAcQRr1BM5Hf1evQroFYBI5gLV8vhowwh/p
Wyv4/JvtOjQCOVUiALc7Sk8vlBU42yv9kzJT3F6vXw8otbtuDjfKqrxxN1cUBsTC
Gvr88vMmSiBkglsJUjkgbcMcgIVM+bWl3XlsVRlq8aK5M8UUqpei2h4wB5/x/AZ2
9bm1KZOrroMMVzmnnXbkTue8VPkgAt2jynsu8P4jwSm4K5kaK54CqzI0Bi9QcrSn
4Sdg6AHtZzAis/3TJjej231+4ufgPvsn++Wz8xV5iPvKc0447LFRVIaN811AFmVG
7J3S0zTVL8pU0T1MMq6NuzBYPr1hfv2F23GE/uwu62CJ1IZWx3+cXMgMrULy1sm2
4TKJo3v/reYBdi9n7LFq85uniuAXDRdFRns368QYat3PfyevRAYQaTz3q89nZIu4
OgPx4ABKsx74j5cE2CqBJFw2kCv4112yenZzlyqda1AnCbZma1iuvb2pB8GMkhNI
twr1xl9WUbT0bxDZO4QzwIv4QmMd+0byBy8bpXkuceBMWJbh/69UkZtYXwssepZg
cZYzIq7oz790+3WNlsRi3EYejbqlnPvZEkjRsQ0CA4BSd3aywV3iFCPMKOWps9De
flYNuNWcTjkSgAkoHdMDF1N+6DrQ8Rj5aUb739UfAqyuuSPDcj/gAY6v+A0deaWZ
+3ntV37w83b+214VrpwJSej82xLx9cIlhfJdiBCxYZbLZmgp5BIfb6kD0dDM2XTv
wUyfY4dM/E561qC2f1Ii84Xg/lnVLIBVY4Cz4yWXfp3+9F9OQGJ3auLW2OluLZo8
a+3k6t0DCYO9GG/SoiglwSoZ4KACaNgZGl2lV6QgpXRIgE+y2ymSQNycmcSY13Ad
5FZeLQNTMBvJudGKa55O3YTuPGMislTgnkT140dosC1EI+0ZohwRUerR3lqo/tnK
TPJwiiGaEVkt/bYV2UlMa1t7FjFqL1kLjG/cquN9RdQrLH7JDfqS0Vg8/C3dTYUc
KXe8EdfLYONjjpsbZqOzBSdH9y1/4HObt3ekdCdf6cVFfQc+ZovUAAaGKA9uLEEl
rp+ziNTXrb7P+Z6e9M8n6YkH0ce8/j6LtZ7LKvy6L+5Tweqwbxtp6bTDxRsbzfWR
9iqrGiQLNsucPQ4UV/MNjqjVuh8QYkdbq+glKpOOxOSnQVHCqkQv7c8hI44yqNCV
VxbDZAKPru59/9O+PR79sr2hPzptY4lBABHkWYMW9nznWSOX87TALkYGtezPgRBy
b6c9ecv/gWeisF4Wx0o6KyN1ckDRzt1uJkkzcZdrQ5WFZzp7zFGrSszlHYwqZ8S2
HzkwAONzQqKGwX+8cCyCwg3kRwGunhKYSD/BGiU/nWtyf3l1C2GGuCzKtgZIqQ/U
5AysmVZuAIlUpx5/pwgbpFqGV+YdqrUyrogKdPn/1/Gn0IhDZzLjp7TcfMRRkEV1
pnoTDLkOzQz0qMbaeSrjAQwTbso/ClDHRjPifniL7VmGckEGB0LMY3wxezsCCtga
Drtc8TpHWAPa7aDxK2yXIZIIwyzOb58NtmK7etVjxVXuhygp/sPO46q0HvpaS9vQ
uNeMwL7L8MN+E6rawt5o+6jnhgv2wQKyq1kYHuERDsAcr4F013lzwdNx387mi1Ms
Z4GuSlUmk4HfsSfsDiuHBW0j/CuXjsqUjACQFq4qPstH7ro9biXIzBdkZQ0cumNa
8GJhxaI/SAEJ0vnphT7dOMXrzVTIw+7IYd0XPw0JzQkibyHnWla+HR9jdCfG4w3F
Lck5sC50qnAn35Ua2uQYjyE+Hres79tcBYsvlHHzYph/lQInXGYtYHO5tBFzKDct
ACb2bNtoPrKx+R65BpbL5pNl7+36qByX4C3bsDnYLFmOP0Q2YDGZ8zn5ttbOxUS2
Oy1UFp5Z5QbVKjjuhUyJyP/09fMPc57ECPi4OBJgZ4Y0c3d19MexL7wUktlCoFDp
etzKdNhaqkjIYnUm4PZI3/9xpdGTPc5SpWFKKnM1DUE+xFxv/zca/ofkbIVDfaIM
dBLU0WDyJ+EOLJEkVhOxr7B4kndqTWL6B7OmytSL7+8AUv3pOVGRoHQJV8dhYcHe
4RrLnS/mSmTPz1y7/UmYygLBV7E1e3FkrQ1f6g+hpWwKwPCm7/Bv4CgUoRHJUXpf
0222CpVDDx/+RYHjHaeCQ7Td+mptALIN0ymMgzZdKxA3N69965m1W8CMzhxIGIJl
t62P2gHvOpEmfP4nXEHcdjvBRepqr37+7zk8sLHCVJwiUc4MXsJwXPbbyfOP5nPs
dVNvmnrF7L+MgIL87nSg8/ENbmZiSfu3U5eZOUowLrDPseMk35OCTrpJMYsXAUWF
MBsSef58W5YQV5wIAgbxLNOlF2RqZrlezhzNDMzMlHIptoTPh5LvEZViubN7HYCv
TCn20YvpBMq7+LuirP482ymXQtLgIngmekx1Uybtc+/smBOfE5pF2U6r+tQXOXGG
JSKeVS2y4Uf4tkfqpWmtNqzB9xx8yOYhEttEpRUTf9E8Bf+reYVXeQ2q7u8GO83W
oDy2tIryaomm562l+QtJiH8JGVlkHDy8u5ZX9B9MQf6UUAxxxdAGbsNnAYo8Bgol
hVtbEr+3hvok45CFm7hZqAw90gUiBbLgDZ1ZRaa+z4Ki3x9wZzYAhq0G4nqIUX7g
b3KNKgjqb7vCpapWhU/96GIsoaFAMuXtWVBfRGJ3YJWKXpRGLg/+z5CCn55U6Rc7
LrElcIluPdBq5kvYJej3jJxnIPCI7toeXRDyN6wn3y95A3OUExj9bVSQhxr4Lphn
L4nLaAm44YusyDvMrVrMKWJGvHgsfJLskPXS8K4Lbyn70yEy8ayC1bRK27l1A8sd
3IXZ3XVNJ7gff3A0qWtJKw3XI311C8jc/iOA4E5tGwNSN+t4D26jfl5CxXw/tBX0
wXjyPHUiNhCkc6SgZ/ZxxCBp8l/Ugp75tzKVmbJdMa08drtIjBsbdzKLkczj8x1k
2XaOR+VHNLPX+0zdXG/ILf1oAeoHaP6u2FCxsd793MZUab3aSh9YW+IE1yWAzesX
K2wVa2w7txivyVLwGKhXjC7Xxb1vc+xRX7s9+o/3XdmdcmAgKCNdg0n0A7F2sSVs
q6qbURfT0Y5XU260u3zBQcjnjQIEzVf8qjW3FSF5nNd2qMuiuDWg6Yz0HYMuzwRC
4hHz8pPb8qlYPREIW8YqwfJWh9GVpZd6kn/Ou58lyl3XAS45oTOb4syT/lL8fNTo
8JJa/KOVwWedjb5Q8giJ+peXrW9R4Q7ZFTVrhzRXU6CTTFsjMxZMba/mvnZehF4W
jLEb6n6I4dBTfz/MCqkVg1cIVD8c238AskET541lAzZ5ucvfHJlc9TgWZlC2G9u1
hStmoDPqo4ziKZrGyNn/aZ6Q57kKVxgnBJ2DaHG25HrITpp9IPmnEBaBe9ppN+sJ
ZMd22xFJh9MTJmsyEXqYui5nKsQyMgQkv72dxe5m2hvncTAZTQDNzTVgH4R3fMLO
p5BYXx+WjSdwmHBN/pvEPdHdwFwbaYL/zjxqBzazL3htnGqJ8T24K+3KdN6a/sr/
XcL/rAd8jt8Q4tv5a8oUQpFGtABeVQ1U7qG00O81IeLlUZ3tImbUAbAJaxEykQLc
5VJ4z7DPE3ZED/4QL/8akmz0LroXf/Lj7FGDVxCa+2SZxJuP+KlfDIxEZ5LHbom2
fFFxBUZNA0WgaZ9CS58wwexG52Qb418tqOyd/XFBx6eDEhuum613tMr+sfD5NoOP
p43z/rwcSpk0hqz9++QVWlWODDVW+nmOtZnNNBgVOwzUQPwPqjPJh+c36sREsajS
oHftUsgSiZrB1NH00YUZt7iE/zG0L9F1GN5zalSvhuGWnuEDy7LCLXRun8LN3/Ep
sDn66hy//y5kX30izRxXtgHQtp26v0INcAH7yI7Pk2+GAA4MrRbZIOPz20e8KpAS
ObKZVCWPxydhit2QxU25A4nVrpP27i3Q2akqZab6rZ4tcNFJk+m98mObYKS3RdjS
Uwd4ks5yxmJVtiB7mskJUcu8Kyr9AvoiNUogQOGtF2ctT/3YA+1EkUpVeZun04mY
U3eFZG7f82dwiEAXqnfmSDJYWUjeIt/1+2OrvP12cHjtLuZqFy7F4q2OD7VTiGAR
dDo8vGdCjh5FeXYLI+Yj3E7L5eaJsJGAxstsUM+BQYv3RkfmkQf0mW6l0BfIgszk
HAb8Wp4rc5/DImKV/YRML9dgkVFruXTBki3xT3UrLolnuYz2qgNV6+swqrixuqVQ
WVVENDm98cUqSuAcoUhzNy4OZeXzAsW2t23ZHFbNNB+/9zFDtzz3zoIYtvalIL9h
dg+AI+mKoIWQoZYnL85nLBIg5/EX99rYD+xwz5hFpCvEorY4FPsvmmCglKSorDMz
KC7dfiCh4xQ1zcGxUVAxYfimkacDWATiLY0cU0PkUoo7i7AUGLVl1Q0LnmJQG/0/
ZqfKYSIErxpEdMa1OdJIcMwGv/UUiEdxIh+UtXiWEPFwBjIV3B3niYYl0lNFHQsc
ohppbclZCxwR5osUTlLJMtkQ+VQXwvBffT46xEeo5d1PVHTIE2lXSSjSgSQnQpLo
/PIGugc+T1DIZvf1kFqkxVFmfLQmB6nMJ94Gd5Gu7rx4Kts3MvIrYA6BZvRWu+Gl
qESlRjb8WRNwLf5aQ9hoA53S8eBtSw4AKAF8Djc6zjV/uCFu9KVictNAa99t9SCY
X1VFKQzfRUwyAOAlpe1SZPMzcr6FGXAoapFtpTLygHhr2oe7SG6kkDRnVlnU5EIQ
+U8dTdFbAaGf87a50VqKn7QDgMdMmgWjEpeQMC/yH30ix3g5WE+d2yksvFx6+gbn
TmIwhhq35WQw8gyqrbfUqlwNgZDMZ/OqtS5a5/4E8W0JNgLx//M/uvU8Rtj+4fVr
EX7cH4WIwHag7gOSI0ivrizSsDfX42yv48J/YcRZs2oTGED4dyLTkShwYBmIM95J
579C+eXDpPm4uZty3dnFR0mU48jdHiN1ZIBI8vPRuzr4NGbOnCCto/MZwgDw5ZRL
+bXmJ+hRBWwAHVNOgFHmfXAstDDpuTTzMefP88IucO19EVbfQh+e6y+DubDa34ez
zC/iJCrMBldM8RRixTaUIoNd8/YG0zGcwse/+6P3/HDGzwYH4bcvPd+/AUA+ZJYe
aiH8QF5CtUfv6d/f2/CKiza4cm8Yty1nqlgONHh6NEvWyn0OK563Iq5Sb+X6PZ0X
JuX7K9eSnhwqTs7Qd/masSm76/pP9wn1CL56pGcnXr4Lfch7YfCRRSEBK87kyPcM
A0xBl32qYQJpy4I8L+NGfrbfenBJKNoh93oX6NHMWMYETUPNsr7RpJ2Hdigfs+1l
khIsv+VzvHlU7UWSi0T6JMf75OzRRWCBkYCSZR91HYVUjloQU6sCasa73IjVa88W
foIUcPjuPlNLEuftHoOn7KAsEFiAj2gb22wLZLEeV4aL4tBmlFBVX7TcCnTJZaYz
a3UrRVLtYhWzJfx8XufBg98sgGB8VcHVztHWvzQ2hwu+cL8EPEnfC+jeh4lqHmT+
Qhs7Tvlg9adHmdXXvWb+aOt/0mmQVDEp41mxzfhIIHOH1G4XJR9rM7bB8YwSpXVi
4YzfaBd6FbxgWjvFvvlTScS6SRRwKc9ofM989WqiAqbGM9CjG+Ao9iEU5tnglavu
KGUN3LEft3vc0myU0GHYSshmNJKgbnUnV9Mt0VT2b5Tz6ExTmp6F857L5tfpfJMo
tJVxOzLbClLGEFqsbXnW8DtaR9EDVfvw81oDFU8EeFf4+l9HWxnVnU9Hfgg12sZz
P53VWf9EQDg3cN36KEP8IlmXcyaX3Kqow+/e3JalXmE9EElj/ikoCDTST6zv3lJ3
rY/+91/jucP5okem6/YOlsw1wTMjfHDUtyLiEFsVpFO7eX2Aya9Avq1YplYVG0IZ
p+batZdiginpvDFoOAzr7aRtuzW+XeWE166WYqSshZKAkcFQ3VUXF9FGhgjOUeQc
JjTza716YhGLoOKXI7X0r41XZSD68d3u8XycrsnmLBlSkJoQYx46b+CXAfbkL2SC
zvnQQOuN6Va1h+sALN5aL145yOGEAhUQa11rL79d1+BLPDMl4IE84QXOpLGll0aS
lwPZ/L9Vnom529OjUMuCsiT9eTAZqHEYohSjUPXa38UlbJqE5nvycEosNG/SYV8G
P07WLOxt0N8NAS4qw27uL48WCIC2vBid57K7yqKi/FKjwRaIU8LgfcPhi4RFDWY6
X74oQ1Jg2aeTjunbopIsn4HvcXICDSwj+2bc1R3NaxLEDNEGWa/YI1ft50f3VnYc
t5a01ZBS7OsV2b+6jDsY6ApxB1YeJM46z5afgD6aL89iRSlLtSF1asgdlwlHIQn7
WTtC5SW7zKeLefHVfGr4wODUikqR0WcCO82wghm1HP34k+pgP3XDsdqsMRThXKcs
E2aFnwUeICw593oq09LepaaFH0O1wUUnojh97Q4ShqZWOR06Id7/nl2j/3e3+gDA
78Gm0Q50OfagLu0aBTTYZFBvhAhYsIiek0aIWaNoAOoDPvGZOeZ7t7TrLopN39dB
Vr3EFcZTN8vnjM6UkBaQd5c2B9hh2DdwYMn8L4Y5Xi9oUKlna/rf9HbQDHSDtUPv
92xLMHYaOVM4cc2uMmAWmII5ogdkjq91newbzfFK0xLcZTtfPMzIifgg8TYFhx1P
2ik8UyR+CQ8j07yyd/6uUVZIdCP/IQfJQezYfKGpOTJTOvhGZXR14URTj4ZPMiEz
autrcdMqvdNzI27DwEGF7FA92vgJ1okSsXWicJqj3ETIUUqjr8nIRVVReAeRb5O/
3ch6zaWpW7hDuKhZQ2UN3mBehPjr0DPjAVJcByqqKdn/2/UiKpJPAxyFlRTyg4sA
5nYmF/Hk5wEsePIMYTUSFW2ChwnCcqOdAYrHw0TXp8cbgMbEF4bWzJ1TmfQnVSTQ
dbADtIASMWxOmdmm09dmWnHdoIganRf2vGVGVGZDlHgxmpq5FChsOelu8i+6AKzZ
tLEportRpNvtBik4Bezq/H7nHVTbXU6Pz+JAHl6g5mf/11jgqLSxwsAf+8Sq8pYd
osTbrnozvz7qCwvBR/OijyIjkNdM6kuGWI0fqcCIZn6jLrmOcnbTj/cD7PmrFqhX
NMYkUpw3MjoJhseZvaBd50jqrm/0k7s0xg/za6gUJf92gnRos79LVYgutFKkvXmO
ZLvZh/ATRhN+nr9x3VktHGw7GyPfPGtAqjldgK3H23Dw6wGyOK70RZPd3nkt6isG
3ypqCI9RJWUI4nSEOCH41eUrdYNSkNxZ36t9lcUVuGP4og0nXXaVwxEHV2LBMZHj
ZJBWfmRODceK4CmGdxj6w/Pmx/IhXdBoKb5ffKnsPwl95rS6a25cDvHFW0UeWhOI
S9tzjn6syx57jKNZ1KsiVNFIXmXyy2bH3gUwbkN8MyH9x3v6SUnIpgz5qy7nVxFc
IFsNmduhEopiUu4QcuUaR2B6Qj1nLpp1+Uxs8hKknzcvi3rVk3UP/8kILg35tSgk
4+c/b35uFfutWs/qZiJgNe9LbjLAK6QrQ+B4x2KaAzSlDQzudbRdZ8uw8QaX9yT4
GZ67Q3uemSkfYQ3LX+fDmXxZXcfmVbJ8ocFOcmNGjtNkzL6vp5KyMHQhemHkD43a
wJW7ifXAiQJqQ6p7FwKgMHpqSqYysxtD5a7JJGHWvKOXH1vCwlSymU4If2Q2JB20
72Pns2Kskeeua7mg8nCpt0HFbyZx4rHEfXWlvtBALB1MaF7ErzFLYa8bpV5KmhqT
pqDq0uVgzPSinFkYOBKEqHgRUhwZkmz6lq2K2VAe0gkMndt9e2i/CV7pHT2KYB1w
uEQpt/bIoyX7I6t0yEoV/PLEZkX8w3s9R1RnN3kJxl2jVX0zrt+1c4dauM+XkPma
WxQbKzVhkKjEe4QaAc1LFPHqg4Q6x3CpDlyqPATDEmufJjQjKdcDXIIGP+o5P25/
qOXbPTPhMDe36cJoRQ3UfLZYuz3L+VWeP2rJzc6EPaPsLyfRI17bp/hZshDaipoY
eaFDtLwd1UeQ2DpNDHKlQom6n3Sx5NiTSNnLKqgdkYE40naH7HXuHT0CXzHSC3wZ
j/aFEgu5dKXRRKRiu7P7P1YaFG/V+CXPv/85pVXnAZ1B+spVs6O2sSZKXZCN2qzK
VqiPs7wTD4OtZXqILbu63Iu9XsyVnpk8NYdaggd3aYe5fSq8t6RIMdWGb7ZNR9uK
OtkdUBZb98GUGmdO4T9wRwlkPqA4eZ3XmexAL6+xAGJHx10D4/VMwzPOh5JRxBY/
4w+66Z2SiKKGqbqCYWkBZlcxRsvh2Bo6uxU4LQs5dsGmN/l47CPX8StlEK6myHqG
Cv98H0dJ4789k26z8CsSLyHiG5fXhadehCZ6QZcXSnDEZS+zuuYX6fHLG3Xeh+rM
YNCbjkeZTN3n4fykGhXv/ud0eqFW4j/b11tcmA5GWbQYxIG91Tit3uxWIE/56MnS
pTgA02DMLAZ9R6zDYbT3LWfDl6NWPcU4AIR62Pf35iHddZTM7yyC56RtrHq/vFXA
GDTkkl7Bd9fhV++hk7Rzr3eyjvbIGclGuYDnuBYQqXcHABezmYs/VQg4qYg8fVaA
3QpdfM61H6WeD5UBy0n85mD81gLtcjfh6I4N3CRoYM9tnbczsdVjxHNJGdGGuWZ2
Wtr3yWKSURO0y7hNkJBTQvKPjk2mpiCLMk0ycVh57u7CSDTPgiS++nBefVik4Cd7
SdIUYnXSEuE0Qg17CdgP5cyXDRPfSTFd8GGYhkfTHHDbmgxcVJ6XK6bfwPEF1w9W
PpXngUMfi4mdp+uDEG56Iz6fYYUTIrf8aAWtv/4Z6x+pMfakRgoVsREg6VTc0prM
2vNxJk6USHiZcyBQBpATX0TlYlylrleCyljTHBWFTXK1gVP414RqJWM98QUnydJ2
SjqNoL9nu4rkBUBBXYW6AhcJex8cphNgzfr5ncc1vF5+cp2SgJQUwINsq3AygxbE
OR849iKTy2+E0waVOz0qapWE8e3QoBgq2t/08yvji+1oo8UrcLN9/l3IMeNKEKLg
BxI3HguIAUNNtY8FCnDz8BVhAuW21Bz2WUFghxIYOPLaAL3Av7R4dVRAaPWicJkk
7TmHiCQDwz40Z83syPssKsCiI3L7/njytNhls9vvtnRBo9yFuzHYm5i5OfXKCtVx
aqqc+/AAYhkoisPchHxvdDDwAHFOK4lfD4u20GNaDAKaiyqN+6mpDIN//5+y2AST
CAWtoersrDdAYj5tju3H3MqKtZA+Ck2uFgHmMKWSZkp78U3c7qik6ZvFF8dHYw4/
/dbDFTx7aIYsnXNj66neY+XAL5xg8ZDA3AlMDsszzwivXkHlL+VH3K/rnYqwLhqA
hnD+9MlBt7Ho9bWrdKHM8tQyXBXnQ4luOeF32OAXFgSFUZyy/Oi+UidSUq7QRlJ4
corBl+0gIzCDx9o6sH3K7Fld2Xat3SQLUIcJcl5gPMvcz5HQ3b/ByyVGOQmI76hA
DD5zpE66lJ/gYAScSHfJdBPwZiON3DvcxfC92HaCgqSOwksounrgn7XR17YFL4Rk
J5ZHrU94bGQUgvuarqUNYyUyjrzZyTVEA6aVdMDhKLe5WUrNdx16RK4fHtxa+/ij
i2TzjAUCq2oIJp3je769vB+cTETqfyHGXt7VzBtk8Rqhg1X7q9ZTcu7luXFF5d5C
wSdOLwhXAdSyiZHwInT/IPFP6zlCzGcQkiQFIIVLJAq6CP4wY3WwY54ubVo91ltx
pBl/CYqEUDfOBHzx9Co3cznAc64+ibahCekWJ0kQaq5SJZS0JRUrCty3LnTigqfY
F1aCJMgH5wkLmWjveFHM/VC27pWtlERdMZuP7ps4Wzo984XvBf/3H70OJOy2tNl9
Qi0fRnv5f98FNSpfnCRpj7GVX1wERd+37V7XV8jqxc6ljn2uwVRaMrxfi1uH3qZz
2IOAsvyOO5vzfqvpLK/uoz19VBIEqpQuFRSpJxrAmvgVBJLBU1DWJ+u8DBD1wtrK
r9VmGvjN+BhAgI4H+K++o8gEKGdhEijWvrS9dcMp974DJiJeydeCFO0X4bHxRbno
0qt3AFmgsOFULBRXZxbj6i1/mLZwjb/EgjmvJNQoSYdBGROkxhIPSuAr+QGqeQRh
GYb2nEAEUhqfZW+LJ8QXYj+FrqnQJcv78A6qoJ5AlW9itNFxkJfmJCgJFHbyrf41
ZVeDcXUwjutCsuzWqyNxxXARr5HQJSH+5MHm7PJX4SPrJTu9Xhpu+EHBYXJGqRNn
h1t31O7CIidhOyWdjPZqnxYb6VbyKmpoEI3u5HFsYL69afEPvs/4F/g9WxEzXTuD
lmHlNLnG07vVEntIzEg+1t1VvSTlljISJG8Q4CaDDtRYh2l/vl2G0juJge3tdfQ1
yoLo3TyUB/dJWtcmaJhQGnZcT6O8+P4rKNhnACTXH8EHxOXnXIt2g/rYKa1lhYje
+vXkEj8Pd8pG/UdjymnNbZ7JWvrkO/HTznCKIOdqC6PoAitSkFVzpY8NE/EYfadh
41vrsV81F7OTlmzcInC24ksP0geAYiP/Y3XhBeXHS8GEgbWstPrVbf2W3sfNFk0n
NEF7S2qCHzULcWjXNh9sLZJMD4ADrvpjRdHmniRr+DOTOf4I48AaYWPqpk1ilaMG
fErBbXMVAyLa8vn6GSBBNajIVXBjKPTD3phIKzoui+sV1X9cCmypbk0AUuKCGpIT
VjyX3u7WrGkrMi3mboayIXF2KShjANuKE6Nh+zgAlkCI37aGKZ/7kodMa0IsladG
nB9XD0wgRFbdLrPeQrYYLwWDl3Q8PWz5KNZlQkMZrgrNUipCyZCNKn07k+xy/HBy
nhkNQznvfqfHVNonhd9rzlQpwRd4loPzRK7M9gZP9FM1Wc1Dt/VtiK6ydTCx8Pg8
GrxJ2nrqs1PK6i+GIClZjiHN14Z1O11XJBKY82grWkIV8Dp217/2tRGxvlzDK4fR
wI+tUqqvfLdVtBDJU48MgVrW4tJuV6F0w+u6Aj1fM66XVMIJOBi6N9APLhIdepeM
etQAZuY8LNcJx4d2vcoTTLuUmHCUlDOFtLf5+iHLhSy+akEPt2ugcmnbny3+si56
ykTxR5CKGX7p3oLRYNZsjcBQ/05kKS16ACcYc8WfV8xdfrNXUw0QB3rpPGfTipmx
yFtsuSQiUlUPI5jQJrVbgTVVcR8GGgEn9Z67jcM1Ig9BwiQac6ZSwst6A/rsPIUN
Azvxs2wZ9qPmxs9ZhNWEHBpNmQcrN5619zv+fINw+TgGNVeXd1jSQ5Xr+HYoSxu2
CFk1NDAva2tSeckEsCWyCDJfTrbGFsMg+j7dVpNL9LtwVga3Gr8pUMBoW1nmTARs
CMf/Xwm9EZnXSFn37CkF3NGIyAYNBZ0Xv3wVKkKitCjd3xUwe/LYFKYN2L0mp4Ep
6uv0JHNdY7fUV96ZqNf3NKj98fvwrGaKwJ3I7ISkGEXx52jc/Q6kKJ/ezQcOoG8s
us3Yrf8N0cROEUrC1OnvZzVVb9X4A7+jm56SSnOKu037Ya8D42X9txkezw91uyjF
+3q7HZXhL2YW0L7AqO/OzdM0rYjUhKjRau/vLfByIdpkcbik580lbjlK+/plyeXK
maXjPTO6pcAu+HwlAbONGpCZ+Vc3Hah0sOn7QJIQ8Tw++lcZNPH09P2O468n8+WZ
QGMWkn5BZrFxsZVl3WFP7Xs0+fVqY7r+FNjfDcmttN302kQOkMfkOLX1NtyFGwcx
8zgVk43suJWSvn3amiZ4T/DdAARYM5DLZ/fXd2+Fsql/+s4yQu9I8F2i+MiXYLQL
uKSqu9/sOUSQmkLg0/4KJP8Ulk1tR/Rp31ouAZioXupFJYsVwJvjcEIJLsbqZYh/
KNOlG66GDmGtixV+3p7YCcMwkTQK5aRWyezFWbhbD6Wp+2JmSVJTKGM/jqKGMVjc
NY3rpBI905K5P5Fj9KhPcYSoM+Mt1vMSqVsUTZJeSnvfdb3ad8YmlULgcTCflDLN
Q8Kt1zn15ZYut/tlqsDXaBi1eWve6gocU2VDigh95fJ14HgMflc2SAuUOvHgjcG8
lpWC6asgaeKZKHZX0biLzuYsydkHGkGPUVgKWKQk43Pjxz3AQdsCpPNGhmrqmeyg
GSB6iTVLKMtDxFEA8TK86iKoRTagFyeyZ7W2JppitalPWaX7Bo3TQqysCq63hA4S
VhkoZ/1CLhzgdRMxHBM0A/n/I3ZokWiSJpMt9BcmI54TFBrnEPf811XY482l+j+M
tuWDq7Ue6pVMpn71Dzm8KKEs/JkjpdEv3YIrfO0YeT0XgESAYe1KvIXJvP0yQpvr
EF5w3M2f5zw1eiVt4tEA8AAGLClOucZi4g3pOEA5ad6dayze00fqQLT8iqzdx4nG
5JyVj1aQ9UdBqOgdxutQUhSrwEgXW2kW9w0FDlrCsR+gLo+aI61sjBICNhzHnaqe
bP6UMA8zBhWIP6Ctba0c4QAYQMiDktyAKFfE9idfLEZDNKgXnhqt02bGNRM5wHPo
nzuchbqaEw4H3q+FONWX8/nyWtpCb0JL3VDQGFAGYwyAGrj5SapIZs91PGVPsX1f
K0DBHwZpq11NJ1HJbnhkqfLNk3eCMaoeJ0fLWtEvnQmSEB3RK5EzRF4K+PzSV0Hf
zUKnOJCURUpaMLqJ8KkW+hb6eUJIM235wN5ERt3OqrWTNNl7tSL97mBucD5cyDYx
KaP06/WdmIRNpiaWXL511oSApzKJcpkgDPkHMptpmTGdjNLDNhcVxmoiW45FAqzl
qKT8EOPgLaq3g8mI1d6hd3Ab/q34vixbjnP+E+2rQwfBZWCC9z7+TvXENV57MiI0
yW/WLk39TuLVceIrVMmfjTj/QQdu4ZH6nuqwBqrAJjdofh+EkssqBCyBePH/t3KL
3gvZIHNUQjqHM4lmAJqgbDJvJPAZT8GWRcrOToK0sH+FRalDpNtFqwDLvgC57IFR
yHhrX3XbIB5C9e/d3w7YHlkNRSMJAeFaj60X1SDQ7In9EoNMNFdHLF+F8a5pfSEP
wggn2hjOXlf/tfihiOZCmYt660aDgduheidWUYpX4tWkYvrgJokWsai521FIPJNs
QBDldhIYTJDJfmsV/VZZ/fKfaQz2i0GnOMYMaQv6DIX0tJNwjcrew0BrFReo68qk
sU9yofWswDtOzS48nVL3UpFGi2sSkpXzXXvv54Vsdr9wjgXaUFnNkikaTklBMU3j
XxeNSvEyO71dCfbTEJhMpYXLrC+omntx3Qw8QF8rC7ABpV2w94Vs8v+YonRcys07
HBsCjZbW1mwtgcDTxqEEeGIjU0x/EVGAu16buvpvgHY/UZmJsIezETHrpBaEoB4y
NNkB2vW2hhJoSwHKzJMpZQEA0SCksIXN+hV+sfoWa6VrdqpECN64uBLwGDs/gjB+
IH46cYO4jFQxOUpHHkBjs7qv0dYUvKaJNrJy1PDdF891H1MeO7nz4T/CKSbcnb6g
RxJ29GoMDRJsT/7kI152nzu7DGnB/vQFwIJpWyN8V45wJ2LyQhOdPxG+TVGXIup/
KlDqHY5ZNn7liRl07UWilSW0Si9p27BbrdGCMs20qH31IvtDKGQ2UNX+iYH+aEJ9
VL0Sxv862gSxDzPPSABwsBKoJkGFt4s7dR07on+v+uW3+9/qnO3+2vlZg07uIarA
VKLC7tdTgdiA9b0k0pCcYFRJO/B/3eg7x3yKz0XWyhPkzvKudXT0hJD08MLECgYq
idyWCr+RmECw17nFkV/RkPirvZHJNWRKVdvcVX9d/y2crGth3fHb62uh83SLJrx2
yCPv27KhafyjkPg2lO3bN3PmaBRvN7g3x4sxiE/xIwWciZg/16gi3NRrvn7G726e
4yxvIdygLN+RzO7/JVsANX7abW9U6pQ3ZKZEKl/WJmRzIbtp+8CmZofuIxXu6qLL
IKGvEwUe+tslFvYFuSbUOopvajz7zozv/oiTJS/RhBI5Og6WsP1kK3Z1F3mCMsVp
KBt78JiONW/v2igpVy+mz0/ujoiMgavd1/3ISo8rzfw2dKYsibuFe+esjT5ofRqR
oFdJKkBfhprl7UoLypzJArpQSmSypN0nHuuVDPhfBrYuUVxYTn7NjaYs1lowP0/q
FzRENVbe0vHC+0EepGoKodOFrWHMNCeQcum45x10kpj5wxXoDwdsPhrNiyZcS+rr
mAGMf9K2QbnSo7rhdkdoN+KuFAHb5zJCT8IdDatTGOFXtD8Gk3ZvNWnrsLa1VeX0
tU95+ueqV9Pk4UkR7CXZnyAI42vsluj0gq617/rP1NVTLvAm8sGoEVMakSQWNKPj
m3Fg3JIsUDapNXY88BGXbcWcfWHZV6zFj+EDNPuccxDPonQncdhqWMqj8z67eBgg
OEFnNcfqfiXeWEqIfxbUhjGARokKkrPGd5nFHiVZDT4zTVmxZ8/W35tZ3ks86iZC
B83KXuWy6s9EVUASdMbDOzzdrxUV+a/gCUJ8NDYmBzYHTh1Oto1863Ogsaq2QsH8
K2fu1Ki1DlQMRQ4SQv7rbSCc7VvgkOikncI+YYX7xWp7hRP9OPBTbAOJrl2ydluF
8PGZ9g5W19A7sbw0inBwX5jqRGqsvycHkTB2vROVDr1UqYhZIAfMEujYBjkewxXM
UqJcKWXeQOhZ7vlb9obUpXsYSBxyc65XqEgHuTLElJpyXs3aLr1lGqUTpwPnPVpz
YFRvLokOa3NvoZcfqYdSi+42tQR5gbesGzH0BQZdHb+Xi5UnyJ7Do3//FAGgvPJr
QrOh8JJzS1gLwfd+igMCTOtaxw8iO0EZWsb2SoVEgsmfZhp6F3Zx8rwRGnmYx85e
6ecS0EZxdcR7SpCYCutSnPw6POEzefc3PUI3BtfOte+3AoVLADfzBvlIwjf0ze6F
zpcD8zr9C2cq71BawnPBdND/9QINEqGw8j+JluaRcKAt26XEWoFDyeAzJVkE5E5d
KLYnHYHugiS31qbnXcwnt5/q3vk8sfkdTQ9bZr+Ys5EUuAhWrMx65BJvJBhj8vC3
2oeFOYNP+bhdXsZ1GIctd/zgay0AkRVc2JbdILvhQAOPh8ZIwepuOutzBWC9UyBF
J8Ng8GfL4R0O214hUbSoL++n2FvJT6vm3iLS68wxoZY8vILwL6oOwh9Jqx0B8sUE
akDbHD7qPjWaWm+zCgNqKfhzSjJgTQuVIObaKD5FJ7VCkhfeeiuBkRE/Xe4em677
Up2XOsPoCP5oLyTXCLSG2RyyEF6WAn8A18Y5XRSq519MGq/E4l4t6ZjSFpN6941g
DahCENQQ92GdjR2yqTIK86z6MIuOECsiAPsulNaCvTID+3S2/sM4mqjLd1Te1djH
cgaF2LmMyHsgA+kpJ23f7IhHurnDvgpqKYrQf3XY06vy7rDPNTgFIVd+JzJ+Hwdt
vfjpMg/wr+iX5R+lP6uJmu6IJ8P90lC8IffzPtxcdtsiuTZKPNdzdfTjb5Sdt37E
/N2WiIi/wPrf1INznzq7aZUuADA3YfqKxNQpAqTII9ECYvC48RAn+aHnvhgSmKD7
/enefQOK2t7soq2OCDhj51mT5w5ZXs2nFhMXXLXl095GZJ4ad8ZOOCiqoxLVmEuA
OIWoi5Jb0mGadPF6dD274Cddk/4945JohI5gGcSo/a79a55F9BISI2tpGZ695a2m
FYBblxOgu8vT7ZyllA2qKKUJ/iz8LpAy9VYPlJkVM70nvfl5RcgxsWDCXf++PY4c
OhAIHXfzKd7zc3X7hXuXdKhKQfGNfQEeZQifEGj8z0om0HdGoEzQiSPIgsmigLWU
hXAnLafHfoTkRGVR0Uz80rYylfYQs7se14vBwghQG1jB/Prz8EnSwidUsWoYx9xY
EXC5VWtLwa2oAxEcpgCn5F1gFZJsJ3ZRmRWg+WQ3PXqWr7ALFfPnFNQ88jwAYNQD
Tqs/U2FjBkWneyGEecxKk5Ufc7ZfFCazm5IRIt+6lxwr4aXViMn9boJOv1obDehB
I3KXsLtbJmsxTEXPvigxin2l3tHyVHAD1Bu0CpNfdmG3GRuG5GvrnlWPyh32PF0w
mHlKHZpk0H2WqYgSwbed/3W+W8fXRVDqEyTAfC8NqyjCZKiJDOM6aVfj7Rap3epJ
cGIdN4Ua2uq108c1OCj3l2O797aVtI8tGLHN8nQ71o7Zfx6eo2RZ7Jc0o7aRhoOb
ZqveK0nqgBoh6Mvivd9gYqk5HqstlTby4fr/6eCbnnR+pw1pC7V68c3lQa8KrttQ
OcQrj++xIWiKLTuhtJEZ75gjP1xjKCQ0+TjmFop8T+PWO1sQ1mCO1ZOXXAS2H61y
5mU9J6ieCGukIgxysVEiMcSlj0mIGwTtIJ/pkLtYjs3MhOsXHxFJcNXx2ZAW19ni
Jcb6Z986xPJJvtV+6oIQ3hi9R56Qx+DzBzAUR6NeRPiQrUhahvA5OoRhDT8TsefL
+Zh9ITZvJzW3nL0RxD4F4aux6O2tg0OxfUUJjLnTr1Nrx+E5gGcuVvh8WHPnTaVg
lDljsVVzmuAJV4vPHWnX8NEuYyVhfbuw7vNS5WdripQE4kRC5cXY3b55qbG0FHnb
Dpdy6hBiHXT1qNs2D4Z68mTXAA3nzpgf6p+CA9N/kSQEdiGMUyIiY3EgQFPt3maQ
fwitP3Ddk2oOWGeX7PXRIkwDgoTr9vOR1olnyiUDvNlFZ2OYrc/jJfDExA+ivRNv
6f2p7QXq3cqElt1NTa2GdCmI2IHQKdRPYiNfwYsAhTZN7iE3GoohpuHE3ogv9tW5
1xvj+GLJ+PREH6cjS/rHoCfXcPLF67Oik/NegJCgYnJqcvoAl5VvqrOXiZoqEdWx
4uqRuKFb+Mwh7hnWZluBLv/L+U7t7bwnlSsQUp6CGDjUOSQC7LfOeqAMF4UroEOF
0kACMSJHzaVz5iLveXtf1BTQuxClnRp6C8vgmO7bPuOd2eUWR/2kDAfccGd5lhtI
G6RANQx9E3ByTAr2EarH7KexmuSXwJAJyh35mXs6YT4PXoDhZQM4f7vSwlzdUL1d
RYknwO0P7ERCFSkzXJci8bTbNNV8pSc4TIADCQFUd6rcTEzPX6WDy7Cfd6u45Cus
WUUjv7jhslK03bprGt70ZMOIHpe7qB1Kf6peqEfllQJVIk7rWCM/j2WJv04dwoy6
Z+ziU8opAr55pnxEAv9qvK14ETeaExJD2j4K0LBIR/vqmdxPJHt79ANCGwj8cpqf
T/Ey5fYByiTVoThYOKJFhNoD/PS9Pq1adRfiQKZf+NpAbYb+lgVhwH6o2onutKat
Qq/y1WLXgZwhdNcCKfH3dxiegcEbBTR82Jub8s96kYqU5ZGwiRpTP1kuofBwkvT8
OHn9f2Rs+gP5H6MY4ZEUkjtpDXXo9HAhWCyLY/xESogJf1z8bi+59Z3L9N+ftobu
s44F72QCmYO/+XH/gIvsvY9bjj2zyqETCI2gSh8wAobem5JskOA62pXL3OZW/ccZ
TARESuSOXl5gsKlxY1Vnne56dbLF51mgjXwXfOCDmwHTfQ9V7QISjrZ20x1/yVOD
DgI+pcvSTiIwinczwN4tevZny06JtHwdCwZq1K+adJjYMBCxZHsTl/AFsybFUtuo
UWfgpoUg+bpmcAe9RjLEBJoHULjxu2wy+UscPMGkEqvBagVBu2mW3w0O5SvTMhRd
bU8PxckBDdzd+kzpyCytMvSBaUOYw05Evrdh4KQnvGa6LeKpTOUCm7pup9RJ0d0M
15Qd8/CKTKrclWQ8k6eQGY/Ya/cZjq5Ee/4TL9rZuGrONeelB4qeKj8lyw4yxpEj
Y0bTzTMaLqYLnDRUGu67VQdTjQngg6Xw/3RQdFzU8Q2WtI2RliJzjxz1X1nkZfiq
2nPTanRzE3kSiotXfFB1JjHn0wa7PeMW0UvJZQR0FVN6vsHph1m7kqM3iaZwHFm3
Sl2vsgxhPmYBCg2RuA86nYCIDh0xjmsA0sJ7x6GqI6eXdIbJWIq2Xy7HQU01VojU
INjpc6LV/Owwwh+59raTxunwxPKL9VmEmiIFoGZqZVrejucErW6UKhd5VZY/Bm3r
jEWupDqnazUC8MDF+0IyGMD+LRE4tBpgvOp2Z8glzdJ7WmsKmucPdtBVPbyVy/vx
gVzLenjTt+eRZwYrDre1mh3ij3s6fqpxnsUawhhfdsiEbjR6D+1w9e+k76171aGK
iqK8goPDFGFcju2vm7U5VDzpw8Bc/bcth7jhKB/IJgxNojKfLeMcY+yrRiltCoGo
qtYF+feQTLVH8TQXqbZPFf3gPZZtsi7krxcfJXZ+I2wi/QdUc5jG+ehoR09vBpG5
OzqeENLmU1Lty2ZGc8W0aPxpYpHxYyBOH8/xU41kyOTNLscNij/RxTJgFRf0NNb0
VDhgtpKLHKrpDwL2LHy0PmzfTM+vkXwfEVCLTqF3L4/2j8xeHVqxNuR481bzNgeF
T6ak95eUkRwhLh2UXm1ZQYiRGocFyDffu5oxUt6E58ogq/QJRYBeV1qwCGBpren7
5QZwKAID/zhwFVPOuh9N7XzwaQifxtcDxeCbjNVkWm8SLYieasxXUexl0uo/bzaC
m1LkTq8b+ZXmYRUq1ERrxePIEO995QtPIswqDF54I1t2z+OQyJxJNip9VMQ9+Le4
DN/HKM4PrsHkCdI4TS6fNZqLjHFj9BzfvpLvN2OEo071+4ZGSeNV9p5k4saah86f
PzauhghJRSiHCSCD3QhwVVN+SM4VI/H8qonNLClMDNgc8hclyGx4BMWLe7i7roAg
94R1kzEEVw7Y5/73rSlAuAw/rjUINE3lM2y6Uifj4fXpqtwacWtyYXSDRfbvca/2
+ZZcXTD3ynHouAg0N/F/8JZbmDpVKOCOiKzqebVLhP7TeB0vXjf0LTZto4jFkE96
Vc881R5pXlRA3+sqq10Bnnv5hv+qsJc5s6FzVwmeb4KVfgs26D9aIIp3TUIo4daZ
JbmU6VEDK5w/ffsKD+oYM3oF5msKLuBpLDWYgwuNCoPkOaeHFWfwWaT+PIpcO3yn
LTeqwy8x29bHDvfX7xFkmNSj87n42rxVTopzsqES0R8JdbGrV6MviBXiMrUtCUD0
1zmjMI0iSu4cnPciw4XAxnl2a7pbbbgVpfu59ZgkRTe+M1iIaMZgXsCSt0ojx/z9
JrW+soDIpUoJdLTT1Onjc2z1CT+Z1zxVKqxAh+3sslgxb80edkS21tbNBsfPD2zb
FvO3BToMzfhnozpgHqZZV2U75JENqFATGwfJYya+tcfzdUp3RxfVqDDC+oak96Vj
cATx4QPOFTmKDcrYW2s/ZfVofCDwQlduiCdWEk2hNV4pJgWDidIY/8BSqfzbUUaC
8FyKN/yA5OKDjT46Z+fpgwNdRst8yAbuhRsnBa3rcJqGnrTpJs7I5hIpndB+g8SG
kD8S/7TtgNJqFS4XLnOc629JxEdCTMtgaApEvkyBtvHD5TqUCJZP3mWeGt6iHfLf
0qA9kirjLLh7IuazH9ZtvuTgvsety4Ylz64EOyHPvtZ14/OSxBiyoKpZwu20JOSm
F/ASmVO4VivqHEekjMsvxOE/4ZlCVwbmxAZIJz0KJU27AX2WqAAurVX5opCZzQMZ
pSEioQyvsjCY18JGbVqMklZcqCc8AfYbj0e9XFD0oSylR26p03+m7rPAcJ9A0L27
t70gkIGf6FoGBU+D1e/Vor/RD9heKpS4jp8pgDW3g13XBmCNlJJsHaZ3bdJjYL5r
7z9Kg3oXcb/6TiKJrNohTz/Gn7W1hSF+y1BNxqMoCTSRnzF09rTgkIGcN3tw6Sx2
/grRwXBDSMsTYqk6YFD3X6nKj0O23jbAc6oGfaYMWYt/6oOI3Bm077v1atPueGXo
+jWBzTL7LGhYQSF9sWrahBMQE5CqdkQAhzJzCEdRY2Nuo6RHoTn8F0Qhk4nRIj8E
A3pjidS3/AhnKOJVobYaMA2Dpa5vkwtlqa6BJ8WOlZmQxXhlrRWUxuY4uKC6FSvN
kghxpX3o0nyX3anHwcJoJH0tKkpFGLpPk7xuse+mG9T7kUyKBWintw9LeAyDxkot
ddKbAjZJ/krKcO5eoVQ8WfAoFEuWXkf8OM0+kUZSdh5n6uLSJYo+yHaPzj5aDSKF
L4w/yn3u7pb7JIMuQ8fal+OQBdY2dy6UdpG0Pzd9sM4wrhPfzS17lsV4Iw7OztwK
8MU2zYrQTytg6FiffmnzXvDVFKXZ+EQNS2jsOH4/88X2zHvU2pum9btITodbjKF4
gUDvHfODD9ClEvKLZAnpsvGy1hNHFaQjP3u+d4ws/m0TmtpRDc13hheFp17Mo7SF
7FpvSbw+LVXi1HCuEYUZyuGVvqsGkFCSDRMcT5x3sfWffUpWx1ei1VCT0WuiKRvF
S3HyduLDIFkjWQ1AfGVDN3vVdx/0TNgqYbJmuiZZAk4appnsnI7FAsJtWnWxFyui
NtIJluspyfKfGtJGeNn0m4gCcVTBCiUDmk+8tNI/GMy3LKvxOaeH+RYgx+bN2zva
Tam3Au52nPBlaUbMVGiivhnG/14HwL2SEgG4qWK4YBgk7havvQsuDiuS1U7nEWIy
ej/KDTF7JxvAuuXRTUWW48Y6sBS8W0pg9rOzmHg220eYo+aMw8ytxVuHsDfseMcu
qCtURdIaRVMynp9fVKrnlz6ieyz3FlZKUz4ngyaJk5HM4ykHJy6Kj3BtWAPHn5Xk
JQR5a6MfaR9oSwvBUNQNlsbhjOnN1ulfpSYL74VAOpvXC98j+w10PmQA33z4ONm4
J/7MlzMODOCQmKD8PEeappR5ppOVfuf+IAb/kYqeOKGfVNyWQeRklOiM++UWVM3K
KvRzQKIrqN6hPxABuswdlzEVI5zqiyCIp3Yk/h5pjhKTOX7IdPB+spiZNCVlCvGd
eJeu1t0hFoKK/+CuNcF1IA5xvxIusjKz9mtChOl3PtuoWuGvA5BNFQebXSBUP496
wEnJBa6WputREDq+8Cve/xoBREyTU6PpwtsBrlP7kkG5P+zeRSVs+82TgZAMcAVI
5yMXShqqN22IBpORanbCjz5WMn5hLrnP4/sODLN/OYjOAWNu6NKX2ebmR+2RB88Z
5HjRnfdnk0m3hRwPo5qDviirxCa31hqPsewA+l788z3Rq8YtRmt/JYjMcgoZKj9d
JguEN9K6bq1E00tr05NZ8gGNJM0cFBDtGFAA0dfSQ4daqlFASDYxBxOARAAxNw3a
Ty0q4cleZA4NS5WaRWXlzCxZfwLoGhG1ZgXOyTlq138FQz5N8w9ppgL3nIW0yE/6
mR8ix2eaaYJDT4lRxja/bE00VZpaYsd/sTLbMNmWWa5ys6ToEprW9I3tIdZEFu3V
O9w6ukXIm0pyLqWlXGXKPza2kqutppNDe1WoPQ3PQ5jbbDvAmjnOmc/MZwZL8Kxq
/UWshdT4Ti/twUIMJj41157/amdrQOb41KWu6P3pgy+EwR6HlScSq44m58ssPq0M
x9TzaMEO/dLNX4w2VWRtjMGPrEJhFX0RTV1wZfhAK83XPA5eve9leOJkqhbXeK3L
J2Qf6e/frHwoTbnviPMo9DXglAJZPxqTHyqH9Yu1iQR0zgKRUoK+dapCQuakK0BN
pKBQX07A+YCF3jHN1ZjWL36Cbi7rTY6mlhA2LbHHKwp4Cxh/KMv4I+0/tU5n5W7x
1TqqZutQeL0pqeNeHz/E/V/js7nZ91irXPdBUYQnIyo4O6lWeEIPjv4zPtrutMtD
xfdRwn4UJBf5bXcM0PIXxtH+jcWdswoOPmT1RrqqpibSyVW8qVS1EjI1HrxV/H1A
tQ9KlZtH4WePyF2wy2eid0qGWIIPkS7LOdaexfjUMN7puW97OsuEu0THWNGGMRuC
z0spn4OHdczUq79eI84ObmwvSM35W5oxq/owPc4TjcmgvSZZjVINOXEvyffXtX17
r/1GMuHDyhx8g+ZhZ3f2UxnKUbRrUgd2hNi3Lps8D7KSMbT7jQtGX1EOLP/weKp0
+XyI7lBk4Ing+l4kqocy6ZvmQURFA5Zsr76fv0JBwgA84fx8/e0lz3w/hbNPfhpK
sumu2yTROxMAnsgycwHFB/de6Pwc55W4sV6ruh0/KxIuL0aobOnvFO4G5VUhHwfh
qBIit+1N42eMjVMTICiblYuvX05VCwgFhGgTELjtjYsKy3AlvNREvgUW2vIp3qmH
AtCaRNIGCUy2/mWSYPeqiO/TwTdz9ccll7tq0Cwp+gaRwKsolvJg9W4mcP2nSVUc
yhF78s/Ej0mWTqAhu/dcY6I2swG2mWRK27VotJpSlDyk8Tph5XQBrpIodY1MNaxG
rKiS9d+mLf63Rjm2ur62dxDl4+9u6AwRQUEB6h0evf17NAiYB92c+oHmsMueqGNm
UMel+F7TARj1FAYzIJk2rUWbxhiDncsbzmh8st3OKRVcNdBXcU67LX8J9W0QDn6b
LsfHsnWBMVGMpu2q0lb0rKQmmfIkuVPy+HbyqAWm/dpcbfyxb2fh78FX8yRjM/em
Pa1hq75iB0uG+idSvNuIQ7tng1hWoG6YgEvsNXRQXgO/rIrjYYNDZZOi5m8byhxR
vVHblatT/zz1V9F6YUvJrJu9HNexs47uGdg+7SbQtlxUQkyr8y/0hEczcIhZUIzO
Tf9DuLsZMRNblXr6oQdWk/XUPWD8qeL5mJ0vRkcuFVpoOS2/4Yr1IWIOpDgtcuZA
tiS2eIzX+UGHDYGflU4Gj8IttRLFojdMPfqqlvNSEaki+Qx9tLISV6iBta28Qr7I
nUfD7Esh3aoE+TXMR+CttNJ2MtIIOYcfT+3vaHcMigU4aqsa2DHJQd62W0c/BucT
dc4eZmXg2vydm2kS+Utr8anUhj5UWDmds9ncs/ttScBH9+73h4AEdQJ5vOIe93ee
FuwGR4JAc8vIiJsTBm6cSp46idrkqaIFleucpmNrLHhkCpJj2A+vuxlwb4pGpLyy
yNfRjb3k9XCbEqdN83XUQ6aRtJyKiJg2DZSCyKDlCXp9QJ8PbWJ1cNCHO4qI1psh
tAwxTkyJtnzEsoJ0OIBRJgsAJyJiz26x1spV30m5ECpyglRMvhSI7rfouAMekElU
9DJod9tR98S58lGERFzV8VJjEf9oIpShiz/X8Q6J4blhx37+A2UzGSRqzPZyjBKn
2zsaDBEn97nK0fJL9rPREu4OwNAiq5ds+0Xs2tVRR7i/ST0TnbgjqJzWSS3O+hyZ
6wTR3AG/L/gp+cNy5MbmR9V5bhZ1rLmMoTeScU3rxVblYEDB9VC+6pqhtUJrOxAq
dbKsbbuO3fzLLD3xf57sX+pC4dnN9lLMMYnQ47azkBUHGmKWaUOleneLavVq4QuL
KlnzZQA+bWZMzJQnhZ0LCaV19lKbhT1RPh2rhqLSnqntXNGZEEQG0aLTKFxpd3VQ
tIbKLjiDvRoRK8RrzhF2pP8W+EoOvqGJIa6S4vHED8JTIoVZ272m9sVZwcxs485h
F6gbRWW89SFObbyS1tmPWEwGa2A+shCA/QKRSdKSlrOumuK7tu2TVLDZLlZnYm5K
Q7Xn8r4ySBWAefLwbCqIuWJW5wmoC39f5xYGji3Pyu3iRKkAbqg+Z4MNJ19JU0gN
zBVVMdIqrIiTONkSJrH2K/7pCphX/Go9vvd4elIorstKlpX//JZuG714SdhPYZ1e
tZS6hr2OAw7Vt1OR6bPam5sNu8yvikSBmZ1BHsqoV8+DG0nYw83vgXsUo5kRxnrd
tjtlzC1g7NhtsAhMhOLWyhmCrAXyobfIF7kJIXVhyVCRS0VDaFNxk+3v2X0515R6
3mb27oKb/b6pBqPVv+choe95Ep2F35Wf5AOI2GbfQQSyTWIyZKwE1i0wrJ9OZZKV
JlnH7AHA1ggQ8N38lwjiL265iMtUIqhGTSllaqYQUKA3481FE0+jOOzkBrBDtYTl
fMUsBn31n10724J2FaZ8coaShB4vQg/Hj5CaI19dDJYRNUGu3ioqBmZa5qdLfIU9
h9fCbLlZZxMuaS5hC9f7uMZ6YU6Gt2E3TyNVzRyWfDFIvVL9ggyzzYRGTCNLHcgF
H1OoPGgFGqNIdBE3NvxxRtM4JX10JfIz07/aUQadpfVA51RTJ19Fofzb7BE9ipeU
bshuDjPNeT7AEjOqBNWpWiYoNIt9Kj0cmbE/NT1k/VIoc4reLVd1NRcjj402yWp+
46wI+EMm0ZpC/K64sBKhBtripJtS7hXxZKiuL8rkdDjT6Ieu9Jc4KVFVV4YRP1zt
3deUmEAp+LcVi3r3afPxd9T1lBPeI/EiYVi9Wg2fxYiSVFrJe33d6P3j2sy+u1Cw
YLdqM/j1wg8/9oTNRmOrY9+QOJIau9cQPd4p/5XwwZN6W6YlI3GFxNnwWvNBhgmC
DFgp9jBTucqQJXj0NgfgqmE2whDEIJ4JnXf03fPQM3qTDapptin50CPpMC8gWtLX
T/qlKYqV30kkilnDOX5MxX20SNZvBm5b3Grzr+UHKtT/bklH/2Jo3RaK+p6TMo/M
ZIKBjK8A5u1KtsBKPUsm/7/+drPdbwKoJPieMGab4zekP+N5ARSyPwQSp6y91FJU
AaiklTXT/eM1PkE2yXjxG8hmYw+bPlf+FflnoB4O7muf+6Xk1NzHAPLzTU9swKrb
uJZi4SCeYRjWkUdWM/xE9vk+iYmTOR/bLLLiLOZFhDbO5UYlOxXbPoYDwCo83u15
hy75gCmGIc4+GTBA2LvyBDnIaVGwVr+exAPaCbrMxIiR87rbyDuzTwEcAnIU0FkF
Y0XW5XbPsitExC6lpnZVW3vLuYA1gotkfU+IldlagNGl/H8cpphHZKOHjJZF7eKW
DujtbsI/FDR+bu3kEMRcd1vUPJG4GRTlumPeQRVeU/MgH6qRc1OrfxPb0NF45nyb
cwRevwJW151nxJNJ0CtLggouy9tMFnAHj4WXQk/fcwf9eV/sSqh4lKqUv6Ne4mop
vhE/GDDAZLn1SpC49sxhpc1J4qyBU0IkYQ8Md34g0Yl6N6iXdYN3YDo0ymZJaUwk
RCj4KExm/Z6wYdl4Pmjc37CNcC7FpBw25mbcEOHeEdJdNnLZ3FhSSCH/x+XgGxEi
o4E/rKNeMZc+f1AsCVIwJTJ5rBBOIq1A7BkI31v/gavvEKQ0pRxpkzkhMeAnRTQM
N1Duqfk93moQDsPPlYs/atAcZ11DH53PUO8uZabtiK3+SovLYCpfgpgjFWHNtxNH
CrIXSufu9g9sFwfdltZKU+wjb8K19FS2dhSXm2BHB7pq3krk9/PQWj74lAJPL9hY
DjiQaobILp+JBdW1UdZSlHF/hJnXh7pFCRh9FVZLtezjEymy1zUKWKc3/ZLojQ97
jLYTbry/HY2gmd59HBh34NPeYDqtxT8KKVpHUyaWieTGSYxgTKWTK/HW57DIh790
9tn+ml/Bcccrwx3dFYFlAgBiEualWSq0+tmrIw7qF9ifOa5r1LoqSTjGHiME3zBM
G0qZ2+k/UQP4t75WXtwzC/DQ53TUa2Ds0vuLAqnT4sol8yBzbkUKgqnB8jzmERfa
1YOmL955NL7f0FTf4oUAJWitob+8ZEdoq+lTdIrAEdMz/1Nv/fFSmaOEYsZan5JV
ZfM0TcGebyyvhFC4ze+GXT2Na/ZdNRCZcPqg7pa9HtvWeYwNQKCO3APqnzB++RYa
G07XUU3RUzyysrGGinsv2aCo8NzY7tnugXLd0dJvaTCZi9IM3057lswXYfqiM4kl
Ai2kxFgiNNMrRHg9FnRfVvbbi+YyJ7pjCkDpO8vBqwCJ31NQkeWjTLb/WAQOnH3X
++auQnbuGWJ/YChDDwQ3r1M0dOvkE5htn3K5i8TCLAXRfJZqmFVRmowfz+Lox3wa
8TcxgE8GA2/50m6JtGx90AIEYjA0CFV41KeNk5rwrfVMmX5VnpI6mNs0cBb9ktvI
/7oZVtf7sHK+7s/nv9Hdg9AQwnwnsafp+kcICP7PZnwZVPJ+Dey5PV3P/n63MM5X
vxcrJxtoswXSSgYpgmps6LGz6wrjCURUei+E3NP96DzE9Bl2GyKVGrkohNiQaKvO
vp3L4XI45B+uAKCflIpjFT/yH3GRqtqgE6KHM3Evc8t7aca4fHzPIjVU7BnRqc4x
sdq6ZNKdj9DBltDFz1ofa+4aXTsIn4ETOPH+IkHCd/g9BOTsSeyuHig+JfkSwz38
+Awlc7mm/n8O/ZgeV+Y6+HKc0U98HkJsYbWNhOYykyBLo6bfEA3N31GmRZsQbvxM
uSh6pegvN+dKRxsQZ7/sbJzPcHmFiTXhnY7OF1CVW8Nyfb9Z4avfUU31aYGziJrw
WUT5WJGHJjMGt9wr1J3u80SQPLughBXUB6rOtGNO78yJiEjs9iag61p7wRJsJ2rh
cj7zQdALW7uu0iykRF4XcDJHZkN1/RDnRka380MnyVb6H+2FX6+Zw2xLbVVlpMFU
d4zsW6GuzYIOiYgtlRXBpuQr0+f6tVy47Ov4pjyAZw3DQngdyoGtjr6Pj91YQW38
NUF30KeOjqXY9mH5uo/M5wzhUQeeF726I59g3s2CCm2jZWXqBH24+5S9oyPxC1hN
OimMtU2bLbYP/bXdj2QfKSix7KbwESVIKVZFu8BdjphKfldvwqNps6+Ng6/eQxlN
YpnO6mRTLnuUnHwoUkiMkeHj/iDWuM2zQwckGqY+nrm/8dl4L6PdbCkEFmwwZKuk
GOsSXGRxygzjI07ZsrAFN1CNDQ+O3On4e9gH/nCP3iG4roGeE1f0jYCN5lRSBnnO
/DKSCQ5QCslzKbbMbCf6LiOv2rkLSCuBdoyeFkwSZH6ZefImBShXnGG/osqvvEIs
a4L4e58Q+IHn5vxlsH0UlRyOUh5I1pYTcZUfMvd3ybzXRDEPmADnLqDvwIgdar/F
CTDsSN+FgT7HJAxHdDja3aclEO5QiOrQYYq0HdS644J2KI1zURg+7p5+/X0qf5FT
OB7y1IZCIlFYR7ZhtKwVOlFMspXiZ4RYyg95yGrgA32pjhN7gHbyhq3ZcrEL9Wtg
TY09SqKKFjkZALXJ3imw8lh+2Pvl2RzmZPWxg46cWbG6LH0pnRwh7wRqEdXTePsI
zDI6E3OtvGSQPLJxdW4Quc/SmXhGRqeVzB0IXplRwv2uMFq1LyQEAZNsRdbH3CpL
rwQtdofVAq3v0nEdBHr5+p5TlSODDLCJYONoHDEv3lcCKdmYxqYhnoFpUsGJUppb
D1iXVM3AayRmOOvD9W3PvCjQt6AO+jJh6Z9J4kURcklbFwhK+buOKqcsItfAxoY1
Sv1Bymrn4Yqp3JUbzGLc31h4udpBf5djrwCJyJbUaUWVs3hld47ZtNl+9PgNF8m3
blWI3/eCHWCa4y7jpVv16xfqakUY9omd0HETjNTiGmtCMP+e5Xcg0LcvsnV3B4q9
p+5Y4gFB7n6t5vzimwx0Dsbty1+c5XnyYsGtlwrBwMJ2idspqWuMzmPDZu6TBVfq
0aTTEUQdFQ01+PtFS+pMui11hgBi3ji/dF8RDHeju0fzVLuHP/VhCtOZ+GlqAw/P
XnrA22SUoyIXxl8kUfQrdO0V+tQU0lca9ElX0OapCqNeDR0hsRPBROR4e9TrTZ79
H5Wbw6vcuOu/ABAMGh2K4rUt962Mi0C7vS7Fd0rsyMMn36JOgYQDwmFI5MgtN/34
D5DZHLv1s4JAWvoo65gQ1AUvOOc0JnvUFAPLpGu9/fwaaFPE8AuN9dqzwyijV2/M
trSLneHQAtJTSewlaeXqlieuB6Iw9+AfD6XpC602RD4HsrlTQlZabeLxpq56g8Pt
tkUcWBCz9Gt+UmOzKltgU3CB2M3AMd4QES+PfidlCVOFavAgOOd1omshwhG+CewT
fsoZqJaRjtb3nwcAGCGkNigzOWdt5wY8HtI7SDMctTy5kQmWKve+tP3UeeZhlGfT
qlq2P+TGVto9adJYCIyjjn+LBKxwnZfIXBkFJdoVyr1umViIRf25I5xG7S9HQzgu
Qg7iyfLzpNw3UlCxHQQSY7USAHSyJ3aX9lkwq9274nz7XeJEEYoa2+MrWwPjT3ig
UQDxrxkjqH3puaS+ozqoAZYQeu4pVaF9ejBQHdaWrNiNvSkam8Ayi5nWsTc+l7a1
1jIrZJjUEu2/HZTwPCGlarEFAeZnvrl+f3ccgk1JlhnqITd6UjKoyfH17oSschUg
7RK7zt/t8sw9NKf6fhmoCoG/OuXgN6Ri2nknNA14Irb4wAblF5/yK0Q10f3lhvre
tdyyZRKSVHSaoOh/pysqo8XhpJtZx76z+exZghHXqYjjAzaGJWOwx+m2yMVmPJCU
njXmHELJkqn2k0hYt9koLnp/2iTqw90QmSCexNzrncIsPGRIAfzp1Ty09n++DrGW
IMtFbRRaZAXV+b9SzzG1z2orNc2r+ORsVs4d46d9+fk1T6aZRH0iYySBl+AjEF6s
gm2h5TegRqaG/VpwjVvq7OrU6/ENxxQt87y4h/DcveY00vvFO3fVxWqFJ7Id7k2o
ednCg2EkrkcwdHwziZumHcddtIJziPWaHkBnO+aRbZteRcYScnmWNqGJNob+SO2S
SESfMhFcUhDof6qw4xtMvjNr2R1gEICvirlxpw3LT3TzZhdvrqE98lb9/42ylsIa
UkCbyrX3NNGDGnmKIx7nSNcYVfBdMV9r8niJldaGDA7GuaHYhE2ALLfEde6l1ULA
9IiA9duNPJ0lYVv+Eh+H363rDdWAAIV/R3LMn8cBmZrXvXJ8u7l83cn+5NRKO0H3
sr0nv7JZSiFCcStT2vj6l02lodrDhzr4XRLsXT1TOQJgoN0CUkBUXIWSrzrnCKcv
kVDItbPoWMuzxgiJbq81+MVff/12LpPg3Us0IATHfIqeOFrGjcCvMzLoBLPhIpzM
peDWM5ZSA3vITvvbGRKpzBmaYmIrM25zKQzYGRFMy+N7uic69lJb/3YszswfvxcP
87yyplM/IRw8XOmYQJKjoSdHsbh0iJpmZIPk32tndequzL2rJMSSN5CQQGeaz4nh
73onT05G//6XrNoKa0wSEvcFQ45M6EQbR/XaCd8yNzsc3PjL7k4mH/e8pj2IgWN+
8saoPHdSD38ETAWpM+cfUuFsNv2ydfokpeAgN4waUZf0jAojqVeZP+WilLCd36mt
vOltXLallM2ct8iCAlLlhTgLSmjfS5w5g8ZF1yJT3SknS+Q6pJIK06d+67YcraWF
p0ZTUQ+6K1B1pMDC1e8/QMPrggx/uMhQQywqgK6UNvGlmDkjVV7uHArviBVTEGA+
EBblPnZ7nbqGH+g4zszWLFdhEGJXQwuCyYd3bOY1Tn2g1N4GYltaGosiS5o1kRZH
4LZv5aFoGwe43VvxN5tnl0f5zT34h2G06MyXV0cEuaJyw0hmnPffHILFMPKl9otA
C47kRoHE1fd5yAbDIGU3JFrQ62SGBWsM5MS7MUxLJ9VAuPR/fd5NxovCgW4UiYsh
HyjGfi3Q/bRR2eWxMjyp2l48plOwIQTs7yKkqnHZsHPfjI7ZFN1LvcvcFPMYmyCw
/m7+5qL32Q/Fm53bRq8q0BlRlFxG6WcBGrWeO4w2sd8BXIEB1pfILIGDiEcFuNlZ
z45VZrV2q9h9inicR9o691UiJliIGcpi8LxSBJFAUsPc7qtcE2q2D4Chaap4NMDx
R1w4fx3IjCx36vmo3PP2Dyd3SUPNVwqSW2WrL2lbpjBgCzlTZmzOZ8Q6Rzx7KfSq
Y9vOeOK7K84Kt7nULqnpXw0oo7Pnga09IepXgpKv+67UhfBjD7OKJF8HW1wbOBlN
fXv3IvVbPe9cuUMSe2uYXBxQjzR13arc5KOPlhYnXl9p0C96cTxtKrgaTtar8WKS
NtyOoN4OZ6eAp0huGCzo47bqftyOnaTop0SRCHzRWMPN3O963DdIww96sug6FULB
oe8yLn2KUM/s5CR00r5qjnar65rmQkQ04ARPhvygqaKTjd6f4fGX3RPDK4eBbuUw
ZOV4VdbY+JOFkR9dETlKDq/DdAznM+3uxRLCJHzIKXHJZIwNoQbEpUujWBgQwwrn
co4yyEvC+tsj8DRW5Y9uEuuAAXaHStDi5gruR/HHYVXlenTbw7xRcUWbmVYACpMk
r2Snxoi83OubMVS4qRSbOlXFMw5b6DNuy0tyD2zMxtaGFD4Eh0gLcaYzFmczQHOu
+tqmPXqa+4bPHMHb+dWjxxEK/IuWj9oDkU38FJX7W4i1RUmN0R7EWjIlcP7KdDov
T0YDxMYrINpgUVwtmKQdvoEnyGav3OWbeNxb4VOzb1sFUZiihGpP8J1oEgKn2//D
L7rOcGtpq4FDxp2ZB5GV1jSWLguvmmMAIqWWP0xZYjLaChNH0Pv8Cvn5m8dgK6Mi
0nlXDXgtKHew0ez1ReNyYPgBCLPOOHMTHitv1aiXfVHtBk9R/ycpjq1Hc4XI0wZ5
h+6/tGQ9ok/X0ASDAcvYLXUHMkPZ9VSO/NHGPvntbw5+9qSfTPtuyipkoQjNeP2k
/u/lY/8ggMRzgkMc06XgqGSU4hXw47dx48PlKoXieTPUCqp7DMpyBJ+so1JCvKlu
JQqiLeuNoSIlpEsN0LKnRBw2/18dVcbmztXRoEDNGT4NKgbmJUfBhJIOWGl9YjYo
oqZVZIiMvwLzeju08SIelBfmZGd7gEK3+O97ke1neKPVR87TYNr64sAH+YjtLZJY
MUloCc+HzxGRvhAHYa8HdI6HvuQGdWe3xjDeLzcVW+wC48wLYyotlg+yDxglW8my
NEKVJx2BUDA+JX8n/YWB/U0CVwQEYD2dFJJmfPdu3pFzC7t5oNZKwnG+GmMcZxYn
b6UpTyafQCWmsUtm3kJeaWlAoimjyNrXXACm8TvQ/rNr5zfnAmGC2geSSVrXYT7b
0DG9SVFfLokJhNlbh0q3VSrTKkh6cLdmVPsEndZTKjAgcan6amCEDaF27Aut3HEZ
fnFSxtDX3NgmBOjB6EzOgOFZJdVcEsM9D4Z/25GW6hnqt0CIoixvyrR4ROhNMP7y
nuoUbfm45LY8CC1L0mArjl0Vx96/IBIISO6kAK49gNtw+mDENRoHaoqIpajEaofO
ooDuywsiN/H8ooaYovtrAWnEzy6r5Pyhp2/5ijpz5rUyiF5EM1v/OP+swAJDLRmm
oMgWH5pjRtMYLxeHHeMbBOJhKFe780LRGBc4E5mf7tSXhc2X8BpB/pN6ZRh69gky
ChTpfTusn2a9SxedNSf7GWy/r4rIyYjkLYk+uVJHklhGLoI+7loJvHurPS4AE7BB
mujLJAKcJKAtHUmpgyXzQV1lyRl83dUfXKlbPQ2m+ZRdVCqV6IZu/AHXGVaFrO+4
THn+8hAXVD2VTwmUnRuf9EM4iJCukFbW6zOpKndBUudj4mWcdbUDtNWpMUqogn4L
CRAOXhl8oxspEib/bAjoIzl1xY5o1P4qAtdu6/GWEh4wUrGkPEI1jJ7YFM0F+PR6
Zk8MnHubxRamLROJs/kjCo1nydcX2/OMe7xD0XZwZ2PuF3krFlnPEbFu0xsqfHbt
aZocZNSexMM7t4z+7I/rECyP4zaZyGIt5nfBprhjyQpdA24QsHe7/EPihVJBsB4y
380OauWHGhnVB0RhhRRc1SOS+6l1OzKNqU6NMYjRfH3oAbNRaBtL8bFzn8M9DAMT
YgphU1NBWUjc3RYw+ABAv8/kLKrW8av08Y/Foo0RQ7CHWQNnVzhCcTDuzPovTf5V
R3CYDMx9HpMs4dW9fMoiZGVFJe4kirUWSY8zr9hLFiFCR+6rpdK3u4GXN1sxjd86
yyNAA5a5nOFWW9c3rDM64ViXc/AR2iYyKMfnwOTDJt70Q9MFGLtTNDxgjkZFoda0
W8/w7xjtAuLH4a4XVCJl2tv6rM4m7jzF7MXFvs+Xv/6qSC2SGdWyfZ496XszeXLg
quLS1mXgwXT73bUyf/oPzZfcZf9LaLWVPVe/zGDeI4EeKDIkPATnliycbVXYIuW8
GPfYWmgsd4UmJ7qq0WxzI6r1tv2+l3ps6TJLwMaaijLT6n01hh0bA9PgCsZK3qSv
2bjN3s3AESoF+kV12Y+hl/nD+Ge4+/YwIDCmYw0ylk/d1Htp0YtG2r6hcS/7ZXCo
tCxp6Kkkd7z+5xmjZt0ofyvDh1iAXuOekNDR2/N306NsO0xDfkr3OUYyLckwr2y3
dxIPJGvi5rMCw/d5/3DmOCfGQCKv2IicDjYoPBSviE2TxyZh7KRn9jCG6PFSOLAJ
brNU/+qaTPSU8gJjKqb+no3DxcPtbaO0O+u41m/vxtOtwYhAQPEbgI5gFBA7viZa
nygqAKnfrBFxSWgY8eY7WT/ci0mH5W7oJahFEc8XuNpsBJor1Gvz2t02PhFbNfMi
zAvxfsKU/dEYZv2sKNkfs4vIESRKwA4ycYxTrvFHoX+hJFXIdA/LfDhFfl8LHcYR
PZBNLdgMbhXyVBjoEAz0ZeZ9dAdLI4NSlDowVlLLg2JGmN2I5VmoWxoPGBTPaH0i
t/bXcUCvFGeYmSD+YU+FH/4uaY9ncuLS0aqP6H8lLUiiTR1u99h6mZUpypXoMg/K
dS1IY8M+N37ok1Cn2mMdG8J7KUimY5TeXjJrsEIMekvcGB+T+j6ZIgSSNBstIBDZ
UNubDtl6VvlZVdiPcKHZZWHsWuaXw0N962ObLyGI1dkkMNNZDWs/ySy6cQmgPyu2
s44BeGmMURJJtIQvq9Bva7m362nxA8HoxBobp20uD6udSz8KLUY2lfA98gSUvvJF
95VKkUIKpZ1Pt7gS8/uDuFcQkXG2kKsezOUpioktAqCy4wTTCbl95TX+HiFhQ/mM
Iv+Pa9BqQ45l9c48gNxxzRCewN7OjD6Y3fWxsclj47BOmDiMDg47jiyI2w+0tXGg
kFJvVy9q7FJsyPDLY6o5KpyNM3krjB0MSXGRVRmZgJDBLv3qV579E/TCU8OZY2hn
uWNKVWqrkPIXVZZPfRsE1lTZcWFpVrZLi3aHWFv7RpzvudDsnCQJtfKdFmYyImZj
ILXNwoQ2ml2RVHAGnzJuJ46UiiqEIqyN4FEnySwnTrUHt3EpYNbV383Or6GGNV+I
F5qJjaiXJKQbCBk7WjQmnUrhQs7n/5bDYw9LogmoAQFy9wBU4B/hTfFcQ2p2+4uA
kfVfaV5blZO5AQUqHD8rxNT6RJcUH0XR5uoQ3jUhaS99F1wMzJ6yFgFddHqXFPJK
jE2iEaJyPGIjIY8fNUstwMStdJeK67fVRFi4ArBSRACF7d9x4B/loFYOlBCcnAVj
AT1p1wpDwCWbdK0eIV3FA1DDIaVT9GvlxZR8egWng2P5K1XIDhqxT9/EfkjYgC65
eAwYjqvmeLrQrRuiyJhq6R9ICcm03fQO0i1B9EO3LaTU/YdOVxpmCQ4YkyzatDr4
f9o0ybzePp4uimHxLBK/St6vD8VFo1h2RM7H1V4a/7JAf41WQMtrnkrjqdzaskGf
/yjpL3pd5+sM+/d48iJIx8ntzJ92srN8OfzzgBXLVHTuEAxK8fqLSNNmqCdPU6k7
IYpbD8T9Q/U9fGwUEgL0wOf/tCr4/RdhHF+bRgpvhI1LHtEbcQulxbyVK83fin+p
ldxeyHoeLU3sr4YkLOWG7ESKvuNMkpOzSPiI37thZ5moyH7/ncCH30ZCtSqy1dBp
kMYYnPuritjkKxH5Xt6z64XWw4qJYtZXBl/OkQjZ1qAYTQ4h2yrE//n/8L8rC/QY
1atenMd34jhD71z+xsNqZRGianJCN9RvoV3f3zBT3sYq3+mGwSs3S4ci+zQ4Pk4X
IdSqTLHGwbsktw1JnDiSSzd6s5jEP0VbW1iMyx6AH84EEW3WOVxFDQUspy0npriP
Ck2yX8mqllawbfe3iAMfefPnjZSniyamnDjDd6ORdYXM0huwK3lwPK8R8U+tBxfF
R+foRphGwKZeFWVM4vRqxWy+V8diA9sprQcLNDV+qLrzDFpq9DUE8WIcPp1cAotn
nPSLID6L2J3ly+4FfXkMVGBFZEI4KWEq+9k0IG2ESYQZ0mUrlAhjTTbMb+OAOm1n
L9XzX+7cQMhZ8atLDuxPyH1P6h139LvDFU1jZODkHn9Hlr/5HqmmF3WG9Ky2/rpe
FuumOh12LwCpJFMlBcVXJuX7+hrmLRboiugskgrTFKbYEUjhJOvWzp8wRj5zKVTh
j8Q69eBIe427i2GsBpWN0cogKbWp5gC0N4OTWc11TUQ53bp5fW6YGAju+GDE15Xt
y53oOHaP3JM8OAjpzfXmdmbPCN8cg3+uirWJ8H5shP0NM8ZuPSCOBKIUBU9/QvMc
QiggMCF+iB0gafoGlLCbOLEwUFn61IjVEt/jp81ZfY9mZzWEiIUo9ZDbmPbb4vax
eV0ff4IyU8XocZFfiWFEsMqH0zzyWlOlmFymBN6MtJsku9p6SsHxGwCLIE9EG4n5
lCGkq1h0Qhdggr++3EvjdkSBV3Afzyce+uwunYy6mQbXO1KB8E7rONGDX8xT9jkQ
Dq7Cotyw5gLrNBzotWYrl5DhvEPWU3M5HHVkFIYjRa3g2z5+aX0z/DEDIBYE4ifO
1/7KFuNwcqkDoEMDF6gnmAY+yPKpq/h2X6dDQVRJNFwPE+C0Cm47+zRZfad6QMGm
aWtXZ8h+K2Oe795YFLnrHnkOe9xm9KZg4VOY8+STCq1dZD46Q7heWhb3/1KxfyPG
gWRcFy+LvRHlZUDbkHVzyqTO5RJoE5CLojQt8QJZ9LQpvwBblq2uHbMvXDpXfU/T
mYYCAM2uvI268y56yEB3BArXo76rzRmdVhInbUvWF77UXm7JgDHuanT4lHYoMOzG
rGqqFW+vJ0GbMwM/VPTOsYPzcnmg7CoRfhk3vk3+C3TdqKWhj1id5jOVrBRJQRHv
zLN/IDqQgJaWFBtymoXZ1ni+y+ZiaaDbFva6iq1gO1fHeu8FITS2ZDLA4cY/J582
t9G6ajBnYQ5beqEIYgBYzxTgMP5Db8Wz0QYKXnZRh0FyWIqSVt74m5jc5PlYZLTs
KfCEVySBG5jW8wR3GF7Ylp/e5/qQ2j7Fsa5TwDNEduCotSEHWLxFp1xm8oI5mTU5
wYsy7MwlJ6Ug0N4s6/Vt9+54rlAG+suOdmzi9H+wsLMPZ0debrf9TJU4ydiuu3k8
9T320qdEoCIXpFIviKTkkeuFSFzCZ9YU+LcdXyuMO7EcCG1HOZlTz2cpWoDmr9Gz
cxQ3z8ITlli3nqZPNmbFgxuHcCUD+8J6ix7Uj72S50qoDuaZUlS9ZHLBzg4u6zUo
/2ym1FO/+oGC9b4P8ZpLGv3qELNwXoVkCAa5g/jS5X5/8LqgsmdFq951kLkzUCQX
XRwF7xgPlYwjvbRNtdsNSDg6TogxW3SFj/sW19OgPf5rQzNjDq27XXZIgoKKYqEh
2CYWues6jlzI96YMvMGphEDFPS6jnMsOqP0CUZ3Je9LfUvxi8KgQrb/HQlcaRgDN
qfkHxWkSP5pnw7+HMq2lo6Fqzg7EF4nSz0z660lYu/+uU+iX9RUyznNYXfyV5IWa
FUkwg3haX2edEjLoQGYBKML7g7V4XNnb0lw+K3WwMurG7DEpKATXP8zZn98KUsHL
ftmZabar1/B8IFOPJtvauxlNS2NT7yRLZ9hkTaFGq9T058VRqTLsD2xXtFQq/hs7
7cPDJSSpLh3TlOw5GVWlY3QAV8wQo2vHfwsuQ4/BJBfuZDL63Few0PxavPPFH7eE
Jh81KYOmE+D+LtPuf5dfsUL09XsRBlKaQ6v2MOYoVP1EOMCy3RStaS27zlEdlwJ9
fm/hqh5IfgbrIObTLFP96uMb4Izj8KfqRzFtQSycScPOmAgsxdBUSPbjnCIwwLqN
EZqr1E2cfLp1AB2BFb2b8gV6GIBV0UzvgzP138BjZpgLFKFbCIjLnLLtIZUTyzrv
4TPFfMLhvQcn1JLsqrbHZKW+cR7NGvmCM5didsxHnk8BvwGOdtp/HgtmBksqT8Ni
2ze6LrWg3zSIqvcozrKmj2nPJukDsfUUgKBMW7cZc19ZO9L+mnyTH6LMDPq0QtGI
ttWeJJKWUu3ozERzsTXUHTCbKv8dEvE7eWjo+Ukop/FI+2kbQ1OVYnU7sbuXJjYo
MiN6uFkS2KWsjUWJQeaZ2K1WaMoTeivApmwJIsgOGUwqGn4Al27r01BpFg+KKqct
p/DgZGLCj0DWSga7azGfPpPwpkq+zXfPHxQlefW9VxE8ASjXOGE9/AA5tEiNMbev
SDx/NJjC95I1vGYYoR5nnv8swsPscK/X/oC4ZBysXkZdJTl1vJvs5VS2vxiISO8E
rW3+x8aSLlPvEW//njrIAFETYpD24NlZB3kZtoPSgfy1VVo7F7LFCaZbngMRYmfm
98HmMZhEjStBBhbgs4ce/5h33cH6afOpmkLi7nO4Akxn6JgktSqQrru0wETdAxSo
AnYpOYUIZ/cjThyDRU0QS8HhYKpVYIU9dRhUqwhAAs92vXKj9dfm5c+M79XTgby/
iBPMldJRr8s2Nr3f5Yo7riuSnix4TP5gGXv1MhRjTvnyR5VxTbWY/CbtF7a6xpo9
wkWELgB5b75XBrZchXhlnyg6fX/GV+aKqQulDNwibkmtPqsCVRTsh7C378WSONkv
HGnNfPViBfixhK15yF5m8uxg06/exAHPTLjcHPJIVuLOHeXt36+miAGOVuWJWWdB
C/aeWZTX9T4RrVRCEFNXzRXpQitg2ypDQJuKERi9+nEGMOLxypsI/s31E95wfyO3
UFn30lnsVs5qmbm0kOnQdhodgOeItbEzA940Rk1xxj4T6YAxxISv6JgdKMckPNlp
nURH5ev6dDEyK/pyateYi5HBpa0UMOezapwH4rRIkXGuANCc3uB1iMlwCxiHOHUH
QmKDmFdt8ynssEOsA4B2yNTBghdjfZyhmYmZBA5Nf2oa/kSIzdBLu2s5lnwWbXuD
dRDzUa9z7bq5ya1FOxlNy8cw4QGEN2M6PshJYgk407qmklWowFhbYi1wWamLWXRo
BVVE+1qK8DYkbQRWSKmPOGeuxZEAMV8YUU1APZeduWti/fhiRRpmKqWmD3hkV8Lt
5P+VN1UTgguAXehKu/THvud+cVhpyAPqWJVTeyYUZr9w2EsuP8Sqao9qeoftgQR+
xYmnIPWkHCJ/Emzzfu5M2VPF7xQp8sQak/6CWcjBQ4Xg1X2o2sGyjRPxhqAXPChH
/fnxUPYys25uwfzKOKX9keIHPAr65uMRqX950nr/icNqvS4waw970aXBF/aAUaCU
EOz/umhLiE/6Tc41oCoMdDYBHwhy2BWglYdhuprb1cQ9KCHtZo4+vKi7RB+CGiW+
mnl2+LJ55J66dFn7inoslUOJMyWPwx++I1efT6cZu1gp43YLCYWWpkU5e0Pb+Sbw
7XMClIx/68K96pVGkUpsy1LFkkfyMApjFTMjR3wA6X0ONk1+DQqBblOPpdqqty8F
qZaC/11HYDDGWsSAR1lQRfcF6ciwZVLvfVOx393rEhKDHmQWdB/enYL3cwxwxy8+
KYaUJo0ajPAwtz2+jysxUBa+i8T+R3UCJIHlooDZTaq3VgnyUJ8DzDrPGeyOkJ0k
XnPnMpdx8EfA2G8pccJ2L30pC7YAo2h63zbvi8gAZ2GSXVfuC/G3nXQhEagpFkjU
olDW+y+LdhHSnrrPF6ugjgo5Ea2cwHfHqkO2KJHk0/xtO0FT+wU8Sejh70nSTpnO
lIQAZSshYTDxeoA9gVUrfd/1GvzHeS9sHBSt0+NR5oI6dZJIwWLsExa7baklL8vR
DOwb1+/pGBPXbSFQCuCOtF1ROQGLOlSRcNsRj+1zsPfFIAek97anljUMrRw/tOl3
+/SlZnBPwwUvSKbaYo/KpTA34LDM0EzYkPIVqCB/XUgxhp80h+SgxyuIvqCqdzdR
i/zJUj7DK6hYKvss5IfbH02696zZfJJL8zqZl2Ud5plD4iPZKetQcFY0HHbYXIWz
Bg6J4e06h/u3eAPUolWMjI/DuAzz3Wk3Q25SFR7H5gZMtOAQKOG7q0HEBIw2Y/Fa
4Gkql9h5kFKPgp1D7ELPKOjMrKgVFKtgl+q8ponIOuDZrIxBxBWQkkh+Z9m2qvHi
uUuECp+mjVlTIa0dZK8156TzdVLaw72CadNtU3+0hyENGvkfmVm+MTwsr6DG+XIa
bilSbzVg7CQlaoRbq4e41ZAVaZwrpjdAli2sQ9uczaFgeRfn2+BDXelEm0wrSdLs
BMqOFYRSmHlikhSwNfcrjTkCH45fypuFqh+YGAJnXf87/QwUyoDNbdqamV0jlIso
fxqpsVbwDnAg9iYKWRAfO7ziBreNw8/OUn+9pzETxR99WEQzjFlx+Tx7g2Ose/JW
eIGPCMfi3rBi67N/4n4EoAWJEqFT8oU7AhJdC+7tN+Tx8ni6VcMzhA2/O37aJmrb
oF/EOE+0Bskk0T19S2UuF14Y/LtOlLsayMsWD7FOQ9Xgq73vjOc5C3CWe8PQ2hY/
1WhANIfHKG7LoSDyLUsDx0KhdfY2U4QWqsHTXAl8qtBvBWWWxfBUe5FKQIOstp+5
FbdxwsmK8nKH9cCDYWpjT8nC4GFio9WeV8MhQTkJJA+jPvo8nNcui1Rat7osANX6
P7NRyCfPj8xPaAmuzjtCe4lj9N17PFTjIpEXaifKUrQDxxp0OpYYUeEmaXOdY0O2
P+qQRLd5zuWPJz+zBavWZ/4AHMIL0cy4DWj43K1xg/Q9cSjrfImc/ehylKhRpkqU
aJ0cYZHULiEB+GLURhXwRfM3+gnjR2E7Ye0w1tHjunK6oe9k5WZEUHz28XVuEL80
NSJeekrwOtrJB70+vWt5HvLoI1fhynvMeGer+IO+vh+MEq6zyOS137HoHIKzT0f6
BnY5qnaOHsIOkPsyubOWZDen/KYilW2r7p36+PaIJSEGj/2CBbgyqsRlBttmHUVe
4syaRN0TxPfLcFRI3ZLk4nX9H5YbkTc3Zz7ibUsfXjw2HvjplJZ43DZXwWaxUAbq
I7L/DlaCWWUWwvQQn8I4wCpR9VSg1ICh/55OzgOtWtehSdecNW1Udh6vA5WI8a6u
L/8o6pa8vgXfb104BLS+P5DPNWZmzP8d59m+y2Z9tkecTg502Su4q9shOYgh7ViF
21aDtoxbpPfSFZd7hwwYWJroHGs/o8ikdJXH+0Ubiepdlmku2SOkiBeMVDsHXoud
Uxo0vtY9xPV1MWubO1/en7rZdIiNnzl4YesYAeLwanIbksRDlx48FViCDaqZXI2T
mibzO60ON/YThaH20oyfLj+euGr4dBp/NTr/8x0wACSXWdnWwr56Cg+K3s4C6gt2
R61noEdNtpN25SaPMOi+Ah9Du0NvvGcNQEWqd17Shs5bsql/JF0vj8z/fh0pWPub
7QaePgmS5RqA85D7lhwvqSfljWCpxUghzWxHpS4T0LdiFe+P49vUopm+TsyHIoBg
hmysTX6ZH4u5SfQ6qbTv7It2IFxa8jRxPZsbSkdr9jx3PRCNmQZ9whNj/0KxgNZi
B0z56TDO+xWVxq9tPGK0GeGDQQ8olkv66tRy49lLlpoKLXcPynjwlrIxHLWcl+El
Yfy/DMEVVVYHesDwTJ1/Kk4qCK2E8AWz4maMzfN/f2f2KP15Hh//ZjlCe0NhuAGs
hnj7O2+Sx77Nxapi8nGaTwA41MfeCMfdy1PiWzton7pnumNYDcBseBNLPXFGiEw4
ADHPS98+rW+QfzwwcQjjRZoedOp8r3BisQrju+mM+YhxL9qeaVqxLgdzkAHaF0Fx
KIBKg3uJ7EZ2yfcCW82pP55BpVQQ+bdxDcXcp5LY4YgNd9jHvFupeYsnOA5kViCB
r1nmyse5v7RCQVaE+HfU6KoitsJEqOjIwPqIY0UWNEoU/qNzOWTt55vREDSlluEN
hRGWWzyuvh6Wu14eFyYF3jCWB99YJZkUy7jiupByUbPE+U6hdBhXqb8Ok7WVhQy5
sU3sAUFZiIlrLJw6uwnKSXR3Bxi2n99EdXYJauwmk3oIE9qAkcgXFS09aWcRcZFz
mwHOKqtwp5DfxKepI7CGCUQWwF+o1tIoawwTuABVCXYh/svtCKZ4UBBNIy6zhjqK
pKETVGBY+V7nLES4OmXx6cD8BTUVGsGqiyKE8yaxx2b6PhWpJdHzWJyFInL0Gkgm
6lLwp+r8HOeQnPpwx/rf1A/E2ipTaN14xNIS55ebS5irhZi4FkveNNaG7gObPsBA
Tu+ahxysvtDEXLK1IZ99kIFn4amrQWIUGbCrACBMeJ6lwIxeAMStD6vRrR3ZC4R7
dYMq2R/i90a7E9bjps4o6lltE+52TQcm4i57PWpBClEVHtcJv4oNfwFgJabzrkf0
wlsy7FM4CGS/8u5Gz+BzyU5msJ/sdHQ7A2XsLfMS+kc/PA8gNs6kI1mO2knO2zCW
ueSkLK23xNWqWwiwK6OwjnATrXBFyom/NRjzeED80PHTeCIYyXNaRFaKhqqU5M4r
gFXj2BfQWlL6six5aEBXZOcsnUfGyPWgIlVxT76oLNs3o44tiAYFTvEz1kEH1tAr
dU/kHpiDZ618bAf7ZNIpVpwtqI+8c2GlsX5wc6brHD3O/HhOluC5AdCp0RLh6ZjC
3UBiuvTeOZkJXqaWvHV4vCqiG5GY5JSV6lE43SxTQO67eTUg7FsYyRakjw0VM4cq
JAj1nxuMQnCT/snTran0R7pGVWwlBGl8R5CqpvmhRIBp+f8kbTUW4CP/VILaMWQE
Ppy4dZVsdwPi7EH9uHH6ANDQ1Ze+zeCqG2sWN+XTKSxIvaKV/9Jsot4ciEler9/A
gcYWh4tD9vtTApIiumWtxbdCFvoQdppTt7xC2V0uo4+wWn5kozRoVEbp5e8yuLwB
Il7chnYiJA1hnRC2tdvgG1zwEzQDV/dxnAQpY2CSBHZIGfSZLasTYC7kIlTs6aJm
kzn+JsxFrHXkpKWu+3L/SaCjUJszG/7XoCs82bwdSs+pCkk08Sv7SaB6Qb2or8ME
VSs49TjjaEnnCowmkjnLtAlEKGG5DThHoJ4Us/yxzR6hjCtqo1AEb8lr8SIytbW1
HVw/9YgZoeCBfzMY8Ie1qtnyb7IuW2hZunX99tiLAZAeobGeIgCNgzu4ZBar72VH
QDaY9MVjacyy/gss3FK0XaznwX+5XyPts4ZhX4lefEriDQxXZPaPwtk5DqGIt5vN
DPzfddHK0vZhFriNLqEpTKv2JkvOxTVaaR2o0HAoDmX/W1KMgd1J6q/8D/blS2uV
5gIKQxv6oUDiJX9HJkO21VZhx35VKomjcxnPIbWkOrMTmymO68oMaf4JnuFVmPB4
3uK0xeyoEb0+WRFnMnUJySt1t/Bczjbn5WWOZq9u2cTzQ+KRz9iMEWYedWQmMy4p
c1e0oflg5VaGU4BNnHIHLtA+Be7SyyPmkZuvmlhR7/VoAsLt1vxzwm94h4UjyusV
LNU758r/cCOzxbRRPS09iv7H28a2BWHkNn8Hfidik82lNVrbE19IXbdmU+X1Ow+S
UA5h1upUoGAnMmnvzSw8p8A6Ai+ny79Wqmlhtsy6D8IRUOI8+C599dnl5B8alXtY
zYGlI2I9DR1D3nfxDJ/zwlK8P4ey83rLRMIE3QeHYk4XdMiy450Nc16t7+HQSL1b
L3d3WLelIxmsH0TDW1XXzMzhjHGRVzRTm6kKjqVjqXbUG/H0tLosIv6gFwzgxJik
TiKqdYM5R3z1nFxjbdHQyIoIfRv69NaigHs8VdTRON8yQoVXwhHB0crxZbtLk469
YDbKRxusBjo9sNhHlspQul/iU7SxtIR2DDT+HVZgd1XiGpFhg5+aXIXvq0Rb229U
nimwzm6L8WNDaRNFOIDb5GCoyvZCQjqoBAeGVvmqzc5PXb/ouh9cv+WAyQwYNGKI
5NVw/vzpPxza1wivdzAdTf2KkrPJ/GvDqy35v48HKIhLrY6ZvmKxH+3NWPlKxvAq
ATsrnEsQT+/sbp7xeVyP3BvInXmnfkUqwTDK+ozt+dnl9gSsQCt7VpnWRWTAHqPt
MVVj0KtXEOGygvQEsp2yyroPSuME396/0j3CTw6XbyGM+fz8fU0LwFehgX4TJZnk
xardg2z15qwxW95uYEUPw1QPsJflwDHFYgNeoQrz4KUTO1JFrX6MgOTRr4Gq8iOp
hlcymxbkO9iVSQsppFusiid4ot9G7S0rM/5DbjawZ5BmS9NlkvSQ1D5Krf7mBhXb
2MTX/4t78zwU8bTC1ckpGWXXLlElTgAK8qpuxmjVjZZLP4nE9ul0s8XY6rDP4yuV
357qV98dNCypqH/NZrb1G4ZeXkLA2n+TKZenyoFFD5PrUWggJfjyRT4N0lkMbzwC
qL3Sv3UALplsOhIUe15O/CsQHJw9J8mlb6w2ISjudGZ6DBwS2qhKlZjij/64cSjP
nLY//b96FaM7V+FHTffCNOwWtpF/X4JvVCFX6Kqn75+q+BDoMnj73pt9jNBwpExe
nKDASnMGA3AjmuNm20vkBWgwVNeC7Ocd7beNs+RRkaBiQlCz90SBCCB/7nZRHTsE
WF0s34YTg6mXpV56+Ty+DusCxdWpVv/f/KtVdSeIw4Kn3qIoOav/E+qJ41VZGzlY
wQwLmxzqc1Rh3+2acySmMGOEH5qOh7K7eb0KCjzftkueX+kfLkikeqLQHeyf8TtL
Ops4PXX4dFwisQxz6A8KDn6t6/SqDpQ1UXm/Xch349h1N8QjZJQLvPDPA5WF+ue/
KidlwOcUncOCUNiZUDUTKtySehaAI+/fYnYgHjOYHd01R4kVdI2zc/dv0QAFLXTh
qRUfLtqjuUlMDVPaQWxi+OmK29gbtwm43RUR7qOpBpPkao+VDoajmb91ai6JuNTI
c/IVjUXvbONg4DtM0if4tkGZtuMaIPTg40FC3ODTjwsPGANcOwhN6xuk8zPBnnZe
gDFd5udPKVV0axT4nO9Jf60+wqP/itoLzEE5bgQlB1aVMH821H/v1INE4CuqG+D/
NJJFayDM6Fw78wMTBRAL9BOwTrZLo+DTtpwteP0ncmebhPOd20kCm4aJvnsmO1OL
W3K60vTnZURl4KWM/PIiXONxQ1tFKJAJn+f74jush79HK3hQGec27X6F1Dllt2+z
doCc7TSeQGUWZ5sJC4PVEPAVIQNFe2JMlWVZPxmLOSSEK04pRsB27sptT0kvsjNk
jriwDcA/VaCusMZWy60LlCXmTjKQw5O2uFP6z5ztD5XSXEBnEzDxL42W7qjDf+qP
sIug3WAzGudiRr2IacYhuzliyPbAdKIGWTpTd8xrBsaDkqn7HigyyhlZ/5VhPlO1
B4HjoIqZVlvirQ9Y+fOCCejOcadVDO05lSmtKqC8QlyBd3rtpzLxuEVmb31g7Z4o
H17FTVU3kLavOxV9kdVr4V3+hY6etg1KCcP7JBpdVF41z44XqmoOExDOlUNx4aks
gp8jF0lmdeuDYTA7dKYmI+tzdc0SBtbqQli5ha0Y51TVZP8KwRZOeGveJLNBCJEf
A8cEaULRjyo4O2QJPbuTfyjOKY7E56x5M/hCufUyHJyytjPELoZlNMB7ENsaFJ5Q
+UMGZ8ARRCWk26KhhObYkiPrDaVvDoe+2M2jPeY7bnsgDiIccRE8XamJ4B4fJ0LK
f4903Tp8i5H+2GLzx5fS5DEtazTjeq8KD6RytSp9wIjzfF4sve+h0pDaJwMY4v0H
9buAu1utwDGQ1IFKOpcHQgOzNbbE2PgCDNdxy22FzSwG0Aafm+7acwEzryawVA8D
8mdod7FgGRSWgWaKRCnz59WOWWLwgDhWZ7RinqDkorh7B9k8Tpzoe3n8PwVuoEpx
+6jrSYdilQvjr5OpvQSteDQFw+5U08ir8+9OpjWXOqp42qoLXuJeGjT5kaxiQZAz
72CaPSyzIMkmfpDnB4cU9cE9+uUMAEqj/F88ELZE1qZb6slqMHi8KRYEumM8AsL2
yuTBiY4YstNrLjBRrfaae5AaVP7XdyIz3f9IdL/SEwcK9PaPVuehIzZkFNOM5X99
PeAXUwBHMvlafBvwevJEuX00zvJD0w6eiydH/s7csYiMDQCIzopBs59+fUU+Xztu
sKBqAnbqlwjoQ1scVwaxSNffhWZrJRPdljwH1UU6p9NBFqLBi4G79DEJVD5E2isc
FlgH15b6aPXCTFsUKn5jYFtww+SSBf29zrLf3JJ0IOF24/sZxK4tCVrq0uKlXoz6
yeYqwsdO2/w/1Vwf9+8mqK5Hp9Vhz2vjBI3MS0vjbRvE6a3kRPpgfxR0nl6oAHgu
IpIihSc5EJDGtXjRM6uHP3fIuNbKnLDeJmmRUq7r8HhBkj4Xo6RJLadB9Q3MVPMK
PJ3dke75IaYOCzNfsqR/Qah77FP+RLvaR72WJYauItXTkkIRiSIiOO6j+o7rc6o4
k7n2AlYYX3jWKPAs8PyrGwI4P1QksiQ2GtHPa+wO7qX8nn+hlSv1GJ0BprybIbV9
YNSSIdaKcsU8G+Q/ViyHkcv6JAwNuy08uSkPx+jc3BljS2r3p2TFk7UFqjaxYiYG
UZj5usa2n1mxfHeVAUwAaNr5d0ZqRagsIKGGkEHFXUVGLJ1w+lI9jtAP9zbYgvgY
wsfGLEBy4BkY5KBDSxjtjbK7Y+EzHORacGc/rZrv0gO+aDTO+yaFQOAD47Vz30jt
+lFTbIenJEbihzkPRaGGueEFFMhtRGn3/mloKCj5YNULqe+BQF+Bs3JEVSdNJ5/D
aK6PS/R5siV/iqhTzwfYMKo8BHrw+Ig4yU0pGbiXEXX7v2rMLr7nnaeMyGixGgd8
L80fWJpOzkRGT2ia+VG4gFm7fILG+I28TH3aKkOyAH6B/ZFvxo5CqunqMUL+QPWP
NatWbfICNeI2sEcHIwUPj3eIFJXnwiodTgcns78jj13EhguGZETlFxIt6SyriJwy
MncnJBWDBmb9MfwxVebRU++jsiEaaLvqagWQ2a4JlulLbF8+7lgJeCefYO2ti/7+
XFJXL+oTiCtw08awv1syxMTlqSJmPDXfBERo0CyVPS6cLa51wIHrT4NY82rKH+2R
plYJJvkXrOtpCfO5RGb54/lioFX37A8TMuyr8sVpsW/8vgnJ5D0xLAYM8tedQdIC
If90Ndg2MEO9iZiEl72I20Z0JWJEKhF068MdhZ79VC9sei7lE8jS2CXaW8xf6AxR
I8GeImnxBd/wu5PjzTzb1gk2Ral7Um1whrJStwbFSWfr4GNvcsHc6rOuV8kQc4EQ
6AF932YapcjWyrcu5KDtoiqPzF5fWfhlvpjyA1a69DEDjpyHh6yo7vCOnblvZa/A
mqfJvl/ZUMz4SQ13BNlpN4tS3N3t6Rg2tt9Ruy6P+JIV14sr6VUzketneU6tj4cV
Uvs1IrRMX+QhkXTyvBGYU70dmI1snGAzpVt8MI1Z8hWgyzz/H95C/el8wW1GFzbS
PCfFG03r6VtuoNPpsfV7JA+0mJm3wxQqMoGFBdd7T4ppdOLhldKun81vZZAFF50L
WlD7busneX6TawZ3X2UFEGUaFRL5ACZWL8WsiuYsblbGhwBubczbhS4LOwKLZXmB
9WYaC+wiaHCgUBUfrmL/K6g2whXbKRT4SPLt5ogdcXl5/2FriseTAc+D3cOeQpAM
ROBfSpS/HMO4jiVqi1ksxivjgcJBpapvaCkoywvZ7oXgcBn+61KGSgCwCBCaobvN
c0Dggp4Hx4+gaQUc4UyjJTj75qWeiUtBoSPh1bGFRYT18ZL2zTC5mOrXOrgLWNeF
PGm+CC4Nl7avSG74YEi6cMTQI6ddpUhvvFxDcJ/LVbBC1d9bbsoNA3rVwh8z/gso
3UJeDW0EIrMemv7QyyXldmdkuyDcFkBO6LwFTCBCMBVpA0SUP0ej0GGo1VrZnXLX
mJbo6oTE9gWq9iRgd7D1r03nDa1z1TjXulgAgyDb+AdhJ7JYOVv+2MvrILBPPOWT
oUG5i6N2fjJDKEzWy3v5hiqqhafywVoZHN5aoTnJGiPEqmUcbhKOGeVC0wh9mNh2
lhi1e/pI5MhJpU/O1fHYTQYkGUNjep2dOOkLLr3oJvvv5Twf+cHn59jLzhdRfaeR
FWpUHmvd/cluSd94CtFLbiSp+pJqVDe2sHUwoJRM3Cp6SBSQ2Za+DxfpvpnWGl9l
A/4UTualE7zlzgrQm7+N4NGAkZV33u1zzkWZ2flwVBsmYJtScokEskzF+WdrVm/H
OytnmJLIG+cQ1m2zPl2CT5nQM5P3HfR0RIfFEKuOUBLkDd4BI72TJh19gtbo+B23
JoUcNHLLF179FWRDHWw+uVi9aKnwGOKCBNNSQsUJM3U5BbEWkYVJcxEhATuITP/m
iPxIoCWLASO4MYviCy+X/52SpOZuP06qbqL6Mv9vxOsWo2jWnf/9VX3oOEvIl6QR
8XBkjhFeXCuE8rMXVe0PgEEaDJXCBOpjNm5ffQf4F8lnhzU7Bdxzi1Y+Sk9Swtzt
vTUxvOAJybYnhKttMjNovWj5B6wR4eBeYmf3tC2Xab5hsUnC4nDvZcgb3r/mr0Xe
OfzsDvdFagVDu7hxm/bECo1wb7nTxF449bZM9euqFywGEkSVlMkVPzOBOQBaykVA
DBwUgaFa0mW1WLwWyemgy3Lk5o/3Za4GQnqnto521r2ZVlV+cJ0MaCQ8UvuZNRaU
NwMn6rEsC7XFhZI5yf91RXA96ZGXbumJ15dCAkV5aemYnfYpI3mBiJpCCUspl2us
eGeKRk5QrjaMW3lcVaXjkqPrECRJA8aW+fdReu5nswBaDU/ZoVgjLGBBF5I1y27H
7DNTpaYiiINMwxC8/WQByhHevehlxOJyPB5OX86goPLG4JbM9iTnMlhFP5blbx5F
MSAwUng80s3jeNrFGZhy63mv+1qpbtNlDuRaYIvm+pZ2EMVjOOK9wOVyGEG5BIcb
fdEFFSTL06g67+UScCKcv1ekgogNp1+CsEaxaOrMJF4FAFrQKfTvaagxLyZ0ZdQJ
M48yh0MRicOGei6+aWhrt+v35a7EFTFDBoIB8Bca72eNDRjTt3omxDSB0mUUpi8c
fwCTkzoNHtH7mJZcChr8lPKweB+QOdjCRVKdNT/HGgMcf8gjfKq22Frf46L/YUDq
khJifF7rIIAcv8NMHsbEb7mUsS6opFKzFdWZpQ406f5B9ZGDvPueU+NU8yv3hkqE
0iXRngaO6Oov/TLF1mMTf6rki2pbI/YZ0JzW3umheH1Xe/uX+DbnJ7IbLLBegNdC
v5orT1mVYGReyci6xtWN0pFOM3q5JpopY7LF18qGsEP++al+BUKb8A8Q1KqQrZtE
4PMRX1OZsFz2HRf6gHDXtbftB9WTlXyzD1emYj1KTUzAL0XCE6mzs7WSYJPdNUqY
FGGO5GC0tnkZL0IpvR1mk+R9/zDY+DKSmGWUbwykhmyTWhNPpxDKmN8U8owVPYma
ZbqjzqlhUN62FoXVF+Th70egyTf6PfGfaBkA61zoMlF1o0/OrLasbY3xoNGEgYji
7YvA08VmVm/qSTDW2OZzgfRxG7VXQyhCYd8NdLmX21/tGZCON9yzD754BRH9amXZ
9bzyD0eNV8fKKs7958MUOMCszMEcjHx4yMOuDgUveYvcyUoWBto1BsNbOwuMQ9UR
lBwYmhgM0pqX3wTbQPoa4NRCeW7qslHjUy7WCwcAWfkwNFxMTRpIoLpBLwjwFrr8
06p0Hb/bvoYNDmwBvcp4Yn1/duAIm2qwMDGzLTvYrcahQGDrtRdthVEh9Y7NTo9N
xfyPg/wlscghyyV7lT9hGrAwb9i5USkIsjIuj8gELQDbgE/WxM5I80RNwR9W5nsR
pJkRl124gHq+8qjK1IFgmaW5GMhbd0E+bdrRtZK0End0/ykmpZplo3+RpLc9TACf
IarB+yIqT69T5sm3V5nfZ8oxbbWLPr3iX6u3VnFkVDZxxX933I5Tz/pezGb4lxZj
lsWOW4Y1vDKk+jCRSR8y82tzWeqs5kF3iPygaPnFdW3Ay0NLjTrEIO6wqjE3YSSL
VU8RvIKRFebh7QRfHhj93i1r8RxLT691kf62t/B6i+91+Mjq8AqAaywMt272oDPD
/K52DgCQobHQawIa4ZZpX8GwUWmvG+xfl7OsFE3nlSMF4RZDF3X4sbhgSqO+kp8y
QX5C1tsCHmA0cGWndcio6tY6SYhmWoiCdElbkLsfPOmsCQp/s65nO62N7qLeN6uc
zACMKYRh1agBgkyK7Wm539PmggABnQaD+ZV1u5B63PqdPKwf24l+UifsKqFCu5S2
HrUuyN/usjB4tJlF7tt2XYhwpi6YbwUwnZ5kOG2wofFcBuBZVLkCO5N9K9C6UL6b
GKv1thoI9C+/KmOj/8ONcVgLrOaddbO481Yq7neiC+Q0vx8BQpEXXgATTU6w/OQd
rkUYX8XzGRat6cHYqxnkYjSHeG3DDJ8LrhcHhFVTVXYDzJs8LC082vgPZoC8cEyS
g/ud0Kdhf9ZEr+Q0MXbMbchvk63LxgvpT93tZNOu+WanWINBEqlL6iSJw9qVlEEJ
Z20lHue+6vrFEXBH6dQjBXZP2YOKVQ/fmI5Z4LawUyaM6R3ac6ZIgsLznIHJmUFP
Z2ijinCN23cJ0wlsbcCypd38fDEjaHZ8gAiUUDmvJs61uwo8ofXbNQYY2cao7WTo
kijkjfSvnSzKacyMOCTYpBzMdN2AUMUrQYyL4gN/OBFVJupv3t1ogeiwwUYRZcy7
O5i9oEzOKepAQDClMO1q+5/jgxdSaQ8J2bWErmVIrLEQa18gwAGx5rAwqOD22pqB
AgWdIiIfTYlipOvMTBWYmLHoOXtBh2TehcPXq4730oR5JZrmEwMP8P77AhT0OC2f
6U6lmuE9JvHcuHJV+mDwLkkYK/V0KJVM3HVqkCA+3RiZPWCAvrfV1zI/UCNaLk7S
yXeBiw/vDlFcIcJD6tGHr6tvCKkcBjb/u5TxRm/T07RkDS4dXjKjBDcIhhK1Yoyv
wjET93zogy+THRAjhFFK1qNqgXemzFlG7r5xi8YGmi7aVO92kqDf7fwm490rCf3g
UHQFEmuYXvx0TJr6M7rkZX/1DHMXKorGEsMrGcQoTrNzR1FDDzw5CI8VsjA/O5z/
i4brQKrnlBsha+AEceM4jQLF9JVd4AcOL/MfRZZTXtfcu35XrqiJu8Q6WVHuBetf
WvQGQUyJuohQ1hGld+doVN5WaWSxiRpNRMP+XHd4r4EROUKc3R8+CLcqme96+7gv
AlA8zIEANY3iERx5vOMXwxWC+zszf4CiWj3KQvcu99Q+pSmRS9O6dSkv0H2Dx+6j
o+aEq7wAa39VDtr/xvJp8qUN1TrU+bvQip3++2ieuLEUeLppevX/WIpzeXtDEEfa
0WTuC7+6lF+ZoRQRHvZWac1fYYWUvj6H8qSHJ08aN9KmNDAa4DTYGgltd3N46m4h
5o+HLFdAu6Q+0oyQgkuAupFfeb5bIVYsAnGRxbfFkCqGUT5dOLlLQDW4i+3LcKOv
eS073ZnIZS2+P5HCFquPSlLRKVssQvZgCvpx+drwdxovTUm2g7qUdmcmuDpHAcSD
gejPF2T7mcZWRF1O+CHR8JQtUZvrMfbUcEL73wrosAHOvYq60yahYuzA+Xgkxzw6
Sq2dmFe18AHlIu9fV17jtVlSa18/lLtcad+QckhhTu6x4JfnOg1THiL7U38jQqjJ
B4BFi+wMDNuBn0Gcfk0ZVPLU2X4S8fxIuQ9mA9ZkfUHDV5UTeS07Y0xLPbZoI5fI
6Yhy6vkpr3UbMjJmwdX7KvE4JnzmOSibLeLkBoEkH+u3i95AhOKnUDOyHwAC9xDW
wQZgbrVBkOnzwI3XaeU1xgUZOx1pPoomvlHWoYawsqu5MAgx/ZHEjNOykoJGwA2i
li4lwiO/RQMlFVzJMoux5UNv0SeFlx/zVZQKMtXnaUGgtFDchjFv1eag/ghGiJCw
oL5r3Ay69Xw0n/MxRNJO+8bdzSjfckg5nA7GW8Fe9q4E4qhjl939A8FQa1st8Vn7
gLFHMLY4FQaXqNwxpvy+ML4JmoLDVGd9dJR8wDfknpsOHYj5Q3+kReIJpmNQ8mYR
17FFyosv+YUhu+BH4rLp4Ml1LDFu4V1z0JkM5cVRpOAJfIOYTUXXGM+E1iQt11IF
DW+oyG34MdgJQWqK4Vx6qZ3gX27+tH5tYV3Jg56gzcD52PDCg6kklUKLu4y752Qr
hpN+Df0MJsMcZ+LkgzNLezttKpVq3fJaWCpHdyCx/HXYc/DYqeCUq04MX3XkpcKA
TazBx6uXR6xp/7OJY1e2X8FuGjX6bxGlUtqupOn0Lw4u4S94KvNF17IKMiUk8Sql
VglC+ntHhA35HqE2/lz9qOHnG817gmSZBfrZqAutydNE7MyAeau1swWHblek2JCR
hD4Gymcid5Yg3Sxbu/MmD9BZNP8mShRzQ7oAywnynUg0v1E5j5srQi5MHBZ9phgv
KGGw/skQu5TDL+C2IdFTen/NE5TgtCZdvDkB7VRO4czI3JFJeeVGJRbecRkj6OZF
uP3p1x4L2FLeV8dic6pvvuy6C2ReG4ly8TQuneysREcu+DCG/JGF4LpGvA+ZlvQl
wTYt+4mKqMbiyfbnFMhXaG9bHDQNAib6qPdEoDqDi2yEF6TsuCKvQuzJiOD1v9wT
gNwqS54s7oMSXmjNtCdeTeUaUeV5hbIsZP1qSQA4Mep9UWtlmL5LQbjdLiyLa+1u
nvSAw7vNIMeJUY/OIc3+4iZYNA4MEfd35OgYjDgvCkHEj9kRM8tRsWd/DCe7shcW
XPZmxw0LAj51bEyqBkpWc3+5dFIBZfqvxBNk5wX16EsrIfCprbkt37e8On5Iz3w4
TSMLhIQkqgw2ToC7IWRMQBJUa+g8i3gmz49+w+TeQ4leq/5cQX4InOMyI9YzR16+
UOxB71xqBjc2j4CTXukwYt12wBXZH/vD/Ixbez52TF6J78TeQf8Dg9QQjNKW1QMK
khzQzaR5K8Rrr4bBko+31FZV7FTIlx4CjU6qihsmaImm2vbAVrxVrVSnOtGAHJa4
EXWxGWUXrDdI0c0R9xq2Iu5YdwSjiKW6kUUc07qFUEQhiGkJWOO1nxZzTMGfiOYB
QOzDf+gEQhKz8pQE/6kgHbz8flCwCpoRfzK4yfpJtfbbTywMUGuSSG0zz9R7BBDC
G36awu8GHYxhEq/sM9bz0k39g04bPauD8YW5to9ypg9H16EU9HXfPQfmrj+agsUY
k1Btf5Zav4BBcNU8WNPfASts8DYfWl4h2ptPI9vRgEpkoqYePtVNJ9KHBvqdoNVa
vcv8zaSVrQBexDL9PRyir8pBlZ3cdUybR2iDmJUj/ZkWkKSa2PKQXuo/H2/5g/pO
GGvtPTkVKiuhOxnQoesLWy0EDdL0mmk/5mny5ABK7ReF8wo2tEYHMincDMYYCTpu
ANOZdiuKRz09avvriirycH5Zg74gZd/rHVo47SRNLuuS8M6UAG6qLjYWShueC/Cc
2C5KLRUhXtjkcTNodbmhMt7YVdB6sZ4EUe5r6ncAJsBCLC1Et3SCgrQAVH8IuXMZ
VEcj3hR9bWxiJNM4EqV1lkqIGPHAiYuuS0fAMuOR4OxVCBoryZRaVVDGBySdNnsc
OGzb8Hz9s3QPNoOTXnJO/OLPE2UFn4uW4eFRiHxq04uJb0697yAyTqlb7M/Lb8St
KEyfEEXc8NyPmpHEye4lV5fK64y9be8FWHK2g8po57zTk3R6UOovgIg1GAK0hvfE
5FZGZ6muWQgO4CGEeNJILSoU4HMC1zijyH3K9RPpmZxjfVaJHNMonNEad3Grh251
aXAfoH10HWCRPGINWC0bGVL8xZvEG4VgainxlNekzEetA1ewdDEffnMCHZIhKjPn
m3rwGtp+Cr708hxePlk1w9RP3w1brFPqqiFaYRIDk5yqaSP3+a5r4kfPhnW1JDKW
bpK75BCdvILsjFmYucHafVS24BzTu4Lup9lNL/vABafJ3kcKgmNU6TM01lWQaBxq
3+FGtatWYx9Z+1IgFmzk5Vjwbd7YM8ZciaR/JETgWTidReojrAADVVCEZ5WZf5Du
gWl56zDa1Szruj7tbYsV/d8ZqgNcVT+7bYKYOlN3NcmSMqVh8QSlya8MUn9dHtrJ
B/62hHXLxru9vCsELPg2dYobKUE/RbKvbLAl4YsRLTbadEJO4wzwvP/uwE6lDPox
xtl+cjd6uxbQTXc0Opcq9Y0NS5VhWcpGjMSL/uWuuoKQ11O3zTcaNRtJT9CzN+Ox
OS6Qr6agsNhtAA8K3liMerdX+gvSQtIEVJm6eamh71HWl9h4f+Xv2VKKd2sjN52i
GhTX6X5PJoy7Fzb/nEsKFr9R2myaShw51lSdVAtXzSb6UqOlJcX35HyyPVrYEBtF
9LPStlvlrpVJNmRKeXOrTK+GtdrMPBeieFv9Ef71BAaYHZkadejgnu2byY80yioj
JNaKyGoZ9z7xlhMateDZb5I6zi4hiuEc/5O0PRw7+KKFIM/X5l0Q0w6odK+4jnO2
511FeRsWhG2xBq6CMWuEW3VXKbL/BqZI7NTSy7rbaj8/oVymZkFficOupBN3tVYf
InrN6tT/mrAXtJtW4+lpHS3rT+nXMqEa8PgrkyYi6CAiilJtr6fI3ylDNHqlSKGN
mCa6XcNqU2L7xQlJzGBT176Dy0CQ8PGDpdVYzEyLFQKvu7AOBlW2bpWG7fhScs/E
+F7YCl3+J4WImkKM0eioo9dv1ga9R+8MoiGO02hPmvnUrQXyUwtMf3havixYzRfv
Pepp56Dt9Civ+Nl56+9V3tsK8/bfFfzImlD9Sx4iyY7exO8AtN2awSAltH2HewqL
mm5tZ5U1MxRUt0ky3+EzG9QX8Dp/TUVRbAWzBX0Zh6qszYAgcRitExBuZT2VVHDM
me8A2zIpQGhrNBdLBiLGwDO34TejhmVnKH55XMbFKeNFOwjF9SUhac0KG3OQDEwD
nUSY50IHbknbhMyn4+gqWUBszWGQqx/4YacUf9COu/Ref5kJoQA5WhLUZBcdZyRN
hFQLEHuNgpDxlLIj0tOs7FQNpX2nUDm0KhutvV+Ew/KjZ6VNwEc26SZtyDPD1bLn
zLkYDISNQav/GjMmmu1tfT/KYB42hIQGe1AUmONozIEbX5rn+2xP0UhM7lDy0XGV
5JrkuvFYKXmiDLvjUzm8f3p6zkgDisUUdrmgatTb6AaGBcpXyz3yD139mi1sZGxm
sEGoHltFlNjk1YDf+9/pfyJipLy7dr9KyMqJwNG6YSr+XDYmCNbaHvT/BkEW0za1
aAFDPbToTITRhbxuDz3mYDI8gMfVmKDgT+BTfgfaaKWatWOBpcyQotRjtZJ/SRiN
R36lTOwHxoqgkJ22fRLjkz253yQEJmBcH9e0ZFaCesmxOruk5JLoFAORl1eYuqva
0g9/3o2SsDMVnGjFxuwMtbCpLxiPBoKCq4gswKQ2IkXpjQET4eMReb6DPZZoOkKo
F8iUz6TNdyGkQSUhicfjO12fOzj7Iyxys0n59aio3mfanuC4nh6NxrK338tidWkr
9zw+FTtdYSvcpEBUDD1j2P2dm+Mk1kZT9EPc8lddJZy8BqAlVqlk9dkimqwuaHqM
/hhnpaysrLfyYEr98W8/lThEd3kVvEVckn7h84TVr7mMPJxVypMp5rvA+s6ua0el
Eyfer7655aBH4ASa3ClnD2vAqjwshNP9slcadrAbSRpBrAZX9rDICmzu1SYE4UCE
j4EoT1C20F10qmLIF5tGyLWVBTbbncj/gFQh2x2QqLeIelbO0IPwlZ8IhyJOm1pP
WSrZDmRaOYwG3eTB+kF5ki5g5Nal9SjjAXkrUb02tzl/xbX9ejFqPXsqlXaI08CR
EKYGpmZKC7YzTMx2UcC8cWOCtT1sxiJcNSK55xsFM23q2cTux4UQDZJKVCvD71CZ
2MAIMkr6MrezIvmFTmvQ3Z4NVDUk/Jv9Hwzx463umDJ3NPZCUFNu6o+Ns1vg9FZ3
Thug+jnEdbiy+PbDDEObbu5u8mJNklavRNsHFL+ohOK6jBXkdavEXN/HjtEBVRwR
In0buL6bp/MDTucwuhLHsojO9H86rbK7FwaLJAMRLBSR3G1qNDiK5XHEYwc5utss
2PaCCwXi69VxvsPTQrd3c+Hs0V3uE9ZseRXecyWu3sc2e7S8INq0TGHy54XMKkEP
dPKTjD5d9ZMDtwoyuLpes81HGIRUb7ia3VNQAJo34qrXQursFiWmgdm+vQZBNZ1U
zJJC42NrWOpntTTLORmnNdMYNMxNSfiPjFZ4okv+iRZSzuT/PE3+JJxpH+yZBQF1
VgXqBxn79VnaYn4Yiis5g/acbl+hMRcQYUTW0UsZYIHMeSrlbqgitzWZRN5NkN+y
G3CUgTmXEX9QaWM5ZH2ONVO3FztwdHyeFjXHSQJFmaS1xQh6ShBDlj/LjQ8ZavnQ
HkYMzNa0Fob0hRcJj2pTqXXd/F0e/Ou/QO/3ewz7pVNKs0Blf7DjY4HlIPU73qf8
HLsElznFGBhS0WdFUPWntB9CFg1Vo4Tsr2ByHkBgRUVl8hXz4i6/Z+NFxr4ph4xL
KWnzNVPPhV2D4BTmN0WdBHts6oFOpKwYoaMtWnqk5f5/NcnA8Z43VsTe9zMemXwV
zvc445A7ukwKMkPdHTaVJGwopG1YEOqBpZMZMWj2RZBXkMGIobRuJnbxzAe3B1rl
TeF5DpHYSIiTa/QntoGyOTonwxnxfsrrMBRq4TSI2uKSaNWaLU59JpBsp28bgoRm
U0essdvULnHIqgOtrU382nyWDM/lLSu+1+Rpz8Urb7qDW8NcYr066Ayha/GF9XdO
R2p0N37iRa6I/10lPLD6X3s8n55mKTgvv6NJeuiEsTIEEN57Goq5tXj32EajEMAu
pa31AFnq7hMZOJRjUnzMxcumZq+m89c3eyHrKP+N1bHgAQXSKx6F3dQiw+EVzoIA
6UloP0vDiKrdEiGiq5pI/PPysDjAhKwbWLmAg46TeW4fGZNNsS0ytysjpugspnQ1
xze21lois5ciesa33NG+mwh8tqEPsBzssEQf5D2CoZejV0p/wnpuvYXc++Ecodd1
JAJAxACxBkXewAS92VSQwE1GtFw2YD72OcR7ZPcae+M4HX3yQDTDQH21hYgMyWsE
f+Ud57zxvrXwHaDHI8rI8o779NZ9Qsu3tbGD8GuC9c2ElmQJk2Rc6AzgtRC9bmme
eALmtG9E7jWhTbTNU+ppGc+qzDffoigPCjamccdlVj8VhXZc866j2NFQwx1zFGqx
gBfjkdU3yRyp/bM8jpZQBlv9iDPW9EYDRhDAwgZVUosfnw8AdKRb8JdQgBVgd+Bi
5o2DTyvJKkA31f14ehf1r7lOUVUTY7jJkaAIRywgssVNjtSUdEb9tyo2iua7iOFl
mD0JqINYJHgJkPxOtiLnoQGea/eB3etI6y+uD7r4oEQzguUGTAJfn2CGkiDRX73/
PqRp1+ir6SzD34iy4KxOZAnnTeHGftJurczIgRKJDR+pXLiM/v0fewi2VGP4pvTK
rzKJTkTp6SJEnJWhAs2e6+fA1RkxHG45IjX/cqwSjaxBFgQAH3TIcjteSTW9n8SH
eGa6ctUsdeNrnG77n3P8ESjPB3BkhSlccDeFU6iEzPLaEsm72hInho+DOOICnPhe
7/HT5miA7qDhvlTJtGlPMfCix9cY9X1gfVmhVjaGUsidOGz1h1g/t8YbK1nnfFzH
VLWAej40TA2cJOJwZXD/jIy/l3zcT2fHC92+/V1dYPhMzyIW9+ipcNuM0GzftIMV
V+jlQmQyykBUsTbavIq93+TbZzrWC9O5wxAkHxMiaVPWJfto34TBdRjYIHwBUvcb
Kh0iL1lVxTcNT1fPFZKsmqeEpvwDn3VdVbLLFIf1EeynIaozxtvKmyEOk566EfMl
QH2Kg6HlBmvRx8uT2gzqpQCMAqGBA82Te6x5VArb3xK5eBpQ6HtuMPAWr+PHsSQH
1qj+lDi69AaOlyiUZXigxQ4eUQYkjNluEDQe/DaTcS9KT+74qMCHjAEA8Aw7LdPS
Vl+mYmb2Sv+4eBorIhNLtZdn8vn6m1X86dMGchSI8dU6VbaW/xEr3SyGXvSjRVfs
RVHbfxTnAPyg2kUrhPruJwLIRXMWN6SVeZWt4ZVyWekq3vqg1cto1kNke85/Pr/h
2Sqdy4hq6OH/j4ICBKuT9eEJiQnH9KMEzDVoOnoMLqWPNhkUiEzUcKSzLJX+A3LL
ZvzUT7i3p/kHHnhlarc9D57ms4RHsRgOEIs40PNfP8jkFwu9LG/RUsh4UmD3ONyH
3Cbje7Ge7VXMc+cbXItLHmf5nu7JPJGe3OqNbhY3ckn9aV6CpRP+XXLI6WQ3MSSS
t/3ClD57d3vp8zBXxastk2I5YMfAuimzSfcOD5uKfw0PlPg22jQ4MhCpaif+L5Gc
Hc/LVG0pix6e+0JSzsJaE5zG+0ju95y1d4QBpRWzo+6SKOfgYK/PRU/zCCUgxvCD
/g5IfUvcMCVJw331UasywcLEnhtD+xznxQJcwRN+1jUEwrHG2rCtd4c24QyYjSB2
6cNwfYXD3WRAXkDnqqMivz5RZEH3c2+xf18G8VPlCTQINROuA0OaJV30NONN4f10
9jVGxEuHts+8JHoGMHx+BISqJn9myVsjo58IA+p6eET1NrNL68OtDI+A0w3oOMo9
B6IkEFBCUFqq+hSI3unJC072+znRI/Ue8b5n/rx1GbxcNQflGG42xIrYkkunvwlw
QOjXGiYf4YcVUqvkeytjNYOOhNocA3CTXRGdTTSqzlTnroHm8N6/II5vycCfVD70
X5AetXxNDBsP/vivWuEOeCuHN6C+Fald61Ed0HcCQHoRmByJmRwbt/IOeS/qpQM5
qfrWxweneC2q8CYFd2ks8WInwmgXhG3mvYU+csHb7G6Lb+bn0vYLBgyiy4U2xyIK
6sT9NKMpHtLC65HNnIYyEiH2VBd7nNOTvWyogiRtCtF+CezQqQ/tThK/Nxa+NVhJ
V/gyoDwqh5wO/ShAJR3yBSh/B4hOkG1A7zAorv6AbFKzuG7Jc63L71RbL//SGFhh
y2/QqNbMA+9xLRsTH31ahJTGimaA0r8LGUku41vU/zXfIloXTw/YkwNWrzCMGMHy
4kSzvShFMnPO6x2zzvl4EASiYuAzlu9k/E6wczKXIl5vZrIhbxD0mjo5yyB0pXrt
mYFJGIAaF6dXES1FYfynqmZVzXf4ecMY5neJLP5LVN73jYPeaRNPe0AiGY6hIAVg
qivMJxI7W/weWoig6v0mBWSRJ4id4d6YFrKo/C2fdhDJz8zMMz/WEQ0FpWcJHuiz
dpEI6NnPpDgNEdJTlWWuSRfD8X36g7Bx2CpzPvWOtAZQVz0Z7SJJEZnDrIXYfZtc
9ie52oLBaJLmZrl3bNgjgzIRfVXbITBz8/N84SBIvwMJbCtadnDkeFHUhFJawLNM
aI+NGKUuxX4f0PIud2U8v670ui+nx+Ewuk9Cxq3pcol7caihQq51Cd3ArpN76xqq
0baF4NuN7W/S+WRP0s99104uhB5QaPVxjhKx4AbEs89ZRAON6FZCsNqxoxcERx0i
pjnfC7QEBgupgFWOXuu8I/fsi8wInVOYenJ6ryGYMfYQ1xMzxAFiEpbsdwPtjBgY
hYAGcCQZMwGZShdfDtMy4ITE2cXPoa0qt3ph1jt0ekrkhaP2g1qShoCqmkaEs4xQ
hq7dVX+4zShx2/wvVLkiEv7iFGlcHt8Bwp3uLQpNfRBc0wHf26hJnYePqN4rNPId
yjM2CJd3VLQBHaJBMH6fTn4MxTV6wCWmoB8zuWbHh2eu2M7X7d3Wfq7+yVRMaFCV
NrwJt7i8HUb6B40dj69z3kXVIWanjS8MUgRMNhRA482tkWecVHvoZZa2QPZOCb1P
HpjbDwwScw2j0dpdGmTG6Gds0gCxpl/dr7grvZsXcNBDOPBo50yW6V+YeshvTasY
7nADK6uhuuwpp83Z/6G+vyIhiJPuKYZyvNgvJl593/tPT01dgthXFgNodpUsWUCv
3X/ABfBg2dhfVrPUIhvKq/g79IxoWcJfnOUdH4kC6aN3Zki6C/nO3WtLa7TdDb94
03yuHnSwYH6hlehUeMOOAEW/Km1sDIDFwKzm7gBhaqH2r9j1L5G3sg7rYkk2CrL6
vp5sbMSVBvLiPCKl7bGZzwNXqJEQ+O8yZ7bgQ2IObB6hzgYdU3AqAZS5GHD50+Jn
VUlBXBrDf0Lu1sFNgBYipDFg+c+o+ajeQInv41tKueo9nRWa2bJZ0uGsxZihaRVM
X2tq0rswqB2e4sHteNEYgKLHT1zMZFxU9OYJFk+6KEBJgHqYFTnl/7h6T0+d2tYL
2Jh50lyresQ4SdmTwod1MrgW8cP3Q+wTPfN1q/3DGIybxGoF6F/WfiGj2U/IdR0H
7Chl5R3SmO+WrcxYlI5KgRvGXckqwIrWDmyIJh5RkCKiU8LETmgnEg91ZSVk4MPM
oTpXrdrrnxpoVM49Ol/nNW23g1cLymKigEkKCrb4yPdtjqdm9EijH71qt3pygVm8
WmZ/wFUiO2nyp7l7qoqmCZlRnX+9K3Y+L7D6SI4321Zin1nNLYNj9zTf8e2tgU85
2lYstwuPs9cDhsHw3gWKcLHTwGsRoKcF3vvf5YLZzvLmvLqjGpLc28kBEmiDYuGU
EM4fKzh686FXyOhdVRIYlPXYJlrR4/Dpo9lvgoLW4+irsmTvOCAyS6MgCq79ycox
mByXouUHB34b4YTFv6urnSzDMzXLq6UvrjZ6Rw9LuCKpaVE6SkwYdRSSMfSQ0kZT
o9dCW59oLS3LdL3t/TCvYso7YAJ/JyvuuGbKFklZH9h00/IPPar2OMXPRsiSSzGv
CmB5gBe1wteqjnCzmVWiUTSohsk9UtsPEAwtrfsZllQM8M01wL4SbRjIaGOXJaGB
2XmoZWx9ZrWpiO0dlhyZLUBOhhXUeaBI450fZnMpGAlZoHqJS7+l5e785E2NJ99v
hRC6vlldFHhMomMVutOdJ40HSovd5nJ5nueynINId+CMYJdiysTkT+/xsf5Lop/y
ue/b8z0GSllqIdUxSnA6wNYU/0LfvF/3x/09CbUiak0oilxxDODAixiNqXt/8L8N
qdnQAKCELauzNaFd80xY+Y1FuWOgYyTkAXeUUEarJUurUyPAHRNyxwClAZhtXmXC
4CKKckl7g9gvY7q5TR2FAA2wyyabmazv5AY131oN+RWcvyxHyaKBPLzuJzz2fKo4
3vwgphXXkDlyWvU2pk0TCkO7kI4g6pn6Ju7fuaEoe/XYQzmwEjLQ4ItBNaAqxbJN
CbGGy7Bz9SLLcUQZgbVkW15estRqWeULDvwvWfWM9MRUeAFTKOG6uiw8TIncV+pj
2vnqZVrJX9AAFFYUVFByXsYOHVwveU6t9owgiAc8M9dx4i1tgl7kMdTuGFv1Kb89
hthP09qd9OkJpLzj5ZeFh4xiNfwBOiJzeOd6uTcZR+WZuy6o0ONVQYI1j9VjOSV/
pvutabjo17mQi0FIQWy5+N4eDIo9Jr/DS8dsL3j/AAvDKwmq3P8QI/PT0qsg0S+0
CqQTgtgvyGsXTetOIkmmKgPHWVckVH7+RCiNyum27PS4ZgvEI/89OM3w3MdKlFY+
e5LewF3Qpi6w7dJy/b7pouLvNsYqCf7zZGKHfEy1bS7i/YKzjPAjFesqpB5P5pVF
wELRyJE+bXas7TbdPDShgh7xcFYltmAQ/QdtMtqSV8S7uVZ7TFtBZurdxkZNUDmu
zyqFSNfOWBuvzUBeSYyjsob4n1G6BJpUMHmmWCql4QhP4H2HtJ8Kv8pgkO4h345r
daCIfN4aEKqTOoyKxpXZ6IXt2f9DEYtG8eJ6bulDqxXob1eNcmv1A6oEq+7e7J9O
NXwdbRlfEA7gNFWo+SngxX3edr2QkmQ0GiCCeEBsqWnAv0rS5o3NuEFeLdimYcKg
Xq0PJv5Xc9oE0rEIW8VY6kYeDjd9uDR9j45EJhtCIz0gLw9ZQQTqlK6hKUUDeilK
/nQCbf3vdMJRBBFIlmHD1U7U1l9BWOzy/KLq3zaH8Vu2a3kEXQvxiIbgh/esUnm7
7UAiEgs5BXtw1iIzGitWlQmWK/mxI+OIWSCnnabi462PMaxbXTpM1Jy4GqaztahY
ltlJhIJUoM/xTBP8sEwR92aaKHuMXwL4ZPRfX3qEHbos0DQLdayrkR6B/eOJ1qO4
HoQ+eaHrG1Xv39h/iNrs0fssswGbX3rr3IErCuRgKFfaMtk/nSSZGBADqYOaYU7b
AFg+5CSSORA9kERDEyDYVhrL3CMo1mWR4mxMqAhLNdsBw90k9qmpPdfRPfs4HWZR
wQVXPn0iNH6JUZoTIZmlTEZAoH2wIXNlKdDIBX5o8vHbXX+3KA+wUNwqAaBhIyoV
6zVuE0+DEjDixwlfE286cMGpzwQPbrsNxQNe/JAKKm/WaQ8caWycTwCjm6J7wxIq
SG/i06d1YU8llTVHREfYE/UAmWaTWywPl/hUHcnk4TgUXCXdNIiR51eFNHLQGj7v
hWOjw5NuOWKk54QUihZ+S9QcEtXexbk30XQslEpgTWvugrTUDeSXeuJqhj+bsePy
Cq/UGNSsuTrjpuCBTSTKGq6Nwv3SjJXEUAH37r5MCggBpK+noPOFP0yvIdjQA+jU
Z2r+X0dok05phjFp7wlO0w/SmXo+DyR1OrcXZCmicvn5UGzQmQIi3FfrPLD13fNV
FTUur1ot48aqKV6So7MXdv9ShLuuzIXynSbtevzFr+YHfER2bzh3lgeLxCHAAhEU
ALegD3n0dAvDB1r8MB16n7kxUJ2AMgsjckgdXP/jEP16OuKJXxEOQxUWygf4aIdO
wV4+uDop6EiRMl2qLWmSQxi/I3XWn+pvmAxuVYA7rkqo5R9XGGnxXR0GCLtUv4Sg
oWu2ubG4GJSmkUmWb9IDREoQx5F32/1+t4Uu7LhgpRJ5DbnApJzfJ60DvLlWYqYz
RFU7MtaWm6lJWqPJzN49JvqNiZKvsLeORku8Au3nB1iTaMeKowiLC0/LZdwnETAy
bD2mm4ScXNSg89j3T6sz3Rt7YjHrU3dMRaII1sTEJ2iBOqZvLCuXc5tKvJrNnpPC
mEBAmecVcr5fpL4d0VdTXtt0QEsxhZXl3KANhKKShKpnts2I2rPYeBqi1Y4MQbzJ
WdCL8ZRyXIjpuAOn17T/khvCLQB90mhvC8C3i5KfiNZghYd8/wjTMRbZx0Rbi15K
NIMYrEt3hAH5HhJ779YEcM1wqQLebxEuzPKmWOJ0gMsaBjQxK1xPo8MYppc0xjcm
GDPjXjKOtkGTYPVh4uLMQ0jLZ57Ho0XJAa34S7trMrXTz5J+8ty8JFR+Zf4ETpIa
PUe2ZQkJm8BN0wg0hcYDUli/V2/k+Q7D1rffzKyAHV/hcNapcTcLaq6S6TK5gK1P
T7f1JE1iMNMfC8mA1S9T7lowJ372OZHPjKwYPXfn4G4esaasNB2jt6vnLxlwMCkq
vF9XG275yk4OBBaVncRJGGqS+zHwDUPWXem7lMMNMVbwpXy1ECykOJnaOvVijDau
jysktYwBTl9GL3+ID+ps1D6Z3x4srDz5nJCMobVVHcj/6IHY8uCmKkKH0fb1k1ap
h+DcGj72EyeJmE+IGPPXJGVldXRGEji4lcBMjPcqryE1A8xXd6+AbYygyDxVdEbx
PWqxD5aFUnXGspHcLXc1bUhopBcxWxl/1QJjBPZmwNEy5R8mDy1JUvfPSQuaVH4G
fg8RoUKPlGs7fL+I5v8yuVDMmnpChbgJ7iwFPCunEm2U+cz7l6TdYGJB5gczwfI3
ISg3Q0xCFfce8Tfw+E+lWsXX9BEnMW+BTcH2trRKZnBNej74QhF3MB4xJLArO2tf
o/+/NdiKZPY5uE0eqBn00fxv7irXaCM7fW7Xb0CAZz+R7zUDf/dWQaGpdnLjvJn1
+Trk6eyRppYgwa1T2kTNycYpW1OOnywMRMQoNEvTs0QGqYU7FZXhgn4j5S/bdRjF
OfswvibHKUJRmQwgRW/mTJ28VLsYYah5zVhA5J3YZoKI8BQju7wKonpnXPLxhGjO
f4mkPykRogn+tndLRYm0Z2Kk4m6qtknDeassnj0I4Y4ZLJLOp8PfsFXHcp1kSNv3
USXzM8JbANCIOx+iINZ6/IbETdDwYEiPH0+mzB9v2YxLt8WKPBujoLff2v5WVxuf
nlMlE05qLAQHkK3M7H4KeJCQ/1b0GYMpuDMalQFod3DYqjBv1ox1pR3pBYpTw+dx
pT6Qvhc/yQPLflLOPH+KOqfsMbPLR37EhSxlVfHF255bFHl1D7iCDbaroUIjKmP/
GzP9yUfc/wW21nElxAXt1xgM17ZohymJ4F+noPBieFA4NMkLuoIYBqBSVOPIq7rg
YddtEPBFN3XWnITCuK7uzZ0LaqllauvB250YlUgpcQ1nxk9CRxrivDeQxxhv8tB/
TRfFfy779x2VMZRA04Vy7I/M5g9MDwyZVAbEQMqGufgezA6EreGC16lEecXU/Dot
HCOWvY9Qud9Qn90jfcjX7SnCo0cxEJy+RyjqJYaIADlamWgNuUdSNd23nwRs2atP
yZAz87rzkBIeQIvIYOOBr/mQjO4qncjIgd3p99DJq3W6wA32fFucyJspyBa6q6Ho
v/Qt5j5zMPESOjIPKtvXVT9yuuurqoHmz1z3EFzqp/Cb29Q1COhklWku0aIPU7XD
tEwarOeGBghvZi6+r+gCOnSbHtJcO9QGLf+gT7ZmTwaeFe9FjHvk75IDh80UaVxn
w3bHxVLSJAfBQWNnHN+AZB3LMyAfu2gV4WBE5A9PPLGHkDd7m/8+pmrOSz0fDCNI
kmQ4N0CO+ynGC62cfuEg7uL6CK+WlSjRCvw/0TxdgFSO1cYH9Bj4y8JCPOEOG499
9Lw6Gp4WxbXlOOOl4zmlYnXq+Q8dAM2HgcfxOg78WGi0+21kON/ZvPvElCqvuvje
ljLWqASpbAuWgMhPvocHbRjohtGYwhy1GUmYyYh7pwGqSXuqdDdEn3jPd7LBHT1n
/uIKC+AClzuzhcCBs2Wa4qLCGywiLVnLprh90sQad92TzgFLS9lX273c5l4bvhJX
jbIVic1XzIOLLDf9K5ztFIy2TLID8WAK+kgMQTymuqtWPrDXKO9ENJpMTaCf/ExG
vPaEOsREGIa2nZM88EnDFfN19ptNC9Rk47EqLmsUy8XdygcVGTXLOsoN/ukFk8lo
3R8BwwViIxAK88+pqZTnfB67VSsQoiJ6OrbvrcuPp7JNEFmEFD3Zxh4tMc7C7Fpf
P3gqyKXZ7oTmMbwRy0lkrxE8xppy51vzGUJt5U951FR6xxtE3H4l/GvsSbBxsvj6
lguuuyW539KexwMLT0Y+80JwTY4vzflrBGK2MKRQP4k7dnY3WOCLnV3BEJ9Gg4/U
J1l53QUohL389oEqqBTULFxlFJ836u2uAzj7YzkG7UvunlCGGCX73TLxHxZnrbqG
Yu4SH/4z1zxShDhGjhBPdbqUnyg5UfEMawYtRMUf8F6ZhWUG+plpL8SYsq1HSowo
CVAu9H3z9x/eveGTJFuKpCcxhjC2fonUsAucUpx+Xm4t2I48/VxnTsJmuUgQqk4o
Ybyukw52Dbzhdl/91S4+1CnVQG/7wnSINlyu+v6XzojmbC9N9g0j3tCakyJIWImo
WbZuptTOYEDdD8J1CPf0Izl7SZcva3jfavCEN0JekaQBlpWlUdyE/lvuM8luwkm0
NHgqEQv4pBkknZjL5HRxm/PFsxYua8P9NamJYbfjr/INpB4lVCtliV3H81ARb4HT
QI9+68svBKbrtvvXQPmeypfI3Luaqhz2ftN+VTCz9MDtXRx4YNWjYWxmKlTsn/aR
th3IJbOYLbFdAhb0CwUm5y/cnJwsVw57siWNUYO2unaK7M5w/hggmzUbUIGV5RpH
hmt0yr3saM5YPOKXi7C35eRHGt/S6xTus0NUOxDJCDeQpJZ+2mdSO19pj0CRLJhq
qo2NPLtvsrw6OfH8MapniilmwHuR5agK5t8vQvwnYSyzE3LXT7Zi5NKCh+tY5eOr
PoAKk7BiDeY8ktZ8va2byXgotzkwJB8IkvG46EddgVffXO+IUSkO/P6b3411nu4k
txgYuBpeJ8sNszoWJAtFX4SNlqHdFY3TYbqLikghjsH32a2vW4s5ahLpZrEbrNzL
9CYBBfSCAfhYJGaBdUTvWvrffsJWcebyLQK/25VUx7WbX1jZ3WgWpzpPYOY3VXlj
dCpb+zNn2QqjOp1BwOft0OrBgH8UMvTrcU8wjwAMubSml6WUL2AvmAnEz76ltdX/
cOc4LNEg66lqjSw1uOHCU3k/YU/uNfB6QcBrpTmCqiZGxsmo8H9HhLoUzpmK9xgg
r8cRuFt+rFS4iSl/L3Xtif4gpmpo9au9dSPMKHpiGXpGZhFBoHtZHUTx0FlaSPn6
m3DlNvo7AK47lTYyZP5nUwnyvcIi784LUVT2kShkZJHZ89NOzQYlHNR4UuFafTm5
nGo6n8hf6fh/MAw1W9UiyIettHJ3ZiLIYu+DNxKD5t/utg415O21GcG4KrduMP1U
PhsIl5fDj6dWOEUMNET4PaPtFfIbXuBeZegi16Gz7/105rNt1N8Pksko25L+tG2J
JqbJrZivjHoubIwgcNq31Pkw3/rY4fsk/8SjdhTq3oHxRHZlG3tygbeuvyuXq/EG
LFbMJ7y7LvoP1Hq89jyOAskXiTuxjNwflmpsWgTP9/53amAZ/1E01zco5KaES2jO
aKrCCQRIph/ltzfXbfbwnNwC2chSsS33HWMahngSDV3mALB8npUB5msFHZkI0H+d
mEXc9udfWgjyXTW4KC1Gc6MWq1BPVw9fLrY3AJgmakLjeEXbsMe2DdkqM4T/MkpU
A4bC+X2PUdG4gMMFXrehDV+1o07S0h0MVpZSkZFxdx4IvEVIhkl5OObv8SpfOYeE
RP+0jJw6b0SDqTW+qOMIXAoEDVo8kJddnBgYu9DYEz5ak9Zpaf8Sa2RI3psMQUk2
pb3KHXYpXHf4Bth49c1DvlIE7vjR4btEjYtJ32Mh6A35Ch0h5h/uTleG+ocrbhJ5
HN1sYgwPo4iHb9Fd/KJmTJSoIfMQRVKvs3ajXI6pAUvyIAXvAUJ+IK7Pqy2MN4RV
lsps4XZ2oqQUPAhRHNU5nyyC4aqeDncMEM4rqaZN6N+DcGfPvhVRUQ197WpgJv+C
hnAe2lhZ8yBJfwSGcg7tGPowO/ZNX2RT8JgyX0W5/KdFj9Yty75rvF6xfBxSYvFa
3ziltFsXxUls3dcVeKkzeyo0JO6bTuS2JtVc50pv73RiBxN1YLJg0poqyhJ8QSrx
MMtTXqWjXlsyiPlUcsGM4ReONCcLLUJy+vR8iQY18ED/ADlycraNHItVERvXxHc4
iEWRHhy/qT8qjs+SoCnybr5BNWdcWM/Tj+EzTelMVJmSd0gSDfE9kXu8BWrs7v0X
cVPLmvVR/Jh8u2qFCpAcBnfnZGjapLFU4pT7QRdrdP96iPYQFkV9u1gmuTsVbFNu
qNCkypEYUoWE04cPNBTPtjqdKq593DH4qr8DeenLKCr/7od/jHWwG6ET5hQ/FHJ8
70QYZ6qMn9ZOwJS0Jn8+HvcCIudHXQf4a8XzW7eC/VPZpekCqxC8RHNj5GkQDQMD
k4hM3jK+CMBDLd2n+s7rZpcscSFRUoMvS0mVUPUUDEhlC0GUOamBTrMScErjsK3z
pg5OqxdUYpCcR8fdq8CdYWuCmwK5v/jfF+dxkHwWIY7TX4OwOxhrCh/UeeeRObQF
xNLuozFX2xw7fKtzGDdsmxH/OuNpZSiKD+blITMaDHCxxz3/ob9JZfJqYn+aCd4Q
rSO/5VwgrmpJEbfE7wqnjY8WCjeKTi69YQ73O7yGWAXr/kyM38vLixKsFNAFS0wy
0aS2Ra0Zn2jPwMz1+0pqKZ5cI8wpnvQKpSXnFLph3xtoWO9QidbQ7DaImxyltfF/
W58kwAA+zIOoHDZYK513o9dkicK2wpF1OlUGaymDh3qX0xHKvv4dP0L9PcT1dmn9
q5riZFNXjRcReNQ3l499LfZg36oi7lUcqZwi7SsJ1tm3z3vO3fuRPm4fk2ydCAEZ
c0phhnMaiYcmAeXulO9DZh1PMZ6YMZkgPxadtokDN3jbkhvcgt56d72GmwZMUd5W
FrrNyGVE9siu76ILrBE2IIx0mhzyuaQycmBF+J02PQm3g2x0b05WAAP/qJigdS+l
jcpsj7Ux6iV5b+T8HSOkzuBD1zffcESwkJgIp0q2lcc+DKBVZl0sWpjvs0FmvTuF
0gkos2FgNMU0IuxC+vrTPhI2u+CbN8M4zKSteptxN0bpIQZmUduEyJ/erR3nWMrP
C8lDFEw9z63FsyLDZCdCYf2ubiJXRuJF74DaazwCmkJiMVW3Qu0DF8cMdOupKrMT
Cm4vT3KHYR6nHiGioNASkhqWqaYHYnKTGWxmNNKa/7Qnv98VAHsvmqk3UujhBgyE
YF6NvxVKIJgS+AnZLHXk9/nWQ5Q7XTBe+Rcxy/OEKXikeUH60sr3Fiuhr9ZTTtcX
HER7vKrnRa8e59163/EitAa4fshPVO3GD7xWL8GSQYsY8QfU8gu6xto6KPIxIiz2
mcXDerEZ9pZUiQzN2ZN7VGK/vEN0a27tYnPBorMN6g6PFgdhSWhTaTOOt4UEhWFf
OpPAO8hPRAdCtxL4zOlulPF+7H3Cb3DxDBMoyw6t9y8NHKO2VPf4GWhxSH0eyxI1
sg68MBXCjq1wIOVdKkgtOPTtmZB/LLBWbhhL8nJ/9NeINEMpkpt011aujdPxgzgI
ML9zOSaN/qrubktwoBGq8jmA27bO7jRJuy/1oBYO10LgBsNhj7C25ULaiq363t21
v40wXlgCX7l12OufET8Je1UFPa3BP3EszRKhimMZY6PeTNLZaff84gA8z4Utlbzl
IHlkkKfCxfa0nzaiT6sNHALfFsjfdWOzvSUDwormGtyWZ2cuEgUOCBA8qWtA6w65
C2t8KtEoNW1ZSIie3YvFrntPoW1LOamZ0jwWWD+uFGgojxbrvrkw5kzpOJmHEI1y
s69ntvN+aL3STFWe1YwcCO1Lr5vCzlc+5M0GWeH898/393Bnd/rG6ErhMB7wWy4a
/5AOYmv1aKKOqNFlwjmLseEW8Nz7TR8Sa+WN9+0aX6zBSoA4IBZ/PKgPlzJOmcdl
Ql39SL9xOHWKsW1X+JEC7H71QJ2uXxPyxKLTFmw0K7RQdDbjNSf3G+jhwJwFhxg7
zSK38AxLMuyl715qs5WZbnjtBb0DkZDS7w6Ly5QlZbuNv3HJzMKnupQOhigZmlq2
W+SKfBQIJK67/J1o/dJBLe1KcR7xrveELQp1nl6ipe9ZBPjshBfWzzabKP1fC/p6
twNEmvqxONFWXUzbmiFweRRY0WvsZ7x9HmK2J8Vq7XZ4AAhFjm3Qzd3SxyJY6Ha3
CFCOTh8zeF9NhzsLCCjuxIL+N5YcKTa1giYXEEuHk091cCDF6ViTYSjNgaRnNHum
ibbopcqBn+mOF8ZBr9z+jkXaCwYh3owGxDCSmeu9TLGIg2nA88/WvDk5/NrtGVdN
YzwJZM/LRHg6dXHMVNjpnxs4K/F503cLBEOJZm2wDtvvFUK6rhoYzSYPuF+EV9Zz
pxO8bFCHoCyEQbteTG5jR0iD2x5gjdRCyu2xryGodgNEasFSo5lUa1mnT7ltq27S
L6ZF19lz4yZqFlxiDoyHfUKNAewuj/f3e/EWCQbo4ppFCqUAi0B+/Pb5Whpp7U4l
rBAmTidP3cCbIt0M22QLStQXMKcR44nw0FJS4FKRIqeWPGxfJNDeSORsjCBLJrrL
5e+p5FJgM0K3DosGhd41XOIild1ALXfD2m2RwJn+t35bsI1UedMIuvGcToOPMimX
dcS++crV37mzzYYaTcNzPLoV5Arw2qt7UE9cunoN2Js+dbXzc2icVPpFEgjLxBeB
4vPfV4dEizt3Dv7PRh0uCrY7gQYr+bj16iX+/ayabEHjNAwH6Cw6Sg9RSVcs8FGi
STuIZoeNtIMFoR6NFI7gBApnOoPoKtUsd+ncS7+lZNYtuPn+E7Vpfm7/nBToed3H
VaVE6/jP92XQdFojK6YKBN02D3WkIWAvIu6iDWdF0X+4CxSuePx8VUJB2R6czdBO
/Df1R1Slu+7NENtiCl/FiW8PNU1rJV/TtMw2u+Aw3+nUIRuevOEQ+Y+BzHhvIH8E
af15Ssgt+MJUDf+vOWp49k37X0izhM0X1DIN6c39HOxDqI2mz/Y8s/jj4TPgNVtq
6MvQqMCbaQRYtIEtkr/HFlC6WOy/m1JfdlY3rqgJ9HSmNd7cZQD8UBMq76QcNZPY
LyxeHW3MzUITobSrKsBicnTn2ioxhk/PwXsbKtEOPMAugcgoJoJNbN6yuvWbUmcL
NSJhfPHRtXQtSYNwNrPxnhTbtP9ZMWNHdiaKYS/Sqm5K8foiEJpYaWQOP+tFT6i6
Ofr3MSM+YxwkMiUMYPKKoh9Wcit4K6KDcl7gTQXqQ19iKXXqz5IHuY1aWDAfteLX
OhD9ebvdjvEEhd7PCdfMqawQcLDWab/sbxdHsq6ldiH9xsYuwXSAFEm+BGFIUDUu
aNk9epNqeTQjLhq/4FsOgBJd/Qx/BSL5c7BYX7IHgIZmAbOXg7NGtYlxrJFSKdIs
uTOTvy+rJQaJbzmwPyUzSaetnTtBV6FMQsb77IijLFaZu4yZTiY+ilm4bCMVz9Yw
WN+r4qaSR8efrDrk/lWN90ZaLfbWgweboDuMe5NlDfXnQhmSxKMG7D0sIgJWSLzR
cL64U5JpDbPir5rMzykW1GxrlV42/qBGtK0V3uALmuKjfZVGbaKt8FT6xZO+P7YQ
4x5xprrZMBuzun5iDC13gQsHHuFQDHjmAOJXkSktTgisoeUDaWtd8YV0Bd6LN8xw
E2Fb7sXwMI8G99AFzOsqq1YmwuZFku92ovqD8JDfjnJqhYitLx6fxGoKSg7yp09A
ZGUFzThsAROpqptdEQJACjyzCJVAUNkOhEzl0+Jh6tFwa6ADoPGM4kGE2G986JQT
geKE94tA7SZHJ9XkX7tdKdpKbilJWc75E9zGLjKaFlkPU76GMPgKtVVRVtZNCVgy
zQeJFf+EZI9QBJNoEnfBFCmLyDEQAoRO5AaIo5bM2wRsuTX+GrobGWn5pOOuxLlc
cAWp5CVNJK595D1Z1D3m8HWHipmFT7BUwVDgoMmZIj8N8LoVaW7e2vFwI1Tbv2Xy
Oll+Tzrdce2ooIJRp/iT5TVFoaNoQQmBWkCitUDolBE4wT6ixoO+Oe+R0Myb+1ih
NxEbL5bvNDTeXvVfzNeIdIAmDyxJXIkaoOS8aIC8INlzi5DTVd9LWv719NdSpVkr
TVdtJvh20kmVEf6SB/zuphlA4yJKxyZ8vJRJ8Jlw90kjIQPVAPE3HM23qxf9h3IR
JIQGuBtecndtDqrX49ErkL+2hv9mYZ/2nNLsU4L91xB7pjTgoWNRyPyrnXPbzBUw
xyfyP0mioH9Frdowem/1RWuBjfA0p2gBUVI8M2C7pHxumi797t2OTUWSFvY0yo67
O2BR2DDLFJ26/hHwPe3jUXbkFi/4ggyhYpQyBtG3eH0cJzP0kGjQGDAZaKe6SeWe
QwwzW39D2BiIA3l+MFoGCEnBbm52AnCc1D5TFTIJ1eqsnfCEe2m7ePZbQobfjCXE
jInZfivqyAQwhXaLNyqmNJmFwGBw+/okMyvuG3PxdiQ2Eb3rXYGvLszq5EiMBUjl
JxqnTkrIoe8GWtMIKcUHVlHsIlueYOcnpnioB5Fv/R2hSJrREf21woxjDSPGx9jA
FIRCEyFZTrXOzNxalzspcLJ3DPLamD7UrX1OTHauiyaY1q+J8eHQwWAXnLOLD/Py
dyfcWn2kA8y+V4jzj/d5j9zqV37BZkfBKwP9a17cH8QfwFZ+u+tNljuX8gSrO5GR
eVfcBV5KfKqQ81C27nW1NUzY2YLBvCx7o5K60krAeRUu+tK5YvtILchvRViYdkBW
8CE4fqgnMqJ6cJCpDNJXQzshTdBFBQcdJ+UXZeJeQj7UauHDyFQR0+W74O4Cslaw
Cd/s4CKhUd8OR7HRwYbUDb/ExhyaGgZ6mqWdVL5A7xq4gY+5EKNMVSgrJIu2iAw1
uzeCP5lPpnBjExtSf2C/OQnWPCt5Wypzg3moXGkLKE69QLLWXUgyK0AwC8NWVFCJ
yJXlR73NnG8d9vEtK2rLbWZxXKXJs0dGyUZ5WJgfapHGhJvmHdSd650Zdm4UrGHA
mkK6fBDBmmTcVPJIX8AvqZZjtw9fTILzI0gq2Oy5II6NqzfG7I47m5zRW0VJJ/c3
eH4LF0gefmaHpthtLCRXXZyj7+Gqfhbu5snBGV9ZypbUGgQkef2G3QL3CgCC/Ubs
KRZsxAQ4XuxMSqFw7daP8WxNWfFgsf3IOUOmiFm/ljOolO/UW6nz5nMwvOVdS5hg
x1qURxfJartI8ewVtaEPpiMG/1UKwOuFGZiDMO0Yio+8dz/1uuVs99CQhm/lEkjZ
gJ0SR8z7Xidy6dAMoMbb5VYx5enQNSrqa1iY+JG7NjBOlhj4Wp6UpPpfHZsh72lJ
Ohb/mxOJWuIAF208IjqJPC1gIlNboY5kCn8tIWdt/dMb2btHlabY3JdCShRUTH5x
pUUhG1bQL3M71R2MYbQl+RegNcztCN07T6338VsySVw2qYbJnuWsqJruVb/dBqv8
2jU0ADqV+OwveKBBgiwS5xsu65kQA5SFsjLCc+s+RV3rVG6qrLxOypMI7JXEDD9w
Ui8DgE2IWUG8SqyOmWxHdaqSDYCtySD0qegBIKatOvRschQKkR2dmPG/6EmP/AvR
HAlhfAc3h/dwG3Cn6tFIoHc0tnQW06o99WUmcff2jQ6ld5XkvEmRGB+vg85l/WKI
6PFTuen2lkrLZHjUTi2N5kGWO+S7CmWTbZMLxAtOX9jiS5wpPZSeVcNVpoj6k9G2
SP/4rd3F6aDjkoA6GgpUdYJnwlZU3cvOrW4w55mOq1r2LfHSLSPIgVBs5SQ0SFZy
YFXWVn6UcrrKs+iFTZhg07uIZAS5FtBfu1HA5mdeh3gPBTxa9agGPixhCnSTLYGW
rLgZBSwdT78RYbePbj4gi+MqI2euVQtcC/X78xLDFk8HD9Bk/dHFifQcBRVUSQ+J
CSIYp1WpDcFKrYMX+TrSWs7/UjekPVALC5nBEsJkHe5EF9OkdR22eRs/3SItih/H
cRHkUcZH22eGHcv+GOCmJS0g2Da51SR7Cfb/Y1zRuLVHKRHSNEuiBK5sCbnA3jr5
hhc5e+Bc49G/PdO++Q9poC5AN9L8UicBwVoW2WSoh8yg6L81RIVvZ1v0N2dkNtXX
cCYNFArd4aPibHbM+qs0SAqdu1l47YSA2w1c+yp7JeBBoM5GuwsXsNNQt7/cn7xe
Yoz9QOUtTh1SGWnjnJ9UBpI8zX8k1PKyrfLZSF+rRzq1EXgjt+6fNJKTyEZMNhWd
LLBYLLaocD0g5C5k+Vu81CjRGNgJ5oYkcMznjANvhPdZIehLdlHDUrG4BQSWUJHq
Yzf6YtjGcjt4mbsp+0q6A1j++ARxVr6oT6lx9oaCZRFiThSnBid1f0oxSjid49ro
TaS+ewrUJ4R+TB3Cyo0g0+/fY4875sGg1CwWPRHSxRi4HwC5UWpUxjl9nZn+gVgG
8Ej8LyWbQ0B6B8iU6ST4MSBww+tBiGRviX3AHeQXU/XsbDNkSbWHojgUgpvPwFtY
vjiwmhsmjcJLe1xt+gUGH7wpgFhzAUPFlyGXqXxI8bL8njcr2LPBfd8B0BzDf83U
p53FNtvsSaX9227po66Tzv/Zox/O40YgnzBaB6rIaQyZfZ1ccxmbz2RxYP6s3Z4D
k/X/spdOhgrI+UV+JNp4FF0UohNm1hl7pb5dsEhs+rzbGPEnuT5tKiffPV2zvZ75
SS31bEtRHzjb3bS1gkKKyjCL+FNuPQwwTmbSYUldsUkdh9e2EIN25fXxy/7IT/5j
O7rwBlOzLv1VE149KZ77g7tpY3oeuAdhYD92w6WGCkF9ANIIjyoWSsUkKFnFj31r
ayS+mLVcAA+XVupeWPONoaxG0wyEwvfq9BMWbphNLQcYyXAVN4lncHTHOCDt8EXw
K1p0MXvf5upjnQQMNA/8o9rwhph/5aQTZtFbcyXIcTffNxUg3ixvtAZrID25dwxV
nsdK2b98I10iVdqvUxvbk8ebzd5UxrogVPgGlG9JtmZONu2/e4g5dUA1mWlQpIdz
vGgoNm82G0oO1XauFm14YKAIyIEnA2vdq9kzechDgGxj3QmfYcyZV9RF8GMBV7+P
lhZkddl6SvUAcHSug9AJj7DaqircTdekHn/+7vjR/l/F7JUX4dmtfGJ/uTo12uI4
Znu2HlX2yCKorb4oUlLiWHb9PXOzmSGeoNmw5ibUvI1n84Gv75ki+VHSNY5+D9mn
N6ZMg0xatMYrmmFgG5q9PAOx/a4+75z+DQBQu8sfUZW2uEhU6Epywl/cvY/F0bRT
ufB1aRJK7fdDTUOGO+SYTTHdAWOSj7AEqfygMKLdoVTAWHhORoIa0eSydzeFnZzP
cvJ7Y2wHUNpg6sDZnXdnjjzVfJ+HQx8WdL4zvQhMxpPKOMuhKBM96nAfq6yXd4fl
WfcgpKHRbXY5ne9RU9DZ2AnNJp9jeeQfspVl5qSpCIv0dKl3QdWhSwbBsoVDs0eH
6wlt5/N8KDdZTADRSmrK+LY4B526jufue4Brs0N5YgikhKQDpsaIBmc6IBkkfDNH
gxI2aMGiRTRh5ZDDfZTZAC+6tHCjJDI3dE246qfnh2tDFD/pwhc7oHhCbc2bxwtA
rPvjx7t68shelh8AzjC1wmvobzz6qKgFik6ZNj0YmU4QtdG1Y9dbAF9Tw436rowu
phsuGHhGxP4XspSymICrd+eWPpzBwVpfC++QHkXn6CB+RbZskK1LYVzJlmdksfrt
/hg+H3lUcGIpz+dYCdpV6q2UKghPdaJq6Nt5Cq32JzV7Ie0vvlachUd8BByCfQh0
0fo5SIAeNEX+YOhBscKtIOpOsdbYGgV1RsjWe29TaiciXBBUtAaX44xxNLpg5i+3
QFcwNMDgadTJN0Zs3a2lARilMDHgiN2C5LsiZkwk1iXg3x91oj8c7ctfr15GkmgC
mi+CY/qL9tIT75TirLUEgFZo3ykFBYSNwk6waCw/UVUMNqog9fc5B/B455j6+fGN
y0pjwZ1rqvVwQj3nIgQB3ABd+JtOZgMXw6/3buGekMsIdC5EcSdY8JOeXOdZwMTG
qeHXWCFF325ivqzzOwRXUeLVbtLOTZBwC28VmC6080soPAQLijFMDPZuN9j4f00r
6XHnTeHxw+Nbe66D8RkW6AKtnFtoxj3MOakKnPIKNv8loMCrOovxJO0YwLnGBF5t
rvLVD7gW3yIx4mAH6DcUFu7++9qfvvBjYog0TMUY+bQ2nn1puvLZ4PM/KdZkZZ/b
qppwNSzPF2OA8TaMHrI64jPXkWXPUZObkjPRrAs+BvTJ51UahAMrM65NTAge1BVb
aIR4vblixwyRi892SHZuBkDudVcFYbjJur5f03TCfTDsNnp+2VZjO3ZHjNaVx2VA
UvextvQT7SQG1gl6Amwx4YtFi9Ju+hy2RvDgjiBNQHYD2PPe86cHTNFApvwp5owp
Nq/fV6wXh13N5XGz5EL1wY6VjHluj6uZYUpVhMD9en/FwSCABPWhKSkNpqhO+bbh
FxkfbdUTa2Yb1YyfwJN3gh2qRpGyzZPJphD4RlxqVL7DFuvLh3Zoagkl5hkSSpYj
MsYXbtuBvIzHstPSHC1mge3qZluk13rFLKkoQU4Cw9pGybkfIrZC52WWevblrXPl
u8k6QobPz7Lo1mQRVCOPu8jntFtVqaqKVCRPszUGLPMtl6lhED+F688CS65cTALw
6zcs4e3lcHY78VAMvkmsNs6sPNx8DxrfXe3v7XnWqi+ngrSFRIFfjJzwKiqF+9im
/CIsdxEIE+9JwBB2tQCFmqFNroug3kNdjWv5iKy9ewAWTHmPUnksI/9L4rFpqWq9
SBkd4a/n451trD/DumMz1bPfywXXbt1dnSSbqrCENw9ef8rKqJQ+W8mgI8HSHSNU
XLpbps4VUjo/YAc3Mrn4tkrBlEFNy9N/6IT6qtAgEVNhPVCjVZGCRcZA5Pb1hnDH
M/4HQTRWkSdP/V/C2THa1GK0SUX6JTaDm4QCOWH3P/wa1EAaXPKYUqz73qA4vZfC
O4mqEnCVixbi68cw9F19ctXRyidTtBU+EgunMTD4X96D+gEwPGAAeueAAjzjAp84
hrMQz3QYiLIhKa9fT/GS+CEwSTbOSv3Vhl7wCoTBRTGEO+M/aIN40b+Iy8TfOICG
np2NCyOZ963WI1QbquU9xPuGHWZjQQDFVSVj3YdXlikF3tLXQM9DfjAt61tL4GoA
5c9yO11W7Z2nL/g1jo7CElxo+HN8XBtmRah234jBjoa3wVaBDYo0MOPEhdkEEBKL
toPJOqDEGxKQzM9vNjbK26WRLkcQ1qr5kS4xqxKOz2l5+DEq08xqO3V7IzjUTvYg
Gi907KAWz6c0oJBzJ6S1l4RhgYxt4GVP7RVxHhr4DxyLMD1HLSK2bzrxfdss/4SW
U3aQ+nNmC4EXG4Ovv8aTWwnD7ywBy4xmJhpBLBIRV3zV2PfHPcyr8y2wyKC6rCNm
7w7iSXiDc4IeN15lSF4VVsGVWoJdEc1FZXE3wkLGCyaqO7HZ3bTNP0jidOM5Koo9
ZkhySslWTT1XWvZnF8znl8hftc+SXZB5ewvTAhKWqRbdIgbK45ULnB9T3bsZqA71
vSXoXxTdnBhpv3b22B/9hmzfLek5+LptAWrIwLUV2UuJ9dSvwFPRMXnPxhdqOG9j
iAzN+gvTucB6rQGawA3Gja4As9cSjQOwZi6E+3V5fW2RNBgnQrBPoqpYk2wc2Bih
AodtvfJ8a5q5LDIUp1kAZ/MZRdU24/G3E98PfmTE7E5tl0QBpYEGYIsrDK2263kA
CCto3RswQ/Q/VY8P2R0TCSXfF3bnt2cfBvaJX+hZ0XLzXdc2j6sQ6VxA+lkVj7eo
hL8hO1BlcyvQwiKGXI5ntnlrWGS4hArGuEdzgaLTVxGjMOcsXKyrDd0cOPjzpx6n
+j+FLj1KDhS2XPqc7m45JUZk9rLAn5jmGg4lGo2ODYkPyAN3nNqGTldeNqybUUfa
ub1I2UhqvFJ28HJxdFJI+kDK4geSGo0VRZ/uGsYGJjspCB/R6NN1g85S8ttBHuWw
QMswRyVUfbkQJ3nrV256GEEajk0FTUXWEMACOzf8ij6IDrYdmE/waOAuj7dGQnFj
3m/VxatQHVnbqfe4HDqICn0ObFNmWj1dtI6tM8UEiuWVoVHhTfne9VU7styNkxte
APEiMM7irjD/0P5Aj/8V7DTp/DB94C1skzrrarUxy3G1r4NuLB9hEkRXukh/EB8p
VbOmtRD/rOeoBySrfTaF4qLncg7nkFy27zPgzLmCE8zOsuo9nENVk8RCosGzEcKR
nbemDiAFm6JdSTPLrN61ekTtfpQSMyZBkZxWECCreLLmymyKYv974bJYnY6bD3Bb
4N5z6h/paCuxRqLRpmx9k+cWFpXF/Q/3JLWKdm7VhoNlJbKhiq18xCY6vm61BKRC
288ApaYocYT2UzHuwYAsgyPMwnS62QEtbBG47jZ8CCo4H1UtP8ldqjnQEhGCtBga
Dz+5/wu3g8qAgj4MBqPpJuXxLbRPCjIFU4VCx79xtk+KQJHDb+niGlTZJ/hgDfaU
ItOIU6RctmoJl4VKl1F+RW+lMFaETX0TYCXY3lr42TfP2g1AwtkjDBnRrGwNg/2X
2ltB4UAB7C7lvntXL0Yi2z3SwLj4BQnVTcRkoUzwP8MedFFVLL8mGxws70urWkWq
e5v2wgna8YRA+022vjVy5VGxu2yskWY1rul5ph3czUtsRfUBOOi23oOvLWIWkhqk
GhvhxaTWIAqRxCxF4DKV2zHLnBWHmb+myPv2h7qBBHwHY+5SXjj9ChvE5ASJ6Il8
q3TWo014ZdWEXm5LzLUqVQ16ZpjEVqXfqru7rsqdNVfkVsEnV/MdUO5P9hjqCLL3
fZcWPELwiwcgxLJw/TVqCb6CxMaRY197EuqHNE6wL4adup75MgIarcGae1ozSuxO
YDBp0OmfXCQzGVDeZxG+jG7qVsRykqZCo4D+p2GjZDPTkvUscYPNjTK90uI5FUgN
p54Hr79ZEDOtapiiSV+opafCKHEsUj6OXun1E3/I02/lzaR4D0oENeuZ+jRoYcCs
l8xYPzY8RN6NPcXGn4XAKjJYftpdhA0888teedD8BbEcwaQfOS49gh8EJmIgdaVb
k22/6DZ1yyaR3sVdzUiS23e58PC4NnQw9ZHzCrHMDDv/NtxbzpJLSVK9qjgg8nlH
7OfhkRqhFhIzHE0X1dnFBQXqtOraRzbyasLus52SEjalvW763ZS4efx2FLTm8eoT
cycgT7Kz2Hk6x65M+6W7NGm1w7vKvKNK4c5n9sYae33qwhnc2sxsvAgfYhDtt+PF
fIdB0sWd2461JriaN8n6U9dclArhhhUlTtqxYL4Zp3QbRO5kBpDcWZnf0GNcbyUN
mpL/QVvvvEmoaCL6SsVJTkwnUisXbzcRAybZVryGxNLKn5n0Mv46Y9bFF9BJ78dN
Fg9ULIS5Wz/7OQ5ne/+bkTWoOuKGzGQk5/TkjI5z6R6L2fh2qMptuxcO7RvNMZ8y
hfw4vToiB3EBa0csZOk+LQhZCaJkahkSOXG2cW+z44KKW/wsWeg3GYfACHmh+TQp
k5H27NmsXFNm/xj8o8ieCzFalDuP+rGMuF5Lh6rhvJqwODwbrbmBGR2/t/7bahiQ
owyzSJmLACUjPwjBF1+QJt61dTd6OYxENbpOqv0Y+cJW80edbxm1/I/ProuWyVYb
XtBTU+l/nYHbdNhWX9CKNuDt0pFDNB5VN2M8GO/oJUPL+BlYTaCHXuSdt2iaQLzh
EWWV92y/27k92JjQ/R75L9gE9GhwA825qjT0uGSUVQy2fAiWsaL3SgZcO3XX8n7h
1l/ozfblabIdEGm6VEjh5VLRe57FYXlMFosnkEHZHmOSTCzkDswRyI4nlXj1ydRW
7Npi3P4CR6kdAENLzkVJp/ONnZc/3vt+92IeMP2AqWaA1KFOA55KcOuA53VWquzY
KMQCqVF3mrldnZ7e2LoaP/6uUoUax+rU90Lr51rJl+6fCsEn+yy/kZNj7zlmgnaR
FuQ06VBuEpguSdCxjrYL2X73OW6SveQCb5Uc2/o8sZk/gjFj+70eHWd96/D33wzA
FkgzGx217tUJr8nqLL0WseQktj4cKJ6SQejLQQUxvtn35neTn9CBypYwUfNR8rhH
wozwtM3+g6o7/1iJ4aZPn7FuY6qtmVoFX9hn0gePZE68OUw3yI5iafDxgR9hh7/L
eSUK0LUAK5GrrVQz/y9so9NI9v63P/mlO8+LThZGaqANcPPtThbp2rZcnCqYEPR5
ttE8/p9/DCLUVzaEZTNkhofPF1W7UkQZBgEySTsib3X26cGhhH3WuRkw9BkewGsc
ybEVPDoOGIF84IjBKQK1WAhZUzCUfx6BSxwJH2iUyLUUFKqihpRzNxXJ+4Z/FpsO
AFpRwkF4QKsqgDIormFSDijS/ZKIxCpIsUyBYmzde9PEtnTX388TwQfSbcFTu7ua
jXQCo3PcCSnJA3TeRvCarcUrO6VL3PpUYbHMG8GSByDht7/LMwv0DrFnNAiFEYNk
UaI6Ae1WkmobhtJpSvcjzUYSlXsA/Q2VWNCLP3gqcnmqX4T+THNCj7GfoZL+LWVo
Zy1wfVoAYD1m7nfIHDeDgLXqlgCGoJJF2TNeN/tDkcbP1wCUwYlIcO1iVgYLH+Bq
h1DjaTznoKvHdOYIkqJXEmyWRh1CKmsU85UIRZJ/B29SBVp/6tHYgcFvu/HsLPm9
jS75t4LR5tgqGiC85v2Zo6rbjaW1Y8iu86Hdjcp+WQkNqOB2vzGyVNRaiWfNrdhN
zaVSs+P7D1Kk1SdW9933hTYX7xHsqip0ytGaTA0kZzSnWTwKYnT2nz3HuvizfPtz
enMFV9zWpqztdecwQlzkBWwdi/eTJaV4UQksL71wvufDVDfDrSKtwXAHmfwR+Ary
5zqJZ+8BLSME2BhoP/u0DNyM67xd2/AnOFo0izoEwH3++c0Nnub3v9pdU6lBTyvy
n3IBxLKeXuZCDrB5vI+YCDXyeaRv9vByn25irij+4KasvNrk2A2qrF8K16mPVWa+
Qjop7xNRxuACqCdnYfeGfe3YuxOm+zunHWtdbKfRX1AXYUmsSW1sc+/IBoY5uSaG
FP3bRUWd4z/PzvX8Es9fCKQgVSXIUjVz2T1T+o3peTHaYz6YWpBGtN5iOyhxFxmA
Ipp79n9uUANE52+KltYU5rHbKqp9nK9sbiy90PTC3ILAkgirxwELbT96J4UnAO3o
w/xmUNum850QXC/9FOv4fW+8GaFi7rbP18ST2GiFc7/GXDC2P3Yu2l3y8Cm+Zroz
S2+LKp4VCE6Jrt4nEMeM8kFjI5gRXbwCa0m6Mf1td02jJeWhSsKyyd5Jt5w0F7WN
ME9UVtewIkMUz0NHIN+XTFfoRTrG8WR810YZAp208u/vuRm77ee89OrI3e3HzZrC
/lsTi2pwo4QQuctdPr+69JVsb9RXzHP5kkK6HsbBN2j3TznBbHNax5hRXXayComI
0hx9fFHGctb2WjQy6lvzNgYzVrEq8ancKYWARVuh6SRZ9mpFSc8Ll5UF09nenE/D
j0YfA1sWkcfK5PjKTy7NF5ZaTs+i0FEK/uXsFN5L+VNikDzeBbgKX4ZhrZ9WRgp5
ldjzBBOGz/Ug76e7RIVaaj7O1zOGVnLCr9KlK+HwwyPRDmtmBT3AqCS4m/Zvdjq+
tVJbca7PiCF+j6OZg9daH87BcVJ6k5g704YkEcHk2g+w1xLBcE2Hpo5ZMLyCZE5C
Rb08H8/oPzfLFmeaYH8EJNI9G/YT74oLuww5A3xxv4P/Byv0JKZ9yg2vKtZc3M9q
Z6eR/YnmGULcXSUd738EHpfDUW2Q3RqnZSxN8Q4nSU9Pmnqfp6ykmVuTi4LY5Nih
34LoGHY/1P3x+zTQ6fNwG6NqLbJqSqSdWTv9a2roBj0SElNNEwvkhkCJfiIOOFFm
t2y//LX0GYR97UJJEl7QFAAf45jmEFxAfB0J3tF1Kgi2NTHnde+sSxcV+vwoIs8N
ZlujlLQIeoUSHWxnPGXZJyVoGbKx3D1c2USc+Zo+wGKa3IxFCjDPWp3/rybENN7w
a3grmP9ll5Ta3KEbKJbJC5l747aejP1snL+633PifKoPZtz5TryW973/MkATJDb6
IRFKzBCwbPmaO2kqkQ3LS6l1yGNSB3ojQCb34cTrFd1PeLQTTlJRqocp1/X/V5PJ
rtoQvYEnHPYo7J/PjtAJIdnpcs+FMKpNz7J2vdHCtf9KjS/6Drc4MYbiGePnIRry
bmqbAU+x8RiJE1nXtYlLO4V/GoJKo2TjHxF287KPNeTQS++k/MtLdeLBJb25UwpB
EAhQVtRXk4+YDOC3N51lWLlI1l/XxC4A3BjLSvDq0WXXgJkieqKbpw7k8gs4iwsV
JEIIHl9+9z2v3gnwGOEvS0TjsPUqT5tRuKeOGiCQ8wD0WCqLcqEF0Iml3nvukS9a
4KNn31Bs768iTMWIP+h5Bwj2YAmE71m4P2hU/SyA14BUOfYhYBFpnLB3b0UYd90U
IrUWHmcl3EFlFvD7FMCE0GmuAGbVLLpzB6Kkjbea3WGlx9MkHuXFoRXEVan2F7Cb
veLiVzMsB4diFSGRTjGXubJx79icaCWlD0Y1QEUTjNMcQZ65guVHsbLFJj2Vun5i
at60VJ722tzR+F1nH6sMmmMGHW3MD1DUXnkRIF/j/Pkpr2PAVKnLQoMBMNmG2vQb
QV2Qmkjc0D6B+50i4fZecPSA4u4sq2jiDAgHx/2QJvLPl8EJv4FZHlOw44onsEri
PAdTON2ggkltVq7dGHi/o5N38xGt7ueJHoY+ZXnAXD15pBzqw1wxwKm0XtWapKU6
YgcIHMTxcEYRZ6+j85O1emY4kvXQDxFC3qJ5dNcVp01ZsP7UV/U59x7LWnx0IFfL
CSqUljzDrkgfv8JBW565hZvquojkRI54i/JK1bO/pUFrG95QIDZKCSqQUMs+xj/C
pG6/7RSDCR5CK88K/F+7M04qKoQrMdoFmF+bMRwaOEZQqwNbNkR7Z3awoYBhI9Or
r8OqGcB5PlSLbUMwfqSGV6VOMpiL5zdEzKqBo7hnkVPelHcA4uR+gRKjIufNs573
FJXXeCY2QxsImpo4sTE1Uw8pog1QL8Kf3ZjdHl4a9RwK0QZ0XQgALx806ogL3gCS
e4x/JJfalare8Q4DI/L7l47LJgK1vKk4q33Fb3u8XJvkFwNJRcowk8g7YbQ2EEkL
5VFoCz2khR9SE2+bcUONH5Hggx3TGc8uOFtGaL+p5vXLPudRvhPu8C+la+rY1+r6
fFMceWqPBsms3uQ+3TRE6SlRJcg+2XwsE7JMroJZRueh/1zQwkmPlcA+xbLcg9J+
9OovdQGgc2DoRTqGRD3MxPa2z7RUgTd702DdOoollRrYckeCmlbNFXr+L7MDuvh3
hDwVRahShbSMkkOqq81Zfy8YQ3+wPDgG3fsliXPdnKybyLVkAkd5yEiRhE2oMTzV
3zDgSgEFJ6YcTZBGRI9vQdFouRvgFmtiL2jHorkI0d/scWG+Lnk9OmWIoL9QS/fY
HkpF45BPHdMSbBLl+XgFR1VlU6+eI1jEHIhsE74awx4Q69LTI27hbFF2qOWB29WW
USeTNsu9DeapOoNWLGGUj85WmHEwfV/UBTE57iVkatBU1JoWO2xWdVng0Q8/z5o3
Hc2m0NNUYTzVRevuj1o+3b+by8M0/dxyint6nqMWRbFofc67PUFGqCTu4UJNyxqL
bT19391i7jx3eVdDCFn8VDYGklNCxACIMWSHJgKonJx27NU3roWi0zk5zXyBuHVb
fV0UMEg8ZJx7W+d6AjmH6Mtq9PHCQOc/EVXahzxlpCxexoJRs4Bv9yysLCxJnmys
ZtSti1MHuSSKebijqqLg27DsVUPBG61A64bZtKIkFAE2x86OBMPOQBnF2E9XwNuK
JNZJ8F3vo0sXNcsdPaAo30DFv9Sdf+A4JNJSGbzobNf2GyXt8yj0Jb3o+KPjqXjS
3Nfika5FVyzh569eaK0DnqHrL+bhuFzyj3U1eLBbIq7DJnHcYRy+StiUEjBP5Ft+
6PvcBZlJStCcv9oCP0waHXbiH5Yru/rBMXAc0cUGNBwh4DhEzfOQQTYCgPBi1oF3
IJeM8rzfCd5G2eSjNJcr3nA9ovpIjEFPSnjNUEVqOfoCPapJnQG5Iee7EIJgn8nX
6rBqOSuuYhCPK9alJPnjznw45y1zpXVpv5ZayN1uVr97RwGs7K0k5BJEmSSgDeF/
AHykFxQueMb3E5IyawDMTmYp267WUbHqjPwydSSUpbBS5bBkrowVelBswMOG58iL
Zv11fjvupQIT6lflRi+0M/wkLgLWg+ag2shBogDLngMmgBDlenWjiOHhdRQJVkFi
QpoK6XRjM6FIIz900PCmIIHdQRjer+v4pOydYVTA+0l71+XNo7CP6f84G8noXbVd
+DONk2SzvcDowZ2QmY+KGBvIJCFOUqC0MriF9sUNmbUnezyCOvReee47PEnA+PqD
tLWAEmUOAWcp8MQ4/9MXKKdBJUwU01/vV/or5kS2/yDh2zjjCC1XKIKjZ2UqGngf
+tXLG5yWZK0oIiqeURFb90OMtSolpQJrlntMtIj8FuFRrc3OdpRF5orx5wV7AGhA
npcNJmfv8zrhxao7UTClfwJMq2GwerCiNIewph/I6rzu78iKSKyiSdJ17vGyD1Gx
1N1RahUh3A5j5d3ApA67SsdkJJI1Z5l0w9oFGh4fUEpUlUDa24aYehafiqqLMpjf
qBJtxOy5rx7UzQdK6RnQYlTiyUw0/OPPDdgVSxVeAwxE7HGctdQCS4vG0cZkUVju
A4zdmuT0DsVTppftzPCM0To7w9iy8mUQQ+02QtQ22MVsegJAzJFP2WFHRDipu3Kx
uKG9QXmudo7iu1BJpkziAhl1qC1tOZEoQvwdXbkM7mksXYYorsyLE/eelY9aPEXA
9/h1A9OaenhCiwxLy5m7w33cWVmmci+NdugNMWDW6T8iWJmUYpg13g16DBXjv3On
t62raHhPvS/+OHkymND2dOthiMNhWbh7iymCbx9b96H/91JWIYSJYIA4IOSgjX9d
+a5U/ZV+aZukMYICyYWWCM05xGbfXJZprcaSP2jM+DAg/z0n2MyInaSUxXd7ne9x
mxtLdEyzlHZCoHOcvUDlg+1QCaqAh9w+hJcli3idU6LAcY0ka350v/C00G4Qgi6e
rrKWAzDOh4eKNdp4w2II+VBxKPnTsiVlKA508q+TVw/tcSAFaMehM2jG1yW041Cl
Ag30Xl+Qr3cQcf+H6jyBF3T5UC0f8JE0UrdAcZId8iui/Q4uN2abufKlS1alvjQD
3KSTMHAjc7V+3xHYxnujM+NTNpQyxC8Z5+iM1fFgAY4So+NXbWyny7OG3TS6ejCs
9J9xiimygj4iBjI6cEH3XQnbYzQXP7L0GJbryjepzuvFCrF/BreOUf8i5xpjOvp7
kNjaY5sb23wnC+4OTLPAW+4LygRAMplM0st0OKtQQrL2oaw5IHzx1CwdX4NFu684
fuOPD/M1EOEl0EbogUGYts0wfY44av2bXZAPbf/lUpEZMYm+IxnokdOhA89PuSsS
0BmhSZ1lp7mfNfetV0LIiGypH3RC4rMvMsnpzL7dPSHTARMNU7QQhyUqUY4fZnjU
QuJGEkmDQCgv4rxR64LiTlxto9e6FZaiNQO7LI8XQv+x8eyIH0CIe6cLRF1Mq6V+
GOENHJ44ELeoO5YCWfidI3jq+13RuQtjNnlbP6neouoBULQohXHDcOgunBz8pkYP
oJh2xrwJxWo9XidsmOK3H6svjX279BBcogDhB11Inru67EQCg6Mifh0s8ACp5d8g
Rhsep5bf1e7tef1Q/7dBIInNuqDwL02NLZ+KFXAfRs3sFWa2Kadoxp+3mHHflreE
tm1z7cO4LFl0RWcncZ2HpT1GMevV6QTmLkzYCQ4KwoN4B2qQzU/dbT3Rk30Sx2MA
DqoUGK8Aq89a/a/DHZRupKDBRwwEsZWf/ock3egTqQhBH+bhjXfOLG2NVKLzUY2K
oVSbv69EvxJenBaOPTCZRAbpkUR/PgT96IjO0DGgZMOqfXJGl7Z/Drj0QpOF8T9M
yLEjpF9eILNrLss4rwdJfLxRuoI6YTps93BFXThOasPrvE+QZhZ6KgKtH04531NO
HEsnqNGGb3qWQPzqLLXoQAO6zKaF7mZ/5SuC3YuVrYC7XeQTg372VPBDdptssk1b
OSUQ8Ep3ndh76Nay8/rDoU1x7DzoOHLufB4mgBDm7RYuoEZyghWDR8oaBiVsLIYM
T3gjNsJq5SpICqkQ0G3rtqwzB00tRYwSPV5SIYieiayEfkgylg1meJ1ZOkhPCtke
Zcy3751zlF0Jcv2VAxI5Evg3h8u5SUh4eFZ0J1BJeBsN9RsJ4mzv2gOdZ0J+c4w/
7D4aNsCxvNny+xbaBSeMmm5mx8aAZz2YFcJmHH2G0mpqafCI6pM+yxhViGOvsObK
aszUsSEHpFC3/SPl2XphipQ7sOxaqDQODKyjCA6n/7G8xzeRTY2V/D6A1ErCZich
6FZVH0sGyDbY7Wq2PArOrUw6W6HUaRC2hypHta36x3ONyTKlI9cpT3TSfa6jss+x
6zQIP1g20n1XKc/EVtXENdMwvZbkOcmRgWl9tfYStkMJ8t4eRf/EXs9LdQwV60wG
VXudDoaRBzVo4Nh/ko6GyJKteK2351X+eGMwCicF0fzuCo1meDfQ7ssZlUGeWkKF
m1oS46xmnMIuXYGzRJRgxaVi7zY+LkkTIzCXvNg1iQWaJTEmIFHds7EA8vmEDDXt
aDIBIAQpv24+sjxmZFVZi+9yMbLFIse0v8v7cPvexJ1n3l7llulNu8J7I6BlXGlK
Ldsa/jnVxrtqgORWgrIHwzdicEnelCfH+H1jTX8t3hC2AcGu83HDEnh2CIfGXlsZ
gsAwqs9PCKpkzloNsbIAKiYp1S0vXo3YCDqWVjgaOHnyEty3R/Q+h86O5+n0+/R+
Vo6rmXHMukoVUVAwlvjvCimDu5Dq9yFeKZbP72NEgMIXougBFY9tToRhjJEL0XvD
rTxvFFp+xktg5cGUEIRecGatK9QDVqbcTqvlUJfKDWUf+U3uZJRf4QvYmds7D77K
w5DKgT5o6dODvvajIROiHNbwTi4fuBcUVth2PnsMkFlcMXcXEZNPhARAqpiaK9FV
uep0FZrS/R1S+4v+Z0HgJ8hdO5U6jNoagRrIOG+gukYVUtsLfO7Jim8xjCQ2iEwN
YSAWwnUzdXwOzy9D+wLr5mVv74dg5dNSbWoQ3YxPe+ntmkuNV60DJTCapj5U5CET
RHOguQLREPy26IMd4BGFULY2+vMmEGFgNa4kOd0nRlbwweUxhrtv7zyMskZm2Tnb
nSXd1SjPB70Vb+zHwED8+/jK2b/U/iQc2QeGLuPJThdYOPXclNYPSASp4733eCuF
v8pqayUbG4AoL26SqFxgEn1UM55656S+AHoX1s5xQm1RnD4ndwS0qHEvnU4EY7ST
xjqKVqxMSz4kmERns8ON/X/oj18tVAmn2MKhOAPay1W5ISB712tVfnRVRDeAfD9m
+V6FZMUwDZUmwyVZlK2IqGqDOMl1FyrWf7dyZ11nBfAu0/oj/Qj+2VK2cs1zsBlZ
MB0x+6dCsEMFg9IkNJVTd2APoFDR+1qLXOic96hJMMON8B35vYMFlqSWIohuyY+F
UNe5dtBywbV7ql2xGiHk3dEkMNkxt3/Pp0ptKI2PJckZsdzHzxQPoTDSuHHg+RlS
cixPZvZ+ZRXflVBXBu6Qr9/6f4Vjb2JDkV0e5k16Qgs3zlkh6lz0kiUoQJ8vKT1C
aVGRNCsxYCbTL1vxaqh2/zZoml7C0/R6tOisZ17v0v09K1ff4mhaRoUgnpV4wU31
meOIoQH6XeWCEDJrXdplPOZIEjOTQ9fAHiQdVLLPJTJR3ShjCAJiG96ZxiaL+KGW
2WmoGD2txbDvkNN4VNJoAFz6nZIR5kYg+xu87yy+iSBmri8NblLxb/KtO1bik1/i
QVt6PfGPMrUGe6HfR0vftxHpwweOB9WyidpydVKXO+L5ivpB0NBrm5gWPYKvAW2L
XoKPaSzljs6YupZ3C1Z7q4aRiEelYefpOVCqcGAnEfLARBOaCHh6H7zsD3WS0VVu
I4fWcckfnu99PeahwQaYOt8a+ere79qIvxZpWaWfwNy2xEHZeCJXzfl1vOHScSjG
8KCWJsKhDXuwjooQliUqO2oob7r0AOwlGih1e2HugoP6Q2v139xbZataZoxHYfOn
HDu4uqi9daylYq7voOeDowF26EnEEuN34ecpJ4ok2L5JctAXwBWiabcqvYDVP0jI
kB44b3+MjRhZJhUUzxAZcGjBlveTnNyAmzb2wUTd5pofH3LfxTbVILkhbZmBINpJ
QbKATBdREV5NuNjp3o0g0ZX9keyDCD3wCuaKrKCj/AWPIMhr05m+BSsWjXCePwAm
PCjtWbSpXkcf2uirOvrPXz3mDI+LHTYAomTM3baCOntay0cSnaCLUBOAkiNEQzUZ
tl+ObEAfFtGXQY9j+6UccSyXIpvxYniAwldSrDMxYDwE3gYLmdYESu1itURGGk0X
pBCSEw5JgZFRGyG2mo2pSRf1QX9L173AOunzI7uewydvUkbPWYYBBCkWyuLewTOO
pk/1x0Xk+QTv4P7uJ6uOM7rOkRLVRYXWM401jiq4Y+kryyWjjeUURt4OQ7bV/eBn
yg2tx6POi1L+BEKL5vkPt+RG+DewLEwKBuiYcy+DH7ZfrwTGmGH4Cckab0zPNgkx
udNvoKmqZ/kkFJ/7ZNjrbBro7NePCNdceQdMG96gBUVFfamhXNxEJKrIwe65K867
TQm9iMlF9y08FYJzC8v4OI6a/XR8Bz6EyTXNhClPpS6WwzPQgOIbMFzd/bSD+wVn
RJ/c/+l7dJjwbfAt/drkFHOytst4PlAle8WeLflMqT9N74zuoiJQnhhJg05T2+88
bOdCNUXmKg0Sei6iW6/UKmhga2aJ4XBCdbRItULyqqGlPtt9zP7/Opq1vEyODqbW
4PVMH8coBBb/SoH8GM/nR1m0QLjprscuL69Z8yDDh0Id+yxbhUS/U1ze/36FYafZ
++42DSUJ9r8rsEinIgS+z5lCilW1mcGaTihXwg3hQG7ug+OEiR/uPbiQDvTsk/Nn
nEfQV9o7RIOXEQXZN4anc6i5v/czdwx5cPATy9qHp55kv4dh99vQmW8fSwUqvYC7
9xTeBUeNVSA8ANsFBHwWDhENArZ/e5dnTxXOhJ2qCwOoHWaxTuhf+TR1M/H4dUc3
ZGdpSZEl01U4cq/I/atJnTdFj9apZyLUOtbCXU6H0r7RFmkVy3Y8PdG6yLC8aJ54
4jhRnB7CH1cE8BKeYDooVNOVlN1WG9YYNcii6qLa6Wm79FY5NynkvXPaM5xluuMc
bgLrrgaQpnijWezL9uGQABJh0Mo2otdNpJmgYqcUK6Aq/rVch52nXiOp6l0T5bpt
fZ8voOnwPQMGBP3k0an3I933bx4tUD4KaIMYET/NzHMck0TlHrBYm0lb43AmERL2
dgsR3FEtj0K+vMrJs1s4iPd1fvptB/TdT5rkCXjK2B6f1F/Pv0EtuoaanyfCW2XU
ZB1RthGd/N6N4dthEVL+Jge77FSrWKVOCYn9+XBBbQKrXN0fX/I8NwZuO/e6A0bU
Cx7oNE8DBBbrs5kOG/d/rE29WOS7lG543/V+s4v2saK790MiVG1zl2rIb5/AuNj/
p/tSfLkx+PmeTh3b+CCeDIAeGjBFUcRBthPmcOM4ItqHwRnqXulHlEMsnX+c/AgU
nGwoHbO6F9JTvRFQ2mAWTBAhlfFrkGafjPPzCR/cdYIiz8iRgZXxgJOpKow7MNmN
cbYpOJaLRxqFXTGxLTVPm1iwB/760WBS940olSlMpJ6j/YkcM2pgBXDusx6G17QB
P95mSLxeRc+yj7BM1bL+Xkq1oerUeiY9Ag8nCk7gwVRzc+830rBuc5rdXVEHUQFL
weO1DyjQ4k9jT+Z96spMqI3rS+qEMczS7sj4Z9M15xXXZSDd2WgXmVrU7z1phjHg
r/J/6+za3JIT2qBIiT/RraPWs9DGjQyb2yU4yDA7c+srF1B9jo53a9K5HyRyaRZB
qnyb0gP5/L9Xz/aqg9IYXkyKu2wqmcjpQe9/zPDRMBqNOqgywPfSGoINAERLcLFL
Eo+XzRi46rf9e9a/lOvSDHv/kRg+pop+HOkzFWoeccB1x615wpzJKNxh7PSi70qb
uBFbrKmteJjLrt8dzlRLD/t8cZyQlhIhu6FB+UA/rnwUvvj214l2JOwaKld87gn8
kqbRn1akDqNkreoOfJnl8xv6/aLdo8CfswxpPVq2STMO2ubZPrLMjM6tr0XLmmyn
N+Hx07zEcvz+aOtqC56+4aVPDLvcK18gASc2VUu8DIVomgH2BMJtckfCf/aaW82P
YtbGAhiJvh14InXeHMp2jLoxz3vgwMF9FbSk082zeC4OhRERLMPunzGsmeN7emj5
rSHRG9k4yTe14rnwmLug1ADlARUcQ1vtxNcpoqsmjp5GJ/6ZFNwpESZNoQV0IpZT
HzuXC4VyVP3cwe025mo3edplmFpeYSVAlpX445u6DqTFvBdlSf1AQn3h8TjZpSp6
ZjKBPlmaxMKGJKjSl9O4iSzFgz/uxmQm8A8BeSzeBcg8MwS3vLEYXVN9rayT15Jj
aLLqIudcUYatzsyWaHXmAdtJ3aNhxzv/184R83T30meSh3uSUkAAhMrU/JaKJoFD
SikzRTG0vQ2bv5IT4vD1+Nfi6tYDszn7kqq+Ri3DvfV3Mz19UgWVTWGCfdoCkkBL
QrAs1Q9bHODUbf2k9ckp6Loqe0sPJ4Wjm0dcRiEdjuQ2WBXrBoCTK4OC6DrtYBe4
DcM1oK5uuIKWpFcjpYpjbA2ff133Mh025Jf96GPGZYGOy8zJA0xL1UpkhqZ78xtk
BeQ3iJ9p/4f1OLiYJnKswuPXO6Ipnfx00aB6/qNXOZk4zxtFNKmEXU2DqNargvd8
kd6SOEvfShLcwi03SGST6QoxkqBIcVd9MdqSP09JzbAl2JJquJipGXOBFii/OqNR
lQcacf2JZyf9xe+NmwxZTOoLCzRvxWAd89J5yYbCya204tu0BYEWqG+BKp7/ERw/
TX3YNNbWVNdrjwEsRb75tCAxiw9HFMoTW+0vgZr/Ec9cCKouq0761lNe77PRnenP
cntiN+bEBS4A+zS8V6366n4AoQ+hxPYMWGQfqFRDzoBNp0QqfYUVwqjq71G6o9vg
q3w0Pr/EI+ha1OEMjozDLfilHJNiTpdDs2xYtWpb6i9oNSjcNQ4+h/bDpDuEbPed
iRTNUdTvRymBPDKaSBEwkg1ujNRcy1GJ4ByCTAh3W7jtTvJ+q6vOOqz4z2t7bepy
kK8vy5DdwN0KNPP61APnH0p6QHmuxpk2q3snmZ00y5CA1oSjiBQa1Bch9AanaxWY
XBbMf86CPnqvKDoOK5NhBD7m7aswYclA9iGFQ5YzYtTpFG3izdrfyvYp4xzVK3BT
gn0sKsnzn5fNCr7psEU3GJ5LWla6O/aiuq9LuiTHTRwKQwE41dfF5F4ogoVg4DoT
zG3nbYo6/unaKfbhrhhs8WTH3dSungE/QIHbPK7Yhd8NSl93JExYlJ/tklTZFEi6
ldFBxgoA89vKUyEKwkDGNJq1B+GrMDDkqg8VfdcBihPuoVYE6c5JhtUIpRTzCEaR
cLG4ESFk6G+sBF49sqm4tPI+2bVdPJsar5ONJVorI5mjhi6K8Rl846MrmHPK1urb
wK+7sqKe5+LyxbIL8sEAiWeVAYJv/Vk+D5Vrkqd4Ik7l0Uo3Gxka6gJScf4WZiMO
ycLnEZqVvkOQlmc7JQHtHF1hQHGHTIlR5vkmZKofVwAyoBwasaUdYFBEdZ/Vg3iv
IlhpnFDmyVJv0KjLo4Zqbg2Kkz2vwoJcoR9dxL53U6j/jkRAh0jyxE462Hzao/7h
4YKkTZwqCx8MxkVd1Y7jGZhRXzD5oG7VXSeOpAFeImAmqKDValRb59OlheYzflzD
ZA+uvjQeVwAgNVatGTNuCcROB/PG5R5hEXS6ZFG882LmGZ+oy7UByKz4Q/EcBws7
+Y97uacDFDScx6TW/E6qJV9tI4WkWA6r9WQYN5t76ADJ8NxyO+5l3kdbTquL6Rbh
kdxe5lZCMjan419xg3cQyu+kwVwXLPF414rdoCzKLhMOThZ30Vk1h1DrCQk0vXwa
n1VAhb8eF5tHG6jFpGmLcmtI72cozMRHygmb+iJfWjXiU2G8N27wfDGiFuES2eFk
+n1pikA0MNXfkBuFIFtXU7IohaFEaskHd4uq81k0cWdmIF7TdTSQMG5bMOMITCrM
ZBGzTuMp/dMxDFf3xRJ932R5KUWMmEEy3nRKX23lxIl6Es9WuStna8LSbUY2XXvv
phUAEh/p/GaY27zQrYZikxgNQzllShJvhJrJ3njZBj3cYaCRHkoAbDqssTlbn4/P
Fn5R473Z3cbqCRJmcQtmSA5Rpaep7dx1buuFwmZYl3hxX7MnML0NWKMpMov27wBl
OTOFUBdQ3C+fb1lsf8m6jzD4KA9DBXhuHI100JQTe8vQXyXiHulAccVsOJAF4ACx
rl6gd47ZjGZvuy3ng8TFYePQ9tNNEhATLRvr5n9l52McfnMIFYfIjrO6a4lKS3la
iQaB9ZYKRxlvEZn21S2WSXBVzlgkp0714DxyyyufHgB2rBlXaEviVgmOtS1/eXfU
3VM6WnQ8mXaXR4alOtn2wNv5MIhKHJKqeKBQ37NRlZ7IK4JYbnBkORo+76gq7RUA
XvShscVwgCLB6FkWg4Gyjat5Y71i3IV83lWxxvneR0Pb6SB9XA22Yq9oIXG/ZQU7
YDNAUDQGpGn+gUdo6HC2+/88lk909jONPXOqn7sahwOcOFUWivEG8pKGacfnYL/u
SxyEkDP9VWZitxcM9VK98Nmz6+TgXIKrgNo4fiZSRKiFx/nD6AoGS0E7BTwLzldK
rS9f37FnOlIpr86YTSfsSlZ28zd1Fi7KaPxddkjCvpPK70tW9eRZe/HKhpVLjxHM
B0tmh+QO/ymGr/XJrYoVXLbtflyYCE0Vs1YPfxGnluEb1VUB9Gr771+PBH4qTkzQ
SpusuCZAgJXA1g5a+3so4wKIndan7AuBL6tfztjZ6k5+efIJzhSPfQkIsE6f2WSG
Ve07BnBK7gsgWhxi+idlhy0ESd4/hOSAwuRVTuWNS3/6xCL6APlBhvCnNj6bxTGw
U7EfP/T+oyUdwfxo4jCL5MtXVDHRxzbfTkRporZtOJnRbLj8prFSh4Xg5D5qzneP
RfGULL4aZ9rBUc3iQOucmIAi1KfU1LtGt3mR/Ks9/K6lVluJrYtrkS9X2ROUjb3S
puYhmHgBrSlCdqLCivf0EY2+5dcYfWEqH06Pchql9cbxoLea208FiY8dTn4EkDmE
McjzhzaYgaGJODI56GtjMEn47RJ9jFgbrVciZapDgXGYW2pmMlCCO04+lMzNEkdY
KYa/cNiyvrKCsy9VrT1SDB/+M4+Qw2t0zg/AZcluxQHFWLIRb99c7ru/elx3t75g
9XIkhK/dLe7pp2SJ1dBR/lDcmPgIod1JFDI6x/pY1xoWVgPOOpn2mMJ4TuH7bhxU
CrkbvlJdnI1J/CfLUL1c6Iy6PySqoGaElFjYubHbyUC8DlbiIwHxGhPmOYEPocEc
FrGbi3CP1/JtKo8uj7TV8CIG5MGJmjx3LzeY7KolrFvYrQAEQzdGq2YUK9ORbxoz
bQAt2pU1cerqZn6NLrFJFRMFLgRe1XPVXKuK3meGlKQnn3iVsWmE7TFtFGw6abRI
OZMKWKH10CPnWm/joaBvbFIeDAWRRF+j57kWSEdNv8yMNeoQtmLk+tQ06VdXvv65
UWbdy90qZramd8BDS4jBHnHWIqkSU17jGCj6F4lzFHySqCc3VeZV8npqkdVbM/gf
ZWXrMJluvxppoPl98zmEKjUR+sZP8uVPqG5YccJBiI/M+Nv8AWYuH2CJKMplsJDY
inNEInldq83xrR0ugyx6E6Svhw0Lp4k8Z90Y9Yx4Ydn+9Wfu+jxiaYQBsFrjMV35
XOFj0j4xhbT5M/OUqnQ+zESw7xckhttXHOm0++34k/kcyrL0UeOoqClLYplm5IKy
xRQ0vhVJkp6VWPd8QaQsAE38rVQpBi35iSJsm8LAJHhK8+3z37V1oem3dJ8fyBI9
HANRu+jtWyyaldAtu2kO53B6eXu/Njx2iveiuXjN4FXWtDFkejJ+oVuoDH6FKJz0
sVl0Nkm1Ot1EcaZPly/bOWe3fA2YNhl/e9DXOnfQmPgFFpy0d/CXqITGnG3aZCY/
yK0/jYpx3rIRFJhULeyX2PVnJsjWbROXAMSb25tiTsqxU/gGpMD9m99I6JewgMyl
EC+fVjB46KWJHpWFZvDl1Ri8+wkUivlaL0f/8Mn/FN0qDGWXus8hmT6zjlpYUAmV
3p4logbWT5RLsTBTQpzD8mk897lsoDiDFb1OKOp5ZKjeFfWybWMx7FHwV5mukcwa
5UjYr0v8F0xw+dCKkMpPV5nncHbN83qvTNss7ABJzr5UjH/2Qi0ySskM50UFsirx
J30nnkYLQ4favaHBrAC4DJwy1fp+y2vHd75jLxkKJEFtRkbaKE05EJ+T+hDyuvxk
iHdrP+Hut+bSaaeyQ0qTaxkilYjFKmDSfXJoM+61n8uX3kVNIZ++lFTUPFl9dEpv
NXbrPi8pnG9011ABuhEjXeXgVe8bj+TekyyDy3WTZrYlXwimkKCbwsenCaBNxX3y
xWYjaMqPtpmScvUCgYPh+sY7fN9DfYT9cqjo+7DAG6P/PkUCcg3+mNN8xs30GbZ3
Ppx0934Jh3ps9Kxru4pOVy14+jiu9oBMQPxGHiHIKE6K5cyu4jYlP11R6Ue9/a23
iXtK3ld/JmAimCiC7NMwc3lbOO1xdKmoQZ7nlcy+hi9VPYusEQ0K3AjfOEaMOKt9
UIMI1vW4VYBo68MI/JciyNu84fw4YbahxU78B8fyU3m2QUPwMp5CiD/4SGjpNAn9
U/B+k/lr4WtvzVJwxGMs/oYL9vfQshMZn+28i/3QL32j/u4iA8vEOfDLVvSucafN
6YVIuwySQRgpzL1kmzh1r8/arn9fbz0Kz6H1C0PlrhbJplg3wHWtDGGQckQlKQ/d
Fh98QbqJotSKxKb3uzPvVx+1QcaM/y6fnCYR/8vAKQBLJAAEjxXWVolhQaKlyOhI
YcI+BXBX2UExRTFz+Hrj021uPczFcVubO2/nQmz6qf8hCApmDL25hMiNJqflGWKg
I4490ItlcGLKy+5i1bq2b4LvJxsqa8Yu+o1mzc4dyt1oAHCCJR969rz7xChqJfVE
C4sQHmHLrTCP8DKni/Im6B2Xz4s5xHJolHNwrqQ+v4xciUzRskvCgQ4h6IVsjuEJ
EzWT4Wk0QynPfvFCtO1nlpwelc7bqlZWs/+CjmFy/xag22lmFRhbpOtXRe4xdJJZ
iO7MIc9won4AV7+xUsxE/AWyRjGOZzJCGO2dOhinEkYRtw9jPwvlSbFhtv2hWyZF
CcZ7OmitZGHzTGOs0qzUr8Tq1/UsaGKSmarn5ZXQLFuZvKoXDQGJtM6UR64sjtmX
SduyPgVmD7WwjLq6oKWqulDe4hPzD/TWN+yaBCKrrp3iGw9AyvEkkEiYCf+LdUhi
uHZyTtladxD5MDFa2yXC74mMihFvlZy+tvNojpArhv/6w7OTO9OFZNfLnVHQ22nq
buUwFUXG57UmbR2mU3N4LwaRGIrWWtUeyyTY4ANV7EpooaxtNpYl/mF5HZHDMUYN
MG5XqfD71/wnlWZnv45/WMPWSTGDB0bft/t2zplpnnywKvm9mUGKX2/jBM8pdaPk
/Alw3IsYDSD2rr1UM2/q7JYj3562MA6gzNlBLhufEviiRuwtrv7BQBCeezwHYbPw
poulaFjLU+DfiqiyQ+tDSfFNvwjv6toSBq4LFOsu/g79oILIEcw96qSIqG0PUBAi
WAlPi+GS9SdreJ0Yvm+4oFpN/GLpkS72Yn4DuLamII7TTHwNjjtCfpCxggPUPWO9
mhANZPSKNX8K0oFkwzUq+hH1SFkhyiC9eh5d/fS1wR0lPgpfqWbonaJALXeLCL9a
LUeNvvZ9HWuDVWI0Jbu54lplI2lwz9yZz4u/qfhpORr1RdEsxmLh4OibfpoftPAx
P+yzOI+59tSnZc0zt1H1AK8u29yH+bxAV9xbgJvVyNeZ2j9AErVdw+YvKre0Szie
DRrA6w193XxHH1gETrag5AudISioo5Vz+6zYyUaP4AiFWhF5w3c37IKjfXXcNqJL
l3/nWJhh1E5iItn4bLSxVX/1HXOqozHWlH2/T8jyxVMbnmnu4EMTBprc54PPQZkr
4vEkmAP9F4BPBJZLFHNK2NNiUx/SKYznfZ6h1JJGhCXjKZs0Neve6T7tA2yDYAUH
JH98qcjq+EWLkv+mpJlPfk8Z1g5EhFz6tCzF27APDBtM8PEwLhDTjA/jT9ti/cwf
/w1vSMRDoQlrmRerditUnO/6lw86K887IatZrRo30ThJ/U4DmRuWoITVzYkmVlMa
gaFGFN5HhlCaV4pvIV3LcDJSuRPT+2HkxZGGzDPjfllnhiPL3a1ugXCXSM34QRJ/
b/8MIMGXCxP/OQAk3vXW6hJItdWYaCvE2gP/mACjzAd/OvLvtoumCs36FO+02kWp
D1ZnA6L+rTGHEBmjTfzy6q/Wx3GcfU0FSDm15/wL+bKmXdlpWzK5pu/GgIlVshHg
1vB7txZt01pfU/SRR2x/KRMZZeFsUMcVylCRaJhRnKFelZa6ZSBlrkcg5yVzsoKM
yDCud5fZDwzgX8nV86HE9ptRPVdHbUHBOYZinK/4u+DUW+ap8KPNDLMDVLqv7HE1
snZrDMPDQYHrWYXkjZCogEPFmiCEo6q40vxAVfTebH94RUNdufUi+erxeG3wkvOU
44GfcPJGDV2tfy9MgbgH9NPqHN3WKMIPy0PJk0y5ZgyaliZQp4IJMIqhXrfvtBdV
CnGrc3DBPpQSKzM0c0IkiMxg94gKJvAISPZvHr5N2/nF6uR+6EDpT6c316/a30ti
P9+lCP1CIgkfF6pG6hP4XtXpM4oMVw46rYBoE62+eCBetOGCiKrp0WQgqkPRJmYD
FiellXG9TPhI96JXcUvCUZs6Symu95ypFPff/sGdg8yaWYjjk/vtp4kbnMOtNu7R
ARJTwkuMCCmrljQ+FwC+ho6TUVf22aCLZ2YnuGeBjxA/kh7OnKS3zp+WD4BomzrY
kTMg276I0H4EsVzDCOUgUT46rnFswSF7CaazVkfq6ysIrGsSlyu9dP0K/m5uKHwv
+8lIaUq4pSmZPVsQnPrnTL8tAlYFKu0V6ZqssV+mMHpKCmKqdTnEtpZOtqQukr14
eD8/r04XSZ4HrJAchke/X63YBL77QyHAHkpy/IEIzroTCH6shed2GhmHgEe0/K3y
nXoZlq+G6nb4LDeEL1y67LV+Ug23PFrdxJMgsp3S/gbyoBcV4710advH09ogprBo
aVRzdMBKrj8GRKgmy9MtRBrOHlkbI1K6iIDmlQ2QpWx3niFllcsi/i0vTsjJdA+q
VGNKZVKKqNHOlKzJPY9F7LJ/xvWN4uv07JqljVb6IEt4FoIUgS3Fc25dnqTMPJ8g
WRaFO1gTG73byZv2ZzOz+YNcE/H914MHf2UR2V3FQ7rimT+lgKf4AR9mYhOsXkVu
i/MaP6xDF2bRlX2tIalBGq3B1t2h7HAeGh+cfnMyrWZAN4Jp6qB8yLDTn1V6UNgM
mts4o4Af6iZlwc/kc5Chpyi1SnmFvFzB8Fl4eP3FXcQ9i1uT/4ImKlss9JYtxmoZ
cMn5HJQ2bLW14QgwjtPCOSOE1TB95ZuAw5oHlnzWHQt2brQQ0uv4jOp+Ybvszqh1
0SAFk3vOsAZsD0LSJmYfzFLzXVDhn7kJyCUNNvQy3x/+x3/6Lq51IO/xMASwduMy
CFD//0o7WvzWJ239X60S3S96p1kJYC8vjmR5hHe1DkoFRgvvlthG0IndslvXpRQ1
eyGS+S4DWxJy9W6Eb6brB5RFtamhsS7DzkQgB5bmNGgOtbGrV9uE5f9aRBJKJHpT
ejBI+60k2k+GGTqPtP2+1sOtwz/f8VQvXPs74IzIkoKniA0ZDLdczy2BTSddcY3d
URpTO6uB+p13NkONRGvrLFhZg2hXKYghuA1neltuw2oQs8ZQ73CI96C3r7dyVRjZ
RCBGI+tg+SnwzUX8oA3oQaQC4O34ssy9+vs2Jpp6oJ++hZ1xq3v5cI0rMoziO6wt
E3Aavq6nT0mpUHyzi6klXKOTxoQFH9K6SmRLawAA4BzIJmiX4QO5Vu9UEPqbLYn9
ZwGGVSgD2nSPk0CCCIUSqvJl48S8aRChw6ZFzC8qUdT7/gNwDY2d9TO+VN7ZpHWl
W/7HOyOX3MJRBpaCBplkhj1qvdij+R6twKIuK5kYzY+PCnpufPgdQ2gMTB6Ga+EJ
sPlLGko4RKZCpOnr4uUoOCpKovJi0OtSiG48ySpIESysd4AkdF1jZz8RRcdT7U/p
YpSOPGLch9t+skXi/egA+atTKphCVAKTeRyFHQwJ/qzPiDIotrL3zenQYF3YHVef
abgukj61t4upHUCf3Vfwd9WnAgz8KT6kur3I64e3OEi8v+h2Xxj0OCBGA96K+nSk
Zfi2BkbcgTU5KjbZ78OX9YE16rL87OwjWnMs93VENEbhAF8erc6hwAH5DjPrRgcJ
RUH3Nyp4QU+FrU/vH7U0AwF4rpbJGoX3NhqCcwLqWuEWJtlAU1n9XyqoAZRSz/Uk
eJausLysIPHO0dM0Ewmj2eL4tkqgc81hTtCxJ3Z5iYVcp+C0Zyt6zy6MSfJ7iU1g
igggfyKOuoqSil5XqGyxZs6p7OFUGU4a+v0r3rABJHLFbPvxIpbMHo9UDhP7l48u
ISOzPSBvWq6MHJ+3LbMNvgrnSzRWkiV+CMSu3g2NgXQUs8yctdO+OwTuOd3N3XUT
mIdJIubJeUHpKX5tckUTeNp+O/9Hjwqa+xVovHfFyA7LCzYP4fWQ1CIxEB7q22p7
5nTuGQaVm9i4J7W64XmJEz+IlaPvpHRBcbKbe0H9reRGPvW1vWqH/atGr2MfKeuw
m8xC7h0Tsxma/PJa6rfUqCJik0fH1DNKKRmXbsImrJSCTSjMEiLHrl0gWcG50JdC
bfOPYwT34RO15H87OPeti+goVtZFkkpeZhex0BBPXb30PbbpHhAgzvzPypKalAG9
gSWYEs1cpEEsxU14QVLFdPUzusSM4grIDvG2WVwUxiW2Hn9rv7jaXZrllHHxRlQ5
1KfiM8v2X52r0sy1E4uiObQd6X8UhkdjwY/xC/LcWcF8dGVyDnRNUKDrooHfVCUM
BAxJIzAnar83lwVuM/3NAqLLeneT5e+IhAMeUAHgbbV+RTBEyB75vxBQkSJGH5ms
MI8mHqZdsKtBnhqBxT+YxjED4nzglRar944LQ0gxthdhJIBlwvWFu2EjM/VQtOJL
qEOk85xwMsy8vgsWNOUp3mMXh/vV5livlL4XDgnQ0CLyafvZc8OuGdoByAOVORyw
K5GxvbX7AYYfmNoukj6P4HooFEqwduF/x8i7JmnPVXY2kl4afKh1YM1SI2asxRQu
DbE9KnNYLtzsrELbD1DFK4HuTuTICLvP7xN1swIS91of1amGj5sDlv0nUdprlj/a
JlGyGLtgTVhOibkiGsK657QSSSjntUZw8191R/SDBOobrjkBr4k9tB7wp/yI5CAB
xHVZmmfItc7CxNBZbCPRTRe8eTaScY460VR86KvuRENjrJRV+NPERog06yrm388g
Ij1svbtQzVHVX99YBXIJST82lgwGfoJWIgIJbE2if/HuqXdkMd94ADYVMA7oTxmc
YX1ep9XalX1svlPqlOx5/IbT0Lzm+9SZSYErE9CYyRQvzVpI4pcAeToMfPjNwt9U
XIZrsYGp4XMqKjOkJXIQjCThlVfIpEELXX7BQ8m0PIASr+p4bo1eTuPxgFvpv6JG
mfLGg0YGBZK1wDwSnKwDKwpTjkc97u8TATvEzyh9npLwPumcxWNZSdi3WdDxCZp5
U7BWzdNzPVRD0V/3N0ycob6RrwRKC0hsOI6zvVlDQMKfepy7XgUSlGvSTPVk8RsJ
CVeX3isW61spllXX4FqFex+v2AzkdLdhJD68YTfSU/ABglPvf3XK2lIadlvD2wMl
m4YGbLdyy1Vr/34aFHDM+Rd5dXx6oEI6I/ciPJ2/zbzM9O7XfoWfhm7IC9vomhic
U7ABJKECpdaA0oWEMcJ1doAqsuwv9wCil4U+wxnRu772aQ1dibgyTjfGrvc368sH
M9+kftdOVYEzOqIxf0j3nt0i2Ics6811lTP46CCTAkdxEN5YAupW8XA4+otO6WZ9
MAbrDL8+30jcngCaqCXsdSKwYLwkUhtQgo+RxBamgO+cEvvNckUnoLVMf1x9DwmI
8tiM39+QEIscIUOE5NO3IkcKz4p9fmQF/lxO5XXsNdLRXjxpPOknBQnPViA+f5uC
AFuCoc4WWcChlCkCtUYvkqhKzz1gYSQlaVj5ZrIDnTK+7PyYb0mF+WlKCV7VGe7i
PmIAgtc9HWnJ49BYDihouxarfe2KUYgl++80fiIm/6E+yAMI1cZJjXXNwYV4zffb
pcZxvM7OknH3SVLW2lF+wtyAB+k3zxEY0Tjh9FKuKRMCRr22jsu5nCXu9ptRMENy
eXyyTFAc8Y/UbRPdPBGJs/nFynzipUSoHC24SRncdUXZSNONJ9psH96cqzoTeukW
FReTbMczoQ4iCFRm9K5xTOjkCVAjl60E1RTgRHtQ5fDzP5fc9HKyEt8qS/dAZhPl
tj9gYRq9xrc/htj1JG3BTlGBhD59GjFOFHvRpAy2C3SF0HSH4x9SA1Wm5Wj27uE6
NaWERdUidleflo2IfHNrzRzXRvkyjQ9f4mgLuEEkGfpM7w5N9Rqe1xTqdKAtnqeL
22dvPR5NLxtwTxFZnaOBEH+tjEKQld9dNvX1trXsPHdE0fuGU8OsIXwM/hR52oy3
c9rS48cCGASKe2yXm2PErcfElP5jXLGIXUEDTbo4TreGsZ6xqOU3NGqm8favBwUN
/Odpfm+emSwDEeAHHhn6/nF/roZIY4t9utGUcrKvKUX0273U40Lg5L7YkZSXfoGA
blmEulG7bcIMwD5Iup2XMnIWKa78fYpJrnE0KAUq8FwjpsYQLJAnuWp9LIWNwafD
qmY2xYUMSXMES7tyDgsAIq0xF2mIPAsCFHvBSJovHt3UHTXLc7YTWjxCRB2MDpF2
5YcDWdyOUrI65ZDupjsDa9Ctm4zgTE2HXY9FS2Nk5jtsl7myZawhbVscrBKVLXWI
E8aIn1EZC1/bjkK9tfHmDya1azEMqTl1FwsGaDUhL175Tg6VkhAG3ufeKiWudqGU
d2zH3KdOYwmU+VOqXXo/x9PdAZZMw85V9r+UVxSacvr2lfDgUnaTrRjDUB/xeFqt
Q2IE3Wdjg2FlwE2gsD/I9sUzDDrjsUMY9GPbdB7CWq+6RiGdKo5/SjxuusQSW+gL
pFXrJFUNIaWcXQTwfcv+EE18LgBYqg14Dqzsi0nUTgcYldJyPa/E0AWkpamRyMt1
itySgjRZkU6Kh6XwCxHXr6h+YDl6z378e3faOK208CwL/fdTkMYXbggUDQRZuoG/
/BzcoIiyXHj54lEDXsDbwrwkooLrX/jgzBvCpWDCqqbH27FC8O/LDt6hkQ2Dqnji
AO06we5Nk8GBokBGeOXamCMyjgpjToNUzPkKLd/AuhZcNi8kQxAcKvoEZ83KTrRw
G2hU3n7JEbAHM6asidkBSlNYyd1tE+zrL8gtxOWIc/KnI49XB9XmnwjAaVi/dFQC
1kD+/ZBvGk/GnWC2yAAjJBfAkVLXbj75MN1Xyhwj1Mx3zulg+QcCADK/x9stAWbm
V9MpzepRwv51ueulyaTVU9sCZwbY8o55PN31HTDlF9ID9iUo+MDEUByu2KlExj0C
yVdICVowq9qj66utL4bHVZmDDmXgnVDJT2D7/qQh0rQjmSaYzruqBgiqCGxwpB15
+TK1iTdzjgOCNIEGyHzf2urCRWp90YEdeAxv1cHCPpIaWcJMkf1xUFwPLCE0aSot
zxlj6mHljFaYhh/MUNTl7DDJ3uqWs8sojogg0OT/chdv3ckjtrgGIB+w9vJuYx6h
0ZRY9cqBtBXED52CcXLTnDviKQe/s0FRv8u9lm3Ss7IFyRrTCKmGTIFAdqiiBAXo
bcOGweDcnLAKMw1lcD4+1LJ2XUAHdbae/Z2xHNHL4KxoovCYl010KVmktYp28U01
UhCz+K76d/gemAN8wkZL+9tjLi4/Wnp1VJtp0pv4pJGS55gmSSaQYHR1E7DvvJB1
mgS7r6t5YvZLXKdXWtGIARNjesDbqokfWNe7rjPNeJrzBbULc/UyusIIrRZ81/dh
nl6Mm5egEu2vMVA1Ejhp07QEJrh4L33DlfRnAm+JHc7k84O9r4MWoRmeeOkq6MCB
PII14ExprKAp4wXJr97SxDtGHdtD8aQG7B+DfyHurUNXZTSjOUFJ1E7AbTabxHx2
ydhgGvxANPlG+R8zWCRut2/UStSRxbFH7H+cHXcmXv2FtpYObn9y9WSNiwIU1zLB
lD2oxEDWUx8M2veiJjPCXHT7XUvz5l+5fUWZHpvws6Dylx3ZzkUff2npTPBHaIBv
kkPj/EEdN5zbI5LotAPTuVxSRgNZcdnWrDVnNtAUTLTR0bCQUIJ0A//gsW9kI4lo
TEznGHVccJMjTX9ZLrNg8gwqb6NpJgCr1CF4mcAGBTeaUuWtZ/uMMPDDVuAc37Lt
xpxNOWMhmO6aSZ8tGB1T0QXCsm0RN/zMsjYNqq2L0+023njeDTcDJM15kegU3H3D
XJ+9C/JqH8axT+4Oz9hQFAK9nkWrCCSTXUueXQ/QJe7RRZMoTuSgawOoWneLwvgv
NAFDpDbdnfh24LmoxTufz/A1Me7xZ9CYk9v+ROlJn6gBeJuFWyJM8RASfqQLhmlx
9Kk9O1g9g7f0vLC3QXI+6W+kR8LAovGOBur0bmtacRTgJzVoIMnVbHEN6p0h+GGM
R9yxQ5B3+6jXVepLNFxCKGEFa/N9nJYskZoQjxKEH0klW710aFrBkf9JlZ4UAaMc
vak4J42CRgLJ20sDqboXLvhcc9iJouYWGKJ/DWxY9sruPlgAKVKbmI+Lut9Ufu+W
A68a8jPocJcmrC++O4oJzfKuese2OkBiuYNjj+QogKdL0i4BTstkG5pFzSMjF8Ic
Gy40EnTKKXN3wgLfIR+WH24B/tJVwvhF+ba11vUDO49MMArIgX2orTfLErK9kgxu
6VaKkvSBTYlzOR8cO8UZD6Spl7RKA5Un/SfaCUq9c02O+SV6UG35AOOfVxs5us6k
IXr9CdQh0o9Aaq0TvQghWEu0nxR8rN9zz8hCuTD9UhkqJjH/gXDwnZXUTC/bk3Gx
cP+9ep1u99B0zZEcCu/t2vcofBdvIEMot4dfuDYCOIfH4conNVIlzY4eq3MQ9kz8
xUlQleQ32BBGcRABSfhif3T6t1L3hgjEtTiJgKtEi3IWLjkJyEAexuupfV99uH/i
SC0+N0f9eR4AbyaoAww4L217/du5g6JkBULqcc0PAzjJcatrJcVJwIsErHYyI73l
/2xyW9aDQ6TUN5uunQDnJzKp5+IZLH4mEl6ffNxMKY4v84YhBYF2NapHHFSjOVPw
mdoSFNM+oao3t/NWYmN3qNeq+JcNnX6rxuMdm03SIljuWF5L9g/LzuINs8VVxqC1
PjCYibCXU6NUGjbcDt430TTmf+f8XTC1ilvE1K2XWvp6yE2YT6l+J5XbZ4dcQKpW
A2GW+6qFPFhETbjDDGzne3kk3XXYXZtDTlQFqQhV50+qaPbqOpKijpSBQITh96fG
piA4TsP3OMQXQTGYZWpDVl7wK/nwZry5ZTHZ3WiIdVPKU50pT0GEp/lTFG1wy5OI
3vdPCtdM/f7l/icZUW0HkHil8DzCYKfrMzduIJJt8nEwOfE1G+1OzWPqz50AmvoA
SUWGyz/clWB5CEQFBySVtgJ6enuWIL7hr1AqjRHIl6M/E294T8TEel6AHgd5mb36
cA9jokZvFIQ4VZ5tSqPP7pqF6hSUCyFcKPFmLd/FPA6/pfPJSmLe2IBrW/RL631w
7rjsPrzd6GA1AUITyFEBqvct/FMH4W7F4KM+DF8mVjw/0k8kwcl6tPOxkOyWjEVM
M+tZb3EFjpe7aPqu03C3YzP/Dy3sUXDqXc2pKtpPc7hslVPO6hmrsousFSqqhtlC
U3NpUpwef3TVwnhCes4XyEQoSI8z6JXCReoCt7/PKqrC8Vs3m4y9YwzwvIgj5/iT
ANN8dCZIqwbganHAlIvtWAzYKgiQEkggduMRdl/txV2iaZhyxf3T8NrPFaf+RWMQ
VTKYllkIwOg+9D5kIf0JFssiclSQrxhrKSOVp6tjzuO4Bl7IASc5+MNRO1gpZi/M
+9NiEje10Fowv4HM9ijrKI0kL/qsokBf8R3r/JzwmddmEc6/UvZCwl/nIp3q5gQ/
mvWa0vDw0I1FK2hSC4mmKAJijkSHmLBurq9no7VrLDISum7YBJ8N7w1QffV21e3B
ulEuMnjmeP7hZKu9YHFmhm8oxMVN7PnJASywjzhXUAm+RXzTmh7YeEH1sOBNdUG3
typuq/OH21XXxNAIliEZdxvr/nRJiPHBAuHXaTzsh0LWtWTjkKtcUPUirfSnBqi2
7pJbCFeFVAZFnxpgO5DHG/6SjyjMO9KNly44nraPZWFycMonFeXCYMkiSaegXMix
SSR7xGT8htB1CYjiFK8MfsdOWiUX1hn6Hl3Et9p9k/dN7l+5jWQZIswF2Hkg42OE
pOcH1MvzgJRSTFnL5HyIdVu/Z3fnwEQEm4w6ET+zUY90yg078g+jjKZm6lpmLj28
WLDxAlr2bCwSkeWXFbQkSSMh2eEljDykFu6ORfeCsTevwJyozIrsQaRg8Jp19Ssr
Z4lV1uMKMFTBQYEtt4sUIVCvk7rmsijRsqquUKFrSeqes2r//D0XnErVjroc+hBe
GTFmY9eFWgTCvUGo+Gf//OGBxnO0s2NSua9daASRGYBAQWDd0j98o0fLNk+sMlbg
HddetnV8s390+cW1AdUSwrW+1dQxGcxD8n/mG4XFHlgmiH7yA/lFfqOVU25Yu1Z/
6t7yJjKVcBmYevVPqrSSPNQXG0GFwZcryexVMu7Etgs+htOzyu3ybTd5zEVH/2re
jfEEls9t2yyq0AkxDMzg5NwF8Ey04F4CfsXYNJi55UBUaJ97tKut+cgin3FCDBoJ
pj7ropomXE+f2x5sgJd+6BIN3CCkX1PV05Iszd7IgX7xbJ2JU8p8Ap+xzSfZJ11V
hoVPyMqVcm97kFdNhwQdwdeVe9OG18E0f+Oytq9+fRAByASW2ns3IPw8IRZJMj6M
bck8S1R8hbphwWNqbdzQz+V6MycSRi5KzKc6OLcRr4TLtvNgeVzaaBVwWzcUAhce
39hoKrmAKjbKMwlSupDB+eidYVIAIdj8/0yQt/z9ufqCVPdX7cWhmX6oUQc14Nob
c/UBJWXa6bLu820OXITT/InsKQ0cIsuEDQVocf2dMM12xx1P3KouPbnhnOOHuYMi
2gIVHPsThihCNlDoWX5RNlDvWYZDiqjqWSx2b6sZT25sEG1k26VjFJVpb83rOTKf
KC1tq1LIlEWXFadI8kZOQYtPoTVLhXdR5SVxS7j3F/4/H5DUZH9wVBJRHibOs5b1
vf2ROSUK2xBqOf6CVLbn5qBhWkyCoTfKXLTQVFUvUoungrYveXhOV5mdoJB2+tk0
sODrWOpQXjkkRKXEiQuz9Gu8jv+br8E58epz15VhZN9jmiXwAjl2NLuYW+PrI9XI
/IXL5pVHNgbwe+ThuuKI6gxw3YQzZsDw9mcPlHpxX4dof/ts9G3HoOndxokQB0Jb
SKXpd4R/EGmwq/ZJuHNV6c1vqPWSgQS9G4vYAXZZWqeYYgQsY87tGTAqcA+jflfJ
QEO9cEW4uUX0Yb+LRrBEUdh27SP2W0Iw16Hl8FAKwtT/+KIlrmoCMxbxBK1uqm8M
oi9j+C4Le9sUh2NpQOD8XBUk+G8yFbHOBviC+v0CJAnIZJF0XGtXpMGvaxPTyh1J
h66i4GWd2C1v6RdA/C3idCgzXXOWVG69vNEw8+9+AXE0oT9zUgUypxxI8Rd4QXoO
b9lbG8kPx++Sli1fJYCX6ixjQ8kmHCRhq5IX43VxvXfW7RX+Ct+q9V81OTijgHST
AB4GaRuL0kRRGI38j+3QrPWQ/ZO86m2qs8ovNYMENHCF0R5VRSXW9lr2aa3C/aQ/
dtAm4+YJfimccFKJaqMe6HyFplFj0joJNm+BatLjZxkY1E0X1ZejZ2SDcQRNsIMb
uVbosG/R2MQK31C3Vkfj4mK8Ty+Q5IoA0mVO+SvUkwtuqZZvYeRwNjVw1DfTDxY5
1SV6OkBmtM+0qIQQeqLF6mGTiUShvtndWgxBuafVZHjSQwxLvZj/VZZFCU5yCZ4H
ImRDPoVagQH3SX821SwxP6HiimlAIDMPQ9a5s9zOIsb3kjMtmLKgHGu8xLKvdjx8
YdyxOzSYU0n5gr2gSuSm/VZvy6Dkv753SmGtl96YknZVsGMjwJI0vOSEJdRQAg0V
eGm1VzAZw5F0vUhn+gsxe9WxLUUQMitleQF8774BTHdHp8j3CvumjTY4bX3LpKbn
B4ltI1rryzd4JzaekqESU8SBteM9NBcYdn2FnAAWf5cU3Ix1p6/jC3zwVKMbZ9jw
54/9i94jToFXpJVtswwHJsni9EUpPFM8cmba/1hNDLjI6x8x+UKJfZzXUvGLWnKm
yJD30skvMY+ut8rbUpYCAGdJkxizQlbF1bPz0uw1n2htRuiifjgsGyN+yFAmADRU
9L30Y9qR+8yKXfHCFoYT8PLE3yb2gRFEJcRw47Wd2+CAUkq3hHJMpBCoL86Abidx
5WA7FSpNrgay+vIveM2bIuE/EyX3uVHisgCHYYiqNZO2Pap2/uNxcyqisQ4kVBkT
w4vY1MUExlBzIsBXbBlkE0XnYuYluFx08DHLt6UnHGGebXGt5bEVsKaxFMDwBbK2
0V5OM6HkGKMJxWhVRbTAAWTd74GQRL7KLkYDF0kzArw4vzwnYeB99SGMFFLvFK4f
Fe32R45IVnVMtbFr5+V6m8OtTIoaRrqg/lwivjumQefEzJH0lU3EyUAT2xVHrazj
BjP1WjqJso2FSn41ReOZmhkifd6jW2BAbYmvaRP2q8akLYopfqyHXWwN2wgZzHwp
w01ToyUy31v5LGFxhfINr2V72MCzXVPnwX/h120tswcs8CxGx41AMBSUgdg1Y7nb
4qdtQrFet8b7NhAOW28XWQOWKZVVqqVzH9fmTGNtshNJmJNS+5u33NvDqi5+BcQ/
BFLkZKVs/KamPk1X5gfc5D/VG69Yeo0DEIqwKdd7nztVqhkQMjmRMBf8pI27y3xe
pGZX3PbgTJaF09xHddk0GV9urBTQv08zi4jtQLtZ0U2IiCECNxO246F+gqNnZLDM
PsInft7IOsqsWDbClWhMQwx7voR/qWz0gWrbwG5pBIjyno5afYU4EVo/oKzrm5qQ
3t/5GceoWV3ELZyOHM50Xk7KqHHYvDezNjsB4HFX1JFc+Z/4G6VYXMdT3eIEJUOk
daJmn3GuYxIkIiiOZihSUnb4iAa+vnicPUa/9duE8RSZvm9w0Uz2U1BNdUBjdYh7
2kmDZqRZKfq3vW83n9XWwSIfA5naR60hqmMTjlzbW/gkOuWblnSLl2KZZd/+VM89
CLCYouPTtXozdem6LEm9sC84Z+GJIJO+9vMV52j6njcTJgR3qC52aB4xcN4YHvBb
rfgq0qLw0R/lAyanSw952dq741AjGo4M9XSqow4cgjAU1v0vlAU/XrJx1EngK5dz
UUtHS4/ZY/Pe4DKO/zmY41B+XTFerpY1Z+Cfq+VWHKlCKI1rx5R2uU6RbNIp92CT
fg32e0lKJGroj+pEPFukNbLIVSTdhjCCGmW54X8D13dJtbb5zDK+7Tg1thm+UE7I
7mWuEY7/AJqrjcFz69gSRMtMy2dQwJYBVrcVz+EMQeen6y0j3ZzwTFjI/SaxWeG9
jL+rqjZvF1zMfBgEu5E78INDpFIfCDWkgkfNL7kimFEc6A2q0xRmlywqhiDxvlI4
oArrBQh7XDKGR7zccPs+v3TFSVXg+Bq5x7tyNT7U+WJtw6bZgW8XfS7RIonV4lYV
VZhLhrd7nLZQTGLg+3HYItWAQkO+JI4kOe4GraklPJeRiEhQJzk+pWoh8HEse4UQ
n0NNwpP6Nl/MynmeZhnHWiAPZS0Tj6MKr8W9YFMBIDUbN6vpzxL1aaTeDm1reH7i
B+MbAimebU00/gvtBV3/0clBUXEl33Utt1jCNlcV67As4aSnSJj9GhHiu8aZXo7h
KSxsS1qMR0zuXpGsM9bctCJKssJlmbjSveJzNC710C+3l/ISjiRn/QYtZQGyL4FN
MgcaJ3ZOC/DNI1wvI+nDomKuLHFVAS0a28YT4Q0JYCuhjIAglrQlvMh4Vh+7wCqr
SJ+wRXSjy2Lfz3D8i1wEMp/C5Nf+N1ogGPvjE4VIxKTX3EZrgQVky+pqFvW31srs
opjsFvutexkh17ElCudtsU+D4jong/GiW5hjKTAgw9IMxtGOzjCAQH9qeTKKDmKb
+HIcRJUzbbf0dskZZcoEpkdywVxUwOQShi7fnx4Nb1qt0Gfot2+ojrFxttKAMu2F
OYo72/SJvhlL7Gb84mSWcWZpBTL+yCAUazgbYflD086s4UmCzpMsiD4CJn3dYlUh
tlku8G+OyAzCiNrOCR8IC9edb7qX9suNrfJNnWQqZjaZCCVYmUeIrdKrtIpmDK7d
2YekdwszpndS6h++IErsM5m3k7seSUmew834eADKembRy8SvAonU0GxmAQLBMYeT
om33HX5jHj8HJiD/AGW2yhYCzciy8Vx8CqOoxBMnvOzGVoJ+TA94h8t/TD5Q5G4L
vI67XcmkvwJDRL1CQWSVlMyS3lUoaAwZmGIxCD5l1fDbLVsfws13vsxIRdyYzQxJ
WoKxdlVzoAc31hy62v4O3Lb0vVpL8pbO+FsGAm7jFpU6gn8R6Z+JFlJm/a8sQboM
0zSBVRAbGP+mXysWtqeBo1jqjT1RBQ0ioofc/W1WXmZvHjcVZKbbI0XwuFITf5M+
mIkKMmmc+fxmx+4Evq/p04DCmsqQO1x/FFj7YyAdXTiZScGwjVrCaxkEJEi7lTMf
YUwns5oW+zl1mL5Qr8tS4fyxiP2sRk2zV+JjOJd2ihCsIoNArrd15U9h/wu3fFQe
8dEQGmJ0CT1UBXIDqKq+w4rpz05XQcq+CoQyFHLSFK91h73t4XjRXBaMq+gRoPxn
DpkwVsI0ThVZu9RwjnHyofPgkQj4GhpXQ5vsX6mTk14f4KDOZQJi9KMLhFAIBjeZ
szd5Tk3JZh1fFqq+2LK5gZHRteEOIHr577M+gwrKzOgPzF4ZTgVEtYz1s03CvSQo
Kulbetx0SKxY0VPsoz8D0Mc4SshI076G3eg2cz+BVI3GzjxQ3fkAPQpZlFJ6yZ1D
wmMsmfP5dwC7e6f4QBouolwfJchW1pYesIAgLxbHf6rXFpNhgnTvKJueoUIk9JSO
weDpgciyiz5By+7gXaby5UyDx0l9ocUJ94re0R9Buh1DrV4DyuU0E2dbbW40NYyU
O//YSW0znNov8OFYmiLnaAC6oaE/NU9TjbHzSsgDvJdRKk6+ZXGA9OIXVGh0MJ2o
/gK030U4Do4J78gJtLhP3duaddy8lVwyMg2SxCqvl26uwYocEvoBznQBe5HDQpgQ
vvIBKMrKMhEz+9pKVfvzBLkeFtgXtLnJFU0d1ZWcGvVys15UwLdo1VifKVuWxevo
3yyPJtfZn9DZTWpNq7bm/mJAQW/OOKX4j490bOs526xGO8EDyzs5A1R9lU2bvcUy
fHBJGIHE5SUZbIIUW+AVncWZLx2UcaVV3/FIdelB2MelAZrh9bZ+55e2GFBFyz+o
nJz9c35on0hptD/NlHm3RdoRWRYJg+Ig/zWyOE4IurFYLKsHYzh8PMvHrwqCh5sG
KLvcaCtIX4CZlYhCxl4pYt7YgIDYquDnRSQfHiuFZuIgzGK7WKWNvxyJfEjLNi0L
Z/4St5yuG/dQnjSHR5JnN8uZNImzS+ebt46F6jj4WLaBjoE9PzDc5WFjfMzOqS7G
u77ity0mzIgeYF/3IuP/ljPaE1ZdltO0KAR3XJXezOH8xxcd8cYjmBIcDyj8Scgo
KR6r8IinwBGf+VJsHyaOnNJV8zCkDGC5LqhZM6Q9HcyfjznkY0paUJJKKOe8LYE+
X0sA/nxlI+cnx/Fk8SWOrITwntmfMRrmmQLDDBQeWsS/PtvGoOZv/Y/OpVnSjGEV
SSoGW1BqI0XUJkyjw/kQ9bJSUYb67VTzsMvfJBuBX1Od8YvLP56+0J1BVFbEP+Tu
6w3znqc0wLkpEPmna5xwEkzFhSXR6ar10p5wnBM3dJs3QgRbGtGzb/Ufu3wPKGod
6k5DgwNp3PvCJMDjcH0yENZ+0ec66DW66+Qwrl0HhljRUcjZjGV7M8tFvtnk6uxA
VRjwIHTf9kBQ6RoT0gfn13pr/js7JWw9DaEDSYLVDxnc3PG2jE/D6ucnR9WHIFkz
GhU0l0kZaZdsWRvdKkGOHzZO6qMcCNbwPFCY90poDgJGwYiLIV2+NGVaiqc+E36f
k8wIAb6vzi8L/Sgv9dU2ulo4uDRzboYFgiYwRvcd6Bvv5Vc1KXYMU8vhgNmLesRI
qb1If0vXWomYeg6b+O3lJtmHsNctb2R/PlJfQeCwXNvOTj6N1mIpUl4KmqgLfU3A
C/glsixUNCQv4lio3gBqyWPYP220huGZ4TuVL9HfETP3e6k+CAATW9/fDVOJsoqZ
0sjh6g3sElRrpfk4O+Lvyc4JOtPQB2RBuTxR1ewrWaqcAwHdefDSoP0v8ZQZsRb7
AEEVxLy8Itg1EdvNShEfBhB2Af7w+HGq5aPHKfn8kO4I/Y2SKVPwQ3LOyZk8lH7L
sfs3OxiA31r3lg4hfQ/KRfRAk8rHdcf3gimHTUqfAIjjBg2iVqBgqtckM+PvWJPD
PEGOEOjf4dq65h686revC9OD4DGkZd6/Hf/jQiq248+hMsFMh1jpqlqNRYxI57Tc
hLNaaEw46jh3A8jw4l0I2fkPZ7sFqyNeeb9aqwvQ0uXF//Xck9t4dPYnQQ7jh4mq
gFGWVy9dYEs/fE07SmQ9mcGDdXPuhKkhw/zUJFUbx/E4vRFljjJrh6GvNxt5cKN4
+lZigrEY7Eq6yOg1Tlva8Quk0eHO7C1KE8ds0d3BgJciSsBOTId20g6glJyAUV61
5pUCK0PyD1LfQH5xJRSZ1E9DjmZe3vDVP3L+fbdNA8Yg9XTNjIsrhLIUH6sfWzHS
Dytyh12Cars1ryXa3tk7VNY8MbWM0i1p+rcE4VYrLc+Y2lXCxVFjjXNQl5/bEijQ
lTxfMX/UQbIpeJDvMrIEpwTrKLldbL01f5wtGOejjWASOWSmOzxpatGOJyQ4gsk6
zLbWB5MqJRmbcjacQ846ZhaeXLettRfx4UVcCx84OTMyLhE1NxkpOG0x+TlmLO2K
PsMomRgICTQvBo8nWcsuuvDLETyXTg8YWS6iR9Ri6GKC0BYLKQKyWas20a86UvDe
Mt/Az/MQHnr0yg4vhvNh622eVCx6ym9qCyujAIYuZgncMfZGuLURQmfkvNAo3iev
8u/k4vupe7rtLAXnx/IY9R3EzjWnFgIAgt65LLnnLeNnWi25yE8rjKfC5DYKU2bA
jYu6vyiKqIM4V/20ZRxBi7B+MmjmZ+6LdQhC1zG8tpgt0SiHppxSRuygkkMnZ8Z6
ddbODdkc0MrAGWYD6LHOAOC9nz/HCXko6s9JjjzZE+rV7Pt6YRO8eCmTLNlg1LIb
M5RzH/DoY0xkTq3R1X4ONR8wp1Ta40Gx0m+N5GhlqI4rvFMkV87zPByh4+f9xmtr
gfadD67o6cWDG9ujsnWo2Fhzc5luK/hrfIZdl+lTeikbjsraPeQPyZJYOtmdgTz7
kMgrQY8i21buiG1I4gEiX/amW0I/U0J1OiR9pQ+TORhHuXKb+vg/po95C1mtoVKq
S3gQdOtu6tPo/zDZPq822bGcHdiaW6NZjU9rv3yAfd42CiBZHaL0wOm1YzDIdizx
9/EA2FzOwAD4TzqTgHTGAi2IEa4bdDBi8LM0SStx4AK1bIqBfjs+fzFFQCVM7klQ
Fp+655/R39WmW37mfWiAePp1OsoXfEU/JfveonffrownFaQPTfJ1ZIDhyqyf/5ZE
qxkoj3xoHAXfw1gErm7h2HoXYcsgv2FVmTCnA4NNRTA3IdH8XXN1qzlYYHnPCkDD
Q1C0Gca7VV0PhdbjZmB3TTaq4FdwFe7oWUU+arwz6HMDdKdWsEHD2hAJ8Tys0NGw
sXDSZF/O+awtvPmiNazFkRu6jRQ9RorSq82dxpSfr8am7UMvkqtlc2mGGtwSsBbW
za4czTEY5PMjNh7CDoVLMjPIPDh2HuBE+leARy7EP/aSlma9WjVuKtjDK6X+UBJt
8plnZJLZJAdRwCwAenEnapHVEbj2NQQwEAA2qnpsjS5UKQ2mB3LZNUFbA0xgPEZh
4DSCLbzfbTnq5tremohdS+qTg9vM0b4WvrQLA3hOOQJ3ivRMgrCctP6XfHpZ6wOF
BCLqDNSBL30hjYfnL/CEssf1n6umTWukOCQITJQB4s0PG3zspjvxJzUfqbKOG2Rj
V4CW5LmSDzM8RVeKfmiiCaPfSEDcEDrH4rD3fMsjNNoU8PjNM4WrdEmIq7BiZn+i
nlgbI5hjXqbUN4ttSpC4sRhD5ntGMkuT+UnUWmLF/lHMZVGvWq/jcjabMRBJ48sc
Vod4QBA/EN+cRMiV6Ni0y6CoKzcL3PV2fllcprbs50FESNSFP/6xJhxCYlKf1quz
eJ6cZ7MuPxubp1BkmC3NQKmm1e9CXR7RQeHen3tJXRaMYExkAD21GmLjKP+foleJ
gHsS3RkDI9BYyxJmvG9nvuMzgxdttUKSAY4RPs3xCQFR/XqxW5ZlFim9qH5MPAeu
YGb/4BUVQEIlunkronpCRg8S4eQ72LiAACEEYO3IYPh1NhTA3/3DsMBeFXwrGsLg
RCnBo9zrwWpCI2cy5N21aaMRYszuJa9A83A0cx8mkS6nGWPQv0nScc2WXXK5Zfhr
jzHQu7ToQXjAN8gJtCP5+a6qgpduw/47aV2oBBw1sUekvpyJiTZC+RW0Gp23p3f3
N5HITnNETOKackwMgZn5ZLhe8x8VMWaFzE7kyU1+a1mJaxTucL5AAN+mLg94gdcE
OHsuywyg7gWhmc7im2QXAEYYYljdiz3Y49QQOLWKWRLdpimSaqCKeNHYoTxapdzI
ciCopKnIu+5aXLFpLALd9I+3vqpr7LrQxsuCpk3F5OxDhSyN7EUWjDQH6DcnUR9i
sxseiCr3Z/8g/jEHeAEktrK5tDbPoP5zseFib1m9ZfcbYGMI4AFr9jC+99hLNNQZ
lIVpYo0cYfTKg/r5yZNSxmDS4Q4UikV2gxhrxCKLg0pdUmo/H2ausmDCyvgB4cT0
EQ/tEiE7p+hrArEYV9LrZpa8FvDFz5U5l8U8OclKGv7g+yXSlo5fQTSk6RaEaEoI
PEI5Ce2U8GiJT3vXM8FxGVXBVGmiohh0qOlV8hjiujm8/RJFdZD6C8t5V1kVBNVS
mNRXJ/bmboO4U3K6iaxgH3lcR76Wo+fa/CbILuhTIP6SWj41X/wRAhLfJ5kEvzor
w2o0BtgIJqTh7sKUhCuO/GtBQhZefavPB4LGZ+Qjw5y03gALuwMTFjowvnraF2f1
chz05TIRxFNxdBEPuwQ/waNrwDwG+7LRaAdFL/krKd4ep+gyzGOYdBRchS9r4XOQ
GXaxOJ1/daI9gA42Q0PLsbZRcWqTkUN3Hega0X8O4WrE3THGPxX3MZVLjpl1qdf9
ckFBNSV4O/FBWh44katDZf4eKU9ui4ZaNZfqdcvd2qtNd3rUDdq6iaytD/ihBt5h
fK7sNY4rR95uZaD0AIsRdvgZRKXXkiz69egy55kVMIjr7K7r4cLDLj3iQiV5dvWA
fRx4DJfH/0dKa7p/fEPslkg6hUUjcuDdswYgBiW5j3ZDZUBPAartwzntsoVOGwzz
2zebYk/CHIt0ngrDgIzS7rt/3FN2S230CWqJcmODNfG9hJ4D0KmU3XoO8COL5lza
qvJTeT+9MQ03ia7aZdTzZP2/JzXNm9NLW8o0PDfmqPkvdf56BsyiTKIZDmZvQCbs
uAEh7QqLuTvficLtzgxZIc6qru+DhUr4G/Knv8DYTf5FXklh9GHHN/TwrQHILVlo
WHmK6SVF1vKxVSVDmBIx8cWO7dlRDbgI6mTMu7MBRH7pVqRgW50OVAzQTFoLVlQ8
JDclLog+EMYAbo8QTRVSGD1loLTIobeIqxoB/K3+z8XaRS+8qIX92FGotGosqb6Z
pVyHVfwV22EnX3wlo9/5SmMWY4s6flvg0GLT1ltqPoB61SRttJr+tqbeOq4OCxjd
PeXl820IHs7H63WRjdzMdF/NMJocyCWPOl14fBSUG02OKJC32nzO7k7QzzVtTmwW
1q3GhY+yMs10pUCyqExR9RlJ5Ggw2er7nnfcS32NCK4INNJqfieLNf7twrm0zmEG
XjzW39bGjr9yv7FEAt3nI7KQ3Tbn/zbOR5SHzp9MlXXfuwbHJkkFEClo+RDfvs6/
eCCarahs8wqWsn6X4SXZXO45wMLK8JBoBAMXIkggoOadMey8T4p552ufm3oKFqoH
3JGzLtSVHcg3rhWPj9fIp2s+L9keMvhlTtkoV7/Igahi3aHavzvGMyMiSr7b4a0n
+SJnjF3Lw3Peg48EoXD4sfXTqNomiNaOr24c0ZRXPaMFTK90qtE5H3Pl/V8gQKZ2
Gc/MlUhQwg7rMDXa2cp23jN3ehuLFKub2t8zlu+E6qhzKkvQ8e570mVpPPXQTcsC
yooREpSJ16xsJIKvgR8WMVcFYpd/jkI1W1RV9Rwqmc3cU/Jxz00MnO4s3A3iDQaK
yhkNnbNfagXFFwvhICDsQpF5qqUujnpqbF1+jjtUhNQBiBpybVN4CR35MBDeYMng
rAHhjRwaMCUnwemN+k7qgqkiEX3nZS3wdZ+MBJv8dJrsJNz8c4NnUvIssN0W3h9a
QYzAiFH9BaCom9mDNB4W7vwNLocULNDT0qAYbEYDZiYcND/dyIO+ZO4w8tRbsQV+
WDJKikEE71Qwq3AgUQO+emRJpyfBJk6D5vPuKOs1vg/hYB/6sjGa7+4tAGjafXeP
LlDaSJEYvfKOU+gP3AgqV4JkBnxnrN+hqfDlJNIX5tjYGroM4EaRWgpuLW4pp2kr
1RuGP3kIXpv9Zm83lUpolxU7+CMwUvCqFS7JbjCbA3xEPvvd68yUyoAPsqC2pt31
NV5xs7FgdWrb6LpLzTtJzkTH+2oZr1Pwu6dj3CroyfpPQPvzHjqjG7NtSumiZSFS
XqM/AZ1SGzz/IywkokxX8KrS9/df64w45Nud4UVrNB/e9S919FZMc7XwzQCzzhdJ
lkUIzT9bRXB/bIxcGeaQaWFQ7oHdetmOZps6hUtXlzTUIkc1hYOO2expX5b6B9Cg
uNR1pwJIgIcE/y6F7fNsYv3ZNkcSg6QaoP5c8ZEYmpK8Y+4QAoKXoshjs8CNDmYV
xdlqFd6Jco6/alVo6t61Ee26y7lvPiyh7TcG+36EuSR9ClKuvY1JLuyVDumEEMSG
m1SIjLonHmLruHftvPagT+Vqr2eEwZkw9w4eACmwfxctmzlORlkRICpXWJBEZwpB
5IQV5Vzg4hDgSTC7gVLixQ1vAQpagzSH8aHzX20o0a8tdTwGbc0Nl28aj8gP/s/8
EduhU0D/WsPLTUn66xwDxNsBSZAKItf4PJcLjoUZpqOsCwqpEZeawP7Ckqs7zFuN
lwBFrva45hRx4+sAKGm4SObJRzmScL0+Qq6F2M1brn6BPsgIecJ4qcKj29NgeyEm
W23mgZ/cDBGM6pbVVhAT7PE50JlqqAv1ARheLXPCr9I1TfAtNnZ/RWrvBposVc/u
fx9w7GICWxls0aYyiT1L4dmErzTBmRcjNynwvQ98hQRIoGvwqo501E0FlPrSSseo
2YOW/Whcchgd5DLeA4Ox+KCAlU+izOEJEWFz68mg7FhQ3+dYJLL2wLmkCmsFy2gC
XyozVLBVtEL0GRYHWWp7LEUcWliMPAAUUtqE9mOQgr3azYb9wxRovXIhC9CFOYab
JkYvtOPK6yDJxuvuxzWfjfA1hZSuR5wm2/zhV3OwU5P6JiiR3c8vwBL3KZUb8e52
OD2KSBogMayyQD+wpQgwpMo/O3XprNyxLpZRs0aOSFndPkV21AaTy5lhcQ+8IUvm
QfDUh/0KTbySiRglauOfKUmgnTitkRohCuWmaJLrjAK7vVSlAR9k28+/9b1Jh1xp
Nn3/bj9q6DxmMbwNkbDpV1dmQewPQFAV4lY1UNwJ/oJPobgFzztOGhP0fs/K+ZjI
uyIMRJb4OTL3KOeTLlulYvPNU8MOxy529XbrMJW6o89zplO7BpaWTp/s4LpZM6X0
3dnTG3MlUVSiIR6gRcDSGZ4eukVAPel/jE0TTFYbsPHavvbWWnhvJQSbYlBlzO5P
yr8hCmv9jTO2Q2G91hDJCRnGh09ErvgWlm19kNVSxfeg1aFpLbhx8j1LyciRKPvw
rD6GRB6ZZQDw/x0JnuhjyGyX0z8ky89CeOgM25vsOZgI84Ub55l7X8rKe6c0XbYW
rn/J9Wv5tWZ5SFNJM5vjhlCOH95c6LYpLtiBGQ+W1OfR6g7SdZrPfQsiixAZFMYY
VXO6OX9FngQUZEGTGuA13PPcaPEt0bF4K9aoH/c/ub65oLPOEe0JxdOY20ajN5Nk
ErKh2+OTCAWN2i87Cw57emDglFyHZ9AQYfdiIaZgN90BJ6mz4pi2+BefY1BN2D6K
8vxPuPmRtQ6eRyEptQYEmq6VqlCqssdbMQNdBuGr3CI/P94lNS2KNg0tN4TULnFx
AmV1viqYHcC5+ruZO3cyeVp++584rwo21AufmPlaqfdG3MNjfmKjMsX25cFpg7OD
Hch+N3N2yi6BFTKeLWwG8H4AMXdxOB0k8IKFf31wHFi99vysKqR/x2Ajp2FUVAl2
i82MK2G/WgBL8Prd6UPlqVWlM9a4kRIwrUQ0D+ayzWL4YzlQNkhYmIQuMrJsXFdv
MAfiDzVbbloHjCxVM0sqJR4ib0cQoez/Ln2e7yIhkmGrHNSNjTr4nTrMicKAFB9Q
bJgLNDovrUkMqr8hHWxMddhalIhkBNlrlavUIxy5EqRdYvgAL1iMl8gIlwJbwi+I
dxB+sUGVGD2+1c3BCkgjwuDO6yylOC7jqJ2qibxWf4RgRmACN8LnGqG/24nS3TVD
B1IIPYtawwrOiXNaLVjgoVhuuYo2gQxr7sO/r62jc/pbY6aaI9uBQ3GcjP0L9bAk
M4zGWBotezC0MlzaAO7v6yZcYalu+HGWQ5+8LKK5ebwlY+l3Cny+cYIBjMnfZB9t
XfaAaQpf6M/E86VkVIGnX59OAGJrPu0/iG6TYV8fp+jIiyIOUiBRnn9cHhJCCcQV
GLBTUpozokUzQB4yOVwxxw1mFuiagDXTF4HafARqIp0goxceYwpN59QjNdkko6Je
CvmKWfZtJyX4g5TH38lVrvhgG0iPIhFD0L7cnSp5m1Pf68yvZGCHrAMTN1Hv2XPq
Gb3p8KEC82q0JvD6VUV9yQQWt33ilXNxKEm6xxmTpC0+GLiiN4GO7vf/675Myu37
PHsjI4JFDFgh3bby1eT8mOLk/smODEMl1vk37VW8r9ZC21Z2SDsiG5EyWh5IL24N
TvIn8AiZNcaoQooz/qZnLXkSdbyII0Pzul8SwnT73TU8DiJBoCEPBHLf7wIzfTEE
eTRBCvy9RMV0YKFalOQNTvQcCdqcn5vCR4HfslpSE1X5HORa0ArZvDyqh9NFapqF
sMqVQLnYWHx8u8170oH5glbPD3RL4Ac1baBSykV231F36S5dEgjwQJ8nVF2OV9Df
Ykl8JNp69G8geB8qBMk3hLFruhuntXjMDR4BQspOQkX15uEbXSUvrv2Rz7i4929f
xyaB5SUgjeOZUMOw/9Z2DYW7oaknWXnvbpMOhuxkmR/bwUL6ZmeGUCWh8e0PqqRT
MKfURJ/cEKKkOZQfCazUhOc6hxDdNfRsZVfnpuCwyTH3WviyvZzfYWNN+w/2pSQA
noM8l3TVc71ZgZue0l50bi2I9Mk8F+0crQV465AytdLsY/d8i7jX3+tYD4uRdXYq
bemY7LYD50F09GHJNPTwRIWmISdGArY/6hEZzUgWatOnHtHZ8N63VP1/Cn1H6m53
+4yk7CNqFaNpsEDC4Nctyx/sXv2XaFYdrlr2r2EJyQ89XUONwqRLjc00uQZvCbzG
FX/A9coHO328rRYblxUcr5rm7KphpDWsLkClhDHT3zFbSC/y8LbohgweozZCz8OM
i492CUB89xyD7rCY0jBgDOg+ExgtfMFYIQL67KyaLhoXY4gzw5Jj8MR/C618MX8X
D6ONp8lx4XGIa1ie9HI1yQgXz2xaV43pjBhfb/ql3rZjPVGboBrVBcysZI28Y5XH
xvK9xr6iLIHyA4d6iIrJFXZbcuuqSgPdBNKsp9lijvEUUdhnTBEq1rYCnd1SHSr4
S0oSXDax3mvs2DNtm5tyF8Xcrj8NFSlpR2qy1VYbjUuQLFKOqyTE192sjWVFlPAT
V9IedEJKdKraYLWu+rQfTqCBJxn5ao0tg7g+BpwTQzezdFrJ4Vz3htWFp5i5FF9a
AnIycQBzufGNt5klnXLbd69gSwHYpXZtARYumG7Vc2hlgjiZr6hA2QxUQRUh692L
KsH/0PZny4jOV3L5CnFnJPBoITfIHPv4KyBrFjkzPAGTsMJBqNxWSL5AUxytcRFL
mAeHLXuYlA68IVwxF9GjICVawAoz8mOMlShBPIjOHppgr1o0OJ2CBerSIeVr4lqT
bisVL1Q1IoCs5USZS4t7qIz99jg/elI6waQ6jTLylvknFqU18+VbJVtyvpaXmq+8
aFxxE0PpvCVG6hfVEGCjASqqQEdtt9cpbIj9CVjcyg3oB+NgKZOohGhOfRMpLUdp
EoP5laNjCP1y/sBGb8EK5apmNjKtACbJB+dTZPsaHHDNzuJmKs+RtOo33EQP01X/
hLU2O9tNCtgvYHRr0KF6d/+B1TE2YRjLyWhJAY4WDQ+ECjG5bbTjL6WNiIL3oaJW
SarCpTjN3JNiYte4F12D7TDFMEEVBG+dK3LxGicNLm95XpzvLjwiwb6CRgi6jUJp
WL6GsnABl6P3WadntjpEUZT0u1sCClrJ5dGKZTULsaVmoiuRuqPogT1hue6RP+Bx
S3iPU43aimjivWDElyiZCD1Uxna2qD0J6vsUvBPtx0XyhZ245AnTJRiYsOjOAbTd
QQUgxXYdM33QWqvYNm6xhYrtOlG7xkuy5/uvk4BYtHq/t5mFt9CHVriFhooueL/s
SYGf5g4lr9M7bsDHWw1H6yp9bIKItErh+2cHbEQHXdsL/FoSXHkq+NIQrvEl+Bq3
1bZHesQkA0Gp6ZuInZgsmK2wby8ss2bycEzigJ34NZJtO8ZKKjuQvxRAdWmgtmcB
3C0eGJpd7g49dUhlE9qhc3a5BMANUj0yoVGWDtQUUJgLgY42NdXbJrT53AIXx8FQ
J3tt2LbRizhEwmZlh/rvoUVQhg60ZHbE+r/s+LCmKQCDfYHzRkDKzLkxPpUQR3Xz
PZEbBPtLUuEyEY8L0wo8zuQIBTi3pzcoq7CDaQgEr0YV+vDzXn7qb0/ghsyecnHx
r8fvHcwXjp2QlGVxzRIcMYc2paJKdXXZslZ/AQlOjqg7WJHO6F4IPEWepcXGG/gy
eYwPFGQDfUfLDL3RY94vRgfYV9TsNKZwOmRe1+uldJyhuTxMCzv3xy8s2Io4qI9A
3OZoyboe9/5qLpRIUdilJs7l5rbhpyVhxNTJABviM0R/OpRoomsKdLQ1iHeC85iq
XeSOPAC3VSRdqZ8gnhxSByhJdqwlphs5vobsWsQL+V0iFUCIbu7ITN+pnRlylN9y
1UdAJhWag1LkxMavrSX1Qby+w4/Dj0O9VKcHTCA6LnBHicy+gXx/KpiZiCzXBgoT
xBTt7eS+nhEpGyxe1LheB1I/7Q1HAkZwcHrey4Vwvg/V0pLuPLucFXxOG+ucHU9j
ZF0rkObqfjEGjQDWX6RTk8xmVB2koBaBDU7/P1G9FvKkDbcX8LiKcIh+10354oGw
FHcTjtWD+UlLfKyFrvlpNn+Y7OAP/DDUiXdvRTBhCvm5WVqkvgpItDfVm7IXSpO8
2AzUBdURwg1o1lzJnhD0vNABDtm/y90Oy6HSdse64FjTcI112sfGnt8CB59GxtaY
szlPMuAjj58ak87j/S2pZ7IGihPkeL6IcYWwrK6BIKKbxgls/EjVzwcoLz5fxyb2
I3jinJ2LQ50SVxPWqODA5tCygoj1V1jcSB15KuRAVN33FP04rAcwdW7ojQlUqtbt
t627LccEq7NQVr9WgorJMdaUJS668QaQjBrVt/OzMK4N48juLeRCWSUZmTnmbxO9
C5cwkBvETPkDodlW4B2xKrSOZzOUQHwE7FrZ5jSYDG5MbnWgoOCBY2Cv7DQmjHQj
NIGlJBtUi0p4dNxRu6McDABV8OZiFTXK/YhGwTtBhzXUjIOVh3Vfpe+tGpPr5I5z
vwSVWPtMPdXlsyvGjD/pU7RFw00NRFCV5sIEr5+/k/Gi9U+L/H4ofzTMdHMs22g3
CVZaT+eFjsLJJZvGP2Syo1y4qs4GlORqH37WAFatlVm7l4wpfQ27fIxJPxOQiJWJ
OOctIfaPoz+rU4EMlZHf6pXeFp8NMHEQCvJPO4I/W2TDJsjuQOInMYTRa7rww0l1
IMnacRGqeN97xNJRjsa1/8Un1Kq3Omr7V5iBUMhMzr+U1lpx3LjEur66sLGzRxGK
MKO7lXCKXfEnxFYhtjGvFTMCpeX5AKpph86JxB836PBr0RImLDJlIo8oj6Ky5+lp
h+wq5e+QpSA9R3CqoF/QqDNoM4xLNDO07yPjZgpV/ZQ8PQ/2eAhWtxVgwBzRlS7M
rdA4PAYi0rZEVB0EnKQu5669G7bLbcQ6csnEwBddYIP5u87ZUDkpWo+0wMq5TGM0
vWVu5k5SAHmygW1QtH2DricE36ABYmtW3266FRffKNa9iiV+MCNlSBcXAjRQUju9
JrrOenIzitV2wQUh7QCEQJpqfGMsXMqqfLnBMFoabDMLPiKESCJRLfcy1CLBvW2G
xSqjG3EaOwXa68LNB5RaFTKDtoiAylGf4wborPz21/my9W//Q/znwHxe1vavrCg3
HboGlWjTPKPq0G1co3rjCXLPYhnDc5M3PDoQ1I0YMzVmiYbJq7sa4z0asKKEp/+/
iC8arpWNJozsgSRVzZpvhOhaAbSk0XMTpRtRNWuN/JOj0jy7+avp8GBHDisIU/cC
7qNr6IOE+ivhg3+UAkAAFyoCnbao8xoBj8YZ38mJ2TMD8ynL3+OYCu4oGt4zlXrM
lV9hR3nrI355YYMfK8jCySLTMN1MyaB/3XzsikI8o0fwL7ZdWatbkMGS6VZh8G8W
k2KWN81GfMkB6JZidZzqsOXfgLXb7fNBlKTY5xIG2aUNgLc+XCS7HtFJl8+gcUdd
XZvPsG9svEON2J2ByIp9khfuO52YNqnnYSIDtGDjMRfKxCQ/9WYk+tpREIgH+F/0
Pj3YjG30Z5ypKtpEgrtzGAnwe/MNx3Nmrc2CsUPUOo4zdzjqRCnLjk36x7pnhVc4
OXykmBrqf16JDILFlMKgCSypaBOHhx89xWScnw7eOMQwz2vj4wspw53xrg7Tjb0u
dbdFgVrzOUKRKcJtnr8zPYVUhgAliooNy5eFZjwQpjgHGEJUF97RgTSc+Q/+5jVY
TdF9C2vMEOwcoBUlRsnxJ8mSDdQAVv6mEJ378JKoOhHXzqJGzdcalFjo+cgxCBoU
UzmO8SLYLtT7phjqs9sx3eeelg4yyHDe7rJw24z8VQXR9rUiZAiVh/PU9F/mPxvs
ZdnKvlKpNsxenbfFBAER9vyJFoGZ2eIiTdz2zuD3xre8eK/hvQD2YgOd9jKI1EAd
nVc6aK95J3xwh9SDssmyyB2bBhb5yr1oJBBsawIbE/DyBk0zdkbpY5Du2bF7uOOn
2fexoc+AeH3TiKsf4S3xnuEkUTyLSr4osN8/CuSFonPw8U1hJIg3XBEaixlbHvRc
2EJl2PGxHTjPa3pYj/odU5n5CgwaCcPFdwsaWp9xZHqp1Q3oYbLjVZL49+faXps7
hZ/Im2rByUnVEPbLnfhxAzLTbAqeIFRdeWeSOVg6f4AINOA4BNS2UTZDWBDuYouU
F65rspog2wy6/XN1hhyVTaiiCVIg6L0P/F82co3Hp2SmZKRZ2aXCzydC4ijKW+ok
NtXH/nrMHJ9Yb1MWSDUbsLhc6h/hSTeRfkZhtE0zO7zXj6qcNtnRmEZ4VWr5oJHL
qGK6r7X3EAyuCflzBR4VcRL/Wb5GGLNRvEMeTUtWwmjMung7e/D7F/Tp4v3ZgIhQ
fqh1CJfgFGS2vcYRGcGIl429+JdaK5KR4dtuJrdEvaBtWPATw9TVaUuvVxz+Fp4Z
9K/fqDwX3Fn4Xc8rVP2fkuMnXuaHoQJfVWb2+h0KX3+V7LxjQ/Xr69pLTWRvtuuj
q5gnw6YOFXffGDmZg/B+jI6+yNQfltZye1JV8Wg1IurtET/tPFPhmEVGEbEXieLS
/pnHyvuWsVu+8COazI91ljTzsJM7v+d7WcKO9M5GwNRhE0eSrce4Ch9gSY34LHFq
mrjgOMUmdTaiOiMq8pBJQqqB3pwJzR220JHs2ExaPFhtlHSbBdf1V3M+0Em4K3hN
k8+9Ec/QVtdF3UmFknItt8CpKmavZ2oRGjCe0HEh2MU4sSQhVghnemIYnLsTa65L
b2MqOX3dMoQ0bdWIs7GlJb0pAO3s7/xhguxsx6yit4K8QLnR+3UQb/9+aClko/1o
/a53JEr3jEuc+Xs0VGPMvSUUiEJ103b2UoVr5PjgO8BVkQUFL/6j9yvedASZ/4hP
UV+3Y2icjbymgJR0if7JsBb5Uj5nQwt9yYLyWbRoIZhDE9u23fLNgemJ4l5hHe7X
fwL0Czb8amB1HUEEeyecW4wjJBoFHFnTniQRWin43NPe++KumCONbsUwTaP3X6Ci
7M4mmjPiGsykVI568NO0zVP3XDQRZ2245JvkejFMKZRFbBMFc919qQDSAVaPI8qJ
H5uxNzgp3QLO5pGc8evQFLmyqJ/q5BdyuMmMxpu1BOqeWEQcuQB3EuaT7aLbHSNK
p4yAmxvN1E3cQuGWvQXMWQkxJNwN9NAUDsvFqOq3WVRqBafqRcJWTssHSHuLl9nJ
lzdx/DHNFnkdX5V0EdP24CDKbgWEhafqHchMPhcdAYC6FOiF99MHM/VLNevGjifO
SdUiMrBjNA1eAKk3i2N9W67kId9QJs9jHLXbLy3y1hjQ8rQIFs9A0UWzc8Uno6As
zOKHmGmdXAg5NyI+3xNno7/gGNPvsOAmu+RYtBwXFKlTlr2g7AguQxTgkzTU97p7
vKG3qFJdaKnyGQv02S8VB5Jby/L5j3BsapoTXFEc98ZooCQ/ULGba4m49TeZXWPk
PMACpm7nr9Ud61dQElhpD8JAaP7CtEIPd1A8aC52C0S8QROvfCcPx6gt4QZL3n7h
wlcltmfPBSsIUjLASathGhfIHHwi905K6n5TqJ/eIrPg1Vb6Q6Ek1A9AqzL0pK5q
S4hFmgC9WNmNJPy0urreOoIezoJ1Vqbx73HbvyaKcMaL2mGzjZaZiHvzSXwqXVOY
7IAqjVNuc4fHwepLtxJ6UXD6Fh/Onh5eT1kjtV87Eh+Dj69xbLXrq5y/WJk+ljEV
JyHX+qj78Fxc/rEAyWpcOXZQ8QqoHCv99T0S6+op/VMcT+1lkea/ZY0HC4L287Fv
EQrNfkJt/y9I5g2Ox4h1pEJKKiKPhG2phqJKMLpdBJZy3sijizzbw9PPCRXByubp
zU6TeKXd8I9Llvgk0Yv5vupWqgRFteAMm6L3sig1iB6xhr3uk7pTEKezub254WvT
FSfzUsF9MDjuhGmmNoY5FhAgn4sPKUX3KcCsxpzSPn/TDUOLdo274kW31UUQJoRl
aarpxHArYddOwwrCiEZa6Z/oRYQAo5YsgW4+oT8qFCoBRGBAd0VHD+hLozIf9Ba9
0Bsqn6QOAOGcVYn74EOk7nUNP1ZW0O7lPxm5Ibjf3BW+Xe4LK7I0XHR8Ht7rNH7u
BBJwsUlB29ttwh+FWfOYYGbKyZg4Ji8Vryop5gX/pjTtKPYG5aJsVVBJCNN079NU
+VoaNA3mes5MF3vRQqrDYgOi6PJ8hcFYQkI5QoxdNT1f7bNldGUHAadKFllVnKML
SDhbqZQmeQicqMFdx1kCJB56AOrjDIxk0zyQJUn0JDnBgX1mGKW49orCZtnvYtoq
XCbOt8dTGtxDgnT4cjL5cIFlIGrg746rYSqomhucA6ThcOXngR3y9kQfBwMdlTRS
oGWOcn1bXrDlmhgTcGVCmMt5q02UULwEGyP/OTLCjMzRiqkYawlJZa+M1+4alOOa
3WPqAhvdH8BR8/CPSrTMWNOHfgKPCJ6oA02my3qHOqoG2dh5O42/ITS0cP8p7BBH
5F0uGy6i4ktcKqrenO2sJejvmVCGfAztQgtAtDWileO4Zif4mMPeb8OzAzWUp/zB
PJK+qa6FLkcWHBp1Y7TvgSdShtA3XYDwySdwPz8uGor9EiefDDDpat58e5Kbtb+e
UyY/h4bh7YeB6QFlucNpl7I9cs7vQ2Gc64yTqVJs4F53Pmb7PIWcWMaFka2yvTUO
wHXEGkijmlG8jZF/f6kL2gZzh8mAKaJ7lD9aTOghek3gEF+Vi3VvCH/NWBfbogbt
x9dcJX5y3SNvIZhTNk8dHOs8kPpgtnbP6k9Hjm9l3WO5kY0CBo0DoVziMyn5pZnA
aOt0U2Gi2QDgfqfiwofCBc1pEPz2Iud+VIPwrSvZ9UsyZbpppucFq0h1js+qE8wv
UddES/fOwfGmD86JeGZFoy8OyMv/VXwW+AjyYUb4R24vVxaavbV5mxLPrpdyjsdS
53Dg7ZAwzN5bY75A2UbO2gyU9C+WWYBDH98oJD4Mt1SKs8FmzGoorVNhbPmTGD3Z
TCK0nh5cI5u5Ao+BabubLBBat2fCZLepIzpoJ7Tf/XzfuDdej6ZzaODN7/LVDc+a
mF0qg5wyC6jkClBMFje2HldK/zHXCZ0wHv2E4jG8eO5ptRQrJj46bl4rOTA+h8k4
bR1c97pAlsjPJxCsYbvkM0EWeTIAm0jTdEPwWoJuVNKcJWSCSOXC7f+j3S+N+Btf
1sErtkOcarVUJLwfZ68etUYEMllvkYC/8fOhlUbFrgYeAkPNhjLdpYgGb+Uph32h
ZTF87vnzSJWPGzZNcDkC327V2k8PEv+EZ5I8+dOyowow735SbX4hHdqacU2SJnkP
hPd1F5rQz4VnAgSJ0DlOGdiAqww+lW3eGhWEWdmS5RMRDqE9RDop5ppqvcCOsjOw
FE8b2b/n1cFEg15XaEDJThC7R7+K9+L6yBAohwLnPxIczy+ZkL/FpPryfKJ56BdP
xf+UNuCd300KzkqewyAN6unQP3rx26HJ0lSJEG5/0Y5HPeWV9Y+2IeZTNIYB8lPA
M0O7saothzLeIsLB4Zzw5NhBBF6RmNSLNRIYhEr6CAg1OSEvVhjYV3MYZ0yVF/GQ
xMwa4gsUvxuJWqZtuAXs5LL0GJdXe93aGUfUKdrLmkB3qvpBsCVYea4h7w3KXvic
Br60gdvomWhQzJOwe3s89RBQgnU5mdM6AOReT0AGBGzNIeUAwWwV7leqTp0uh9uF
jv5QvYJB0xUil27vk95mkLZFgCQ5B+Gnr6D71FqPxT2PBwJBzs0JVpxvV3TqfadS
/tjCPs+tPL0/nT+GE+JrCRD6w8ljLnWGdpNu168PHnExyk9PxerlTWaaxxEvJs62
VJYgwesoTTVHQ7a5nYZPNKtd1i/K3WLw8VgRuYWuCBQhM/RTs7J9dtVbkXbMGi5t
G7AkD3wGq9n5iNoc6pSVpZEBluvtVjkAofi6oktZklruCPm9IBVD8yXGklakfqQA
Y56T2xBk/kywOHotx9W3jAEXnk5EEe+i4ugGFCuNkfa0C+DstWqYoaEBuDI0FXPM
lLCZJlqCmsw0nazoW0oxWds1P0YmA9+eQNl8rWEfNLOfN0jm+OytBf1isHEX8OgN
CeXC7i4xUpNkadRycvFUKvz8/WoXokc+JM6dd75poLzpWxTBfoAKrK0CUb9LeEE1
v8/878hVSy5Sl09JYtrPCdC8STBjltZ0qB0NX7SAsrcIdtQ0bZBDAPk6M0ghoWTX
ujcBTs7suRfS31nRL2oFw9FaqipsqlS4leWFmyKQ7vt+zfam0D6yEu98uGRhGiED
kwHTcGz32ujLVmo/RA9mGeWWgVhBuGOcYgYCPJbga38VSLleV6XOSz+nveD0aqqn
pp1Ay1srnVbOvUGYgW6WyHISXU1IGScLcYMxYcL0segv8V1KmbvDjeGpVNSCyzqb
/YgBtzfKNuApp6AMFDwBztur6FUzSPvTMH4v+HtQbm6CORm5XxQGi8bzbD+82Mkr
MkM+sXFIp1UYcd9exGev3zoqEslxMgYHmSiw1iH7P1iSeYpROpDoYwWppLtFsy5X
sq1wGz4CLVydHQUpZwei5+DLnGInRDNmDHN2BJTmDcpZoUnLqn7ui+4YMznLvyMo
L/w3ymA0B0W8ZCClVeAi9npEP/rk/ywgNWd75MPv7ixfZCMSfikS+VTl8qAWycMy
AUnjouUwf1+gjvsXgXXqIuJp9XiZqWmNkZELesqcNLVSWHcRuHtbzXnIrrfQaBUU
8LVA0N9ufS/h/Ens6IYTIC8zyUSZeoIJb1fMo5sEYWU9M/XbmDHfrUmfHoB1gZjk
xfh/jhhIjcsH5NeCoPVk+HYWIoxyq575v1q0S6R6cSvmd+KL+CygHR4X0FI6TvcT
ZQUr9NmjN8pr4wlrNgcAY8vg0yNlaIpslq59K5uBdB3eRerAvS9XyNhdmPSILogj
CL/qFxiC+oxyGSnLmg+FiL1b7Wm5PO2W1k9fw6bX3suOkcaNvsb2NGyhU2GDNmd+
DJst8JMlF1/6U/6DS6Vu1OTAq9UYcJRDT10+GR9og7PrBfQA/IEoreEhTOA1kohG
ttjV0J39m0IxE0q+d2xcHPk3afrhCsdNXwTblIk0MSo1aG2B55nTEdaqp90nXNyH
kpzjCMYOuQqY/CSuDNURqa5IRPEHbWKz5g9LFtvebPq6KmSfizJwEe78EQataIRa
c9A+hnTsxsZSAG1anqOlAzQMz/nLlAe8kBru8qyNfALMQPaJQt9nrjE8to2gf29U
8h+hGogFTGkcPrn9ieX8Anb1qWO5sfzeMqD8QbKVdwL04g0SFuZCjRs0TbQN5jmi
oDpjYNKu65vl7ZhxY5kpDeGY5V3NgsXI9ltvP5ckOt6C4gWK8h6Hotu0xRNpaz/9
ms02Yc6T4q6ZeMohs2PetjdL6Mdy7KhcR2W2B8sPsX7k7cbRD9Hnucp8rzTw573u
HgF6ZdKqCtG8aOG/lnZvmQ2ucQhf/dDwezcEZeWYSzRYoTXFRiZo68lrN6P+OpJP
Iz5UNJp5XtMQiWtV5REOYft7jHma+4fBuOCgZo3RzOhOAz7OA/iWXxo+oKSdsoY2
kakWAqUlnhZ6h+9v0KnFX04GcOzKpmibZnrWBKVPtCvWB6wzY4hX3mOsHas++2sX
YxT8WTD/sptRBfzGOD855SOLVeDYTWlyaTZxFXUXoE06mQQ52B3dODoKyrNy5HHa
QxKpDht82j9uJaeelwjbg77vsNa+D9fmPUGYEfg8nzPztJZmVvCysY1nAs6v4E6o
C1K0aoZhrxFyHaWiwa5KXh7ZTLKY+CjIL2sbJ5u3xVmowLurFdbxq7nZ0OMO8p75
CGe1te3KWy89y3OZLRa1OegYU0YSAfU6tGdtG7XeCrBVJbB6s8dSmqmB9iINlOd9
19dhr5devDmyLsVQpRKTB/CCRl1f1C861YqZS4Wn/wq2vbCse6WEVXhurhA9PnK0
ZoJ1mRpGvpEkk+02qzNW56xUfpd4PW0M3Is9+s5IWZQKHr62Tox7rwPyyuFQeA3X
pySC4XzWNogCdBTAhcKI/5j5Qu+bZpsEz4pKALqwg1EEC0LfaLulGkm87gwWBHgl
22JVLTt+BcDIU7/QcUnh1SxqRZ+3h6doi2p6HvQJEty2uFo3wUUOxqezv00V9e1D
enQdcTMNy3uifFeJiKGR3NtuLZX8M2LddVHI5Rg2S3iOjMc3AkmkYkoeguMzRCOM
RomYlRSoko60T8fSEgpytB6P29G/eQxptb1Y9b/shedAf70Z9h1JPTQnrcuxD3D/
q/s/FgxFzmer3fZfAS50FlKhSVgN9npQwhexh3DQkSn6oayOTwJJvrjop7H0Eucf
tR1MqG4Ttl9Vw2vRKBOCallqAinGojex02aQjzu+VIz0o0SoZst/JBlE+X2PJ3WF
kVjkSXp/02Gvi8pwVdSa8ZmBzhtTXKlYH9itdc3AfgJgUwM/TBxt/52XdL/VlSHl
1xHMW17VuiROAxd03KxuwlbMYd478jtYquM1Mrl94spdlwFH8ckeKi6H1tOudF+G
VaZPx4LKkGpZTsnhNxcs0jLHsr2FcTdCD88a0wqCbripKQ83+3KSZucL1k0GIaip
nHRE9kk0WulaepuJ5wZdL6gaSyr0l+r8vw1Im1FDxiru3rax7vYf45r14BErC3Xb
iZ/R9teyB9Ly//wGKaGHja+guotT6BDZ2oIH4F4jmVR8hJE1gis2BJrH+htG1sHH
UKuJ+R2tueYTpfme2ReapttiuulNBn+NpIo3H9/VBRXd30MLly7Eob1++P54rPeG
wFN5xDPnToGQ6eL/Tg13bGBpxNdUDh5S6wVjWg+DqdaKubIThj81GmE3cxZkcASf
mdakvzvOTaRQdnh63RJ/o6BxNcv/zCZaxgi9TOszp60uTwFYpoPFRHxWiJKUUK84
loAj80OVGyUMBg4zbiaXyIv+VFIzegvbJxCpQhmK07oqvBury6QTITnNzJxieD++
/BLSbHay7o2audRw5h/xfjbBIIR/mUhrPp7l30VcgfmNFWn02IZfhbh48LFTVxMp
XdgSyE+w7MlHgl4cPmtQLlaCk7170tVIwpXoZxc2j9YTXoMuITpLptWuZNwzK689
xTa8dt+CLPOTz5ro27SLtBQrcIOjM4xdq4J3M4IyVFjwfsykh/0QrDmb06EXRaHo
jQiuGXX74KJYvL6XrkXmKQgSoBtx2dzy3BdnYWqh9SFrqrv5pdtKUntRqpA/oNg0
VPuXeH30fkakSIAVxdnK7y8foPZ8XxEZTccfMEGPaQCrRCACY3N54zBXjBuoHia7
bSfZ5rHQDvcUzXJKruIUI8gjM3WsdkEvX6ozHA1l0l3jgREnsPnR00W1r/gxP0f+
jjwho3OSNND+QqsOGvFdEGFWQ0dep0tFwfnNYkj3nlslMOYZMYk4jy0MbyAbxy9H
O0ilMGalKhwAUCbRg1JTsJgElYHzIuyisGnxwrVufKbqcCBUG1mJ8hWwl4Fr2Utr
H3/+wRoKkOHfPMnw+uobM+5YMzWluSPs/x3kqLy0mzZP/5GJY9MZjfFmgJ9umdAt
zl6r9duTkhIl2hXKgh/quJaC+yQt2e4rrNCXfEnoexIm+BB5bYXeQa4sOAvOAMRu
K8oAnwQM+dtG9MS48WnCmsbVVpU/d4HdsViK267TCknt4RaYt+9IPg4zdTyPhf3P
sm85+dMy3lsx+D1Af0/tO8P8xKXBVvR8tLiKH4I4IooLFVFTrbBslUSlv4cx/4el
RJNGTrFxBCt2Jkx//lr+zU4e/AbnyPjW6giOO518XFnjmAZO974zsQ7dEeF9KJ5f
wGURr0CydY8Bfwjz9BBAJ0B9L4npSrZXH+ILDkHtF7l/JhPub5JMp5FCPfYIqS14
5XWCLQntucoDwz4LSF7YZpGYxij2qD3BzdbaPbtZi+HPWSjsgFHWHdLazxT8lsPb
EJPEz35OxBSkdWmWNUk9FPLh1EhYBor2+Hhy6O9AuMMi4q14RclKKYW3JmZZphXn
Njda/s5dgbRjpBRw+3WWdPwRYOIw0/IxOcIuI8nVCJU0frwFI8LKZE9m8JJOGGtk
YjAW3uHJWf5VWEtA0XVciu19LZukSGM5bq6JiuFjPTZF7MGUe2CMk/G2Wk0PUxFP
w9W4YW70fYowipq4qyl6TRtXIIMgCr16nmKUsF80Tx0yGjH7BsoYXvCJAUvd0tAk
GzV12DjzsTIOr7oyXZ8GQCW093RbnZKs+kD0EdnTU8AdDjEdZkvnCAnDUactuisn
5/15CuPvNQsXqO8I8NReushMr1bEyl48+93al6OxBOeluCTqx7UstxlDsMcg5Y/j
ZUvxJVK4aqFlZbrQXfP07T5jQfWepx75Z52elmP09UAx91Wn59PXqO8H2iarEePQ
Al1yjuqi8cUCvM9pMmDeIRUy3YRZHxLk0WmQZCAffsFmzRuHbppyILJSplf0EFTY
RvpxQMIiRQnoM5S33Q7rmamdJFmyNMkYCeH8Ou/I5xdiR9dkIQtdGxcT2TMU/kef
zRRVh6OAnB2Szm0LpQuOSx6B6coiFoYGxGkTEc8C7g/lkrM2biy4auWRw5JlM12Y
aTyR6VhFObUKh2SweY2kjc2S7EYt4CYG3cBe0lHsxkFfcWLpjmtBqgZ+U9wJhsvi
iMPexGOVbEAMwZmhzBmBkZ4E508t9kHe649XLUQzMWOTbo9+Z2b2VzsabLKSt4yx
kBfdxsGgpCU7MdAQ7hNm7Gl6y4bweXjv8xdk5P9A04yj9wM4x6WwCauXmO1tSJyS
Z1q9YyY9nCvlFvjtZMTnZpfJHEYQC5BWZipFUMApt3eiuTu4qZp1S7kW57kLcZW0
LXhG3kBP0URmodls0Q34dZs1wjw53IJDw/jsZMSGpMUfOE2yHz7mVVyrimKEdK6a
xgI55CxoGb8A8fdpGSPYzYKFA+0xP4VIoF6Q1r/EbyCq5Pa55zn104l7/jf0UyQv
h7/OvJODyIXMiyHwUt6X5lwCEX8+YSKr/NE8+WkWkmZ3EiPNqvuNzxP3JVXQFlD6
U6uTPFWRZRs8Km5csM/iEc2Ac6TOE7dZ3jEc+LxGRovq3883U7zEY1TqH3pePpBX
icC23fKzKGpYyY2A0Rqj+cRPZAeg+2TnimyurZbgTXflX9O9eqWx5yUbHDUZsoO2
tbnZuNmY7h9SaM1423Jbxwgwazch0fTgrAw0uPKliprgBcN8U5A5rIyHM0qLULY0
hAIjiK+6y1DXKH6p8TehROfNBtdopEYMHndMwpmMz95bUDFItBpT1gi/5XzFX0Ol
ZBwQtnT+cZyhl+q3V/1hYFIoFnkkZYiUNxH1rep+kCBhtzTRd1Nqg33sHXQHlu/z
KELtcN4CLQIo+57gC0S1EBXoGgSi+uiiEFL89bIymlGr6NesO0Aj5WjHAJQOfsRp
TY1PmqwZjDPyP3BX3F8+wZO99OI1B3a77ogW3gVrfLoni1CKeFbb7KXMc4z3yoNs
n0Mn4J7Bes5hbIQK6tahqbj6bfjz5NIJe/+BqTakjqCz6jcJp15ZM53FLGVCbLqM
N5Qy7NvZoTSzWiVh1AZS9jXo49hs6iLr4O3jg6WfneqH+CREcnfVYLHxlQ1Lj0Nh
vyU0PzYTv5MlCsltPczGTvBVKRdfFTUghQknqvocgGqqPwvhegL3X9WcaGdKBdbI
dY+t8UlvwTZ8ir4S4pLWY5cBg6aLyKbHog5YUs6jPLce1F2me7T1KcNrlmWBmMaQ
t49jtOxS7gWuSqmSVrIhX6B8N8bIXgvujp/19OWYZgeF7vfTaKObxIihgB5tnHcr
Gcc9+ukw8sxKCMm4PGt4+ATynfkvU3DNwODmRfnCTs8Fv5JF15P7AU1/NViOgFS2
GVjEHxh82LZVXmtkGDhblyPl65RJjyhm1UflAiWRAyLQgWRC8vC170nyxtIrvlm4
Mf+iGr37+Ok2UoTkdAkcqn/9YebXCy12OrKjzPQizxVSYYIUkWZt1pdbtq41IMT4
ACM6fmQQ2GFWj1fqH/qIkRsxcBakUEkQyODkFuTLYwS3r8IIUxGRLN423BBunlYS
cuG5st1+NYRXWlRf/f8lF4wHPFMSKfIkv41PRsrKrGN2nrMeY3EE+9OHyEKFqPpi
keTTSj3DD7RuK4V7/dS97VJzOYNFTzvmyKfQBJIAqNblZfCmjB+Xm0SyNOpCglzF
PvdjKpPWOc004fPWnzNfJTdjyKEX2ROe2sGWoq9zJLqqY5r5xCsaNcGr+oV0+2df
r3ir0MaJht+rYs6iUnbgNs9oqn4vAh8Ik7DHnfebMC1JHpiLwxvNWo0/ZJOZwvXj
/UCPi36MnsJ3AqeIEkl/9OreFf2s6WVoGVfibnLnASYrohZgf3jjUrIJZ0WOq+5I
oSHpEfAVAKT4yKCuhMRutjDmMS8uEpzB2w8T3MYoC1FPMrBfjd5F1YR917AhPzx1
wD6+3zQk41rXOCgFGxjSEE4EK42Y8A4P1nrpV0akZnbVl7iEsH231rzXPqa9lJJ6
BgkDeCV5TVFFklijEFexTg6eqHXwf8DWMAg6tg3wZkLoM9UC6fkuej/NovJqwkqx
yj6enKfYzJ67VeVugASycvDiDzixrjNEI1CzCetbZrKGnqL6IcrdihiuA9jwcV3X
IoA83N2CwHq86wN/GSuxCsjIScUPmaNop2OrB26AZUkyhSymQW16TWoMvaKRagT+
1KIOl/oU3BowfSdReTHM7/9eLuwGz8O1JWs5kWP6eIzZ7kr4MViFcCN9V5R+wAkf
ouZPe9Gf/LOtZogxUnyh+XwmfO/2ss1kZTXrr6lcQxcQj2AKzAjCkLs6jDl0Jmwu
8jBbAoLvfor11XsvWIVAiXaKnAberxydw5YpxPmjyDb8+ABeghXMi5zUrS61LNaZ
+YFBRX4wfvtPtASG2HQs/57Qvr5A+1oTVfX712xUkAiDxDOvUy/EU1G/5LOv1Oe4
ijfPUfFmleuZlICpCzuBpr/7QJMTqGYsalRnWX3c0XZJm1/TP7tt86HoPXY/BUSg
hsR5Z8uupVpP978XnxFzhEnhf5ccK4+3cCvlGN/BiU6yVcEjmTJ86YgyJlAE/w/L
LM/WgGZFYnPLRxczPt8aJckYzp3XzM19vIUybGh0DC3ktS/MyxPtppZ1fY2aGjxO
mcSHXlfwU+l1AqlxjETbgna51VYFlIeSMAwu1lChigmYx7/iKfuCZXtM3dhNFfua
mpqIfwDWpvWzX9eV66TVz0PaV9+dE5qm0Dl8Q76/w4o+uMeRMy7tSgkgw5m6jV3y
s7uieRiAA5vYYWJGkWTgk31C7z+GYuVP9cAq1xIUQCHL4j4dSpR7OUd1Ov2B5Poj
0MZdEQKcbAPx55Th965/3E0Qp8kSOWSj1IoAcOFzk61TQn7y+i+t3bOLhAR+aTcI
L9Qmy+7EMu6xgGfrbu0/GFi9ij7h6IRX54XQWSh9xPDnIHZDIf5+n8fzkhGSbAWQ
QOYxE68dqlzAa3qykfeCnVcVY9mX5Nn40mq0MnzsvcXiun9yRhKOkiaYSwxv8wOh
3B6WfB4fa0YuxtLVdglxdhTkByIoiRqMGbvOcNhXA8RwiCYbaTASf5C8edApgxgU
7DTAb3fZsBowYWVjUjQXeX5hhcG8afFlssL/OSRKl5e6elc6NiKdS0/gVhlOj9HR
mx5Ch7icei7+QafmUt2x+BWzHGDmFlLNr5QCrVIIdK6JdLxTN1APiQI5n/XiYE+6
aetluFpOJiwuMLzfVZFjvX8j6gqB/9mXD1tI5mnOOLC5L32AdAO2dVfbBgSPzfSL
2nDChrlElJ3sfEQNSarrhiVzV13t4nkSCGs2gejhIpBh365hsQW//RXLV79mkcZ9
wAfIwRTjmDEBZpcEHUlA+BEdwcr8h7y0PlI1BZMVQsd6l4FeNTK7FXLoSrCYJU/C
Tyiv5p1kK0e9ENIaZCRHh1HgFJ4o4C+wV8YPut8nkdKSiCnwbQh0tOvks4vH7khp
s5BH7VizdDfR8GnHwtG9f2Mz4Y9r8Le1AYhco/DQL5qN8g6+E7o5fRK87Xhtblsd
YQWw8J7iaGxzHyoY2qch2zbv1Sum15klvWL14DTzVk+BZkZgQ5Qf+OIsoT86Obml
hoDi/WjRRBKqOlHHuWlT0KTis+cm9OPldbr9XtV9PZJUU4K8kStUM9ORvUeorT0o
1FyNoBFz0NgFp9Nc13Mm6ngO9HeAJGCQ3kkGo1DiF/xV0d2Ku3ZA8LoCp9NDnH/D
SXlf+1wS3KzEGq1krDU2TsyD41UCPgxj0fuOzySNiwPhHWUBMYA0e6RkaYbphM3P
MG6+Hgg8Qtj1DsOSz+fcwDfVzFa4GxiGg9hBD1AQszfqGcR6qw4KqrLwDXulCHO6
v9OIsiqPk5gCYiDhHImdGUsnTtm2aEoV//VuwzL/Od8aBVzK0JP7z+ucyErLARhL
RSKOwLNXVsnxjNaRPdAKDTkDmCg/biDJAca+lMSiV8laFjCP4euM7GCL4T05a/QP
XDFOK6tfYzhqjU9/cJOKUvB3X3zyA6fmfnFdoPFU/x9tfOVwSGPFc5S1kEG+Js49
gWsv4Ow/b0PkQCuTgsRo8D2Zi+633+wLJP7D4Iz3jiV7s0l7Jcc/+ozPT/UnABKi
8dOfc1AKKvkYIdv180wqXPY8+YqxNEMn7w3YwMU95sQSpvqDy0RVpBmK27XdZgbm
UgsMfDacLtdty0YF5AU3MDM/eb1uMEBhVGfuet+h5DHEzEH2AoJYYGJVRho43shD
FtDvNySVfrMxhowYc73QJKbtLNXtTPaOf/DSIWmhi8xbr7YUmfxlEB+sQkEsRINg
rfeFdqVpdjMISjJ0yAZladKo+6jXC5jBlmoe9y9BWE20r7KyFZR2ZrSrgurv7G4/
xgDDIqr/Nj3tqjDfm3znPbv7ov9BM6zZRYluf1VeoIBpkHkSfrEMyOrhhB9YSZML
FWEIp1RJWww2vsS92xA7sddQ7TA35hr6VlZ+dJmudHgizg+aHFL0nWK7zETIpE9h
uk09q9EdYKlS6nWbEvsE9kA5n8xdWRu3T3Ydzaijh1hDmHAGQbwQj9m8AZ8QlKWx
Vk3xanMt5yz43Du0RGwwmAQ6MkS4llNG0jKfSflKG+fHMf74Ku71F+sp7O4Z19uq
CqO16cZFLfngptdfi/0z02YbBJRk+1izpwoMZKmVZ8saQ2muPlnmfv1YeKRpf3nR
CJWY1d9ALMQ0lueHCECWx9++xuctwb3swJ8EBDyFAJENCkVCw0A7yz+TqyDqhEjh
qDIbNLqIdE/8Y1TCYrf6awbNx2PVuiWptM/yUVuCas9hTjp2MLwmrwe/BI7PJHyv
w++qJUPBKYeq/iUMWkMHU8Y4C8bVJla7AsWiWVH3XKmR3/ofuQjmb3GpKyzzhIPl
Tss17YySGl7MfPYeMAXh3yEMHEyy9tA+scV+U62v+A22Jwn5CsgB5L+ivswZkg3d
qBZ16gsocdH3I/ZGuy1LAYPHEGsoc9yCWUguwMhHyBmjAiqas25ryR6WItR19CSB
WU+b4q4KEqSq49Sq2DUA+3wxcVdfNwrG2FrnhveeHmMzpWCI4MMIwPupTtPgKb/V
H7yr2kDBWy7hWxcOQljB/VA8Ke3zs0bnZ3WkSkqEaBg042lqW25tlSOXVxxgcp6/
Ts0k1dViTf6tCv5kRPYbx3Ys85Kk5lkDe9sIdZWYpXIQMSkIImynSe3RqgNgpejD
j9vRyRAyMkynFbrzhLaBpM1UmyA+415+OxtVpDr2kB5nbmGnNBGBTxmV0XhktBDS
cWDPUSPj3SriezgVHP0GSqNIPsm1/37rnrXTlbpVD0UBDFQvUf8dhMoAVdTYSUou
TnLX9jCYZukOUC+txms5rIJC9q3BudDyptDuO5BX9ssHbWYrkyAXPwn2jodKXwHR
fdLSJ+p2IZB1sB9K6r2eE/PNYB1O+Pd8ltZCXcaGo1mLlG2etuJdm3YNQaVOP2Xz
BTPYCByKkUwG3ufg1SXC+RIYThrWNeJD42fB68iSU0X4atAiYSfjOGzzOVMb0uHO
Q4gl2teqKbsYP1TX6X8SSbGC4CfF+ABVvbjZBuJY5Y/5lcbNXLAA22jEJ7IVM7hM
/6tq8hfGom6jwyVL97BFIVGNdeUmvpdaHON8/UNkwdJ8XJW0M0eJ20toVFDjIN0q
N2HkcoqdfQsN6dujGgWq/eqx5SkhMaSqWnZFkHj09cPiXpTDfNxiqFpGH0+EpcHD
r1xm07TWD0WiFKxLuVjblVQcPZ2B6eMdqGVkrDGjB2tC0FyEnJ/YbzWYUWlrOJ/l
9iTTvUELCS7bzdhwSdi7NUJxg57LarmNcV0GeY5e6tfP2GVO0UsOQZlX6Dz8Qo08
TjjeXzvrnWb7T6aVlHdWHZ0iX+PRMIWYf6UwGKvaCmJg8/gYEZbe8KGfpWIB580w
Sg0Glypq+07bFelODPloimcNc9U0SP58hb/x4LB8k4LAHzsgycQvt2YH5KH4YtLw
AE6jfePcbqWV+51d9wcpLeo/IVkYdBpAPkEtuTQBaXjbZ+d2hRXbhsD0DZ5FyoAy
eLRCpRijjNUpKWasSc3GhPDOtNzzhnSdp/JVob+kRShZDjIR5nnqko45nbXb8YeJ
CxY2NgSv5Unqv4dwUgBs95Hz1BRnmHQmQzfcSbljPqOGXLie/Zkm4C7ffuS4gF4b
KvSbiqe3y1tujSr3Uj4RhM2jLpbT0BB18qRDGbbL7Y5BCIifc7SIwEiSt03irYnE
L247e1AFPfUc6Rb+sW4auQJMixSWaurDtjyywsHWZkMKreD5kEbi2kUH2mJRvAjo
1v++SNroSto399JfC8cjQJw7wbZOYd4J1uu4iEKExZNikZVmNYWZj4BPvJ38MpgZ
8fitaO7HlJQ/S+UI+jBe9RDnTR9nzM0FUxMq+Wxqs62GN5zEgfETAaVoM/61fDYd
MOlWOcAumiHXi6sVxrTz1PCUMCb0XA9G9H9l0gkdRhNs3ZpPPu/WEE+U9bsC+Ggz
0bvqy2aD7vE0LMEENosyOL/TXxnei+Ax7JUx42RFNH6MSImVlzCp9509bxUZoLxV
hH+47Dfw2Aa0Uvt8NICQFgsEuj1RHQWMggxSqsAlHM5zzbM5B3yJnslDt++MVp/c
mrk9d67pRNC0jI5cPPNWYOat8Hnqj8LdZ5hDc3NwZ+xw2Tz0iVUjqRy0tkFMs+Rg
hrH5TGEkp5iJpK8bKepcDVUfwhwepWUK1eP2UYLoMVmqYIQhIc3KRYTP+JYewxyK
4Nzex183Qhws6kLZR7s6kss9zWtmWmJr8y1dZaq0H4wYMbg8C6G47aBY7dmqVhVF
dK5SSLyqNKuZafKGEgs75BEI9k1/tEV43G3iDkt+PPcyIH2nOn011gbADCamJpeZ
MROULi/y2HfG0Xa0x3RXxrqaEMQOuD8vPTrL2yxF0LCpF6VWk7f6Tf4/xJtwFTN7
QGMWG1OwNjxswun8FY0v/feKVYst4yGtYiyDAPVvezG/6Sm3xxu5W58Xq4aSuHah
mijKwQiFQWgPYKKvIecLiValkjfKNt5hMnWEF49G4fRJOz4Kjpf3857QUa/pvrm3
gt/fjlKDkm931d8EcSehcSKJ+qQIbC8/exU/9EdF+GPwfwkbptpLWFOsTwWjQZlI
iVIke88wyvDqIQ2ltxdOvrHqYAGpqjrkEmn4Vt58Ls6DTLl1FL7rsHBAYuf+8cNJ
HiQmbPI3RBUB0e4Nao1+SaUuo31Z9rLaQKh9QfH79lZb2eNXYzTXu07hefnGMAYD
dZVqymub86vI2IAxozTov6GS4sOLX5qNS5Jt3YeS1pT5kpc1eTCK6YZqQh4Avz/d
kQqA7HNOadSamBGo93XTcjq6vnLStVar0exZqDq5zVvVoZIbhbnbz7JuXMq05gmQ
XV0NH8GGc8iuLceSn/O2b4IgVHv4oJDFQP1Rhi5rAGYvSMRqwKrlj6rFVsFo170P
L6DdxK/36IMMU7ytzpfei+nI7WhrS/HYhx8F9tsddc82y0S9rT+1S+LGVD0ldRM2
QbsZsa1dwGkBXrLZDQwasLm4i1fE3JyniHZ2i0PNpadb1GkEQiqJ+ij0aDz9MHjB
RxGZsI7FICBB7gBM4BTvbPU2xw5zX5+w7jdS274GIay79IFYNFoo7UxGMcgZGJRG
Ci81N0Dz7q3PZ2fuiPUV+YqQhkCBtydA6e8X4NQxejnRAHjpyWvgzG2DscJ2MxCm
qdfOvYJixVqQdvIS7TiZUhtM4rFrAxbeeyNIZO4mHSMInUFhiu6md6a4fx8ugyzU
dmJg20OSxmRnrS94cMWRCrPLjGyUBrfpW+eXAmffoghokxwrhgbeH+Pf7cLky/9O
wBUFkIO4WWGipspGQjHKjtoq+1nBe2/p7DzQ3bXEcsScQP6CfT2Oywv/LvG0o+Wp
cZtDWgOsdG9f8vCuAjOk7Mgdrv2q6vLLP+0Wgvf9biW2Wl5GW96vO8TfwYWkvp3/
bdXX3IT6G5O+ILC5fMbmeQF00WkgvMDDN1xRcyQ0jDYVYrNg/7dbF8WZECCY0SPt
skm5X70Twea08QR8iAe8YTafEfGr2S3txstvwMqKr+gRZDGfMffLLsgk9Dj/d9d0
8TLYXFzsLX8tQLJ1BAU+M48jOSopBkDurSWkIdPRDhYltrH6OZmzKU5abWsxZYOe
6B6lfd0DbA3fiJ+kxFL/eNORQ0+fEy6MjtWxvahDyviikBtCtOmG0xY6DloWpfua
Mlybsv5IagL7rjnN2dtgE7xPeXmvkCIkpzIrCXE22phM+u0VG05/U8mCtTPtW6+d
0yDa86edqB9uXWBEBQIgedwQqxEv6mRtYcHFbt8YnOwnAy/SwKhVJRn03ASnd3a/
yA7dU53/+Ko8c5zIpKt7B5ijKR3vqXWKdxFPsO2/EKIFeXHVDMw9EQtzAnySvCCo
dUHAeeg1LU7jZI6fRutuYkbsq+VwCyJFoZ16Mx1cP9TL13B4bhZSWSU2YEBq4RkZ
qRGAb7ko894lH2a00fkR3CXGbc+XKSCK2Y4NTb702mZ2v62yNGH4hnqLCBYwsZBG
bjbv/DVZa0RDhlwIw9I3qICoVzeWKZWk5roLQMR1N95nRGt23QsHfVU24r254G8k
2kJnP5VMA9vyEuL8iZWucNZBv5H01RC5BOtqfYtBLLzq/dq5atGpGQBVdCiKrcsh
q0OTd/PYJACflRfakLCtZB3Bq6vZ6tn1Faq4vtm4vmfAwluLXJmBQtayRnB712Mo
Sb/x9chQONHgfqEwRTYATD6qGsdsS3vLrq6S2EcXgKrYVIOUqWEX0FQosLW88wIm
ij6j4XWOwfIIWxPQQLT86duSVIPxMGvog3QhF6I0lYJ5F8iL/WC8iDE5VZ7Pj282
JO7T7JLRb6ANMSgQODEqIiA3lEPG5XHXlJJIuqW9pD0E5XYXP8CKx6xkaRK2Go5a
tHzqtquuGBRBet6jyz3jT7Vy6nSIAxkHb4gwm4GNNWC0+pMS6AjvDru+hbIndovK
S38Podi8TLudMmNbN9WNNMKcltrhr1PdxNQlT2aXYICkxBXlGzGH/2i+Sw47ra/D
dP4nKQ2z7tsreaEf3gPeraWPibKOniCmPd55QhHcfn5NHIdrVGsPGXRrHk0cyNOO
Nz6akRYZglo0iRnDigHJ/iBYB5CwZE5vV8jP2C5lz1wiq8PT06UDFA/9clcAfmLw
Fj5t8rcpi7bRQIm7eVCDDpgw61vwJlsjm4LfWQb0HZHR2AZI+iRMMgEzGEcpYagP
CN2coWES7Gy5bI/iPV1eDmkFHwLNcFiu94496KnNEakMbSoQqcMUWnjAkx3TDBoc
aIgCtLeYcMIputIy41rUH3Y0X9EZDMkc4pxz2Z0BN4RYdgL0y0+/HT1NVQFPcg8k
krK9OOoiL6lQR0Ko1ya1Nzkjl2+BG9m0NMVYZaaFLrR/9oIpNigSw5N89xI1dJ1l
bhH3KMlLza+se5IUAYn9W/vAyEkM0f7Vxq+jTAX2pwioP9doL4FPNKndMIrWpq38
JPtcBg87ze5XNtq0DsCMH2Nb6xnJdz1hUOPOBQSwrPCGhco75FDj+vPypEykBQ4x
4E8Go+guf4/+nOVkV/89rGEcbSkW3D/MxavOLhtbdK5Wh1Ppvy4e6/rWT4D/uidW
iG18p621tgu2mQfA0Ah5MeXrbFPIUjjAM2EmZbDuyCYfxEshwDNT8ZtxzvVFuqrr
hGEuftuW4pdvC/ckMMo/HjJ7rJvgoU6TvR/KZuBc60aBqVhGsTQlDGob05EW+Kno
cmviwJ5HvWUbJSTfNlTJlR5fMtH1tlyw3EK0gOoTl9QrzbIHXLIw6iK/WYR9EqW1
iNNNORxV/qvK85/voyF6HXj4K8hg5sE4SmpFNmDLnCp2ETb+DKQEvuEE8MSAe+T6
d8uiNRSSJmPZnpBkClz9sfCqc+xrau97yF1m73EPDqdhiAIBe5m4LULPQzkm96f0
RLywWNxXgrXRbwrEhCH4HtnJ3B8bN7prBShS14OeqGOcvWMih6joUSf7nFN19mH9
1FG/b+F56xinPd0ysJ6iJioPD8+rfzMY/SWalY9HK32RodC61MyaXi36ssoNKAjT
+1AsjIS9FdI7A++L0l2LH8oEQaL2J3h5F+3/NxVala0Kt4horXm22+kIEpCLpeBt
o46E9/LhHhDsWPZI6Ik80+Usi+apwdbWqwL/I/6PKCYZrEsK62OYuqqNLMMQqTBS
ae1kYpiJVTUjUyIe1LEzSpsQ2dB9EWZFw4/xtFsLnXES3i2FZBQEmryyU24qL0jC
9flWM3DpnTHEwUwPbXDVePa7yr23b24D9mH5H4UL5ADfbTBnllpdU1Y+fxly6iic
zoFY8t5vwT650iEVbMxKsSuFiCsT/La9iRBhDNahrcjWOGq7aLQLHAkjCruVkE+f
FIkyVSGQju601Kij7Yr6QE37zocqSDnJJfFUoSKuV3UWf5L2W2qTH6d4YTV7139d
MvPHrqJDM3543JMRgmFUA8citfTJlz1QqLqTZvXeRJXsVpcytASKq7qrJ+KRp3rw
Ir2Qfgbl7RTi61ITTWuLB9hYU93iPlJa1mSOZHiJtkt9ET5io0OnC5R8DfUFqMxy
TnP0FENOI+gT4+Zzq7rMz5kG5xwNqdNu5e5PQFNn2gL+Gd3nHJoLz79ixHyJEx4R
6lVxlyA1tBu/l8EJr4lWCmX6PCHXL3/6eUOZyaz0VjwsWU5USeQHkneNzJFwkQCC
thvQP8LlRIM7PrdKeceIYjqa4gXr28zn5vWJ0cWtM5BXg6I1Ol00wcnrYP5Nh/Wl
N8bSJLqAQ2NuFkS9TpgGhUk6yJ1jagd+JM7QEpHOr6X8mfaZjHY5h0d0tQI0ht//
X5z4rVU+A3CqKCm6xAa1MfFfuct9I/QV9KwfgLvuLGxlJtm+yoLM3vmuf34LAwDY
AzS3HO4QvGHZ1tbSW61bcKIuL7mkvsjU67KjODWaDyOIX/10Z6VBl0V24pW+AKIb
uXzDBEzI9jSJLym+SGp9iAI6MFmCzdJBMKMzKySlj7Bz8MZWlzYIql7k7bLQ+qHL
9Cqvbk1f9eEmkWPvWW4NDL6WUp4k9A9mDV4HtTmj5CGj6DpaJgbb5MPUHQnSg/CN
eTQH0E1BwmLpXDDzYr0vhPwjNH6P/G6zul9JGHNle1Jiq2IPXwmn5B7g7UL2j0qR
vtMyxIATvVcEMPtQD73k/7OnPxqZopXSvp6DgeLtgfAGI86ibiRbwL2Uun/evIz9
V8bIRsIpLqrNjo4TUnTQonucSYQO0piI+ACr/OlS0zVI8FrdMxN9Q9CelZxHH5V+
BFjGHBRJ2Fp1XGwpw1so32De0B4h7a+yI6gJct/4mFb0EOYu/1f5YYaZ6EKgOXv0
7+8OwJ4rNGGhNntTUSQIS3sPyAqdx5eb2/TtDQr7yuIflkWsZ3UZM1d/Hq70VAk8
X+X1RXEycypm9JDMV86+Bt36qkIZ2i9f6PBVbvRlUDXmqF4sKiZtM7BYiWgUTsHl
hIvyA23NU8n8hbbrE/JDY83YnVvPNqt+YPqPyWDlTX30xU1rdawiN0DVJLEBQEnc
bQ+tWFPSivHcR9oWh7gQd7oobwvzRpRr3Jcprkn5U8TaemhenaqOMwxjENEpk+VJ
crShoRBgk2x4B/ZY4wPOJL6GuWsQKZfUJZBSZj+LN05YMXOg5sDPX1bUveVs0xm9
eHfIrquJYBoBAZTrdtX54n0ZKMyk8PppccAICcft1PtckpfBsWuqM8TksOtdnOh3
wk5mePMecJHkAkKtYSboaoGTkv2vrmpWOIPD1SPej2PSrfGdHJnCy5Uik0EhYENi
l8/E7SSmW3xuEGqDsFupMLkZ8uRyUgm007GbFB9/xgOLQcmQdZktBTcvu92M5y/q
2xGfkN49moA9xGGGMb2QTb1pGaji6MsWamXGyc9SpzTVyeW87HKH8wVrXUCsj7Lx
lJItkGYEsEhw7Nle4SlV2Yz7Qy/sxJpDq0Uockkv1m4jwswamrEnEP0pbmGATPbI
GkYTjtRTmlcHG+w04nB7ORv7ioJvCKfxWy1fGAEi1HHohdnXeTZ5gYwp+spkw7Yh
6kyUPxxmjNXAuZEFRh3YuilFav7jt9T2b5piafvhvky3CIbwgwnVnQ0v1FiDSVxi
UbjnLNWocjg5gw78hagfHsMUK0cMZG6qiD6h3tejD9rJehOCWh8DC2pE6wtK/SKO
2jC7F6lS+al1H1X9vwRQ2ecqKh2mI4qNw+5isFWmgK3C1nYBIbLLRKRHiu6rNnlM
syF5QdQW8/yIUvD7Zk7ua6FMqikYD6oyCibMMD81/Zp7qIhmbiuzsaj8AyLcB+eT
guXgtRsf8a21r6CcVw8cQHSn74y4VtAXRTiNzYu9phgw4S7D8YpBuzr4jrL2FGjQ
JB41RdmlIRpL6lM2PAG0sVrCSDSRrMe+uVDhxFaMGDcxtBFj6RQJ9B60dKMCNr+a
/P6y47f/u7lxinzNRzIEo+7LIL10bt7BEMX8d/OHR716JnYqVVg1lHKPZDPUgitu
e7p5L+RARTLLJc2pRZ4w1vgVmPAbW5j5fTuHM8ZGE3gePK0J3+ZMZ9OpbP5OCyBC
82Ab6bELtsyASO3te2qtpxOLclhrviBLSt6e6ev/XexOfh8buhMPkSD/cfRPMR6a
ysvFb4pxtzjesF3cyq+j6uvuXufgIZBap7+cEXCa8ZTnv4iWZR3xJoQuJ5mz7BH4
apuzcJD8oe7VwtzfGqpctSet1ncYBfbgymwrMv2uyVxx/LM50qQwiaOpYjUDUcZb
zA88dnLuiUJpUurEn9NQvbhSDacFIWVSTsV5BrZOL1WdOu1rGWitodMcz8H+19iX
SF2/7EVVKmIiwMlYjv8ePyZLSaAzBUCKypyFUmutrZSX0RV40n271DLiaw2+hJaq
K4JqB8up5hlF3STM8wzwPBr6eg6xco9+ayE1ZjSkcW/VDzQ0o8C2pI5Cj0JBwcBn
hgcVRR/0UTH2R4m6OjjbP3QjbbYnv4fEnDl09Dl3ZagoLFgU1+PY/+k1OJ/riqtY
hDUKq5kTqt8yTje2ELqFKAag35FM2u2jOk5zVvXVMBM2ftfZI5dMFOJP5rIfqzwZ
kRARgc3MghHFZpEQELrPC2OA08XwcqsDnQISIDGq02YihdlAyGkHuoUGI9SDpvpT
83l1DxB5J16jcEMmLHrdPd7TYmxLudCguDWoLuHPLcIApHtEE2i7+Se5pLgq1cDZ
UzG+vSoBWvJlIYh7bNUZV9lMYu8c5kJRIlHTzvf5jRhiYZ2LGQzWGldSDUGXm+/7
XyNnTNHXp/61IDxwUGMtG/rcEWPwtNC4hNneO58nGp8wp09sAtYGnpnAsSk9Hz1j
hxI3gTrFYCWYHI9SHAILW8WzDOn1OEeSmG4a5AY2F2rKQtNj5S39Ad8Gcpnf/A7b
tv9HL2ZNbqjBhHZGSodav2S53oq1eidTlEQD7ZBzLNWRDCOiKEWrpnYViSpad1qg
vsja4reKljzLhbtrRFR+YLQwbp75Sd3nPNK7A+8gsPpNfEmb0Fs74THZhzo0o4W1
r55u1VUwb+XUJK8w8HybiWjHnfXagBbbeF76cW8Z991uH29qgfJOZB9DbbHQif3s
nY74Dhea0EU5KD1inxQMQyvIdTvBopI930brQtS0SbqQOW4PqSE/qJtmfXTx6pHs
Pdryq8x6R6v3R2wOyt2FR5zQcPf5l4HRdSHlcl52xmEJqYBzledaE2IRJzpICxdN
ZVqY8+s0d3B+2YngvmlJ84anTQSxpP3Gwyfv5E+Cviif/3H0Kcu21yLQfk+M4QSS
j9lZROYh99XupFxUKjxjr62HBPXP1plkyczA9ev0fzwMV5jBn1c/CiqUhlmPDkGc
L3CKh0cX7qf9cJvQr+tItxOPgr2NM2YkknwBs9Daa0W0+k9cz6eKSRMZAfgGWg51
np2FAZ10ABhfaKXTGIFzuKrjyqN6isRRa+OPty9W9MrB8l69lezuDZELbfBqqwnN
9zJJsoGAVd5nhc2oCv0+I9l4+EjcvWHYk2tw+Q9omVc7ax/Lw4AW4mn96P9caWpC
sLYjbiMkVN8paWtz1tyDnu2saHOqfgSQj5oiZe2f3/0W5IRQzHDKKmdOtbgYZlRr
gzbKidBghGc/Eaz6XgW9O68kY64zh8s1B1L3vZPosj1UgoL8B20iE6MCZNXsbadT
tp0V/e2++e5YPybkszwJoJ8v4J/H6LFgVQ3rztCBsDED/+HIYqYbOvWXCVVk/tki
HtbjjuiSvGZEOcostlhK9VcH2/VujSPNjs2FM3olOuLFTa54NJrrgllCTlacfAfE
wtFM/c9y1AHH+ihdPu3o4Mm5Cx1n6TtOr79z+I2/gCcQylkMNXtJhlYjpmF6OIhe
oAZOfNOqFsldadvCvINbxAm8ShOVZaYNqgKuCwxibiHgs+Su7wnMIcSx0r6/jc9c
Tt9NNEWtmOipeAjcZozVq4EyIvsWrz3Kz/UP/nYUS4ry0oYiRvc73Lm356lKJoSm
jOtdGChb2t4O2ndEJdnTaUGSG8FXuLpfIlf1U39iKCga+6FyA/3sFB14fe70fj5T
SDLxT4QqWsWGHp0xKaV//ROQ2z8883gc7/xDdokzIvatWlaKYC/gwNKEBBSLzjwF
j3Sq3pSogM0xUoanxC6y+1o7egS8l0giu7xJQ5bRyaAs4RRJ+hUkbP6uWLzltimX
unlUEC6rbCztFPSVb8GM4gnK723+8KC1q89DDOlb1PG3bkHI2mwNuqpFwVhqz9Bo
AYcS+lggQbm3MR+vvCIhtH9vNTUyGyxnI3sw6grP8q848802jEeV0GKe7oXSWyx8
MvgyegT65RdkbVGDK1hzXnvqsJ5m+C7kOahRf+8Swyh2tuqT6n2BfPCPcW3ZglBK
JaDpGaJ5Hb4skNpHjPLwZ6JjMSi9ElXQS1kIq/9CLx6xac5AHowSSNLF3Gpeu1uP
3nIaXVwJpXtIco43jcLJdXvUyveptEYpLG1l1gZ2UPF32Q58MqJv7gx9n3Iqasci
G7TQZ2zaQfOToEGZJ2MkfGKB/UjIpJvCr1jZDMCW2rY2YQewgg8OxKZxY4hPeVjT
SvfJV+em2RV0WB24SluQYc2Iyi06/NK7k33Yxmy8GoCKtRvtueyKFufKM4/X7GHo
68wrwCQNrrAps8BHZj+73yDTW6JV4gRf9Z7a/bhKBK4n0lBA7jhD/jHctHLS30Bi
Bda4Fa92Z3Icd5+DzvzmJ6f05/nrBJf8flapwJ3lGT8F8Ct4o5t2LUOeclS63WSK
ByumCojkeTQeoYSC/2VdijLJZ8BRjxmjXtU3WjmFi3N2C+Hvq0kqh9va/1u3Sx+u
FHIcj/sHVodyhV7MSC5cBzTs7W/yrZYO21wIlLawTPEKs91MDjPZ+b661+4gZaVq
Jq06/mcyhoK65BlBnj970rYNdMDesH9ZRvw1D0AJTHHXCcoHiaps6NDbi5orhdAs
LMU1qT8hndNVxvX+NEfmkTyvd5wJaEtf2u9J7+JkomcgXFyrtK0ObrQWg4E0jegp
CHkeY+T9//paEZsxyOpUsGjl2KTT3UKqnDXgRzGVvOPDpjn+JHz6hgxMOX11V9+j
7lUXfnvUrAbDeWg18ck63+E4yaSAG2/nyfMAlEw4Y43rGNWwfhXrl9NaJGJSbn62
aeOp9o0u/m7Su39DrZvfQJEVI7KXm4NmBTYQ1xXAU58q/uNIOuqb7PtOyZ7i/Fik
12zKL35L3u/vaemcxcP2QfMPSeChnq/UUvuDRL2j9bwX/LqeigD21aCLpqi3pcer
ih1SeXCGMuWPDbG7QWUKosPvPdw3Y/HNo17z04U8J/G4kqjG2lk4FwDCQ95dSKP3
LrD/ycw5bQIG0qYNpxzyHNGVM5mMqAWJtFvcD6EiHGZQl773uk4R8wSuoevKVZAy
mtoJ4n0yJJCpG+fRcVmqHGJnJS6NJoN9SQpz2PwWw7exVX18LEoyQ0S5Tp55sb1J
GFnRtiqjbYHM/WNP2GMH1mtP9vCd6Y5tCzZMUOsOAAHxEA6WTrwNMMlrOWJgwUpQ
ubygpnLLo73JF6P6mKFUNMsVkKR1xfKP2oe8Rr7ry7JGKVj4nHZ/6cjAO6JCmfx/
umwRLNAm7HGEbZs6P/cLApWdvf7yYcSFoXPBKHFygvijYeWxwXE4N5ML1+9uAhrZ
sceAEf6WdI5qbp1+Mey3IfzjUTaIhwMAoT+yH2wFEbnFLHdxDRrc9uCb4X1to8NU
lrjBuRRbq1Mzpjxsi103HhHlO55R4hYfAbHcE5TKGK6D0dz+IcydjWSkdaWBndgo
LPvuDNFzeoq386bKDCJj+uXfD5ku3i4EM+x8cY3D9Q9CKWFf+PS5sqk9yut4GdhG
7Z+CHpGdWV7Bve+brS4ZQA5fFwq+CIkwoXx3O+TG0NtdSXhc3vQfpTwoGJoySHr1
tq1rmj9laZ+tM4QsXF8cG2QORb8G8YrjLAE+moPULao50+Im/N1EDy+u239NnCuU
0BY5UC0lwPgvGR4wBbPOhIYfA2B09KumqjsD2m/zPpgmtNoFV5FtE+cYmJsM+UGb
RGj1wWuD1S01G8db17um8E552Pj/GoSgnxDz8KVPNHBr24yXLIWmtbEkjduHWSFi
KscfIBs42CO+6zAmQ42UrX32zWve2Olql9kaySiEKggQWKYi4KAty5THkiYNQJfj
UmpyOpAKa93L5GMAQsLgjuZATmYKjV4+we5rU70/jP5hi2O4b9Ty6zvCbH6zGKN0
g0vz4Jbs5tbytaKIVMxRLXmbSEVeDMONDbfys2ATbT1UzoRMsrcpm+ftySBbxyo/
I6a5pTMeyyhMAZ63VAJYPSQexjcW/TxXMoxizxCrq5vCgYiBz9mD0bXDAXPRq8jL
VytEfLV9Uzq3sHy3fSiR+4V9XuN6f6mA3zAv2aiV+tK+TPt7Q2G6U52l7PEjRWUv
I4CqhpA4eDewgOvUul+bBsMnkXt2HKmPbQqgliQkizZo00D/sM2UTtvzHTTP1MQW
1OeYWLuJTlKgsDH6/LPt7IzF/TL3H5L9N7BOS/PP+CTR5zJs7lUSyai8M8cIVKQJ
pB1nnPRbXDM8N15dVezxq+kNyRGZJHTNaZ/lFmpr1f93wPo/Tc58IFygUZ270YQx
TDthujFKz86TUjYfMuHMp+8Zke4Q7UAUBq+8Z8KDkNHOl9Jh8x7YgpP65PH5yW7a
fxdo+aU0XnAugV9zRDhdRB8hrqdQtp0HZcw8RJMPofAXeUEsyPd34bKOf/OfiU0h
gU88mBpZpAdP5wPVrJmghuEk4IL6IFs6Sewtskw71DurnHpr8XMb9EC5VfVte3og
CFm/y5llk+rfkLgFpEVUPAxUXz8ZmWkaKcl+NpX/PfGz/8xHjhA3RYR93cQfHkk/
Cre201F8WoIyW5GEuCk5dM/7TDREhOOuEzUf10o+b3q8qfhVRtKTEKhG8t0YncCz
iD53ZWKrKVRYXGFN2P5f4IugsJf+zbi5U0ziUME41GFBzJZByl6EpMF0o3++5MxD
xUP4WE/xjm0K1Vsb+gIP/P8VrOOKPICI97Z0Hp1dlfSkAcaNg8CyyxA494pEvYpS
wlU/YPtj19O8P9ghg5GXpDd8+lcmUes56ujcnfs0yO4AYOhq2yX6ivD5Abgc83uV
NmBjS9oRukVzDBuq2wPzJeQmnfPzL5f5T92hus52zGXJre/w0bt7/xvfHlODT83z
rFgn7RTCh2LLWORtT6eRr5cla0yTZm3UUPGg6pgcItGxpH9Z8jbZfZbSGP7LJZCV
D/ixSYZv4eztRd0W8/3+ocYTT99+vLwHxecYMIqsTxcNvtUgFQobn7cm58WZdQwL
Nx+igV0yi1TZm2SYb+I1JtjYq0Mf7/dz9ANayWdMduOR5cX6jwURs6XhvuEM/+SQ
tEmtYYEmRcehzU1htsI9IKybma1kLI3X+huo2EjghjMyC6eHug3Xb+9h649zr2Jw
/THhNqEsVzI3U3IyKQS8S5gkV6ID81yGixs6d+xR7yoDjZT7rOEsVwecrBiA2uK2
y0rXBPpqRleZUjVjN/A/5TJBJ4jUiY1q3LytRDojHVfPYH9QEOglzEaY0xgpgYB0
xEpCBfTxzT75ljBLGot7zM6XGlcGkJ/DN7pilL8VzCpKtD02LiaWlC2l9/WbDn/I
YYzozpldjDivutoEBsrZa2E45mRC0n1emE1D3CvWLl1z6saxyh2/1jk/LZOCsOOj
yH1Iy0iwvK6ZDwIobyopcDzqsDfu4UzU6KDM/XwDemrfJGe4y2/xH8HAd242wxeI
pxAoL6cZSyOX3AA86M214SzNbwNOjJz5HlVxreH7gywFl5YCduLogn7DQQqEXWdc
giTU7HucjQsOm2OUlEZsqA2kZtbylV6jhJUspxM/RPwppLl86wSgSIw2yNBpzIcL
5eI++BxDepjg9wkJhg0cwWD2ZtLLypu9Ld/GFhghDsecMUTwPNz/oE1FzLFRu5Vp
Cezuj7e4Bo8jrGdyZhUoJMQZpvQUXy9f0O0dNBOvAS3651CSx0d8UoKdFvQZqvVR
5NFXsivyWDncPIOFqXXcea88SdftTzla7BQMXPwfB7EwY/lpwOqKBRTbNPgd/LJ9
cyvM3w3xxzFNQw2i0idlXxl8fYex2hy4zc/78OvK4CBEC9DcdFc8OP+U8EzodK3c
cKSB92InFkWXIcjnlaC2KTIJe8S6VY0BRX6YTX6XN6XwiCtQNKdgxPN42X6rZ2BH
O7XtUukMl2Mqui4xaWmruz2IhLokcdG4YG1WuFOC2nItjnVU0iRel7p25BvqKN+m
3oRxvZEVKyESwVCC+XeVbYKMzgNJ6fB9wBixcvxpqdbrqUTD5VJYyYUSubY/aeon
uwFOJlJvLesvwkhjjHezRAGjgFRcmf4n+Mgx14VFXAmqs/mqxwt38C2d37JiUgmH
D4LqEeOP2KGVEMuo+AQ5mFfZas2nywoM1R051UrBXO3YV02GJ5sPV8JeWjgWt+ZC
HySkD4FLnbeKWvdbwiT51AjmY6js+Lb0NWTbbOsweotoqQDX8NdLyhIkTZWn9+Yt
/oZhdgLX5Rchu3IG/tUIviRjBS0xvCaah1LsYRqPQ4VHkgXwTJTjyIl+daBFvcDq
e+cdO1plA31fnJBCG/GPjMgkBKYvvdZvql0xRfzdVgbYAn+lHAw/udyYaKxurDyD
uSA7oSsUCTtcvClQqTjr+rPiexScD4VB406rcYXseSeAM0qUtB/nInUFlJIpu1XY
30E88bT3QBOwL1jeI1Osv3iGuCAhooJ9PTd6AkVbw3hkPphxLu84OSbidkh29Zn4
UWu1+U5xMzmZlu6Mv9sgnvAkIYJ+TyLcbXgT8s1vTJ0bf8WvoWZEIXGIq1o/5bCB
95uYndK03nPxcG9rZoUUW4obG53T7XFZ6VgQ40yj4NJZtETb4sSiBSH5anHki14O
LKPZZFbwcpQfKMmR4IkTENzCe5xBYTqCE00t7ZdZ/mEQ3BP/0QIxPoXGcf1saRO3
ZPqgCunmbAQAevSq2ALkA9UeHu1m/GpOxONAwS1zESsOh2uiuMO2xN6ZslYM9zM7
AXD9oFXL3mxJlvcsfR8sKbBR5v212p+DlqLo950QLnZtWRBe2aeC2XheVwSIhcy8
Utk9Zv0uKTK5HwOEn781Nb92qQpW/ixukvfnby+0tPXMyDEeZRj96wztUS5dAGkc
gHqx2cqi2m/tNyHzUle6Syyr7wUU7qlp0OywpWdta4SgTsn7QH0FdSxGQXSRcvxs
/ZIgTN7YThTMkPUqJn71iy93DCR0R6uKVBEx4xqWVCedV9mpGxVU+euxu/b4QIFQ
l0Zxgs3CIdNwwhxRS1jfySbAg+7edinzo6kohP6TXlA4crL+9a0mDOONpfaqskWo
0IqRJXR/E7Iqei102BZeu+SHsKKJmO9ZehSjue3zR3Ik/P3JSKxp0bw/leNt9s5V
uZjamPKCdoexOu7Bq4ygLwp0z8uaVH5aLAvnPOlqIK/s6fbNO3YzgGA88kvc6CRD
oHam4R5RQ1VOnGOZBzQD5SxMHBsxkmOKIsRn4PSnCfdPnejR68vAAu4U+Dr0UxZl
UJ4RiZUPnezXnhlTWQXmh8ifcdp9wLopTKiUnYD2bUbyjceC4Fu/R82KZ9xg0d2V
fbVUImrQvEkvhSkc+2EbL4FMDS8ptD8qJz46GlpVLiDkKdF7gmxI8M1VKTg3mV++
F5SLKbkxvYr0aHOf/tsEycPJsEy4JLgtGPRoylI5GCbgGAQ+ITyPr6Ym8YpFY+3A
Je1jOg2C+yiYWaNSb6P8000J+P3YnLV5H8WXeKSO5xZON9SLctXlYgKQVLo6jhEp
wm9yRucyWkkmBHDAEajHlH1NO8/JM2uhTyucenXrmJqwk8vMzqaM7TStWENBCjjj
fvqpV6K+3NFQgG7r+GkcwZhtydOmq5zdcKLbBQBCZNbPhgVvs113coSERufEy0pj
i7f+9g73KXEd/YkfifpPNLEY+NN3ldD6pIu7TNDsrzhGGRW3MFUHLEE5TfoM19S+
Zjuhhu7VyxIaMQqsLvHPOFfDWXhiNt06Hpkf8xTkW0ifGOh3GmHQSdmtz7AdjV/c
xIdbdbK7OzHKKwF5iJovpKB3l34VJSvABU06CId6YBJOMIa+iWlILdJngTXA5wEd
x3vbys3OdlemjBur12HaMJQ8iE631cEYAUimgG56nBMqLsnrbVmPeuEFjp1TOhQe
025thFlpiYPo5L+ZoUy+uTkv/YzO9QWHNZ4bpzztRUd9WGA4zVvKenYj+fm0gdbH
N5hQLY05CBfWbHl9u+NQsg1GljdBTmiWRQHMoyWGvKZ/85G1PJoj0uJu/3I1L13b
BQZCyldWLy10K879LOsdfLrmWPs2WbNHFByjxpiMN20zD7+vJrIJF2UgrJr8b4bW
tGcDn5zIRfUZG5O1d07FsB+fllqtEB8TJW0T6p96kguojrP5baEbIJBDMCIrzG8m
u2tLJ/9ERwybMISFah/qV4kL1hCLyyv5mHR3djuIJifVCPCRXj4MP7Qu9iEyJLwr
qePFbpNqQS6o4qfE6XAMSNfQEJ5+PLF+EMWru4gWN5gfuFj1riYyolaDimpxS2Dt
6Cwl1KTj4vRmB+tnnxsqbCMoL8r/E6uLL3RmKvpX01jGw9dBbbyHTA2c+P4UOVov
x/Vgp6lT8yjxzclhh9dFwwtg2FyR1//djOHW5/ezX1oDW2O7W3IOqDhz2B+gtM1F
cCvyhNhG5U/sXYZ7loAp4BcsPssRFNswAhnAFxEwpR1Tp0W4isxC9+FeN0BzpW4E
cby5XqrtKM+ldVbwiFRBF3X7ruM5h8XlgW/nGA+nbsZvFZ9aoHLok+keKvFYq6i8
f6g/Lp5ZbapUpbjShvb5xtJ7LFCTzu+sui+2g0xco0SLVZRoExFUCIxPdmNPBnvk
mrR/HkEUmZH3btYaYq15CCwzrrQNKrdJNdngwBPSIb/IAbVbBM3x8p5U42LFgUPb
wUP3FZzvc5p71HYBKCXlDbeHj9dZuzytOk8mzjac1d4h0Z3qTlRLnQwGoHyKF/Qg
hWXNvYriTUYoQeu0EGqBKbAqbc3n+8ttkHwFppbCodYh6QBEvYH4sREx6G5nBgn3
4anb4xnRaLevHtu/ZX/2XBSKAA0tyvkxg4sPMZMZnh1kOiurm7sLly9qUC+NBweu
3r2gI/7G6c5APzN+2wmv1B8fFVCCzlSHPvbsLIuxQEkAF/eRQ4kirGaJQiZAl5s/
jIXL7ZDD7/hBrSWzR+A4cVulCxzuhFQZC4JwwUu0LgTYm/c0kaQsXlA4RMCLPetO
HHqEEfG7MMvuovbnsetRU5sECeo6rrNNVno6W0PapOfiP3HlDh+SSjiEh34coa1b
sNl4cIwHUFj1zMzQW0sxX1jV1R7aoS4844jQIqtnhWQf8jLwwfMe0w1k5+569B8H
apU9fMIP0LirSUgJj2sglhthAItynM4N0sDDdPSrdKujDLkpgRExe/8BW43GyDhe
no8a4mEv6MDz8bFInzuqXv0RCAY2P3lxf0fPwCvwVg4VdRDuqALQi0RbhZQ14jrK
UbvvSW0r3Z5yvQs2DYUefwFhDAIKRMO3YrSrjqChfSaDrk3WTSRdKyDFddWysfKN
HmLpFFBeThgGIQz75B3YYWt3cWeQgq4akx6ELcJcT0LTfsNKxmQX1MoUUhlm6SOk
FsV6fxCNyUsyXjiGCDeBfL5QWpI0ZlGYD229bSYnFuniYSKCY7/uht+8BCvS2Xbz
nMd29o75z5sEVYeZp9xi2aUwQV1MaiekeB4VYUbLeD7Swq0NyzifPeoIxP4wpGip
Is+bpDn3JbDnMrjVf2Stl1ICSCyED61e/KUt/XKLgzvKnBiuazt9N7PfV9A/T2wM
Q9Pmlth9hj3BSjPxyIPKxISHir0a/DFQwUv7P46/fUz7OkWbuwKBkRa72AWfKlRK
qYRwusObsmazLyIJh8pUNShnVH7QmRLNe1M9m+yXHyZk7/jymWbZWQ7wX8GqTd/k
dw6wPUnAzsDSbVEvN7MvmzJs9ebu6bHVat9tBgLjQSpGVQZEv1BeV5Rr5GuJQILK
eyh6EaonQMMhaDEBGnROmfYUtf0AB7P61y7vVamauo8sVH28/EABq4SyZmpwjqw0
3HrfRQoS5+D82h9UKD9/cZ83LQZRlBfYCF8Bv4snZb04D4dlsBCv11DZExBL8I/p
c4U8x3dY99g5Fyh2TbOyHimzZn8aLyCChlGn/AzvKrLxHUkU81LZBvCheymQf25s
Al+mEvJnEulG3uTFp0GW9uWhJ0ZWHC4dSVu+u+KQGVv2CPpFLTA/LEIzA7oPWvVb
OzA4xBcPoLnWs96J8UKNEgks3tbZHapdAoQYzCQp5GPbrG/+qCTrk1At09U6LpMc
kfcBbQSGnc5fyMzDe/c4UZ3JACjTfcEZ4GVJ+3e6JJKNza3UjNyds9fmOwnAZ4wO
raw/chpGFpKDobvERTVsfb+YZ4didfHrz2g9oGAywOxdaEmbLXd0Y3trhzu+XUSz
v33d+1A4uQLWUaBd48gnfZZWKgb0Y4ghbeqG4BO3jJKZkh47USXwHnN2LfbldpgU
JIBOwcE0exL/TyBqLZElRh5WMnVjD6iON/IVEZRk6FME0Ipe21lIQYBB0UnZxnZG
dbWIQEu5FeQ8dxq+GmnKIAHjXFxNmhaWxVUyCd+4NLTBepE/OB7S47ZhbCY/9gU7
Y5nBdeMsUvP/9jFYKJuRuC/p78A0RSuDuwOYTkmL17ir9VsmmM1geSTU61WsRM7r
XymFjC9m9QGI9OwAnfWnCR+oHQlYbJ6MjaNaXaCIjjgx/X9VxqKtJ0sW/5lxpDcw
KpaA8x/sC4GNIit5rhvACYSHWgli3/yfjO+adaadOar42ol44hSlGiSM9FD7TnRD
GIz/ONJ4MLqWA2D3zJDS1ieSrkT+LvyOCViXj+koIQF/pIvYV9EFN/9pTVbJaBpy
2KXDc1Qz3VemjCwneQMjahQKwjs+M7rMxsnGLLJ9MZ1VKvW0Hb/9OVskWKjnY23d
M9bCuP9h7sA06MdMeMf7LMP5HIPomPyu9sVT6FuqHy+P4ugwOT7B7ezTf2m9tenN
0CE2rgrFE2FxTMlRB4rVKGl2NiZgldvVQAfliUQjCf3f9VOJRSYRnwj3S/h9eFFP
K0BCSpoCmLJNXFgjK5Efv2PaEu4wz29rtEg/+iGex9iwKDCYzZxqdNIRr1clflgM
z4XeZgwNYWaEYT2D7jfogg3Qhdo8j08s6unzrC/UXZl5usZnu4pFUDkBy8lmRYMk
MtgkWGJ16A6cCOd2EfUMwV0Bv+W7/PTdlNHzIvkYQURl6LfqaCmYxd4fBEgMvOGJ
8ANQDkSC1E+iT3ZKUnOvXR6+OxjpnDKoZv8PBOANsPgl/GAr6HHbF+LWQnV9bbxb
99wiyM+spuFZ2kT/Znw16nA55oSxywc0MoBmAFafLyyaIMExg7bnDnVlXrsyvwBH
V12AyjbRPTiAH1ToWjX+xi6o+7zgXPDQVbglAlO2Q5hjqtDTQrQLW9ydbOwrxy8/
g+SY3IQqVHu10Em/xY4YUHPYCLfzl2M2ipw3zlp7IE2adQTBQJBhOatZ5pnhcq7k
yf3BOoMJtk6AJ5K4nYr6oGeYW034lfAu0ue4hn7ik7QN1y7qh2uHkeaoNYBpGMml
FeiUI70sB5Cj1KOe1rhACaAnA3/iYGIMFKN5mpeF9azzqny7wSSRZKPANkFzMb16
gNLAWdcEdcQu9+MGH131SWRDbMAGbbc0HPYqkOBytNAQyzaWJKaKf6bJGFKh4X2R
XdZDbZpVPC/wAxJxUwsvk0B+b0hYHhcsulVfeXlLCTrs8uC9/AJQx5wONWoLVlQ9
UrZwJWO7eTOyPoyv6fXxdUTIIWd72DlJDKCVTOZ09uA6elRU/bROGgK4VFQ9ekMp
AsFrmWh4vZXHQDdFDBB3ql7Zlb67DbuSQrfbYZeF7Wy/Ru6ag3rj673FlJEF6A5Y
g9tDK0rY/5IqvdNpX6V8gCx4d1PLtfBv7kWRQ0dgN03+30sGW2O5/Zfa4ZQnm57B
VglcfsivPe5Ltnk6x5B2awsbvlDoAIc07tkdDRQfbVGSex9x2VLugR5cBexhV0e/
rtRLYO/bg+LjUWX9ecQ7zdf1x+5XYtcH+eF8JmvgR3K60S82t+2QHe8UhiGHD2Qw
rrdJxETQPo1uZqBWy+C/LNON8h7o1SwTFIM26IEDAfW5Fdb8veNE8d8Lx5lqiBfw
VPhi0qKPr4hTf4E80Jb0mkDtG3JVSF7gXlRisoWsUgB+P/N7tCqQqn0+1AfUkYPF
UpuKrH2SEa8vseApmNhGoNPAP3bWapbuKzKA7pOTDRz4suroevCBodcrWljrg0NL
CrS5DOlaSXDoZrqEPB+eI1FXTqBGLbb+dZhC524s48qQH0Kgypdz8Szo6iDFAhUd
v7YBtieTKbbFlrDWJJF1mmYE9NmxZx2w2eDkxB5QFZRworaA6twhYKx122QlxpSG
2WUWbjzMiAXe4VJqGzUI31ey0WJPYTDOCuOEfqFliHRD8sKqgCSJ097WEf8koRLS
b1zGC3UY9Lu8H1mUzwkLOgp7dzDOe9AxqMbbmYX/d9O+trY64f4cbp23n6EuXdoS
pEG9acPc9tvBbqIaH20Dv4Hf0a585wOeIVYiqpUNry0BRLdirM00NlYzssjUuQQV
/51FxVNlTUCPZX/yLCukizkftSaghYwDLKTSC/mr4eHybENog+cc5VORytOT9DFp
FjH/xJZiDVaqCIlurUUFzMfNa/+4xB8X9TZ1Tmi7CT2f7y7Rk7XNx9+/kFpIT8Cz
FgfLMVtF7JIgv4mCiQDtQ0NHhEvttQfVwZ7KNBftzE8hoMPSbAzKRNxgXXgkrfqp
WrHr9qb9oqjxckD4kgQ7A13ZVIRr47bYco9kRx0Feyv5WobH/+ynz8yDAZvyolta
v290V5wAo1ej24NLOMyI9xc+hgov6STgJXB7Q4yuZ8KWS3VieqNYRpd1FowWmDPn
uV/Wi55jHOX6DQjk5zxWHYXXAB7J3a0bhrymZBjjr6rDWDOlGYjK7FLV9BpejhOB
3bLsbpVWpnvj0kVJVwS43d9yQIj2YfNKGPLkUz4VJrlpeR7uyinOYJ0H23PE60HW
vojSAF9CiFiwcYAp+cfaYh7C404NYNuSuF3R+KtKdU95us8F26DKwyJwKF2m0urR
mUQjhpJ/ALBXXryraumeOVuDRstEnn7HOqceOWUII2lLZ728/RKY36Z5BDsM+i+O
ja8aVSC9AEkBgWSSceLZLLWehv0b3MMclHASnAS5YgStAvVFIqvHw+SFwYY4OWJm
eEw7cexGKG2w3qRb5AWqV3VE8VqLaXXv1w5xMFmW3mayLG6a6JLZmXHOurt9Xq+V
xPJVu8rkm4/gUlCxhlUSRj5kEdNSSuebzEsmiZXGf9QnkydyKlqfBf8Oy/OEF/Mu
q0yM6nuIVnDktfyzGls57Rz+XgB5RtKaFHYRIcDtz3KJGx/UJSrAKLP3DR0lN4V1
0qweCQEuj4hBISh5C0lsyHFnIQZVFt5zTNWK6yJOFoRhPYpKP82VyyXvnQnWRmiF
UWoj2KU5FeYTM1N9LtvXBCx0NBnosTue6CRaijj59a+/6foJefoqjwFOfAHim6R7
3OQpIg1lJR8MhUmLjY3fa7Rb1kab+vNpxJa5cm6XY2ziSNMbF2WJbdeEo6SVbWSx
tdfioF8prNDrpiL49kVyP12QwZZPAzJPM/yne2uVddd/Dhp/g8zIgaQinSE4ClzC
R+NP7H2kc6EkT88dlfux/AWb0WsxUPmqsn7pX/SXgfGLwoVaQkp2DG/Oyo8dQDe3
GDVP2icqE92SRSiRb3kSqmSV0C+jPUWfmlgIBU1hYlh75rMLFFL7Ly1zjg6Sp+ho
b5EMgbuJ69ftbBoWovglOMVACahwPD4tdsbbSX6wl0N1jPe5xPJpGEk5xP6fITso
GFoHL/l6wBSJD1K42HYKWFJn1VXPYazKlqyL7ceDvFXWJqUc/Vq+haWXiFxbbr3q
1dQP1lQ0iPUm0KTzZ4oEEhlBEgsfYeiBVXUMgE1Zn1ddqBLeemU0ker6OKZ4Ckbd
nUR+ddWbgOAhTJAZ1KttVUbQ8UZ2iZdps11smEnsmgeo6efEwSG/RONJ1DtHlV/L
zO/ZhYdKUjfYwwPABBTXuDLa4SpRL52KpBxHWihVWm13Z9FwD00gT5IDtV19s2p3
2wtykvLPbf0/KieOVF15wREukdE1JH0pYjKXoEeog8efWps33fnuh3zI84NDb7fT
9McflxXkcgIhcoMtnsihsrzPmQrtQqE8ar2fVJumxSL5l51xEhxiPMBmGgbTXHcF
gIIz+vQ5n6Auv0Bmymyj93OB494ewAqmoHvDWjoz+Iv2+T7yYJVaCTSU7IsRmknw
NDXj8QOq8nW5AW5yjqGzla1TMYHXI8o0d/FIz/TPbhCn/HbjB4pvhXLdQ6aBsXrd
ppombOAeLf0DkFX6fCdJvGRAxbKgpD07RoxNnju6dzoQRFt/x87Bl9bKCm3z8+3k
XQov5mHA1c8ju7PvVlwmKBA5m1K+15RfAYYTYX5B4WaYNXcjeNf+9UP7MXrwFWgQ
8obnh5DinrL5hGZ89MYRZ+DCWLq7Kq87QXOBkiUxZIoJT69ww+6Uk4hC2JFOlapD
vN1nL7gBjp0RjB6g7jjGYyiuHmkX54U35i3N6vB2Fx9PJVIDbd3A+WU04YzTgFhl
4z4LtD6gjr3QLTXvv+8snWzmYlyXByar5Ev2TiXlh/mUFUHtmhp2sgSXdG+9/d1N
i8dLLTWFITKu+Sq3L9TRLLEWSnvm3mmTJhAp/CIOcHGu2WycxMPrG9z9qK8PvENh
MjLmflSjTjmT1Hp07z40951E3Qs76MRMUTTRSIpQ95tMoRqvks21MBjEFI3/5zf1
nyu0ooZ3KJbvFA6Vg0ItnY1JsqtM0R21/IkRxGaOhC2QdiJZZ64uP7iKx/DR+DEZ
Qbe2wrfJiud//bu19sggOF+Hq38HsFjXb5ZIXTD08PPZ0EJSAy3ifJpQ71F8KT/y
dwL4XRjk1Hc9KD95dDIzdVd2e0yetmWf+Q8nPiKeKnFeZUaLWj2wQnqjd04DXJiF
6WAdYUmh9O09EqrRL6E67cwLOyAedv7gJ4/0HfaQ6NQt5Xncr33pjyJPpAL0z8sp
R9kJtuQxc9BEeEX7TtBQ4evCkaa8mp5Ch4kjVdiBj4Mhun5O15LnjyD2G2/JPl2J
Il/2FC72GeZZ9XKGpT/0TUuh1sWcCi84u0atTHFDouqfyaMPT03vBo4N91e/tHJ9
hCq4n+0UbrWHXBa1apvGq3Grbzb/sBYKRa0YV982H06cOWZxmnsyyX3ofmCucKFh
otSLQhpL+cWIrIu4aEUrGi2g9EPJBYGu21cHmcviYV29jRgEnUT7b0R+efxkGI5x
IXORlURlsUssLucpdjbGszM4U142gVyNEYC3v9PbE+9DSgs3aaW1EXIoF6fGXoYr
shBivi3wCMadMSvjVGgLIwQKocIObRz50MLGoVoLPfvEh4rX0SARVe9+bMky5Kb8
QDSrbWsb4FfojsjPREJGehN3an+Ekmtqd9t+CQM84OF5jDNFHM2BqS080AFT3GOZ
StDyODPRx5wV/P7OlEc1L7ZLdBMOxc9NYG/kPHSvEp3376yX3uLEh7Vd0rI+ptXm
egBr5WhXhwTpZ/Cx1iW189QfstSlclBeQRhcxZV2E0sOCFRtRo3qxyB0e1iShjBL
aQBaog9s/fMhIert6SxAcn5k47ZiGMI1zhJH7ZhX/VVR2obCdUmvsFqJQifrWeyT
s6Rfboo/wVmIcCSg4PYn9FB742BX0NuKlwfmweK8yDpBL/1T2g05iHxEpunQrPxW
MqxGKvORtyICh5yIzK7IW/PNhTHBleKFeaPjrp7IM136hD8n1kKYMYV3MfSV9YLy
YUixHl6QFEbW6QhNIskQ0lNqsigPze9tCAc/MNdr8hYtNeJ7a/v0sfiXMwPY4OhN
wCxfBbRUDpeEKM4plCCTfOBJjYgg1lZqprNHySvoO+ea2ZbTxTwHFtFWFQm8tln+
vqNWkbevGTl7vjuNUivW4xi/rUZyZYbH2wc57t19/QsqtVfE0Wi9P5Qg16bDVo6s
7v2F9YWVbxUOUgwv8O5M+NcZaHL+b2x50rT8OAMtp6g4j2nU2bP7D/kmD5uemakR
W7n52V6oz49TxOg1I18Cw+/GFKFb9rnTwJK8J0ZeWbtvKjzSdRqObyO7WTbuRTlZ
G9q2j5YI6dYuBVizvnM2wsTT9ByoO0mOh2//R7eFJHKNGE3+JY5YWPyhp0uxR9jD
6TOQPlaOsXHLIKNB9nbKbMacpIXembMp1Ucg4rh59pYZi851Ngp0oC42mv0tjJ6z
Il7sLOJ+p2EvLlzUFa+oTwJPodHjJow7wJNkNriCGHTfLmaQHmEYP7tZutcmRoBZ
D4X89mPXvQ9ahjf0uSesa1Kbn6TamokEfEICRUB2izbcNKSQkcrLL9jiR5F8vAfw
3Cb2hXO+bBKD2/azOZjrOjuHWhl2gpFtN07YJhuYyMtNa5pmZk+lazo+GyxtUFJ3
NpURstrcsCFjn/2o+Kt5oulaW8Pch2UP3qQA9Ja/LAVVOiHNB26eYiwwPs5y6Mdw
REIl8u9+hER7s+RvZui9eo8gndg/KEVa3xq3Hk5tKk0pB6D2blnn+B3IThzWRQrL
M0lAQMhONSjcWyOf/gY7YkJhMexvS8Qc22e4fpLkYcHJVF3uRubVi3hB46ghDXrQ
2z26lwhnbjMQSUwmgE/scL/X2DMJ0U/NlP+ulIb7ZSqoCEHMmn1BpUqYR0rpYa5R
wEMAORtWz7z3hMotAvSfKky7soko40VojPY79f7ViAj9eOQDnlJVRbGpz4yo88ax
cgb4WIL5ZCKROzYCpO1nGJdBtPH6jH3d7tK0JJKKW1waz6jvejToP6orskFY+uOS
Lw3u4n3fT9kVIkOWWVHhcKUiDel7CcUoUD0RC3tgqHLPntDEpeN+0z7yMU1/P9vL
7NbvS++CSfwfrcpgm3pAto7ctMUdjlXLhm55ramMH3iIITOGYONtWV9NSyx6wxLs
WZTYAdmPTO/pnFM6s1II19utdvyYnrm6XiA3ujIpvJ5TDtJL3JPQ7R9W4ehA4rYX
x/DGFj08reP8Hc2Q2dO0hmHk6t0VR+lZ3G5nkpPIZ2cW8CREH7d9nk/UHRznMIBU
MyijAlFl3gpTuQyJ+G6eXL/TOjX0O4jugg+ltuxosWeu9I5RJeDdq2YnqPgE63FQ
C/mmjVmK2eu/o34Pxk9RTR0tNT5RlhovxNYRgCFJ/QVdMsVVjmZWaZKTYrr8xoCU
gs/5+oK0k50RXSCWH6ebVbHylmdWsK8OnusgzYT0hGhyHeylWXYwrK37n6chh30m
SqDp9kEK4oBQ8rJXjSB4SWQ0Nq3isC41uNLc8dBa9SsRILTiGsc/eGLOl5JRewjr
Q7tMufP+BSUHn7GajpipxA00sUYOfCPWsCMQB18oVaKMxzlPG40oOYaa7YJIY0zk
mADQWkDsyi/kijfFQ6eUAJ0F8KyvYp3TWYuEtbgYKYkkE7nU5VHsDsfHIi68lxB7
dT+XdXXtyCV2lGJOZwe5HweL5+bdK8UARgrIMZrxxJ+uTM5wLKrfz6UAt9UQLcE5
pCLIt10RMbw1I8E3P/3v0i+KWVQ53cSK6oNOFtT1uM6vZZsyDbGFRsb+6X9al6Fu
lUahwARdt9o03mSdMgiisGUeEXbfOszjLdRAUb9WUEMnMWczgZnypD+xfADnAIB2
mhHqObYpBuzlaSbCZqs0WD1hXNuZa3+mEoZgVMJnQCYbHtttctTd+o6yTIpSgQ4k
3nRkvaLk9aPpzriQzjV1rEyIAf2aOKL6DianwXZtdqSerz7EU79vouhlNQD0NLus
UCwAR1L/ncAV6ECKnC5r6OJTZmK1Y8x6Jb8EHRTyfA/m1F0ph9MAql33QnqJ5Rsc
Kd4tmRCB2ovPSlFXmCXREqCnJrnP3F1qAmNuGh75L4n+l1zmsFJgRN8hEnq3Jxvw
7K3Nz9So+61CSEm4eBR81MdginiLvADMyg0pW6R5qam7gvyKXcVYIo9/cYPeBa0l
7IvgUAL+JwE1g6CtjJzVCWTQnECJXGghfZboZ8X3pUU84deXrd3V95BhXic40OgL
dM9sW/VAeoQmbFfPevtif0/kB67mmF3HW6nTc3VSKWyJBfsBFN/xB3yaPOBXi9XI
ldLC3spOrZLshwcs4kXSwoUGLvwcy4HNHvwF1tPk64OhaWQsZovb9RMHA1/qwEUA
jEVecR8uRfXSTYyw3Fnupeh9zfy8efhWjrQRX0h06LUqyLMLbB0+zW9cpa16fr4X
0FDjLUEnyaLBa0lhpLjjQJHP34kLuaEambxZL0tg6Sm5DWe+1WT0S89tQ9ABqmw3
xJsKyxEDE70kD64SIFot90VrUJ/8avc/9hQ8D8FKr+2D/CKb8gcPcnfuQ1kEFXHf
edh9bcj9DTQfpsDrnxbqtVeM6+7CXKO/Gb90fRXM234IdpQqeCVMZZ+gHdbcm6Bk
NyTzR+cRyXYBdAGEDgK9cvS5zQFLT4x3x/GXJC9KPSndTnnv5wxed2rIs5e5/y5E
wCnRHi4Sg79WBIEDu+qyBsLLaEqMn5EoQ5EtNNXw0EX9AOOHLQ8MWjF8wdNkWCg/
BaVWcCi9MDYJGQpx4YrukQFizosloVt6zMkVPYadq1JTRTOfHUwVcpOdvu17nM6q
izNno9/Hq+Q3kopUD4DEARBXo/NkjgxFOS1a3un2MFU7sik01bXJrX6MYb/fIyRZ
lQpa9gGyE5MRzlpcc7TSdvcRNOxdh1Ail0RhZ4EsTLwPJsSZz26992W/7mchyKBD
7Pjh5l2isLTNsEthW8gZl7gREo4bUdoqQkibzOsV175f3D+mRq0IJNjAOa8qnktj
YWRU9QefpLSA+o0cbCjeqgZnAb1BOPI0ye6L4ay+bS1ZpkHYfp6KhtLgVU7W+kxE
n0NaK5sOFn4NjTzgP10EwQahFtE9CrNBFAot1gCwq+LcG+rHY7Ox358i6Wq1dxSG
p2TUJkaBY0M9XqfDJgQm150t0kp0yWb9Yt/a0aetG4x293/9b3RYhudGMqT0lQCw
GzbaiYO3GdD7Qb5IbCDTI/2vAuevQyAy6hvk/hF32xnvWMO00b6Kq2rhbGYhNGlj
z3ggLguGkUwpw73ctS1imAWqts0HFkTFJ6O6DVYR4agXsZAZk1KAGIwf3P8R9Qxr
BAWUNNhyT4LofObVl44JHxQw3nLUdyclylTtUNJdgnMvvtlM0k7P1IiOc+nn52M/
t/hEEGF9gguXcIz/m0pGaIc95RF54poDpD7vpf7JqOxadw0GJ1mb7LxiACSNKcDU
8ph+Rw4Y2t8mOTpmYKTn1NUrXerg5L5gEUVxoY2PIZnWtJiDtV+URkBXK8Axeo9r
rb5uTtmza0QUfTTPis+YGWEpB5vJg9fyuYqhXcT17R4pLp/qBlhMpuc2w/MY+mLi
qpl1EwS3OaFzOh+FZUO8vcif3XsVcqaIgt2SuffFVCqTic2qA2MjRER5kDXY0Zt1
dNHzG2LS4BVePpsqx51SNc0Rvk4EzdqEcc86NTf4cahdOx0eb9Y/iWPeKF+m0zFF
Fs+YrzmNpVWzuJBwcCcvJ7MIu2/bJ+yavjVQuh+bTfZOM0I0FuEJnIB36Yvj2AQD
Jsl4W/rn9DjuQiUr2OFI8ibpzKTMiXrEIQWiVSdykvEePaTqvGYQcccHsMfG/lSt
+wB1+yDdo81J+V7TcRoSYhv/XPPQi93zJP4Ifu0tlf9o3YqMEXouPl/TuAYFnC5e
nl6/348Ca7XUP6SSUoeQs0pyew+jdCpNxXL2qI9YgCJi4JhTfEBLCVhN6KXDUCon
0bThH9WRdzRgfsXZnjCJifDuhGqvAuUSKSu1twjBB0I1jGCsKOu22iUBl/VlJ4GJ
PImk8Ia0DSCP06IW57bNcpXJe0rRHhlvYHoS1GU5p5o0NEV+Z+9KDmpB+oPxQik1
seJML9P2kTslhYdidzPTsdhtof5lPMitDmWcVdNzIC0m5lHXxrFDdWKwnf1YiCJh
L/8+SJfL4kitrK6EOxBqhuM3Tam+9We7/rEknC/YLxg97PL55ClZ0Gaa7qr/T03e
RtIyoEoF5GJ/DHisNrMR+yVO8mfWRz2cklUWICQiaENgkevqyyYVS1lVReWyWnSt
jY65T0g/Hefnz4G1hQbZXeh1CCStNNFRzG7O1YuVhA1wRDS9rfkF3n4esf0eDJLe
9f18NgrWjXf/fQMfWspIyPf1hAStkVLHLEXzhWQnlaaIYnENG7YfcvJq04zXIPSG
5OUmEyDun37xGq0tvjX0vNBYYtTzIpKYwafKHz8XNpZJg7GO3N46XKmQUZB7GQ3U
gS90mGGmYRcHzn8/xGUy9MwlmOEZczpo1ygWRhl3oJV3PWb9XYtZlDJ2RhAointt
QSqq6XQ5KG3bmTQOklErds/tgVrp6Bzj+pXGyHgnGI7BgHLJm9JPop7DqsRO2gyy
5TYyYpLw1mr85vBFIZ8PzrZ54tmcCpSVbXQfW3o0/fzkgSwQEDgx6FZQZv4wWW9G
txb42DHvQq71dYw14f/5/+AaFaRY+ol8OB1Dk/uPLknt96H6tsgPkK5evlNxWwwa
EsEEUnTI4YwMDDO5ZwJALgnfkAdX1lw1Z0WcNUtoQKyyAig4bYJ8XLPjiP4PyJ5T
ySwqFfg7jSnEJB9AA1LpOjwg5r+DJNFuz7EXNcG7td91jQw67GatkGSlKwG395UQ
v9gMbrjD9DCc93VkfvD4cGPpT/ZJEx34e/SrP2kKuiwea3GBtDRpw5ZZpEUPn7oN
9y/7YDY0GEjg6nOAgvi0PgLatxBFzfveLOTAD+7cOB0RZB8YxQ7Mp10yIoHlkq/1
cZW9LEzJIYbBApFUaW0XrdHeiJCjJ+SWsX57aQmGaMOrN8uZbPf8oWT95XEjWeMk
zc6Q5sJy77hjKBRAfa7KArp75Hr72dt7+HELnMgUEGItSu0xQ7zEu1L7Eag8/BZ2
6zs8bFtnn+QJs0wv1baS2BYoEhGb7AXjETOgEH2/JlO6l4Ir8vjmjK9NuAsMkXFI
qaIhvNFkDhcjQenD4disjFYqeB8mxXVwHt3temratbTPjSNJoyMBIR4IO/5rTydf
+a7B1Jp9Ay5nFpe+hM99hktqPbitmhKai+K54d730DhAC2qGMNVIiKQGpvgnZHLh
nctxLC36844HGOkP3lD9YFWX1iIgwJcMSfidzDpYVI3kM5pY7+6VDYAeg0Df/YTT
3KGEk/XNjj7X/I8lh6eV5cUMBwxdFcOTvIHWczfe+0nBYraFWJUitcD6YAGH16SK
ACrUc+dVGb3z7XaPdybJsXiYlBPebTXZ+OdepsGcA22lygIrWi/mnb7nbot6quUc
EqqzBA1VTs8jJ9fipfkv+xrlSsTkyrCs6/oWW4Zx42nh+dXgU7sp5h8oJMKkz5KC
hX5Nu/CRgAtNDH9LTaH7yacpaVrM/Y83VQQkZ9B7TwJZvM9OK8P6SqtAeRvDCkFj
HPZvMM3BcORhC88tL52CDGlz25tyaJf9PGl+iDAiGyW0FYFpwnQiy4jGcbBrKSr7
wqQqmD0PibpAeetUP0w4TVdpk1WarP9f47fxrVEEbTLepFJUQKdMNrVwCyBIFFVp
+PBRneoPix+PlIVlgAdubSqAfWu2oR7eB3k+uDe+P4xNoaoACZhzCozlcZk4QaD+
OEwyLSFdHAfJbAVH3PRy+kg3NsqH2j5G+9RlHIvhmqtyesryZ6Sr9mdFj/iDSBIK
0l/wZldpE3XmHMuhXQTLxcwML5xsGKwvIEFES5o0QEvfQ/nzxKCcJ5U1PzO6H3M6
W/slPEGPH39rWy9uI/sRfZ134N6q/Y39l7aZlq0Ddt3m102Vx4nWNMRqaylQGVfw
LiB0JCEnp5TDYLj0+DJBXhZrTCYeqw6vg7R56j3Yok2LcrODtxi9Ej4/MaG4es+P
TUfCnhtcf7kUNTcsif/6ADBVdYopmDiFJZmJfaC40FHQRZaBofXTemWkpmdUogrJ
tRIajGgjkNaPR9qAAjhcLa2HZ1aQ0RHtBn/YPfKomerz7ac232odC+w8luiEgp0T
GlNZ0xJcsZmmHTeJWVEEcn2OLay74CdDMdcE8Pg7LnPNsitT4HgvEg5gPif4QcWA
zlcfsUUW0zGVXtDR6/3NcQYvW/fgEFqK+dxtShKIytYv8dgEbir87YWeLWjPz5Gn
vC0lhfcu9VcIark1Jl7sIyX3v2jbNPIsM0vgGuHvq3CrsQDDeTdZxoS2wJXEffHA
oAAaAvPyyUs4wSHFmXbHdVeh9lsXnhOoe6Epl2IWjKOkYeOs/iPEreXWcDTkt1Na
TN/IqttpBUjw14puUmktVpcJC41dPU4iC/ZwiufekDIpZpWE922kqkr/0OqCasnZ
zhQijs0HFzkrRGDltc4uKB3cNIyw8thx/RwL8YT2JbRSR+eMb0XkaC1WzCcDJv6c
6cB1Yom+ulRw6NZVx8Tq4fvlsO9kOWkrtLn1r06HLZ+tgkyPbei/ogCRY+Z7mNeH
sJiMirayK1h7Xep9DTqBpfDZ4E5w+xn8ZdmYVP3TMtR6gGz1+BkEsDCfXoUvUWRd
AV5wGkSZx7aUBiCiQurJevMkMSnSfFICydYB1oJ876ym7+3b/9w04B6yQLuEgGEf
ZBJv55eqxq28FTfAlfWaKr3Af8q9533CfmeKlMm2L/JlxLKD12iQYGQWcGxZOGFk
CzrMAxbBEhOX7vznF4sq4asecycXzEbZGdFnjeAjoM/TsRPwDoqk5e1fX5pBItPQ
v6T0R3oL+toqSJaHFMwitP6TMXT7hE60Ha87dUGzKrLltxjcCIq5z4WNJKlnYHNW
rE80UtYlpTTjpEFW8tXDXbDWK5DhJJQvwJy3GIY/vxnChm7tfVBCUG3OwJ3TtkP/
eSdgr0Nwu7mdj7z65ZZg+eRhS+F5J0rY26ICDQG/84XZJmAZZ6O2BmVVBOS39CvO
ezJHvxCuSXl8BSRFDVyPujfRVrHNpTKzsgj8tr1vIybghMO2uWow7OkNnhIJz4M/
J3X/xWRiAnHrsBAdigbVUcCslbWG6TIszD5mveR0EdrldK7WXNkfjhvKENsXF1Fe
9FVe6x4lII8zC3PetCBxpDMbGV1Cmo7IW84t3hM8JXxt9E4P0wkGxne8BzWZauCi
dukbukc+NiPGFJftWE29ToFMsFz5vZowsKDxMt10M4oau2YmUL8+jVRZJpIsrSbM
ruoBZUXLdkFKXC4J2RE9izXRnUTG7+ofqMfHyqBhVJopjr680yqNbsQN09Wh3A3Z
TtlsmE3ZksjasCJYw/X482ysxzHSWgNbscOWbkYp6C5GFTzOP1mOg7hRINpj2pOT
66SIEBWtS04rDW1Wadh7kJylbyzhYSyJ3QIf3LjZQzEV65nUVlr0UJY5Qk0oTfbg
P1ukwIgmghQHZ0seT8emtQvNOw3aTWFZMAMeiHuVvQkIjBiXw9bJYSuKbGaSfZwD
cAN2ovWBh3l+HKTjueEkdDUx1uPG6vKK4ZnPcFzTaEVwecRPr25n/D16ASX6tpxk
n3SzM05aLzU7NMSoTpBZCFw2tBJpSBsTiSlPCRUUt1sXbU6d7lLuqrJt7sbLsPaL
Yhohyc8tUcpsJIm+gJO3GX7g73/h4w+xa63BTH4+IyV1fHS8SwNAaJWsvdFoSb9U
rCf4lsqPFbgDCOb4YuIYtUT/57dmWR4MN6Rul9aM1NzmzTmqciEIjeeKYkJ6ZVo0
1cn0JBJKp3q1gAqgJChFRvCI5R7fcF/A12RAWJp0gkn2G9z4h85JQPlTvwQJqWvT
vTv2jk4w/Lih8aEh7fJvIR6nK4iFvhNszwuojjrgFBLKl+q+AKGfPGIhL0nTyCsE
5TWSkVYHzv/DMdCDVW0CWrMpedXppcjbs7kNd0aUNd8OsK0G1HTAW10m7qm7xRn7
AkyJ3614z4R5IaqS09pUQ1P92CHXwxXE0rO/5oavxOmIEtiVxqLt1X9N3igj0qou
MBUqWBAOWPdDMJB9Jex7m8ouGDtMy2A0E1l7Z1RjiVr10E64+amVlvX+rt/ThQ2v
o/a3K1uhyRHXGg/bFjpNiM/ysJXzG4bTyK+z5Qur9NqVZ7+hpRxsxEDwB9TlVn5a
P9hOs57RJ3waStkTetR4dyd/egH2dR9LbOGTYzqQaJ+23IoYz/pOku6/cUm3VL2j
7m5IUlvglXQ55RBk7My4vHCAhvdgxly0K1QarqMRfM6WTNqKQKIrEyxx7DUxH0VO
9WhWMc9c0XQuTmT5J8ExQ4GlM28gv7Ungx3hJ5eL3zLK7rq9+XD+EoNVMHCfhvTR
CRmchOYipXSdzZnJvRz6/3a89N8cvj3HerHzWmmsPer9dyfbgFM2Q07yJsTUicGb
CglC0hsK2FfcZIQOtKJ2MTPNa/unz2iOGneBsMVjJ0dS/WEmAKF7GDom00pCR040
DSn6ZTe/D7GrmxJwPhcnv8KjJG97wcEj27ziz/5lXYJZFjrFn6TbSWnPtENd32tN
E13/57sCdShEKIia3VxPw1fb+l6gybte9huKIiaI15+hxO35+CungAiJQahMJp8H
VZsWiB3kjwUq9nhRkaay2beTnEothcJqCFjAAp9+XpkBA6eVt4IMMhO6QRECXh0e
JQCeoATBTfo9fbsrQOgOOYd0lKoxU3hNt16b4IU5Kn6qQX2ddJrAmfogv4KOkwPc
wCI5RhxQEGSy9Ift5VG0H2OiktYS24iB0zUxIhew2X1bPotpN1CZ4Lgp/A60fTpv
WQKFB3D77Y8iS9HtpZuT3dFJsbR4ff4VFz8UvNrfnIHxT4/SVNsu2rkqMkw+MOHO
AysqGBYWh5mVR/bh5bGe3PQ4r8doiRmKMe7EDBef+OZDo1UUUfojWkJ0lUYPHU5E
Qzn4Z/eJpozFbtBlhUFYXN4fTevWjQwX5FE1RnMiuDes0CUkSo624bNEaFlEslxp
/8+9dgoayCrf3wlvKlreUbBVOjeCJkirX+QQYGTlatWuXtHc9UIfj4DUy/DnO0jc
NUxbYs5Ootsq5Xrm6AbhTr3Lic7TwuRGDU4Y3PPIKq1nbebHJTbpnegJj8M0BmJa
ayHLEySAVUqp/302nfvZeiYCCHle4tQq373SQo5CX4qv5KtCSQMRaSJpNXNppmbi
//12Fev4+1iKT2jNL684DGMty0spdCaDO0iZeuSWEh2RLzoCWEmHSbRn6vyWPkfm
yqbQoQ9DhA+TN13rYva2S+w1O3gEK4/mY4geYs8P5hUwdN+WNg+6rqPVfuWeYOv8
1bH8UUxM5gY5tYSZZcNnwFt4VQ4IGQCIHYOLuaj6suhaSPSfdXG2AbykViV6h+7h
zJLpbjjUDwzZUkkDe8AzQpH79Ai3ozJgvsCapag2UCw6pVuTQF7hk3S91fiWFwtg
49yIgK3RpfhvCKOnaiK+hBgq8scLZei9jfMPphEg/s5CrzRyYKAu2Tg4c/y9hpcB
rfATnaNnD6rEBUyHlCpB3clbEHeHdG1LarUmBkoL357TF8Z3Py8ug46L/jWSl8i8
s9uD33PFkUlz/ywZ3QQLZXw/2rEzkMHOUgoCueQWNGSj4kMgA6jn8nzxFtEsNdQL
QRnqCVBCwP0lFtAGzzq81RKfA++b2VgF7psrC5RGiqvBZBAuKyr8afuRTxwyHm9y
mvm74y2T5Bq0A1be6oexJ6RqXYHn9mjVSrZlOLgZNe+ZRCvp9iejrMVNS9iTryww
CPoCAnkzceBPvtrSKkqFYVSA9s3eAPX7vLP/ir1xeZ/mfYMvXJoKfDzStlR86oGs
Jd24wW+vB2UCHRlRjNrDCsxFvK+/DzO86LYT5H22xhspizsuEnJGM9GZqQFw4Lfh
VLB+8bEKayYXqn6PnY13pXe7+uu7W/Vpvh9Tw4LXMsVjxqwi17Z0IVK/qzW27wdh
Xkkji0dn0gK6MyYf1Py9K4cdD+CwEf112gcSL7FIQKlT2mLb57IaLl8Cv084JqfB
Ft6IfQSxz9su1rM6Ciy9T6DNxe7nd1VfHyhL95qvpkww+/iqmKdcA2p1P3hjVgqh
EJbyrEMzUbcDxDL1a+q46l/3XKHO9rYuEjPqk1fpk3X298ocbrsioBQlUIA9//+J
d/4/JTBFIbuYZ7dXvqbmeFLkjcS1xrceSHAc19mtHbtsaKfEXtXcvVpOabULclzX
GEMeG2WYfqcf9na5r+HlcW6+aUf6D+ErdIoOWpL93O46OKRCbUsxZGNhV9tlfz8u
n1WwIFZq+chcAS62S7Yx23zeVt7wTj1STn0GtWLN8LHaYwn1gtEN0m5LhEHGvno9
JAX2lbb8y68OUhkLgXPKJFGZQEr/AueGX0XzmqM/WjYzjfkXqhu/xu/MgoVNbr/0
BmijjTKFS1vSja+dqDxhuq5xzt6buXJgDuJsgOe7T7FFRVIf5duGu1nfGily6pUA
+xU+fv/0s6kmjUxYqUfDRcqrtuGMRFoExXmajo6TRCCoaSvXW3Q042t7mDosG1nN
TWMlK1J4auXQxfI2vGflukjAWcMiIXUdYwPOQoZZAQsuyFxa21im5Vwg9beOqTyc
amdlgYZvtbOZrqyT+b9OxGoZJ95lsUJKZH7GgRL4e9mhd9RLVpXka23YMOXjUmzd
XYxtbosJLyjQxBfKugN9qRFSvM0n9IlnYpcGJ5CECxdYgQXJOoT2cf6GCaS6t/nb
g6Ctm8n3Qau6gF2K2tRymx4GhVpX2Ljq2/H6h1zgUZ3h6sr/hc8aNs3wiR3Wx9tG
+yA+53ZsPvuUFPibdMej6TcxG8nDrPk3znceCjqIEzoGbKUJhDH9fg0dk9ttf7ed
W69HHS572kP7l0WyqbvofO5xqVpnYC7knoTEMjzrdkw//obqIGbQr/7jav6iLpUh
FhEzMkPopNK7gwmn1yS8IaQ+SQwl0LvG4WjKqnNplWoBPXMgW1CWdYKFfABB/l2/
VxoFyA7gxc0yAiDntVyGogn10rcQD6fR0TGVWEgPeZQhow+sapByJSfcTT7sVCL9
Lm6/6tWdya4Z/rae7GjjISz92EBj42d1fjDllvhKYx5k+fii+9SwbqwcUefsbSHq
rbRcd+d4XEaHvmDt+v90tCO+mXEq+6JqKn3ibVdD+khZYrKfERtajkbCVa9r2vCE
64n6SbF2lZwa5HJ6zaIEEbosl7kTGCCea7UnudY/R58I1ff58oufE95JEyYZEP58
83Uqg3sdqufjpa1bfOw+tg1+j+P8UoyLCwQoEnrSmysWkSRLnYNAq3pVn4sDe4MV
z7bAQ+LZK4rAYlmsQZax6s2NqIwV2L3bHm8nEmFirys3UDI0BBuJR7g/4MqF1cel
rcGVQzTlhzUN/XthXPM6sgxQ05iG208zDw7p5Ft27p0sZV++kAFvENxIqQleUbvu
Vjg/jSFOobUDUgjaZsldW2wVy9cjpANyg7knor++9KKywnG1GYGqb7WO5DceKrWx
qv8c+TyqwSaCPyaz56Av/r9exep3AvQduwCmwPhExFUYbjViNG7GOYJd1yiEDqTY
fZLoao3gqB3w/C4NJh2dZBMXjF3MoUYPRERiSAcRteQUIKuqFeAFtHyBQ3bI7Sug
j8S/QnuLp0IyOKwB5lREkmCPU5r2Iykm3SBGf+nRJZxDAHH2UL8gFClJC3oQSQUz
HGncnJKzsCuBEILshgAludnVTBG0pfUWYoe03GtH1VQ3kZEq53RvhVEW121ekc4Z
jUOlKGWRjo0rY1YNdpJiPnCNcz38oDYIqYIn6tS0I2SSmY697BIsRjTT61ajxdbQ
sdaJxzs4DvZCykNUI3AcchJzy8pfnCh4weR4Mzv/G1V8STr1xSlTVe7a7JoE/K6q
gdT19kPvkhiq8oEqIjYRw23DGqadxLKJ0iBRjxYssXosozPyAoA8mWEkPFgOEXuL
UAo9olavDTl3qMz0BvpIUSjm8/5BwnGLLpYuYpL5VNzwGFMmoVHpH3OV8n/TgQPT
e9aGR2tS8TBIfk/UEMibpxzV/88M0+Rc88rGlBqF2Njl5bQdCug6ArYvtQF6yFy6
E07gQk6ZbTBjVfUtDcB5QRvdKFExylm0Veg43J2udeCrJjjQBRxyBYZtL4hc/6EK
Y6ByTIIPWlRByzRKgn7X3Xmao9q7DkbzN6wi6IyMq5dcgAQ0kybArQ0L9fy8RZBF
VIKgH69qrsgs1wu7LpNjQ6EHM1vSuxegk/H2NBTjjQWDH8EowDuH3Bp9P6jrlRH8
63Ryw7e1KyJGr863PXS2iLoXfjMB9vm0Vo4rqPl5NVhI6brHa0s4DSf8GapOWGHd
tntxi1QQmoDjP97/bh795QP5XGfw9GXGdJF5oY4zXgW6i7CzOHwEpkMijNCL7Vc7
Ysui5+TTL5IBzBY4AX8TPyKkcz68LMSoyetSeVe1jGzUUCtmN4rUwsytHII1QADZ
Jq+8RjE7EkvlAzP3W2+R4hbm91/BYnSjGWjOh9xf6YvWk4+OlE3Or7ga6nl23Csu
dry+emoJwN1JL9STcLEZKc77yyM+FTmwM6W6AeuY+x8lU4CNe41+UvuJroTxjze4
Fp5mJOP9Zuk9nqaR8wsEEosV1fOKzCv0pQpDlRz1DoM7Ikep2xlFRxVvLNin04Ab
fCgDjBCGB5OznqhwhoJerN+2eLiBTM4IIFkWYUH4ndNcQLQgcfdVYhER+2AYdgc4
BKLbx3+HaOD6uH2npeAASeSRoscslB+Pg0hQVuRqofP4ZHY31kPGifsnQEVLs6va
WEMHzhEJEB+cT2pAsNND1tcLbcfeJFFnEZQgnHfWtzVg5BoXGTEZPAroneemWMZr
Yg7rnpTEiArusCVSAncDWICTOLY6Vd6xA06a9aN41dIr/e59MROwX6FNwx8HosD2
Tn2LRqz8/jU9Lf2Nlh5BpeqZTBPeY+Czou3KpKQhGPE9a/zFNJOA4a8hh7fGKqDI
OBXWywoNOQ3uga3tTT4pPPlmQTQVp+TObvOGhxxP13OuYWo7Vql8FoN9qM/C+/FF
ZRmkVLoCSHKztnxpbk9y0uQ4WSK6q/X5OSsF/fWKkVMeC/olkYwa+Fb3lDcXvWJB
tdIl9gIsnT1gtXxOKomUEpw72BGZ/k4qTviKXAh1vuOwC7kq9L03VFBxcYRQgpJv
aRk8yEEqRQTYJXTmj04yaF0pAV/BxDF+0K+fM63y1Ebpoq8w/QVCGArEW4cnmxdf
WuPiPVMRC0tdFdlDNd20H5fFJqYsusuFkkWG2twV4TKoU8zW30Z3X6581VcTXnzp
w6Fs1NuKJGslI8o9zsTKQsTXXqOCubBKZW/1OmQqqKxQOmzi8C8PjWD6WAHTH3bU
zaHQ3CLU7xCvlCK08SkMwYzuPISwlKzLm9KyiRsLsKaEUL9fOSJEGPcWMEeSmHti
9AYhBnqe8j/m1ad0m1xbHbbiT0T2rkDfPrrovG3eInHyj66cZtNqqw/eqLfLhCi7
mcZ9YoskbhWxg8aUtaQaJC7piUDfpihccahrG7shsPkQCs7H8w17rWL6oM3W6KSu
ljH6axJ3Vvktg9sZZr6PJMY9YNOXAe69EzVCQaXt7DbmoOZCNe/FdYlYL230OA9v
7PVVXTkd/9ClkiIa5fbP4ypy1PIt4Vj3eKKSLXquSuEnBgCcbJyBlI5djZC2LTtk
9md6yo9X33eC8R8C1WNT2teriNcgFD66MhihkEceiaOdQd35X4JeN3fH2eCdiWYa
pF3F4oa7GvsS12bL7IJpFYKIkHyF8dgSuKZC7mA7CgFBoFjzVQnTnjmm8zKTmIrG
/m7wUDKjlaPefwcHH0wCT10D/jI8OhIvn8FPPOntyXsC62Me3T2LQeRQL9GzrRZe
8SSOOxs1fVj7nhU8qfsQH+aDgyYIKBmvdpBIr+y9uv8YOVEBfMKcqiQeUus3hA2K
R1Zxvt2+fQR3CVElICtykGBoPQ+UHx/rZLFfyfF4r/RcXtDWNa07olbG7SrRh+D5
Oz6uvsCCf3/yN1ckZ1J9UngagbztgHdeOgz4g3nayH2gv3/3Q5SIosPTelqofbXA
lcjdH0LVy+bF77rbq9X2QFwaUlAPUI0IzzLi/Vucz2veJEIhzmlLoAxazlgavOGz
kGUGBOsSYKKmXQrLN5kgYDEbuuYC7pLnf5SFDuFkgHrU7Z+8/G5i8NxudW5CpQWo
mgD5jRHGSlByvP8JnUwv2ONv9xwWb7J9saTAeUluri33i+KVY1n32+Q/lIbGcaCI
LPcFiIgLWY3tjVXz7acXfrWc8QNMKvCoy7hvbGegg+VrA8DdsI24z3h1udwf0dMe
5MYmSd6mU/o03dK79el4WPKxKuHBp95qYVHVtvH16Q/ba3Oe0zaVvcFsSRAIuY47
y+cQZ1D+d8Dvu45pW6LLQpby7oDHggci6BpQf2SE0nGhEbqpBk2sX+0u4clF1Xie
k6JiybjQmn8/uinrKontR7n6H3Ihav1qLDoh/EzgZeQSaWzUox0I9A4y6lyGacN7
CHAIxe0I29oSA8Ov1Ha+ySKgRQVeoIQZECoW0po6vayqmHJdBC4jODgZ7xeulHDL
gpWiDG5c6HVQpc4mpdLqJ/zpMzdTiSc5Gljaz8+3fb2LYizFbYq95HXP2exkLUuv
M3sOZv7HJnxcFg9yxH4eA5eSMHVc367u4TFDDZyJJZ2nK5kUaj75VsVGF8pGzD5h
voK5XNql8L+hq2EBTduyxdLxfodl4NHJYNOsTrGKnuSp5uC8WlxASina9Sv9wwre
CQkHGeavcJW8DTWimNue6tuGdhRd9ixtdZj/C1VmvMFkZJqSLYwjoqv/c/VcAOKX
l0NBq/0U7yOg0MQnmyt1emhtEVGVL5mPDPeN5sjnW629P26PrCuzrs5tLLO/uQCp
GoCtccYqGX7Kg13xc3/8sg0ZTiJn/hlrehNGbFOw8YM0/Mk3Jh9yHm/tXh2VcRpI
Z8La/IYSnQp3qzWNiyWdI7ZKRKz7vPOSts1sGYe4QDb2Bc/otnvQRf9G94SLB8NR
vdalTqskElN9IBDXYeoYlhjY6FQAvwZGSZdUD5gNyfk2/3czE6YnDBAkamsCpVUx
pvhx1CyTfXhOhljF/f+FxrH1yPoPzzKQVFxRIdfiBnOJr+mZcn65msKcDIjgWLOo
hHAFk/r6QUVINB6f0eTiYmG33MsPEb93Vi7nZOx/olQszFvrPVYxG050CTzD8tpw
/USYcAgDOkl0AbaHoXk66WeHPrVmsDaUSSZlQsaQa5zSaSuLpApMZHOKws7gOfBp
jV4HTFGqd+FlMYPvN4Ol/nSjhGefl231fjM1jxSAlbS/6Ji8a7bJb58nzscElwAk
qLWmuvdTOsZ4MbGMfNBzqCuisy43fq6CjrQY/19ZgxSiQNZs7tyKhlUEboNqI3Zh
1VzAhxEtLG5/0B3LRa2bTbNj+mIkroMrfEPprvSstbxb3qZaPmoQP3o+lEBw/+2G
9aKUVwldQp9cq461nUrUSycPq+qoNHkK6qnRwBJAl/37IJjuhejE3NFy1SiBkrI/
v3abuab3C5uL5kvH8F8blUOsf8QiuDIuV9HGRgOrIZNLtQB5eBZt3kHNKqbkQWpW
YiVaubfoXcFEq0rpwqlyE38cJ2rmUBflARhsLezSmzweFPtPw4tRQ+ViCZ76QeYi
bST0Bje5uBdxWsGiuwKO+IPe2HNkZYXydvkFP9XweAheMXVUfCKsaHCXU4MR99Ju
iPPqQBqOp2+l9fRHL4r7Ir5tuj5k95GkqM/w8KWCZB8l0nCYHEKso7BMI6/MpubV
SMji77xPjvMieHcFmpkMy20v+cVemBu5eGNFTU3pKMZToNVyf0Wyksuh8HxvfjXh
Au8HOBPdYoWVFqDMrlKHJ/pGXlX7MJAES4PeDvjJKaetaoY7sSXoWRTi63pwqaq1
HBPxokz4m96EbMazVNo0l5o6439XKXwYzHzy3yhshjvW/j3VwVmT2loMXw8SnX6Q
YXGfSxd2lUg8OujO6pnlsMxuGycm22P/d+XC4azp8KdHQURXBaFnfOxuokWXESxB
DrLIdFUXfNABdnPr4neQV2639sjsb3xd2AVxWXh89TbrmH2kVU2ynr0Hp99cFZFO
LpzDY3ppS51hDzK1lIaAP9O9VY4gS2wnwRw7mGexAg/YWtOF2LoWRTdQ2yeuv7Y6
r+M1m1Z/Uo4gJYicQY7h4T44oxT9Jg0F6ZokbDigQhC/1gMOhxnF6cBGpjRKXJWi
MylYxkIgIx0aCkPt7Y58dGNHbxBxJPi6mMNmALOUTIVDjtUToIwFFu94YVVejcpl
tuKXjGCf6jjapvLa63/cKdKxh00euxkQut8y/nlZrHDkHD5m3OYM8thMUR/NFqYz
JJdZVs/SOY3cbi6TGFsE8MWCAXxs5bZinlZUaurqPO5IUOkvQseFCDwglgSqXlFw
Nva1UwaSqzrEWkmgv/lUN+q9INYtuBeC/nZ4SkoGJRdL82fHHJvfD2M92F25/VGQ
Pj6X0c7ua++BbGf2ZQEvToB4dWYcb17dDTRw88tCEKfZuslJWj548wrErwWmX+ZV
L/9qcUNOFZlzip5TLQbAGv3KJGj/OhqZjdO3WJccDrriaYCWfF4p2loM3T/Aq6vT
2/0SKY++ADnv2XyKIMmlXuEVHN+LJh/+/XNYon0IpM+X676PH48xBiv/CZK9dSvx
8urbjam3QePXPqYG58xoRIYvRxsLgpTOum13ESwvHWDBfPZc7kN8yjSVjc1kK64a
fHOmiROtNJqYShHfUNPLBuFZYH85lB+Fa8puN5VYPwseAdPDMDswbX4TJVIh8ePx
AwXDwW56mgCiuiwuD3RIpR3po6XryKgdUDQyunwPvaPAF25ea1ApRjxQI48RI3fs
EWI/IUL2PaEfFB1BoILs9xggi3aQTcZs6ANjBFq3I9SpxZdgd5Uc/d5GcYV/PiMu
3LSNC8QG+2p5YRuvUP2YbrU3pM+CNnxgpyY6bXWjEXPXEV7EaALony/POmNYI4wt
GBkpNCQAVJHC8Sj6apPCHdlDtFu5glmbieLDKpskJaThHnJk20wqWwFO9zbwGQ5o
U1Y78liTpSmLQb2mQcXKIVkskwqSiBCyUjR2y5U20F0sVa8VP8IUDSBR3HSWrO5W
DUGKQjagIMPa6nZCVmZr/4KGHVPGYttGnAgRGGQdg9iUSPgWxZJ/86VofSA26otJ
5uU0/4J2aCNpP/EwGxjyV4OxdROo4BqEu1ny3n3KLo8BqLczAT9zvgpRWaETuR9L
2bcj2Jlp3V6cWj0vVgNXZ5/RmpTCi/DLQTY1rr18kM163j/gdXOvGuqcHRfMB/Xr
Uuj/gyZnSekzmsB/xkXI4pVgSSP1u7cWpNTz7JUnI9tu7kMcgnWPj71pyJb91ZeS
0AeC90/EpSq+D2cFcTmElAEgEmEmfiRKvfAtvUNEg9vUxCp9Zvp3drBKSEQiJ04r
96w9OAb3Ckm6cPPknfHM9gTj8INl5WtZ35Vp+M84G1xkYg3TVDwTS+jxZTXEUSRa
tJ8+68UmDJkOdZ9GN3p7Ilrw7LikiKvvG9w/uKPr/KZ0ztasO8R7Gje9RyeAkz0b
QNdozziVcQZgB2fpzXeX6xQ/smyFt9YsmEQ3U1yFbCJFMYPyF8JRnUVLZ/1+5X+Y
UNjUX/5xWHajwx2OdhcFXQJ0dSXEkUFSSX6OFJIQDB0xbCTlB2DewkegqagpZukQ
zC1dri2sfOSVZLdL+heTEIGwMdqT6JPaB66Hvsh/LbzfjpcBfdM+/eYITMgE9tQ6
/iskFhyUfPlK1hxJ87WQIQCvTvz7LtzkPEQLlvAxFPDoj7f94LRd32o23lmGCRc0
wMG2i8fScjLEw6VU3YgS+VJBm8mWMSIsOJ9tZz22rDWcqULjLO5gvWWv5ibb2lLy
LTen6mKoYSmzzwE8Kdg36G1GTGcJhsRJRMdox0AiHMbg0SdQRUG8vfTqcwmLDq1p
aQUrN+ISG7V7D6noMRmHtNtuDM4C4TyFMdpVLPi+kaWo15DTYUQ27Giqn+XIsLwd
y8m+I4Kjvqdg53RC1wL7hqqIf9u+lR1/ijVkyyHaKdsUMiHd5r6InQx76d3jkzQ5
NFaY2Xfv+qxD3Ar5sLOflpkrZO0tkvc+hTepVOSy8X+WV+1Pzkt7IfLCj5U0z9g9
vVeQ3vyb4IppF/503Tusf3APPpWkwumP0aENUsKMl4sSQMB9WAKyMp15TyC7ryJE
JaPqew/qH8y5uaXUQlAorC8oVOH2awFQJ2BxZnwMfvinqki0e5hBxaFGfBkfZcO3
3Kkh8kyhnz+NG3QdMgQQ0RXXeQa54LlP/Eygk0b59dU70ALA9e17ywMc92UK3PR1
Papy7kfEFmTxZUSLNB6qvdv/6lMA9VP0PzJtofiWRYC3hOk8vu84Ue90B962UHk6
deO7tB+qBU3N15H+VA02B9hmUyum7tPKSTFSia2ZzZWUua2P7w16f7jYXvk+3gBs
prWLetNBeIumiqUTkPZ8p2ILXy7T3NAgq9hECDjKYuwj223+ejjvpZ7j6PMmXtdS
cDeYUQ4nSQsCsB/JFvU/w2JIwjY1ymOMFAd+bdFrkIHGUrcY1nZex+dX8rT9w225
c22eFO/iS9Da2v/atAABWZYdWZIeOU3pAfsqR1ys+LWAS+mrwVw/KqpwCV8RTgWD
0R6ZsMftbDbtorJeVt42rh4GH6QPLmRcRo7CL7FyiVAlrd4dRZRXCSS/kJRbjstq
/xAhOWisYAEBQVuZnLAIoV/iK0Dw1KvV+4Mlqb6teIUhPtnzvitIFQS7exUVbcEF
7hLwLpS3xRdvIWsZR7sqPBbLKMQ3HdFvzOzcR3zxMcE2VokHXMR/iiSbZQKQ/Afe
C3pUQ8+vt3Upc1GU6UreXFnvu5ngvYv8LVruY98sCQRp0YXwGVRObUEgSsIwT875
fgbNM5W6Bq6oIfhhIfarvwtdLn8Oky0Y3LxlJ+KhTRKC8fc56s9TCT28BuiLAux6
mWuBC9RuFYPQnwfGznLrYANItouMRMt0M8+VeRklBZZVnZ7uk3Xl2dmHczFmyC9r
X9zFJ78dE9X0baK3TGeEHLTiYYTxjQ4grZD4o6wJlHuLmaHcBfDfnW1xtep+29/4
bNOH+xkXE/DAg1XbJt2d7WDnpwPKWmmQCUgETVi6dqcC5GIem8VIYPHwi4T5Ykpd
zoYiyHp1QT46v1oj1vsyp0RzW30KmTkCwrS2Uh0xPZ9vBjPIs5BjhdXaHMDOgbMa
l8tp/j0mEFWFnnXVpYfHj1CfCrGkjy9eR0JV2vKFbS6MntOe3bhIEmbjj0HagFs9
wiUNPLbHpa7FMRnSOOED0ZwpUIO6G/O4v5ui7iJw+vAauHj/bOP99NqOZhw07uXq
3o6nmntDM4JjdSqQVud/1g/shTEcd4MzN1tAkkmIWBEnKobTdIuap9w6iDoNObYa
/l+hbf6LKa94BU905/KaDqnHTpFsxNpMuqNny0SM9xo2qfbsYXpqnohNf/gopkom
PRFDBJ5q5PAx8ZtxeqBkoaO8fok7aUunbxrTC9fRinjD8qiTJli+A/XPt0ZDJpXi
+pkHABcp8JlP8XfRptZjl8yNieMmHh+Ahj/nPqJZ86pOEvH+3eUO15ELSTZ8Jekc
YkFhOCWuBvNCnCsIBM+9EXz2V9ATKxaFsb0DojFdfjKa31WSmARj1f0XZJ/Q8Ibd
E4+i4k9+eGokoUzj+EV5VNb/PpQziYHoNX22nJqlfGD5X9zyjb/I0IZBktNo5MR+
tsG+ZWp3tmYwM6L76bvI4vQUnZyCAmIAF8deZosJTA2Ib8X/wsMYRmJFInjr9eRW
PmEfN4VO+qpNj+llWbGYygg1cyFWMvqVvzcFK7p00cErSfVoOAE4U/btRVtZDYU9
w5d+QqNSAj2kLVFb100fSDGqmcu4+fnesgyZc0XOjMCS3DGf4q+jrfV5gDtjUfHI
gV4FZrUbQ9tpPH5y3hu2vxCVM3nNlK4vfWf6yqy178gRcts2DQ4xrnhuN4DFlpve
ljeFOO8cZqfc0qZFIhzb/iXlGPgEujhyNwOgNkLFn0V7LDYK2em9KUZxkaSGyxYx
gEIOFu4tpZbqsPXHwMboMRpYreit4hHUqnAnhYkihbccng5Zbqrm3mGZoNzy6byQ
Jb/xMoaXfwJcsRYnwKtmJlf7nY2VxmJrKtIK2H27Zygq6u3DFwXeLtqCrFOFhQXE
/GGCNYU70d9vVDvX5eHs4JCGFR9MO6WtEKuT66q/vluxhUQYxdNf1RfnuX2QyA/P
kis4N5LdNXPMc38yn9QYHG+trebLaegP6pUNSMNoUZTbXHmZmipn0xsLiT1L1EEf
VAKQr9oQhPKKwl2dDX4gDABFB90VWo5DvGm2J+CtnwxXx1000yYSDNBWMH6hY2w8
70ZA7qdKgoQieVadkQkfVVQUhUm/AKN/gY/g3o65k/36JWXftVgd54Dt/u792mv6
oH0OqxjZpAQjKNY79sabH0bJMBa+KiKSIWDw7clHnV94I5R8ODl8mgI86HkvrSHZ
3aDrADhvwiS8flW7QvS46UvJ+CXdASMd5y9BvuzHczkaA4NI6X6I2QQHSQJorOFF
+afWOJiPWP5YwxlwkwKtrOSbhaBSqtNgSXLHX8q2mpPgeiyWlTN422JAMW2aFuMR
orQ7789LP18i4RA8TmtHAPvWLhi9ARFucn4stjBVgjek25LxOMZrJ/iC/Pyv1fv1
QyLpK+f3EkqAMi2Gs7S09AWB4QOxI5FH58ejge7Agj7FHQJgMG8uCA072+k1bBvY
XHZUl26gF8t7JJLQGzVVrPrvJtdBfh4V09+mwV447FUqVXJN4n2NStzy1+wbeDDR
8nmjFDUDCYiEDfwbmmL5UdbjelHk11ZpQd01uDwMURZ+4I9D0mxvNgrtcAE6EAUX
NZBKt59KevOSBx+5ABq27h+qJOeqTFYp9bYhjDwTQPJKmM2ZatoiBwkouVZ/q2LO
xj4p607qck33MSySCc0UWzqGV4EdgRNYT6uVzn8MgQ7kdSea1oIQlxGRV9GuffCO
t5dNNZIf9ij4SaCkpQ1iGuecsCdDfuO4KqBQukuzbKVzjtDVHUpfLh5gXSFVnBRX
9qsE7yCx81TBFk/PwHB41hmmXRLAO93L1o7bbuaY81iJbjn+OGC+sGtRbbUaYPpm
13ewenhdGY9Thm0RPW3pCJsk8hr2NO/aTgYAZF/dTlCAshpbWgnMClFJW7paDDGy
a41rTOsi+smr4tL1wsvQds+LIPFqi7yRkylPEg0QRSgzssxXivtpcEinrbDQj6Qn
EzUrzoy8STQFCkZDzHd5m7nqcfSDUasPoTeQk2fi2oJ1dogm0onuebSvXaLFdXyt
WcOxrGXrDeqjbDJ0VDZg6wbXi1cvl+BzkTWpu5gFqUjY6dq+cxM/eepy7eHu2FyJ
7g3l2zzLJ/JSIqqRgud65YIgfrgUiT/Gd3zdhTYTVEchmR9G8iRXiprwlDgnr+kU
tAUmKCOEIcqW6NBNDmcohvzUHiHsb5SLVZXFBVtQ0lzXCiYIxbBCwRytOircd/cm
w4nyJKsB/bjiJ1H6i+dquItjzD2BgLv2mSiw2GkaOxpZkuSCTk9x8Pw9uInBy8Bc
8Nd+nJmo+TYcKp4ZspMF67zia5RzPO7N1wgz42dI5AeG5tsIVd3wKRKrUQ5/5vbz
+xXxwxkeUJw4CBWUjhvtT0ehYnKER/peQJs49Mohgj2xP5QzG5iUZXBx/qgPpfoO
OjrHnYh60V0H/NOQzrmxIa+4cnwFIks6LNs/kfzz7c9zhjYoqenrqMWiy3eCfJ7O
MCxIBV7uB66QVNpe3ZWdQys6KXfRYtA6ecyawHtjtbf21fWGY5LFYAK+rDpj++qA
pgv2WbXNm1yTnLqlvPCdONcibztZlK3u/LhBTJ7Sh8qO3xjmAllB2o8GMTEOiLpo
x4lr8HO4mTk96qTCmcd4AhClS39493RhGGp3jfJkXPxZRO8VbLTJx76o+v3rBGUX
e1O9KZ7ylizOQbN6a4/F4rYMdK8Ga8pGhbWj6tJAdbLfiJUv1Oftz3rML0pLBOIV
F6mh8SUYIpu+8I4Oq93ObpCaDuEiNfBKWXNZpuTMcSFLmDsigNzMRMrv5MU3ba0h
qWXMsP30dNreiC1OZyjHSf3EaHEVzUjCnvDLPkpY6fMACD+zGUgD5YCywPblGljd
tUWYk8jdR6Cuk/JYN8S+L8i5OT4fAzoBoeDfbxccInwQ00Z2ZwcHgLVBvQ+3Uydu
XepHE7Mgm/94jP0cy9wNbF63ugMwvBcrQIG6vuLLNKF8SsH+6NvlKirDAW6D/7Ze
V/Cc5S3i/rG3QDAIN4eYkWOGQFie0Bgkylo8r7XVpegQ+UTwIZ2VQeDYFJXNPKen
81FK1bI8eTOFK/licG08IGC6EEBALs2Vi+TNjsgPigkLJAPtWU58kvma9+WMZpaq
JbOJLatwsGti50rBJs9Z+0PDcD4tTd6pYWCg9BQdzn5KMvuXAp95RAuMOP0Tzn6E
dG1d9RjPvZBbSUgn3+NsqvUxZVi6Nr9+HYQ7QtSiRNFP2ZSabs0QWasFMW9R+DSP
kEQMndDR1l1Qs1NwENxgB7Oz1LquuXWLDoxqGmLf28hGGij9W8rUjZaBq5ZTjYcY
uMNdJ0IEOVI6dwZwbuWa1KcGIBHwENxkozafyL7jdGepc199tx145KS9pZpw1Myz
VsrXYt4c3I7IS/l/qkyxFtffIa3myNrbF/m9q/bEG/ElOje2x/yTCRNCl4liZkK8
HSzFC3uDeMg8DI6UU2PmxJB/i1EBj61KFG/yxCFbA/dhEHGzGuqwZldZsNUoqhUS
pyB30XA3r9IL+NKUjMj5aFAvSfJYQiXV8BwXaEClTBd3ZYG7jm1Zw6YyLm02GBHw
SEk7NtAnUzhRjxw4Wozc/LUdEW4c2gcPAzXS4iZqsseM+enNUdFrN14qYvxcn0Ps
S/ZfoIUIRysGq1z8uEpHKRRO+nch7pm6XVsWY8/KciGCGp/5+VysT5JUdJxAZhyQ
xZsVGKqnJBLc4hlpGd8jm1pMIfLM+2Ko9HPkd5ofJZd2PgsFSuh0YOUytLBdmIJ+
yL7iXGQu2Q0Nud5rrBsnEnzdVpAz8fDFKIyXIWjM4Tu27H7Uykes+eRhzztHHVYj
XjmVQCpEwAQSrxO2Gtw7Pv6mACoyKemui1U2psfXzDDrituRTatZYibI5Ll7lON4
85QQePIxcMf8fAYgzk+W0aVmTj+S7LcISvDqhk2kJhv0pG72IGzWGsuxQ2RzXIoZ
XbL21JiQVmnsJXqjrR/mrKJm0ggdS/eimsq9j0hSMUJ/cTyTop8QVjRR+/qEoyoZ
8TmXLx69hMxw7qOLZv0hIn3Q5bfoBJFSjrqcURzbB9Jtnqx4/wQDZUz7mwYy9zb1
rmTetsHKk9RWDa6f0BAPAowL/Va/HRyMGrKYPdwO/hG4sx7sVebHF5Ut5X+f1cRy
0xQtlKguvh3rxWxWbgyy/SApC30AOblJHVjh5+bOtMetq7GKKLq0rQajQivciq1e
RA5TrVwUjyxXoFgbStv5A4zasTOEvUGuhyCYez5EWZ5wmTlXidl0PeDQXCLqwvIH
PYlT1LpNQ6UUTzq44tvk1/duZlnBkeLqe1q5uJvB1PfH4ge7t4xhpP4erOoMVb7V
rTtc7Kzy2l+pE+fuqeOOD8ekuRuH/vMLODwv2p10wm0j9UOtwsHGSnUcRShYnNR3
VorjkL5rg2aglRl4lvGD51WGPS/562UYGLDA+ofYCEg/Kp6bO5GSPQhjjYVxefs3
C7hwpCthZGV2AZPje9+NDQpkOU2NdX02u37+hKrEJJGvaRgDmegF4XAr0WY6849m
9dZVhkSUozFn8y3EBuuwdVb+Fu2uByG33k4S3xDCeg87bLzHossPxmvcTzne+fxY
Dod8GvGB67cFq71adok/j7AMi+s0h71Sy88Hebp0SJahHkc09fWy//KLNtovFBTO
eXgWJhkiwzYvZMRdu1W7v5L33y4GN/+1nM/QoGTRyfwUnSuGsnmjr4KGZ4AgPebM
w+EQ7DpwzwIvLw52nunjlTUBuaIeI+Qq2RGHtJLvAcCraDuDW3yJVufokwm7wLCw
rQ7ecXzq+aJ1u9fhQszch2JlKsre6wrORb1edc/BSf8x9XAsO5Gw+7ZqsgK4E5FA
mUQG0by/WPFdaLw9Ai3lep+YQ4+P1d4KNPC0aVvdlZKlZ86ReJzsQs0LUfiAsRLS
0bfILn9EyioBeYK4z8RP2Q1bTuaElRXRqmkOsEklclStfdILioAED4V12xvgEsVn
y0IUE2zh+ATKlR2IKwsLVXQ3Ac3biDOw9L6fxYHC9cGSJWXCSa4Po4zMlqI8V4fP
GfwaCqixn9Gds6SMdhLWVg1uKQP8P/ftzbXFzzZ9drvvAOxHcFp7L8HV20X0J5C6
8SGmSaHzGLeblkgNEIVb8hGTUvw3cWebXe+b6eHaRMcf9jcz2e81DWLviwgKimiD
m/1iDaHpkePWi3z+sp52N58DkF1/XzJ0Dr7J6WERkMghidaKXaO0w1G/fsk3Asns
rgMxcOuos7qEk0RtLoYEajQaJZzAoXc5xuHKgp5BhbsCmhT+Jhqp0QQ6ddZhhiAE
HCXw+ly2t6S0XOrvOz8XWRuneuGpeLBBCt+M6laXQw2KzU3mww2G58yuTuta7rMy
AkFY5d40QJM3Vle4QJo9ZyVwWz1UcSNIIDXYqbVPKw+WIiGBdQu5BGx4uShZloCL
SUUeeeyv/a4/47Cn/DJOwJw/3ADkSFJoOSkhwFSDVwKUcRsnp6Aa1MBWbJmi6B0U
9PTtDvd6aN3Ou9hwic/VgoIh/SuI7Ao7g09vO/Tf4U6QbuBqtqyEZn5lYamY45rv
9/gMFXdtzulEnzZWq+YgpcFqMV1du4/RuPej8tpEHpg/0yJbuTS6PZ+iTC0/jTrj
RF4VSkDhMjUGB2LOo6ZQj0gx7vMDw5/xDnMZ+oozxm2wjYE881PFCR4+iowxpWBG
WLRQzT9WI0dQKvCEZ1n+ZX8U+WezTo2bZlaJjePGnMO+yhso3jLLA+22qkNPJKaD
4TRiSfcjza2KuYPuaV0pL60j3fSubo/LW06Vgw16V77Gmk+fieFGauUuQr3E34lf
H1wZNvdJKVBQnNTukHO4yLHlkuQ/UqNsogebN0M7uojjPGcxUF2UT1k+yxW9EqU9
B/QK7MA0wI9cQ12DWXnCg2n89HHTP/hM2ut3LTV2+zMd4VgsZ6wkt69ExWIyveXP
3WNy/siJpcc2XuCzYg/BFyHAGwjrWdMahrSE85HnIsZpeKn1o9a8ZAuGjeXwXlva
kQIW3g2VL1Jdemlm7OKCHyL+Mlp57DCWgNn6aM6OJV1OIA4+TWkMIUV8YFxHx/Wv
IEYxKXF0Q4pdc0boEbkaIU5xi+o798532P1I5zFtqLCliyFAo4PDJjygiPUVsKzY
7XkWo+KNb6ImF695Vs9ADFjOyyLncLxKh7UFhFGIFC3KSt8zmqslsctOOkF17k00
faicrBrRnrQ4ui5o/iHmFJ/U+yAYvzylfijfUAFjJiaNASUF40V3S/pmihRTs84F
vI0eDOUS6k4V5oLTIGEzVsLmFEbB9wjikRgJIhmKs/MeW5SgR+C9wsXepBMBiyht
1Bia2jX9uNabE9kyQtPeTmPmHvBzEo6gPT+QdSBMfZYJG/2cACcytyKNs/NXKPkV
w1WrmHG7d7Fqzxd9J8bGGxlI0svj3cKMq3ClEGFiUEYZ74on/Wy+Dh+Ic5SYRJwe
fD2vYyBQhxY5kVqXVj369f+zsoAmrE6IwZnQC+ZKAlYYvzUNB9LdABO4c006j0lC
vMDzEwQ7jD6m7CYijpPYMFePge2NroVIEodT+VKfYfttD4NKwk00zowlm0PL2Pxx
rjmFtZSLW/2BT19N+eqyfNeDoDymZuARq8vpxrOvQH2a3caXSb2TlGFvwmqtyvSW
huHO7zrqUNqQ3g9USUigqG3Uf/mXj8hzP0mCMwSr+3VsQq3pOnmG/yNyGa8M7ivY
cGz9mb+Ggqx5ZOq1FrgF3D3jFpyN8DgOyuYQZO05uHggm+ypI72ozEkl2hjwc7u8
ZX/HQ9qGFWK60OlIVuaLTZzFJ4E75uev3F/FjOxbhbIc/Q2ptUYLXVLB58oqckKI
5S+3cXsrqSqCOWSFsx5Q1jAfmxkUvG359875Il71YI8E8KtbX9s0rEdd7YoDxlAk
AC6hldwFIbW5PHfhNHagtusey7BIVX8Cj3a9W7odpC0BOf6YzglO97HkHz+j48T1
OQWj5G0bVJCv7mZ6hIsHHBuPdfwTZM5T9quuy9kAQoUQ7mw72uU+eiFj3PpeaBuk
/00uawS3bfY0cydIcEDTZdL1Hd3UWydeA+P8NJhy6qBak7IliF0OHjgCgIpLSjMr
JpgdEOgDDtasJn8x00rCeHG8mRrxZ9BumggSnSPI52invi2ffOJ1pwJavd7TQarl
vSuSrEfUJlJPovw9mbjLyHwa9ZNOPUnEHjZelFeenyX8YROvFGJSmN5u/tHrYgXU
IojimMLmbS0fDIOSrff1U4iLfM31LLP5HrMbfVD94YoFIL2lKI526ot+HEcyoK2Z
VTxZDyf8YHi+W/IZ+zCvY1OXT73GYnULODE2j1Bp+633F8y8EOt+87h575LkVxk0
3C2LFms2ovb+9UMxz+0FXMR4ZYrq6d42GXF9y28VChdzNZ8ToTtIixeQDGL5ZruW
9uCdyMc0cJHhdyG0shFZgv1ymNgQriO2f6ExvTgsX6lagcZ7Oa+c0P7QV3XSDSjm
s9ZmOmm862GRgyLaVY9vATIg3rXMPJCbOkf2l9TAPIjl2MJrMZk1dyZNLVlBc2kk
xT/U8otxudCedHRDVm03XmRai6zFpYyIpxc7FT4722h8jRv/xDgdoX4ysEf1D/qb
PiL6NN6BfieiISP+3Pyu1funeA6shk/zz5/mI7hylwRtOOBMEXBAw7ALSjHUUwVD
2fMOE0rraTVr3o+wGXUGDooD8B+g+HFJrxMbv7zoCscyJd7UpWFkfZ5YDHqjzmLw
HcfYGRWt0C5jddO9F5J9H0NyPYaUng9N3RHXyC9b2co5uVhvuiBosp51hcfRhPAa
ALunpLvwXAVnOFj9neIANXC5jMw2mEeIK7FT33lF8TYPI/QDwnGya78997r9BVvA
9QgPHscEvItRbM6zfYSvBsGNs7n5W3PJziiqYd9sLWG7aZVlGfKqE15xbzYHoLka
tYZcDhmAKT6igeKrKQtNCU//3VH93lgpA2QQDMZWCJSnFe1K9zwhu/PPqfK++bN+
ioJXRd/D2LQD6raouZ2wW1KcPmjki4QCzEEbeNMKTcKBs6hO0Xjk/tbBFNCbRkSR
wAbgtm4Llw7EfTCUyfGm+PKUxkscqtZUpGrEefeFm/HEJuY06P9gRXH91lyyEvbu
rYNusNu+5pRI103KZ5CBQRMW+Sdn4WdhiHMVmkiqRp9q3WPDBhy0SvME+XYFum8p
vlzrWSThm0qd2IrU7oEclMsctIYJMhZJTVbqcMBD2roBACExLpksvZL/sf5P3rSs
5vfyWlMcyK06sW5IEOHM7tidEWgvP7aaas8keH8jtub3FAstTZR3kg2AUuup0btx
jGX45nyKCdSBBi1InP+uGzIPdJF9uVhObgF+oU+lsT9ZwUr1RMfFXzlrNzsWPAK3
npDTmznFjun6E1VP3V/mq8nN8AguTTbARvD2Itq0DvT4hxe1boyqjxW56thLGuj3
uG2yOB5ewlwMmmnNRFUbpupdhurW9LTcR7FED5XI73Eh69J9/nntnHJtyP9IxFNV
yKtJ0/BRpDrf19kv3jfnVdsJSiTuFpIuDuunYeGhgAz2t7iZshel4cGiBNK7N2D2
nS+qp5bMeJfbdCIYEHA7teyAEsJu26Kst2r4YMvLfNRdLqv3xk72Y3nvqikfdehb
FQ8zLC31zGteQGk+pWV3fmvHc7F+7W46QJM3jAxaQt7d4SqVXO0MbpT52ptLMTIc
O+FPG32P2TGO7DPAlF22g7V2bV5vwGFWyQ0aEQZEW92nDQMcE2Hdaxtl1KQqJ6Tp
eKlPTEXHMqS7E5bnB0JidfSkACzSR9puO6r7AI0MFh8SGud1lT0/vA9ccmQjRVMR
X5kTx3zXknK4eFgPaOVTKtaTYiEXal9sH9OAJNzW0r6nZM4sEvDm8zULF7Pt2ayN
TY8CespE2S9ZqXjauZ6VBscZXxtJqlS7OSQ4vgzchrkuCmf9WffOcxXZT7VuMXKV
BUqBT4a7UQ3+Yr1LzrVTU2+uSK5gYdE33lD6Hl4H6TIHAMRffR4q3jzydfarrRsf
OB16PY5pDRljqpy6rxta5c5agFRWYuHR6w3L35KtrXe6dIfSHor2S38OBUHJj31D
TcIsLwAe2FF5ijrTgGTyk5WlaTo5QXn8sfH1eBlmOlxD5jAoSBv1gKEzL0uAZpJH
8WW5IelnFO50WL7mkfBndrS22tPUTzBYx6ceHFlY8VLnDesDhUAUdW4mIvm8i2u1
193q7fhlxKDaam97498X3JvBoemNVOQX5Aio1LDIKDZQTw71ePz+l+X8n3CY9UZu
eQ7PNXmUiOCRgtw5UdSdV4/9Rrcg/0wCpG014suOnwsBc+GKNgEXMrGhPZJw2ei/
LGoIuu1qY5CTiIp79r9J3KCdbNHP3dpQDrCzb4b5HxkDihYKqeSlv+NWlNKnhtK9
z7pbMObthiaCGz+2CwsHQg+IQ16WpnWzhkfN6TtwAcZK+/btgLY16hY5ZFGEZuYj
O5Qzq6fXgK3xcdTzfT+eE86XeXHhPxlWGrwtmGndXjhvl2sfZMLV98PkUPyj4T3U
U9zjsmbB20Qht4rWrYXGqMT+cmqgVP5QPpkfMTfMiRWDqwwNlaODdfcqBfVNyfm9
Jgn9iroN7sVt8lsubKHc+mTJzIxdG4Fh1bqYrLsZdqmasbEhJdhoQrG1hUX+tJYZ
RnhwTP4krOT7Pghvdw4fPyK3LEln2itE+JLChxevKN053YFrKeQ8fYNgZa26Dkfk
TkHU3ojRjBMybhVP+ikWYj057f32yyAGyRPe30j+dVQCgylWMe3B2+IgKf33yUEr
q4zUWERY23AqbstsE+vrq5LwvLQ7M0T79GChYGOMks872zHKoojrN8+r59MYsjI6
yRZ+XOwDj1hX8g4nBw9/J6yiExX8vPs++RhXCnSTbDrVCgf64g2pjrYF6SysYZXd
0v6Ld6RIaiRsoMfZT1p2m9csH7XSEd1KyYvWaCdsuz31SLkNPXPHXTzDfeWF6uTx
Zcj+NkQzRw5fgcwBzQsuqWdk/AbTbG2nGbKjiW73EkDR0If7rbEqXCC3uWIpzQgL
xIwqX4lzF4v8ygSM1HRRKOZl4mWO4OYiTK6d6t0iQa0tN5VOMkP/1wOtu+7UoLi6
ocKZiQphphOy9jY1lLbj1m4JSfVzOxOpi+rrcAXwWSzZPEi7nVxhkXh29SHJ9Ukj
3R84BaJIB029V0Kx1dExF9yh0xjRZRXm6f/4xprGA+uxiDOZuZNMwP0DFvWVIpSI
/eT+X6qgQgvv47tvowfqAlEB9U5o9O46TKKwPj0WqPm0AJm/AtRfFbIzU2Far3Td
oyihnrI0sa1yqayJaehH6RoaqTc2NfA6uAHvO+kQppZwwgqeZGLePL2HP55VwZcv
pNXKg00Eq1kCblRwuzhRIWBtFJ8zwU/ltGmuSf7oD9fe5/DLJbtWOyFwZ3xWHsco
6vH6Iq8Oi2tEVFD66/wLggE2mjaDXLrQisnuTMBSFhBRKju8JszVI+CMD2LPg6jG
2yEIM6GXM0swjRrKclOj2Hj9ob9apjULrT1OhfaJ182EhVg6+yCEPYFi9pDktfKx
9Cc+3LEnm9ZcCEV1qmsHQRXEWg+tYMq/H/x7X+ejF1zhY1CN/Q7/M4UlJtxH8rOO
d4MpePRmrzvRPA73j/G5W8ffHpHrPi9TkSTNNuy0egKLGuLKeIBcBZyc/PuVrris
lHeXfrbSxg4v2K8DZF1j95g5QtJw/wTljuRIJAvgcVEkj9IF9UTGnryzqUOPb22f
RtkbvfZ1ldtRSjbIWGnxt+wP9T+Ox7SrV++p4dBtPYO1c/XX3IYilmLWhxgQwzPU
8VOGO29c+9XOW2bUdzr1ueJ5s6DUTaBKy/y521lTLSTRuokLiL+FxpBIHhj9FZCE
H8Znk/JSjOuqHdvi2+ra7Uuu8XqYLeT/+llUeyGCJLfUMaJSPmpfcFDAfmRUTMYS
ybVcuwDu7ey76ZK+VQ3jU0nrsiM6AavEC7u1I0mWKedosb27FTXjOBHBgRlQUlJX
JRDmFtzAwfyz+ZsH2CdYmJ+ToK9jR6RuTmzVWEFE49eK3SgnwPhGhVjcKJUqA9+d
W4jxjvQseWumyh4wdqHecSx0E+QJvPuF4qtvZKbRVScAG2VscOkVMBnQ46aIfmzG
Tu352eyfGD+UF8HFQy5faI/u/5rS8KIW+arInSEq3upzc4BZTLzC75+6eXSHAeQC
y/ndkbsK/RRS2VYZOqF+WUHd1/57GsuqN68fcrlMfAaasLP1E9hH8C6GSB1tYNKi
ClI2RXsRHx7rNoYUQ6b0By+knrjAb1viFJQQbG+tK/qwa3t9YhnWwmKspXyaqfDp
KmLrv7FWc8Vyi6DVikzoUUZgvOZSX8S6C3ZeoQEwRwEPm8rBNd+ExxR8eVsz6ERv
gF2K7hon3/RkwoP7d3vNNuR3wqsaUcLpiCmsorV+L3vCT1DQ1KEKPsm18kp8ZCYU
7Foz8tWajO5WAIff3lewvIQ8CdbKAk1j4B+peLKqrL7KRLOlKfELqptfKFlWEulY
o/B4BFSWPaTSe4TWEa4CLtrspl8OFDLt11tICfwtl+bjnbimBjH/QCRo6bddhv68
xfEJSQJWOR0uc6v5dGr0+7qxAQ7rh5uy0IlzcpYaJkJsbF2eI1tzsM6vr2sutDXE
MTWHfF27yX3lNwOF91nFda0ZGS7NunJNNJIVLANSnSfM/v3RtAXbVt3y2rZHxA5p
LhXL7GpzM0iwJrNw0aMnvZAauSZKmCFOk68886n//BkskORhUvvoqbtrBlvCEvqp
rWKRozZjkDsZ2oYcbamR2OegcydpMn2eXzhiW9c8yTJZ1QoiSZ4XIwPbfn1HzOn/
A7VS40ZBNwVRZ7vYNk9irqseivH+kF6uyoC4/qNwovKaK3n+EFhmy7AVNxpokqqi
vsY+pkxhfK7/rX61DdMM7qtdk+jLj1sCF5xSOmm3Xdd0LNBJQmy+z8xTHvl2dFSs
JmIe06IOZ8r15icaawkjSVx7Fbt7zc4G2speOMfOf+W8pv4kSJDcn7xni3XoK7hb
d+O5j/IqaKluz8t4ZiD1IHEKVN8ODXrU4uX+DWmW8Cr5vPGpLSGgTNIc3cjNpUDY
rI0yAWdOJvLXjImHir7aYN0Y0ozLHDFHBmocXRKqCCR1VQhNCYITj7OVumMJ+INr
TSUvoJQODpHC0/CDYGfYZjF5wa0rO+cHNVRSMuCqy2I6qmJ4LkeIaekUnl7Y36ms
TSjxrvCgeMwrTRTY9oZQ7k64gS+Kysxyv8IAYttXqANv1fW1hd3amYUERGk5FAG3
O+SodDzcQWUyRtIRAphf1zDrdwvnA8PoovaK/yf3Xqqd4AhnPaatfkjstRZejCFn
BUs/eo8QYjhGB/pwdIdfi3aZCg5CSIjUR/BrSbHxhCAV4JjpbxupeztuEU5IZ2gu
TW9Y1Y9G/Aj3nfLeYf0VqeyBl49m+lOo3uoSG4wLd9vnnIdg8BhpIv2bw1FL9M26
IPoRmO1pryK0H5Z2xy8JZasihyoNfLg9nMcdmmR9ax1Lk/mDKPJxYUOk4iy/9S8l
L3bJC5RYL2aHB/4UTZlZaauyoZDyqPfqkmLc+1S1jx1Id14jxtw/MbbyDUKLTlTd
MBSBq2tX/P4qYCYL7i5rBbEBLrhBNnLsEqqgjevh2ivvRZHwumZu99q4Zz4XpgVc
OuESxFT4kJ8EXZrrrANpiljVwksWQ0wWhYV+8LIPYyJgnIAcS/d0oAV1VcjQo+32
EkQ32vvwJ17yxvTFzfbuGj/0utugS4T01JHLd/uO9SVCKJ+qQ7gjcuEZYTRm/AqY
hhAycZsRZqRo8BwAsqw3jdrc6pIbTVuPK3hgk0a34vnFs+OBGPqYK+HPIrEVhcKW
AO9kqMSrVuZpzh7WPvul3KS77X4xIOHbI6KgbRqX6BUk4AWdGM62bXnUnAeNtC59
pKF3s6+sK2bZygiMLZpaVgUxhWymXO6aFpupB4dS3ldE8Npc/NlYklH+KJVqMvmU
PqnaAVJNdMVOlyXXVBBSgAme8oKpgXXwZx+yqQR2aHscTnXog3AgphPvlDJxigj7
ZGHo+GfzmA/tj56/E8LawlNBpnndiHvvOKNySV2oOLkDYm9sbDnXoCamnUfnPalb
7Bn2uvkZsIN/Gku9gvPS38+t/l6zGwzkpmPaBOoxFlY7nztiCoIyOiyYZ+5+/JAq
pDnDLK970LelmnzNr1QFarL9eJGV0MyhNofAXGRqdz7sMzuf+Pjc1QfKf1V2+9u9
HY5FusiC095axK2vtKIaJ1bRo3GgwQvs3mDx/O8sgTl0Vx15+4ua/w0mlpR5M/BP
7ucAzLgiSmuuasC4TRc5fvZhCz/kwSkqGQ2CCZXCZKwNGjbFL10Pxa2DA0hsacSz
uqFFi3g4GA5gL6kTyS8Myaofaw7lN21FVCkdKBrLcSjSVc6GL8fsq8L9OhzATdvR
xbhrPUZSTBVVX4YdKClpu5tGsXXyWvHDO/oVLoOpCZFbIQ05ZWxKh/wSRy1Aa1GR
y4tDhgQmOGmPoBCYkOstvJMYsdyeNOCFf2KxT2PnQ3i1V64IPPIWrObDWCE45CW4
KPkZ6uXN787c98RMki8JrJ8KFXvjLOnnybCjZGmpcxabjU/XRdY7hRvfY6KxjiKY
Hw7oLr3x13EiLCufd9nrNvoSQvWAQ5I2jHDCmAHHGGK6soHTSO1Vh87iS0Bu2BGo
cTTQkZIBBB2Y9bnyH+8HmjZfMgmDlYiA0Zsb5ZN6RliZU7sbsGWkBj57OwPNqTuL
OuufoHovcwF9iMVqXgJX3MDWbNAve5I1h0GL0jZWhmrMtR4J8Y25l26hugqsuYQF
4WjlL80eDEEk7fQ0cHPbZZgzcEsTpQ50ORdTdAyfueTd2XuuoAHclz5i/xKPwI6M
OYbpX89gSE8oMcwx/zJ7S1mPCjxHEccyvF3BOmmxQHu9xPkZzdVjNTosyOBIDIuF
VOSrIUpP4V1iP4giCEPHZb+LB/Ssjldd+v3P62ixE7NKbsGb2Nh2ud1eK0SQwY6E
sAc6V/fL7Iav3qKUyo02FwpNSPUCAw2xxHO0K8YUaPjEo5N/ZSrHeUo+7ornkdNR
o8j4Eg7MZW68GO8a1/BV/UmUyB4YRY8RGQzVkW73wk5YTNQB6PhQ8Ds7/52Tg+xw
0EpfETzgXW+Kl5AGjOiN8pPfVdbzTL0f3ELF1TGwqBMywGAhw7bDVdbF1FKprRL1
vA7O+zA8VP8L6b2/gQJOMZj2zMMaaF/tWdcr+pGO3kxHUke8m6bNqdFkzu8t8fBN
8DsqjIoz0SKVaQPlWeTMcUPrNMy0VXZq9bYMB4Tvztf/iX/75XGtpuxl2PSLHJ9f
u1mm+B7gqWLtEk/uG61u3GAwvmdaNJnmh37W/I5l9Y/C6CavQMgDAAOs1a2AeIsT
O0FAl6iEjrS9G1bW3P87y4LAKHYedP6ns7LJSQ/oGImdw6NrhsNZDUbkzLkQ1SpX
N9ilq4bX+rNsdt98zYGkRTJMqbiz15/FrGKGx2oHjBE6vFJIJUgRttgUBw4QbKM2
Nj8o82ShnPzwLzER+cxg/uMRWIEQRqraKZ1wffazmL5P5k7MZMGnXhuuHUd2L1DR
1WheUgTC2vcZjGYK4aC2uQWMGrs57+gitcfDYxqv2nN8y+k/63XsN+rSXfWIZeU+
c7FnOObmaEJgUx4Nu9ptiVVZGA9K4ozS7ul8AxS/OZvQt+bMQLZJdcyBqcWfIaZ3
thBJIKSxANdsHRKLr0X/i7U8+RUCqe/QFmdTZDFT0XFyrsGtPT/POF1nVMD3FrL0
mrqWFrdGvKw6PuXkpAbEG8qA78QbXO+t7Sclq4o0e+G6L1M4UN5teT55S56i1CtH
/yfHfIfKJf9z93FUk+ekukF9QCL70Ca2taQlgXR2yu1dY1tonJz8PvQJUa93FV8v
NSsqpzTMBdhm9LvrV4auciRxzpyXzOPPXxTi3LenNMNjZ7PKtj+zF960kmRIk/4v
24tBU5D4JO8wn/vzyMKhEEQH8knuMet/8PLI65bLrNrASKI/kpSo8jyBMY2KFIGS
y0U5CJkfpT8YjFQeb6P2sMadou4HflsTcfb7th9Xwhbh1BclXYHpgiaYnwQVLMbw
Ti3eyzEpnXkCbz3tpbpKd3zRcrOLG3EhRnofUCEOMaQGAgo0TRdVZjkClJbTaqGk
1M/I4hVbZxiRe/MKrHsNqxRcyaUleWBCN+vZEOvNnaYsVbDejSDNtTDNlLsEXRUW
JvBapwjKSKhNMv63Cfu20d7fb491U0m6YjBrPxkXM6ThYmIEC7z9Kq5LOrntDwer
LHaVwYxlrFJ1kPiG0LHeZI+OaPoGpM1UPAdWXp5EakCqZiWJN9sL55Nt8kq3t/qc
Kjk4wDMfVFeQ+ojZjePvhdJ/fJh9DxEPTrllDHZvzYpTZ4/q9syIF/SaxqdE4ZqK
Uy4RSmaDOff5ho4AX+fWZhOdAALMly8sgH5weEQXdAeHOwqoBILBdqgn7KOmOAn6
JFv8bpGfLJf77quyYW8nSOaeQXYBTVdM6nsWYr+5FFa1bYAb68bmroWwnBTUTwKb
iOqeArGbDI/4lCsBZP6Sy8OYTa6v0sB4BMMxQOfwWr8utf+7X2y2Wqm1abrPQ3lq
8968GCA9HqlVqm4PiMyGzvbGKZr8QrACvang99ufwS2ktKaieQixfbaLT2fjanMj
W1ieyuzEDmH1+RQwV9HrkIpo8dnLBFBS7p4ESO8/ba7LqD9TPHIxrwXWKeClCxEj
MMyjYr6VwuD8tUnSKFg507CMZaOdJGwDEWERDkV1ZIDzLcWrGFq5ja3xCa/7NWLx
lAHrn3ziN7pqVMHcuHIScQXj7icxKqet0jLoCCtBM/C/G4imt4A4zETeDSa/7waB
jZfHD6QH31wUnfAaxhqc3vLNdJRBGwLhNOuTYmXK8Eo1Yd9QbY+Gfgot8/73eNqC
CWQDpqcAn8k1ZMXJbuS03R53tTLEtwVKRNg/hNMCs1+u6Uq24lP4UkGcLjCTIMNr
8kBANCBZyGL4n6ZswUFBAPGRc7CFsJPBwhrQuPJPm2d9I0gMlR4YIgH65eJAu5Yl
EjPFuEeekIuoek6bC6kfijUpPRIeRni2usqnYneA5FiBhK9CwFnEL5878XlLRxD4
CXRiyMERkRmOs5Al1qcOQ8J/9CeDy4LaiW27lHJ9cjUYjeQpdT4J44AcTDDo5t/S
asPPquv5frzfjYQkAyByou6lYFjbtX+QAzVch2D0oCiDXk1glhxIfrwNy7fHg2H3
277nbPIRvuIAkalnW0zfoxWVMypvyDpEXGhFIoEHnWwXBJCK7YFRNor6IZJ13raD
XDQxUzoJ6cEg6Nv6goyzC2Wi6mInFLk4ksMMiSDOPC0B2hmYCg+x9gLZey6aEYOJ
Im6oyhz2Vhshy0khrBVb0PrZRAHO28Kl8c9pyq6Zs5lAuvWmBZBnOLBdQq5X+2Tw
dm9dRl7MngGpjPUVXGvL+2Dj9a6R6MXmE05N1XfKzdz43EqaHmaMlqT1jyKvNwrs
sMg0HTq67sLt5Sh0psDL3Ajoxol0tqESUNzHx0U11RQH+hvCwz8YKsw4OIJvUX9v
zlfeIIzSO3IWJBeG3kS5bsRiNYsWBALTLiFoPvKCooe+OvI5BW8dMBb1VoA65zZJ
CYAZpv2nABaS7qyPLTIaEKChu0TmuTEftMImOIqGkSDJ1TRXqGu5XrwovidQItt2
sazdOgG3rimCyrKHAADzJZLYhwWrT7oP9WCDKwONov6JzxLY8HF7xGuzEre8+JN9
dl6vqfCGpswrHCv8VQXYqIVZJVKIBXkg0mlUNQsJaIW784VLvhHqugeimkjdl//5
XtM7ePsWVZEaLhOC5yI74pI4/w1oadYSSufkYTJbfBL8HE8+Da13sd80gR7IqGNJ
NIQAGHMulqdx/16Imj0VVURZeolI0/8cg0NWvlP5IiOYe43JKBL8eIk9SUiTu9Wp
KxNwx4IVATv2wBHN5ZrqVAr9tmuOqlqSl6i1zdSA4IUJOuYJuKakUmuF8T/+Sk/9
UD1R3uis6IGEMNn51RvRwliwcVbAfG7n66+a0g9gqdtM8kTagraze9rWgQ9k6S+k
ZvOcnNTUoXcFu75cyF15jgv7sX3cLLmfg7LoSEeb/TVbCai2rpt/m+Qa1Ex+rSxt
G6yDy+FPnZxsEyjZqscaTL5TPjfzkSlDmJmNY1FLaEhC75pksdeY5xIWdOhQmHeN
voDj/wn7oNW1hBIj7Zh+KL65muRRNrk3Pi30fLu1ZH8JxH3OVSfnZw3fqN7I0vca
D33XfTcrfb+Sazk0r2d3THZjS71hDT/DAGYkSGFTskdHxSqgsb+Ng2RhyrRMebCs
EjwuX3vz344uAI8B7wBr32lWK1QGpSKfErKM2C2bZ5aDvi1tZRAxTMp42poUTr3A
K1yDEH45wHyl7hyXU4jD1i1Hhi+HifTkUc4AZVfR39uTy6k+QEK1yxULIKSv4Kp2
HpJWzKX9yoYE/tvckABasKBouKuAiaQf3b2s3rHZ5e08ohOYxdbMgPO2qAkq2VRY
lL2zlC7GdFiwEkBPTowQXSIt8E8C3CQfnQByZ9QycUjOluZEtz40lBc6hNAz09L+
KURtZkwuoM6f08+3lMqvf0E+0rn5D40hfl488OBwn8GcszYG19MysvcvjNZbygpJ
k202tqhj906mcQ4EOO7psMPTg+1yEDTTjxwVa1WLioI3mur9lfK5qd3DqgbSLtJl
8aE9X1UD05o7Bbh9ulKWmBd/+O4nt+WmYAH2dgxZNIpkyofzX3ue5Rx1PnMZM2xN
yq4pVFhwzHouo6vlfQrMuZXD8JOa8w39IEryncslu/6q6uYG94bxztsrLQlNoUAA
j89mmwE4MGyWC6pYwJu7vtED070x1ZcgMh3acniagvlvk5yc5aon3NeJjQc/VZjF
GJGlmTmSFOAYCIa9wsiBIvmJPB9AhadfLJnwvDnZkRUXXWbEypnlDR17LU5YRQoT
xW0E9Gy8ykdlaJQvajG/z3u32IVEHry7DLHU+ButsI/PI6eq2KaqSBsmOub8T+kN
+Vsv7C8D2gYzKIMUg5B9Si8wNW4QmXlx+gOfkX83h0NrKxPmt1S+DYGwgY6Z4fwb
AvmKW/5l6BxvBX87XjD68WYTUCxfvS8Eo+iif/9eaGe5Nx5kH3JBJDX5sVmm/KNH
JD/C5RhZM+1m/5DRnrmCnISmPoQqXIIQCfQ6zLOE6IKqSoeNxp8WxQ9KUeJ8r7bV
vQQrnw1MPN+lLhdigmUhOacih/N8IEL0ouGkgdAv5guS5rry18OzXVRuvJm4kURk
HZ85SRZAVrkoaTYTjzX52/RlD3tebCKnyOC7jli7hbWcYoQMjyd48LANb3Ow3sFD
YU6YrOhJ8kb2WKTQsDc9UWO3P6XBvMee2qsJ1uyf3kzyXCUMPRc5mkk3gbgN8owO
jzWmNwd741PETuwqQsWNr/q0P2gD3UoNzKEP20vhyDtBhc58/Ei0J2KpClfC1cKv
OOk9bVYaY1OSU8fPSGt5v//nZtR3cjmL455SOasbJ/zGlER3EevYE6CK2wA8cgwh
e/NAJyl+OSosQtQKZ/lHqQKQfMlI1G7XITEE51c9Vp6+8tLKYn00VdfN1ZetAFAP
yV7FJXwgf1nlEAZ2emMRJeDJ5+Oe8B33DfupfMWCFlyt0INk7Fzmir1SNMSuBytH
wOLWMyWbo3gnVSibKBh+a//1z3DTbdoW6cXnNLjRzl2Ol09sS38iU0RNWv4v/FXx
kR7gO24lXcDfDLTOOe6KXQFUBntGm6wY6oWQwgAKv8HSYKIojUB2LfCDaxy3+OPC
aa5PnQNt6w+pZZn6tPa5KDbLkZt1kE6Loda+7dNSD2Fq9h3DOBsLlnNXag8qG9T8
XAMID1m2T6/RcVMN3+NMs9EbDbYBqZMM5eWlfDrwcRjBspjt4Cz1phwzwm8x5Pz2
JrMkUejvA4nafZOi/5sx+98yvJcYIpjJyMiin857wdyZPYzlLEocu56Ej2qx4E/8
0vgTS+O3ZzMHTb7h7ktU5tfEe+Q0hRWCMvPb8TYh0CakOjNJkuicK1uT7sQW/CNS
JZl4kiQnKQjvVSPRf1F1Pnhj+857NUKh6HBjR3rPFD57LISbSLxjur9aAvyzVbhM
ZlDCU8L/RfNmI5OTCQ88WVlBCTSEG6LUcQscN4JTmcOeHwEsfRhly54bIRJlojxo
yuN8infO6c0iwmQqHR0MyNAGfXaXUUFDGXrc5UdkGf7YKelgE0jHx89yalZeM4dB
5oTuDtWvh7dXxoc5KG3I8bmhhCfsbbQZ7zstJEaMDuNTpiSpD2MhsBzQUbtPlTIO
hSMtgYKDKGno3ilhEcDS+39Teu/mTeEGWz+duc2ddewdWa1kPDVe+UMFGMw7s1xh
/Zv0FMVkICc0TPMl3zDP3JqnLA/X7wqTtfh0V5m7INQWcYhuQHR89htbxpoWUChh
5U0wRLFI1H8nWoDsWpT4xyev6MoS1lJvxaQR9B1l+nBRUnRy5bZZXG4d8roI9sJf
d1eG7h2pwfRoazcnRaF0W1QC+346CP1a8TNT79e82+2JDHzECWVetEijvvTtR6hq
AUeZ1q1NMWrV+EbGK9wNf5s7/zS6ze7Y7wii71veIj/sscxsWqNkJLB6mhvBAVHL
njBWIeX5CzKUfQYAAOHNVQayw8lRh7y54og8RZgi+hXt660LVjOm9Ne7OwNWDlkR
ldo0XdFau2HpME+ljoukp+nRxv7tvw6An/tQVtsfJMFDWNQG7xbFNxkIYkY+n4QY
jnNHYxp+bu0x7T3qe/dV0jNa+6v56fvpganz8l7tib3M2zd8QZE4zHu0PwXVCVaw
gjwDInZcvlAe5esVqO2ocOsBcQuzN2cWlwSdkWpz54LMWwhCDPvcjFFaGxtj6KaD
nnJGcJd4dQ/MJCyW0cB0SpBEUYOiwjDQDDr1AB8/gTUuXz8b+2nnZ9bI5XWFGpj0
C/fgScu1ARKFYo6w1YV22dh6V2FsVh2slKct5Uyt4QX7c3zG3ZlpBh2PQL3Co4ds
Eja7mDVBgIjs3YlKaU9pTNHTBS2RPKWJC7C7fcj99nsmITzMk41AUuBP96vlRrgP
+F+es94ffcQQZLEu9LnzI6b3MLZGpZXg0K1Lif10T9yg94n3vq6+qPmKJL04MmyZ
r49XjIDoNr+QOqM2FUHtJFV4axfHHPdrcC1r/TrmlL6FnzpjnfOHix1B6CMaL2aH
+R9vO8eBM4UngRT/M4pD+WZeAOM3ZKA7QxIAd7/kr7NVx9bwFq0uYNAlrej/zoFe
4OqY9dGPytvsLSXSCWVUG4NRPcyeFgp3D/coyO4nqEswUjfwgr9aKRrISswB4tLF
YR+ITT9pQdAwEgDtt79sFDK2dkjgVOXmh8EagWqa+4UczpRh71d8m93CoukbLDva
1sOG4RzHGHEygGfSf+W/m0AEKY/W+3NJDcUnm7BES0lli/o6JN4uDtmRfVAGIUov
4Oz60IrkGPze4i6+2E+7HJ6NHOKRi+PmPDiMS4OgNJf/1PQqYfBiJDkHNuJMUssn
vdnhtDFve5C9tOLFc2tbIiOQ7k/1NJ6FbHEaLUan6S7nQbmpFkSOT8RtB6sVZeP1
wwAonIwo0d2Z2Um7y+cY4Ep136Te6toDx/O1QDpILT7n7Tt8Ei/rNeIObJ3ZChEo
GwsnsfgYaCrc9N8y0a6aWqOLEu4i6qPhpmz0CjhKz1PooKcW5QyqloW2jJYJzlgM
stTgj5ec96mKCLbQHzJCu2OvPDPAWW8Ft3xbEQRthP7Ww2r5Ckq4RST5GK0UK36t
OkB9mAK8zgctNtAs7Ak/bWaSQzK4QyYr1UdkBUnS9r8ZODggZt9M+FoB5wK3T/RY
TCCvQYtk7cANsysiDQRo2ucCTDsv0t8YLwEvTL1EU5l0mwkjPRYfQ0Y80wOuISEE
9IH0KhaGzUpIGQ+pKQua2oT02KTTAXAiqQNFuuw2Cb4tAuPoVw6qddWa5e2D7hLZ
EGCKgCe+rzLS8CwS8Ddw/Avv4AR5E/MoMh07MmCClB92wRldNbh7Ong4VgnP87ws
IM0Xoo76YcgAJxeP2cDCNBn5KciPvNypmeCyka//ZNWfSBip3s49CclIar0KlaqO
y6g5MT5l9zlbpUAwJaen+S0c43CZBLEXB7Rq6vb/BtimaOPSuvH0HHXzZH1vtHgQ
nIod8uxTlrkkELfelx6xy13WaA2hY0kAaKJCtt2Hku2ifgRzzgFByO4/+vPaWzAn
Xp/9NLY2nSPMh/SNDTHxYXIBRaCmT1REgT4S1Sg1uRacuUE5fTRZ5p6y+WN+aV2y
XsHkz7DgfryyFhlyfAno2PFyvKJBa1hD6XVplVFMuSEpq82dSTYhmV2zqPaCjNyi
sVSYioGs7x0yU5qH7RJo67Mtafh4QJJw6O4yu8kxc+c28uRZmggRqYDHFTOq3Gdj
UsOl8xpfI5uKljFfF1oi5zzIt6FPplF873utDgKTfsm1lpTZhC3vErx+MoUCc4Il
o16Uknn+9FEfzqozxtXBrUyODztEGSxwbv4mV/lSgqtfQydgU1LADoFnATPtaBzV
Qx7Eh980AbXF4DGNjQ0an9ZUykee7QyYTR3HUCT4+vvFLA4RKlWUKCQM8zoNHGU+
JFAvJ3CmNtliGPJYPdqi7dg2SlOQ2josDytO8Gg8hq83d8eK2qKOcqKF3oLX163E
HcaKLYGAQ+666MhH80oriklBqSllrkteRITTJsyhGFYcehqhZOHM2jnY73DRGpgQ
o8e8W/PYdjvCKmVOKPqrhjCOEgaeWHHCxfQObIr74hdA9QGPf9QFzPc1mj8fiwfm
DPy4zW7RgWNISa9qZ9dQtczGbJCDYCyA5hYkxiDyVxVh4YmkWtIxsrAPQsogHUDg
L1uClkS1z/vFaS1LHtVzaXxUblwSYeF+evtBTeqUxcd//0DsPf7PgMjtLKQ9/XmQ
H7sFpX3afFR0uHac8qck6RUUkF+6UoyI5TybCKr40Q3PtuoOH+uva5JYsKjgKKhH
/WRdgjDz998dF0lf90wTQAaHnDqb/424DL6mWtbK3hJjHqgyNbWQWzT0qIB3sZ6v
hZBamGKXMqZXit+UBNtRS9Vw6EUBjR9vDmWXwhV3quIQVxIH1UkfKAttWdHbqEUg
NYyLbY3w8HgUI+6JSCoNJW4gX+oKhJIogRCC8EA3TTSTJ6TTznATEsuw+8/G8ZHt
HlNLl/cKEDoST6/+LTZcCGoXzPAuzHZbfg6wXswota6nVU/NmSBd3NLRyfBGd410
FXR9+o/i1/rNIrN2lmG//tmcPWOEd5NxrWTcSzHnpV6+GghV+vAX/gEZzWeopTrW
PjX/S2Bc/wDMoJxPJcduUVnNFUVzLU5AoBArECVsvcbfsD1xbV5UdMgCzgXtywid
OngQTRer3GylgQ+z8geasF4/hmYnrbWPFDGqCsNqPGT2HiTMRCNMwdDlOvXfgTfO
25tmH3o9+FAowYh0iPDuYayWLHmlMDCL6UoJNifiyAP7c+vXDprc/n6AOxsyBK3V
8sCwm20hdBSye5tvWHurf8fsuLXmFCPH4XTlOv61bVum3rQxI6wJzPi4LFyKIiB7
I7jvF6pNFmZGT6VuwEAbxqoX6eM/OCjGb6hN19xroLtVbN2yGpUFBaMb8OJAi9Ef
h9dl+NC+dXc/thKzs+zugcrp0UwRq548Bsy1qVTsgAOnuFq+PBo9+ajyfZfVzY+8
X/iYguu/Q7MfzJsiWQTncgrDVIl2vGrQTl3e8gWuGrZ1qll13MX3VTAGmO0C/110
JSiDJTMF56Eh6QMXYbFM3s/etTfl5Fn1pjmgfy0ApRD5k3xX4KObk4m82cAadbBh
TUBN4iT/IBTjxJO2pUw1ZivoaQxb9dU242TwhfmUt4i/jSLiuvDxpCWrPbMRg9ra
9bZpZ/nfLCAF+zKd/1gpf64g4L6kTmcpK0TJM8wYOmV4qc6PcNDDvOxzznrGTS4y
5HXngqCkP/EkuaCyb4Gfp2qUQv7/L0EE3lQB0FOIfLJ2VcRqJE9/Iyw/dJq26oiP
KvmgVo++L4H7ClL+9P44vnN19wACqmNwvzk9C/DIKG0cXqUQmq4Ot6Dec6wSpKya
rMoyVNJxBqGdm2wwGqlKX2EZm53ZwCgCXTq1dJMAR+z6B43H7x/9gxi+pRfO2bzq
HfoaT4h0pC9vwUKkAEzSOW9xwy4704ErEjC4gikV33Bx9BqRLIj7Vpq54Hbp2Wty
RRPU7nh9lXffVHQll2NqfAA5+jjv0ABNmOYHGTOQcYWg57y4WnTwZi+ezcs92QAG
l7nOpexNkOU00mPkC04g3tV60LGq6grSitn/1BGf0KlIihi80EYLFMiepO89LoqU
koQ9ggvMqPb3CLwxiQdFDVPzPgClXxubEu67WXb50ElF94MNUp34ouy+9epJTv7x
Eu6WIPZFkQG7hwKhz1VfHR5IOXbQZVhBoMm1nGAot9ME8bfbI7zN9xIBxvagoXhA
Xtz92g52TRRboCSvuj9UNMw8CEeoPWrozs/eVi2TynnK44uPDe3PojY0a7+byIMB
9lFUh+Mz0HI/+S2oJstiim5tnMcfGL6+ENFI32CaVYKleU3q57s2ApfC9KpJYnI7
HT/WwQ8eaMiIdkOtpw+NjY/Vcwytu7Emr8ouV+wRvGBpVUDMumNNELdOIh3ItYn8
yiZvlqdLmWbUwwdFN2y8+tbXFiN+eaKbeJDliK1oYZHTC9ccp1mpQbBAvCnt9Tzf
z1LMMCstoObRWh1vwMR75ZrkrAcYeXBLBCXtb0CMEND9NEX1GAIBvP3K+aTYJa8w
GR+NVuwR/WgKvhRa2WdkguwbTXp+H4EaDMlEZw/vXRcBgYbatyuQIVXZ9V7yWfM4
d5evvOKltjwuy6B48touFrAQ3sDvPZdgiiJT/Za87Wxo0DZY2YetvNkB+539Eqe2
KVo1yn/al27ln7CYT2bgqJhCyENS4caHZzWNsooMn8FHbwx97KIaDJBhzeH4oMjU
c0Au50cDGPhq26j03+qHXYU/ekcJ89EsbK/J1o5daamOLyZr+H659AX4lxPfV7Fl
w/OuP8Ccz9G0yQE1T2Y35ssG0VfJMwnQzlrfxVXcdI5nvM4K7k9MLGzzkFy1CZv1
FhGJVT/QIbBCjAQYo4HYjhGkDgzmsFnmyiy3ov+4pDfmPFaSoKBNyLTlSFo25UKK
4nKL6pors6sR6nfUiTbrkpRNDrqyAe2j7JTH1Kvk5DKLDNvG7pW5sNkVxldi/IUO
GJbUvnHcErLxsTJSylr3xm3sVnBjSr9ca5lM7ZPlv4PPhvTYmUvLLHtR1qMDUWXP
4jwELQzBVVEVI2faabCGlD11k6EpgaaKncJBgwFcpL5P1k+BcLrGGE+TwpzpZ0xH
RW37L1Qx6kyksNKJJUecRAFb44O8XI7uBLP5EjnySO6vZ+gEu9Z9zATzfivGomiy
scojcc5WSiABFqhWdHDJPyRkhlh8DetOqh2TGajzn1YxRMSnxs8YQo5UgwiMCU5w
sf071/rSLLol9PP9nJxwzEm7oIRnFnuXrpDeUvnZpbdSMNyRgZwSIqCX187ma7KC
W7C2SIAZsaZ1HhVHrMjRcWakyrOKmlg1y3OanIF30dsv1DMxzygWEsKU8Q6ykvvR
uyASncUseBMZE5NhLG0FF1SJZtsFVf5Y70aiVkALQam+E3boeIYQW+JO+U1rVvQA
X+r8jLavm51D+ikFzhdYPISu2RUxGMyfTEcr46ckmsGBsGvdkH7B9vcGcpuIZYiv
kwnM0d4a71UW3UGnIj9OOtdunm1GfVWk/DLfAWnB2Y0ZSTE1yPimvRIALIQqgEIv
2BDi7QcMXbcFJZK5CyNgqdZ67N5OpE2k3eDjAvJWSWwVQ3hBFdJ62CctAdkCDFbu
AiV/ACsK/0o50bzGCmuR3Bg5ylpQicn+MAfot7oEd2zpneQ9101aOChdNgjrh6k+
/yav8ADTShM+5lQ/ib5EUC84CldHQBwiwXEvdppPN6mqVNkdQNLdawXxbUwMwyrC
MTQyvb9UW+QFCzOrljaFE5AQ1V/reeibCmDFFIVP4k8HiUgm8j3cguRBAfSF7kp3
Tmb8xFfcgkDMvXM8w+dgaFRkX9756cjYgORwICXknfe9HdlmlvJYRg9HbLIM43QQ
o5QSzkgYEpivVl1Tt1HyYFMAntHcUFsdHht1JFjNbb4M/cYj72HKdNQYF74owttk
2o7heH/mb6fnx/KTEtXCqLWSCPjsFMUCO94rTl5ycfZ+F6uMXgOwLkqmyr/nXtia
6Qd7gPgpHLERDCzvcg2QC24vSJ/RUIKQlzAzB/+m2xmdmDqZYH8fTeDirCsPTA5q
+OT6yDnwD4MJFLhDxcZPmuHSayQFuEy7xaF4VkFm46uY9GMo3LXnak3jGil1+DiC
n/3IlQPPi039l51DxLwJkyE9+xIrGxOTzqQyPYccJ1aSxULYNsqu6F8jFsaMFyME
ghct6sSRQM38i/bmgHFIQ4vCYcGi5i29qvXwWOy3e7hq6ddchSl37kWHuttZHduW
YRvgg8NeAb4C8Apex4fpetUD1nueKAxD4CEbvYEbNGLlhSuWQfQgJw4yvz877q5D
HqSHt7hPzZQm9rR8r6KowebqZtAJ+08ThXI1RyIDandxpANdjJobRfNkshIhWJst
iwoXG/HsVN8cyOBMaBnl1EKolgF65DXA7DDjYjy42CiWtzTf1xye+vQtckv/TUdf
nQUIEnM9h/op2+VgJ9zMibNTg0DuDL947X7+wCEtU1YH8QUnE6kpbwFscfh05Yhz
KO+2t2RZRYf2DH/O3kHyq23RJO7uzNcUPdD+Uq1E3h76hAQzj0cDTHgLu1icxbjc
VapMqRjKM71ZwEAfyAWeomh8KEEj97VIOw7EpWlgm0UQFd8O5lnNFTBYPrLNqG6l
qRC31O0rMOg20R8xILZ3pI1xD85AyE5Ugubk674N3zo5Lghj0fHoMev2UKnRvlzi
EhKL2QFeoDf3c3FLXsDpX0GoSTE1K2w1i7ilVKoJzHrncFysFImRbORXZoBiu7LY
7tNbmNCgm3l1cn4WiGN6w5qn0udClXPjUEE+QUELezjRSn4JS2tSpFB5CylZtZ3l
cwFqLBU9FUJFejpBMFEoZMeuXQvNEJtIFw1NbOHHjGRbk+a0nemvYtu94W49m/dI
exdhbTYZqY4mJeB3EcMMizqRJd1LxKmK6uL7xyL88e7dT6y46iBqAGhJMP28AmIw
FZCrbs+uFuUBcrBZwRosg5E2tuT17kT2nSVaqc0B+O+ZlrsLfeoFBrGDvffTQp9h
k544k/vGpMaU8jn77RI2+67Uu7DMjcFVmic+WKZ+997/+xrJHQRq22NJ0LPYC4O7
O/3MsntrD/PADc9wEg5uE+Lu/w9ymBdQ7hjAbVpIBbvKdPJzya+vtUytRFu8Vfvf
a1G6FpyFYaupnjqm7i6LCCEt1p7WHDMQUNw60EjFMhRABXOML8gmhJDb5H485Zdy
cJLOhIKWaHHeFdYrVIn/6ayynQGbxxvpHsIuinj7RTtVINH55PczLkMnWJBkZwmC
OjnstHyRLMZidQxPI6Fgj1BnPyo2Ivz28khRFiIwoVchNoXLwYPj9P2JHO9y6Ou5
ov1ea0h3ZpzYM+1nxLeQIlHjbfydZk4A2ilXP2MGIb0ksOCGbAKpePi3vPr7VGaY
MXICSFlxbr/8GeqvNxstUmkKJa0nyRe8hhFuIA64uzekn4ijysqinhCtho6vlxSs
eT96Q/o/cLBNRsejflOwE9N9T89rzEIRgATTBpqzKElgh8KsJPpfmZz+YXN31/gF
R3qLtYTDNsz8stIHHJQt1ZHu5RD3prKC6B3Z4qPuXmqLr9q9tZfGBRWp7COnFVIl
1WQ6bIQqdozxyO6HAFXT6WXiBaEKpq0cazduqmviCnoMENVvUAm80W4EGHOaC8E5
ymrlEhBOfnZLoUFN1KLmb6w2B3aC6QqeLJOqVsybvA7DCubyylwdnvWfOUQcpaUR
NvHnCD7Ot8QM9qCnOVW2Pcvg0O10p7Iiqnzg18OGKUf5y3RnjBughQNYZNR1PbYt
q+O2cPMnkVz3rrENGVOznTsLxiusdu4J3UmQTyt8sqd8CP/5ky504JYQrqEKXkiv
5s7pcyoW5DxvWgNIMnkDKzCkIOESF6DP1lXsbOp/Xo+UZjaamv3gOnmgf10Nyx9/
m3TaSIiynskYxT5Rcf+FiER6eTdIBp9zw8K+qir3Z+jeXH/kSglRyOGeLcheCVR5
RxK74+eukqeWaDMfggA9bhRWDc0mSun5aoyFY+izwRnM3/srEk5lM5Yo82t674YI
UgnkU59ouQuIvAasqE0yRcPJnJ7+tV3ninLJKgQvN6YfzFoXnxP3l4RqwhfZLKd4
TdqKJLVYrYpyK4VkhHUucR9FF5bRbP1D/mJW+sSUHhdcTltMN9XKwtrF0Jf04FAz
MK2GaECoUIm06vaw/OojRxz/QQgTTdsnccS9XlHu8ZKUVbvcKqlggKMJ1JPj1ZMY
9UWO1iZ9hNTbVivvbPHoP7Y9dCrkODQq7LG7Z2zAk8LWtqXcQ8Nk14iB4UDbMyb7
1zcMd6QBM5tJ7TqNSQdH3aZOjzs1628mlU84TIAtZKzvunYAR5frQbj73UsGkfy+
hqRsO46hF/hLy2ReCWOPUjyNO5ll+u0YlU/emYkmzUrVdeXFYSyEfqghGNipxYQJ
FTcQOHnnUW9IFe7eHbaLnO9F6kV/Ax6THPDSbES2A3NKgYSyuYVGGC76gGG/m+8U
RD/ckGJFckfLD4agWXuFpDEtL6U3+x2AXy7tDKIImcc3IWx/JKMUX3TC013g84UC
mE6cooc30ksHrZzRz6CexWwo/+V7NqYlWaI/sVEUT0vLCkY/DYQzoRa5vnW5iycd
qndG3ijFLqzoR6ZOK0eU4AVDtBeZHxXitQYAA2zHLXZrG5jGq52nri8+/27VFkVE
SlRag0AKb4GpBdG/twKv82+bihnGyFeonF3ePTHfsPYo0txdLT9J/OyXB6nXeRNx
j7FNHdwUnYok+KmjPH3JFk4WIFKvKNYmgJ2kSrJfUXTQhogzfchBfVL0IVwkGcVX
3jLojnpB2gDGgzRVFT9BlCHID1zsbWLr8mgHjASk/AX9V8XRVF2NH3w03khPH8kg
47xaFidi5n5ez5GuW6ylPIstxTrqIpnxHF5cPhH9p5Ii2yAl81+QjGVDE5BuvLPo
4R5742NK8TAMxim21keGHEOabh02v/3jASspg8SUJGxE/i8mYKOP7JfTFpS62Nd0
9Hx6W7kDwj9Vagmzgczq1t/LhTnW12DGFRAQYMvwEbvYy6MJOttunQc+hJT3WjRA
k1pQ9YQ2/5Ih00KIwA7odh/u8Rbs2mWzrTbrDw1LbfTPKUbv0mNE6yT4UrrEVUSh
vJfhTBN9t4muiwVQXddMI8yNSNYv9Ac1D0i5NX1Nq51ESAivMABGl0002vm3rwmy
qyKaz17a8FDyd1YrBEAAmAKmvql12aAS+7Sk38RuNVveMir8xwKNF1ToZhbY9hID
SEPqldY0ouI1fpvP45XivmPOJ8PNraRPGAOPQOtrTasnpmy4s6Ql4sHSyNdtaccM
qOMpDjXl/Yd5vxb8CeqH0FpehfTaXVGp7+hOVPnNiV2DhQVDhP4fvZq6OWQxf6Qc
3oLC6E2phAj+d5hVH3jrjDcRUOQx4VoRrMLkgQXNQKhLwXtQfPjMiGa1PVLCnpI5
LNZpxldUE8NluNIWi36tIaciYCDXSx7kUs0qrk94MWF2/Uf2RRq8j5XhYsYlz6VZ
CxCY2ke/cdMK5qLvt9mXnt9Rd3dMKVdq3fabc2jeTvKjF9hBpyNlJSR7rxK+DUSC
MsDYKdAF8ktn2oUR43ueCktugvDY3MoGjNxY5EBMUPkd7DbvMR7aRl/XaJ0JhLZI
jbYYZ50hhidvGk+kepkxzwy0gL0qrD8ZZ8Bmn13mZSBshl7zrk7MJSPHBGFwmPMx
3PKeVQm/ea2an5NFoM3uoGLD2PE0JEpuNM3PZj7nvXu9jde2mzK8gBTKMG0lD3lJ
ZJ5bpErxZxWTRkd01/bP5LE+apCbsv+CcDR6cLy1xrN9RIt87HYnDicbhhI8PdYN
HYuO9xiJE8X/0atjsR0tGB/FSASEvGkcCsi5EB8YcyC3+X51afJJUtMgy5YUiXwR
K9e4DWaEpTEgj/03iaFUq0AA2M8gvtmpGdMPdcjn7+HW9rMTm9qZ52kxg0YNewmj
p6p1eAQGfJ3DAOLUAiv/qz7hRu56XoLs/vY7DftJF+wiiGdVEaaDWI0MQzrOc2US
h/PEgpjvzquNPVTn/7S1QZ0nXaTqzvVUUfLBkr1E0KWAyzBDC4JUnE+mPEixm4mU
DdcMulIFgWXvNRTXt+Xw4oSqnsZjRTBGuyXYYC7jlem/2gX1qE91t3IuOzQwWK+e
eLSRStOtjsTdQ5v9FjKOyCPZXgYA9B9v4KB6Maaii6kLrorwbpE18sz8XGSEtcaQ
AmcAYFxVXPFuqGVtK7gNhOxxivV+o72MJkGz8oSuxf72boVhv088JK1z5gyzWPt4
iYHQ74M1/BYZvAwO6hWz3v1JN5i9YffFueOoQhOIhB9uBM49p+Sbw4FzX8PyIl/t
vztUmDCSDU7Djdz2PIGRNJ7cq0r6KSgTwx9uEgoW/scNYFFgKnMTzD4CEE57ZvBn
KFUdALH+1ZeiUKJJ7i1a7koYJklxwCaoLm9ci4PQxgS/qObbr9QFIGlWEfHvHvAB
S2K3UKaEK8hljOGRRByZJZmH8vXHWHfaj+Ut6sen7HQbSV7smAGxtAg/40VH7Nt5
QOnXHCJoIq/GInE5sF58NiU3gjaPkrlwL3TQtcvsg38s/Doc3KztppnHU48u3L0r
mhlFtoi0jneVlsdQ3EgKUQXFwGqPUiUreeMKxeiEvxqoBtplM1cRSPHwHFwlJ/F7
z7V7VdEIC4Eic7xrAS3vTAGWF18Sk4rQ4Zf4ZQ7bnGadxHk7MxuQE+K/mA4c/QYi
H5jXZiSb/vHQnxNEMo9suTz71clyqOw9D53TWTgPjyeR6tAXgn/VyHLFKRy5baOL
AtxjxC/ct4z/gZqaq3rZuJnxGyhtLszsBb7YK0hs4WS05KZg3s6mezW3FsH4K96z
o3VNJZRVcVQybrMDaWRjk1w8E2pSIyDFh3sx5oyIw91f+3W3IVXxfr08KzafSqik
2yV25+lfm7zhHqmE4sKFiofN1T1AUHNHUYaKAbekdN3p5MEdMomVc8C+TnFs8SkE
ouKn5S3+KW6B0j5b250DcK/lW1N6NEMyK17TO4f3QuC7+liGcfRTgZTkVcWZxYlw
vGxDlbSSRH6CHBIDn4PL9K3ylR91bQy+zsa1uwo8zB5nLVz/OuVxA+ZjJKcnl04y
+slOIcotEeNQuJOveq4yZTvlwOCdNHw5H/2nWGO3NFCj7rFYFeTBAWjXz30QmW/3
BGQYJBBmidbRfmLRlS4n8S/B68EmI2egjONiHj7qACXMpaY0hgZzEbtAt6PCOmcO
wjta22jQxgeZhcASmJ+lgSvO4fyqx8Tj1QQwr7ryzI7IiwZoID2Lh2rhzjXPARLW
7Lr+8kz5aN/DnF8pfqdeK2GV0fsENA4LGB15D+BIFntoZpUNy6F40vX6COEJrYFe
o8/4eDqEku+Rh0P+shrXIvrKHD9mEzAaew0ycr9LdOYvLrr8kcLppz7Pvs8rfAZy
RM0xRPtgf4FK0mykL+RCtPJWASz9TZ36OoyqJCqEw1wYQ9AXwDTaAyuUcPji8MDm
iwSKnfe67ff+0ZQrZhC16Jt7KZF3I3yiILLhSbgTZy7RlGBxEe9/iyE++xTpW5XI
/uetTaiUCQLNYNsQfvflf0e9UhDWPxF+SGs+o5eGBZj+RnFhYVa8bVpUdIw0JfIw
4T3i5kDxRlccOd/BEQK16Diuhb6hVkp9bibN256iearWI5dRbPdCqk1wZcjsa1TJ
qRf6aTDzkpj8FijIKAdcdKGyv+jy9BohfiieY5wVP71p/KRFVUxuoEsgfKThtAIz
+/hWHE9lTGmkSB6Q7zCOUppor0mPBVXQMDs2dCLr3fhlfnxtI1s9lerSVnURwCw5
LIr+vWMF9Nkdn3ZIFlul+eHOo9wmYgkQr7Fp06MxGqMZwGCzwQQ5uLi3pA8yPUw5
tTH4Om5n69O22Fi2QH0X6dqAgZmkw3DmD9Bu70nQO0+XpglgYOJGl1dmgrLRjVxr
EuQgYTOg5aOzh8h0897z0SUC/qbqFduufDh04ADwOkiAM/ly6YcBo090YeMJI+fu
COo9U+rnvspSNdYQ5M5TiLiUuSxse0RCF3t2Qp2aifwFQ1SHHsdPBBZETicix3Gu
JCpjd7WfCwcwGAUtSQ3iGAgJckMM2HQe9CtN8a8GRklX4Yrx0bdJmx9EilHYXTJW
fujWG5P12Zz7Va9ne/oJ3SvrvZKOx0dBRgQV8jWt7lWuJJuZU5Likj1f3IRaEZ8h
npQX429z6u0h9s6TjYccMJqOJjR1cBJugIeQCkQBP/EUGt4K/S0AYflyRTWlp11g
6/JI8/rzfeP5up8NL0WdDZ1NvJI22W0SR9pyYhRI2IkxwHihIqYYJxNcKHsaBwYx
xzEsciCYg/LVjt/4BXtx322n+wG8nhzs9a/+D/kJm6C2hFcrPnRGA8Nl9wuIEFP8
5NCpbL/9agJBTloGHS4S9NdVVrp5GWWIS4S9C0q9536MRz9i8/u3Rh73uGndEmFB
V20MGBrT/HrGbVC3WfgBpmM3aDojgx7obIxGUcANCDHheDEwn9ZyZQAmLZLjDI4J
ZvOa2vDuCZF+KDQrHZFfh3jzzYNGa6SDdKW9R4dsHpW7NOjoQtVpSwuiqx3nqhIt
q1LuBip5EW3v7uFEtyT7CGN6Mnok5VwkAmYQDYEQrj0DDi6mQFkiLXedDCGRJWCL
uOOfXj+mL72NAbzvI0YMQve7DV7lnnX7DKhTCVUvdWLfWKhlNa7XWWnbUmyWbvWR
ZLH9plF03Mt8I86p+YQlCIL+V6RRmKxPonu8wKrzEfJx4fbADC4jnb2A4UWt1BzG
EX1Iu6VlFKOoT0qxU0+HPUc57iys3T5G4pLHdBy9JUTILF+l5D+CjbVWF+AZz7SV
ik1ZjZ83bz8QWOtLsx07DIXecDnH46wSDhObOabHj/uFP1oGvszJr4eARyH7gxgd
ODYSeTJOF1QTbWASKSXIqOy/smf6C/OAQ6ard7AmfE5wZY30QilY2Mge8fVF/FV+
7FiqYulcUw0NjWqYgq298IXAARprJK6IudLlDbyQ0sjNPYj+TElsEyVM41caM2sb
DalmieDKPV5ui0I8YV/tOMQKhTdylyoXKBHNGtlq9r6tn5+aEh0uLj35sk1K2xTn
t5EAIjIUIJvT3rddO4D+TxIg+IK7Mr4giDMIrVQXXvBW5fpj2xbwOl6r6oXaAHdg
xaoxJ7BPNb4vo5fXc3mzHGx4m4RtTNMLianudG9R4T3eArk/KE3voFx1y/VxL7DB
coGPRiw5meP40Z0DLb8JFrXHW0oAyopvHVVRhvqkRxAKaqh02UYBJXq1I7awp+GX
T1SQiTwdCB+qabNPQETS2WoNW1/vHwijuRGdTD5BNTTBndqSTVhVQmlaJlHzpLVB
VTO+cMRbxyiPTlagRST0HfxADX8Ltoyafjyzf7/JekYdVO24gG2KdqhEbKstBefK
ywqVLxcPNxSnAzzbxax5+xBrCVt7p19JRS7AdyKhKNN/iCe7sjOx84+6XhP0qv+M
YQ2z+ujmYmoWvBALtr/rkFicIiCJ7U3teSf3mamPLYUve/fVvVxTZMdClhBZLWrB
EfBqeHJle805c2n8eo/Fzcp5P23IXzkQAkK8bROdh3A9V1hkrRTE/tZdK++IkEqn
FTIiFYSbfdxClw+6Whssbxi+kcHj07RXIilmtHDFWoKacmt8ZPNOskHEc++kBaAn
os/OQ6VSvnogbg7eHfMYsLZX0EFKLV0Aexx8oP2Ylz7pd2vzhBMkjapl4lBzl2qM
8YIEOAGUxu7l5G9vkRCRSoUOIaeAezDqeSZcBGnET9dVb9sSZcYMjKdT6cvh8hUd
ClTlyskNeAQMqf5Ck4FDU6DUs1IMhAPii0VbstCstTDBQUxTADtB65PDLrPLHMo1
TYwAm329GL+oXU8S6FaoEI0iESwSpilHS3iRZfbe47S1Fx3N1sNyqBBs1tJizH+q
snXnaY6oZIyK5Rqwey8kar/hnwuLspb5s4reVZRFzpT3pykqnhMLJvokZUn97Pxy
jBsuHrW4IsdKBFbWtbdFywukTI4FhACmHGxnw8J56Ti+gTmTMEfeGk/W+7+ebNI5
2ePI94cjqFFmVYqZoXZo4hPWlS7jg4Ru9xSfAEE7C6e0XrMk50RWDIxSXHKEAdWV
lOaTURrZWPAbalaXsayH4e9W8e5xznDDFpA2O+u7DMxzNWKgxqXiX3d5/0E9YDj5
hus/aKlVoiiIhUmqRa4Hc6WXB4ljB9kIaoH13MxFY6Hub1+pq95qbH3voOzRUuk6
wjqHM6xGlpy3A4MuGBdiI77EvFUIYThpC21uKlWiW1Ace2lwlN75WnTb//O8NrvN
wTXxxghv4F4pDX7T5NOZ0XeflStQCuPofsEiIhk24KAnn7e4ony4WA+BpdjnRk8t
UzO38mP7T6xdx3tok4cq9D9QYv7OYNKTwZTP5ln3cftETlngB90idLkZzSEuXSC/
+79Ft26f1WkdyFTvU5nOXixZaymhX2/5BB/AtARIqe1bYCJfEu2aegInlHYZtlf+
7X7t9J5/4yaen2aJplO1OVsbFDejpsmPNXqg1DKEBz5OSRcAHOQhgRy5so85Ta39
ACGFHrnJ0ss78hd0EANacxrA6oQ3TtwJWL2jUE7QLqHfx3MFlSiKTLv6cK9zGBKD
OIy/h18KnRiHJXox+tZjPaYkVgULnR4skQt8eko1vN9nPepZ1Yryi1o34x1zJb0q
8vEPo6jKj3zrDH/K9Y1tpR6MCZCSiCIx0CvyR3S+X1Z7c62uLZB/XxP+QI7060JF
h7+4Wc9WGbScmin+L1eyKfCyL5roAf6eLr/Noron/F4olFs8GE+9KKKdafCA5Vk0
GD0CxugtCQsXgLQgteYXDTl33ZhfSQKg5cqcZm/O5ML7Bh0/mKZ0a7yPhm/FOwXC
CNG94iQ46paNuGnG6Nn60x5HQqbk8D1EBMXroSvEXy+6a5oKrlQOJztpGnd9R5Ej
kbnz/Cr7K0inuCN3jKYTz9maoU1FWYMsG1ZbH4a48Na6iKcLsrn00M0/Lacxckz6
0NLTWMEgyCrzMABV+A+YP26iaoUAqEnC7NL5yiO5d48MLHRYvr0BdB/7M+7H/Ao4
VoZzjkvnPsZF2mt1azix1NnAOqSjxlFCu7sU/R0bodL9vQbUq7lLrX1Yx0scJJ/h
r259RPnBcm5HUuh0DmjfHZN3ekX3E8DkvChW6/F/OLBd5obwQDFYj4q7DZSiwzJ2
jCoJWAyEDaPzZdWWYwmdKT7JG6rj2qKTgRzx73vGzP1CJz2RuQKDcwWYmwUxSkGd
ZcWSbsskD6DXzeOiQOrdbOuUsxr8fHRCqKHAdXLWa4d/ocGX41hGaAVZRiK7eGwS
nblYXzlUqnon2/ixiDNSyX5kOqfA/hxVjuyL7jEXR7iAtggeLp1zJoLGLjvcvxmI
HzCH4H6IRgsm6R2cBIN9dQzmS1GnhJDqkfGslIsms6eP41ctkZobNs56LbiRbwFo
vJBnCQki7GB2OCopNwNA5cjRhuBWcnQ80h5TD0mhpDLsJtvoAMrl1b1fw30Owxma
Cj6rYCVRTZaDn7Z0YQcdC+WFlfUSY569PmX8AK8uwZh3M1J187qtIp/+nRakfKTU
l7OXtBpKpmVXY3tGMXv8KVlo/WyS6IY1BKU5J4BTLepGWd5g+YJHbJqtOv00khPT
J/zhBsQD00eAtknQDxjQ3xGk4xU882b+VwDNJoJZcVnHoxuECXmbB0lP7KEdVMgm
BhWkQ/w9afuFvbJPnYbaP/XVT7w7flqjscboDwdJnrkbdGgNwoDexM4ALrusPhpw
yF6IFAjmPpvphQOzmeFo3LxxkSWhMNZCvlZatb2J+tGJ6ft4qCqIroq/53zDuD1C
MsyS7zuRdIr1YVAtA84aKkd8RuYSwBm1KRRjitS5awj6UGF45K6hddP41ieU3tJ8
ydjGFs77upKNMwLiE1T2PUWP3igpL3Xblbwhjxie87L1J65L7hJ7AzumcgNpGHl4
oHqBUhMO7l05TTiBJGgleSmv22UX7XP6n9YgEI4c/IIOhnkXp336MT7s1gfG146N
GcSv9tOHEBDBSHhUGE/xSs4Ea0lJWhA1UzQ+W1/0pRbGcbbTy41J/QjLPJjy9Bpv
8rLAFiuXEYA3RzZ5iSUtX5m75eho+f6n68EvMJlM7sFEMW135rUMSqLYI1XkSSMX
SEWJDagnjrG5+EgTFcACwMBvw8H55Xs1QgZbtgmS78PANKG/zLXN3TckqdgPqtat
Bw2d38K8FK7PYDMByR71igUXMT/SjF5V431PVQBbsIgN/hun7JftUi0QgYxAmD7L
Zp8zjHZec0qwqmIpRY4rEedFWMehjvYjOXYJMAWQUX2t2YKgGR71/icFcy747dEf
ak70hREajE8CjFbzF9JZd7ByFqmZCex27JJeCo/4ckKl0grgeVJHHIVGsPB1/Jvw
g8xwyEk9RM2ywcN2bbmVqy4exlb6xc1TW6tH7mXX5QPgqF7TucI8f8z4JWJEyl5j
RrgiXeUPjVfxXy+F37RynT2JSOEKcxyjPXULqL9EpEoQ7gZLWvMuvbOx6X3v7hDZ
UGPgOR31qMwsiqWZaBOJL5BP6nh08dW7sfxaeuebfajeMMJshmbERxS1TZK7zDF4
Y9WuV8Cg2b3WwtQKpzfjYSgb+BWWc0bxUFKoe7e6xir6pk91I413G3zwJcrQX4Yw
KELofg11jgTvauJxzUfKAJ68jWA6ueMIsLOLwaYVFNV9yFWLLEQ84Dz1maRsf8Gw
Dn9hM6LuJSqPExBnyi+7hzlZHS1qxMpt2h8REiV4HFI1a19EnA0tOPCtzdTEapM+
ELjpyPIUW3qZVyH1ALlHUJbJ1wB2Z22cdOpK2cZFVUJHPJuQ31c2BiAuuiK0YtO1
SjQc0pxS2R3wS2BuloVNxylf2vZH4dtWl8Y/5CQyVRSBkNNsKZag00diOdx23HdM
U3ka7fdY7haRb16AD78gB9walrpVX8ySCGIlvdk/HWEnYjuC7XeY0X/o593ZLBmj
Apb39yN2pWmvK2Xlcwu98gEtMQEssmglI3/NIkBjwL7Ui2sh0N7CETvIagyKYoyZ
CYWl37vJUiXWt/T/NCbrqaGtoxr4+JwPACBMDXp8s89AuoNR16zWfCBXDAg+bMbr
XgrrK+CfpvyGG46nr682z0kbBDrLlsAxx5ZX2QNhqz91gWLeFamXAgljWFt6ukRQ
wym/tYb52bm4yZ9CxilNtJF6jwuzvD12rdFb5FPLQceKdIuKbdyyvEUJj+tTbVSh
ZDRJmB3mbybxODYFJw1HSAP6hmvYl2hliFqGGr/VM33aLnP+sySozV1iBjAxGwMN
JLPGAE+6vvTI+mEIepw4QVQPo6i6sCAKbt5DSmpNPr6s+f9MalBg3o8z/n9U2ItR
kXrpz3PmUyDt/4O+axiDA07I5kT9ae3cXbEWHlSxMaIoc6Ip0QUUhSdA4GKuBATz
RlnwkZ4kbf1KGEQb2MRXumwstonLw5ELBZAJHHQm/g9mby+MdngsddrY2kFaFyfj
8vE+yg8hMI4/TsRB56IvNxPvB9/grBSqUSGOBtxBEK9Cr3lrW3fTtD9JEtOQOkg9
z8HxkpcmM2aIk+KYHTc2coFrekuDWRR/8K397oy7h5zgL5Y2KhQuU5wSSulPDHQs
595mCA+dyYR4AYivt2IgXJOjhv/SDGVJLeobKf8DU8ks1+VxIeS3+HkdYVIlwiwg
rfY8E4AsTB+rMazXZzy6FUUNM8TX7hxnkUdEeAJlpRwibooSsG4KBRJ1IRRqEDJm
SM4XkW4fscRalHrX5J+EQeGYkaYyQS5tV8AxundWlH9/7Fp56o+8tqX81GjQCttF
JBsQsIjyQDiUXxDAbORkM4+GgfeAuJCCT+NoxG3LpkK1oWjPmjaV8YfB5RWwRKFn
+5bHdyYAY1cpQIEFG5xXisL7gWsUROHp/7CJrNKXJ01rIk3LuVpobqC2LQhlIQCo
3sn1/tgEK1z5OPIvdjo2ceLYmdiZ+zNrUAruJys824SplGwEhHCigw/JqVpp/QM1
mC0BHjXCCaiqV9TMQ0ZhOKgMBhAoZIg88kBO69rR3vDyXBv6yRZvqop1E5jX9pKU
UbVtODDYpSs8tsHaf46+yHWmdyC5KwW7Ltol+15wHhAg2yZK9A8Bx/klVZ24XgSG
TnmamU1i4mR4W7KDqfkempwtxwxb+Pl2WyKPboCgdTkkYGKXwmv0C0vaIXvdL4sL
emibJZt8ESXP0s0D1kiqBEIk0PGktLqnRt7grbXIKaa7GQSmJUjIH7o4ulcqw/qw
DhW/N8I8xCea2BOdhfabvDbjec/3lI2dt+6mvN+NP/xrdxvyn8Cqxe0/MeDw7oUY
XGFtic73SXnMMOLb2r7/6ik8LiDsWQnJk6Y/mvSdc+tJKo7DiIrr/Nng/KCW1TUk
tEIm8MLnnlxWgAaRCjKYCv1Jw6kDzzrmYs70ZoeTgnvEcATcnagDGth4MMIm1Qum
r/hFs9lHlXeIOmL3x4fIB81d2I77BFkm3x9jXDLs8NpP9cWS9W/IRCMdHCwInoSK
VGzT0Ga/grJWtHtox7tH3WTVrD2MVlfwI68L2UUWf+Awh+pQNG6kCSEZlKejS57Q
53lJzNCgr4E7yA1tXf5ZKLq0Hn2waHt2acWRW8UewgnAP+eU/v1QozTC7/8FbjUW
vQpMbu/FTZsJaPxFDzKaufp40HelNenwTO4iBYALFZiJAj6URD9Ir9Oo32jPp+Hb
XxacKEGR5zZnXJMo/3eg5F7nIPuKBQobws3Mn13PBItYpSJ3G8slukgMuiPVLJRv
ZCGQy9se7Zy7IDAey47FcJUARJU7k6w7gtPsuobnZZBuvdcYnqcSDMhXdUcjH6O1
cWwL/OAC/SI8Wkp+tlHmJu0xsdfgdfpqq6SHBY/FoKj7m+Irrah/4NjR0/iqHhp+
12ZUGE5gwyvW36o6LYuV05ZBra6Z5R7HaxubOMw60KjDmzUzCqA9YrP41qN0re6b
+lk6PY0Kue3kfMb5+tXOivZ4J6UbThMKE48R3ByQfTnRFKpS/3jXPG/JsCzhQpHM
j8579wBXEEmmkODjFxrGIBzMNlDdr6cB+bt3DcQzem/k2NBIcj6G3AEvJIQeS7P+
+H2/23JmjuOwSa565Z9brPJWQFqfvSajHE1GC8l8TTZMtOcR2Sz+vYyhLNUx/Mey
/qEsuLC9Hfk7bfJ1a2oqDQAJXctMYISjHSx02HONCMD8y6opOxNbGddIGpEtBh1p
Bq2yG13iqQ0DpubCh3MM1Unt2uuY9dd5MJXiKvfen1HkAXHkZeVEjrRZbT+ME5Vo
raS6ZCSPTtAv6bphsM/TYufhprcbhYMo1fATgrTkUBfpnNLtb731S7v8S46jb0Cv
jq8dSZDooCc90M5duu2mlvFiYr5rl7Fcw02HQ6IQvlrXJgovhyvE7PPHX+6XiPST
7K8MUbz7hIom4OSPgLBZkWuj4VYr0GFKXpfddPJWvde1OlwOPJVkbIgFdbR2X0xm
29yqh/upYZRFSQ3e+2YCpx7ldskKyRSwSRRHHhwq0Ygug3BoDbUX/zR35g0VSLsn
dj2kL0xHMjSq1v9jDfIZ0Zd2+IkiVp6mFukzeVNPfEGJrZI5SKTlX+9btEr/poVb
5WJwdzZjiYL9to3N8Rr1Ts67qRhGNsu059Bs9ndl0Na/kFZvYSWt6qWGdrAqm1r9
ADpeNvDNjcm2obAaVfzHDeFOQOWjb8XAZ8VP33I4nw8WdKSiIgCCkNXbqehXFZhm
EkP5c5AwubhJwEvHdM9cZUVr0rDGqozi+rC3cKjUfV8K19L0GUQRslhrroUeKw1/
yU6VLg5Zvtce/vVkuSEAHbIyuh0DCkg3dRqkh9TJLpIr3dk3YW2hKlDpS5g74FCj
XgVM86NO2BeBy28zuJ89hUmWHn+I27pYux9qfWGZo6Vls59Yt/XZmzxuKqsJxAWY
kJ8dyOai1l1rYGXl8zppPHbgd3FJLCjKQTeK0NvAwQfFjny63MshpjENs+a+5xFC
UMC1ZPPtzQaT8s6COtxgH1zVEoouxNDrVB8K3Fbtm5ArF4Kt0YnCDXnQqymnH90d
wW2jwmpI9iKfY3X1T7maO685W5z3ZCYKbKN0Yrahy8jdzMXLIS95sye/wCQdo1Kr
LMMsYl/00jtGGCjveWn6InDF/uCyrbMgfSSIBAuuM92lPDvM3hjjqTJwfuxeRgXk
74gia7qzLCVf4STxSUNyYtuPtaCrmIEIedPYyjttbLK3Yw6i5MC+yYK599jjYQqO
BMiPHVlaPXnkcIi7P7SWJxurexcS99E3nnIjIHEs8dd5iYd8+bkHEy0pA1ReH82z
rW44+EH6FBjBDC/8eXHRqDSXooINltBR/MdSbbqYbWtHqLTg1K7imzY0nNf92wjG
dGko9fZf3+fx6SK3SCWCesDWMN7Ko0nlCYhHYCsi6fyqGT8x8CLSU2PAyPGLoTwj
SswFU+UoiDmw5p1R7AmOhA+42dBe9Q+Zq9e2T9Sko+ehKEdLUTSu9Us2U6Sj1/Zr
sW2q94p7Onw+rsU7plhuj+VpeivKE3rXjv+fsskA7nAf6n+PCkUHDudH7aJKVEKX
mhdsHyKL3AQ5N0P0+faK5cSrH89wWQK3uxU+lreL4dJRd9HTfK7/RAltdCq8zWFL
I7TJxgTP1X61BncHmKwyMim42pjIcKsWJRuoHVkjmXF3YSMDzjs/y15MafYCNF0n
9bJUxjjsOQnpaDjOwOonpkqpY+cmquzYo67bSIfLQyI0PBHVGJ41tOKLexT0vBod
BlnXo50XhWnlDm6D+bzycQf0TWNvDoMV5XrJ3C1KQc8LISL+mN1dK6CXH6GoaUNh
vSeXxUwCZ6mWFYV+pt7BGdqH11WM1VBsJGl/PsdFH137EbSrKUtsDfPzd0iBTNLP
7RskoKLsWmvDPo8V6AIKfcWTJ2702HWlcDWt24mttFZZ3nrW1IabcvARJfHPAQEQ
FfUn4E04NOVUTuSkLfYGB/tE/udIvJpztTviBruXiGYST9p6Bsw1K41R5kWQeUGm
PNYSct4FDnSXpOMqG72yOM2+Wj01O3CrqHH181P4kfWt268ZDeEFSakO1HbDbs/A
TOO1XGoMIISUiSl4d/v/sx4naNMub7hKHMNSYatvNfgjZgbXleAJQBeps8s0eFYE
FNpQQS7sLZEGqwZmIk3Ayt65ji7mih4XD0eInpIs2Bs1WAISj0aqgA/Re8D01lbD
HaO1J2ZmHLnlJGv2VLtsGuNRRADGscjPPEtKT2Ez0XyspCZ4tnbjTS+OU3UCQveM
kjVENhMuiCVJzm52VSVgifGuEFbDtiCY+jCoUzUhhoX4YqrPYOTuAUkPW+6hSRS8
8i2m3d/Jgz1GJLoekYWB8GCe/YOFC/Z4MIhgxCSsB8kqEAHQoiEe1iD6x8YAX3sP
Rukv2plXgwo4ff0dHgaNPYQ8UClQFQL0fABKGj9sJyqcat1jhCjKVSbbi6cn4r/t
/THSyqQk5X+DZobKjbxFRGdEAkD5TglDAFRKvbd5UTwew9rrbW/vd3GOLV9Ith3f
qRUYTPs6z3+5U+b6xArilwYAKECYOX0Aeq5fvKXKYLSUGFFjLVXwo3g1LBpQdUFw
ab9Zb350lXS4YvKFhJGBZo5ey9CitFfDa5kLH1MiFJjqGQWT/MYPf6ktA9NmfNOA
8XA7JD0z09svTdtinY/p0sCS4bvwmi5JTtEIryl50JK1UP3T/S18JQn2vIS3MoUk
Dji0/5VICQi2toUVZkNoL88jvKEpkgJ5keB5Vlb1TYJcKtcXp7KYaYfqCvMTyU2f
spBVt4g8FYF1mWLySEacpG0YGM1s5EFnl36XHjzGTRH2QaWJmmHnqGvkzkfD8ACG
KyCt+EgM3R+JSvUMGKRIqh0C+4tBNEC4H7O9EE/KccsHsvJoI+h3n8Q/LHBOklWO
XFnMKgTpVtOZzcJmupMEa3xQvISFYXC2fGPyShQxBFZlKI+vZxJjk89QiLAh0GAc
cpzA1fPlVajUJx6uM4ZPtJl7kb4+3LMMFH/we7PmpfFSFEPAWxwGrc9BItUhnmN6
1udgckvAqCjFoYL1lIZSRysKcmDKa3B0emTgKjKR0KlLO7DOt/1lg3VT5Yef9Ucz
nzjO+aibbSHzrTJeSvL3QPd3BUTtF2QfvEKyTZj8HAfMA205xiLK9kfJi8tQ2eFH
sLL26Bl/urRDCE5m3TSZId1WMcqDC6SVFwbONbrCJxIFF4fvtCLVD9CNiuJlryd5
TztwhBKSMSM3C87IDl/q8PWHF9SaXWGIGEgcAt/KpgsIJn7LQxazAQMFVcxm+L6i
iOkKgKeqJEQl9IYP48riEs/gaSY48naZya4sIXXBYbZ1kB51aCu+/ancHfMwu4LV
PpedIX7SR1d3QzGOHkZcyF5McAMW2SapnVZ++kgV6rrbyVhR4qTMouBy0RnVoIgk
NA0N0rRhnYn7DhwhXfxOPs0vpFHTs7kCKRim69CggwNHYN2i7ZM+iphKZkqKXluZ
nIQvdanYYmFZ0Qeer58Vf/pzb+c2Teqg/UMeTmpUqTVWqZGDaYoiuxbwvklQDAfT
+7QN7oDB+vkZtQfide2dCPQhbn0+/w+O2gO8Bw5cv0ErwMgTH4Vs/P80A3biOk4W
7YAljp+QLiMbMQf+X0lCTmQpE5h4WyAsQQE23/VTVE9FShdKyBfE2i00uh2rB9EG
OPGpzNtEJCwMbTZWZoOtPtra11G/iWKzL0k1jQZHhvb4CQ0sMNceIGeO7zv5TMRU
r+kfTzBZGUAIBJJPJf7Q4bCSusQilpxhn+Z6NxWCG2Fowt+TdyPVSJLULOAkPGmG
cUDJwqe6dyLwlzYDQdE9myx2+uKMBE9rNrAvcyLxNMfp6bFN/oEh6A/SsxTPHVIe
EdD6p50kOAqO5rf9SWrRZOOjssUOsf0JvjR0K/H2VlsEqMwkKqR/B3/rvNVCgTHm
d+H0v72N5KFgidNk43jHAjpOD9ZBO6G6G9BHKHu9mv/qnhRhAQyVgqFx7ZDBiElG
ahmkjvxrxSo8n2gm41qZCuJ2n/Oplk5ClQRm4eZDth2A/i4tZ6tWxHVPGbqNbfqX
71h+0cIXgkPBrmR8TIDcsEM/KmFYAP8GAAcAZUMYK4B+Qz51+CqNxGzHO2qISTy9
hwutwUmATomtM7zA+wJu3n30HcPHHYik3S8COLmnm/MA5nz5hWVeAJrmMc1gJjnD
NusNaoJ3VRFQ8W6fVM19vtl8XVCdIlU9kBGjYY+F/N/+SItryChAZC1TxSsY/cK6
Yj0KVSfoIVBJolXffE356gaKguUZAof+7SOO2CVU9LdEz9MUDDngXdBAiUR9t95h
HwVHEmDi+HcAqShUlRqtZRNbOqzDQXLUGUF3qjFdKSr0I0wy6ImVnPadL9h2SYB3
GCce58lK/XScKOLWr2rSOn4gQ3Q2R9bab/JFqScoHYqR0wv98yGuSxlV6i9amqun
JJbyCiS+0xPGF2tttaG4WdGji8/EjT03SMOSqu5Faq1bIcQ0lZecKhOirdl+1jZk
o419NuejD4paDUjakbeQ7Qq7braHhlgolkplAVsggT7vZKsOc9k1ruPAJP7zFlTO
6MbpLR9ZheUvoflvY6+CitBL/8a3DCw5goR0yWDpyOH3lAjXRHq9lfA65Yh85bLJ
FA0Wez9bbYFdSCc+41n4PZcMVWLbd/O/Bvztj/5ldQ5ABGWdHoEol8vKfgv3zTk1
lFbBmQ7B2CtEKzx/OCAzma6qWEqML/91tmjoBs8oRguTnq+CT8W6M7v4KOoafxzz
vb8f42QHAlDwQX0qrQ48m1l4Qi+Tt8qr+okEhKql+G5eeWVoRs69N6ZDqsgdm0Pl
9V69Ajpq9r6Xb340zmuASPv5qn5U74QI6BMSF/xKc+Ap+9I4D8DoZf39bqyx7UW2
iGen5QA8wbRULIWW1Nx7dJVbOchQO4vjPa5tvyMk2HmJmODrgQI0lahTbXZkKgr5
DZ7XWELhRWBoZB98LR82XKUtTbC8C0//hdRrvjLqHN6oAI2/nsMkNxBfs99UWfnf
NLnGMkYT8fjf/3Tnls4SFhwmdOY3b3Js0kQ4rHSkZFlWOC2oiQvhXgnppF73mzY4
m/YxXP4FlfHYekA47cmy/97YIuUjlTaxTGha1vbMcgLi7IrVfSITxOrvraRnwCvj
qW7E4pPhyqT/Y9y0Gi/TxEa8M2hEYEcWxlLVfwtLysR15qNkwt89UQdboiiM6hiz
PF+gi8fxPoGV0anfnXhoLpyZjAseggoh6xMXrlmBrIztl6wZxHDtc5iSdQ1J1ZVr
9idZlEHUucbNMOsunObxvW5v3ziStMInEuG/QSiGqVFss8HR1pulhri7alMkd/AN
CuyVH81OhuOyNGPeyWQfWG0QES7eOaEJYGtJYWdD5uQgivnMMEDyBK8BZQF8BdUF
PV7edVBkU+kC93IF9pZby1oaw3YwpgHwufHc7SSnESB3P4o5SCr6ve5bscfM+pqp
9pr7H6TarN5iR541Br1LZD1jBRulp21IhyGWmIEwQYPUoPdGh4+Cffnm2fc4cMT1
NazfqWRuiSjcvpFJyIM2t1Iykdbd6zC/ZNPzUdBTdr6EQSKD/oHxpfT1rcdycGy9
u+5SnqubA2PKu/RCbSxcXW2rzND8ScwkddeWmQPE76hH1pvvCmYsLLD+lfrRWiAZ
WFFGotnIXvu72PB4wWi9Nwc9ZW7Z+4Qi47fjhq5JLayTOAic9kpF1fkIZD3Kq6bQ
y/xg8ulol8nzsBcyCnEgiESQv1cbHIJSXQbx7/lty1FijQkGdz6r/vOi2tdHeY9J
IJz3wbkpJ3qUWqdOQiDl17gD4PyUAfw7aIDUIcIbBjmen/vtfOtjgatAfHZjI7yA
1j2mGoNrtaLt1FxqokY27YOI2ReWNfGudI/3zFR/NlnvZpBYKEAF+1PEmueWKHMj
wB8aIXd6jqqEDGODYRAahH2GQDmamP6QcEq43iTHn8sv0DksWoWgTbKFiwM+mVZF
kiu5KAgPBx4HJ032qzOqRVwIOxYkAHYpKgyvsQDPj2qERAE9a0olQKWiSO2T+SDe
DwnWekoHUHYZIxyzwMaCyE5E/LFB3OmYF4gqfO+O0nv2Q7GMzA6d4dG9CIu1Md8c
P/IoEdWAFMrACKVgp+u9b9ZHppwiO2NHXzW+3yhHTIdkbOueu7hG/RQfaCupcG2v
JbN8FHDxsTsf/3jBG5HE71k+8h4IzYEUTcFZfaKZbI1EgSorrsLD05zI+Z6RmZqK
oPxEfn+ly7VGQXG1pq0gjalNLXGRmV8WOpW1Re6jv/yMBc0OobvNuGrP9Jgf8/AR
CPcayxzASg+CyRvTodcZiofZ6SDx0h282LyNey+HFLl3uD0ql+JSOZnR1SO3TLhw
n7sFjCkfTPfOXWWiKyH1HHehSa3iq1zNY5tI1Sod8dEGyXoqlY6JrKYMetA1shHz
Pc54lQcMe00OOmfPqP7KQrWAiqc2nk8VHAA1vO1+dDjTY3xIIXqXDTABwWiBBkcj
fpVSjcFoaaRgWEanL+jfngLJT6Up4fCSBITmEu5nIjR/udyDWHUnloJpfWNtfbFJ
z4eJKUGwshwmq0MaA93KcJzEvYj27IbTM/wqIW4Z2mru2LEpU7AaETM8FObF5wJO
q1uNZikB1iIme5PXG1+3BTBrv1JApV621MboXb9xSh2sDz5UPept1ntrepdC1WtK
HZFC9/jLcTcra+iUUhZbfFSVg4u55+49fEEjMjfzfjqd7AEVr9XyhcMQl5KUNsw8
Kc3xp+s7eGLcfarDJf5Q7HUw2jSk3GdDnmcyXXkrHpIDuKk6uKD4Cz4kVnz8R/bp
v7wXWffCKDMeeheSKsOtp0IkTEazjqbqqhqEzENBIyQ1ki8kyxOQr0/px/DBnUH1
5wlSsq+dnhaHHSCu517r3PnwDPF6nX1WSTAFtM63luuM9tNOyNxGlWLNvf9rexzC
izAz5rplbCRm71H3tezp0CWjKt8gor4nrYJPbLgOJEBLY1KWVEb357BeanJHADQg
NLcEqBCpOOAWfqI0GQ2+NTmxjUZLt+poUbna7HUeW5zM99gBU285ZGOFKTV1bUgN
bBbBE4R9hAPQySZKnzjjU65HOcaXqctaq0y8jd10O4laKymR1QzrSCxJTJ+smXG7
s2teHIiee57GgF89WgF+6+WF+57Og1i6khU1SgXUYBZbXkwivaC4neFrMUs5IUfC
xfipRH1FcnKbzVeGvOujruPX3R0j59/WGbFtzzRYKG3aE9B3u+JYijiQaRr/4ur7
3xdQUk2xoZJljsTtK1KCYgfxJMPT+WWeB6gP2Rwb6deT2FyZa0FJqcFvwmZFEZkx
GzymsSOrHlh26qzKWjhP/k5/pbdV7d6WWfE2Mv1DrXGCsopo34CCwPyqodXO8lwv
90fVE++2gsRemmbJ1AZQCxgZL9yvUmZaklfnuSUzcX6YZmeKRv9vOB77NoUuYnWs
qhjn8LiB+VyhOjJwAWi3EfTY7XbQ/nEVZhiqbz/lLQsOf3LYhD35Jz0WviHDXLwJ
BC+zvXLagImH/cs13RQzhvxKLyTjB7Sw1DRWjsobDCP5OQTfoEpOSCxLqQhWkIWL
p7XnoPC0XJfTeeFNr7RIPy4Xp/FWsISRPo83/eoUge68vGzKN8ercbUKDYSenIQ8
nA4yLz5Gx/QBGMToeECil34skGyToYhUoZ+Vqoxqn5tskdVgVu8JfvrhypDJlNV7
2KZs+Jlbx53ZjVbCoLtlR5OmEI7KEJsym9t1+KuSSyIi9nvg2IZk1wQGXNkfvrU+
d+tc1aqF+05VGu4FLT1IdmuNzTessXT4DsX9D1BAZZ0EZNYXk5lBxqU1XE9jPshR
4IOHguOtRH2NC2LtY92Wo35JjW5XeR3KIcd6O0N7fppUdojuATtO9s32QRkFu6Se
RSCzS05asgurhJb8ImWHfdFJyhQZ2VsB9oU/C/4jpDOs3ffJvtKtfRO2msqISnaE
yNnV5Dw7YOPdwNFbN6VVHC6CY5JBs8VP2UrhnLaPc78uqpm37Ne6wB+giuZ3R21J
hHW149tqa1cCJsFCZHtTcYjT53LcHx6B+Iv5nwSIQzzNqOoUv+W27NbLWsrcbD+R
rrrahcHE7KqIXHTbPGClf8E9uGIgLpo4Mn9Y0wCoVNKTDWWgrHqbGA1hbwUaXw3z
efji0ouuFlnzLbxW+nbmcddKtE54N6PcgrIUW11X+dB6/qeF+6Ws37Ifwi+2eSwu
pqNFg8UdaLXO+cYkC7za5B0AmQ354LI9sHtIe5cvBzNrks4LRGuI1oEXT+WvyOJH
eyhPw8oksA+GEJxg3nAIufukvS+PWAu6L1hl4BMPZmNbGERkU6O8lU9mNCxl/E0w
2KaHHwEHIuCfQ82UwOCxbQpzHOeBMOWuV2y8z4If5BhixM8O4mWtTBBRw9tThyox
vA9WUOJbLaaRxdgQyfHlg6+B6h8vVQUAYfSSMyEO9BXkI7gJL9U3jblVZk6Fuy70
k/3QxOMpV5zgFzC2HmJEKWSrpUeTSCZ14IzyXrIFiu4tp614so4c18QzFO4MKTBz
j/tYNUdBkm5MlYRRmwmmKP9RyVwuDUncvXozdt6tj86Mjjf0e6ps3qV/OGXUGKC/
CnQh3X/nnEgySaTTWVCitSEQBAFO1jo8zdDfew54jG7L0neFNi91pQxyOwVYYkAE
ZH6iG1rJ8HiT6mWLapi2uSc2Mo1Epevp2P7570Z9f8rl4LU65oVr1vBBvEoaDasz
xplntrWAb1mCW7o/VfQbjnsRoVjiM+6Sd7u+TtswSxojIdoR8ZtlQwTgDAxPDqd3
G+4VSchVDtvkgAOD7xuM6jbfXZ2QH/nOcTKLaVPfxq3Hm689nd4MOqWGnDilfKVa
MFK6u1epubIQCydK/5CPySBPCWNinPfXAeNDPEnPP5TCJskjx+gGu9+qRwiuWyA0
hip0+KW5eMNXSnwwsLeyjearM7OKB2K2c9MiVlakIbBrNfTsPxiaM/OiqphywjSl
AbW9ZBrFIulda0daB/XNpcIAcu3IruyoXLJWX2YcfYlexBp6x2TijhK2ryR1elV6
wFSBSTqDseCL14xpxJVg2OQpF48ukaTcuoBdmy4+VjW6O9PX/Owz9aEV0N7Dllaa
yS6FVkJmj9yOzX+KNCNP82lHtnKtn7ZWpZn4M7kttmr+Zs5FHmpO4KIjRFW5bFRL
ev9GRtI9pAYoiXths4sYnHHtlRN4LSQWDdEyd1dVHPY0iI/v70jYAplTgKdIMPdy
tmljEJH3Fjd0snSL0PMrB/DpmHWgM84a4MLqdV95y+qGUCIBXZFu9Q4yIvVr6gxX
xRe6Fe4/1Liy3jjLHQybTORshMwyLfTrb1XgF8nhcSa2yYIH7gGTsrzNxC8xMy+C
tETJoTKs4Bly0rzb7GEhT3h81tTOSYUckpBcOpW6+pfYpZIXDjDzz3lNw2ALJ4ki
Vpolh0RZJVOube3xWC4FlhwxnS36lsRJt0Ume6q6QsQ+fXmUoEuHPq3ZKYldTze7
NlgePaZIV34IYJOxwuD6tSQIxNn2eZ9Slyc+0VO3BAPI50jVP/7ha4XPEYUutytZ
Hvxy6+ZRTS6RUlJgbNu84B8eyswVwW+5/vbU1FmYMJHL7IGuQfDM6jnoJcubts4Q
5QRIuNuiHYXzWGHtkKUaQ7D26Hy+cffAo49xHKixAYNmJnPQYVDz7X0ZaOiOBIgh
zxUXi6EPZM8UQfVBkJt6HvtklNqIAwlcFXgqG4+5AQdya3arLOr+PAEZMlCSyMNx
4KVFCeO4S0cpbCXh71hP9vahH4AJs508HvdJ154CG8ljoj9N7iKQGxRDb3K/+iJK
kdtrUj6PsTm/kMPri3VsUCA1qZSHr34P3z1aoWrg8DqYKVymQo+CCUuf1DPXpo9N
S8bF+Z1k+CTfCg95GBHPli3jFFQf5tZGs9SRiauny3WIOOcKMFgpM44tqprTvIt7
cSPPBJOZ1subiFPvw9t5ebQolcGxS30t7DcueA17lzXt5X4cz2wtQOFKH+t/ybm0
BUZbQrup6vSzKq3gMHY2r0cT9U24CZmm5EVpYKegvT6Aga4oyPjKB+g2oj9P8Ybl
vU8EiKYtFBBlcTg4MVXC3R0FLP2GMZZt25iJyJZ90hPHMYoyEmBeAFOCjFtpLTek
kqR6582UDjAM25xRMuxg18zg5yfMn+s1Mafi2DRXVzcBsK3iDRs0zo3hFfv88iyo
0XYZNbCc85jq/HrJLEM0Opg+FC9eB6oDM68U3/k0Ro9Ehf6fvEu/fFvpiWZQSSMX
Vn86cQWo1odCj3EwUXR+OJRp/ioGDUT8U17TMYetkIZ5BDJYpVnfdDtWApvVWYP/
+U//v7RKQqUAtBgP8RzC40d/5irSzKqrOzlqbBBNNNsQirp0szP8Q1YJcLFqQ+eJ
ISI94IOLhvi5rBRdj4DcZhbxv24E9/s8v08agohs/TsBhEb54Pc78oPNUGRZgVzP
36zGLOsS0F+ECDCVD/3VgJ9CVBxYGPujEzi1QB/dnCe+9ZYlraB130nGgSeF/sGR
p0Q849ZQ16T84alWuwZ8QkHpCt3ekFLkHyCnqhzKotZD9poeUzY5OisiW0RLBYx4
u2LMB1jrsti5JwbwcAuJQRBbmvzmG3pS8A16s5G1iJokHG4CxzfhbAFxknnJm7cS
3ATBEXlRNrK68tjnRklSqD3pXgibbKdgB+/cZx650CImHXnOSCIt5KfWhDxa4Cr0
06yx5gYdnVKKUMB54/IjICUx0a5Kfs+HyY7ZSRYGvQu17mCbxf40b1kipIpR1gJR
0axgCgv6Nx/0vtE6xhpRivJpdFcG1Q1nsKm9h6CPnvLdYcJ+w+wDXktYtQFK+v0J
826IebSvvN1KR4Lu+dkm4N3F78LfaNnYZfnJYJaX2yTOtd2crsHjiOerDOo1oSmh
vXm7B3Uc7DFMwojiBtvilyGktejNAVMzMjhOVwXFxIaeqSQ2NaoLKUoBc9PB2jCZ
PpTm5ISDX4TpcAcIue9edcPuq3rgsD4Vt+w/UXABknChaR8imjsI6dNRdiPHtohj
DXBxfUjP7W7GZTOJmFwCY5vE2wc04BD57mGR72oOaPtXPg7L5Q7JnOT31EHaLE7H
VBY8KJg62mmv2zZEs0F823D04TN6kNts5VptAxsVwWG3pMmUz6ET3Y4W6QgRUgWQ
Fj2axtKlMirLZeI68u5wwjXYpm0Fj/ld00IdmVOrEypFT0pgt6l8IjempfmtJYyk
xI2OI2nbco8B4mhJKH0ClGRCLursmoseqc3wjR7Zq/VJ0freTYUBDSNdoInBOCFm
gwBT63OY/rlg6ZeEjDnMZouWqd1l2lnzLasjr+aLIOkqqc7RmaFl7IDbXVq/TI6S
WjAhGTS5oPVuoxwa0W1IJRhuYYJDnflTGlMPYLk0ixXFtpNuvAbEwg+Z+VVugQC9
oCkBbLlQl1FwY8afPuX8fSCClFLd+uolPGFN5iRogW35P2I4SFN7ZcXKG0rIsc/1
CDIQG9UqMcvG7APT3o11FFkvI+PwqpR4N0xnQAZBo8KBGubGoEuos1yX+82aMEmW
K0dNvyF2xU/oKLhp+zYvPDX/A+meLX+cAUuiytGc64WXmfjmCeUJ2Ha1vHLyRG5f
/1hF3odBVlRvkM84FBmhaYp7j0ax7ZSzHA56VTnAhQZsYp2wsGoPvcR+Vpeg4dP4
ma9k8cb+kqHQmq480Ms7vgGK/zoWKbV9x8b7c1kZVX8rHqUwUjmrLyO3/LFaQfak
gansxEApE77tQSdLQ3yPMjazPXLbw3FiVzWuXgOWsvvyFvRBfHRDHyzX+b0wxe/y
13AEjKax32tEuAhka0/lGb7lItALpEIIHU18pE1lA1qWRJjOvD/kGbhhKTJP1Ilc
Yxi+ltwzcycQiMAmSpwoICJLeyfZqqgH7ISvnkShVOODm/pZFIAbYqNBPeckX+jJ
HdeKUTnt6NXxPs4XcI6FgcxEGHjJdMOH/rtxQIw3rvwKg0NzSjxFSXEIZ7g5YYtC
EzObcdmGg9tuLZC3pziYAvKadK9J2dR32MMSi0Fb+xF2MV4JpeW7fhTvyzBzrCPw
B7eyPc+L3C/ZoNklRojjU9p/lY1uN5yAQZe6O2I0lYpN7XX0K2kD/VbPSbM6yBnK
5RYbzNVyi1kjFo5B+Ej7w5vKzEq9rUB2L/qZ9JXlmm1f5xVm/W/nAtzJUA+pwmTL
QH1bO5ob2H8H/nHr96ErLZO0OuduLxYvSymYZz6dxGvcgazUcfLRcYaCiMcwdz1U
Q/E2g9STQv762Xw9sL0wCRO/MH5puTc4WKnzprecImXySV8Q4a22h4wQykr0g3tv
iYQvDMNBVUDJTOCwPF0ySY2pJ2D3D/008NJUqzaEcnvzJtocYDgP2bEqnrZmyMs9
5V5JYh8Mnv27M8Qp9FokZhp4K2MeFYeSGf6JD8+5k2W/T7c7mO3S3pn/HrahYn1k
K0oYLeIaZSvgOaWoRab9gUINWMglwtcKjqx1htCxLx4x1tPV/W4kGosBn1JhVl8d
fn7hKBhp5XNgXWto9zYGPqi48OC0yE9yscPN9QUAMrCHcUR1ecMrxrsn88NEFL8H
a2QFcmMtH8XmyCSfg6J1/8vxsjqT11oeiO6IudXq4xmR/sfbCs1FmPDgx8YaCVSe
W0N52uRRymVXW/HfPt5WKkQ0nxZspPSmiGu/GahpOPlqzRYGGc497NFyFOVbZB+D
llQ2/7Xy45qU8HIzMp9sL1+e7xRnui2QDKOzRF2W03/LhEEqK7WBILYLD+WFL3m+
IB8YgQQ78Tzkwf9u9SiVcSkXFB3rScCJw3hDvMvRIwgHys2syqfFq0dexFB5Lr5j
v0OAhxkoe5UdThKiP/X6pHjf+aO/18bN+AYB+kOoWbCs7VX+6Er2fBYaZhIRWLIg
Xe20WA36+N225UIpRyaROBE9cyeqqhcG6Ld4mgBk0V4DDO6zT+uPveTkW/6jVpc6
PLVSrnZERoFh+7AH+vLdy5icTc1kTB1vnq6/us8m+bdsXyINQD/Frjx35YpCU9xG
YkCkcoqb7VCgwxc6Pc1gw3OzuPvDY43jvWA2audlHKEtguVWmApyaOJ9oGkTU8ap
20ex8UqbP/l7qKWK5t0fSr+YvLghcOTwo1D6KaDojhxlJ06hzvR2m9mniQ4Ce40e
sheUoD6fHeC04T3qEFpeJoh3IYJISvp3VQ5/NCNXqZTqO9cHg6hnAiNMlIbyDW5t
nG4JUbdM/c1qm9Ae5ppZkEY1iKEK+25x/5NW9wzlfTcT8ammv/yGc8UJ0LZ3kSn5
pesUeTb1gUepr80Q21wePMEws6INBaiCCiIuB6yG35cyc6fvvdDTbiLrmUo0+PAZ
g31mQocjPqL/vxP5ZWy5NcO6/kn8esvB7mgyMC5bV6/8GkXbCUxJ2VpJuskHtnyS
WYSz+EAd87uYuDS33hCL9H3UQROUdYzYjLHy6eMHC68h7MicNdS8Zk7nyEpIKp7y
D/vSt7I0NpP6y08TvT2YE0QRMl5R4ytOiPEcrg3rcgafEJUPc/jnZp6PuKwwQM16
BmX1TOXhluKTGh7ZTh0to2iKoS5ScMrpVjQtagkLSwP8U09V27Fbw3DeCr8X48D9
MWQL04x3UZUXor0yEsVy7oEp4JmU+V1Km9klNdEV+Ih3QigXPcNZP5tA5yg7NzU/
ZezFKm14B63baVsRwG/ZXAJcnLQeHxFdv+gzvL1TkJAQAS6GREwqTD5ijr9Ckl7E
+KQFdqTowElSq7pwQrTvGarTnOi29z3f0AtQz9gmE4ksptvwqSztCuWbg4r57y/f
FRcO6DO/+q//CG2rRt7Jdu65lcb7HfxCEEI5pl9pYJ+o5MIeNEsOihA7IEQN4TNd
+PcJMbjQbx1G1VsX3BGWnghI4jfvOjFPYt2dZgcjyBz6V8yEMA1FdO6MECfE/Rfg
L1vjvP44wABO3ZIg1tHfCOJjv9TkftQX5BX9iKTK+ipHHn5VVosGnW7an+sZp9Sm
g4B60mY6Rh9nZMVakwW/2miLDnYGJyLMfD8ZqR7U7QI7Uk4E+cFAfQcaGdwpHOru
ZAu52EGNDo9D31hjsiwsPWx7IxDOd7PiUGJJeKzUozEEP3ptMVUHbTBzHeIgu9vg
scyLfPCGl7uY2o016OXE3swjxAQGarkvbU8QZJt/qjbC1OorrhN/NvxqaOFbCMTI
ipc6XqnbhzC+h6LSr0R6kjdlhD3E5lj5dKLrVyn5sM0sNq6DkZqGR27SUORZV+hs
a0QJeB+S4kWmIUXLaUWXxIL38kLD56pYW/t6do3BHTqpfAOXRQZ7/J2rx1Sf4Gxt
GnnCC7qmvM+CYQjAqZmSWyfmEobon6weMVdNluDL5CPVqqvA+dEKn29cQ32GZk25
yr1hrDaFUC6ISC100wpqgftreBfeqximnEPvJlYoqOgMlNOTQTdxKmlX0GdxCzcV
s3aq8ilGh95d2kVnRG2Jyt+mQ+mRLx/bblvF2FF+kCAN9og2eeEfiZ4VVqB1fwOE
Y7YEq921cTHrt+56p4L14ztUoBrdpnOIOU/fz+V8/K2mjhjYtmuLqrSkfpHQnSIG
16IqwJykgStMU+I5vIQ4d5sC83RKfWg25n7/GWQSA5m0k1ieDyWSxvNC1xdV/DsX
qTUa4a3mtyfe1zeVy3UxSkgBf26PgLDGW/OLsG5Ick0aMBn7Dw6I/DI8YfUxL4Uj
0E7uiYNqMB6CIeO2Sgu5E16sC6+Jt1shohZkyaNDM6Yw/V8ZG4uScVK1nJ/nuWIg
KDzo3s/K/EzWwttNMjNm6PJGT24FHrAY5RUm0S4pLiNzpfJtKc4UusY8OAKhyBrf
bfnVAhgdHgFZ7WilSHJyAG1jz471sqmSprZA9xmlgn184IxCj8/YRcxAJmebZjVO
TM3WshCSapnuHju80beKUszfnVFkcQue2eOUAtus9c8QXUMhuhK4ssI+/wV1KtFs
zDi2Zb43wYJ+TiDzNT7GUEPmJWoRdKoLcajuuLsEjMrly4bgICI3om5x/RCTpJhv
eDAklukOX+xi+h8cj+tHk9oBHCvwu64XvcKpQube3U7wpG5CunzKHuWXwNPACGvh
2s/vj+1ExAOsJlOZG7JahhYgI3FS7ftHIr5vrM3N/xD1q7j49CYBUz0RXqLP1RLd
O+0t0fhtZ3KNQ2U/OsBXJ/rkdN9242LNpQRQpn64/q8078LjSkS3fri11+/RMGWO
8cGqCPYQ/UdZz3yy8Wn8eB0J2RGbuhCSd1KvZIyAYS4z0Soy9c2ZTfp2yen+LUHj
cfyzwqmL9tFEo1yMpGuMIDc3m0/kuONzijn0uUvczgXjXGzvVzVrWo0hmOX1tWGD
z+JMTmDccdq12dm21xn/5MwI+dnVznD9bIs+tdSNgWSmhONz8BrWpXfIjk5HRYp9
IAV3sbqc8koym9wqYp2LjN1WgS3bc4GYsA4YWNTHC1YblDs5V1EE3p9VPh1LUrCS
Zs9xeo8Rcl41RsfwqeiXCxfzTYrZs6b6/s0kex83PVoFloaC2Imw88eMv4LUqhr2
EBEFSqKBM5GO/QdpNKomr/YeboMKicuAbHyPKz8UBAIm9nH5ydb31j+RMxMQAxii
vpWrFecQWe2X91W4HKBa4egTBb5Tk4ASMf0KvNiR5nGe/kELG13W38Kznyg/U3IK
OFcRsKBanj3uLmcGGi18i46dz16m9LQFqKwLWiyZg1N5oyeme2g34TXttCW5Szf6
TQ593fKT9mCTkBscj3zXnLgNkF5kzgpYbIEY/ZCI0xDRxUXN/jweIDLlxOebRHOE
GjTBa9Jep2PQdRxJInUFW2CPn32uNf39AuZBi6tNx9V1XUf24CLAyxLhYnAM6Vaj
Q6xPgoVIUBxjCpmlJnTHqMXc9TebB6vf5R9ElPTNm3/b3T71GITxg7uvYzY0Bd1j
geESFN+qzfy0m3AhjVvTxH+IB4g+unRnxOCJJQ6pubDWBjKpARghaYB4CgQd8ZHr
CpqRqzWwx8e+YFZUaEpZUbjDGYHfWMut7BS170dVXB8USP8jVnRUm9yweCdaakWH
UVPYAaPr98ptuI2jop/vmwgbGyRQPNCUl8PdX867bPfbPYTIDGfBiRiqqEpkabGG
406pw7NbnXIqDAwIht44FtofYVzrv4eXrhmWpGQMdPErW6xmPM9VXfPlEIchIQ7G
YPllm7Czoojru7AZXCrNvltue1/vyMJpRcwJhTkxC0C9odfk3qVqWBQdatcr8MeO
CkeOQZYyWzbuGUwZcYoJte+kSZoaqayWVR9TOIBTGnWqJegdmhh3N7nw5yjnzf3j
dN6fZhGa2NCJB0U/ugIx+eQKqTROKxy9CCANc8iOAuHcjDJYq5QchSqTQzLNLXGW
OncW+Survp+1Q36EcIEfGXGa7emuLgHv0q/ORHEuspc/oCUHSeVWFgRt2mJYgkp6
/JDJvjyFUfzoJ5ag2DRtKGf+LsLqEePigMZR8y2ZGkSuOtrg+OFlM0vkDJVPoLFZ
L/PGPANTLb0CfE+g5xybeMIvvjzCH5utAizlA0LRnaz5SzOlLEpTzodh3gcqH2N9
N/RGtJG7vcg4L+pTxfzI2YLdMgaVmiY+nphOHgSdcgJe1fMKvElM8IhbD0X1i6Li
U4awsrGkl4eXZ+GA0+/4osHttPVkRZ9GnZD8KjIe1RkYK/LNXFsTbcOtKvQzyo+J
TRrW49xApkHnlum2RRQJp4e4f6QB7vK+OoInvVGscVK+e6PbRqMiAeuvqrq0ZRZo
mGIZuZJxDX8OEtopaMavJrcvI4TYtX3/Jgq43LP6NL/xHwHwQEFyKUnM44SAN9nJ
gHB1JrOuyzMVVN7QfTpw7qyShDn/GFwmppVV2Oa3qjgBcWKwHjxsyhJORiy+7Xir
i3UbS0h2gyJGY2OwS4IhE6UBE6vGq6FaiYxVzC14+Hj/fqeqTQK1/skT7kIkqaqH
Z37x9RU9yPwgo72nNSQTR/YRATrrPKhweFjzTNQ24YEsSYF13RL0oSdYDkcl5Qbj
V5UcDRKZAicKO+1ybAa00v6O7sAZ6ETxkr8JL4m1tpJUzUb7vxzFjVPAydSN/RX9
5/C1tRp90PLj6ljMDg4WYMsbjrW64Z2aa5z4QmPIwXp5ZlKA850FJpg1zoLW+TDn
JFAIG599YJSNgEnPPm74qeCCm5CgF+rj1Y276hLI3PEqoDbsft6I00meqB5X786H
Obnxw85wmY/EJI/ZFWEDZK8UvwfMwu8e20wNFcZmfYEjt6AzWoDNlT9/+DB+GafD
90BEEI9IOUBG5Nuz5meTJqfnaFBkobV1fhrJjZtleCGZUun5OLRfugU/Mgx6L0U6
YzVTiCaq4bC80DVY7VSwyUIyoQbCo993FI1lnfx8PatM9cIbbYZd9CG64EypHOdY
9XUL/GRJmcu4rlnqsrg6HelQwYCDYnFQ7aVyIK+62bB18cXYmacdh3dXSZA1rlQ/
Srolx/h3vjwybRUJ6m3S+VSihGpQ+h+Y5v8/HSuv2tfeaGcDp/pE6zS4xNNLfVmF
IoApVKncfKNXxKFt8R8pQ7rCqC3u1qyg5nnodkl5IsawQksOcuoXnypbO7cKl6+U
+b38xTa+EZjxotgDhTe4malLI8wz7kTbLu5IL0enluAGkzGM1IuwnlzETrZiYgsy
Qbu/rd6Zvm8bqREBmjL7mJ0iBMvXcS9NyyTdb4V8nH7xQLyJO4e/TAS/klRQ/7yH
h5mwOcit6lmUYTkqDcfMrLN8uwXSVrlARgKQ+nwygha0tDxPmBsCSRaifzB+jTCD
BxVjugdKg4QzpnFfEOCjDN75qFwNtmsJ16LokdBeSN7dyQBCNI1YcbLRc7bpHfxs
uvw5+0HzUtvU9ZC4nMTzAz8FymLgCfCRNyww+9WpsCZcv7ueGjQJxpf5jvvuCo5K
X8kGiX0rF+E2jN5cwEXKbemdx5x82GLeqFyPtEMLcaRgy1wXGgxloSUReAVO5IXk
qC4GsaKlp5xb5ScSC6sbk0lj4ie4R0iP/ce8aTcRIicC6mzzmCa49I24CrEalsZJ
XrNYNxCQ9hR0y5+droj7RwwUfnNJSAD3zWxIuZf/ut4CDHGeAX/tVdoXr+bqsgtU
DsbEA74UYmtCRCnlUujdILP05+91DPuGMwa6K6OeqAyKuyXWOHq2t9mz5baxLG/E
I3n3q8Cz98a91OMUMvN7Gixvkeu0khgrZqLyhkbR8P0J0AvmJHvhlZJdGZV2C9uJ
XOFhoA44l6arHvReWHo3hhNLSwXlkAin+Qfodzb7LIWjWGheyWFZl2s/6Xxnj/tR
kJ+rsuvrpJl05im8y+HoLFpKUMuvFimAvz9rCqMeslQTRFyGO5Pxrlg7/ICmBOUZ
5ZGBaomoVY2XdYUwogaEBc1k1JGf3MSVQfQJ4hH7/2KyymdCSKEl/fy+VDpFcFwb
+1P/5ESyTk1eMtuVS0LPFmdLwJfuJ9bk4tj7guT8e+GV1da4AsrnFEAY4su53fUc
JnB95Hhw4FW+8WE5S+z7EppozCzUbsCXl6KUDeb8wNQbZhF2Pwe5lAZhCeq97W0V
ZpkbX3PdIcfIjVnOaSlLxtHzVawKPnGETQ+z5hqWzeUliUHjbxTAdOy5zuNv/gI0
1I1FIdkAiFDDe8VsmmO/+LeadC2b6q3BMTE86upotJauu4StsmSwzJZiIUAG+QNW
EDv2sbaxem7ElQb39zg8ER48CR7B22wy4mygFO97QvDaj43SXjXIPd8t4TYtLgGb
K1uNbjFWIHIOxC+qa4lLInk7597CWcrNiG/mLTmAXCVl2p17BWCGXkY3kKxNBO4U
SsTn1SW43Hbusxl1D2zhP8378hynjTHEHxTZ5ky07/vxXbxzMbqzP/wXx3x4fiEo
Ig4DPysTyeLhwgbVJW4KGEfE67+dK/Uqc+gPj8r+1g9MjCq3CG9DYMddd6MMGxx0
D14F6xh4sk1wzRV2OO3EuhHjwhDvMZD2j0F6STPk9j3MI6xf9nFom/c/3GoHARgf
FAp1Na4C1YbHuCxp0GfQzdrG4hggDmbrx76x34ViXNejXZIvXTL5NPx+9a3Yii/X
Dv1W6MDAa5EmUgFU/fC1B4Tt4TQyREFX6e0IYLWP+z1btVP/6hpx/8b/89lo/uNg
UrM22/tCfyAGh0XWr+KjBjl8oQstU0ksclq2+VXjlyO3CEqq+NByXDNj1yfDT0i5
0kxMPabwjD4m/X5lRF38A/cn6kZ1z5Mq/5POcLv+LcLNJ3r5xkhc7TjYpj2Ke5/m
JXCEbdscN3Bh83S/ptu+lqgwdodT10llKYXeDzwuaYlThzxHW6h6Tz4ItLzJAh8J
MBaexNorY4Y/WqZy3g4S3EM/ot5QprH7OQ0y/sBVzjr0Q9EizIVn1BYV6Dv2aJwg
yWTm7bSiH4BooAkzlSxCnFZ9JtbHhF5qw3N8fYiSvOcflK2u8ZTg6fdcIJz0IOqs
jm8ETVu4fzHNWFhyDI2Pp3Oji5pA1kcSv9wUmFGnUGA6TDKRoyHXiQ1y+C+CRaDQ
iGY8MOenyX5Mko9AocK58qWM89uYU6H6dKT7a32eBPa8sMe4dvigAE7lxGWXp7uV
0/JKbLOHwNHrTGXn1fIaqEP4+KeUTB5vaH7n9Q32CvKOv+vuoRq/7xureWiYom7b
7Bs9VjgbDMf7oiLJ7NZXAxJtuDZYFcGMG9e5frMYIw2Z6rh+qhdy+8jlUZMwbCGd
njfOmiIt975RIBrE2ClTRAu5+8Jxq/ell6CWwTItiGs/ubsvMEj/I9WpSenwjKuV
f6jeKH/7ud3QHO8WwljzNzbdKcufXFIVAC+JRjg7roKyQ1JgamLUdl2oDCG/zm7k
+QH58er4vMVHdP+zS0PWvBt59v2BNsCyKs76yWvuZix+SRgtZPkWCVbuftKxwI4u
UtMyUEHB9t2oPOIwiio6vcgcUB1dSj/ikoNevTDCcsIz9pRroOAC96Wx0wTg1tQl
aXRZUPPkttA/l3o95AHnbn02j39C5UtG7exfamSr/ZwxTc4aLPTV3BHsNILDq6KE
1rbLjSJKea09RZFiOBj8oPJfU0wC0gq4fnZAHSS7o3jvgTwv1TJke/SZ0+KH6LDh
koJBJr0N0W7twWK/vkl2GvmNPg1/12AgFeQRWKPQXmyb4v7kfv6dRpPAXe22DEG4
p8q8FKH2sKoSv/gyjjeuepRX8XHnZ0CHXaE3ouELlTOVGrCwL1n6GqEarxGbjaqT
mQTV7agwqE15jKr86CC1zB92jJz721VbDh/7LnrFWtVq0x/zQI8UK+CIZbPl0kEz
loecIoyAJ2twJJCcAOv0n0E+lWgGFYc4lUjuAjqEiT5uoLA1kLNwElG7E2vrgKo9
RNIUd6gl2hp8hG0SerjIEZcRwEP+Rl8gx+ZqukzpnVfPsyul2uKJ1P9TYncC7Ugw
b4w6e1KbbnrNxpNK9Pf/A9kP6zAbQEz6QS76gw3XGmrRdrwlV9nTyuqupzFYBy48
EEE0wAWKE14Oerl4lwKMaUkzArlK2YI1JBM0MWQZvlMb4BkFroUYYMAnwwXQrWQf
DEeTd8UjwH/RgPeOFDEn2RCzHxUOrgtssqjxQz5lk+zxHgr50t+OBhTMpImHLhyM
awOZIOvw+UyZSTvLwqYDhUPOc28xnlCzFi5NN16wUYYu1+xjhfxF1HDFwE1jGrOY
yThjh+7W8YmMaJz0iNbFifnaciciwIJVOwPaaY0NmmHxGR3jgh/Kj1kf7yYVtnwY
TzgpGt5A3JXO+5vJynLtlNcFJdD+dLqfXO9BN1gKcsm0ocrmlnwsgHNhZVl8wj0r
3cDsCeQ7holj2iyr7W+vR7cBDbW03rLPz9pMGtez5AnswaQXnO2xn0DKcFK+yD62
xmm73JrkiDsULku+bAGTDF9B2dXAnQfAfSt54zZOwFi6ysDimCLu0ligu0q0OJZW
D7p+o7QjXXd83AyjpgD90pVsMbzfX8IANwQs6L1brfHgmELpsRcZgnkk0bSpj31v
oy+abJfDPuFkvmp2ND2e3mkYOT5ayC/FAZONuSy/gCpVx7850I4FzuTsVyJfc4h+
DC23mE8O7vaQtDW4B7Xt1NG0NmSkkWsif1+6C2vQwr2bxq4dbvicFOijoU8/LNPp
M+/pJNed0smq86jQG2HhPhSYsU38ptLg6Hn9PcnfHHWVQxcJtvIa0wvXyat0MnMV
kbsA3gnUrUcxK9m6LDoPV/Ln/NANYRtanx1tEVuz6GZuvj0dzsC1zY1hEUC2WHNF
VPnjpCIi8o8lo7+hv515X2e4THnz0a5LQJs9xZbumax5BJQ6VgG1Tr2AlzEnBt0S
2wHPNR79O39ek+ld2Q4aePrdMMRI2EE6aXOJVZUHBQn4sE3SkG5hUmIEAxC5c8bG
kL1shyaWfWNpmYiil9uBq03FyrJjmuexoym5eEeyRMd9Ydxm96wP7tMmW5195872
QNgFZk1zCqbBXhyomHdIy/zfBkdsmFtwIEAXDPg0tSYfZwlp9g7xsREVh7Ty7gBv
N4ilmMWXb3I7Zz4GZFUBXeSZlJ2DxCHEehzjvvSfy3kntBFiVLKsjncW929PYmR2
tLBXCCCd56ZXVQWRdr5EdM8Pi8mYQybk2ii3XNHmx/YsHM/RIphn4Llaqi28eaPm
J31WznjH0glgK205yFe4yoK66z9v2JVzQkV6A4lwyi+UZUjlokmUExKAL6GrjDIV
Rgldtas/OCgi7MoKQgmP5D5rcOO/0l35wOeTX6D7d3vWXR5jExqFlffY4MG0seVs
LO35BXp7gb7UUMF70tJL+I3zx7fBltndTc6EkBuS6iB72+G+6/F206MJ9FR5tFYd
p+fPOR93TvwrgAaI2oMkykSr+OonIsZ3demtvNliXbCxeunelyGcvG4qD/oyNEw8
4yh5j0iJxoXSJm05w2W3eatrSzb/NTWRaSFIKGXjnQpFQIvcUmlBgsKBezmpzNk2
M3XcHvchptQ7SdwPj2bBkYAkhYL71lAcx3CYqwA++VjQiu6LbeYsZ+Ts1dNVWPMq
RsumOdDcJStbbCY2DhpcnZUA2g8J/r5A+lwnRCa9lSGHu5Srx09CujNOOC92kqCu
u856bFmScnM6WGSKx1iHsLm0GlqxYggdEcmJ65oqaSmL1n1bNePkeGvByMF7psoT
3foIDlgR272WQlpeAFxdDO0NINTc1YQbiDxr/Z8dTEUvHom60lOH+n6F0Xg6RuGK
5LB9pBoKADpXdqVYixKM+1zSR6irEYBctLuxBJqS+CPXEPkRvKWhRFj7rHB6Gy64
KiUKOYC1kZ/eWMWu0iSeMvBeUM0beZBq84c741xJlHNxC+N4t7h/qljoy8LOAr21
w6Bf8EpIa/qchh/crpKhSllCdxwVoqY5MXOI++gRbXgs/g70QZJel5H/P9eZ1Lvz
Se9SVs3duoO+kxWdi98sHa1R7Bg5aLX+eVRYu5onF8QntqoY7GcmYG6JLoQ9o7/1
9luNFUh/UGtleWLPaKNGc3HI/4Ai7Id6/l4DL0g+rHVxdU29jZEPDy1w4W1t3fZ8
SxcUtEPVAHYj9IxaweKp2/0kReEOIY26nMQo+oz/fY/oaBpNTxnV08N5gVPnVIT0
96qcGZb9A3kb6sLzU55QW5lQwMUVYDpccSFxpoFntQqOywYixdO3lETvvpkqmyYA
QU2XvuQmSXg1iaxuT1N99a9HQE8863W69Zitt0OlFISKFTTF7+WznW7CjH6KaWnl
5rM7aUgOyqjHU0Gfevs/kM1ZMIlMO5nhdv92Od2ToZy+LUTFhSwU+CSjx8PG7tgp
hJYWiUDYe36pfWdL5gpAmG8Tvx30DkiWoSZ405bTvc1uytsLs4dBq3IlS4O1EV9T
qzUGElCpRon3ZTo7XYHG4U3KEy8Z6aVt4lrmZ0lePNRsGDquC411Qiw0enxk4wRd
KpGJWfidhIjM7JbjerHYmqZTw9rc8xRETHYhFOu9Muho97whUb4SXleBPq+C4E+V
YksUPWsnYthczNzquO16WcDF+D11J0GJxg9p8vxHq6AvuZAsvcWkJEy9SQHedq/7
VTjTnICZTA9lH35LitjUcNX4hVvzs+1u6d6ag8pQwQ/51RwGnLmORYUMO2fTThgZ
JTLSkxVO4IYVrgBsXR1bihC8F/yKDi2e7Y+ZbBHjW6vqhnau8Ba/QYWXxUKxgfag
UJ5VTcyniT5sV5cfTQhKx7bSg/NafSlJ6wvrEFU8kDMYxEKioDohK4N+dW0XW1zl
EBtKrO48fa9ptY594a7Jedh6M7NL0XswkdKWj9HGumMcrvY7JqBKugB7AqlfjCq+
uq6TTL57pEp6KBBm3F5LsGnoXNCCNst0JrdjUF6Tu82f9/7Rs+AImBPejaPNrl7b
05qB76QnJbOmICaTVPXMEB+DW5oA8a8EfOg4O8eJR05LYF6P5u8l/Cnw/J3zbWkZ
EJv2W5TPVUB2Ut+6oM62W4UUvDMUExRuSrgyazoGWnyJPHl4PjdZst73Bt1rAhCU
hIVsB391ywyBQpVrIjcXfUUhsHxxAdW2a8GcJ9ph+5vpd2fTbzuw3DntjndFy8QQ
cKB68yG8TB9Zsorpa3E3e+j/VHeE9HNt8DlOjP6lT2R6RoNH0jvpLqemLotMd/L+
Zf8kduf+oFJ3wQJ4nfLY1HgS7cnlbpChXNldUGWPdCzWziu6qDo/lXl1a39zM9KU
4OdcJfgKQKmORxPb1Ek0BfN8gczYXWh0SDscAjip91zmfOiHnlYK9UMgwL0GgTsL
lYQYvmaGpGXXkQNhFRAKEDzYLlrr2WuymcQyP+HG+bSwL6zAKArTiD3vNWV5MtfX
ilqOfkYNC7JJXADMa/b/KTE+AcQCwTZQjIar0BxaP9kWEbcnsmMj3auPmxdz2b4H
Z6Czmwh+uCfwX1LKW8Q8/vIlOyu0PyXRjXN7kXY3w6j/TfARCCRKLd6zXE0nIOAz
ClrH50gWeX1OB0CjSuTSX459gAdAg8FRqBF5mIJukfyI2Q5S54n+XHVcuO+cv/wO
8Fl5qCNwJgCefmLtx1dldN5SwUWhCOldAFVgTs9edBt12HyHWckhi2M70ChAwbSH
yWDSuWJPaadXvIgwCz69o5sSzm7sgirCAA2+E29vjb/RZ0eXKzklWneAI/Z60mpt
Qbjy9ffpN3lMe61b8AAuBf0L2Iu/vynriMqL5sdrDLoB4WlhmWjkGI8VZj5XoSoZ
QBqRIisUJh6D0H7dlRJJkJ5ZOiWuXA4h1g97HgPtniKLyTZc1Yr5/NEXpkBrSDVx
tV3At2J23Elgh4UOhrcVdOgqO1py9+aoltyHvqqK0a7xNIAmEOMnbAptu5OnTEvQ
dnvlq3VqCCI8jIv2yCQINCC/Ao6PY8QzBt2duWkGe4ieC35e/7YocBKynAiUHF9h
48xgh/x2Gvuk6/wpMfAMxMF/AerCA7qcgy6GOiVNqNJsN8E00Te0Rq3m5OR4yQ7U
RbrRWgqZ6zH4gVej9SAxSSEsArvElMt8e1XvkKNIHIF3jSqQIRbTw9Vg+rOPS+PS
4kLLPD/iUAsOOzL5o3STCsj/9vufI/ls3r2tz9QcVRQgUOg1E7ACOj2FHZyimlcH
SvSC222VBTfGqBFTzUMutsBsnjUdOt8ypkW/xhaY8vadcdt79I674O12SHKDSyYy
c3DncpWjvmpgcNHH8eKvM4qhMVyBWHQ1XdtwbA/HUk+kkpP1RP4Ddd28uuDZZcMz
MKAtqjxBgVeUiEdqscehxoQk4ABZzo43dJZra4DpWJ1vb/PD1WW27KUKCZ3XnOgM
3sjZHXoeBEKFTxlOQ2d0SyI4W2cGRTh3HOCiSfObGKZx20Yq8WCB4CGZMhttJ2+p
WI/x3x8Cf8nU8yqxXBLxF/RizvkocTdMLca7BThagbhOGRfMy+dAKGUsNpd05Gt+
QuLTmpcT7bttOHoU9HhqRvzYpobvnJBHVVpLrZ+p6y2oH00549zVMpb1pNklOkW/
G6JeKyXOcMNTI6FF4VUUde5SjGC1chSvmCrdgKspEtH9NmmRcBSiEuleQ9HSriya
YtBBtcUHmI6JzQJQxM9yaWpNIRb3JUtGRkvOkoUkn4j/E6PX4E00Odbtp3V7CC/N
Ridl1eMzik+f8uptQG6bXMMPPP6RT7NMazqBBR3aNJPuPLC2XbXVT01jr3mb3Y/c
4GStGJjEPsExsIFzzLPdJaNZsG30kPMo2PWYtSgSoLJmRtimI75y9ZksoAXUrkoe
vu7ZbSQ9VVfeUkaAN8HLNfZONTVvBEUs81ywMQAdyQmUuPVvzbIhkg3gwNrjzmsN
e6g/8Ar6Z49cHAB2UTRmNpjYIcSdDgX99hYnnq1AWQN9vylmHXurnV+XIin8DhGE
iNk/t1rDBbDFd/FnqAhXLnksSuEOiiRH5/Sa9JS49sIpVrIoRRpoYMcBqR+PXFK8
qz11Itt9lM/73r0i+vcGGHnL14ORHorQ9bzIkpI+dMgus9kCrcSpRXTfuIwALa+B
NMuynTk0NRRyPRIneXJwQPzWFjNJLdvpZiP9SW1h6PGJEPtgGSGGd73dK4+xrlO6
O/tFY54MG5262jgJFP3ETZB6zlqrywVYg8wNjLPcIvakPGBTgG5SYQ9Eoqn9GnpJ
/73nUyPwMGjbOOnxpXFb0oKpU4/vkrH5y1uK/zxLU3hzCvRU5qYpN/GdQEApehXt
jQvy7daeggMBQyWifFTfEOsxYd3rak2Rt1xoyVQE8TbR5tTGG8lodC0hK+T+xsBv
3YzV+m4T56ZfLdiqKHCZFo7qkXgfd2NAcnWY3qxUDgMAAjPTWAOFrorw+TF76bls
VIMwhotTRUHrGPVhVFUYcsIRpW/X1Kt+ZTM1BAkWKSH+pR59+OnX5PzSDE9Roz3H
yKddDb8lZyJcwXwB3A+js1pzh0X5UtN77hD8UvxuVfivrbr30Z1TJeio1IPT0e+V
V0U+BSojE20V25cEndJyRCDDSnrzLiW7kYTvSkS5E2hDTk382xKtNRgDVwXuLelB
8yO5m/OwIgX7JjqM2fpStv0refhWz2aBKjcMfuINpOTROJ7SWPyvGagzJN8i/8Bu
wmPf1CNtyYqvoqzwSd20CNVRHVQc7B6KaUOCyidBNXPesBCmEDxNVbH51lr55NA6
Sad50XPIWMhtsAaqICqDldPR2cEEkPcGJ9lFoq9YzepdOFHD9lDlZwOdtq6aJgdo
JIfFQszrC/eeY9ZXqfd138BT94QdQApZucFLxtgBVjfG+X6plitcLs2TxVewoXcB
LvMFpHRfdqdBeMkpKxdEEoQiAk/wrDJbmwH1MPbljRQ/u0Elr7kC4bxxHX/7JqcR
6saJSDp8hI8K2N0nlC6HRDHuZqtrm00qGRm5OZO2p9LSB/bsWrdM9K0jqFwfYPyB
UVBm/KS2uDrhusMWHARMXN2/HAwV07G50/77FSRnhvy906D/XFt6CI48UAMej9EK
eRJGsUCijEjg1CcyGojAUF5g3vfijEpx9DTMKojBT6MSr3ikOb2755STPiLuI7Cu
Q0cWZQ2fQh/gqADlkgfVa7sdfkUyhSo/ULtD80Ae8kBqA7OvyXphJq2tIDS3ySst
BJtSDBBWwSIPR/SMuRW7PVg0T9u765+AUag4szAnlkb+tHVD7nUFdemnHPorWBMH
1ZSUSom5Hb8I013rVmNYTB1CM+/qtBPsDf1sUPXvoNSThr4qAch0aL4gcKChq8Bp
EgXxmJcO0x5iOjBFRcz8kl8VTkPcN2+meMQtn/vcZYsOkgMrTv65l1FViue9SOef
yhfBh58lJKfEu9+APgKCXkhLbQoMuz0lnZ9fBAAlhpsONIoXDDJXd5Q+Yb+lQpGW
1ZFNQplTHwDop51jfCT1cwq0amB1XECkxZHhUNnigshBLKT0xI7irQQR/gByd0Vb
osziZfcZqLfME1PwdqTAUZI4/W2A+D+KaQuUnKYJj/Oj9eMJZZz+HN9HOYSXQJwB
1axtpFvDJKvrCk9vNAwbLTVIHauY+tVw/6KuMW5Ym/hPsnezBMftGxIjjjC9p7x2
80YFmoXKV7lgBDjNWnx1wjEhRGY7EeROwU/a3qKk8bYWosL6KLRMjhiUHC9n7Iif
hu2l5KsSAbV6GPXfqsgvHKKmQJron6h3VvrqTJDF01QtORDRdjhqMgyvv7B4chMj
g5QAbSKL4XPrLtPv0wWip7o3zeL5dA4uIRcilQdHJ8egvl84Eiw1MRjxfAhfm1/S
qwTmt77dbn0kwBjjFsiBEZE98bi/MgHHLME7kKuXPrM/4t7miZZgRvRORF5KXog0
rsv2oOzV7r2KihAw8/9q/VE24da1lnhFdnW3J+2n85bdQEDWfM1eMrAW1PdaCQS7
l8MrnENKGox/EvZPn5+YeY3M+HEQ6xOF8fE+eYcKFPANEV+qLfTaoUrHThKqtnbw
DaGk27yds3PvJWYRPS0pCMkZKSrRf9Txl0APGtM7+bpxbT6YKh0JC2TNp65Ubrdi
WOH5+OjPhc2WsN9cSf/xN9qDC95OzW7JK4ahD7q73873Yh1cEauBI9CEeesJs4S9
Lw31I3V6DD26oEKjTcmvA5yKtksMvPSziaYbLzhEcht0PkJd1zLwZa40hRp5w1tO
Enqpzmfk1xqQJI/kWaMhqpTI5bEkBvwl/s5KxkjrefLi601pp2iyX+KQn1SM7cdn
EMKEzS0pVXN/ykB8bAaOy3RmonjlzFH9Jv7XkCEfOJTMNLU80RGR5BPCh2PgqUs1
c8E0U/7H3kM9hlcXkMULKNmULWxz69trG7Ydaex0SKjXcha7+R8wNGaVNn0nqIKY
jy3lY0G0miSy/qSFvAt8kyvciugSa2Og0eOsjgWRoG+1q9fEtHldlVIBbUIGvnB3
DMzZWzyCGsXwMDD+HK+cnNEBZ1uAABZMO74BGQlTfFIG4mpIsezPyGGxhMPHJ5Xy
e5irOBpYNUu49hWLFN/794MUR+D9WGYz3sMfm5DqmzPgYwV8c7khLov2yEzvM++H
MdYeKpr6MvWt7MR0B/ArAURhhm+fSSj5f6guXRlTENBCKswQ5x5ZnBjLEcysqwB6
PBCCwLY0ARkKPKXIyx9eOwEG5D3gItsBlY+yjSwuZxHzBGVA+1Z89O7Eja16Qhsb
gbB4YSieiDwci0s511Ock/B3rtmeNJr81FnbHDvR+cU8yfacFJm9WXuq/pFLPHkC
YCj6+AYq9Cl8+vdIGXk+nro+C2AuLwt+gSirg+71iaR9ojZsIVJrL2m6apj1W7vx
nDARNu6kwBxUJcCG2xBIcF2fcjuTzG7bcCVH/eaACJq89Em/wCX5CiVmaq17Uk8W
Bf6J79KpThrdSgvtUIdvz4Qc1RPUFk5DCBLlwIwylIjEhkPib2WPt6SJIQz4eNNU
jbXiWUMw7Sh7vfu8iZo7n45dL5ds3IKJQ0rp8gn3u/8tw8OUmxJK5zCT1IX+34aA
zqgBpSEXMN9Sa2KGsE9eWBJs++upGVO7rWHBY0YMau7oZ64cBFrOVarDUiJZdT37
0sUNQvqJXMjtqWpi8iFHqePH0/HUHVBp5cAF/r7IGOlnkT5KvK29NjBq1UT3bKNI
F/Oo5gxyKxUVncxwZdOAGXMlqCxyBVpvU36R66HdP858KtF5QCn1xKwfmjcJEIgq
2RiReFjbNDMVJfrT3kF7Xu5hzLhwLje1HJauVRw+AabidYFrcopDqVYm3aKrxqNc
H26Xsew/zAWm/BSsrR3bepf5YtN+4PiyKTN5uHn2CvxdhBaRO6+ztGtMkoCgiQXN
Oz8IrWBZUvqqwAMHpWhjI2Y+4hjUR3J5xyDvveQKSq0EJ5Zq2aGeGOh9osllOs1L
7FzWVT9NY6wG6YNZ1MEmNmi6p5XfRETZCcZoCNUVySzg5r4dAlaNeUlaCkDPahiI
xH6ZHmBHjBFdND31oirWkposACas4RUUjLqRxcStDCnQNE9Kw3b7Qgr8Um9S6I8b
H/Icz9TF712uvB/XKckoY3JIxmfKM+6AuXZkidkQAgzfQEFj75a8ZxANbWmOvRtA
W5pd0m0sBFs5qOmeylYjMLh1Im6CJnFJAerxD+t8bKuM8yGqlnQ3GuGgMWUcPffY
hz/T2dCkPMRe2bBqxKLRqdD3RpL53uzoH5e2VykaSgMhnKLxgDume8ehZVTUTXFK
MrRuuqptnMDHuRgJInyXkBe+57+xtS0wX9H0YFFseZm7RGqNPvUxWlITgh7DZ4YD
KjGsYYPBdR92TAi6OjSdopf3UrvqVUBJKksYntYRoz4UwbjSmhQSuTcOTlIDlM1p
Nam7WBO6KlpjWqMS9SfVwaKp4EY0A3ex/O3wdZjJqA/EwkxAzgyxOMJic4y1bzBo
ECqCtpUJleWybGjK6A2XUQ9PIgszxrAHfXei0yi9KT6cS7Hb474vOewn/fnhXgGI
4eTAUqF/9FkozVmUbJTjvDqzNVMSEfnHlMx9ran7JxtyjK/VCzc3sAIK/sjN5yWY
CXzOpQa6ycIjRQp5fXuOSq4iRZttERcB5SF8Yo4tJ8y5x+y3M81u/Q701aGHa8Cc
3BfznJ7DmWSE87iQ547jmGIp4myNGskqLy5bG3M45C88BujgjCWglOvRO83aqoPJ
wcyogbuQMn1zokvhUkxpiPGMBvuhcjTmNgnYM2u8eZeMatUR2dJjq4wT6+IBcA/d
M595UqwpnQfwAFL7y9bNP61G9XK1decIbBNsrXwD1G/OljF+Jx6l4zVlghbEQvzv
6gOuB4BmeE5/3MGAY4Q/L+YJxO2ec5ZNJ0ledrP5UdfwXMSE6o+dIxRJlVyUmgBD
yNO4W7B05tcDo6rDnCaYSNaP+MFQ74mitnY7NfNPdzapiMiozUVWmYQqF2kg9pmj
xInXaG+y31CA9QwLQr/FT2+XchNgxhQbu4xS9miLAL6xdcJUaMw4NtlbZzEuboH0
aq/D9oK6EhjkGyeGKFZhqNoSJwFJmW7zPbrklpBvn++oUbhLp0xFrsVVkLV0oofo
Zgz7YUGwP8DEfYrGLkqeMNFkBpIHX3DFqXQP1dcuRoI0rswzYVyfYX/RA+fJP8JP
6qyLoc108YKGP+l+wOn9zIkrMwEjCL7n50vvx+qy/Y8NuIkAMOXuJ2St2AbQtX1a
tRNoJ6EpF8tzzd0vp9+Uq92bZvdX3EDblwPeRG9yrEbgb+wFv3tUhmJurSaMz36B
2vqsM5SMRljS+qTMdmpGFRy1WQdK58MN60/qb7+b3qgiSH1PRSLtT4msUw9PA8pD
+s/97bC6u/XRuh43nCWh6UsJKdOPns/kOyA9TxKuey6oGcXbFyCsDj0TGLRjTNJV
yD379+EbnhnJztpIR50Rg1RYe6hqRvaPKI9pg0JsgmXc0kIyydi2E2qJQc0LFgCd
TPj7Zx9VCgdt/ssVi5J8SNPcaaPaj9Eca3xTpqTF7goG0BMkXb0+nrkxfv9asUcm
eaghi8qNd8OvlzTtEMikBtJjJELn1jxfCUpQdW7Ut7a0RmNE067jQpIb97EVlWq6
UXu1q2bvUE6cLDVWJhRCSOmBst2UPyT9vDpqeMk9lPhtpMbvNdMrCe0+c6QzdRDZ
xQLrzI9Hu8Bre05vQ46vqjg/up9vuF/Z/mjCxStKis6LZByKxGF3/n2dXqYm2FCj
E92ANyVENCrc47SE+jenr81sF6XQ/64Vjlp3BCy+cYbM7bt+l/qCNmcn1is3Qnht
/usZNG7DHQwACFOjU93hEuBQY4VFqrA0rmufrGLkSe1mYrOFc0qJoLqvklPQo0hR
nHpqcaNQGt48d7ij87l06mCSVoGeWyPikHk1mpz02sVvjCIWxLKxrbBWYTzRvXLU
OVQkIuc27QJL1TmbkhqCozwbAZNtplOLAPo1VxvObERkWAQWuDGZzqYLb4D+yulj
lhpxs4jNJZ+f83AD/c7oUzgLGSFF3sVAakNRfVBc8ky2yKqfnzy/PxtWIszFHZ02
2xidSpD64j4SIU06bm0U00Zp/ohVxAZBZ1QZIkTr095oChErt+B2/6YhvN63p9+f
jV5G5K8hORu8orkhCXlLbs1yAVCtuTd6Fb2t7Eir+J/PcgbDGBLoLAHOnnElUkqv
ava8vDo6vTYg/ODb0nbXYJ/sM+6vVuxBsykb/uSc8uI/cdcV3uVp3eb3c8MZljCU
+MzNgl8q4CEYBm1u1oJ3vUlTJCcIWZqssACxE3TqqkC4rn4lk5aPHnNg+VKuz0zP
XtLZCUrxoWjHEalHFGEkfT+sKSgD5FoJgKp9+EaKriM8kR2vDJPcVGHakEQgUTYn
OUzd65wyw9UW40nO2TLfNIeQU3eMO7W8SBxXwXM+R118PBjJFpLl//g8xRrCmdLN
wDAhnxqDEv8QCRZDb4gQeCuqAxWyoLhOZouXwgZbQTGRUYdC5eOCmsZI8mbKdiz7
tREst4wMlcnijkY9V8CseaGA/wB6Uzs2wlNtAeGf9z4e/zLTLYYxvek59oUXT4k8
uhjQF2Z2+xvokvHJcm+wlu9vwWpMtNSG+LiPoAf89k2u3DxYTjWZQkYQrrbwNX5O
ABaG1VKT/OpYmXmgZOHI0eFM5hLvmE+NaYMfW7alwmV4ksm1t1F63p4q1KJ+/dED
3AHf8nMHHEOkg+kS8Nl39J0gnoSJ5Mf6sdpwEGdn/1mZmCe/yIzHSxNgnzohgH80
qk006NpnlQcug2+gJnqOQrO1rqFU29qhoLDwQTpeldql2aGhqkmVtbLo8lT5yo7M
eJktH4KhQ3gw4i/hyMif3BOpOSsS+2MLrMnjPhaR/tXVbQAYR9KKadwIZRzbBIm9
wZfVDX9RVPs68DClPCi1ZZQA3UUcEMS89AWVNqxn3eem1QvlxThQbpE6PmfRdF1X
2uybWdDu8cQjBS4MrtCUcvGBijmVMWxs7hwEFpmmsUX3Jm+2mYwFUSryhVZfbOHW
eyAt5YbnQpA67rdTH+5DpM5NSJnXiriQFH2Tds7z0fcyTXbmzXCABNljK1o3KpIv
I8xnk8j3BGe3JCo5rAneC8taFFg0McUZFmPQOZPCqqPn+bkNrk63zNs305IlpV0V
1fXq5wXs+nnZJ7QsWWlAZC2rU4+qqmts5w/0F+vkH6LqPrTjfDHh95yD7WS4Xh6o
LmddsF0oHXgZE7xjnrIXIt2RGcgijvP3mfCKe9V4wNRucCFLcNsonnFSgFaVInol
4HdG7v4JQ1voKuAlJtlZHc2Ax4NHTvIjMmJA/jRXkBNJ2FKDYwZm3LYmmHRZIwhE
1mBaCyuCXZ6p2FcVQaL5uk/NK3EbhEsyjnaBQlotZ8s+6uA3YLQg2E9wKLDXrMkU
mf/tm4vD5jIJ+eeDft7y8p6a7jACHC7DY9/Ns5LrF6HKpbJxZTQg6eNJci9dnKaM
QZaxu3R2E7s6KoKVmPKutaBFgY7rCgPo4QK8UplqgOAcKIls/ar5Mh3iRgUQoa0/
RI7VT5BSQq/8t3zCSuHXHUFWFsLbnetXc4FZCCo10ahOKUz05NCDfDe9MdT4VBcE
RhD3IUPPuIh1CbLMiG8TxJZBL0XyJanCgHtr7AC/KvFBUFbe8uHwEyrenmFxrzpH
UyQ+MYflXCAUkY6EA6Ovi5ibAEl1gFCJR7jB0qHuipMl2ko8NScE1E5PLSREKzq1
m1P6KsHDETaIEHnkjXNYITXJWt65oVvxICir0X8KMtBWCA0pPscB5+T5UyT+LaZ8
dWOMgJ1MiTusf+ELov/w8IZj4QJnUjn0pj23mFqkkDPecRGzrlkF27kxUKJB1bnd
6OpTDV+nk2FX/yOpWSLpXzR9E4lFGVFZWRsRj+XHFH1lo9MbGeraoQjFfgE6OfR9
H7L/m2gTzRMLcXycqEDC6CyRhUtRBr2wInuFLsuUMsiucBj1cx8ll0jrAW8x7Je7
kqjljgtGGLloKXCt0Cx7i19y8653FgjOP9V5BnXFt2PRqkz2EOwgb1Qnamk81Ukr
jy+ylhW3IBgns8em0GmwpnU4WjFzdOX4+GUMPxV2UPe99bqF/pMYBmTgDzTCLI+1
/BkQ/8SLFKi21lmf4JgoCBOFFH208jZYlGTAsbZRvuouBgFcI/4tyqIgB3HqcKiN
B4Z6onreiIkmqG/8nnekkN3vdg933ar5/MHR8LRFoKh3DQDZuBfl87NkAlUDwE42
5RYiW62Zelhmkd4/NBbUY1O+UiRyuplVvQbdc1GzIM9djzBCoDdwCaWxNpL19Wwx
J1WZ5UHTOBNHy4EdFQxPHunnzwxjs6xG5P4HzYlcRydDVx52WfPvWU8hP2CDhe3f
kCWQzLZTnxn6GNtY8XFV+4K5XGF/z5bKPXJ2btFYc44mSlCRGNUyrE0BvKJTFZ1b
Ox9gwAhWfC6diGbJJFvAYx+/sxYIfMDsKSuMdS10STYboSm3FUqzDopz8RyZrstl
gk79/nlQ7F5HluC3fsnpzi/+k42oo9REvXParDdP9AINzduFQMshD4d8Do8rGvmN
Wr6053vvxnesdxf6CoJ2QuJYcn+SvyCSLbyAaqOPVgALVb2OnM4o7hWNOiJuitiF
Y/1J4gwkFPFv70MBKr3xcNDNexqX1R2/XDYIg2fyJuB+vYfX1MILh+76Pfct83Nn
el5dWRbxRD6LQ9Wk49tqEhDcWSmJ2IXEeMOr1PH/rBpstOrnlh1WIkWiMlC6s+qD
H05UIJAGeunbXN6Phs/HfxJxsV55iIohUc9vX6CS5h8seDNdPLLpwCsdVSMIz+ST
DRrT0/L0+wj1ptepPFSY9jQid1k/TM88X2h165+tDQWJJxJIMO7IZzYGtzWvJ7Ir
ttozBDbf0Cfar34yYvIfUxZWkuw9eDGNsUFZ6+Z4QeO3dER2PKbv08j/nfxQBdiW
AsYiEWdVEBA4OBRL3iiC4uhvevwOk6djE2ZCtvTxwsbCt4oI352/3erQ7PohN04g
vEXChGAKEdXw8whe6oKRnALLRKBEsQj4b0IDd4BI3Aiy7iAfjC+I9fVh8K2y6Dbk
voclmg1f2+gW32HufNt5BGp8FCQ2iXicE1mXNUuRnCsRkoU//g41TfVQvd02Adcn
vNXXKK5VoRQO47iSsrwFDbl9q5Yw1oESz8XtE6o0zP1YHkqewKIiAdYp1aPD+UgK
xU7AUJ0WxMogXjtPejtkovZGYXV7Q+wIxIx8dmuuZNFtZ6MpQroD7J4GfD4QIAaf
nTRbLCibI9aMBExXnfMUoNUdYYBs4VpQk7WryIJO5YPJp/ZW/7+t2NXSBXEsTydg
nav4d04CckFCYz8/vLVyDPIZqY4mWgWQ+J97goAbDFYDI5Ou7QOdNRe9kCuNzeeR
1R497RzI1HQi1LPFLvFb9isv9hGZI+T/3zA04nKoI04NR1GFaqjUpY5KukmkCdjL
lJG6eOOxzcx9tk4inWoA/ao8crK6tLcfe5GlepN7OIZZAEtelHwU4ilYjsyfmN4m
sWZKuCeK++hJU/VElBWd7RpGxgUpXQnP0LPQYNpnfEvL8ugdzpFKm5uxJ2Mp+Z6O
gBp4t/UXnWlryF4+zt6femCI+SiWMHGLc8NZLcvgV/8O0HvHEVqwOeY7KsZosNoI
QLP1ZKs2WPDCYa+WAPcyCsYpMAhpeX4HxBE8pYDiObHbpcY/uIS4rnFauc1u8rGv
BXhehZO79E4mFzyBFsGbB9JjPm+st81jY2gpaZPyEolVRShcODurnFjRAMcKuPxb
RGTaOROPM2kz9pqC/MGcZW05LF0LSWSvqvseYtbLGGnSXzixYy2wgBsadyRf/gKl
+p9ngkp2FG9gq7GZyyz2eozIZLvSGdw+urp523oz9bGPjWWU7dbsES6LTSboBy/8
81k2AlCCt1Sq+QXxzaiPT/t2c8mtrMRz5yvMFVUew8Cs3Uysz5HTdcjUaM8vqmss
esLv5MiEUzE8NdjaQ/GUfsiz0561ox8vOxgyUZNI0MID2sagWqABTnMt2ALmIlBW
3FZ/BgdvXxQfwBvvu32dwT3zaQJez6IC5HmLzI5Nx8uJty3YMkTvU6x34BL3oO1x
wGqext7c5mJiflN7T0qkMURq5LCueU96u+AdrUnj+Bk0a7CjZo84lm2nEuLvBJgX
raxGG73KwUNpovrsAK97huVhQ88suAgORLiAXmI3GPCWNR3hT4UsLHHsdJFyPgi/
U01D+z+sOHeUbpujgMu69xq6NN1nZL7AQyYcc5M55YculgBug1ZVjL0SEcC8Ycga
f81tBMQ2Ze1foCGIz2FS2/IHXdlUaNYms0Z8s3WEqy8KdJSFV+R1YCpjp+GZXEAR
coN85ez6VpqvR3PmPGbCs+QKJpyj5FDB270rv1DWbIlq0kDeCcDteG4y17hGkHJ/
vpenhLSEaxnVCc8MgmaZGXKx93CcMuDHJH0oUh/6ETaV1LvzJdWtjlUF0yc1/BVd
R7esvZHvOmkTB+s5F+KxKVlJQRbbXiWwHQklFguCtZktocx7IHVua9rZ3dwD/Hvu
blH7VfUglt9GenfShUY8CiEeH3AGfTA3kJDfXZoKC5d8Eh0x/ZhBBJzQxZE7ggGS
DsymoMtBp6UYHj5j4vmt3ag27YRw+b+zVjtUxuiFp6pebbfAboqIe+VGe0/6WqLK
zqo4ldVTRSvVtwnVSVXUbTGk3k8S29kfJq4jC5a+mt6EQegrwzyiQuD3UUTVwDlS
R9yoRbGT9TH4tNkGW8HAYEcai+iHCAu89FFGHCfhnp72vqOrh6pUg20PLV7W06mc
26Q/SbRGfZSB8ZnNlrl472YYHgJfo8/getZKawQwl/AGmWfHtsAabtETnDqookAa
nhbqgEhCEwnlbQS3rSI5pP1Y9WkV7kppTD8qgIaFi2EtBWxenHvxwnFNMOmMcG+r
fn15WMDjGaL9kWd51g01FUwjlaJgQORfzClnME/kBtK9jSDOw/HzPeCAae8amxrc
7OhlLsXAhfcN9flgd/99pSnn3mwXfgoOfqBN8oZG3L8NA63A9GEGYW2AytHBESMe
gztznqUyUbPBT3w4jj4s25mnkyf0YdA0fdcZjYVcB8CD9ILmUkvIVcR26gBPLQ71
1xE0JQBJ3yO+/BB02whCJuRHXQ/9d7alS/iV7M2wD90j3uqB6PVPlBDN6ezAJyAq
KDA5FFNXXHFgJzT2eqijNBbRYOqhm3EkfavJtFjB3vj5u71NPbwas+O7KbQ+WbmY
Zmb+GbVG7zP4CSv6M3YEp9nc4XbiV7g2P2RlLFXTg7QcX5J7jdNE2f1yLoULzJV6
GE1jq7GeHFm36V2avx07/dv1d+s9UJi51IADS3+lMrcxLMx8Ibrv8dzTAO0mahQ3
OL7AP4VmYS+klcAfXgYELSNuVtJ+3g1Ct+4ChrYt9ybyw7/k0Xa970N7bB+GY2j8
QuHSpaiOIFIGi/hK5FlYEVWUceyj8iwjJ2garH81tpo0vANQMq0nlYjrd4QYRbVL
xY0/42quRAEH3ajPA3cjuiJwlosULQzQdu9Jow6ly7J6U33zyrB34BUrvbFjsAmd
tR5LJI/CP/wpl3cY/fhuUrC8V1uG9oeujS0NjgH6Q0ifWYr84JyY2ac2FDrjyck7
lZkk0L70ilnhURzRryAjtEUQ1pC63DC9iYxi9boc5KiZciPcj3whvS0s/X2beaWh
Y9rn70XXmB6dZiemfY2T+HinkZJ9hmLlYdou1yxG9Ibj6JByYjLRCwXJRHjhpA4t
gpN18cr/Mu/O3hEPyEM0+gEL5wXAiBi7JsBBr26Ywg6ZSMxuYYW26nh9WyOg+2iY
pFU3pQ8FAeAEZadoRz4rHeGxX0yKbBTQcGSOvQasUQAmQZxV7w61H/NEd5s2Gheq
3vh0ub/OeJlpy2SibpIFXm6ABNRYYBgGARI5FYRzI3sMLilOWcVCvlUunvwg7YZU
rW/Wgk71Xz+qUUZuFQpQWTpobX8WA+rfOCAQqdOoTxholejOeT7Y393JIPLm6RQv
PTfsyv9mhbsKa9BT8gmVpCW9BwSEVsdQf1F2LIQIoB3IV2bKGD3kGwlOj6LZ6sRZ
Ue4C1WQQl5ib3juh+cB5FUs/OVP0f3FhsUGLFpzmUFihbWZxps9V5PKLcf07BSad
+3c9Z/FK0epHnUTOP25jGLSFzfkWgmKz5ROLJlObVIyQx+VgoG7NtkO/nxsAzj5b
VFHJK/WTmVcIZqI2AuO544ko/SZX56FK2/SghB4psgQhlNNCVWcLWnLsGhUJrt8Y
9fPOdtHx4rzHl9H5r3fmavD1zcCz6Xq3z3e0i4xhhfhqh1a1EUsx4gtBOqQ/Byd/
XlPRrh0Bl7TyNsl+mg24PFH4a5hsIBxMFWs2ooTfClFUb93RZYX7q8CI+YQk80Nl
jJTvnPdlJrQE1Catwg/gB9geaZecuDj7KEfHHxll425PNLBpjW9SrCQum/m6hD6y
gC9oznhy4A0KGh6B4z+cPvHOYpHmfSvqmrXZRvXT3zJCanaATkbCftgp2sXM6Gb+
1Jmn9+w0qlkWcjWCF5efu58GJlOKQqvKMP0kH2ut0d9aI6GlP6EHq5bXhkCL0aVl
ZwWLU6II2u9LguNM7Inq/dikU2A94SQ27NQDzLGRx3z26ez8mkMuvoksh4Bf9lVX
fQnLeGt11guUoLAK4ZADovq5rYEMXhKlDGy5MYrU2xM07qkVWzM4Z+9AC5kV8pHO
6e3rqy9XUAMDA7eE1KB9rE6vY6pjCk+ZWB78CnS2qriDVDVRYkvDeLqEOtBsmhn3
NpFsajOcKKu61UFvpXpTYm7h2Z96sermQrhKyDauuor7UHsDd46hzf/L64JeQoKV
5QllH5FRqWiUENJXQoQvvsznx24N/okMNEUREsm56q5ekxjHz8xvBZCQ1bnpDY9u
Xf+xwQH+HgjAPHXijCFyu3t4wbGArkq2uwtvFedU5UccmfPxEmU61WPZ6fjZSUvS
biGo2Z8okqm2BA0Red/mCYlhLv6mRIthHM3P+dJi3SXWDQybcEURWqiFPpdvD1/k
cfemrkJbw9WLMTJLDo/IbR1/1wJTy60Z7Mlpiw8oh+EgHKVVakbzzHcL6fMXOcLD
1TxIT2i72j398PG9agpsuj31s8iCq5lBKYtDOAcXKuiN8FrcKEg5UylqpkZsmE7f
xFsJaHJdm7hHnFN1nPlRzqcowEbfoFk1CaVnKk4vKK1R+fDRUmDmgyMNfFF4eWIV
Ant7/I/zlzSf/0Ar1GogrpvG3JjFu6WENjYAjd1cH+5HsFCuLJdAFMRrUdRgOxcP
GO2ReuBNWchcO3P45ZRjMeM32AEYNbe7ujlNvlamSiYmm3DRdfXIL/Ib2XlocDOh
ot71aix2sozL91xw4XoJE27UbkJY6YxcnkBFgTXepJ4gq1G0juG7wgfHbpAa6bmc
YfqvZui4FSlQm71uymovfHKXl7iuZIagruOMjG/o+vPNBwqinlaOm1ajXM6K0RSk
jpqvF2FzY80pvIzlCKPimikzUzevF2oD1beLKmHZ1XfxATZTxFZywfZ7O5M7JGLv
ssRAPp6uB1aX8Dg0O9eUCpqjMehRupX2tjel+O1as9iAaZ1+NXhPAHfjOvoVbWMh
cTzjOMm/AdjOcMrfInZ+1DmdNAX1ckOSg/wV4ogqZkxxVdj/8BJNXwursocULPST
qd7uop3l4QA2/DcSoBxjix9tFEcc/DsVBcfjJlrRvYB6/1eRxvWCGlCGLY3KwS09
NHZaVHkr0Gob1Z/6Rp+qWkQVMuD+SqSGMlCPkQhGqf5HUrPQU643aE55Di60h7PT
7RKUq6e6PZ/BUg8zbDAnMPBgBFcIHjm/dmXi/1whKn+/kzSfB/HYLqhgP2FCgedm
OtQa2g/SFouTazipikmD/C8pXBLXb/PWuK8XAeKDFqIn7FkaovcGcN/Is1Bd0nM9
jefHCONZ4I3UokAfkI51qSAzORNHufSL6p12Xiug4vO7vzXYiTGbTchkMkRWtBPo
K4VhegX9mXVduoAAQRoQJmOJqCT1yH2qI2zwmxuXrmRGBPNlAOQPspgwWJ1EovII
ZVTy3bTrbGrG+Q3+xhLlimQqJt3sa+8nAiHwLG7EQHJpsbUwIEgiwiroekk2I8Zd
uoxRblWlrpZjkAnwBxcxS3IrL/ehvbKEYdBB4NYA8E8NjWB5hD4957zksoqB7muy
H+Z+/g95LKr7WTEO0UHm4ISnHoaPnITNmoJvPecvMjHl310BsrB0a8/yZC5PbKeN
hBk7lf+xSbiBE2ooLV46dL3TLOluOdWhvdWbzmJaC0969LO6C1TuHb+1HD00mwBw
GxeG81AUACczr/btrQ5PT+I+1Gi8jf/48/OVcypPVFK9KCz3xHaFF5r8T4nWBPKZ
uUIsChA7E7zGvJdzrShCt5XbPGc0eszZ4+WubCSIaLox1LyFiAN3YeA5Afo1M6D5
+NxPfvQ8biX0uBXRyiXMcBWvrd8K0aoRO3b/6qqUZZlC8QmGfUsqwKTOHg68lTDH
Y23/gFtTjejM+pBdfHnDE8gLfv/N30f6yThNEgzaRIQ9J44fec1WVMeSTCnZLR4i
eRtPJAWEOrGar0OBmiwuK8O5tba3tFLl+z/OCfqS2oUd3pe/bISDoEqPUsgvf2Fy
uu3vTFAlHTHfW3iD1cO0VL7fVagJRsmh1URDySnNlCPz8uPkb5h+5TmdF6oK5MFO
V+eJ6rAKvDDczdJrrPxy1N3tta9NrBPZUCI5+hXJK9u0nzRYBXSP9Ka0Il5Ppn2r
LIXhuYqXCWapWV42xYvaQbAZfWnsEHOni2I451LD6PzQKZyN0YwDaLRDvGfxP4gq
nlK41BKmDJ/Bc0b02LDLdG8YEx1gq8D3Kjjs7VUFV2CQZ3IiZueygRdl9qTDJRZq
OLq0qkgky1rSp//GiTgWe7/V6rOzQj96x4PEA4yyQGsZyOFqRg/LRm/C0Dktbm1i
Bs7cOcqscYhjvjnM6ruevco7N5CWKCdRrDxqNE5uY78xjVqk1EhN/Kp8j86dFbqM
LB0MvKlLvPbIVNFXhGHihjX5a8F+ZPidGncycBH/7zNXxLlSRSIo/xc4/hYHWE4R
BG3X7AV7U9xtxXi+9iNtOUTz04eK2OMd3kHyORk0b23UBwGqXEl504Z6CtKnqNVk
0T7ofN+CDDYaF4w4G2OHPt3q2/4qtINeNa0eqGVo+MlFTmElFwYZcAq0ZyAwGyLO
krcYpcizUYCnghTRQ5mNVB5G9R1fzzcI05ci2XYsacFg8xjfxRVG9e/A93zhK/Ra
ozJRck9eRJVes0ay2AdK6+EKPjnmIWncpMb0h91IhT9JQGdw3zVQkJNLbXhlBIdT
9O3h2wcIPSvX3/VoHwD7SFwL5cphm/obruvHXzOAZXxnHjz66JEEFf8HQv/xcwfu
+E9Jt3wkAEk5vJvBf/+YGIEpkaMb7ybYxTBlI9TfjMS0Du+b7qJ/vW+aC3VQi9Su
fP33s4FqBU5uaAQ0x/xZ7PuJP4459br+3jTTmFwekXF8MRIuLpgrmQyQ+8UYHq0w
+aXTGMbS1NbjkaeAY9GFV1xYEzaJplp3l7FKS3WCiyFjHARtq3mYadkVBiHY1rSA
adfYf/zpWvGvU1eT9dGtawjKcDdMLR1uhINzdZlrwzq7Ex09tZR97PPy59YwNpHq
q3xx0Gb8L2Isx1DMit8zfEfv/4xZCiyvE/kpnIuceN1LbaeP9I7IUyl1W17Vhokc
e/7sLqIGUZoIbNxKX0Xmjrx/0GDMU4jCRmlVex2Pf5ZTUqxqhv3Xn4mPP0/cUFRF
R/0J63AHXZYs6qcdCGP3m4pJIhsv8B6tfpqgbrAkoFxUtuQlLR1uc5gmmCyuG4eC
sr+MUAYPbfXoZ0wrPDmMWAaFBUQkngWPj4PYTCQ+aR53Hxm1Rei1HdPtnuhWLfi5
XE46ctHl2kcgSfJ5koZv2y4wL2VUN4j+6NtR6zetd5hDdfUgI81bJ7jurFmtFlEU
qblHZLrKBqJCl8x/g2NHt2smPfs6DlECF0P9q1FTaiNQoXZnsXP78X3QTLtAx8EE
KHqpoB7oXxVUbX3ia2MiY9JCDkfjS+iyaXXvLQKlE6rrwzLFXG8nUoSm8dwWawaZ
Qxz6Jt6CLy8dK6dslnNcC02/A3SURp66gwm8mWGnqRFBiTKsMCykDhZORLD3X1OE
qycq7yrFH41PX05DKBwUxuthOz/IxDWh+sHHYWFf+++yzOSCNXCNdwPmpwNjovpy
rJLt0GhX5yzgf1kdjQix1kaGc5kiOCR+wySK+JkIZghAL6PB1v7oxRyHjGbfaTvu
clukpm4Sz4aZeA8HlXt+m3z9Atst+lMfedIoIYSC1EROYBRc5CXS09MEA4Xg6HRK
Z/G6jUx2LvLsuVn1ZJpymXj4rHK0iX7l1dOutBx5lRci1pC6clHF4r8fnv7jt6Ch
vxilKF7qG/fNH2wrUSIL9gJXdJv6W17HwTZpMAKXpqrj5U508ATg0W9nVNm0C6Gr
SRNc03XeD4t5DTLS0QZNeN7vhjCT5q1L0wX/GUK0Y0pj1iTrDMU5lNzNSMamV39z
YfSV75/AyV53uV5jPwTzNtXtEknNTAvx6ytCot3TJuKgIztJ/2hKlnb4mX6C324Y
2FLC/wA568R1HMj/OAOUG36IFtcYUazZMQwcsYPS+joT+P9uKgh9CHjENxktMvsL
bEobTu4Zh1e7NyIGG/wMhVSxzolOwZR28yuR5ID6fRKSDzEUR7vjLgjEXnvx5JRN
TJKKR8hccaUJmP4P+53EPar95Kqb21WX3QjO/GUOH3BTm3gBw94gfmQ0hDF1mhcU
HcfikoUyEmACZ+ldeXzH+JZx+Oj8kO3gsHy9OW8pCpurkNojq6wP+85ZzFJKlKqn
XuXYtNULLwycrs6sXE3AVkQ814LupUnuztanYhPfRQxfU2k0oImVoVVfdLHrXcKP
sfppdp2U7HMTqvkfCheUmyjQphi1g5DDUEM7zSAYs6dcL4IVi277ipZntvplmMw4
lzFbGLZtOeLyCNzwEF1zd7dXD7TRwrN+XAq+JXwrS0XKtK4ZGH8sWrmkULS6yJMH
EpyFnZ07qqEZP9vJ6G55ubbfFTGblGHnbjfPfIbYw7LuuKBUsPm69ukz9XBMXnN2
U71iHceYG60u9LKPgfOcdgRl6J8ZYNRFPTJvZ9YrSMAV+IHvn5/jWlchKV5faN7M
JFoIGcfZnhCXqTsxmE7nk0j23HxS1MWbq6j/gvpM76E991bnUvq7yUP0LVZHrzmS
uqckvLHlxkW4XDnkEXQ2v803bfS9PH894mQWp4q8TmsUtT82ysn1AE624xM2DGda
TotbAY4Kcg9xAL3YrK/xN6UL2rlMhlFRhgdL60cL4BXueM1eU3RBN9D3QXuk2mDe
3G/6QZF5iy9RxS7VHrfnSXOn/55/XT873EkC8U/prMhKzr/Z2EfERMpvVL5Xd2Pe
DCG6a2IhdQF5LCRF1S/9IBqZ7I83tNQLLjRihJrWC/XAmAMVN54wznBVpKLq0GvA
Xv7eHJImIzyuCmwzZztGNEalIzw9hdspzyhflWNE7U2VOd1Uw0jbufOkjVAtPDpT
6AVj/jChMHsG1MMSiL4XjVlF4UtW1WdMvil2SxKsvO/rypi/M1g1V6ilb8qQTjiT
oyUUewqMHC6IScdebzfSd7Rj241XG/k/SGcw/Q8fYCuA56+BimLDDABOVDzky8FY
JwmTn8xnC8vQIgWvB8VMGM9AHlbuigCoG9RuzBpWXad7mcNrzC4f8thvVChzUsDI
YJsO33K+eNHCyHUJTkwaHmveKMrFkHqGaeEn6YwixLrqw3O4eHjoqj5evlsZKOzb
AaJXQ4lXRxNhEbgPjXtbO1qiu8UPvdg7oGDLjrDfr+/MujdDf0qN3W4kq8GIlAZh
5lRVinWrPGk+9EUBUD3FE1vMilzwmPDT2agNUFMl7/YyG5mW9NUjXo1wLytddL36
HIej3Zomtdvh4jdUDAbWrbYYxD8i/E4x1EmTcViSWOKcmnsXhgQc25U7uT8sjfd9
CMKufpelJvEzAsuDxpkzJYnjOpNli6qDtMsAk/3OTQN32TWc969xrT+x/1FMqikU
1OHZuu7hNl9mg5plKzv3RJqTu5afGQ3Po/kwtrN0rfbaJpNYlbWhuaNvFvG8EJDW
f8yHPFsYFJX5CCct3O3RdwWtQnK6PBw95YbstQJzsDsofNDOCnb104XxiP61ZT6i
i1AXAiHi5QfJWwoz/5UKln0DPvQi/OjZsgYSVRhHV+LZNQ6ONaEfmrRQpyzs8iN5
YyrLItBZHfFNR3ghNdpRd4DvOy0HZ+ETRUmrozx4xga3BFZ6iT9uyn92Leo0nlpE
24iWM41SlWJE0RzaMJL1aEGdgfPsAhzedLEOwAfpnrMSJWbJYnEgKW3xpzAKeQwz
Tl9IRTPy3s5X2Ogz+Er0V5utZQJScLC5+H/BT2rvv6qkt+R0924ruelN8GgJG3IA
suRSLS9KYMrQ3UOEiILmforUYrHACRbogQMauxsNuSrNHE5ta9ncGyDL1+Qo217c
38xrw0TL/W5Rw7fFY5x3QLBbaH8CJHwVpXYzqTtSiLALiIjspHDyUwf269awfBUq
Gb13s2CKu3v2Rxq7tVyCjvFtMAfDQ1djRvJwS55gMP+A5Osq5saaOrB2JWqfey34
Jk8gVwvjwZM60ovIa3Oe88uJf8eiBLVNkpmttPXHc/E0C5mLvkiyfLxHWG1m8hNP
utLxknJ8AlRIMUiDiQjO4Rdy2onaYoo29H0I7LIiCy/j4iRyhFEnJEgFH8Pucqpj
369MWjrWAipsWr7mVXMBYLZJvI05dZc3oWDDnQVRNL513fNX30kfuGI3UHeE0lt4
zayqEKBWf0p4cBnuh1XSAR0nANaC8sOUkLeiaNWAuPnC8n5HpBVJnf2RV/E4fH1y
ifwlSvLUEYHM2QrUA6VrDi+V8pz+QOXwso//Ldb/7Mh1XL0J3KK4Er/K5JH+d4qT
rvT1ybxVs+FtzrawmMBAeN8gc+eSeT3T0yjiTlRMpoxAQV+z3k5e24wxNMWkyyys
7VMxRhC7vHS8KGtBZWF1qKo2+heylyQ1AvY+OmcSsccA7A/ZiGcpn4+r58bHtOdd
Mano84uVAT31zo0RFrQzPXTWBWWpDf0g3K08ZRglr2weSDL17qXjdKOJcu3LzAKD
QJq5bx2bJLjsxfDAljml+KLGZF05g1vekSiIUOrzwCeAoOXNHOKOll9zNQoUAGp/
3tZ+Ee/Z4woyVyj0DTwY/RSY//R6Ew/yi47RVEnxxRoT07crf7MgCCNLEfgcJCps
IdU5Gfk9iHhoxb+/lCA5i/GGVhqu5uJ8mos/ea62Dw/3dGe+29/b8lHceR57yyVd
hskUkHCFpRdzZEciQQzH835Ik/WLUnYvo2R1gJKnSICpg6FczmvyZuJXaA40lzDS
PUxvphUyqYthRJ6DqjzVlOzdf7F/dofGaqBwNK0RyASfDsRXHe0EgscFI5vBOEeQ
PJ2R5L2lSuJOqALpoGotPvOtBZ4mfVdCF0yjsKr4fh1QezkMKWma767nML+tg6ha
zEsP6z0dJULvQQ2593wv25vhZyB1ZH/qPxu/jiBxO1QH4IGfpWZVTtj7Nj4UWQnC
JAZsKMMxPqWvpT0rB8MtoKyNucmqC2KMpBXdi13gcY2lZP0Mk/08L+mJcePpNYXR
bcJC9yFBU6Kzk7mIUy2ZtD0IA6CNRq3ZmSaA6feJ56TCcuGMl0167+0yX7CowRqa
BCVuVZ54rBaif8CkVEeEjk/gYSgn3HFIP9q6o6XA7b4uObu6E/QiekLNvtwjqvhB
NNjmEFB3moO36CVxGjbh1mAkBNrQ+FUpdTnLXyetX6pY79Krx+mwqfzgMTEis7X0
atTSDOmNWUN/2f8c+N4ahj4x/Gfjhh4gpx2TISQcS+WCgX2LF98Ylu44buW7w8M7
TnBUB0IU9zlpVCrEq27aXlwUFaLvHwYsRvBFfP0HOXl7Gatt/VyKtdjkIANcUucy
nrDS3MuumCg5fCkmu0vpqwrENMqa3ioOTW/zvUaBF0Fn+3VSg63Ihih8uQMtAgfy
WJ7e0/FN2IX6+TLekeu85Ver57IIvEZNFlBrBNNv34fYF6IgLxYkve3VlRFosIkz
5w3yZVliHYAmj6QhsTJNWA06l5TLqLPlF4WVDAh+9BRfa5LKDgbCgBkV6JBD5u7q
K6b/P+j1OgbjWM5t1O9FqfYJt3fAOHWIl1FAyC7o2OHf/BGAAY4ox36BVFi3f2y+
pSyiWl0zPVXqVuHGGmCuwabmRQvHPRaBDho/s6JOBpPdGc0ezT2MCOnArmL9sGl8
mRPBYlZUPKYOg5heif0cgspqiR4jM6SZmenqsXIb3yqfe4XgFr3syEnA+VQ+4KS9
rne90g/Mrpv8HBsviLXqIrHOD6uwQmPeTU+DzCPblFhgA8azzRIFuhn+10nfYYHd
zh0hRecHTLl/nglylW/GcVkNKvEfGT++hZd6xflnKW/ddrvGgVpulLBQOBZurDo3
nK4v6xU19KFGdCReCyMnBokkf60Xg888/gHz4bFzhRUXk+PFxfzaiv9/akus2XfI
7yu1OS0c7H162SuMS0QzNCchsOKYuJrj3IIn5aOYxA44KOzcz6b3OR4sd3O0L+p/
zJNCaH9yYhf2ZT1Zoke1Q7F8pFWeQrLxT+xDWMTeqtGlY9C19kcKS7vgNzwEAI2M
7wxIsBFUT4+40KOKgcjGYVcFfYTZfQ1K3dkt4lUfnsk9WO6oqJYPXajKjCroVHyy
awgJC67mBtcVCXDDRzHWloD8/u1K/nQYDr34JwV4/zKf2fI9lx07/Rpy4xWt0dhP
T/+nggbViko4n2C2B6JzvarrFMgzsCB7Rcf8ssNBOfDbJE1GRsU/pQjb0JP84kEQ
eupH/htmCIbXNU2suh40UXq71jUNl25KdPlNZ35yPOplLs/IcJcmFN1RKh/zqc/Q
/j3wW0CpOFuME0WVzhzfZlZOsC084vbMsfjknfjbUMkgdXnrY8y6SLsGrf5PSF6I
+PBp9JfjADOewbzeUoB/VMzAHR2b2ZMx+kXeDRba3mbk2Ls/MRP8p6HRMWCTfOwq
l3XQlCKYmvhptc+X59YYbCvTMAwnF/XRGrCp4mSP+AfF+14kvIJQaYfSyFl5A7dK
GBuyF7TfCVYxbpDoVb6psDEBa/C18s2JZPqa7/AabFHddZkXjtLgj3jYCGf+nlwn
3bt35WSBbTUQKTaAhMZ/LmJKqmoI8RWzXehtq2RlivgHca30YJdYSnsdkl682cTq
lwnVK4t9zJYHZYXwNumOEEI8FtN+jpJTTeFnZTulAIEFAoCE21QuhDiQ6vUEeTld
3Cx19W24KxIVt5cI0qJ7o00S3H+FSvDM7sZgsxeGAFYbFFUajAqxPsy6TS1R4m6j
l8heGVgJkGpuamubYhRVWTKoKDVjwE6g6ppGFvtpHMJgVD6K7wcA6am9VQzVLUtq
44p4HZDialX0mob5/C+Gphi2q+ns4NeHCIUZU+l3yMkAtRFlkPv80V2mgoU4baO6
pFCeYTtzS4/fxugfWdiAKGeT1NVo/pgWjRyjoRedoFERTF84D/4owr82CAECPSVw
Bs8vQm+VpF9b+zAltQTq55kUYXhBCx2UDRqAFsarjHTmIa2Dj+tIklXSoC3SeMzC
W6xNa7VP6WP/O9Q9rc0OVhG1KnpBjJSSgvUtbGO4eUMg4Ij3aQ+1Hcw0YzUQNJV2
btNn9xrS17rGBWWtGHe5Lw56+a1AnTK7hdhawHaHKoptgmbG+HE/1Lw5gyZ1Oi6j
7XKSRNos+WsQFXJKCq0cEEJG9wN1+xu1cq/1HqacXJY3btTvEx7zYVATNU+MNQN1
ZnAjaUV1iCHq5c4wOfBkg5T5IY86wP1WXMcObyOAAyoioxk/u3wDZjjuhj7uXIQn
WwauD7I3bUN135ozmxcrbovsmVrYVomXOxnAHEWC4jwHNHTSAbpMyMEHc1m+b3LI
zuyvNDwInUhNQTgHpwt4xU0jhm9TA48nRC0xHv2EMPXKIxhLc0gPyrMgrevVNmPE
xiXBpgjjSiXGXqxHhL+yHWZjIVbSsqfDuc5HJPVj+0paCFKSfYpuBQ16hGGxo1CI
mr7ckEwT8GjlVnC2rmcuGQ2nJ+Di0Cp9IfXXcDEqQeHwMymIwWhQlbhdkATGUgnQ
WQ5zzAbZjYzfs9p5VBqrXoLh4I2llcMtI5vFeVQRcRxeKSSHdiE42wGoJM2BDTod
nPX9i3irVBQaiAaCz0CLWql1dANusR5842fDbczWV1wypl5LuIcXqQ79CrKtrTxk
i/H1CgwXlBHS5ayw1DzmU3Pdgw22VyiEifqfLOSbLAW6GpsXMwvNovFdYF50wESG
4i64UAf54i88UfEynTk2/tp8NpqZg/gXqp2qatizo69SJJuzVyWhmx0vA0U0ta+D
fufHEsVGZ/PVo6634J0JleTvxU2e7BnRrYnUHRpGBDp044Ra05m7QYtgsqM7FNJ2
HxmP1R7iuuarDiKzsTOxaLrddTMn4Cb/flE2dU47xN5pOfbC37IEkm4jre8tdgEq
g5BkjvNCerExGIBkqFFXQq2Ek1WrDkw0CAL4fjcNe0pvT2JPhrjz9XXTsBiphRuF
8p8s+8NbW9dJQuOmxblGyxQ/bxr2GeQCyFYZu4SECHIDRaKqko6mKG4QxMAdg3Qz
Ujs0D0cA8b3+XY99lUip72f5+kq5Vej8ewu11k4OTC5wcaWQ138f6FYYI8ELcGY+
WZ5ic4j3Yx1BUt12nndZWhJJLoUUBwTKNkqHrv15Y6uCEyqo2wwKzJgbffOxVBIo
OrVWtjtYoML3/sErVR1PKwAyMCqw+oWQSE+feGMnLdek5FatANrwLSta8fDTbtWa
GDVFfjwb2Dv8f0gKC2t+my88Iv2pVTbyZvhD2PKiZ60I6Whx5TVkBgcCEYiM99pI
QdEfcS51dbeTPR1kEFJ+FTKv1UcCFrphKLPipN4FPXW1fPJatu1BCbXIpu4/SpWE
NdWEqSVhPDeF5COtyQ44Ai065VatL242TztsBOwD5u78sH39sz98jTq/H2ykXcCe
X95LQlINH2YCVfmeJjpVIGMABcKWTynrZ66I/uWDq/anGLHf7qOE/CvpRA/iEVsE
i/uyzCogH9uPeC7rjRoYdMQzy4lqSFhY2eSk32rzz8twRsQzP+N2GC65n7d1+AnD
HaLDm3EE9VratuCHNu/Nzqr4xeWuFSF4FRCs4ubxCUMG8nVOQUMyrBu9cWvy4TZI
eJMT64fXFpI5g7YZ5uy7s9S2oHeTtcmHrbZiRUtqdVM3SYwG+RIWl+ZSC2l/Oxrr
h7ESkd8ueV8MHcEtZOixO2fuj2arJz90jjdl6+bW3LnZi/T3vIFYzJYjGxBkcbfe
ZhtfBOlTR21YkgpVXQz3T7Lk8BUu23H8e+ccDoFBVxICK0GtKTzoPUkRxvaPm0NN
qDj+snC4Fcy5aQZjWvbsrPArAm0vkmMJKO/VRpGHYGhh4ka4w8o5c80JS8cjOvlE
xF9vSzUlhQ2h6eeb29nUBeW0fQMze4cvpDy2jMTaHHAj//2uI8fZHi/KnONwRZ17
xDE2/pdcoSOas7/mVHsWzBdP2Aif7vxTpPw0dS3bI2qlGcdPwgJu/w56zj5IfeOA
KEQtVwG+rm5RAEugUNUh2+S1wzjfepv/wSCBG8bbJ4d1fRONnz55zXsjZwXA4StD
Chd1Y1jjOpcpTO71iWnYXoN2JHTB15tJ5fdb3D6KIboeS3Ugve4r/yhDvTaUtgUZ
zXKeAyF8UGzmrXA2MjiEtjIn3Jn6mXEl9p1OIpcguZvzv28zk+8e7tHNERkJMGjb
hPvm4y4O7vbf/vVPaclJCtTKmoHsDJ+2zo2CSsW+oJx8tpCVDi+TB/EBILeZewBf
IJkL66RDkUbQ0JI6vZYrmAgmxAYjOC9V/3iBwMiIxgBOtrt4xTai1HMY2jeecfyK
f3EmqUHoVpjlAQi3JykpNZB4KMT2sfj/a7wy7qwGa7m0eXAIKFcsHIIfeXweiEmp
hbbj/U8CVzkfVtfpxW3SdqvAUBO/tNnYiRVH6XA+bGHzx7xFkuCz13bTxLSc26Ge
OP2BeQfWhF20zx4CdzA7ZoefFZ0/lDJBcCFGGo+NQc006FUpp7i2pcxjrHNNF3Lb
C7wx94uzjCBRdpeVlg7oqxt0cA5n9BrCCSZfZsfMnHI+aRGd91so/LrCtmNUa5SW
81vhIct9+34FhznlF8ZB2g1/peBLZVp8078HSLiB9DlKK/PoTRZVu7r1cNlhafGk
v9vZIZl+wfY4bvl6BruRDxjnKbzXstpHnXhNUA3QrS3HdjrKyK9FbtwZDybt9lhl
V/uRpJ1MBW+WP+4L/RDIYr31FaDU9DpzrocdYZ10kSXKU+Vti/oQA2ivMva8mHey
Qd5ja0QhfOBEsjwiNX0BeefwNTB3Z0JTx+Q/lhXcsdNS8VVbvYnP3gH8rVmQiorS
tk4sOPihW6dK9V6hbZCIa+EyKqCTW4jjBbgDsQq+Jpsd0VmGAGgnxRq2mMyFY1ct
i7R6plUpzIilTFgySzRYsWYYPvrOGV4NVGWIeH1al3QNUMjJiix+NZ44rnwihmfh
o0nJb0fGyV4HTTZmYMZyKVO1rmdzO8hagkySW2iLnsg7MHEqaNA0eKQq1UWPe3Sr
zL0F8h9CAWZrULTTa1JQJuSJfJ1MO32oe0JKUDH1BD5ZJZyukZjq/VPk1USsYdPY
aeFDqiHPKlA4ucTuSNa/J6lhZKRlHMJlzYa+M4xaDirZ+V6QrPv4p4auJGflo0sI
EKkTtReft6dnX7s6o2cchugb5ywp1nnxkClb6LJrmGh1v36Tfdbay0cRwAMTUHGf
1byycEp18/Vl/QTCvcKfriZPOGF+gD6nf/UAuWL+fdstDD2iHOfMaKZZkPG613zi
exqAfv1IuIh7lDsl3KGJWocF+MfOtj7ocm39mVc9b2PHyCCo8s5jXTUngsZ8ysvo
KJkvML47ajQ0rEAwN7AgHom4I9eSCWdw2nQn8gsZlIu1aAkVp7M5jJ7Ei7QZUm2X
LWnJ0o0ekw5iHjgarmSBBWkO3kRe3AWeVAxBP+x2jULHpLlZswIZxemcDbPQ/V/D
qpiP8pGsq6hJ4guAw1SWIkLxbgO2zfOpZ+2QzMv00advhB8yU/XOFJXC+l+9l1Ao
dBfcEG87VWVI49WX8E+PDMR9QXp5pIJjzMbfHoZQNgHMuOJBDMtu7wFBSWWGXRKk
oSqe+OiE0s4SAdDQRaneJhPbZ/frcPgH9sBz42V6Zmp5TGS234C/SQCm/0C+YmBG
nNkuzkB42pmHYwK2YstaObwQ6NagxIxfnkXC8Esiu6NJZTxQNPrVsQ7lz/YaETn3
ons6oHuQjs58ufozTaZGCJEXS4bPFuKmeShuuXplknF1yndh3MNLsWq+hloK1YE+
JMukMtEhTYZPeEgcF8ETVRTSQRPzfUtPDhoUosFEVJ1MCQF/pXSJAql1bcsoqr8+
7jmFmAPpmJYcM4eeULy/M7Wj57dKdl897f/soabIaTU8Fe/3VH8PFJn0XE09Nczs
3MxVOKIsEs/kBY9ZM2f86K4SP6FiC2q/5FeCuG5zncuAm7sGWumVoxr8UCaMr/aH
j3hl9T0Hx5+qugGevKh2u/VnjggD9Ng0798aHLCg1z1c0uNqfnPY1xk3AA6OscxF
Vhz2M+LTZo2Arwm3+E5furHDyGDxR8bpIIKUy6+5v4kztTnOlKYsN3GPKU+XX/rY
RTPLNIZhixSjUxk7myb7imJdTo9XrKtgP5ik9LX4B3hsoNMhtzIolPocUJrvL+Kn
7E0J93dGfiYXa8r/QEbjanquHMIpsdZPNKbTXI8HdSOkBI/NB4hhER6OiNKLTz+c
rLoWhCbIN5U2yKkGfl9ZW2nSzgXOC+xJFhsKXqggRKbCKoale+2zbjC8t8htmyL5
B6WsncsGBQpZR+y8HmJL9Mj2PgNHWrEU3laO038hFJHUd0jX7c/b0CGkcAaRfrVU
/nwuwFvj41s6eEd1505wMhhcfqAvhpAwRXBsjpwKq1dXkXfgfI8sHKqXC+aRlWp3
1Ie0PlajoXMQTsCwl4OXk9eDHg9FTyct7iNIjONWMQ0bB/iYXrVL3rYCVW1/AOP9
UEHMR51ntm0F+aTSl93rLortiumFeRSF9SC/+E+9TOtxKvfxmiezXCT+vmRKp9XR
LXmWl6wG10mVtqc+pB5yP33qBSaFV7gzUjzs+E+Xczu8+QqGuQqWDmupIX0yMZLn
FDJ4XgwM1ZfPsodM/5EJ25GtiiB2O2Q94rB8p6Gh/sJwp0Yw7FXLuBhnnEopDZLQ
k0q+NSQlvngknf9oedV2lURpFtle4Cl/JY/ea5p4qsVX1e+jRppZefc+r5XcSnVY
sE2MueD46XeWeraj3ecabAWTXr2RV11+Bri5nbtkBgS8zKjR1AfvHOtqSJmsgZzO
EyKBoeIIRzvxWG05n+Q3sQVHo2ZuD3uWZtQvolOqvt0Im8sZ8RYz16i4fguqWaVx
SQkDn3dkGZmrzSjHBlMxUFUhSv+PlISOw6yBZv+/6TOTtKqGz+z1PVz7m6YfkwBz
/flU17PNmaTdJ/BTMwhsSgSAQmhpEoIzaepqFBcdP/QVjY40kRtLm7Lkp2yui5S2
WjtpnWe8TtjV0YlWKsGgHLpGUUdPzUgmXvtJ27qwrG04vLvg18eq/uVbh5AWlUPV
K24FPVgTSElpTi2A2Bm8zN7JlqXCAs2Oqgs6JyRpOX2Bag7i02NFRGaYi5CjMn9n
jBPF/zFx7GFbRus61HKrnoezOqjcAxANS20pR1WWkHirL7s1b2AGD1eOUB+7fEqu
FWG/NhGeI5Fr5owj1vACP8z0WBPS3ESfKbesuaCLkO4y0a/3ZV0HsRSdxIUwk5XK
R0vKDYZrG6c+YzB8gYefebAMzEvTZMoHEG+28BZ1ixAe4BkBMCgQXc0xk4SmmHyj
ETieE8nAJcVus/N6jv0I7w14yR9UZQmkqrSxHP7xRiILN4XJzxhBdWDfBGaV2slE
4I0Pf6lcS1BGezLuEzseHByXd1LeKmkOsxIo87fxJj2Tz7K3+XHGL9kg0dPjCvM+
+9NoZzRD6wrlVf19wcasAvHYaofSMb3h/N4VbfhA7FA7HCfh3xhByHz4DzcccXGf
PWwsW4uv2v7JG2HZEZxxYKmjO30tvhyTuVZNjuhPJoOVH8jQAUVL9xBmSrtBQWnI
GsJQUzWlWGT3sGS7KtOM+0CPR0iU2GtZlIcFuP4OhMAoOQ0NKbzDFevnJFp0hT79
J42+lrIqwf/mi3imvODvav4mxWWBhG71FWqF9v/SyCSDl5Z7YJ7p9WsvSevngWSZ
4gHtMM4TlyKjQUyPdono+yYsX4AJc3vIORdEeyhkjM16C8SGF0TPBI9TRPxzm726
ffZhazFI6QmHhGUAsz1tthbeEnJKKXVbohpGNxy0wZhPeIKyiuJjkC/7z7iAMv45
+4VpIv073dLRZ7kQyAMgS4dLThG91gk6gskSaOy85DXN6yI+E7m8k9ZY5wVCc0rZ
L6xrOI6DkQSKX/Z7C9dDjGNWaPmYqAFSe08Xf4ncEgoCHLthTIn4pDtHnYy4f7Rn
IbjF/6BzEyRltuL9qERbo7oraxSvhaDDHy3VCd0WGrGxdc8tTXrsjckOIlUgonPb
9oFIuO+jeNRCcqpg98ae/ArNxFrHNryxyemJRJeuH8QVSkrupqipZFuUlvZ2mPSg
0gZV8lvHeefbjrTWwqsUDuRJDCDpyiThqkD8XPiNAvVjLG0C1Ngmvv6npvNrbQyL
d1tELTGDw8Bp0IXA5z12yf6/q1GVi1gQ9hu14FHBOCTGiEUAuwUlKNhFVCVWb8vc
A9a4B/gmWqgU15zXTKR+yAw3Ibx11PfO6ni9nxQLi5YI2kKqDpa+e/GOgvm+F+En
feHxQk3i5HV2gxHjU1k2nxo24k8iRFNqjOOsA3g5KG87aBEGBYOnfo8tNfREXfnM
7B5Ac0tN8oYjdnF56ZG+bjnygZOH9JDPiHGhOjCc9j2aWguRcR0NRrUTL9ZIf/jj
cCSBXIyYxX7OeU0ndhTQfZtnkjPm+kZx2YM82VvqKRoZ0zTE6jIxWnK1NrsKte6P
m2UFDla+9r8jZB6LKHNRtGxmSk/VS4wo+jJsL8gdXx8XF+8+4AjZY9hIJankU9cQ
nnbHsG3a435f0/jNpAb9zQSpcbaHc5O+rQK6efbD+X6Y+vPedzin0KP8Ph6mfLIa
dtYu/Bxeqkr69T64s3DFFnhLGAC/HxZnSBG2vi/tdYP2FEqQg/SapvdoqM/xCF82
5lKRAMiuxvqlZegyiNPRDsaENcEArxPODYUtFMZiUpHizlHMn1lSK/Vsz75pxFJ9
kleom4g9QjmID/STripG67mOwUqq1r+1lp+H509UoASZt+nfT5AW7Xo+/W+IusJS
xFCEg2zku+Gk4c9uV5/tyTAXE+1jgNEeq6aMUnutXSHeCZtnrkZUxnGpcGgU+XxB
4PdFyumus7IL2pdGqsmqzxUd3aXoNN3XQMSK7+5bjscVkXgPE3zZhjue/VtOCTy0
fcNZfgop/3V7e/ea5S4ZWikBtnFDkq8pahMpOJj4WaFItr2tLxgElwqbreGEEYic
qdveAP7RScFuhqxFqP31rvgpKmfI0xN/X1fIvANsEp9JgqUwaZsLKYw0djJmUhPk
7t6jQ8FUzeEDiAgYFgzk/LeAa3ZVu5oPPnSRYA9At2C6eKKD/y2FbzIIZIdJdCYQ
LNZqcuS390jwbqYVLREUBWfi0BoTmHVgCtWosmEP4Mdw2cZqcrfjEVdx+o9oNMbT
qnmQqFcJ5Mx/r6JBP2RcOApcH/9yUu+QfD4qzLEDs0OCOA1aara4qy98Gw22wUPt
KXmcODOCav1gQmhQqYsKdUg6QUbHWLbZUxCGX73NF76wF9A0kntLJ+Wj4X+CKbBa
Bcr8IDaTKhbsmhCBLNPT2WJoFOgOZ16RxRX1LVL60WpiT1T30lUWVkzwZh7QHdiY
plLmJN8Ql+FtM13hu1s6jHKQN9Ui36cEPKQmq+PxVba+Pl3dw5awl5HFR4wJKjtf
HGaa+48M+0JSaYAzx9LSL6p2q8zHkkm/J6p/OfL17wu8XP1RVHZPg0dZjEdAqkii
Mt1dqDLyrbEerYbK/7CKridhFXf558BUbA5RqKZ3pBCBxdks7SnrndZTx6swpt/1
c6lBZIz164aPnAKbLDY+KfM43+G8S/oh6xeU5b4EKfNwrnLV68IHgjPCgN4adWDQ
aABBKc7/cr2uTvBnlBAWLem/li5jo91qQgGmbctBrSkkcy96pItHdkZEIYFmLOvY
p2vEZ7Oid2R15ySK3YI+8MZ1XLzV4ZUok0nLw8hWUBMPa4izMSvYppFAl0CUGB+w
mPvvZ3RM0f4eFy9PO8RZLfhBZog+h+RVlYCbCIqBFcRWlLxs/BKr9OYotIEkEYWY
qMvamUmJGH3BpC9R9JdFn4d3kaAh4Y2msJvpRkwR7tG6duMpDQp9/MLS0LNEs1ON
EbFlRz/+Xc0xUiWf5+HYZXAUIlh6PiCbwfkdoCo64k1YXsOjQBuVCj3j9F3H+CGn
Ate2nPV8MBp307QvIgQn+K2J/5FZjpzoERrnM0vJACWA+FdDGupR5TMTMF6LFKQ+
2pA2AoiK6C2TzyVTWypu7gCcFbj1ABlTK6eXndkGWOejP5tsbqq/wiWHKRt2dGJF
9AQC74FJW4HOwuZgQPYf0RLO7fLlxbLIAztaFPcoEHMqVVSoyN+FYq1xsK8bc36a
JoDjsPAjsGqSLChDJzWlGi8rFbXrXjf0NErXYZJRjJVAajFnTVK3t2wO6jSyKpXY
DziWWpxZuZBPgBha9GCkns9eFRr+rOcB3CK4QzEDwEmem5kCNKTg8QXAcG1J69DV
j6nBXh1D6aVkf1X74JyYYWYiMxPSMl2PhBwdYAkJ9j/uugqiqvc308KbRPhMCz+t
a/lKz3ePelWPv730QYNwCWFmKeMQiCO5UZTwtYzpO31++bMkSl0ETAv9k7q41Hk9
3FqgEtWg+Lzs4KehkgJnoY79r+MJEoQ9H01Q9jL7bdtOfaSVR+hHsqqvql/EWlVx
n9yzmz/znrc76gcDSiU2+9pjovmagtlJCpM69sz1L5Ydv6fu4d2LOl3D0h5x+Sq0
Q48CKg/2HjMZuOVgvuTnNdGhMzvHex4Jj/L5w3n60vBDT+ZZaKbz3eU8osyU9Tp8
N33tO8bMAAqGntvjRTmlyix0IJFDl+5WHFMv6uSEySnjAJZCYNcGBvJ2Em/OEB3e
DbTR+2Fx1Du33bZGlP506gfHcrCeyxEBr+1hro/+zX7E0BVWpYIFs/9R0xSQdo/O
SSuLpKk4c38eQv2nwug/9gI+DrYcGX5VYO+JR/s6aLzacb11q8vgLHMT0lFQ+vsr
9AXHVd9s510TF7jwLGP44blOzkBo44Y8DyDkwjIRsoK7cTNEO8fVWmVl2t67ljW1
/gvnDvJDpq13NxcW2ix1SnJNW1YXJkr0IlLpV9/J32Q6NU4FKd8vpZrt6CZYvXl3
zDvDtxW7df6zwPMqDlhg8Jr7M4DZTFf0+8Xa9/Ek42hM7WTuAaDVkaeKgKtZyfXx
MWeACFS4+zowVPg3ozri43TlaHNt+XTLnXiZXLUQtX5ufl/55m1ITsD7/21IVL7B
oJlE7tR3A/o6zp/uZF0rX/p+L/3vNEZi6goBcLvWP3apGFWNvfz/YGyyUT3ItVU1
SR27eYFbkPTGyVShRpUc0S0r6XuOjyKDoJPGfW0W3/7yiJ/boy8vI5KO6esZ06nN
uaaKqXpE3FzxJiaijcM3DhECQvK+b+6s7EoMissvwSmEh71BpmtG9fLH/4HXqJ9p
rqizqWznzS9QmsYRRh9o0/yaDSKXHyh/yrkDm8oO9tTOPt7Wjptf7xsG6IOSXjEk
JgUM6ifrFYsBv5BwfopCX+PB1x6KWnWjP+ZjOmyRvAcS6DfeUr5QY4xbRNLgJ1MO
wQAdhqXUCFlbRki5Iw+FQvSipNCNTiCfHdKR7cfwzxgyzwRZFxBun3h6zKnDvPc0
sugZ1b5XBZAR2wtz1rlZFbBaoCgH8PmRhlSeffRQVqDIEoXv/qZN+qioOpsjr+Yp
k4z9P8poV6KmEUP9VFJFhh0kQYDWkOCYxXCHpMj2/96HC8HXO30CNh8ADjAB1/Z1
QEpVGckigQA5ADiBuK2YHQhMcHiA5+iG2IEYD4qqiI7gAFXkbEdNQ4aIYmAUaLkP
OBz0bhCxDDKYZldrzyGRnlTlPFUDjOo4M9WycOO7in59jseYVvCAI6ClkPmgX5Ja
lck0JvXX/ibopL+9om0AYvSyjCHqYJIM94ZcQ8DHGDdwNIihZtwA4IDkg+Tre5hv
hsY4ltgxpSEII5bgH3I4Y98zN/WT8bs5F+ktut5IlAT0/CBK9s1n4JB5DATKCFxk
1IPAuOxnx+6eEIHmUcsw782w96xvKGceWYN/2K8aPteyEPLV4yhWEMo3LvfDdve/
84iPM6gkzKeae/0APFP/y+kSupLxDMmMcHY1AuFYN4hGF5RYFWgCDXJSVe30gKRx
KNvgJqnhp8qgLpcoMXF5wlc/gueA0lZpUxS4QTzeYPLcAta4BG5N9Ijny9SneffJ
UU6PLxooctWrAbSUmZtzt9RZy2KWaiR4HpSRMrjI+lrgL5yThdAYgok14eiZoN1w
qaQdyGVdvbfnVl3OY0otSE1E1RpcGqUvngZO5XmYhTN0JfFaSIhNrAsR2RBqT7F0
vPGD1CXlFhnkHSe14fXOqY0xjy+jnXUYYGEBR+5puBfabaJYQPFmWv8qwf3L5umU
c2sZ3Er8hQz4JJ16fwPsAgE+F0LXdXTHXbbpncmjLDY03gIePwY/MhmeSPb/WtqS
4mi0wRAtxjp5VM263fIh8POWDPSn+12mBC6trVDtgZGEXTkeB5xne0bXlGCFGLJy
ZzmxXH1nYRHk3PwnI3f/wM+o9DiJA95EKHbc2twixjljOvTk+ymfHrz57T5nZY1m
eDW7acEtFNwe135jMrmABSB8NR+vyFonuguQjpgQAKH70TPyJgg7JlZYwIB0sVGh
Y4F3N+xhhKLI0srx9+nJZIGvYKK0Bq68Sti6+TGMl8Uq+0AeO1AyUf3mgb8dhObl
yfHgcvTYoLYJq/tozd1IOecW+1W0I2mQt3gY+poONfhJx8MnuySyS7N3EA0r/gFy
23gwmB/37zw86Ji36oI1nNV4nPU8Web34OWhKkeztzm5QA1TsZqJDTprRI5anhgN
0lHoIQcjl5KyCWmGwG1lB/i3TI3PvqdDjj81VBVnxTUvrKNxPmAvWH+Ga/vYdHC7
Uroq4jeEcxdVFEpuCpmXiUPEPePlGy9RTU69deunf8dAhmHh2eDcIiMp1Z1gNdk3
SYLbr3OyHAh9Df6oQHQVIOwPkB6NZ0CyrnJJ1AQ9sGKGkzKS3c+aLMFfGB1P+t38
/Ge8qeN14Fb/gwnV/2OYD1Yq/TaC1zWvHpxslsoNcHam6rgKPxmcP5mjzc6oiQ5f
iw/yUCesVFYTLiusSsTPtSXdPEbCZYBRgOMpj+A1s747TUZCuPvW16c0zS7kMWEJ
My/KVRPnynRcLlvb8qsMyIHtah6brzSo2UO0Qz+RD3ZY87A2fGasUXLEwcQ4UBet
nVroWL9PpopQkhN4cb9a+6pR+dYWoZXT/w9CczTprbHeKRs+TpQJBwA9esCWHQdZ
AV+SwjqK81nWbQND2XBw9OQfG3gqpydvHFlh7LiBZ9G5jjFZ/MxNDPJVcGPRW40b
7tySmxwFU+44plaVLN9MgmLys6iG6S4e4nZ20hIZPmggo8TKyLLW4dFfPVFfr4zV
hFvunGT+Z1g+SSvM7mZ2Hv7EEn7pD3wOOgYNWJTNUL1BUSdjBwSTtg5alWIm05Jm
3erb5p7AzO6vJK+2PizvVXh/4DGGinoGjx0dfl6iyd8Cz123zGsffMyfKRGWMvab
Nri4kii9z1Mot5N0iA8ex0b6ND7POm1WhJpoHSU55PiGVrPFkUhBsBgLcQs6m7Rx
C1Q6RI4CmJ06eW4jGyeeYTkDuPHuFXd9RcCjrciAPRN7uTR5ErD+hkFHWfm6TrFq
i5ySLvyeQX7I30KvB/uztITQClqlqwj5liiIOw+uNnRFo6oJtcdYgZ6rAQCoWgOr
8eWzwk5TZwfPxHqv+5TwtfQoKbYd7HuBeJ04wWzVACah6tRh3/4uPkuym3Lk5UCn
uSrNN43jSdmyZohPJImPJxNFdSgYmO/2xClprUXQPhjKG8PVR6ZaslL7zQjZ9xlB
I48bG5kM2N97PQSie88tXYX5OfNcx7Z+H3uZGb/RnWFEqJ/bVLKbwWNgCdqGJm5s
sD/tWE40DT6u+iz+SE1qFTYTdmh0j/hvkYRwHB6tpvkWkMntI1pSUUyzYXDyk1Ge
gWpsIG2yj9hS7ZIBRH7M1RKQeJW5hXWcNfBUiSdeHdsNo/lr4mC6FBNyGMlpNotM
UXjxkL7lJXXNg6LlIWkYL79RzJ6G0bmM6pmCyijat7UsAy3gN4J9tmQJs5bNoz5Y
Zbh7HOW3/QQDgbeLzGiD54q41Ci4eNSXZD3jFS/ECzY/WUi5TbEpnmqq83TJiGQp
BFsfxLKUB4OAVPm4lcp42trPFwkUH/HfbrEVCGoOcnraDhuJLbTQs/rG9Ruj0ONV
w/3M34/NebQrbHnTU0EASLGjAcXPd7SghnoURHxUh06zYpw/1qbFgYGeqbA06lxv
I9HfZVqnawLxulVzOLoOHgII7S2QuCZUYxQEgfnVqR7nD6wC1TA978zIua02uz0K
/++a8/e9CaccTtC7sKgetfnvlb3xqFoe5kIkj6E52mMqHivmmI8L3obRfeJCrsCQ
UNiBWvMhlseia36NeutIZl6b7+5JXcsqkir+MZTKzEYVBYepcuW0Do1vzgSAb9i8
okYGt5FkrwTAA61x5Bl5xlgnVH4qsGykoX4InaBgTpnG5zcHyhR6kYxpg+b9ILD/
yIURZwpSe6yJSUws3b/L1IfcIjQzmfKwWnWJ5KlRie6jAev+Ywi2VL+4jp2lF21t
0VbqgdW3Z5JqTJQ3+2gnXR1YHPmXBlktu5/1x1L/Nagu0kGtGhJyWoRVYv+V59O1
nrLGIpx3HXl2mLg+nLPkRZyDA6rHksxQhpOEy7vz6J2XBpEfZm7xnV0HHqrWOOM6
8L/DRS8CeIlyMJQqFH5dEmc2nJQs9Nob98gFrJrXkL2iLa7MUb1e6tAAEsCmufTl
Ap6B3deva6D7Ij5P2xAExGUkqNF/2vkCoWBoKRySYMUX7Mrpnx6wiLZIhTokuS7Q
o1jVLMl8fDzZjroRHyxvX+2bgfMh1lyhIsGS+sxAPukbuS+NGWAqKTOAKy4qgwR+
g2vVbOjrQWZnkyNU3vp9aNrZmWrn+WzNnJHGfl+RtxN+mvpAW0g5AZtwJfy6r8SL
MuHYf84sxCIP8dKUZvIlJVBrYEAj6spUsI2EBmStyISrGP5zXK3PaPsPsDJf2AEW
gYd1bKAjc+Dt+7RIke9UZPDa+VPWey30wx8nQIs4bCZj48f5uzVI5465pspZnLMx
/2prsN6HG1PVThhlqGiqoor+1vrBlW+UiW/DRt7Nq7bPWrJ3E2N6T4+d5bFaBjtc
SF44x3i06suMcIOW9TyJoRcf/zbXDaH/23TIwDQ/ezln/cdBh0gnRPzni5MJ+Ra8
8KTHP+dU859eD85QcRHgbD/6e4vbFVKaTVKVxY2Sn74LFmnq5QusJgztS09wruMT
mMMgoEgqu9X5fuM2cENOVZD3/lNyKr2GARN5JQh2thrRx7gT+eY6fsTxRx6RCTU6
tMakhM76zG/nWZ/dKlYLZSyoCJNC0fifuVkh6RsCuVr7uTKDUg7UDVOGYCGyDImO
zMd2yvOy0j+4xGDqEQNryJtwFYX3vltvIRPB7jmtiUk5AOpk1VYOwldlOPDWHtjI
q7hlt9H4cOE9EPsPLi3AaNLN5gNKwV6K4Mm+o8X4kdWEwt4frWbMQAgxRESH3c3q
siWAGWXzmOvYHjq7E2ZbEAaIhPWwnlHHUEebzEet8xboVoy2FDfwrG5PasJmKbJ7
kcbF5E10r/tQY2+i9VNL/Kd0CgJ9rKvlkWkvHRuzn0+xNeZvKEc3xFfRHPX5YeQP
0itOwQIkJGhsGKHLXjc1alFm8Y75y1W6AGBNsbXv3GQnGoEDikSxzM8ZZKHPVeWj
B1NtlzsOWIP7H8qRLoJfJ/h5wlArnx8DFIwSHAM3UmhZcTaRMaqCTc/SI5m8adRw
GakdEdx9tvO+pD/MoGDsjSzUV0O2k0Fj/9JdZYca/1cH5omZlR6Tikx4B6ZWRHKR
RfMYDx/WH/FDlSPK20dC0S8su8XV1NhUFgH9y6WVddL0BrhKzWRFtJ+KUwXAdBXL
tM03mWzf6mSdrwLfhOkwYaTx9srKdfEoefJDUVIQgXmtx96fJqk2iqQ5TcmiRI5c
jr5Zef6XqcUgPVOt7R3UVb/6QCdz5oxUnEHiJKcAi8EuHIsQEK3nbyMKU34NRDrw
/QAEUfNi3VYd6Y2LoMmX3q2f5tN6xNkJIQwVPNTATQ5DWUTj14LsaGWR0S57UJUd
hK9iNfSTRFZgCAX5ZOo0oyBkvy6TdmzGJCCkzPx9cD78BETzAvWbmSKgntHe/AdN
BzmW4bA8ftHmNPx4XDqWO280JsOG6b24sUZrEFMduWX09addhs44d1FV4aV4Efgy
fXOe4PK2ir+cbGXY4pdLQkilnVXq307LHXBMY5Y5w+da5FJVTv18J8ALyV5AlfVY
WKokwKNcdZTU23Akf1+pnpYzqZ0U3RT9nJmEWZs2HWuvtPbwXhS7Z5aaTWocEuv6
shg80CmCtVBlOzQBqC5zvQOabqzAVGYhB/OiqBbwQmpLRy5+IUDj6i76qUxP8uAr
jG+T9obLij2rKvvZa7AwKURSKuJ6QwOJ5ReNjCpG+vXWh+egDUVjmDbIFcHFylFA
0nDksN00bEA3qMcizM3cJDyVmElhoRd9dfDC/EtLzn5kpki+BCKjI9Titjj237A3
rrCdrLegs561selzH5qOXh8u2Oqiih3XHE2EFLVoulzdmrovACc932VATqqPiTYY
h4UbHe35CyRBcfe6Yhz92WyLhhOWAXyLn5YkuEsKkjNUxcHS2A0vW7w3JqkZrwot
htigN6zq5m0cXpfNmNmCufL/yCftMUDZv7eZdlyEHNjgsTHeFCL62OJ06SMGE0R7
AfzOnWGbb8gUY87k7IFTutF1jgQbazepUIOpmbw74Zj+9Caasbo9jG8AYnZphTW+
aPU2ZEIuIKw/X009ieZMfc96dW5qqO6mGBMKg/aDmguXjzdz4qsEbDAwxPW10PUr
pcdqHGdfVKVqqbI8T91oJFfrXscHH97LzkYNWTwm/1bgJcHeIe/4zQ65RbJDBZx8
hCpRqkKVoDSotXtCrHWj6Y9fJNG1VgSRgExUOeyKLwBuW97BGZXEEh74qwLmSEzZ
cujiDNjqFMvIcu1DicbbDo0fnG0rB55k+SFdJvw1sytmqpA/4QMb3dwA9DlaBYvq
+nZNq/JPSr32yr/Bwwd925Qz290Q96lAE+4z+Jsbz/d9sraBJrgxlAEtdA6LQabS
5vSzKvJZmBI9D/Nsb/r/X2oM6PnASUdAYxitPU3k4PxX5MbqTUoGedAgTCMYjOpk
/CLZ7nbly2XZSv8k10NKCKT3iyB+eiNQupi0Ieytdh5klgzPQcptp2JYYb7uUTNd
YDS5UrCs+Lcj+FoZAUUMPCwildm0z7Wo0ckUR547FHmFDAA1aVxVt69a78GI5fKE
GHvVAq/ZcTexXJfH2kK3vYCSqt+5+hOdqba6sr1+FRlnV4OqnvBLH7TcXv2WyoR7
C4fb7W7ZcIDH5nxtXe1FY8Ww71kLLUXcvp0kgIQUJ9UMVzga9SpFTQyZV7j5khRv
3cQ4kzvtVf1uIF2KfYA7h6th0xCJM+yRnWICmnL5lKSygfIJMBkfP18BhNs6Ax70
gZ+hr0fWR8MH0dYBZAKJmAzPo4qxQiW5w7ZtGYD8Cs3ZmDnZNfHj3p7ZTTDoml67
7U7ZdEZzShh2KXLt2nay3zqvjjXJIoVlHWBRh4GQU4Avpc+Z/mVa6/iQXoUpzI3q
Ee1jCkyM3YLMwnXcwpEvDLwWrYpHKSG05TTwcOt9aUkLlWKv4kZA+6TUnOEehBbJ
F8B5vbjLWFMLWx2Lrj7OWGw723AU3cuDG2juKL+OwAxWr5zGyrEBA2zZYw5KT9vo
4lVcBgt6qc5cn87OPOj3HGNOJ1CINsBzK5HdNwRJl/tmJL55C4THIF9a4rb9z1TE
ltZ8SI3T/rnDTYpqPCoXYtUi6gpSG24jyS33JlzCrSTqp05GzhXZEv92OHetczEG
aQsOHT+wzIk47HooU2E0FNyKzd1Q/Ea1MSQa800J7CcpxVSO0+SMi2JKo4GUPrtV
qjpLB8Ooo0diQ3OHPQSRFdCXuNe9bGe8R7iAFj0QtQFaRhYjIHVLpv6UmiuAi03h
EJukrwsUALWcayiZ3zzrzbWkHMskqU8HEi9mFSAN39cfgUx0JTXvSwEE7ks9QXOe
4+NrfHh95G3uOpV64Fjdyu1A+DVs95lMfrKJ54LW88J74+Lpg+JLMzT1A3XZpkba
7QI37BwcGRfKqW8gS7nPU19ntAkjTM3j/HIKx2CWfujANcYqJEyjCOPafBOCjd7p
hSZz/mquP/MLd43CIXBzt70dWQfL+judmgnZUtVtrDpMDJEVeblW6jhm9BVr3ZX8
7E0bHnHuWHQpvyZ+To4ZUx/7UxAkwZLPmkBYBBxAE8Zt6t81HRJPI2ZSQAZRH2eL
2iAc9wCLwS4uhqTa5yxURt7UJQ1Vryn1c5C343LdNMP4zCHj/HLBeUkyVVwcGMvF
8EJXyBT5vOzVS/PycPH8xkGcUIEtSrntYBlMOS7yuRczkRPKqe2iuK3JhEhRRn3k
O17qIwwNhfMg+L7nMI1tdzL7wqSgxtIqMmdJsJSO4grPs46FlYTKchpqtbrED9Rg
RrHS6YD/Nae3A3c7csXAA5h2eiIhjAswVsvtHu+ZNEJd/hDQVr1hCfFLq0YLVpk1
kq8sqqU9AH98rnWaqK3RQcbZFmHoYqsSiTngqVcc8QG9h/Pej1R5hrMH14iPBv4l
juILaJpeXstl9p2S7VCWh/X2XZx074X0h1JeRr0iOYQPe0qHvDYUUPy0tf7IArdJ
5O80vGE7n7g57jmidMZUVwp7/GqRzjqMfZR01qFICVM7BXozA8xJMmATfZAgb1Z1
0S8X+qvS0PAp3FcPoy1NeU8c1CBcQAycvrYKLj4fnSd2Z1Aky4RIQgsRnKLXNuty
ZezmYgrNFfFn9ZvJ7kprSTOPF1OMUWIOhimcqo2XlmG4u/r4k/8BdnQhVoqb83iG
0UtDey0MUmNxlvTtFoZmh7KJ+wAmpMprhqgMkeOGVTxjQcK/jdh390HGttI2lpsh
jxmcLDExJTHUHlkATa+0WxXkXtkv3KPF1Mj42Pv+oqX9/+03jUm+IvE1Ba9DJtHV
qD505TcIUQlqA7kHo+UfFitSQ8mFe9KxOEBRGqOc61nk4xtpyFwl9/w/UifPkyHu
sQFP9/hCHQprNchVclMIKl2rpOaT/D7pkk0Fyrrw17JrqTJRLLWtzXLrY7aoj9EN
zIvTbstNYUtf+7ykIFVzb20+6iLM3z2XxzWHC3nNYvUUHc6VpQCOhWIbLkEH+IMP
TLvYg2LdoSFY3QGI/1oriR03SzXw/uZXkiwBvmHE+gL0+iejr+9iWhjxPeCYGx/+
IFTFSZyLK2/Pmzq5AJQvcD68P9FvdtRC8fKUG+VKLGdnC0evlIyPm8rswfoVBHHC
+H8l3spTqy/ZkWQl7lWUCRJuevlpqZfWKV+TUIOuWlOnUvRh50Jaw3Nd3eWqITN1
z7Cnvnzh4o1Bi7kl7sZ43mMfCx1TZJSf/34YAdRWiQIoGnMCuBDOphWOi9xSWwrD
/nSE7vxaeIq1QlZ1mU6skVQjosQrEkaIC9gaTRUuyUn46WbXm7oVlk2ajkL63KWi
yIenJhhjIi72ZNOu9MMaEu2sogNJecjqGDJF5WN60KRdtvmYXksBJnDmq3Xk/M2J
qgWSIIAmzV+ESxc+W42vx6ezZ/jHhUSOKgHPWbmVHRSeH3ks0wU3mtTm1xWOMvv7
qF/6CSMt6W88Ee+E/P4wqwbwz1LlrSUUzxaECKOJYK7ywlPajEYAB5csyYA8YoCL
/5x20jm+lJriBOETMtofxMc4W7r+MCHCrQFx1DZ071jzEiiFs2YMfpgvuG7Bu1QV
AIB5/HItylb8Ya+AWATt9jI5vdyrjFcR1fKzwFHOZCsyJhxMxJComvmKgyR5hzPS
u19xoRqLXIuI7nUj0JjsNG93nv76u2f97nRTfD21xfQbgPrKuQotnwiOMoNMmkK8
0dEaPQZUlfE+Veba6sgCdvFAcP9g/ahBqWelaA2tbyCrTIFjzvTmtkb7yhSZis3L
ju7VP00bfIZLsCS2YqV8EkEPQPs6mAgCNl5HOkhHjzzKFzCiSvkJOWb41ZHQYNX+
a6dJLGT1sKRwKwejz2ik+Rr4d9KVdbHor1USL9pb5UikNDA+PhzGFxFOtke6OB0j
atF8OziJ6ISgvGZlQb8yXkc5+0bHg1uFxs0BpsomfhAy6SszX9xiCnMUH5AW9uOO
n5j7GVJjcKEytEgHcKvdTi7sDUBPFLlMHTapCnjswSFmtSOt7CarAwzvHuby0r6G
7JED0v10T4eE/1dwss3kLW1OFegvzEVpX0jpSLM3SsPiYmFI072zTciyuASL+gwF
IzbbOt3bxGZMV7ir/7ItFdH/EzfSXGPE5rl67eSsjYGJF6EHEjYNIZCxAwWj/lyB
WybfBniByHKZy0xNaeV9DeIJi9Y9PE3p21Hn4+ahXE8PEwIwpKIH3/2E9OGzrr9v
vupAWBjCC9UJ3UJv0tcS2WmR/AmL8dJhC0QipeDZpgje5zosphKMYnHukVbJyYhf
eUsDLJHJOcgY/Rv1TYdSyWFDXqbQ0zxLUjVY14qqIumpSWieT/tY1xasLPGFdSqn
f1lLh50gJ+H4tjSflvC0AglXP3Tr9iheNN/vRhTG5BHhvmP1qbX95Z6eewLW1n+D
KKUxQAw8AZe14vw/a46eGBsF+n+hlEpjQMs94d0/A0j2Zg+Bg+s389/9Oue+b9Oi
5qBAMJOzzR40J4qvg62M+86y06gdJ5jJz99vuzjpMoWlP0LvY2wVUwlk/+mKcHHj
+ILv7EDkpq+7EgXIOZLb/aN0y1Px4hfxaTB+wKsdGnBSuP1gelJMSH7gSv7YZVTP
xA4WjyEaCZcruINDZAqGzNCutNn1TT35gU+zEDrotQ1U5jUgpl8g5bvXIiICayrt
vSgcLS5eQzwG7uIlbWn2bj0FynnZAPjLEPUpTD4wsQS4HlZDGzXSxYCwiiDHy8fO
ILbRavieoCpXKWiBWIvnHV+DJ/M0JPirHhJAKRohNPzIVMmacwc+OuvnFd8Os9k0
HMtkAwR0Y/3fPNWcgMB6f2052WFlWTJoIo2r9v3/LnbX/yDwXuENyoVsOf/QOYA6
1YsUg+wZCS+mR5qFyaiXgFOOCJdMtNVJvmivcamFuMv92E6oeoEnxW2o+D5BSELj
ZI4wq0/h37qAsdMW3MHDZMF4Heh+nj1M00dqE5hsL2Bq+Eqb4Eq+DG8wozPATalg
ziTjF6rOHewNf2NTbBMzPQ1NZEM685zU69nlz8S32yxQQJNV8Tyz9M8f5n+Zxtmb
teXYEszj4V01jd8jOVgFPCbyprnbvy0y3HE6sdZzS/QXOZ6oaN7ef1wu8h8hUH8q
EKyjbn4Af4F7MCdwLVugwQgpkCHcEu5/nGe2jeRumQXmrHtDli4k/WZwyzJW8Zhm
5h3D+fENyx6JIGiuk4fAaRHeWluvOMrM2pqFWOAnlQ3q0EwTVl95i36HzxAFZtsg
Yd4Ga8mMYSNU8olbEW5YKU4pH/B8pwRLYDhgnZWWb/ZAg/kDePAJhBJLXA9ohRCl
KPyeg4TTYjBgb5dMwmRM2gmJvWxViFDbv3nJMOOkiR9OZGF88JdUN6B+R7OwYjQy
3GVHLx6NBQZAKkaYv60T1ekZ4xQfRXyu/KlayrQA+HoXp9atcelwRonyz49OJCvK
ot6UFGfHgI54L6xYoxP/fAN5Fpbh4XIAGzPD4r8XjBxxHU4fUN8Ipw5JvmEypCXc
KBaw1H+cw+vzst1K8U2PO2yMPffbMw9HvNl4fnknwuQrdJYAXWmmy8F92uP6oSYr
OW25ZQNpqcMc7gzYX8KSBqRMU4VtR5u6u4OhmkVAAPM6D0MtfYb1gzSELEUUWg/+
SR7+sS3ymYIn/6HqHo0jHwFuw10xmOr+0BCdm+5vxNTqko910Y/greKR6STg/bL8
HSDJinl4GfX3vUurT8oPoOeZW6RA+ztDBm44/4O69FwUULKSGWnf8uW7BLTjKeLX
btGSOivs398Eog8pd4XaktyxwSV9IiP0i/uaUU8sZr6izfoRrdS/ssmn78RZfFFs
0a0MY225C6Zj9UEkyPjx69qkDyrnAv9HGsZrw9GPpIaT4AGN4vVHzlAL6zy2jKSX
+zl6YOFze8OnCBpEJj4rDJFUD2FHeAN4IRVQIx6FDao3np+Wgjt13s1KEp8RMHxb
scKx+7I1AxcQtUP6oNfr6S3Yhzvv287kNHzYo67PsFONeu1LAHOAf4cxcTem5SLA
8Ii5W/gUv4KFTcbFVX+n/8EgheQZ407+K1CVbGB94Z1kfbHY+Ko65Qv1vcsY/dFN
2cSmQsJCTJtnK0BU924++hEl6P4SqMIVTu6be4xo9LD5KfjMvpNk6pdb8vNDFA5x
1k0s+FIr8g2UTi0v1uVjMyln7fpWuSfET/NY30CP+CUw+PvdKlUUldVStblrtHAM
Fi0+99qM8JTmI/dPZKoAn9tpeKE0IO+UifPhKULhHAu50R1Rh20QKJKOsjwQv3o1
PxvitWsssOefnzrRtKmWMYqU44Xgm5bmHAwUfqd9wR5mDI11q1Ia7eS08oUbEbyt
hsVjdFK87dGMCRme/ns/K5r48neGpPHxNCtwq0ptnFfucQsZkBemQiRCawVRqv8I
UWTQ3GVXTRK3CXffnmYH/XK6yxToO3Wk2CjngEvqIwpRhoNhgFMHkBDAf1MHAH3p
2TbfigtTxWQ+DNB+Q6cFwvv3Vv44zaV4BllrR/J5aLXGV3cD8EYmjRN6PgsXpmUE
w1WCa3N31W5YlFoFh0UIcXstM2uc5br+jcKnNPpQ9mU6bSDd12y+EIQ38fp/jHZG
u7eN4e1QecYS5AxGn0T97c3jbd018JhnroJ+tf7f1B/EGussnqTE6LRXOiIELMCV
piaHTJ+eXSDEZ39QAvrv5ARcB8igLN51f0PahA3AATyM4R2uu2kk3fP4r8FruD13
Z+9QRnjdoPEcOzeYvhp6P14Nk1/nJkdQtFD8ApU8WYj2m+C17zFrMjnsxXex+4fY
5hkHnk3BXsA0PkcD4B4Di931oNQH37LAlJqsttIUzj0ttCJKKVBIVP2XN2sWHmKl
iHUvTYM4FNno10XY0ak/3QsDWkkHZTb/IGDgSmLgDcm8jwmszO73VnnYWPTm8bHK
s/3NsYQB85UThq3IFItID+P1kC3PT5LSfN4Lb8Ub8cmyRSD2jUMsgN46OhazoDvE
5RmyBAzn0dQXe8zpF5TLQawDPr7H9q3enTaMX0sxxGN2sBzsFauKl6jZWQ9wyo/1
lmYT5XUpesxIh6uQeZQ9bDvk5Yr+bkyioDSeQo/gY4s2QKwLmT/IlkvHSrGpOFmF
G1OUkuAoEJojK0T5k7RkGH0m+/IyvP1i9/4Mfi6gK3Igk+QoV+c7Dl9hMU4xCTe4
YvN15IYUQcvXtj8GNUXB4X/o6c+A8gE31py+PoK2JTF9t84DtonBb2N1WDkRV5IE
KezFCras8UE8wC6YDLa69E1bLCoX5NLNG2QRxvVQEQTz3rspcH8VFhT5nbc0NH0r
YxBk0f/4ntMXFVqFln2KOHZcsXbf0nKjPzD0UDqyeBEt9tfvEGQ41Msa2KO6bxyj
v5sQqXEA0ZqI8TVfpzmUmb/+BOEtHrIwvmZqsc5yHdmuxqhiQ4cuquwR5QWlFw9S
GynMi7Fzc4usqgIM3cu4vwwMgzenSw9ROka6D5h25CACZWa2udp+y45lrywJbSHz
SSfej4MBpm/9d7fvKJmr8VjHZ9Rgv4mBVa6mJrzavYfPhy1JeaGOdTqLhRw+Jqg4
l2i2L/2HXkF3JvTEBCYTsXdN9VW5KOSEmGIbt4luOdj0YFoQkfXg//pqBodeFCv1
nqRpFdYcWh4M/QZMsKldWDITGvveHub95ayRlDan6F0FxPunfpzd9+/w9+v0sGk5
xv4CHuP0fg49fk/MqZ4jP/Vs0inomiahX5IVsBVXbZBl3mwUsFbRudcv/7XuEw5/
mOobJoGhO1M5jF9Iwhe1J3OJZqg9moaiHXD1IT6swN4ytYDwnRZvnb1KQG5YrFmE
lOZpEwzz5hoXw+ycAsNDh510YB8+Cj0jb+5SOVBPi33Lp7u7MYCXUC4C/8DxVhzl
og5w27W0mHAbFxwzJR95G79u7J7TktfMEDkkaIHvv0JO0+RyFVJ2bog+bMfezP26
WDYGX6A1PfEiXRvm0PBPqvKMzS+4HNIawagFHhJoL8+H83d7eHgRWP5mDNF0gqhJ
r7SzkVxOMI3Oiluff4ClUJuaKz4bfodrDo5ERvLF3LporqH8nOV678Ys+afdX3ZJ
QvcfdLF8Adz4GEvuMPTRc7nkBHIPbYzeH8eU4i5uKcRf/aACdlck/0SO1RBK2YRp
k3GV1dmqTzAmUfnyxHWPGGCYXH6C47ZRcX/1rhM9ZOHEx7ArVD9F0jfIL7iPCj2u
umryYmfsYlu5B0t349zQRONBFgV97EaRMq4UZQ3zi73fBTf7IVky/2Y5IZl3tDys
AHQ+iih6u4WunCJm4NJINuEP/IXrNhjQI7++87XyA0FqGh8L+ppyYCGyDmXsQmzw
3QJyJbk/1WZdcWMqJ0ZEPgmPcKpedwFgfGQgYAWEyl2c/M0W1gHzw0fr/6doSy4r
p2ovzEidcUUpz/AvoA3N5Sdziiar1WuoFptZLOl4xWrYNT4KxhafcXklGoLILLY4
RQZPNSwGvMvO3xDs+PoNdMnMPY92OEjPJaZN4jxIwDgM+q+46yl2yO+iiasoy83T
kUdUeGINm14NoU2i6Bks7d07In7qF6+7wiSECfYaHZ0SRIglXQtyD94Os95sWyrc
79DPbA6oKymKX595Qv+27H94ZaflFuXThyF1xHpI/HGxjnWlpa7ASztci4Y0Le07
cQJsvkAAeYl6nI9HmZNCnLzuisXjtKHBqmiAAB1g63qQaS90fqazwZGvAxcAj1mk
1DbDSj54T6z9MvBYLo9QNkZm45rrJuQnnJs1fkTkTuKWWAYgKn8jiWYm4Fhbm9YC
xg59m+sccfb0At/T12nY/CxYWYzr0yS+TZTIoCVpQbQPDAnf8roRO6AL2ExEUxpC
H+xFjVAWXa8+CJKB0tUTHWdwmCYu6B//fN9z/97hHVQhOh5MyZ9xX/W4kjcHrr4y
sczXf2Ik2lBHsVBRsabZ08Z0ThmCF/bY3z/psUf84AeuftswSeF9VAgV2R4nFHHt
mhX4SPn3MxfTZ5UljJ3AUqrD9gphQ9p2YbwzwZZnnEL7JHg5M68Er1zJY4Ik3mQ2
mnS3l97aHyJSJaiOPUzSf4XoxbhRAyCi2ZI8Rk4WUS0jqCYmSWVFcLqIJbJRpeFP
a+a4xh3++GD4YkPcpq/cxUS/vpMqKPbFY0abvQeZnB9zxkb7jsoa0wFgOXrfWngH
4qRi79zBuE8blsGp1oEIFzHitGv7H3j4M/spI7BAkk553+x3RcgvMiZ9GC4eiFJ2
xF3jbZelREcv7BplEsRtOi20j8It5gydrpDpQ30SQyCwCBmZjrjTk1ie2GJu/HVQ
EzehbG1DACxS2+n0ZWmCCDlme3zmGXf4u5d96AA1ObLjxrFsLYjdDgY2zoDMVVxW
LfRLHIJvYlGeU/P+ZzZzNG3VI16gjVv6bcA+iSgVywKiA2mcEzc323LWHZye6DJ+
I2Om+x7PZNxx1C8vJwwjvff4VpgKXWIyezkOuIDAjWuIkCoru6KFIE8A4r5sIbV4
f5SnAXfxQ4Aboc9vrYfd6yl7A3tMQCUKXhzFKz+HoiUdoLZdahMjM1uvml1/Upcj
nl0GOFgiObm9hFyn+WxyB4Q6GZI7tT83jJFT1JBhfVLJfDBQXe4ef2n/7yr/7I3J
5ef0Og186uQXFH4pYsCbq2qq/DBZPmLVggApkIrqYUaieXuNn4H2UvexEglazaGR
qAxJcFDRNdJ7NXYY0AA8XPRHCNHoKMDpA2Hue5WlKUJwgalFhiIjMdvZZlphoUvW
08mx2Jroz7g4WjYpj+251s+z5sdgEzQEcUiCILC1f2Cxaoro0Z/VSf5Zjk4qpp6R
enlRZSf06WJ3A3Ja+OJCI9qjSa7Yf5o909um+sMztcQlmsSzE9vJMX9c1hxyz4dN
NsO5fh1tU6dFbYKQMhG+cY/3hSFROJSkcf1CCF1DU0F6Z+mavUWJjt53dAYRKKQZ
FoWTfgmSzXKaa8Zk2FUJ+n2L6HyLzoKiKXTS8QEcu7d8k3uCyl/xyEyoEiLKls2e
ctqHgm/eAaZuil8ujGd9NDgktSaZ2pFM+jg6ee5sALoM19zk/H8ffevzcHNkK8YJ
ssnilckWxIkM7anfB5lGnJFR83FuLq9elxd7noSBBKt0D5jH9ekxn8/2IQ0PHYjS
KtcsFR81tI5CL+pwpu6/NGddndyum9s1gcAqPG6GmipDVttkf2+SED+FXUnAiaG8
VU7fNiUMIlMMD0gLZ7KwMH5tgPDrXBf+au3SCX6J22Zn5+iQ1bbxjUtogj3Zuk3W
dzSUraxtzv0NFMyE+wXy7zUSvHm3/HAsSKqvdcdGdS21bzTPa3SoVSCjv3+cra6G
ZijEFTupt6ARFvesSlzk7LWQLZrEOxy7TjXWANzNe0MDOy2aOZtxSDCAcH6ofp32
L11uRhY1ed0h+lYW7yhx2qTAGgbmWsTbGxdnO3xE3fqknhdX8x/5VtBd6n1TIv5w
CKuJ/djWIXCDp658FgQW+btY3PG92xqlCLrHe9eDOPK1P99tSGAKU8i+xrmbC8k4
chFf1kX7Ungqg71IJGqws+xKhIfMtL/o4WI6CAn8S4jat+EFBX6ohw/aKaWbHruq
QbxnbVpPKcTO5Wulf+VYKxvOaR0NyDEkgcNGdnKSyX/oWTfv8hpmym+OBECNZ67q
/A7JTVOGd+raJplybMorae15Pd/mED4TTxaY7MQElO67o46LXOQnGZgyTYwlGji3
JFrj6jgaDm30WLk4KvMdPfTIzYe6bzh+J9Y5a5fH4mVMOPiqvQETGD8zk+R/M0/Y
XLN9SYWeFlGodvI0mvTQiG2gCoPyV5v0Pik+L29xPZT0PTxYsU+yb2aPE/R/qNFE
whD4JJ19N81EQOudSj53lrCmvNiN3YygozYIIYJKA2Td3YxKQvkHLn8snMVk4imh
cFWZTpR81g0kyrQDgFltIWprDAwmj/GYqi/Hwf7GpeoGE6JEgTfiKYAzeJ4dPDqP
VUmM/YPic3NTvxzITjlNz27sIgVu8E7mN6y9/9jH8x6WXFzWaeM4ntubKBg3bGY6
B6vH0aRGdl4mWi0Oal0D3Mj5oN65S99W9SsUFm4fBOQLX2N1GCcpNS+X1W3dnGRZ
Iwn8lOLdpsKAJ3lgwHzCtTdxIb/l8lt5v+l0Bg1R/prXjQObqxUr70XICaaJ+NVI
5wUZG9OeCY4Wft6pEs1t8wzT3jmOdgMr2Zt2A/UxlwUG/sTzlejwZDpJed0mKe3e
jo8qGpUBX3kSzjdJP6zwy4DyoURuAA3XtXijK9FKdYXbOLFObHIzZP3qSjGYfuhn
ZKOgAcA9ZTxb61jmU+DsGlhpV0YsyVSn0d1qmVzyLGocsEWmTqqPK4PDsW3JFl6W
abOue/CwKk0wRtXHwF9untVsY6ww70lu/gw03qCT+St83qkhRcpjs0sdJq7/c1dB
yIYuLgif65cPNZZqirqMUNQMhb1aWDWkuvjZTKb3uaZigU/GIcJglwsnpjCBI6IT
l/4NeHGHnp2NBnkk2Tk3ML0YVHhI6fWYwFVj4xBay1FBOMf+toP8NbHo930ybQPU
82pu4Zp5m4dEpIOhOaPhwHK0rpXdOuN6Q3dtTnG4LwJlkyNxW1twoM8LXwE4knQM
dhmdK3Ip7RUaf/TIUHsR/gjjFD8a/g5gxZfGO9e4XcIZx/uAobyZIGfqEdC2xMvs
kNzdGGBTBbOOhJgFMkVqSaaQREFs8TdkDFEaUiJYTzrRo9/vlt16OA74yjig1hz4
baS921mIGnh6Pv7hJ8ykCSBHxjWQfoTfhD0F2o9WcGNLAZDXbg6A5JMWZ/MFmxLq
JfFd43/OXdeRUFA1RQghy5R7APzFjlvWrsC19Tg/adI5CcuurC9bUu/uluW594HA
OpoyzzqZ8CznAydCGY8yj8zzBgZy2cl/dW7dPWIGX0ymLreTJfyVBv4QVCeMbMxJ
oZPo9SXEyJOIpvip5aKNI2g91jBD1JeW6Gii/0eAbAZC6OUaRxRVy0OgoQmRpJmI
a9KSkhRt8jkQNSYxXQ6X8gMchIaxnDLGhlmYlzVh2wK3198046GUjxwyu0q4bwSH
4N0xXiGVnE1J6V+XaY+4LdofZmkk2HUHb6fRvfXcrS2o4QbDfX4RyLj9rOCeuWjJ
Vk7k6j4c/k3AvrAnlFJlIyeatZjYnR+ZiqyNrC2rKiXAaVg4j/LAPKZc5uMDxiDW
3sGDeTDtoQ8QBpAi7ZI/w9k73DO86Sdmrh95vK9C85Gh3FyQvDzcVofJ/lf5pijj
oqi34l5Bd/VqNuYnXNRvGhWNCAtfswQJ93kpxPH+gPwIBElW1WxjPJ3K14uSyR3+
BVaRnxDEEWYoqlSvidSEx0zNrcn6ktF8lKhZvyQKXzUDHwulQqJtnmr1LTyYzV8v
nJSLhoL+sV1ZdpUgz+OnSxK3Qv9bzlW1qTL/tbA2xeDp2pFN0e92Yv+S13h2p/VY
NY9I2MefTItSQLIeihRozDrc/jG/oRy1kcdI7XDdg4BIv6Tt4l/s6jLUBvnTbphP
uW2WgI3UR2zAPMHhGimIVKKQRh/yhpbv/zOjXm21OL6CoIjXMOV1hxD5exl0Eyh+
Kb74yosraoYGtYWdJjQ4sguf4lpPU/rySNSaCMI3qpD/tVlnY2gvrsVedzMqfpMN
pgGxufVA5fhnQdWUYVWQFvs3weaZlNahbRItQO1RQ5u2T+OY7LXILmWtJDa8baP2
GbusEDcofnVLs3Dr2DwUJh4HCJtLx5eCz2OUGSC2RGLRr9EaDwqk6G8ty1ceoLGB
9V4FQl5ruuOku6BS+PyFLNlUEdiJJuhQUkBJf/31DggYqDKkqXM6gSPUL6r2k1j3
eDVHB/mA6NnATezSfy0cYO+LwRu3MHuIuxys9TzHB496yS3G2hw36Ivk5X5ZetW0
NrP6mghP/BudywXR1lKWI5IevZ4lGrTMmToykXzQ0pQJk2uCPAvzIM3wmrzKf+zf
/pflE0gQnVfijM4PIIzXCfnlGLR5zH4Hlt2D1WKwQjPOKtsNJsmMoUPZG7VaOe/p
JcFPOJmAu/3jkq5MbLIzKj5U8SQs131+tA3LpoAuQItG2furm7RfbK9rc7P+eBeD
YVMYC3GMyLs6pDkeWqkPeBql+WSdgixQJHSg4n3UUjhELo/WbQU5UfKrDiJVXR9f
e9mS3kgrv24n9kOinBTvMCPGp5tGGe/O/pdQIoWhTf8vMGnIX+gjaYPwA5NueZWP
uU/kknxM7r8te7kjvh3Q4EcDexThRnn5K7STNpuBUH2YpMqE4hAF/FMPKuqYY2YD
nGK4CMAlGJGEXmE1SUUsGV06UbcR76Na9ZtW6JlTfw5qTwQGzz3qCOtSmDCJkLaN
Ivm6c1zKKLw9/DQDXmKzCjsQOoQCfLYFHetSvjvAu8K9Sn5M7gn4L1+3bjNp7tl3
oodSFIGgEG3tz8MiRW5NSxLWkdkZ1p49FPEkxGKliecHOvUXOr77WkB3x3aTfD2u
MY2P/Gksi35JtmMDrNaGxhL7w79x6Ws68UzBQYX46ryMx2Y6H3taP6pRJw+vLWg/
eiJtgNLxY8LNmBFbj4yoCEVdifEZWG75qsIzhY+czKA8o3o6leNgQcRi7vQbLvO6
8piIY7MVigEyTzKYz9TkyHmEdWrEgbm5mrdDUJCyVRVXpWDt3yp2DGwNapuuVlA8
2vVCbq5nLJ31utEnKoiK9hslZf8y3KmTmYStE872I14rDgt9wQJB3z9Gtx0N2SHE
fbI2KO9UPRXuJLIjU8F4m5ZFCEQb1SCD0eoHydZCdVbaSNTFx9wcUbcmHvwG7Jki
O7nRY0YkJGKv2NTa8s9pJQiixqSzAfOEw238xhdAdilooXqdw1T6UwOTOsX5hp21
Ej74cvZqke5pFU9vdrYtH7GwgNvzdjl5Zab/1Cl7MGAw1qr9/9F4ecMgfcprMNXE
UTO3uBpadU2VXJ1FXYPDOW3AeWRV+pw402ou7rWyt7T5D3fcX1Jolqa23f7+b53x
5OooUdhVD/WGpkn+GohAnjygPg4AEnIKK0IBBA9FNTvuhgp/bcK4jYspHvtvckun
clyOQcHt+dApbQCJVpYCoI35oWDAWZV2nAU1/Tec2dVo3+SbchEAlvhwBY253W40
/w+ohV/xXneTg5xdZ4cdK6p4um3GB8cMKBzWY95qnbl4He+my3jgCLTP7165owY8
P9I00OBoxLVTed/sjTDF+gdd1EDyHUfS3FrMljLwQ/7wYNFit34Kosj19SwAK5Nj
YpO04qxCU0iXiF9NhdVFVwQvaNyITC26zcx0G7JGibTdZzVzng1Tz7OhyKbDWqLc
XTQ8t3QmsWGQwUQ/QrNMSvlAcj+dvcRdOmletZLsffajzv9fhntQ8FnlVKc2zNu1
aVn0vNCjYVL0DVVRk4f2UMbjsP7h+eZKjqviRgStRWLQYkN3WpQJz0c1BpP4CDeb
N+Imw5IKGiWKWjMHqmOPN64+Ggo5ZgHTLPLO0HIxtfWKsGOoFan0/fLOqyCS1EYp
CMB3SEQcCBt9eAKiOGBMKBk5VIg58iM/OQmOUec+ad/D08UnTVCHuBD0mKvYDHaA
JyKbempwLe4477sSMLlUTxsyr7NDfAOefzgJW/jvBpo/WsmLhTwyOfdXiTpbVUsF
kjtn8v8wIEr4Bs5z+MPu1TSNdRmiZ6/IRRueC3yB2oyNf4yeKL1tBdN56GqC6AAG
Bnzw09RXV6i2rsW/5qp2aXRLhYa2WD8kz0UsatcmKldm9d9eMF6cO57IJpEj2Bue
ZtMY0oi2etrXz/F9ubCRR2V7j8Zn2JsY9RXn+xFEG29MRN/qxQonxHaeNEZBeLvD
b6ffPYw2W11fOar2tYIrSXJQmbyc0h2RAcXdQMMtw9x4D2xl7nH97B22GBgNA2Ri
7DLj00tuvBmnVoUWYKetVUHvUc18JFawHNo9X7Kfnz1KI5QtGQwrAgnYaWorUUlh
co8qInfs6Jn0tZguRtmtxaV6pFAGDDKbtWZWQAptihEnO9g5hNzJ45SOtMc3FLkH
RBQH1ke9DjowX5TgsYhpOq/cdFydFBnfJ0B8ENUM8qIZz9iTO4rtz6GtWjUHcO6S
fipo5zkfNqjseeNT3dUhRPI5Bl324QfObK74ijFtSgb9196vw/q6hHnUMMcVwWKZ
yGAtMfRvObnR9EIx0q/+qF3jWP8f+ntcOSVjwfTu9PkD1LUifqef2h/KgleIm0M6
SEPzNkV4iEOgZLOIcj47rM5dk5BE99qBrY5Ye9BxeC6bKsbRBSGhKc8iybRatEHb
WJp7txbn6p43gWVkRFXuu2uSdGb5de4NHDWYKUO/yOzzLTFiySnggPrO/doRVvil
bLBTAtqxFW25qVFsVCSLo7tfGI+khN2oBWezoh/ffrjbs8rNMKBJryNJCei9pcUj
Td/A0uGT5fsyHvWVr8tCxCGTioZglusMVFqH9DFGyhMKKtPHOMjrGD0vqBaCyUkn
NHu1Ph4Prwn9VkOuQh++0JXm9+Erig7lS7YBzeodgT4pD1wFgtfCFEdZ0Bib8eBA
eQ4uMGtlsj6jdvMgZPKQBO+TpeYa1E2/ow2OOQ+6DTKkJEZ/PUIQp943NKUWLyLW
CEtWnIojE90YE9oyJF/X9pdQd7GKLAx8jvh1dsgJOLUgCbh+b1xAuit50geRjIlA
zK0aSFAbNin+EzGr2h1udR74ni0Hcy41W1HDV3sIlUkJPMMEDSD0TRyMNfap0BAH
5hrnU32MO/qBT7M4oxir3ZKwpk01llZnDn/60BXMB35tcktN0cXC/387cjResYTp
XmOo6rUrL/LLN7sthTMn/abrUa9+ZperwB6dlnkwjtF2W49MheojxpeMYQuCacfC
gYPwRlUvJE/bLXj9mQpSAg2vWWoFmUQlvU0tkeYFBPipmL2Cv+WK/DFnQm653Hn7
HDVb7Z36DFontJjr6DzwGhtdP+iqWvLyuwF+CmMWpSaX6bKEzIqvQ9acEOomrz7X
gXYR0ymwnXvtFrOOG6uwwMAR5nxzMKPhgxQ63SxZuzZSH4JQzolCyGdglcSwNyk6
ukAwRYRfHF4nV7EIpHIYifP07uV8kGLrinBOeVx+qu/eZFLBdHM3BLaYUJkw/yZy
Wrtxc6akQOf9CaxUmAkGQnNbGbaicxUqFNECskw+chnfHZuoEMJ8z0OUlOLYweLh
+GMRZnciKygDZJ375W2LcKHCOQgm2ZuxZp60L0VWeD8eVPHRs9vgy6lICtcQiv/0
YTjGfAHYP4CbuTNfkPBfaFV9OVLKldX+TWv6zdKAXbM8WM7NWlKlb3tff3X/YFvA
8THYoxuHWiCNXN6UB4j9JL80N6g6/4eKCjCoBcRqtCVXiXpzn6deOoPd3sk/itNR
cCRLydfZEGQrf96Y6CRmw1yNircgFLy0ADaP9PiZkqi1Adz1YeBBHE5sWsPDz5T6
wOqijQN2BQAQ5+gDsKl/kF9RXnaW5JV+wMno/aswEQi6Z+/XpBScKegwJqdfCGZK
MyITudWtovwu9Ias+5dysw5He9cK80KZERLBw2qn5WXuU54XEzzPBhVecU51085R
KYfHouXPMlp663z/waq23Ne+eO8jPm3VZjLYZjPckZk12/RBKoiEW7zLvFi1NprX
6JAiYA6I+dip/JoE3bef72OerjNawp8DEI1UWnPFoqC+wvKpoJXefZH56P+ekYKs
x+PyEnrSwqJUdZ3b9CE63PVg7lEoLJzPDFTUQpzoxzlfFU4+fgN339RbHEtIX4ym
KYp2gPRQ/0vV7HbYPxPXsYd/70qFFKB64raCUWIZswrMAsmXn/pSNA/9PH6HRbiz
Qpnqi6IgUm+ld64zYIz07AyokalI2X6jHQAigUs1f9kGB/6g5qiy99bmY0ecC1uw
CzTtkEqHLvtYa3RE47D70kX0azicXxwk9BMPOBGLRdrcZI+tupG/1c8huikyqG/I
O108/3rD+hrSz24ShKNHfOoZaKuqEkZcLjQQlpFF3OqYglk3mWfZyFMl7qahBnf0
AFOtupxXqKutkoTi2853x1veZYUAe0HlEiCxpX09n0UVJkhHJTfg1+EVUAydCmji
dbpYDxclBj+X0F2UyVqhdewgapp7PDX6HkKHCyQzOYAA8WvR4DbfxhIbL6P9h6/d
zF7bVMJssDj9k5dOmJcjpkDrvPrdnA8O/lHjOv4zULIpagmJghy5VCiW7GMIfV8C
aZctHpLK9WnBf4+EFNNNAAXySDCfciv9I5fv5IjUiTkQp6yYxJFST06L69WDV7Ko
eZlpWLoaeYSKTe9Q3LCzj+iHUiYssQRhUpDKK5CBkYPLwv2OA4Z8LAm8D01tAEO7
gfR3ZMcP+z7whZ/WqRzqKWGmX9NRdaFPhvc+ieB1oOJSB8RrjdBKMtVmBP5j6202
Bz5x2uNLnBqm2AJrM2XWPv9lWf7CUz6tiBAQ3LPZxcj0I25kSZn0T2Ypy8T7es59
HHt0N6VvZrQs0GqT6siF5RGNvoLLcEpjxuVYE2RztlGbHszzbTdqzroSCoyc2mFw
SH2RjXlvS0UdjScc4axLZuNM8Ff7O0aqg7SIhw3chStYsF18eCnhUcQFTnZxFpEv
jMlTK3RfSh9SKZ0fL9oU0EtZvBmzRy1D+a/vfRnAtlQD215/onhgcAxi3wGUQ90E
9sed3RgG1gQAFvH8zbN5rHjEC4xRgcgZ+xPG9BNCutL5veWAQqQIqlnct/li/Tor
4o5dwHwxxKvWCkQumN0hnYnxTSFkX5YtNGs1LKcNrQsW/UOqYqrulJXthcAH+ZqC
WisVhDbROtwM5wSPYP+bNA3Tc6mmptxfXJ4mD/Kq+J7g7GZh/uhSSlxUV98Rdw6l
5Ngeeue7d+9+B0x6aKgxA9Tj9C+cCg734oDg0+LSncx+3o70yinfdZK6iVtJ0xpM
Tr899q27id/fFfNJvbMYSbgv55jlQJl3pQ1ozsSE2HGxsKd6x2vz6OeqanhxqtiF
lYmL2TsCMSXlUzIE2RnFTcGpN2PaoSWpAiY9SRhk7wWcaTbDxmb4tT1X5GzGkUh4
tgAL1RayO3CKIh9gZriDuZ3hKoYWAGQErux7LpXo1knZaPDCEg08aOfFtDVx6c7w
Mq7tGyjeEiyll7lk8K8GPXqybxxmt57lzVLoaEsqJ3bIVOhhF3qb3am0GZSv7sGg
CLe8BdhDhMQYqCTMp8i7h6l2SYVYeVpk3hcUZYOalXp47DUC+GBBkMt4aqiA/fS6
5iPpwYXAVlzSS2kAkfUoymgKXFchXB9VeFy4YVd4L1mW4C0w43kRUudv/BrNh8IJ
qR37PKstFBvLPm9rZfKrfvhOSevmS8a00XMSlkodLvET5CJdK1cJNafxokJYnbdM
mlkbAEy2hmX048GzEf+swzTTwtBD96HA18wQVRftQV5UXGWMASFGmb+N3livEHIt
t5YI8j2wI6H6QOffTR0x48hWlhH1h3Meq7Fv0SSYSIfQu9lsb0b0q/xUGzl2/oKr
LGlnWQaFddpLUzZaY8uqt3wW5PKUEeD07UoZqC73F4zDkwNL5Eqz5/VpO1L8G9kO
mlJm5WFvmOCrW0+azcrXymKHPGC9ETYV3NeRFjQXHB0MtQlf/E3z8CF9Br5kWdgg
wago7thA1jY3egP4aJdXfOD4C7Ekb867JecK3fpDJRWZMr7xPDS8Cv8NBN0LUc6i
ynivaQ1YoL4ciNQ8BW/Z4gtZvh81IXT8zNTSlTqW6lEM3yy+klc82KWqpSdRgH6S
YUuw2iDX8bxUWMvWHN2KIj8FxPBkmtXmAjBXiJkOf60dN4tEUZ/wZIUq0Cko0Eq2
PG5HXGol24z6XKexf1kYNoct1hH56vcV63LqnneueWJqiv8vDuhemsbIJQXz8QJg
MEZZAQFTHPpJPA0u3GGkeu5OI2xPpKETpXIESbfaqmXCFSt8YND1/wZoh4L/VQG0
Vx0KIiOBWBMphozSijiwQ8NnAvJ3gLQCSlxw5n7ygHi3nK061X6mE4q1/HI7eOX8
qP0bXQvGnVEkzId1Tjy5aJwx5Roubk9YPRjMwp0OUzdVypHDuip3+kssFzazn9a+
9NNGRKxb9fI+ji8NdOvP1TThMF2cE6SPFO43zr5p9KJqS2+j0AT8FcBRYvVe7QHe
bspsyBZF/8xi5xkwywKysN5K/cVqMeZWeVTLGWcwysPukUUybA11s+03V1S0RtzO
X4K5wW5bJyJS4ulF9DINUuiunW5IKvAwkADXQ4BAruj91a9ndY7BtU4kcbQQuoZR
GDvwv7xCn6o+BTDd48BV1m0+fV48DewWOK6gGoFSzGoaAf5m9F7xqpLZQA06676a
icAJk+5LbYYHEXb4/PUBsrgNBSA82emcM7cVckZnjWkWuPsN4cGdcJahCKUPtLbt
YZm5HM1R0EMuy+NBbWu1FSDiiilY0PIL7w+Nc4ncNl2j/Snck818Y4tkYIoGgsG7
UBJkyJMNwiK26Jk3PvglkvxYut1NZ7bjVwsmLOiB0xjWY+iUmDslrFJ/oyOwLRiR
g4s/1FhBbRrCRADWVrTt4ArK70uPyOXjSv5Nyv6esDo3E4thnxDoODhoYEQGH+me
NOSxUSoB/3DlxWTmk/yKQq5/dKL3hZOjg4MvFMPy5Z//lRvrybybEj4KcsLH4zI+
mAWvB/wE75DX7lHslivCRFDJks6hwqr/0G2kj6MoOJBxPOhvBVtqoX94YP5GDZuE
MuMg6O8mFEXoh05Xe/wa+KcGkhCLOTBKsvvt3/4LZEBZjcL4hzw26Z9SEI5dKKDg
r6z/nlhLh8/lvBgAeMuzP50eaP9/U5rbFO2J7QMmG9F9dtwgxQZBczY3wuNEgdFX
fqQFN4eA3FbY0VTexa/CtqnbTwUpsKGMB6IEsXZbxwZhwxALmmHcV+IZLybd9B7e
vPedI9SF8ji2O4MtTZLnqy5WkSbxHnv9Jp304s27+4kz3A3tjV2qysqnOMgfjIZD
X8Cnb20jvT+zhwocQBgpRZMin8redhHY6/nnkQrIAA1U+ECC50QxVmAv648oJmZk
r0KTLytr4v34rd/F+zl5fMOBw3AnBU3bneh22+AAo/KmVT5/BpsMo+bqqDJsWeS7
CZ7TyUMARHSAAzL7uRSoU/u81iuNNNTF2aEbbPm3/EIruyJ8I9S8MkfssJsPDGgx
l40Ld9L+UAhtNkkuYdX9zotF8tFMJ7fDj8vJIiV4iHhIP02x3faI8svrArWBBuqI
EwLx0E5Wfy7bRBTkNTuHov+0aGQnyJOZqcILpYh9x/EIrKDMjmTpOOx+HUZu+/68
0/adV9RYgsZLP2a0nj5dRgq8bzFciCdosffhtKkmKXXHOZCZH3dcGqtu168a2q8S
Ej5A2kYtiFssq7KMvOc1ECd4ef3xV/BxyIU/pZNkWrJLcPqc6txT1oMu7eVa5fC7
1ddQdHc7FHpcHtxAGGbiCRyQ0RNeQMULga1GathLd1eMQjUgbg62vkdZYCsgusmB
Uws4KtbmOK7j4FOYlsSbwIjjmrwMDFGS7qhE64bACq195gecs+t6lBFFuhJRDhqw
KHoIntUUjZtkLiDeimkyMG++z2Y/O756un2P13pIck/5xMa7OqTaFuK+Yy8bLXfW
FitVlXGVDd7HLpOGEQ7wn5zQs/BYhDkLK2Pg9TM2yBmKbb6IFDgLTIl2f/GQqg2R
3H1TVQmA9NAohGaHGU00ooPF7KMWXoRLz7eIc83FIx3yF8yoLp7eIyt+yg4AGHlf
0P6sl6cbTraSlO3jdnlMQaKdzr6G08wBnYiHDqr39bApHRyniXCb/txu/5SlQDub
2xjXM64BIEI1DULElZmie4TxkEqUHitwPsoJy/y/jna4Uy8+19jxvqK3XnkSIrGf
tzWO0VzmeUDgKF2QziwUjqR1MbruE8x0Dg5jXxlfRdYiko9v6hQ/iQnXnaDKTqT9
Q81yOceXJsU7zbh8P2HppzGQpkwOdUNwVIDL+dd4cqnS8DTRAoqeUFkFs8qDZhhG
BdIatpiZAUM07r66m0IUzuGXwum9iWM6MLEzz23UGBcPfrWgNdfwwNzEG4P8caSb
/XvrX+BQsz0DnWkyL1pBDm3f2flTpNP+WQA4uqDSH12VJBvWhI1nwNP9/D3DIFYu
UyH88y0suRC8WGkBXcpo39RCuLCJaidIzoMQu2OVBpnqlrQVib6AFy4evyH9NUmi
7iqpjHLxUcTalzknfvT5JE0I0g4/aPUBevEkAksvqWQRTlGfiP/i6qESF1ska5wS
vWognvCUEfFbv5wOZld5C0560K7gToSiWZE+UwR+BZwphyCQGEsQaVL42nfAtowb
tMom9wsl1f0WP4+DXqupYcwV5F6N5/ZBF9QK9w98JAxXszDNTyLWCh+WH0RbpMQB
iOn5ZoJ1rZm9WP29cc1mSDKOVe+P2x9N2uLdiFh4XYRTHDHLIG4iWNUFrjn5MwfZ
pC0r7KHytnDKyK4F4P1PzhUR1IYPukv9uIMp3Mpccsy6NDhGBKBae6ao4bhZh1yM
yguXinXrphyMVVD5doif1cUnjwq1yiwZMilFDSGDLQAoigaEJNeV/TQfckGFgXgt
KrLnG7qfNRi2uFJXe7Xun8hJZMepXy2PrPx66d2NMTSJHeBWS2v0V03PgXud9sTs
A7wA+YtmgEaZhqqldf3pSXBzlMGPcWqozmBhVO0InbOZEcbSXAcYfn5rMca09Xvj
kFpT/jGVcTLlCqWquQbzvPmI5XB+k2XTAl4noJjGxw7KXgfENelGq2rvY0vp7aev
g8iElcBep6H5QsKjRcX7wa9D4LwGJNGIWeI6tYYULHefY2Ox5CKnhfcYESAXQmod
ViMsuvsDaBQ/+8dQxwnBomthyICTJUntlgUChPcnaP/Xw+JZjsadLOADbgI6scKw
fNu2Gmschc5sMtun0pJEdh56yKTM8QzXFKfSyeK+Y/Vdb/D1boL9D/gGWsKjNl0h
yhpojK0gVw6MbuAzm684TpznLRjreCFJ1qHEgHhm31fIjVHiZUv38bC0tEgi31Qb
GZUikgnoKBqsXkn/Mh74TAWU8LCQvK3a2LrSxBJH0EFOHUG2fmnzAsLEkt9cr3Zb
yXRCebzDcicNPSXYKuzXL15Snr6HvScFV3VnAbo2LLmt8ynynDBj29Z4R70hC6aH
FdD5THItsJZwe0qtZQOgFSlZh5cD+3BwMQ7vc+hPISKJBJV7/GbxgWWSMQPatS6u
ZtekqGHkKqOb6g1r6KLP+waMESvSOtJERyLCTO3OCScwL0SlV8IRsKt2F9fCphT/
YgFiJikpTYNVbvIMVA3DAtKlxu0jwO0KK777AQTzrZROK3/N7nUu2viBojvjK6p3
d95ARiMgx2mBfG6UqgLFlPJNVWaijPQNXh2MV25gapdTuiB2zC3m4r/lv14GJfXc
gYyhWeG/5zLnekzCzAamza4Yox3f7RMpuACZb7LTgN49atthO+wwm/uKVgDQG4Jn
XkbrAgm72hYrqT1UH3sjecceLTWkTzdvz1aIuSQDUoRwW7AyICG1dM2t5yzLVEZ0
4jDLg4rfSjubKOVtuVYy6wC3aH4XulM8MuVbobUOnLgYyeFcec1h0ZGe9GTZynG5
kKQJAtkzXtcCR43we7pz+RgISx9U7hMzRJmpRD24YnbAeerwPLbeR8AYj/JVVn2D
MV9mr1dIcUvEmlUbizL8gWtxTyc10ansV6o9Bh9/AfyP6kufdow+WqZJo+JyL2PC
1mpNY+5BTCyQZA5U/QD27gSTx/M0jrdJl+6zitUT7YjzSPSQf3AkqecnIey1FebU
bYrPu5zCo3kj+HroXAdhtTNLOsNVD4t+O3Ym+6JYQTmTpxyF1/1tkxQrJsuPRX1m
XznqoitHFhWSujDBuCt7ufnUDKieqJRI6CmJZBjLscMPwQMJmykvHl7rzA2FZGzk
hH31tAUJ9uk/DbRlU8M5tTqBWzGQXx2BvW358HQNXhxH0ctJiWod8mdYeUb+NNOE
U2/3Chzpy3UbLZnInIirZtq1Hv9WU9EZUpfMojIIWJK5VaRf9WonAxCEO3T9iFuF
wRO9yIW6cjCZFEvcG02+146RJc1piB/YLCKaPIBTRfUfl/u0tvOWyswJSSs6/fJA
x3Fo4puwY7DdtYyiI5uDB1AcZUi1My9kGoarsTD6OX6QHdIJpnqlcWGRNfXDsUST
/7hCMwBBWf6r/oTqp+LhBoObE9FdkQSf1JfHqy+RJm63LGc5pbDmMMAJ3RdxKY7o
HgUJB0OZIykL5jPMkEQEkn2/Q3qHoIYzT25AlvjYGhbwAVmIuZxF1FO45VjKl9aE
9toowzg+ZXgmIDmC+rLnP8id8y8xNkcRjnKiHjgakldDbUFTydwh4rFxrXndjgnS
Nhy+dWulq0VnDTVeDDlcbLRzF1QYw9qV2SjqE50yqOSBFHBeQItyhgL8+tNvnNtr
WtMwc8MC1hZL3RSOJIxkJdnT1MwSJvf89j32SybRjFWJ8/1jLiuHZWOp581Rs/r0
WAsTf1T9DpBIC4jpIUWWVymip3b1stdt1lgRR8W5MJmmaqSYypjzz74lIspAopAc
elj7zpQsKkyqNGxy+EdDYaO/VeFjQzqIFhvny1ugu5y5iSjhiGPWcxkqnLBep0FK
E0xbVfobi1nsgnwa0m4QnPVH4Rag/xbBfUzlBJnP2wE+AU4XKX3TXYQwcGs688ih
+rhVrc8ddnzvla5vt145xaW6NomkHeye3dGw5MdgNyDXUm1m1au9HEhYdD2zowg+
/ryCkbCdq5GByGNtiC4LmK60uyUWn1CYEkLVUMfBT8QcSCnxXADAnoQIFFU5cJUS
4RQBqHbXUeUf9vV28d48Mcqkaap8qWXHHJh5quVFfgkSWDJVoFJ6T7VhTEmlWl3/
xsWdFfBWMCQ5Y7+vhJgJ4K9z7KTjvxKJMh3D6TZORq8D4JIlA0KluyScqqpiaBuD
cUtm2bbTDoNYV9LwL8+kUwaF7ffbC6Z/vMl21ZPGDsjZwciPGpy88cJikn0dx4OL
z29hphEymWzSavpRaI3IrO45xiwuKVM0+dKqsxjfOu/HR4hLg7teuZzLyPCmmc/u
RGwg6me52jS6ef4Evm/584qBtBoyhFvUfJtrg0X49JBV7NxxTJ70KG37My7EzgJL
Pgd7XcXo4jWHi3jOdvohqVW8CBmo22Da6xwSeAzwWxJxDxP5IG55gFVgSN59FXDF
jVlc3f1U+Qhy5u2aTPc72VVfEfngajjqG7yxeoC9QhhyR38PO/ZoPtHICwyrFSy1
vRxldwcZnBdv1OH9XCDpMizdpLvEbHgXh3fxl79/chKNUu9V3yhN9VU3eDD8OzxL
2hT0nHP17VPhhat9OdmvCzVKOcYVX8gY5jAYnhR/oeWnRf+YKHqyEddt+3zwF+Ad
7whtVGzcfvgDh/yRrRBfw10AY5Zc3EzWMoZeagezSlpsCivH+oAv6qdKuxUmzcUN
FUHdqOvt1aOQyVhYEZvxYYEtvEGSAueS/c4GddMqK6VIERxpd5llBhSXzTyvESpo
EbDUtQZvLncim5ELm/c9EFRtxqjGOtHdDa+surlk4InYCGPY6Arxe+/7ZskDJd9c
HPILIpz9z3jw5d9I1NZK15BFqMJ4srBhbfHCPnO6YFjz77gE8HxRS5gDnGtLHmHa
qV3EJVL4pzg0YQVbmbgatWeGgrvlxlZ+eEaP6Mq2nkWp7buHYUO5rJVC7cufsM0B
ZyrHI635A1B9rZk3Cn/S7HbwTLF/Gky5zbJ+ffivtWNzVx5fORPngCBQcS/jJdGC
pv3oBhh4c5AQcxxa8SJ10CTd5YGfVmLNuj0wzLYyrJw1Bx2kSNcvvk2m1p3LNXK0
+/IdE+OKVZnGLpZPLt0yFchmV/s9XNHUyKxVIKnJhKH9U9Vop8xAWfELnp4VoE6E
H0hp+AIR6byKyTHROLjH4DgZNON2e+mdc1Ry0k0akA0qvb867MnMNtEYHmhuZSQ4
r67XN2Tiu+lxMx3PLQYle6l5zFhKDDRGuUCcLAyNm/zWxSQa19HXuP7gHTMKl0/x
QzkYZL0r3gz3K0SjdZ6pSE5AXFrE773Ymfa1zfFVDZG+vYNsk1JM1D38Aa0xnGG+
lD2Be64hUJI0jAclN7S0xaWPVtmfLGFNnEitGm20iC9ID2DufD4SiTeObSBVX8mF
rNUBh9QbhNt5kC5cXmiaTTpFZxBdA/3A2RrO/xxjj7qZXjHZR+IXDwuhGnBeHvVb
iVI0DYlAfX5DEyaGleI71R0D4Nl0IO78wwKzF601ULlogqJjlXkuq7PG4capuDGz
rRBKB3dxjdWxrNS/qoloI3JvSNq1Py6gHtce+bBCX1egx6bfXbv4Lp7MjDU9INOz
45kZXqfv3g4LSLEdi04GxuSrPF3yd6KFr0PQDOUwvawxeH0ncjxNPACTtdBg4cfQ
ocSyFjsDuoWXgdB1rrC5z0bNtJ/1EduB7oVP9+YXOi6/L42DPgiDtkpEzwhKrvXX
8IQ2jXTypPoMb6ToZRWRl8X0u+5kNktWjpIfqVkZ4pn4NsBjj+a6jy5cQ5Svgvgo
nYm8TRh3xVxPjq3fTA9UoDloQfk5xVTJiphRbDabiDs0X3QMuu/pVCUFjbOuvdrF
MaBCXYHRavK/E6S71o+Ph1RztAGPQY8+EoZV7XybsSuuQdgR/n7z81l0nzNDzEUK
MTdasJ+70Pz3AhjAmmPbgSvFlmZkWzL0D3aGfFUBMjw6Qyoo4OT6BY2NVhKXD9h1
4hunBnxOk6OKixvrE66blN26IZQtDOZui+6Aj8X67u5cveNe/BUorcxFTazH9BIa
dwevdI8aDpNIKUK6bBJqi4W9QrrsKCnidOshsuNEYTpcB9SFw0RbfO/TkfXKCTRy
MNfSC98l8jYtXHuAd0ThPEyjJf58LnCggxP+o9+IFGrnRgMlZ1TVrZ8zE7dHZfFs
foWgdYu6hFUm+ri1As4Yh49U0HZC3yM/cDNdf3j23Qq0Hk4Q6E/YBeDLmlbyF5BK
jreTUOTcuk6U/hY1jD5hI+v3qxW/a3OWdvE74Y65UmtHNR7NLFAeNeDGXS+hv3UU
zw/nDc+dQXOmb8tjim2pwK7bLVY4wbm7h7209gwsHCVENwlQzzMB/IHNHDVbALX0
XummsEZpqMBrksBiJRLLFaNxYBP16/i0RoTbpP0sAZGIWAdvzWw8MHTSPDaBnJhC
8a57tFIDk9z1984VdGTliXYPDQLJVaKOlyE49qm5Qkus9flNZgjd2M7PZQArbC63
r+gJ07EzkTcxDnPaieq2c0SN+Q32Ejqm72UZRdz9x8Hdg4GmVRLW5nwqhN/zxtGx
VC5xUdz2NNTwvFU0D56uZPoHPaFIyvkro3a8Rs0tCl0em3LFNU3/gTaL42EJdUKB
dBcd6M/AA6Z8qwOBbTWthPNIvb9T1dpAMdGF41vTGCjwx2fEIBxh+GwZaMsGVvax
5biEWxUR5WY8pfP26HzugpCK5M/H/eJowbuScMidoqJ1LDLS9m+7JIYJPFdJRYUQ
7Z7rRrzt/6W++t764WMtCxB3G2zLwLQ+g6/5i+l7a4FeyHcYTBWgiJ2C5D3ulq4Z
cBvreLILCivGFCPiIOQreh0x5BpXNHX7tnWgtvMhaqzLrJWkrg6TVhVvCnh3SU4S
DSi41CdcWu4uaIaN46AW+jl4hL//ObqWlgvtZmb1RRKMS0GeA91S5rhDiLuTj+HB
IEsBRM8piprbKBNgMuiD+PELtf6fmmya96vAtwkv0A5YicuAwqBDHbIiXLkDnat9
5fiTblAt9gifKFKcOWhPG/QVjWnMgVw/ekJ7pzskH4EoUD8x/097Z+iAKKhuNgJt
dPgwtUwHkWPwsCBPCHrePdtfgie0ea7qJjw9blwvczlC2sGVIK553BYtSsI7JhAi
win9IoY9OC/9k/ol737cayQMJKS6Jwomc7W9i52tZ+4kpPvM6C7okQc/nTDwNEZt
YFJ25Kx4N7O/9wB9WXvJUALQh3JbSWo61taF/R27EUp2I2ZIB5Z2Ir8cwyOwKiai
DTzy5ffOV6QimEg52wfmpKdHcDoB4UGc/aQaiMJQD1me+MUDRwoksVf2Vm/fdPCh
XbmvyqrCeqoJqOStoTifk1Nik2OVJBmdQtUUmnV87sn69SCICMcpL80/hDyomJlU
JFtiBNkC0ITU2rEVXlKMH/YeRNlSz6Tu4ZFMhcq8RIdRjuN9ISzeC7rzVxr/PoaQ
AEnpJLVo0ar7pC2dAMxh6t/FiYdlb1rl69CpK0zOoINAAwhsoX3W1wdHC3rGGmgM
Oe57TolPD1htuKVoi6pNXlpbvfELLkTxXjxwKPgt83m02ECJJkG+CV00SY+2WanH
mgmSlWHOxL4Kw1Ov9TteZ+JKO0AjySH/YceIU5Db/sTnztGxQKSsskt9Zmlo17KS
O6my0b/Ma6gjk0TQtelfh9E/mRiEB4qUAJH36RoR03gvWmmRl+WsTTS+u7Dqu6Is
fyMcHDl5FrMr37FHkbmvapOGMrW8VdS7IyVmgUnYDawlfpve/BATKskh08gLwZ3M
B6113XrlSLWEBtwwk1VlU3pSqjnLj59TXwXzfJXF+xxujzXx+KuZ8fy8UCqy2285
YIwt49krTldYd2wBvYfHM9JG0OfYwL+irA8z7mIdNzJPtr/wNWB5SUwrvMDrdoCS
THmjJB6zPJ9zlWTytSeGjXtLvUdj3HRfqrwcwR9WrW7ksschr9SAkAXkNc2odWQP
eoodFzcV7lLzJRCD0cgkD+P0A4BSoA22K1fN2PlvWuGD2OmMZjDKV6Bzn2XsHYYx
KeKr8n212Iw7tZUS03oE4k2Ua+HrfUwf1vN3SSiU9SaxlY8EJ2HVm6Y+StWDYUXt
3dM/NTtrNskquE4pW5ptwuozYOA5+WH6tpD4vujkZhT6r9IyPZqP0PMALXsnL7nb
r+tDIw1BBwpe6jJ/3nTDY0eqpfdeNIKAJm8DiuMXzpG+UAxJfw9PsHxC3YFSeLWF
+YfMq66jFs2c+BWsOaNDsUOk2PX///FAYdYOpu8l4C2lxCH1Kp1kr4wkxUEvLHZj
hwm2f8LUHq0UuSGGSfG2XiKXUlWxvrJRTo1JRctDCkm/fG4cfoZXfqLATrf2SXOs
V+5zYBfwGH5wjO/dXGo/p3utp2VoULjcfw3ngrqguAsNakGy0c81mdOhXUOttSUM
c2UUM3B+zFzLSrKiR5vdzqAKnCE40aaIMgRCowWP69dMqfa/nk+YGAZjj63/9uBT
8w02DtoaiXNzMKlUf0scWcIqMM04bMLiMcVCFEnckxgGsQh+kqhPyK0eeRVg8M37
caBcPKXyRnR0oLqIRFk31LT1f3YX9ksoexWajSolm5Rvw5xtNHfCqM/L3pzVLNbh
CCeehgDW95OTy15F9cEuFslqOPy0j19Ntdp9pHzOpHU25N7geN8Sp46HxHH04mcL
SbD0mpFgXYfHsotgahFeL/DQdC0i2JUN1BjMRB+A7ViM4iHto3aHcAIqGmwkXvuQ
whCRCWul/BVLtQRN+DhXAs6yCOQRSK0usqFoopOCGdMG3I113N+FE4MIaHbPp3MO
zLy9XnDyAo3T7SBLwQHjG/QAqq1mKsS+2LICLZPX7PaC2jvFiWTM3qfBPLn6ff4i
2FXtjUwd/W9vhrQR3AuQrSin384ZNzwCmUrZO5ja2I94juMSuBDpkjomHrvDMKq9
NxeIKg25Te1OVZ+Weg8aOegglHui3ihZcR+dwWYMOfFc3AGoWIqeaEH8+0cjDcTP
2mu+JAV6F4KofTY80ZRGzvwigZsAokekYJ1Jh8Jq5Wk3l95LZ69QUYRsYa1msZl8
X+X/CC/V6etJTw23hcZ08MrGpMCzIxMeugsuomno5w1xaPIe2YTUFORc1HirrnBp
yd1vKBJz2ooBlLW3ag4Mn7x1T5k6Vxj5+SEVrmVx3jxoZqW+Kw4vwD5ymnZf4zyI
pJFWKD/XU711B3m8ky6azHSKz6SWUGEahfRZocsfVQg3ZMEMM6wuXazAzdA7m4aA
XijNwkWqHDw9JDXtelSCB9qinZ1W5lD7C7E+AeLyLZU62ViRkrNgNzOadn3Iugox
Cw3kwTcQLdIir/WsrQhG4ubLlIalH1fGlN590r4aHiuAGzRNJBUmci5x+10PpARr
rGxfRGUMqM6oamGJAtmy5Y8Lvnkl3ZXufS04apQOVbldZc67qx/onjisTC4VVReV
z8OtcyN6+slwzSO8LdOjZ/NK8pW4Q7nCmu/dU3h+/4/zH2ffh2clElN0qWKsvBld
f+qtU1nmsASIT0rmALQ1M/7obCH8xPscibj8b9YfT0kWFd4lF7lga+9ox8ycnKPt
pD4wCBEagAS/wgGTL8noi2G9ovYygel7fPqz6jyw0sihDHlDnoh+flv1+w1zcema
9ZhuFXoNlZbaOa0HGre3dwimswyDjbSa0bVRhmmylyI1QqCb18g/oXi+lZapsmx5
FehINYXJGxQ8kxKUMx3Y3AZC99XWcCbQY56h51spa2tG2wHz6mtxWsAIYjpSMTHY
gl4H5xOgnKIFLtdDTgbscGeLKeWyPIUklaXnhO55+wVWepkSuyjppCufF16uSzFb
42QjuxV/lpIWk4ARw43HeGZproSi5gIHWDc2x/P6mRUp5KoGgSgkGDRVyWHDKoIe
Wla6KJU4CcBcCGslWz+YF2WO9nw1jJC1fbV8E7ohl5+bTLJWcmidXscM1dAxnsC/
f+HWCyW89orV4DwPicvdLPhDnCOiqphTVdUe6RUwTso8CGuUUthEaluF5bkM9scR
tlvJmpKoGwX8Yx+O/CvD1iGPGKYd8+G4H/dnHb942VvsnnADobo98R2mulCFdH0y
W4YBGTpS5x9/hGJLSAHpwF+M4Fg67e7NptbSe43sWyYcvHVagrap0QCi3Sn5BWCF
khRoMtgqSnJwpQ3SKTph7pBWjQut/fpQo1KoIiegwoQPUhubuWxNjpvRT85Dllyd
PG2yBoHDj3UgLvozvFpMmg/d1IhhGNHaSI3Q18Ys2w+mMlNOmk4SQexSGKasGauu
g4jsWexatFWsnNnA1OKZVjpVAXuYkeM2B1nEqTsR7NckORQgOGeBmuMb4WD7nmgp
pGdon6KFstW62X8zbXeVwlLzAVVBCXkwh2p3BF29SNjMu4VOobf7xjZtPSelpw9t
rLKNTUWs//hcF7OkQMeQaZxqEnsHbm5BGqa4cmAxJP15IGijDKKi880ylzisTCml
c3AC6gISSxshtQnKurfU5K++G6diyTJ6hsitIp4VDbvUiCi/OXDEIQ504/jgrllx
uYtUNGbO3SoDATlsrU2VXYl+PQ/SiExCDNzB46he12lFSb7qL1wq5GWW3FtkMP/G
iJXune1nicOFq0w/2v+5ayTBKqu29T+eXIQtyLfvuplMzXu6+fNqhDCj6BTajyMd
8RNZxmhdm6iL2d2E9dSdsUOTMVlXxltdVFwdtzZa4kMlTcQaH4er5gNB/qrqvNF0
eBrWz6/ZxM5ZrIKE6tKQc1aZloz1Jd44+uY1AnjbV22SfAw7flzdSJBsugCupGuW
mI6qzVFHlZZFE+xbeM3UlEOuz03ZfKSUAgvhNRyMK+sTKLgFI+0MvmVThR2/rAdH
JsiI3mzcvfcspOaCB/ZcH0KHPtcmEP50fzIs8101t2A1lgMWrvcCu9v0X7I+bXz5
4m4EkuDsEWVXvD6kzyDcF8Cp4nJb9mY0VMkLY88Ex9Jn4hKJMSSUb0Wpsw3VkTe9
COLdQFB9FErhupOcJkHEWSGWsiu6Lqf21bN4rlvTSaAJSNZ7/0ler2SNII9rnlwi
M6hlWm4Nscf6oqzAgkvQz126oCNqCTb8tl6WHS4990GlNag9dc8KIsuBfm4IuFge
oi3kN2EsPxP+O2wA/xweL6b84FgNbVp0ubnZ61O1OdsjDM6XrdJJddjihDFWclg0
wQ4agmDceZVvzpphja18gZtiLKMg+Msupsi7pIpbgI4aoShaGk4CNQ58AsjVYEbs
YjRjp2Ie1Dmo1lh08IRMomvDsSCSz9PwBJuxmOyHiK8+V4+PVF8kSJit/xRUx6GO
6emSPRO67aehtuDwMFPnIlZ+PDMW1FAjIntoiM0ECRNk/rGMJ/dr3zNhAxwkOLoP
mtOU5ANd9lkYdy2SUpKcbOrQohQgtdKEp8olgpi6GQ1Bpec4RZ5TL05OIKMcJwM4
d3dN9RUY+SJC2lAj/7xcBttW7VthJcWHWr7MVEct9XRQAchFBLwf0xrrM1WcxiHa
I/nQhRAhpyYtBA/i1htMQUbhOyNFWCK2ER+f6tnosEzDxhs+QnWI89BFf+YwUjVH
Gb8/XMyxzjZMH52mWlJ4Mb8jx8c7+VIxDQNa/Vik3Ew93ujx6eSt2LwZaBzi+qeu
hCm0VO0+rn5xSocLJEdjDeLqEzDg7D3qw/v7ew1YtosBjxB7U3eq82wScru81h6e
FFPJi2Z8NBYTqy3pTwnvxWY7XPuKc4bYYvi9Q9nfa2HuWHSfctqSTzMWIJUxpCSd
1vqQLyVRGJdauDwctbCUO+8x6rg+3RfdMB9LAkfzIuuiT40wXPhX6FRmK19VwfLN
Zt8G0KRIF9c2KvS3ATHC1RRda/hZ+PmEQSmv6hwSiAGmOnE2n0OYsOPgq+9UW4Bb
WcuFkeeR2fu87/rhhxwScod6NVqF9G5nZa9h7v//v2SFroctrraX6RFOVE6DlcL2
MW+br2JE/4gf8L7C6Azs4UhJLw3incOc52zk10K4Ig5NTOVbb6Ll6uVWckXvF48D
jbE4WfOYRMoAm0IQvorRP4vEr2Y3MkDxkhDv+X29/yKSP5nZrUDaN1Su9XYKq2ow
w5Ug9xzj1Wo6IlkqAo9t5GfXZJ1odbSuvLEZGpty1RAY3S7yVOxO0FEQeMa7/5JF
xk9pvKtTy6fdyjZ4np+X9jgKnaEh17Ttcwk4sEHlxYifZPAZwqBf/oDQjKSg9apH
udAB6qVQT9w9l3zIwVSzmKXk9Oq4S3Y8SRr6Jj+If8o0Om408wZXMTc4ngCYIhe+
sNX3buTF1k8RvuGnVVltjw8Iio/g0UuWxjVWGDSrqB3QqucZP9oH1p+TcsnxiKrA
gzFaCxfmh694DM5YfpgCXxZ32mqUdBGvI/ybz6YTuMCxPR2QB3cbdSk9SJ1saHQt
99+dps/hfqEmfzM3Z7Bet2lkpyjGi/aUduySheDKi0Oa/oEKLozGQ1kNot4MfymP
1C0XvucKXYPffJYf9vUVEMc+gV1zLtqLXxViHCD+VkEE7vdxY1GIIL6MDwHQnyOD
b7xeD+EGCaMUjx4B/+vuL99jDvdwLs3Bziul4dWV5tQ4YRmVdZdOnYwWS83r9eBs
7YuqdNQCUyp+4E+Qcv1FkZrdDxr/mC074YQ3mjq/FzCVIDnhQGTFIzg4pVjmWdng
jZoY69jpls6gbqnN3RhfEPPBOqO631IhoWciYm2Yf1MI7DzuKUvZ6+YBc64yi1wX
L4e3OTC4K2OzXtWtgxbHEhL8utRjhF0eMg3s77UB5yt/FtBmafwIKr4LUn138M2W
g19NoddreRBBsO1g/V5URH4tMCp4eNxePZ0Tuy0GvorhBUt1LCyqRVqM3hbb8bmX
ySPSEOFFuc0J83886aBFIT4izx4Po5JgMoGQ1Om9Kds75b3arZvihr/Cs8SZRS+u
nKDdq278RgzCoAtAeUN/XlYVr46DGfor+Tgb2kGJHR4MjuCuxlou2pfW/Zi34hvq
I63eqyy17AXQpDR6z1lh7LG0bNpocDeM60LNgRPTjp+xRmaIKukxxN0LMdSVvFNF
wHeZtG4qfFdS/PEPk9XtAtSTA6fwzbbKz3zXWyskcWMpSanSd6PwHyaVu8xqDvuB
BVRLwA3KCEQp2iSB7Q1Oq1H7/40Or6cowCxfzyoNxkUk4ZnfMGaB5jR06cZyiMBV
Gr+qmG/LAgRmVSgrmKtbYmOf+13dHq7RkR3ppzylDMwDq200jAZVWFl1lN8gfXbD
DER5m39SJK04PmMs2yqh5o9xJ4ZLYUfa1dzf7uReiCbeWWHJHCBR0amr2Z0NgPLP
ksaJS8iSgNyQZO/kgy+xgk34tiBUbo7QGUb2hQxTednDlPMB+HFa6Uw0yXCprsej
qSLj+4vT6xC9yHk4DZ2EmzJXIUtaBkU2vBCU+AwLDROpHKbFLXoJLx1gBj2RFYzH
9M1EvSXKXWYwhguzNIQqE8ksoocQ7cWyKgm9EBlO17DWwCA7r81KRgnEUBF2Wv5q
zLy9gXbNJTwk2l5QorOgcGRVXd5Lri3ZjgPPjBOYLv8bM/7B9HQhthNp4XuzMgDd
mAv9Kd+/rnktiFOMWHwDNWu+Dhno8wD9BN4DZySG8qmmAgoAiyXMUFb69ihTzMqW
KdZBiawNR1RHqbdWxxIL7I9qFJLa2mRq2EY3rpggfMtlX7DD/0890nryp8QVeZmQ
E8e98LZCEsusiFxdWt3Xbbxd9KAgCWVu1KCMxuWLBaFAz5OPfovh+qfhvRkiq/si
LBc1M3ANuFnAjhB1fdP3kbEjgTwlvWDzCqGvmYhVU/Fq+SD+ymI839IbAyJ1H/vU
vVhABh3HckG9y3S+njD1PO1vlbnKUDExMF6YrfpXcn3eTKQ1VZKxQNPlLe9z6qsu
zoYOFtPBdUqHLy4+BKCQUVi2GEP+Ov+o+eWhfNR7JrkwsvNwkFvzn43YGhuIwQs7
AkkbMyfxTiavN8ue+XBtF9XBH2TZ+nG4xdjlPR/J89VCYngqtxzDGiGXTVIiobXr
oEQry3SWeGC/Ty391AsqCP+g53j+EE0j9Fbmg4SxihA7hLFYyZuPTBERIqQm7QdV
nr0L+HhK3ndV/P0AcvqFIF9OO3BwYgHyCxc5BSvBiREBRqQG/rCcweYHVQxHKcOG
2pnjOmiz39AZGA2vsRLGEaUGjoDmaUKmzx/jSJu9iEqlI7O+Nj8XhNrVMYYVTFnS
U8rWTlACJzdu1mWpWSuMRn31F+QIp28GPbb7EWeG1UlvyJzsxIpI+7hLK7F+N08y
3UPHoQF6ZGP3y3iQe1yqcydqOzZHNFp9x727WSjY/fPAVjXjUWxVWBGvhIvNYmzD
zQBMOOR2/r16ZrGyiA6YNgwH59BYB24ucSlvV9kktX4IstXcwYndVw8EnCDcRvqV
SOy1GcLK/yLnrERPy4rGyhnWHko3whdOGZaX1/YsVzKbsQEuAi7E4EC+SMyfJFQj
fUX0p+aAlWD+rVgMPnTuEYVNPvkgXP4KCjivmJOE9NyamexEYq/3lyonFNAEWmzj
V6c5+YBTbAJWURUblSze6e+Glb8ord0Er3V92lXCYjNUnpXGIOJWhYaQco65T1v4
yAYXXmVD5c6hastXjmm1x3GbwMQco4iuVtiWjqeDnxlVvBafmN3g9WPss6xBn93R
0He1gcD2/ZMAGHY5vABm/mUu73v3Hi8EJ8rWjJgZUFc1O6+u+g8oATwCf1co4Zuo
cDpo3MbuAIJzHl5MnelSdBu4uP78AlP5WnB71UwQ6pd3Qhc1YOM5kIo7MI/MUKwe
DJDELfwcWDSu16/YLBjXw6dyl42jF97GQ05+quaBWSaO6fJjqx4aUdA7jsVr5Ykk
IVL4mLgwCfFnsN45H7EUyeMiTdM6xP4TmbOtOJMcJO4rP4X4HXLqzdKRK5masvq3
NVaIQXTf4Ng7zIoWglnDx54jl/1jC2CkK7revjFCzudde9OBYFL7aylycE4btkPb
8yeKfhfNKuvNG5Uo0ICvHACMRyVBQq6wTTOrTj6LzySvPXZkwpBoexadJ55vsD4x
cWlKIwP2gtPIQ8lW34oSMdRh2iSs2NMY961qpePmPu6xqbNcnFmajbgnArgV3XR7
ury+9Lm2VLJ/6pXnAFxZK2Lfc95NKz1xBPwnCkaCs7EDD+tjQbQV7vS5ioOj/dqX
w2vt/BYQka0+Sw+nOa/H52hQu7qCdecZ8stkxzkOafJm5FdI1kg/+3kpgD5zePgs
Gh3+25skQ5n7wRv/v48f0TDefR+j4zqh2uTjFx0C1h069y5pCyP8W4TU5kOa6TZD
oBfu5hWSpCxrjvA3AK+aoMJPIe/1cx10+ODug3O3fh7SkLLbU2bwBDNa9FChF17H
D6pEyjSokXABQ47E7cH8Uoo7r3CG4PFzuGoj2PttjpDZ+y5XEsC5fZ45kM1dOWRj
AB8w9vHESim4GuQFvyJufAXGhBFOEyyAQNxvpnLHhj6wz+xWOpr+6mqIw9IubzZD
SobnspZGG4z2BNcRngbQzrB57A1ExnyTuOR4X8ZXLRz9Wtd2+7+rujWpf4v9YZ30
etF6DOMUCBjiPy5pwnBrJF/8iZfJg6f7USlHaBlzODuhA80MTS0d1jwkgW53NRz9
yg25mmD78W9LjbUor6blAhjCCsLmoAUGpIagN9OP1YI9j45fpDTXvpMrLEGLVgFr
oQcutXBy8MpFOdiUcT5d5jUBiluDezuTte5Svr5NjzBSfVyRQ66DJYuCeuoa1ZXx
x6Lk4UPr6qmBb1NcjvpeBK7XUAcVlzi9opAiPkBdcBk+o/av8XkOFmnYJRAGXMvF
66yr0ATe3Fz4jU1SR+vzp+gpMLdm1LtlYGnPP2pMhq7Q7t+2pAS38snyw+y9vvuH
SLLLcZPpyeGptIai0WW/gz1aICOu83NKv0GKFOYxNrTajYi5d6833xlKmiHiakCt
ZjhYmfDCCh4HX6XmkbGpts3jCEyeh0IzV0jmCOJvWx2EV2ukznZS6+hshDDZsu4d
LhQT18KbxcARzu0OujKUvJaJHwU5zwcw3UxnKLtR9CmNZMmxR6gQBlh39xSvw7eQ
SaHnxX3i8otYRmmU23+2G7T1sXv7p36NBLczn+oM4eQSWNp3Y32tbA8WfYeIyc2N
YWIL5BqWsk6W4I4V4xOUrPMzsyvUwj1ZpPWeuZ5ZUJDcQtHcWNPbbAsec64lweHU
Yqs3PXsaaJvUp/mDyGcu195sN5OBlgBp43t44itYaKJjZBD6hR2apHkV71/gqSuF
6dT5WZ3luexuyTwKkyYJQhYx1yUknG2eJ0w9/gwPdn9kkz/BIkolMYdtGv/qMYXl
297jSfmpEQRz41H/ZlWORy9I6Ce51D7ypux8mJuKnjizPEbyOH3TcOzxYAk16j43
wfwLMB9pGQp3aRVxeQSPkcOdwqMPJRroSCB5hGpf54FXe4Ib2KzwUiVZBXisecvO
BsfplwnrU6hrxr6JQa4XQBkx/UU0QCC7VnlBIWYo0/tXsV+uEidQ35IggY/7hugJ
b/yXtYg4sul7Zch8qEooXO2O4e8qMUFujsEJIKkVKoCWPJI4yoX2yQRcA8m/yxE4
jhF1vyw4YzKszDxty9523iuRvdzUZfEqJr5O/ZdvhHfNka9SMSKLt+uBFXKq84X6
ZMonh9cwdUp7x2nc8XTws7JsMXUc3N0xszU/biyXWMBZYCMc6niS0jIxXEBoaAVe
PeBIHGS9iJuQSkEwQ2RFQmOtXtBIjPHQrUoU2X92ierZJ3GDSlhZ2W8wKrtEKOlk
N5iOgceHwebwWK5c4HquO/dUhc1484zkS5HLrdc5XmUKfVKX9LcpmozS+g+BM1jz
zk3nSl9jZYPs7JJAoA2gikQG9r22+1AV971wQnLcJVr3APvc4dXQqrehvc9niPfL
MkeRhvp6LsqL9iVSxLg+YW2qaX3ZjjCbhKGCJj1n06ETbXxpDua6plUCW/KTQAvG
Q1/DA+i21WIS7XKYeIUX8nrmaA7TNjFvxdERWlmMGk673Uv+XURz1aAFMDg3JRzl
6HkAku/O8533MxdMf1R67ihO2g/xTXafaTChmTgCmAKOmPLUp52MQXpEGPFN2OCf
XkO8hVxQJPHxwE0iiTY3yVaoQ/vIWXbAwBFlmefDBOlPLhZbslRphKgp6UdF+P+z
UXFwxDfA6pGdWnIL+DqK1GeMJW63dQ2tOCbRXdX+BSUQNpUzllnqRVGO1muj+gqQ
KatPgtCu3gedfqFoNFYdTedTsTWLF78r+g2oNN/LKTtEbBRep9Pql037ftYqFmjc
4uZ9Inkav9Dqs6PFP9s9f+xskO3YJXjy5CrFi5Q9RtgX6wm+lioOMhSvcHfy5tsa
woWjuG5Aa5sO4y/ArGNdd/NLQffwehBHOwBRsDyh6udiHb6EWa4MRUob+KHcDKvY
mrJyVNaxAfcn0DuA8niGH0khvP/eVNRkq8v6OFDJKdmCfYiCu3wiDKR/FEpmedoT
K/8qbN0e7EL4zN9YIX9blUTUmHW0ZblnxBrKfrKUN9n1kM2DR43ywLH/VdfzgsdN
2uomMwpztu/ww80RLuQFv13MdtkZCfxEBRf6BhFXP8EAZ/5kgiSatd1rOZTA2AkB
UCXRqz77naBXaKFJxHwvonsrFh1CeN3a9saV2KqnQfIboiFfdab1Gjy8vg/bG4pe
rvB4kHHj63/P9pM8F+1cQZJdjjxTgRDywH5XuooAhdCqyfFOwKKphPU0T7SDwypR
YmOePqqz+ku01dtAlhGyAE0hue+mMPg/Y0iTm7zKix+Nn4u5z7xoc47t78AnN6FZ
KgPJYMVUU3YKb89tEQ0wd5WPHcwWjlxIZbWyVNwNGfVRQb4fSH9zKczMav5RnnsR
HgrrWjokxCDZxf7WDqr+8jut0jOkoul44G/dTbjEwuJ0nnU8ULMmEDFOOulZ0qLt
GjH7dWklksuNkYGB6ngKiIfOAN+bXnujD0Woi282YI0OrN/WI4i6xfxkWQnUW7fl
1pqDVDl/UaU0gc/HvwqGV1n2G0BuVW+NBTZhHm8VP3nPtX+9offKE20qvARxCGys
Z30UYClGr2l7bbvzJUT9tcg65CmKLorTU6rGYCCz2ymjGBi4+Ikd2vkBkss7ZxrZ
9KyO2dqZHZ1b1xCY20tQH7AbCZXoV+wnDAhtdslD8ZEaeLgIUAag2jD+WF4Elp5n
Gu2VPUAi8gV4rnJC+PBL2NbdN282mQB9kLCrV7f+xWrs5/ezKJyBieM/ZMKHf4TW
/HDoqA6QruxpyZC/OnR9zyDbF/5lOJT4Cm042PYVm8xROt/yp+XfDHAcbjO3aYee
bkuMg0CUqRH22Iu4LEC5loIEma8X2lf+4MPaZjLNa1KOOnHKMSSVV6CcpdbgkIfw
NKiKjpaqdNS3E4P8eAZJNXsWEFkSF+b8M6tn9rTFR09CUlzU1exElwz9vSsbBeRI
GCTm80rLzUfUKeMggCAntfWNw/+nsAPdTToeMY3jN5J3cavWOfNNotlAj4s+RuON
lNyBwTJBESqDxaL6ebD9TscgCFS3QFy+Eyo6h32DKyV2d3e+tUWwBMKLdangH58X
BQ0mEv4rvC+aW2IZO4QgdWmJe9NCqapkIKH3jXn4Vku18nJ3CdhZMAgtSTaSG+tq
xaHAo719EQBqQlndV4c/ks5+ZrxWlv34RLyrsPxytYu4JG6zQwPQ1xVKvo1tBCC9
i7KdQS0pqEg+UCnwlJJCO4QC5cl+GR/YZ1kyaP3y80ADz+aFQfFIQUePtHFMPqeO
3tOtsjJNNV7PKXa4J0GKCRQDNvSg3MWwbkj6GJ6n5yhxB+ALtUZ4wHtb5U48dYKb
YzI2TG62HHPAdXEwRRcbJHY8cNL+ppFfCCq2/1p8UjBFJ++laVK/4NkqlWaMtcYz
Xm1TIALc/+i7OGhtO/TrUtxxli4PjCZhVBH20d8+kwOjMEuPukuKir0m3hv9+VRV
RUJ/EMAAfsk6d7f2jmVQnKoZ3aScNE6j8pzSKEqloB+w1YHAIL7LR6rn+Wx3Fa9q
H6ERl5rY53TRMGeYHpy9/e9HyDMd28eozGrq7vukNqtfKBJ5cKn3C4ypXSfxSJVc
0FKGGfMVy/A4i0BJQ1ifeVg+vfuGfTmJtTPeZsKxeqtgYUfQRcg6PczBr3KLqm7X
Nnqj0TK90FTBFuqDpq9d9WGGTMXSJEds8pWay9afdYKcFhZlFTMxFrVHw+KKd5Zh
qN7BCBzXb1Pp57tAsFaY/E0BmKuMi33Ay2reOpCND/SMqUXPQBHhnUC2iMAPJBS1
GRVMuG0CVFK8jsv6DwRkfLGN1sY8HJRSg+X1BBb91Un4PW+gSFRl+vUlsKs9BOgB
hXS5XdqlCeM7+pI9Atnas5RxGEXiFA7SIBBMXNpLRn6vMrxTXYEUAhFFpAXn7PBL
DuNkn2lzp+rq13QckXfx2QyqEAHOlTE8urS5Uy6CFgEmMGhQ7dlQmCZ7pdD76V6A
LJdFRoI+l+uuskarIqc/VOXPpR8/z+MMIU/XcTmWFOf1/tuj+z4SfiIX5AOx5ZP5
0bsxhXQlZkiJ0tx6Z6D7trOpyet7Uk7qtWqJ4hd8wrBxLrjDJ0zGmCwqp1xu8k0i
PXOI6xw8iHat5MbAuH+XU2NlyMBq8UCYZP3tfxYqIcvXjTxUWU/7VbXPPcspo2ye
JY5sWSmynu4jAbfW63bEu6oRmdcXsdleT0ZswERPnTLMiqAlJwDqynXSFoYQwMVo
IymxIgOhy/d62NBBqaAoa2XX9DQejs115LDGYhM6Y9AZiKk19QkCf8WqIj/mtCcA
u1jRTQXydvxqNXatryfCvq+XehG1n+aVmCcLBGQg77BbDQnH8H6DS07kBynj+Eef
Edh0nh+pi/29q6D1D2C80gjZEDSCxGQAVrAIEGjZaz51rtB11+YkFa9mnjRNuZ5D
DR92jk6XvEPs1LmFO9oZVnRO1lFPyn3PsyVW350Q1nbXfVKx8Ch2ThuckfhIYuv3
8eJf9bqCc9YFB0R1vXAJorEWblG2SL8z81LzhT2dTt2Zk6nPbtWTmF89iUH5RKzs
0qMTwt+uMEZVL9zLEOeyPvaJr5knk9sr0F7lAZUxGGBR/NsaVhInI4niLSVpn4ei
EBfFCtjBpZdBVDYDLF7IvSm1/BxBf85dQgfEDZKsA6rzB1ciTDZBhxD17ShK1jjR
3/5YVY4+8LJLcv6htDFAg06aYhghHo2fmD1/cQv4dbqOP9bsZE9iTap0ft+HYe9H
7YZZzl728a3mZYMGKK8j9bKXeDoHM/zJgklvi3/iYLgXN19EqG+6uNnFgaHzdkkR
aPGXbbEv8+gEkTQaYvrcBXHHoCR2rYyi7EfYi7jdSoNtN/6u++6S4GtEqaHd+Yog
bYIUszcDx/zRxdRSOJsxhbrC61yPoje2N7L68AARVcpRdJW7ZuC5W4u+1vrSlxo6
6d5uwBfhpD0POTCulCKwNMs2ChMRxQZFGaVwalEjlYdO1u4sBgYzhuZgKXuUlGg6
jGbR94+lCES211Bx0e7U2PxPUyi1gK2wOrql5jPjqqAYzcOfS+aLLMxZp5wo9vN8
tBdG9cnl+0xA7oJfHQNRVc9isfx0KE7rEdIdGkybfYWiRrSfpz77akBAaWTcEiQr
LCIKQHniRNeyPRiLk2tY68qfP1jTQx0leb8fdY+2eAlW2hcrRolk0eopB9xaiezE
f8LXhANKY01T9DNIWW5xswelW9MPQ2lBnh77zVBIcMbEkrzGxa7fWr1orDQbRQip
nWmJoaSs8M2mhuX5tJspUAa9WM1aBC0pCzsl/MX4mWqJ4o4UrBeuVEYyCCSN7pXt
Js62R9W7Z1+14AmeH1BZHnE/4pfcyk280kUpqLHVlLpZdpEoQjj8Z0P2nfZ4xdiE
3s9i2C840jXYl8MzpWta6gx3W9BsRg1l+Mna70YanVNH84l4QezTbguAY3JV1xGO
IFnhv8dugF3PB4FnHJae+GBknA9Ahap+fNCA/33zfgjJKAhSKF9KVLmtthJLFJ5F
5/eHtjvbfrBYOKGE62+fsogVn96vqBU0lchkw0wVje9o3I6dvlLNyuXrqmB9DTvk
PAaKjETy+4Evc8v9SFuvVaBOWD4Pg2QKJWVfIPrC+XujK+lRztKBUBgxCSs7aSX3
VgoHToXxghoRQ93ygoXWYez20snYGGwCu8MsdiUxAqT/T1vj+xZEZg1Ihu2wFDYJ
hdyRMLemvfPNoNy0kIIm6G6HxUOkRhgKgqjXV9cpPB3fILIdvk+o+Sy5geabJE9M
bQL84S6LbNCUvFzF3ppvmUiYFJl9yqx7PEyLTYPqWCjtrG1KyVN7Yc9NNlKY+ETo
ECUE+0EuYTBcdNStInvWHE+CBQ3t1y0CwkTSqWLoU4DbCRNO5cE4fQs8d8WvL93N
S8P3ehm+Hh2XQkhRzDhst3jfJ1lDMzbs4rmSV1BN1SBcdKM4dEMWcHAxyUjeSduG
eIh1T0g39Lgl+KB5UijDCy+dKww3nKjs9Z1RFafBJLWef/kx8JZSA+bGlo8kNRNJ
MZlpeVf+o22fjZhRJwm1/Vrmuvif6Xl++H/ybS/ZBc5hvot+L4jvmh8pssrZsiUF
omN3VZy80GiLPb2djIyScxnD8KD2yl13bWfJYtY8RAkDpXCVbY2xRGngWLXWBbbb
F8+5EXge1VWCcMIfDRiVg3vJrxcbqY3pFRQseBInm2kxKHUWjLts2btFaATmxea4
x1hqU763q7nO9iVKTTCuSkm+xhpNd7aO1KRYfRdp6s9ot7CymFxnIYc6XeF7a++e
5PGhwokFgf/rKocAWKgKcrAjwE0+jva25aPecITF4nfDPa/6DOxGDLkbNwVPnetS
q0U1KdXvp/W/Xv6q7cpgVJpE/sPIqL7IkeEllkTQXN0GS9FmjMXEfwXih47N/kep
0dh6hYej8V65Au9iX0GF7ZUnf5J5UVfvTN3QzExePsXEAiznwOkbAgaqbmOSJ3JS
lTxkLBKNjAxJz/dqrGijBRj+9mXES2/b+i1uUfuS+kc528bioVxWyJWU7wh2Y74t
SeKHjkK18o8oiK1/h7GIZTyZ8vUbu9KwDDrSd85utW8SqmRCktlfCrM+FOu1D5lO
7fEFknk/bGQI+t/LElMxOdc675Ht+n458oU5+gWHD+8epsHSWdg+1Ydfxrdp9v24
oYTe0nlUxO3aWevXwJHi51nXeP1S/raAsWit3T7zDPjCzKLiR08lSLKeIX/MMgwg
CjbPqjlLW0tBxZN5bgEOtnIjVSsvCZtYdUc0I5qNkYP4obWL/lnFkMJ04VfZLCtD
ivJHnBMnMuJwu+MiEiO0f9pm0/QGIOqzW6Jhzd00298W2hatvb+T9+fxHHcdkdYL
Rh3Xek78c98GBb0V5ROTvImJrkS4P7BMsk5CTqzusHI9mUkgVAb3Vr9W7Z9V6v7H
gmGSXo0M9XdAMcq+VjQ5Qy1aNR0B8qT0Abzw/lj277rFr+uMk3XnbzmpNTlqi0RM
r8HVstwuVAI+Vl0go5ZbZ4qPTmrBpLN6DWITbfJC84+U7jR7nTAEMBHeHcC6RE76
X6AwssBlzCmnRPXwEhKKevPWGyl8uDOc88WASfXoq5HPA5XoG3AG+jWoPrfFNwY8
FrPuySQC7xyFLHL2CgLGnsIcS87GxkUaUoqFEZAqA0GaLTx06qFbCmas/shFdxke
rospA/uGJHv2kWCDuQ6dkFjkVVNyXqijLAq15VFHBNhKJRJOXUFX/e8REdcL1nsT
IcuVEnfYaSYuUiD9lVT0TqaJOJBgC0E0WvFN4+XKv9oNkqZmt9uMk2LHtnS5RtAL
ma46VFns6UeEx8PYE2FZDhQpDfFJGW73hWRmRmfJE4yJAGpT4yQeHguj8FY+4Ucl
mr3t1704cToa1BVOH6WCaf6U+inLJp2TOz3nMsGiMT6SCf+tV3vjF9QYuXuuELVj
hf0YeVyjwYEHmbgEJqTcxe5jL70QdoO0lz3qteaC6U0QbcdMZrc7oP6QzrNgTOVp
TNeXUScVPlgT78+sgkLtFelH2idhWnB7rib/6Ed2h2L8RSSfAwtmfuN37xak5XN0
VPmf1jASuftMyEl2ziITDySKoVTvj84F0CQYsxKgJYopdNCZuWUyGoPFThLT32jG
GO36D8l+jMCdTHQt47BSIEY9RDxYvhC5baNPgTikuHVb99/zvuMUDdq804wjgStW
XIqPun8UmeRN2N4q2+k+63eTOqPmGiZwnn47S032hqwTWJuPp1kJSWBnFk/++s3a
4HNRU5yDhKASZqGdXiljuCgjJUSKvr7V8jPDtbl5vrOW0dBPSZvpZ9PkrmTJkfGN
hnrx6r8KrcgDlaSIydoVbNol7nvOcbUTRuBDC6b7qZY9HpR5WzfwQl2VYjxfpSCk
6uYsoTNhNAuJvpFhWck9xdpBmOQ1DmF9w0od4Go7AKjViBjqo94lRwd9YE1RC+vc
YPUBybFp0sppDkf+W1JSwCx/xIewhifyfdYEw3NXotZvCLN/nmAUFH1KQ6lYCMc/
4ugwTVyhe3yNWIyYfbmg9+/QM6kWe+4BgdxKAOPhjh5dZMU1CRIVVCpMlyvY8fim
13CILi6uU2juYe5wGpjz2RsxnE2IgrDwi/4dxVrrJHCVUavglxdvyrIskJv8+yIc
gN8UlmH5eiS9HuoS4q4IWU51q3vgnKjiKlA9z25LW8CJEQh2hfOcxho8GONQ1Q0x
Krop7THh/10uR3Jf3PTj2zsfMBMhG5IGmk5aLDklypdeL2oEjALzGuYLRLmbs/hK
/w0HmYbVlxwcLTXjNETRyIF7Q+10VFuPBqz2gpQziOoRZ4hdMcn9s0Slmw1KYENg
83I+1OihdxC+wBa7A+4CRtWD0PBgHf36QjRyK1uogjoiHdcVg4j/LzmyUeAOE4mF
sLEmwosrvM+KhWdPI3AQpaYcOy2D3ZAysMkUWQLN7srFOnBGjpzHWJtryrP81cDn
GQaZ8EB2ACoBKCJ3ob6nIzCeKAhf6lD1z5meAf6q7L20mbqWu0PlGvmCFgTZ8US0
CmaamqpubN0kXwRuswlrMHtXx6+SMBxVqyhkvHOmz3R9BdkHyPJcJCF48hCh9g+3
+LU56wCMY5rEHS+qLwia0rdUeDr82Ztl5pY/mQzkgUJ6pWUKBJd/UuadBj8aBp9b
Wfs8+pmDD5ykwbfd2O1vwDKOLHovy7gwHkhRipaxDrIUwV1EIyf94T5x/v0/1Erf
Xhtc8DfIF1T8Wg9yLXrAZFCvYAkeJ+/cycGgEdFjnakJN5+EL809l7scfU785kDE
cveWn21hPa528afD5FHJ/KYRS3hd8ePS4XCS14WnQTuhMmkk94/zjGcy9c4fLSHu
MMVMyvRwY7ar3jDP1fi6+A+DFrRwPdSjZJcbebF+ymOktx7fRgLXCJeT+qXqONX/
GMl3KygGrf2Yr0aKa0H0K3GAvLN/+0THqA3osyMahWOqQyU+M7JfCUgxKUcht5/S
yJsk7ARpE9Umbb9U+ndEMmk3v/d7u+lnZDDQceBK1qDbaC+NpVMR0S0q2oceoEeD
yU2o0Aj9WXLK/5p/qRXr+yGoJDSh8KQ0NvLUsHruffSE5ov+tDC1/yPjRHx3c+lY
te0CinXmcSEiYXDgR7thLNJ4a8k0IUxUBGmfJXjquF24yrsS74FiqPyfmHsVdJdi
PtK9xcvAVrtIwTHdQPeT+/X8hecCALUP7RAqP2leWrfk3ePoLbKoqK5Nij/6iDH7
FKEMEfw241pZbMStAEcY0zZZRV4293TP3dLayRc1luZjq0s7cdmwVXpbgQT0lV80
78zzjHb0/n+OZzVg/f1e/JXaYlbSrjN9kzJLdAnjkToMFGI6tcs4gY/bBqUOtUY8
WUnjQJ9IU3CD1ZZgPpZUiPL9UuCtOHxZRds4zAxoXnPsr2744kWtAHlGALy+8JBn
X9NXIZeeDAWlUUv7hSSipIWr03Z2uPufjHc60B30f6Rcs/fESQTzpjcemnrA8WwX
iRmLFQAzvDQ0y29JayUXqkJYW2LCLHsFAaVmcwwRWL+9AdTlbKvz1iFCn0GZjASO
YZHTahb11+AxInr7gl3bljZiv+/iQ4/McN2bUDmmF7PcTcZJVC78dSOIttYHggYA
EI7vF/BGk8E3LuHWhFa6FYPrE1SYyJxaEiqVp6K7A0NRqEp/Y14vW7MoRw6Ld+Lv
myv5mrjSk/6mm86n0LkOlGVAR7jjtUF2FeetEC3QpX3eYKWqMhxkZXpOby1qgRDM
15Ue9lStTl0BoHTfj/57X12IatY4XYn+KFsKB6HMXPU0fAjWY4grYJ670PswzPWH
M5u5fxgntikSQK9COvFK2vPocPZSLerPbSp384VWdvkEPsLtJNuC24LsfQHcgxwd
tpbmoW90O5WdqjE0XUilfqmTnllD8y60v4yJ3/2uXpqPBTCNuar0mNiRhpGT3Vms
48E/GkD8Yp2Gqg/4zRrYbeaqPvX+8cwkBjUFOO/eiMAAL6yAIJQjY7cD152cmPOf
4x4/5Zq9WbVMWLYVAbQ/Om4YmvEpIKYCvCc3vaoHMx2hfKZZv7nomN6XVgnCzsd/
oEjse6CExK5/gye3SjyGogPwg3K8OjumuXim3RvNXIuieFkNb61bSfKL+a60IEE7
JJorwCGnBtsJFh3WQCNfVVknI9GS78d2272EBzGzaqrbMgFyJTvXn0/KkXwCRqEg
Vewx4xbsumeeWkJmrjFCQ0BDKdpG0kqCcgsKswF+yqz2J89W0jtJYC6xrTPBoxoW
cGAn03nzJTlS+NKDm9mIDmNxZ18wjK/6Tf8pPhOkvOyfhYQ4nZ3mvLs9rTsgSbRU
gLiAHduK5ZYbhUHHyIJCiFNF1vHl2WevuZOynSfbV8VCvD0gO4gDTH8vWcb5EloW
S09Km/GlMHFA9LhHSdf1MIO9EbTAIPQ7DQk6x87t+094JH+m9BFJVRaIzAeawV+B
x5SDqgm6n4oKdSqPs5aAEVa2jui45W4y1Y0LdTqZBV3oRs6mDBFy15cCy7SDvmBm
iAwOAEh6eTcGfKYjuUWhcPJDyUReyhBxgOLtJe3g4z+EhKOmwvjOqbOUW9p8000P
jqpZy6iXT4axyNWhUH3WhVCUCpdNwijcXKSlC2I8+iVDVWtsKLzbAgVjg87/GIAE
1fg7Bl/Wj3ahMf1gvZwkqyKkrxSP61fOlwoWcVKOPdYlqqxcYYAAP8QmuvHGAC0T
7AzIeQjIfrKYoZkbnOYdcCWtbLrEoocluDwN0YNo4PIOxNwGE3UVsZAiJgVJcFL3
ckQMTWp8PJjrCNXdY+zLMjGmcPjF4w50Ku1y/bnnDsLpR1cN919gQiKKjmpAEN64
YkDsa/xD3kXAqi39Lv0OsV3ZwAnNI2iRhVEXpC/pwuY/GdDwVu8MGuZsVANqOjuL
unHFBj2MzOeNrX8YsqA4Wq2GXLOooIfaqtlPDITVD4q5flhOS1V7nDrE5vFMOVIO
0EZCmepe++M5PAd65KSpOyiGoB3igO/BpqLVk1Rup3iTjCZoGu3F6k5pgEpJJ22a
YcuvWfpg9Dvs4px1JXuw//JSFr2XhLTM/UJc0ivJT6DOU5p46cBFFc2jTMtNh32x
9lz1EBupOykVuznXlmTfyEbbocvp8F1CR9gUxn54OJaNYdGUCVK6g14QuCGJgz8O
NPrjCcAEvjQIDEO/bi3ne1skVVHLLYGn0Uu7s0+SQwFe6AjoHKsopkEeC+zk0iia
OS37PfrhLynd7BnTEzQaJEYYBSi5/KSgRNI+ycWSHPiVbO/PwyI6ke8EUnIbekjn
KCKoQBjIcIdUWUmeusj1X9BzyBRSCuRZj1epItAmxiqoOHTyTPy8ot+0jtRoSO+G
ddCw2FbytBfx6G4QFInGFsEOOZIqDQe2MvHhaDA1WqrvcUB2QDLQ656ST9t8tzV4
/D/MItK9Ww5xFBq+EtpAN5oCMF9epK0vDjND4cJo4CwKVcdzqr1oQLcnM11XDl9S
kjXsx7q43oDcZ4GerN4luWb8rN5IpJjc26akRl3pl5jAWh/9OvqkNE77G2uc97kO
xfL5a3maSa3CxIWc7qneAYzzmKlsx9UTwMFWfVRNb1TRwBfbUUGjuNZDzcYEg1yz
l9H4giqCwkPpAJS8j5C62Ks+NFKkEG1F9EfV8SaptSVwRsf+0O18qCRa4JT9b3XD
975Cgyn209YvXrsGYwp8+s9W0xCoctAWm4BUxpW7b35gwlTeGRZMobrWL34gK7Zh
RHx2cnRbx7zMmzAtnDSfsLQbc70zvPqsUtGWR4jL20n8joVf5SsNox1/J9Ssjfl1
UKNuQwAAmU36OcXt0uQeMJK+KVLKc+dliE4U5smPi2FTHCstzAGICemkZ4ggVf+N
ZJmpuV6USKuPGieFArdIukLGBFNM9HxEDzndftpI3rtEuEtvBgcAnYwQIuOLR38u
dhClGYVneMe10fedeWFVXXn9OhGhZ7tXk+E+qtwEQc/kBl5fyF2M+9/s/RWMKPu4
Rgwc8sv2YU14COCFRizjry/2I25oU0fmAtWgzxezC6lyGy4GaYATsPoP5HZH/Vnr
P/3OFOG5B5z80MLjpmLlj/YxPEjaOKdoV0P2bnRv9k+8VmhfRU3Zx7LPSrqhzPw0
o0FmjXelvl6nXsTiNLky3NgRIyD+jDkxm+44GiM0obTNdoJfm95f0KhhfXvICSO9
FwNJzG8P7YIOTENUmROaGHOt6Fv9Ls99vQkxOKTGXqHQ1umuFYuhdAa6++7I74ZP
foU/Yk3ynXYix7RvGkEPQTmdGoAcIt2rz2QUvJKn6FUpuU6p0rljIHV+P2gwRutr
cG1fKw7NAVv3VOVjj0+ich5jlQmHCr+GPXGprgT1Dxnk/Sae3B4AFLJRs8u8Mzrr
FVx1OLsu5bz9GTNsEe+A7bGP5jWPJgKtdiMMPY0J5Vli0fJj9Q5SPOu/BnpzcwYb
7482wSV8ViP5n+bVGORLpHiIZAUdJUy/J+JZA943ry2Uby8VU3plC31W5086Qcho
UHqp15I066TqCbrlzr1c8BXSoWNg5t6q3hAxI9m3cSLxaW7xyDOh89FKGLSTS16w
jZhoJ2+Avauvyho8lBqHJDhYvlSNwNgXQq0MsxSGJBirYRX4JUT/dMV/NAgLKVlz
6Jx+VfZaBsLGmWov09lS3RlspkjUtfcPfuCkyu5KlczwxU8kIOD4MkgicuWcXehl
ZwzhdbfRX3FXeJUTsatnXlRz42ea4g56pKiZnnvojCxZkOEvvy9ZtXgJOnbfCZd9
LxuAruERfQTgPlTLdfal0fZWRHtq8y3atq+Equ/j9rOFFE3irSyP0DML6RRjr7tZ
YPiIWNp5namsBgcvSpeyx3noYEUJ6dB7YGDMqUM3gzAKmXBs6tC6Rr7atOUGRAAc
vHWWNT8ZMCJ75+QBmlWE6xRjONy4PZ04Tzb+EvnnRQFbhhMTWOriOMTKJwcHO6va
OUOqBKAySnUxzC4ytREw5KPNKi/SWDZ2bFMP9j+TRUWaX9JNPJBgJXKs8B9Y0IgD
zEaX09rg4Thk/O/SCJ3dUY2JneZmHkwsV9OHT1HsJO530xW9jzRVKBNh2JeE26Vk
+iUEFadYpScGri5a9qokhH0pJ1pS/lqmV/cVHxfTWWG97Ika1KDEkxByyHDEA6nJ
Frp+k05tGLajvmhgYLi63ZHHm89XrBO9a6zgUTdL3cSELvre46il+qrKkdGqQK4s
+xUkcRlq1WZhD3xAwm6K0ApIEcbxoyEF/GRCSHyeV7gte+QX/s1GCBzzSI2CwY+1
jANTQ4IH+3eFMqIcsVZ9yABNSGE/JTNT+qrUZWdnutoXlYqFsvBOtCxwx5eDOgRz
Y1oRI4NUnDn+etwKRbHPOHxvWqxaijaAaM9orkRyb2AvLNZZYS3IjZVL9lebDbvX
r+2nbkIi00kJitft7V5jlQb4nlM9h9vBg1ag1Gnv/IzloJPiOXz6KTCv0R92y0IW
Sl5TRl+54RKU/1Cxr4H1endg2DibD6bL85KES55IJNos0sh1/XcHXLVjOQRWSC01
qq7Xwr5Vwpb1eDLw3KpnOyjPf8MSG2OFoUcUaqHEMnvKDgkgToxaatry2Lk0egEw
6nH/E1ewPs+uSVFivFloUV4VQvW7s7LI4kqvbR8nyS5MDoDnSmWuTiL2uzghDuEp
P1C6OZbUW+8xg+LZNy9kk2aApe/aUKfOJOMgAKchyjCBs53JGg7sFnCL332EUtXz
xdvxPT+RNvjh04LxU7Fr2tzRBWPir8cV7aTEVfTr/XQy7EAioz5R3DWY58Alt0qu
PQ7mkFgNvZgNIPGlY+dAadGkbClYIWY8r9QzYPJe/SdwfZUXjYoFYJr6SGtG96my
DHURbtNWYc70Er95IdR8CZ6mpnZ/SitY+RJjDYpXAc2OSCytzFIdFXKExpvr+9Qq
NhGoTVZAMrBZ7WS8601HxnYxxlMNefOxMto69IZUvh9XiU7kfzo9eLf3phOkil2k
3r6F7t1C42F0xQ9r158tGqKaRe5poHf0g+n644TD2BHhxob/A8YvTF8dZWmVckyk
45KyFMemFcg8mm09hvAvC6Lozl4W8zPrs4estJ1JiS707/DdFE33l6fTqAUEJ96s
v4aROEAEvUzhHKVN8Sczy19x1EG8Fh7ATEo0vVb7uksoE4CbsODumwImtKk289lr
hOuXOzM5g3PAQsDE0btuX56MwBc8ZK1gFjx00hSDKmQxAIdi9LfdpmGBqEHUMGg4
ME7hbWhcX6dRQFsnLfOVuHXXIdo94DkVXjFgxnNltkSq09hylSqJKq6oEcSkI/wd
bAZasI4j3spM4Y+I/UUowSsFX9YZSVABpM0I/3o3nDTZIYhgqfIwxEtd2mmwnuMs
9W9FEZ/MG1UgwSlPrf9wxHCiX59UncBqQwA/6H6wq/+zyQqvbCN2nxv3+cRWw930
XnUPYVUMIUSAdh0H9b0A9K1DNO5ZVDIQrqfbYlVffjeUU7faYYHaygiiRpNCZNfe
bE+4PUwJeJnWr/lToDZxWQPKzo5TLTaCFocsUeike+IqBshVGzJt4aQS/xR69Keq
SWEyadBv5+TJWodhrzQ9qpDlLztwDJ5eWWIkQZp58z60h3hPTzCLm3i9iABJr/yM
BOmwopYS/qlFAqfkn+YaGaBDZvJDlcEn8PODD9jSjfP5v1lzEfM0u5tRdpebCkU+
T4S3cYfp6H8v7ezpYWz2kRQlMJdww0+cblXN1vXO9wtnoRmlZ2vV69beJI8mQb+H
QlrYvmuLRpfMYmh690x0Orbsj40t4ruYtKAfbDvRB1wbJ1JyNknXxjmF8UfMUeMx
opvfr/swiivJfQV+nLZtFmYS+vyYOn3Aw2mAQdhadNfuHNDabVuh5Uqn2UI1VYT0
JrghgGcm1ixlWqYFpzr7VBiGy/PCazcbxFWq8eRVVFJiiGT92OtWl092EX2qLRVS
CyzLRZE1vb8yUrA7tk0BfdzBgCF/y7jzEtlnvLGB0TUZPWuKAzDngofJEERTjuIL
2Tmde8wEP/YmqU3K894dFTizEDpaiSD3TA+7L00U03bKCTiYQKjfY+nw7eDEGhYi
Nh0IcA1NvLEDeUiYzsM2M5agao0i2W6bTCRUnHpLVLcLr4QSDhmsMpvQc66XmI1/
keoXKhUEITH1Z9fzBhFE1HF68Zq0BN84Y7IwGGF/I4x3WQnJaO/AOWuIj47JhVpL
KR9vDf60CP1tyljO5swISx1sVdYhLyfs81zjwxyCj1gM8Wg4+3akcLEH+63MKaHw
Qp7rCJdI7gQaEbsH1naMHyGdhuxIJ5t5ve23BI5hWgkC3QCAcEfKNr2eGCAYFPjL
Q/WuCofHSFYX5exnCt0jlZcsEXv2org8xbhkIqFKd9rDy473zORexg0JihFTBbit
vwdTBRdGEwSY+p3qfnUb7+JEW6vFwF6d2edT0lWpGIlLxwTCcgi8ISaB/kXAcOTa
Sp5wfLiPtMT63Am9/sSI2x8OZNTFaWSdScXE0l9uBEgpViGvrAUTziH8q+QBKlEv
eyj6rLhssw+6ewqHzHVYVx5bFeqDBmji3G+RFMfES1sQDiHdx6TtCnpFMbxeryRl
AV/Kmd6kVbSKjL4s+03dxO1fsqYH6PZTKshZZ+T4k69/LpSn98oMTKMd1/UfBdhV
yayIBSOGMiAbWOusI4gVGVLEqoh3b/0aKUxqJ6ApISU47V9cxJBHrL/ieIeH1tjl
jfdtG8M1tYi1py1qRFr6IOIk3eDicf/k7gRx+5DAn5UfE+PQBvw5iKMr74XQxGgY
vsY+XUXHFO5hsvu1FGnHtjFaBPrf4a1dvgsWsjk1VG5kWbP2y8HBxPfx6wDf0kIf
13fxxWLMuoQxj/gryMtJXHPPwPpxsamujvQbdCch3MiZm4YVIaO1puRjbVludjQP
zvKqmOxhfby6QnzbqdsLfuxP47O/GJTJsc2EtuvhvamO76T1cUI+WXGhgjV0JDeE
ms5Xxfymc9aWeXri8aEHCQGS0no3BVv6ouHJyFYTkErAMj+pGeWT42rXTsEPfcP8
Xh7xgs5ByYDLYk8BoVFExBxRdyaj9k6TwHJM+kDvDt9xDML0A35rYV11/TAfjO84
kzdoqgqPu9bhmjsTfsLJ8D4SEV1WLz4Hnz7o88ApfLBn5SHI17E5IAC/BlQFvf/d
UuE5bd4TEKp8ObXpimWQ+lwYH46hJSiVUaZovfkbBY1IVhnru8Lh0mycNuVy7mBd
+HVWCCOIV9yfHaLWWNl7D6YaWTDQceSu+9CV5AKFfpqag1VafXJ47OzKreE91Rrq
2KjjW9nq8NbyverKRM88/fId8O2S1+0Jsqa2VLH8Dp1c8mgyxlF7b15tPKvMhvn/
qfGOIFuxne9VaPEzpzxQF7lawu1IO8gsBmaefP79uz1rZ3nuw/hcCBgZit/nPChy
DqnDfykdcp2X3ksY3wqhasYZWmi2X3tgh4PQyAP/2SnvwvYAqGXr8uFQ4hQpN0tn
8QoUMEpSOfK1FR5bb1opfw31iTZxfhinZWJCqnVZH1lZr/esoS5Lo+yWNmH7yZmt
jcE3AhKEXVTh+rUIAOSlendgX8Lw3mOypBoeco9dR/XNbmqligU37dhwKMXBYLvN
AMjdPNg06qw6C+cMtlq0vY7n3PI6B277z7/j2BPPG7I73xH8rjgQ9Q28wHTl0R8I
1M0utPDuYNybOrgQCRqDgYsrHsg4oKmQScIszuX621G+r1hIMXji0u8IDOYKJi94
9JCved8De2+wEWKJExm3epQqmF6Xc85WaaJO46e8zUtmqS2aruHTcDRYYSG6Rm3p
IGLBwukVT4JtmrBvQuOXNp+vSiW7YduV8qRg1TwMlAgbXGDUz+2hBIffgS0vG56h
lywD8cjt3RLoFTylKKC/43ljYhBUECUsOR2clSmj7gTjm0cQ40YJE1KYh5ie625c
NXkYRS/SdLatHjDT9BH3C9ovG7N1vM9FBODnSgnTNYanz3jSpEl3gvhVz+BJH/wq
V3MJLTQobDP3CeUHmAvsmwOQ8V1OYfQMGZ06T1toH15wQB3W+n78FrtUCIS8e3lR
1NVPy1ekqYqugmNMMmO79eXAEu/G4SEOPEb7NDwJ1c5V2vGc4Us7RBNuGyBTEA9O
cWgNrEnppVkDkAX6tzcCBnspeWNYWqS50KpoMjURT6YwmQZx79AH+RwT9YU9lnN3
z/v0Y1kR7uA6/K7/Gww/3SjXWzgi+OsjeavWHdf0v+6fO5kYiMrJi1uiHJ4bsquz
Ix36/FuT7KvAgJtfOKrQJtynJnhgovTtWi1PdeYqdVAF3k4vCEUqyYRaFGbMI7gW
vB6pNytiuwE3pO2KEN1pDytEZeoKjGQj2f/TXt3ehHsxwX6tUqVHF0YQNdg1u4go
hq23IJC0IXhQAO2ZLXiss4r5G0/RslfVfd1J7Fbvr5H2aMq+PP+X9zIuehINS40s
i6nAA1A8bIUSyunmqeZyKrTge2EvZW6TXYwzBd4TRRF2jq15OzpnQK3mgkqY5P+0
GTwum4RnWsbLmcHgw8pUdDvfDdEFw4aRcFXi13ADa8iLVsQ5Ybkdfp6I/o0GDQ6v
dTSEBEqfJ/joR+MMLayVvZRd8MF3ShSdHvQRWTiIj9Zzw/uxGUMVwL/c9YNfHLnG
SV/VMV3jvWd8DXFb+n0DADRERSRyqNvf+zGkyQUQbW/SwK6JToqr8YTK8qaUYGi8
6JFl7CYiu5ZhGfBDG1pbBPj0tePUHN1oJARnCANfWVWIvdH6qoK9UGhAbepIDipF
7L/2rA0scqcjIk5mben26bVEicUBMU/YuZL2LnOx5ZLj+/TfGaoAUFU2bbmptSpA
AhLjGvL71R1lBQ33IRivia0I8pXaAqPgusqBfuWDLmfoiNcR5fjgJ8y3yT3+tBhU
LbjtpsBizE6jQZU/LvHQ46Q9LiLRYZsEOju4zoWENRzVyaV5YxqyIUET0JyqwNMe
tzFJgOjz4k980ewERakMWSqDVFJofWmm37kMgO0uCw1IUgOKDTr1qQtHck4sgLhu
Om6zHJFY6e9ysS+rqBsr6uD2H1Q0U0et6bY8BmFuXi75Egtug4whfxnDxC2GBT2V
wuY82BXSbQZywo7TVPsy3fb5ZmaVgoMUMQvSaEOanJ8t8CTgI77tj1SSjO/VrL6f
K1EJOOg+DuKtw2LYLVj31TsYPCyHnTEHBhYz0YwucMG+8mrvuMM7slt6rrnT0+Xs
j9/LiMhCXU2xKgRI14Tfv5ZUuI47DczUI3fsgOCIStvJBiseG8ju2vwtTDMi7XVq
Tn2E6HnRCbgwO2PFRFGvGz9BGLUN+cEaM3cmZUlIZjr9TGvJ+m8XJqMlvvRJfhPg
hZROr0bhdnwYxbNOrDcCmCxK6hPNWAWAbNGT+xNNrtbJTWaYNyy1g7FHQLnVHSgU
7GBrP4aJTC5okgHzZEM3fW3hcYdAQCRhL1h/8FeNH+Db1C2lxpDFf9FAhAHqqdR4
0VLRsWNtmHN8tOOl4q/ttC/C6jsFuBe5LlWF1fNKPRQhqcEzzLJiJXI9ryLkqq5k
trJdgLuh/sy6RVBsWqILFYfI9hRqLbyTbe9b/wVUihK0vD5lyZ1LxQyPs783/EZN
hiplfFdq+jXmiv2CHLaHi6OeTWCc2HdzgVh88S2NrUa4IxjPEQetMnfrBxWh9vTB
sf0GamlZ/xqCJ5sAZc20i6g2JTSM7s/YX5uLY/yztt4DwM7aYeY4aUXUGUz9Up/4
lXkB4pyL7M2v1IEHExst5Vn1hlh6921Mv52Seyao3yQLcWxIVh+dJPdIchGXjvuO
l9CFpctvA3XPhyElCSCTFBt5P+mpYj4AK4eaO3bfiYa6+tFUHFcFWvaAUNK5Pn3Y
qmvesnXZcdfqjPZtVsNpAOSVecfT0qCeo7rMa89JMNs6HGYEtQSV675qwmlggCxl
ccPayrvGrDko65SdLDztSXOAWF6PAoyT5MOH9utzBuOc3q0KcV3J8p6GiU2AC4st
noH9McFSiQtiSeuukzfGHugQvBHftPVvEkQT3K6Qq9zmdo1qKV+QcealnWVTzZRV
vGnJOsu/5chgKervXv2CixN+xMc3JCCIk3dxEIXMILAZ3EtTWJpqgq25KPieBqYp
/rO3zICkOGN6xkHXrghQ8z8OsREvscHLMV8zV9Ga68Bq1dk1WFCHWvKOBwEclogK
JhAlxk1QJ3co7fg0HZsU9N3101vqdnjAhogLE3GF8dKTKa1xUTlmSmH7Z3m/Q9M8
K8Y9IqErsJHT8CbMBbabUZ9HxAgCCgsjS7OGndCdeqSLLPfZZu76L+AraEFraAff
m+s62HwPiaRk5y6HSBQ5BxPXDlo8ZdF2JMJe2nGUtWCMQ68koPd/OFiqbCn3Yj5I
hCCbGKLqCR+hSbioUHlpxsKpAyJZcKNMxJR+uoSHJzQavDMXW3Yyp8p9f4G6mxs4
DXyXICfObu2Eb7b6RoL9AI7K3IXY6KeDNR0c3MJCtQYT+mLs9sbYHRVJWz2MIjbg
M9AEb5bGBm0QZCON00Dbcwf3/OH39nIJ8UT6stt5l9KCozv/PSfpkd4mTmNxig2H
pr0nvo5TX2KOB0v89bQb969PAwQx+CE+st4IdEztvOhIYtO+SOYfNQc/txi+Pdra
2yOmuse1PkXeKC5etyFv7phKdnjlGzgdRG4/th2v6d5N+qVIOcYDGepBn7uAPbYo
WgBJB8ZXugUA+WmKXKvW5Sj25HBKbeVOIFuKQt8+ybBDgou2VSDflxOzOQPJSsrZ
kaUJmLWUoqJN0iEjVOPO16ZrOqw1QX4Md9GkNEBI4hWblNNpaiNFafEjxjUL7nYu
w2qn+qffhXT/1gxZmahfXmKuzW0LnEN6N5KXm9Djc73J29HowDDQU/YpbcXLopqJ
0LXOEEqR0vEjuCYwgCKvX7tzRIothbygI/u6TRmyjE9E1Ag8eVdSEHLCnb2prVtO
b+5eg60w6T01Ahk9oLn97YhQPHvExfVnayimM8j9x4vSyVauWjafVjy9t7Zryms1
zdun5yqeuanQslj/vdV82InSPvCSY8m0Y4FGY68glMvBPKqQlCbBWd/y1XBks+N3
LMg0VWijKsfeaxLMTg760OGIEH2Cx+XOLvOHHcl6WY+F2V0ynWX8N7qp4GkymZZa
1GIk+pyPrKTwFVVitk9c2+KL9mnAMlC97TlI5kvUhMmyfLz68OMasKjTbFtHEM1A
RFnl4U6EozzraGAJ8XBjBnr0dRvwdKcKPz8YNIl+B9hSpg9fPRpB0cn5EU9rTnsO
sIXkfA3CbdL79ePN6bjg/SXb8VcmLTpghX7OgWDkhb8jutm4v7apMwTk5nFa82bv
LQdUyyZUfMlmK13eXgugxyUmyhU9dUGrPidQwAjzm0zZxZxqC2EIpDfLdvb0z5eV
gBVL+fPnB9lkRRnLQHRtNDPcIhhRBYmPLXDMlMkxFy/5XtvFyNJr8VDWqt+tmYBX
JIJmCHz0UTzavGpjqDNohBNJtbknPcr40wE4c4c9nTB7D2APXAJ5s/LnJXbDuvB3
3JY1sLK0vMSbPkjd+x+YWHRMnAPHBnteyafbZUjkdQAUNNP4ZjiNa2scwhAwKKvd
jecH7PerRwtUovDiGQ7/IiTZZQpcENzy7FHjSQEHp5kJ88XTygSoCO+JnAWec5Ih
R1wG3iPZB3iX9E4UvdCJ0pwBMxVW/sj/ovuCnZyfFaQJVVDz1pP32bDOFzDBk+z3
z4A5LozogiAUVy+fXjfTYHCSWXV7yw+MwJRYgzC2EAJXGYTJnQgq0QO96u/QOlbi
0MDS473oR6I+cIHT6CZKaN5tjsZnLtyFPV8hJj77nUKrqa0kFwHjm+07kVKIFs9g
n1IvrPK0MW0TMRzFw+bTp2bBaKis/J3NQbZ3KdKKBDSvOsuDYeVwJAWQLZVzgq55
mmHxV8tov72P7fOR9Q65yk/1KsgPLddQ1BDexj5Q8MrAYC/7FPK1Mt8R6Hsk7Ckv
/ruK4rJJUii6tmElI4238FEIm/Kc3MRao3gLU/nbFloPjwWjeMH4tDbrf37bp+qw
nSA/3cQ1ctUeMuhEPAZDyb62pkhuJucl5dSJtyYi8wBiPwt9p2muzldEvzNqssbe
t4YaTTSjodhgfxM00y1StSBAm0FDmhvl3BnPXNSxAAzLu5OZHosT5mC5/8rKJaCJ
b6tW0BHxIkgGSO+v/DlB9J2l+0bqX41aBmLPaqPyRv5yhVh/XI8uj/gnjmGeM+1h
CWpYDqsCWZgmMUXPDcz92qEUav5jC17LNnOthV5j0vbe09s96Y7Wb+z/wPGLHWmt
3R+UudbaoIAyY9PKJ4Toy9dQdIlKaZ14OS3dUfe0TmtUDzi/cCMT1N+/HQYcEcdj
uGXc+U/wIT5mGTeuoU/AR6YD7i+NEszn97MXl6es1EuDUojsfjIeTdzRnfLUrEVT
WnBeA6DvUtB+GTFbDdtfFbtLfQTns+a3Sjmuf696DnUlAZYGyY0JhgKJ1qtrgL6e
LLYazZYrLT1R0uHXDd9P2A3wUYkAuCFym2Csi/KOezCxr8LzvLatGOo3JU3DsEO+
2KYn14fhXZYWPiGoCe8/lzlbTidPROQ5RAg5urPFM5xjzsnDPL1GSk7iU14oEyDq
RnVPYc2KYZ+8wrntI/qZxKphkZVHHBTVVIsWP3yB+/Usom6ZNTEuEn/qyFyhqnVE
g+5BGHuxFR0JAbaE8Zi38zgeJiDLBc3LbmtQ/EjpD0fKY3rWc+HSD4vdbCTv+jY5
tyaPeuspYH4WB/pv7BCVXbMBu5c5xFO0Lb0aGSgIqvhxZOv2Wjd4iaJ8Xd3oslFn
iNdf6uBzNmkzn0Z/LvNl6krSMNMM43CuZOOF5OFaJEothsLIM4c/Cm0qYB0Ep7dx
tSKMOtriWY5ac2PLCNT+dDLFlsJS0ndCN8WgWna1kPCP2FIBnPL7XYMi4QiQ6QlG
ssQ/RJT6qIH84fh0HRCMIFdny1RR4xYXbrewaZad5byNuxKxseCrD7k9ovqiTQQt
12y3Jabtx62783K2lwCeZZduMDNUG48iS9qU9Y1z0Rw8MczUaWQdXjXR19adnBMu
ECo0271k5HjHwZtx4VQWK0VVfs5kGcT+DKfxCsLBgXgE0JSAkXqkYJECgBMzaSOI
u4obxG4rjPhIYDhsvvZgqZyFMf+XjpNH5TQ1sJubkjOf+btl2NVqtGyt0OTxt/lo
ioGlXVWQ4bN/H/wQab4mQBRlpxl958dlW6OeJ/lAxhTIBKtsChlsxxmRty0MKZqj
mGcyEwy2nVQh5dR4tZcV7d9OAyQZ+UCCcKyQX14Iwl1fIahuXM1ivcOXWJZGK41X
uhoRE3X+YATq8NUQocrEOPd1laxa3xKhW9NYPJ/DXh+7XsucCDfrX/0vvGdxNqdp
n8moh4jei1Wuv4PYEt8nZIRBtT7ZvEn4FVSEPQEPbCK2WLgC5QW9cZdD6ssfNZhQ
oXfB4ic08qYR06OZ4pKXFVCUVNZSWf5u18X4Atm8/cnRA3XwfPSgbV4WNcSPh4Xv
+6NElBe1KGsLEkg3hTzqULcs4wjRI+TJ3NEbCI/KKvI6lXyVHwAhGxL+tDj9VSb7
fu/8Pi1FAUjvgykKRKCjmpPVIhktZEPnlcS2IjvSrzowauwGBdQnDOQFpVeYx/cw
sTepsnj+pP6nkXBqNx1MEkUlX7xfdWGyyR+8aL/x6yaWo4h9d/oLf4JshInEflj+
bvg9cmtFWcrfgbAzDBFpM/JXkiCGhtjYe6UsLj7htf3cAZ48GNZXPcgL1f+8v4qM
QzvBUvZWY8JFEHP84HSrhoFZzGL1dkTDkuHCL8iEJuWpjF1d4eLNa9eLIwgUmkUI
O9HMkG/NVvRM+SHRqcAu1FckUncrd4KTZCNGU81GJUaT5HvUBiNq9KqEEIZgVw0/
olHLc/iM+cRTB10yCKRalCQSAkUMvO+Y1rrNi5Ynlijj05WJqC4zw7vK+TnUygNC
mk8/inznSsSIYGS0jmtdq54Dm5jf2X8F6+NiGHzdKWwKq83ejDbux6lcXtxTWtfz
zRSytWmPPtBHUHpXgq34+BegIatSHXOZWp4q2o+w+YsIo1yljjtswel2XHF1BTdt
3vPmBXVySaIzIufd7bbDTxxcqhMD+Mplegbn6FyrUJ1wP0r0zgDM2R2ci/iWBrXF
ftd9sFf9fGrEWp7jknAX0nKBhNHJFWhGyueTCpOtrbBByZe3cFg1CGRffWvFS8rC
Ik+UkCi3DtLZk0U3Cufgi+BGER1oCeF2K6B8Xsn6CxmN5VQD0ldgRGfdNj1ACQp/
Lw+w/5qrLwkd2AdKd37SIzNp411I1N3Bw209iiem6tzF4MuabJYbjXpEKIn3TzRI
ed/df0fgu7IyRZGSpXPcQCVNcBpCBZhVY9VY3tBaTIDXWEgyD1cgJld3oinsqfZ3
2DifGRrzdcq2Ohhha3e4UlRme3VT9322YQUU0IaKHxLtUYt7/GGKuQ8WRoFwF/GZ
7VQkOVbQrrKqMlyS2kVrvTTVk/L8BBH5fPwnSRpBY8BID0DoEFUmdAA1nyaElzMb
H3FgHn8CqYG6X/LZ/5puKbPlLBQH5iPhDuEzi59xjSHr8Y8UFa6cOkyavsW18zNl
RroDJlcySh+2ztZIjYZYWMWRODOc6KW1J4QczgGiEkvBf/RkagJ208do9JXtki8M
kZLybKwDMJ/f8CA9lfE5vcEo/DZtpfKNTbmcBi0uottJf5uvQ6E/bd7mdVnxXADw
QpWqF4dTwcNeuSf48JRwF5RcSMMeElqPsm6iSc3B4L5jxF6j8DO2vOwsjdD9hkvr
yMtUiQjyzaM8MyFluQtt1UN366pSHVpDhlY5E2/DhZauKjXKdSxTX4kfISL5JobG
DaY14pvfX3pkHa5nKgbeOudAsKJbRO9HpgeXCIvieP7X/sBm2cS3ZiBnmZq4Qksq
lOT7A9zwgfGVQ3gaRpIlwYfTlww4jGi8qWvGniFlJqo34Ol5rxVPHTY5G4SNRdgl
gYTrnzOLZldx3Y1hxbfHIa1XMa1l5FASxmyDQgOrt7T5VTfBOvYNS5BgZIXxn5ZX
YH9DfYvXi/in3HRfqd3m9ZfwsBmah51RMMrjVvBAmC4JoBmXhW9xELJU0I5v3zP5
V6HEkLcyb53jNdXooPPTATF4xUQjc215P+YUwLBtgGGzKzUbv4mXwy46xzydSxWP
3XeU9fg4vytXZlZQrPwLrHw49pgf/mZFtsAUndvjujIKH6Y/khraIKnPNMG7uRVf
/YRztnvmk11IO5gQ3Iwx5Jl+TPLidGzPLJq4gKs0ykJi+2YB2RW9P5W6aMohB0tm
7KiQgPbPjYOgOf2KONvlBhq/tVlyT0uHJYRw7lCq7WdWPV6JrOrQVUuOz2puRB1Z
fw2VZAJF+mpAkJWOg3G5C9OBJG5DJ8acofxLV5rcsFRHfGmb7r1GF5BvIl21LjrP
RKDXbm3tiXYR6EGlOp+DDGIwqPN2RcdDft0tuhvR/G2GHiKtFMjkV3F5qhyrWYlq
eJ6wjI4fvEKN9fsXKwE3ooJmDPbc3ddiS3UnQmAagQw7vMO5+pEnfs2rO3kDNpLF
T77a7rz27WReuDTJ4usTsYaZ8ivAbfqJ1QQv1ws0iOyXRUY1sitF0bo2v+xPyWcT
jJZKYWUZzObhg46/LNnv1zGnSISOB2b4XmxzNka2wDIBAKm7fW7Axmlw6J5s/QlL
lZPM2Jj+JjeKR54Wa/uZg298YJEYwvSJmfJA17QYzDz3ifBeCjpyl0qBTbCda/c+
1fxTg85xfwx0dQHO0hVNG61zTU59gHEQKrOPXIZHdiD5dTusNMTsFWpLyxSDP709
s9qELP5ZP5+PVL1NyYDv6U1a6vdO4zu7luxlQPexasNlXhPolImA1NJ76r4tYvNL
CqCUVsO1UeJncZXwbz6Ns+kzLSZf3ij+CfLzTd8/nWDHGPP+Cg3mW1LSvjLHYelb
hj6Jx93paDq/7K6ePDnBe9mBOoK9WT+ksK6SJeEg1D8vQzFedCpKBRDZ9898bw5v
lH1ZGXRvK8v7/HPNIlI088AYnl0q1o+s3lL3cG8o9oE5PTtUm+/gHaPJa2rsCJB0
Mg48Unz4GFhr6JyULMW3lIppNGJj4Aa7ft7APZFWMwIHA58fLkLEgiOyABd1JZWy
HfrwPzcnhXm64PHLkTQ1cMB875WYkn7PUdgg387Zxiul9O8VvUJsOhXvrDZaHOm1
bcJEcu8rAkboCl2YszIKBtXN2vuAfPNcDVAMAT+oxeyyykkKKEXnyNp3eJVzQNwW
tOIOHnLIWRL40oqzFL4CSsvkZgX3gMI6jWAWlj2QAzM0dv5dKic8OVDO4pQP+F9Q
865INOtvxEJCQyzAO9bWnmnFdePTFqN2S8fHK7R0nPn+xK9Z7eHYQDKt9+EJPFr6
3I2M7wwUL4wSaSTKKGMsqhGldDu3Fj2FePDbZpkEJjx8Q0nkOvCvPv5L3ZsjGV4T
Obi8r72eaCh+jrIFj9R3yp6i2QaiIdPzr14BywZmcY4VwomWqfuepZu69ba9Ph0G
8mebbXk+ASYmQ4Pb7bh4AO5msC5Ws0XaRQeg3oaCGvdb5TI/bYarZO1fVLZNqhqb
yLH8+wKAU817ieBbJdbpXZLg9zAKBxoZYLhrMzwASIsP9CtFTL358Dnyss0MIs9k
c1GMfGKHU6xkL2+0iX1mKOQvWDfFM1ELw5+Q8I9TuJDYKIdu1TvWlAR6J1ZVq0Pn
gnipWx9nnO5sG25mIxtyud2J1LY+Eiq1ljBMIw8eNsORwhdaA5q8eLtrjsYxhpt9
r1vA/PGodmAbxXXG0raE7Y1suqUiXyXIKv0oGqWUvStQhAu0Tg39y10jp0ge8eWo
vmLwdcsumksNH074fnQqLMilrsuo5eTobCa3Kj6TItaT2kiU38rfmZCeClu0gIsA
QL26FRgx3Ag1kdlvlGu04M1aBgJ6XqkFeOL26cbzRW/KongDqwIoXaTUTgurY3QE
KEiJQSdFjweg5r6FWdq770HdG8uHVf9smGlrlMeV7DXqJLHK30SgPvSKz95C3oIf
YOBBcDTUANb3B7L+bEPab+YDRohOj8jIZfajmkF1+vyLeGNJQ+LlEbOGdL2NuWFM
SrejhETSqH29ZbkLVqfjsJueSVwzv9Qgpq0pCD8ArBQfEO2MpYLdyCgO4ZL4kP2p
IURqZnqOjqBsTTFPbLc6l0n31VA8wzLOFKL+I8nS2HvAyfsQIKDteSravAc9y4Wy
C4ZmXC6tLjWH3r3+R+8xBzjiIWBhWivL4tiuk1Dq5aK1g+uPc/+askxWxGiOu2OX
C2EMMsCJSsF1jKCoLFMPhlXeihdNxEfcgJDkeKooexjJb1vDtjRLkBbGRdUESjvP
ZZHt7QRMLGZR6e+nHim2d1edArOMI/k1wo53jiTkXGIYhwIrfDZrlGHEyEhE7Enw
2cNTOnahupmtPXsolCJ82qI3icpoq1uzWBDSAtqSMZmxRse4BFYSINHsMcIp0cFy
3crxKZpEJ0IUMNPyadsxpdbqkS9O/irPyvP4aTravsJEVu4N/4Fy1cYgIHSBvKNt
/+TW+8YhldVutRxDMc6SSg2nkx0vQZlo0C2WRWNtCF1J8DERBxUudyvmgpU0m2JP
JA2G/o/azoMJJD4sI2UXuzMa5Rqy8BdiDIOQ83nXkHV+xnyWJS0TNkNnkhnOUM68
R4wiy2qs5NyMJ+iLQZgbw5XZuRGnhMW/TsLYRvgdOWqop9WJ3cpcvQj7KCFO+viK
0PCxALlMF53pn2j+r5BuA6kmpkc3877EyxvnfR4cHfJ4OWruyPWJlBsISsTtcG/u
jFkorORJPEqgQ1N4Q91YqAwfzQQTzq7hC7kr7beh1RVrjCl/Y3kLhQMGsYNy+aC/
02YAtpaMitiNVMblYxDulDi6nS8pXuC1WKhqvXd1+7qW0LoKAjH6hywXs+AINC50
pCxrvd3elTj1m/S5HLTohEb+s3hKt1dXB/WuOPNGdr75hPqcwEnH5J8jqE0uKwEM
q1kqKa4KspEqJ15MGl5rtvGalWLmWVI09HF224vsXNKCF1bIBS2eEDS/Mpd+Fa+k
duIARwOsi5h/vRZYGqrxYdwcKgHeZeGswTzf6shq1GmwaXI6rbQJr7JELgiYdLwT
kmVYAo+eEw5nfTjApTTvePIUWAtTgiJ56BhBmR0K1Kx9IPishSVOTTj0NCfUiKpN
cZxgSIpHa4AleiwNBTSSIyHbswgeFuMwSmKBNOGbcxZSGntMPoACYyqA7egPFAwT
ns1KyfsOcB2ZYjTdTLL4M/AVsQdrvBIaEy/Qlxauxr1nXCOfu8Cu5r0EXAriaAQB
k+HymrB/TeQGGt0tmQMcmd98IqSjVrLFt2vqMk1E8mLGy0masx7JEZmGfmypNtqq
UP905M0gmJ1LKye5C1RcDJcIIFU9Ap6HVEkOxHmUCXvFNwIIwXMboWK7t2i3/rkL
/R80I44EHvjVvzZv004FDWJHlyoLfP+x+IlTP0gYF790hvTUcUVos0S/WiF3W8Jq
SDwAvXh441Cbzq0PLS5F8FUmNn3Mw/yMi/rlMX3H4djwXY8ZOC36wrJSxx8wSJ/r
/qORCk9/mQjmjH1JipVCKuOdMEPckuQ5jaiSqnKb42P5CaA4XIb58mtCOEEIi0/t
lK8tt23J1tflR/NVxKaMVsTLXgvVeqjoiCPWwjT69CKfq3hhiK6mEh1k8Z/xrOT+
CzQ1NerAvL9fw18N3b0FMiFApYFVqem3iFbKg9+i2RVcDW3JkMiMuMVrRp7MGEJL
/r6I4ywP4TQn02hQkFi03TEv78mTP38GoJAtky27QjNtqu+uIcmfhEWFCH+a8LSK
B097z+gsJpSCs/PYMMykFp2sSJ/1kpjRvU8pimSawYFACmmrdl92/L+kN/fra3tZ
dB4lepf7OsU6gPHglcv0hoZgoykVjV+fkYfFYbTP8Bfoycc6Xgs5xOg4XsjLHvsc
7Lp+pfaRP1ztjEvamuG4M1izcUyO/AZiQe759hAGF8PP41h4Fs1aVqsMcfzyU/Wu
oI1nJLkDpc83Fy/9u9hRypizuSxPIEwW5yMQFBbQHDePpMOp1XoxirRzmbSA4l4D
Ic+YGTQ4LBPLKOlQR0f4Yu1XOm7vsyC04hTRu4pibNCa6I70D7WImjvE8xAGQeLs
t5a5OqYytqccrKlIzO/IrEfiSJiYibsJDOFfSGtA9Hq+rMCF2pMIsu2uSiEHXq0S
WBFi3XvE8EvguNWekcD6WinWgDsVIvA45OQe36HriJl/T2LSGftefTovRef1+DhH
L6DYRX9ALCsEhDvKKgIDcp1ibvffKZdBVFfmrSlwhnbItN2VG31ZkTie/7sov2Dr
34MlfhDDTdUXQep6un+8syibzxKugu/n1VKD3giKSAI4o5SvF5GECzqQZasKVkOj
41ws3sAl4EnjteY1jaPf0QZm9MPJ6uIJxQRnyhoOAom7hDg7lYsATGQKFUw81+Mm
yX+IYvhhQdxjG4QZiT6L4MeXdgEoLd63NibHn0+n2p6B6VOhj+CZ4Zy23qO7LvUI
zQsiSpdrKtzsGgzYT/1NzdSjIU/33LAIVNfEw0+rwmVOj7ppvVsmYxPb1RUfmIGQ
0wFa/7FFKxWX+Qp6vzhjlOtURQNoUMXhaLT31lVJBnjKZ/kZIRMnN8ZAhx0uWde0
04Mf8Lj2DEzl1MGKtqDe44Kc955vWKGU3pq3jp8tj7qOaQqr/4PO9V/KAOd0J1OD
iOfk5Lf2XKQ8+Vc518AT0CgTblZ0ApF+4Tmir3C3VpJiEKdlkeFRD5q3Tpa75sea
ukUAdjGPSuzx7B9YpnNpER7nZTvGXaDZUJfK88jR7e8f+lS0LL/V+ZxDMt/QyQva
Z9/d/MuECIlK7G1bq4v1oDUZiRJ4IRX2yhU/l96QVdoxl9FKmyO9JaOTQzp4dWK2
q3yfjPI1TQ5aOxvinOS/1hnrpfqoa3//WN89UvHr6hD7CHHfpQ92hG0pVJDyRe7I
x9PPZa06eoYpHPjYRXWlscV4lxpIQBn0OuPL58O+Td5KFbVbNdOns7MN2vAPAVjL
9x2vjN4fAJvI/78llSR/i141l3kkVfzDBPjwrHS+IjlFkM5+DSQxs8a/BLjsg57q
fPczIzonFaQ8uuwnAQv+NMj6TMagBOfUfr2Lw3SgNFQanlswPLT9wzC3ssJemPWA
1luK5xyNsvo1vWQVpTDV3JSUzr0PttnUlAUGVLC1/q2NUSb+WZiGRKXktnTijBR+
QMLjDVWTrZGewsQiuJ+ZOrs8If++cVEybDjIOxhCa0pExuZpIKzUzv8XB+9ftqMZ
anvEzVdVIdhaJhmb4lNf9BnyR/JY6E2UCSwHRAJkc77Pq2ZSwsIZPxUT7yH7vyRP
6FZ6dT31P0ir3yItDeRpT9gP1m02ikcFYWGRRa2ZEV7k5ZYK79xIDz+I3uhC/wYF
nCrm4fwFJyUxSLx06QFh2pxPgimhGj0MT/i+jkNeLcJxvniGjBUKLgaoCWxwVTBp
mKFN3JUPHV1K3oUyWvlEp1GpfjyAkzD8T4OsF8htrLQQ9QlmOEeFGhC6z9HIennC
qhwlc4Em737hu63qsPd9Yfz+IQZwb9trZSEdkvJW+u84CKSv5Sx0Y9pskfmBQlI2
SEhg03T4HQ2pKRXkGLYZpiIFndBIJjy82nwXuT/WKwPcNeVYjCYrYdZ++CSEpmH2
3EFYwXMeniiJ/nw8Tjg3B6NWs+rBpBaremC5H/z3b6r4oxGvsN/Oh9plTMfbxoHq
/RRzdeBj4hyyJM6MsIFDqQ1qvEj6ImtIb/yN9qXmMOStJ1zEZnUul+HHh4S6oK/P
X6wp744fufZJxs1LzoE2JvQRXa7pI/vce760PYcxZfyHOctUBcLAvhbWY5iL+PBq
FYvq3MRKQLOANSoZN/csU30wNPLnxhXbSEaa4gAqPZtDOg2OfsoJWis4eDDdTVER
QzYpyr+ymW4HYHW0ZXUIQChqY4cMq7zYvTEiklKjfRkwTM0Ao7F1RrqkypSiLmgj
qgdMOv55Hs6Dce++LIntB11Vg2WlGCjCgHk1O0uIGJ4fgT73fMt+dKpB8cL35ZTL
h3r2oBzSuUzEGeIroCWqZKV9kQq27uM9ZztVZbQkK2+s6Z7ovqODGOVPNn9hFMe0
eW6TK1jMQbIX1Y6LEIEO6cBtVl+lyThQKKtVCudLpuiBuVjoGO6tIShe/ncgMLZw
2Kwzd0YnJOZU/p77Qo7f2mMz/ExEaky8svDJDw6UA8e+9QJxQUF0pmAs5zdeoK5S
c4r1eDKUDZnJBT2mgbEpRggct0X3QPqMUlxMvrPZLzw5AIkFhzFvt7FDFaghBqV8
/cdpiOaq8w/YytuquRImky2wpxG5HYi/evFA/JP5MH4D1inKPY+UirQXUgSkAXiI
N0phIwAQJOdo/BOUPAuvUkAlZdQaUjmHC/eRlXpia/aUp9fBiArCYE+OdPmaYqUE
I4/D/IvP9lBpwXC2Ns6KIFzQu3cKLSzqIThGcGJjFAkQnPdOPJzd0qeg5J7jq81c
1ZLpTVOzPpuYVphx0HcHHqNIKEYAxtAsAmCIfwyCeQiH8ZyS+v72eWNDZUaSxFAs
AErn2N3LXrFZBJWLC1++YSWjIuK3Gt74H4btuUcxT7Dit8n0H3jWS7+pVuiEq9bM
PFv6Bv6RLvmava+WADOrqEv6RCwkn4iRhcLyzfIFodzTr5SkRH/evYmzuKYc5O53
C9ulGbEeNeHhjJ3JkcGuHHs5nwONCHtDvN0y0iOvB3uXwJ52xtX3fpl+L/iPlQSo
QMYKf+f37AZH/oD8kBWAYB/4JVhKzqZPBgx3EuUiP20dSqpTDsJd04YTR8ZW9q3N
RRmBUmV2LPHdjTuaK7HfswdKGZ1fSzreJmAnOtHApm/amdkDQ/vJ2gl3r1JGHlVM
bTaXSfNKey+U7g5ZMMo0gwsRDIrgGHiR8lXAVMwzkOOp79+rwlYVuuptvtErnrab
+Otx9MMtFNRpo5Rm8lFP0ZrrOVWtdp+z7qVARN3vqmXmb2Er0O3cA6WZtnzmazs+
kGFmFUTGnOlh4piXKuAbsESxBhO/LH/ZsnNp5pI8GQ11sxMisYpje7x2xtrHAI5B
Wy+zOQV2rRAAVF0O+kqtl0GYBoh64fskE5VQBlWMZVJRH545edRnp92a1MtL85p2
w+LZTIwc1oPFOVUQrLU3p59lUIYE+PlgYV0ldWjLgtbj1xu+uO5Nx/22bB92j0mc
quWrrpLhpCnBcc9CcxkKPJGImVGNxZV5f4+d6MQQWJQMNPhEoaxSNO4OHzzLh/la
f0rdKC8VRtQKd8T6cF9LQElHNTY6a6bRIGAyE59PC8CACjXkAI+Twuqp+ho2zVQN
EIQorYgCixDTMyVenVMr3lIbddeZMAO0fNvn/uMVWqhjU0LAeVRriifrgK0HFEyZ
1LSwau3qlMJxYgFCsB+1HR7G1YsaIjcd6/bdf/TSPGrsYi0y3rY6RRSd24/R9y+u
QHa4Eh89w5SKrSqdK8RV5XhOI94359MEIg9gf1iEXDU12v2YnFRr5FaA1LtT+ZQI
sCZ52ZC2QcrUvhqTA8XpRDa2voSH8qt34eU/tZLOgfg6MOq/OXsaubhn9de74dVo
wiemiegNvJ8F1ulBhJi71N16w2PUU+4HoFRWC1J8TNIOUXBhzUVDPKLE2teT169A
V3xH6ewe6Olk6T0XTDX1jGG4mPA3Nx5LkkM4YsUSxBbUNjERnOBkm0zNRWi77Tdt
xos0Ye6zdcdpHGJxCJ0FPnZMBMoHAYpsDCN5Q8cG1pSCX3RaxkNSlS4T8EAl2SgR
+yZAqEXZqMr9Ztxs178XbztfORgV0SA3GpIhSFA3kc/RAJEaeJ4Vi/7Ly96Kl25/
JnQVvKIV1ZnIQQgz+ArAW6gUTQjteHedCIonDyEqXPDDuiwxAo8pcxaeH9L8vGHe
9ozBn1TRDCCSFXKJ+loG6fp/2DoQM3O0KJEQ2uDcUUeciWzBM4F0WQYJ63KQ3VWZ
o8UM+USmOluXzp0PMQJ92RV3KSN9eYHzCX/JoC9sdMqLGTgBRbK+7tIaS+YTxLzp
nSa52lhzG228npGBW3rgcHaZzSOUq5XUMeR91QFeg6aaokVBhSCfWfLVB0EyUOzK
18ZA8nmVtuv6Cy5XYCRGT7P8enRqvRsZm5Ee5fpsOIsZoRnwvvkK60lb/KD504GM
Lrkg/q2wghksZt9R8hc14Su9OIJsJizjjeGL5Ae6rWkBSYztiD1m9hDOW4TkMUHy
5Sl8gvyDlwPs+4JupG15SWNsvlUWO+5biAOEq2zHlkCIsYkLkwIyqp2AXk9f+IUE
zZvw0rVAXDtCHj0SKueka+3IQGxynlayxvPiq+vjo+JcVLoXV/wqCmg60LY5tjSm
bN+kGHd9K/inSpsk4jyG3ytS9qPDxn0FBKY0cdJmSm80jXMCW3RhvlwxRBzOox0v
UWNo6k6dOtSD/sjlMlTS1UacM7FRQqgLQIPTkzlRMcqkCNePja4sNkD6LUjapuSA
CDEE/BjIT9cHgznMsNf/B/Lo5eb3rW6sGaFuDuwkOdomzHFqnMho9XScRmdMSuEf
DkqZJJU5rUVUAg3I7bD/HEgiQEzXDsK2Xy4t9qHExNjJlMpqZN3eraFHwy0cE79l
PWf5oxUkhW2IZxKunYNwPAYvLV9xLEDUTlUFKVs7SBWLomtHdu7MIgNJbOcJfOZN
faf+QD7EzK+eXEG9nOSpXdXCITi2u/xOzwInP3KKiefrdXQB3cksEbK6RC1jJzJx
IWuenJiuGgy1Fn7I+L7R3nGXH9Njka/m5AuT+Rf30iAqLtOR45daMmY7h/UmXR9X
lKaWVrPyBT9o1HdQHvNqaS5BySgB8SUC9drkvfhX34Es+wC5M2tpGL6qtCsi736F
rhrgyztrJrV1agr+KRSI6h8OES7KWTTs4mxtibdwHQF/M0k5a3TzxofYznPvOUId
eajSicHk5ajdkr18HuBXf/6SLOhwjD/TC0GFCIWGAp0yAf6iIEyJugJk0CFKwyI9
IeR2gYT0sg3n1SJlkQP6cmnqUnuaC/kGgsFvN3B3o9woq9U598ch5BZVhOaW9yZp
Guq6tjabK962j1NsJymGM0xXyrO+Ey1Gz1jIbQtQ9fkqKnRIyNvuUDZ1PtkXN8zQ
gvytW3DtAAeffptmLM+U6mMU4iWo1l0e3RTliN1WeFn6eIav807S2yg6H5cyarBt
fLuOQ3aM8eDuxdaC2cVtjp8Lk9+zn3/tumYQXPBaQv64eRBXcLRMOlc2maKBX+lU
+kHGju/0VS3jDd+aV231zwtskdNvnCm9MhcrIbXHNr/C5nAZayRAKqn2hEu6eQi1
P/BiGh30GYWMIXaBP+6xods0wR/uaSGCnMpryYYVCF7ZaT5zN+SG6PUS2OGpx/JH
6K7iHnucxxXRF1/3MsHpz39clqarVStaqiVL+GHCLACsMNZ8Fe235vo71zLvddqi
IGnZwAdmMGbxaEc+rTGbNH0vyA6xGkD00O/aFVwoTwtagf2UzE7KoJCRpgXWanbi
4mZJ3ObcsBxPWBodogxR8GFtqDE5lGZ/j2i9fY99P5YmvlpD9lQG2db1/B7jJGrX
r80kT4mFPRt85Ky1hRN8U17soVdp/bBBv0gKeXoYy6JKmVlwu9JKm4jwJ0p02qae
d0VnUSBQfccY/76Sk97NijZ74brWjY7I5j82Jeo7AkZ2Dr0rckoS7/mAauvOyQYc
PtOCblrHqpFip1GF1vJB+aWmbbssKD52SqXvsvXTgkFc7QJbtfQvlUXAyME8XN34
rl7hA6iLvnDUPyeeAB4vOKc1+9R4sQe+mrG/hlPPX9qowBnJODLRNj0Cm3WhNE3e
JLa7SblUYL1srD5uxqmTRR5E07iPSM/dhQ/3IUPUjZVfQ1ivBIlluld9P5BJihQb
b3URJmqWlspwVdbMzVUUYBgq1cJOOR0Rfnt8UJws3PwQEFlh94+K1mKuuxdxQJgZ
utaWH7tSfBRl6bOl6JUNbT+mSs2CnSZwPMY/UBz6Njkm+dvEd62JpqeHT+zidi9F
me94Jbevp3WFVvRy9oXOPUDSRa5V2nBSbJcrKjd0IxrMjsbuJDS58DO3MlfNYtZK
haGcy6OKMfMiSYbbhVQKxBk11w6K/5nUqG9rxCbKFkbqt+UThaBulLKq6xSQ7rDE
Jo/OCymqMeL4QHlGCRQCDs13SAZP98N/h5ELRGVKIPfWaCDI8PRvYT7lwpdllWdM
3tRMLje6spnEmbFyADATkkpgv2ayjP7XKogDWM9ZYig//7+cytKorSDEsFZVFabn
kCb4MXYMnTwQyaNW4mVYOPM9NjEU7xKUb1rZ5XgaehoWIdaAPLHz6vvpRJOxgCSC
D6G8iU7AcHSgOwUNwjP6tIrVWHwnUtDN0HEm0iYXDJLcP/n6XIhZIZLpQakukpxZ
g0/zKZeab178lDrBIzKrI+3pEmeApYktErfIR7zX0BIiNQgMubNJ3gYPc92Zfm0Y
JznnVU0bwycy8/MZjh0pMZd08Qw0G72lJyUU1S0W6K9Kj3sFF088sOs45KjMxE+Y
1u35JJuNM09FOlNTY1apA8gtTN1WUZz3S9ABgkKJcx7SaY0DyWiFdlT2f3BMsPUh
JjyExynRFpOVWfadYFVuNZm6cioPdAqeP2RlucvMw1vit5wI0oDVLxnH5pdkN/9+
Bl0+7zEYBiS+mw5uEyJah2dSI2Ow4QTayEV5g1KZzoO4rcIDdiK/yPtveobNCdDg
h3LBIrE0sz0Y1kfluTXUwnYUpxw9DQ69U8csIAsu5kCbAuUORf7tOZlBzXcwxjke
zKrBPaEVFwrq7S1hcwqgredOBcMqClu5AoJK3UEBwlgkLTSOdS8mUXE3fzb5DN/W
DH3MJrVgoM8lsye8yCNA0AwsB1tJT5i/pJ/FNmc2yon/4IuU9Okw5ROpy194X345
K9PtGlVXNZ9x0utDqAhgfUZZ/fMfonOW1207CoJ4RM8uHD+pi2m4YniJ8NuZ3HME
xeSC4mtOd2dGlD0mTxlHbatY2PCaAolkg1UnQ+BzPM+pm+jniDvgWmI6ynan+IKn
P5pgmeI3CpiWgDVdPr9p0OVUg2nZ2Lmaep58KwjbzJMYOTf1oPm5P/NoFyddjB8L
3uLwOdqcBqnHH/QzkXAPnJRViHAhNgvhGAFkQWew+GErNgrBpUVSISHlubvBvinc
HVwivIveehN9hEYTBe7ZWlAhYQP4tslaNsLjg2d6HJ6vovqzOqDnzKw4Zm7+b8LX
9cgM+969NFKke0VTB5m0DaE7CpF4txRgvT3vUkwI9VS+uMYipvQpa3Nsj+PqHNZx
k1wEOC9HqB9KdFqPaOaKBNPZKwrpkfqUnItuSH3gnkBNwuWRcSafyiUEiRpxjBGm
Qo7oio5b0FdMAhvYrDEKE4p1IzGcdA/j3JJm6R+6VKVJE+lTa0RZnGlnzybTo19k
15l4BgHe0x7JaY8+RSz3sHOhMAy+yvH0OS2Y0sgTZQ1UriPsG3At6NIN3MWQ8UdF
SVT19PDyRz0rzneYG8sZeghZo8D1i/ku8Gu3FUjIv26jLJ6T1JDCay+NvWoSbHUZ
mJj+tpo5RqhND2IKvKVDZOQhSVGfQO8n3F+J8DwWH2C69214bM7SRn0Es1qGgGr3
n4AU3VgWyDEle29N34XTD/1W98O+jywy1DX5cApH5vjjTbbFP7nriGNmWOgwFQz/
utRk1HvWFErYXPm43zlbSfXqg7CGl9+Ks//ebQtIkYJxw2kXT/ol8XNzgBHAnqaK
ojymiipzx3DI+SnL/QvKc1ppRX/k6B71k+fOYwBfk39uNaGuoXRo+TYyT1PYsDcn
0mNrCKhhNTLhEPZGUk7CS6H/XC8AZqrmqe5EPeY2XMpaLMxBmEzovjm+GpeReyxs
dXC8V9p0DUqYC58D0Qc0FAyENsXj0znTgN9lQlp2YqK/IWUjQhQhRVr85qGqKVwV
IP5w72Lykelb7tRInkm76uj0ZH2nRb6iP1W3aoYpxhzGzQ/F70d42iCeb2KdYz02
AyRZ++OIoxVX6EN8FXsN0gJqxmTFf7uROQXR8MVIJerEkgmzS3QgqGr9D55l4jk+
Wzm7Dxyt/DPbQ7yZbN9ee0NNbkTEyXcOZIIF04UbqU96us1ZQdJMKVd9vZ5FcdMI
wb/7KbbwDNtw6VV7xkW+ttjOOsoNO+7INFQOvRn7aaST9HHJcNjkiUTqP4zdq/rA
8NFGPc03D7Iln/1WSIS9Ky+03wC5Ug5zm4AI/TwLJ7crCJdLEqu5IA7AX2k+sQh0
fKE2uK6a/KRMgMAjiG8uq2rk9Qm1XZh6GPRM9Fk+eYBo24sBPWXFXmAWoArgEUMX
SaXxz0teQ/mt8JYsL66hN/GO4C9pSKKvbkiL5Stwh1gBGH1yp61EGRvSM8r07qgZ
TKX//mZgA3a0xN7rAO325rDFASxQ17APYr3R3N1YAtLM+/oMmjzYxu4Nz1qb2USv
gmu61A1nTTaY3XLCB0ZqTTWaYBhKYfSK8h5QrTLCFyQ6hDRnqITQ1KKG72oepfz1
mbBjw2UW/U6Fx+tcF1+SjPegV7TR3NtSGc7YVwSfiGTDGsAwCM7JzhQ0Ycww+umM
k+7Fi5hcwhpmkBCFU2JtIPTFdCSxT8rXO1jGKzw73B9f3KKUCPEU6P2SmJ95815o
7v0XnK0mrDbtbAI0A6BpMq3yTe4gbuvqUUTUqmGSGVNPWYpe2DkkiTBNXH/8BcP9
79EuELjBrP6GppL2jEtL5H8wHvI9ua8W39ZCDfo5xAzQRbhvFo+N4CLiPxGOC3HU
dl0o3Fx/8/9ZdPXjrS3gwHcL6SHwTiG2LksGnrtRrRt/7X4U1pCm0wnc5DdHYNtR
KjKJ5yei4lqnuzbW18v3pyZaWac5sdJEEOZqmuABgP2hb3drzHzeqf2RpyOR8Lip
HOMlQvUjB4h5QIxw8yOwI3npXTNFMFHTxw0LbNlh+votZMjNVcfOpNT49O+WZFi+
vQSELeo76cKq/N5fYOnlTZXunJRWklXgp1Zd4EtwcuoM0Z8Eb9kWAae9i257PqK+
Qp/kxBn/vlLn/LO6aeHH+tGYOJVQ1JBWMKfkyMo0eShV+djyGeUW5ih4x7Jm8Jf4
uPfKUSrRvfYCj/FLvZ1haKrYogriAx9DPwtwG/AShhAShQSjaPWyNT6gRUaclHof
291V8vlLzfWFSNqsVWnaOSYM/9L1h3vePZSuDqDQHiXsE199rtCTQSdvCY59BmCi
pwu0/hrE/cu491+hONu0hV2GArSbXQhZn8IlB9r0xKzUy4zGvHNAIZA+56SBKIa3
O5huLj9I3TsDoc2yjRvrkFKLP2Xt8QGMHl02x+x3AQ2JXuLChsBIW5EYcuBLyLhD
oz/1/If70qyqhn1H/t/akLr5VO+KUbqvzuMuzcoWnzX7VIy80pe5XwR4AAOyocMz
aMTvnqs1Zri/HnV7WYRx9cngWHr0+Fdh6JzrBIEHYT1fGtaWDqpaJvqYyP3gsGn7
T3W7KJ9cYuLLYyiQV5faHzp8X7Djw5mRoZaqGGxzJERueVhx9+93Equ707lOxB7y
f3Yib3f/rmZnwmTc0oTLL53dyEIh+1Tt5oVqO7bw89E7dkFPj9+3CVuByKKsV9Au
9q3bQKAmlAhPNxEPKKV3Jp5yHUJxMm8GV94kl3tSTVr6+PBXHatUEd3vnBu8eVZO
ZX9W5aH6KpcBY6N8ncKSzyu4/HftIfiqr3DN5J8u5fbx2vw+ADw53GhSm1mpTFWM
EOWzPC3Xa5WGXChOPDBbeQSxoPErJzdc7m4a8UvRWGHc0TUAPxzclRBsXyra48di
11nyGsGECuz3uCi1zRgL9kqoJMRQd8ia14Q+Vtjns5VGWBiXOiNng/v+squzwEBS
/47duRqa9ECB3G2fVMk1fNj9Pxu9Lce5YXQnv96WT+wjSwnJe88PVRUz/Bd45Qm1
hUwrAOVrhwc9l9+mOFDmy/Kw6XlOug6o43sPCPHtMtLmQ3f1kirzKSALHyIAQk/H
7zQxp9KMAPHjDlHMTvF8fkwrzFetZ1l9jPXcBF6/GhyaavN7Z2UAJNAL2cPA0PoU
sG+tAy99FawhnOWtARzgefFlcGC31IdIxUq3zP4/+GAf4kWCMW+Db23u+rPUgs9p
wQ9m/PvFDC/BsKH/Ytj6zjRQFvrMbso5ic9KHEIfV5kM/j8bBg3n1m0DryixoCU/
NVWaDFifd1xQ6DHd4g5sZmbRwgtNs4V7TBXqIR6RlQFgPcndjw8hP6IWyu7EDqQ+
/vBdxurhNVGsi//UcMnGYsHSs4D2vCWsMq/YaQ5EG31sw5sRVrsVFeO4sj5Jn3ak
5yfGFvTEykklND867eN1VOFPUbHVb/n5oIfy4sm7RLpY58bB9wEa3tBgwwfnuqVf
Le7J2M6zS/n7aidhDTMU9AEAYhTwTK6+eCl03TghVDVWwNfahZXXGZ+l9HZiIKvI
5kSPWo+E7jXR8iUbuCo8wzJaBs4utUkbDUtLx1SkcvOboKOvurEDLTwb4SFHJplq
OhZ+ycSVU6iwjpTtJntFrB4W8aFgjGmbYtyMMBSmYXoSm39XvpyAgTwT4bCNX/Cb
E8+MjK1LXwsC+/n9SRFYFP94cRyvsvA2jJkyllIRQQjo+PU2uA0N4wBfAM4N0yGB
+lIDucpioDiXMDEvr6l8AFrOu36MwRDQm/1VLDz+kBPvf8IkXmXqHczn1xYOFl7l
PJBIUl6+Whl2AxuftzuoqiknMqUr1uPi3iN8b3C6jsCFyPegHU4Qw5as0BvwqBkb
gX7OFkBo/M+s/PCsUUDwtT2M9Y5f8j36kQ+vBO8JApdpZvWSvqq0IG1QmDRHB1vc
3j3LuoVfmEAIEqt/s7Lb5YU2NjIJJEZ+UVFa9QcJtPWprdiXLw84yVGq6sS+Ii7C
ikE1LOcjTlt1PrUi68egyT4govx+LS0qSXFdUNY2ZkJXSBKrMu8vIZHRD6WJEsWt
GprXzidkFln0HjFp8hiptTGPoWtg1A4XBu7FoEnGTbIMNmi6miGWoYJF5/Hsrlxt
lrw7PP4Gl2CFJs1IH43C3ASEISeiBZ7JCnVxIQzKUZIg+7tKnu8x3Oij81YFON3U
X+UtKtaFRsrFwH7KXUbGpYLEdPD9po80gGqrkpU4vkspEJE8k/gq4yeL1zMCl0fK
UqAkF38Cwmkc408DKZ6GK5lcMPd1OnZtEZ64ZOGGUw16pOmvxFzAjb7SOBWk10ls
9BCNSELJqe5G1qubwnRWLWqcA/M6NnybqLEcGzWHEsXCsB5EyUswEcI19Tqzz2nC
sn4vic5Sx1cWQgvzl4Fl04JehJ4WPK4niAYXLN9ifKdejbzwoqPHuVaOqEAQI0nB
5T9ocVRnOwTJNMLZY1BoDLQAuTKzfygezzsXXmr0RgG2Fc85i7sAWsuX3pwx02PI
yYSrJpDvB9r82NfrFEwf1UYla2RqboTV5gaSRd2TEs22U+plxZt43hQMDK1s76v0
lMeTwTFOSEA4lDkGLJxZoZ4LHLms4v/Ve9D93tP2VIaWVKyU86TNpwxnzFyvEOMd
99dK/A56/oMClD0jBh2uEAM+wqqOXADFc6Rbzzo+tNtMXplAlugPZyKifHNpH0hi
qxPWMiyQc9beR701hZSfU7I0227utc1bhXY2ezOCYt9joHOkqu+9KrdSTXxGMivY
PGzT0po0GABbX5WUiMxi7yIQKUIP3c3dEPeYT3hn/VwQS5sbRflsWM0OpBKYha60
R/E1FcSApqMzdnGh4uH3BPWekQPeiDNMGrozvHI8kAZ3msf3r2dAgNQLKeirIR1T
/7ZkEE1zLrBivMCTUyBkx8zR7H7WFzmzuI918LwqFpekFvfPtfQzO8HEvi1nT/Ri
srKQD3ZRVP3UbL8VnMVwkOPlleoF60MwKI5X1I62ImIU8yhU7kHPDgWxnQ5ATRzp
P6AfpuXmJrJDaetSsqzGZGEfdZxVKM3A8fptW39gGCkELznQtUsjsIgdA9q2Y38A
k7nP6Ow6BPnAnZ7UAdpBTxVgZHQwnSMrubrNJvpEuOXlenpVuciYuK841UCSyr45
aDvLjxigP7DgEIE4ExY6phvxF6kLtJiiuz93BzyfEF3v56gJm4K09lPCjbl38sck
GCjhROneOCyqVXH75YKa2X5Mz0EVrNM6qkF4Ly1dVb3zFKOK7FaIpmvAyUcSgyjr
iolpyoC4C6Y457R0izzW83Jsf31mxTBgEYgSuaEHEK0NpH0nwz5uRY6ZrTzS2zT0
o2536t7oCl3HgLGJNNEcMeFxb2eigHX80ntC0621n997mzlhoWoVUVDp64m7b69r
BOGho7G/0H/BOv/hWpOj+sxvII44yNEHAwXRMGl/YtWq+DQMXPqoy8v1Gw5oiF2K
Ba/r8pifOc4gur0kbpXNAr3t9zQk1sJIgbrI/LB7slXBqc+cKln0wBp+LtvvBRIt
dRxbU2kTBb65FwrJyyMjrrsk0rq8Od3PoFx6vL2geKKsLc8u3KI5jUnsfYmNlOBt
beoLYqzs+dnfmfZlSSW5O4OhCUSsZlA9wMFYM2RfKEr0F410WM73vcaRycVW8NJV
AsWZyb+KjrpN0U8MBsLBdhNlcaeoxvNHUbJccjE7CqFOn6bcUywP77xInt0d8Xnd
G8eNl7s9Qrcrj6NtjL+n/LTJhfvVS6RIXJPZqlM7rtgkujYox7Iz2Xn6nPoYy72U
9DOK0Qjj8MQ+HAbOLDwP1CIn9XZKNjETZI1AxIhbQvRcWACaRRPJOawphHLqOs8U
TmbjlI0BTURURhGHogF9ZQ8YYHvz28MzWOKhD81gUPwtQ7ZymnlRin3xBlt0G9gr
icINFypOHmil6ZoSqtpQ8604iMSQcDNtKbqj6IqGOQQRRaeY+w/w5CwwaCw8nwkC
cQBgPodsnIMfqQ7t2tagUGYe5lbvtSzIMKdY+SMMJt4nHemT4+Wo31ev8Zm3w4Hm
XycCV76gqQF/e+pRbBW2xYSOm/VWnmMIUd6KYgvfQyHn3Qeszx1MgMDodt2Zh4Io
9eD1ZLvSr8fyoGXieUrPxVazE1oAMOk/mTbbX7wi3jVmFxmc0D3lHXarwOpHD5WH
VrNd0aPsuU/8Z6zhoP65wLudpGGSN8jslH9nAT/5MzbSIIWddTjSrPtAdacZXphI
/jnVi0Pud25kKnS2tLUNd+EvyiTd/9YXSLv37lryuuqd6gPBw9FzmUkPpmfEkpkN
XK7DSXR6k+4MbMatKkFYuTUpqL+NT8Xo/TNdO2rFeuJRTZk1NuJ8xcZsqHe1EMHP
WSu732NuEsol7/xzkgAE782i2za8ANmG2LTgicodJcd3Mt5ixy56MvtgxEFhQR+x
Pw7CbAIyzd3IwsNDH5SYi0/9cnbhmwBIYU3kO388Hh3mEY1sFh/XKrrZR8gPycbm
zSnQhTafF2pJmfObrM+ejo2hFaN+BcpZy/8kVhrd+cEudo5T52kxVz9GoejI67EI
uOtDIde+U+NwlojVg3q667TpZC3ft1lgogZlwQVQdfaFlvGA9lHWdh+iwh+R6E7b
nsmWw71W1C7kNQSzJBFBKg9XZq/GsP4rFiU6aITQafj5mD5xM4+qB/bc2aCaJYBO
6FJ9laNbNFV1zP6x385K37PnkFUfmff9qA7C/igzdmRVVwCZ+W+t42IqREm9Gko5
iZWfLX3tF1Tyg8vuVT7NQCbgLRDJ2OUB8NanPeD/G5XjJa5kE8Mbf9kARgoc3uvb
D1Nc/2aueFlgL0rxxOIqhZf+go2je83NzcKcua/X0EPrk7SHhd3yO5sjliOulbz7
0g7Ms2fJkRTJBZcbNHaSFFRmK5gWkynTider3lqYiUuE8CfOc1T1zk6mVYlHF9Cp
qjhKqllIcJfhMu8XJulRk1zSSDCBkwGpjKGwAyUhcmz/AocTt0m6gZsL8fKJVdF3
AquGBcX6/Wa4D+DOUOK0Xukocm4MI69q8qUNvNO7EERQFy3LxWTrN+Zrj6nQBkyZ
f/hNCzfw8StgHA0Gkde8q87yN1vihKWHwG9j1bD2aEA/i77Ithz16sz29PiLWimT
f9gZeCEo1q5302jyl5En0+LBuhhxzTy0KFdAKRzOzW26S+kySqjWFRdgLQxnfDXs
tJq88Zvmdd/ooQqHKUfwiutGGy1WSkixwoFgJon6gfxB/0a23vXzdm4kxKbJu0BM
CKWmJPxoV6BRJvUo/m11LkYTj63LTu3dCojKdSh5rrC+D0okOLdsr+x5/0EYo7s8
WD5wVYdEbl6bNpVYMLIShjeiIMH5CgQeF3b9g/nrMrMqLmVTzWdCeUnj3hQBh3vo
e3tMmSEFAS4ozOoVs00e+l8fI+RiK9NfqmIl3u5UuxEWKDU90rMEBwPa8xNLoQ4T
O8oGajpzcjX1AAvPDjpn3dsKWtlAtR8wI+sbUNPShMdK0JlyJbjuKNIbCSN5pFBd
Y3lCbJKP2/+liqclzzWVxkip5cEjO15mmT91B4Sv+cTscy5o8+tw+KwVfV89Z8TV
I0V2dvQJuCyjAqLMQG8tD6+KNFkYujALxB6bjs6AVWIxgQZL1QzpXyyFkWU+XIVX
qYnOclJDhUoTAxJt8B2lo7L/4gu3k4nO+Wnd38P4eNnVyeklfX8lYT0MQRm1i1n6
S8W2ZE8cVSw7ttz9PCJefYeFL82ERLvNEpp94dNV07yMd/qs9zjO7sv6tOqvaY47
d2LCv5sQ5Az/kKFxrLJUYA541Ee7t6wgj8T/QVI9i3FXJtaF4Eo9sCUwWnLs7/b5
0tw8Wcqx6mc2zrCI9rjIQ/68gzmwJTtXFmWIeJzk+VxaEFUzIsyAiRfyz7xz5fYr
T0GKxKQ0VtJvUkls9V1/ANm7OFxAOYqzISKpu+xc5/r/51gjk0VHjIPfXofSQebO
f4H2IBgt94OgaPCH3DI816OKAJLZdh3nj4dRFZlrc7vX2zP/NX7aoATjDyaMu/QO
89rh++KGSzoeQPE5lRkpEKAseJ5XDQOrvjN/aurF7DwDxK/ZcDoEWli6tKzfwggW
fntXcquVu76yb/x+5RnLUYPjLQupeLaDaInb0Ed08sQM5MGxpUw2G2ny8/dBFYNv
SprI6xbXUj7N1D7VbPm+uk13BsBGzMtbgBEAqNy6q/8IXdBDX5gASkIw2m398Ccg
6Ehs7ItRIHFBektr8Hbi0vOBmqL0Nq4NbVFrt8ptmenVrK/w3ioSk5yfvf09if05
Jb8sC99HsVeGUnOE7OmEMpjF403nhEe0/9C9iiUmb2gqDbjanSFpwv1x5ac0CmFb
gAnOlzbeE5ZhjlW4IFheELLHvgpD83bc31xAXTo9M2IheoZ4C9wbm6m5s9gv33/F
aXMbFliiYHSWTqTET3GfUQpOM10msN4cOGhpxpgYVLYJhEJwRGtvTrNH0NC6Np/W
zYL2y5/ZM0clEKPXhmM8BrZhaAuc54qw7zzgMcL6mvc5jCkxfCgW6FLaVOMakO2R
5CfYcQt9MTnhwWiWkkVdRJx3HmrPAlbp77XL3hR2qNyiEuZyV6e3Gv3lqdOJu0F2
avbLzB/R+TwY1UTeNipqoVNTZnalavqsaef+KEQXn+GuuNe+JWGl5FzO11gYwGCc
OZibdKYC7NwjmxCMcmfW3d+KFbhZkdxiEMpHSYXSbCQ1+4ZqymbgmIk+izy/yNeN
XdWeG0a/SvQ4nQd0ou9f5799l4fYh6/C5SzuOdl4dhXu1KdPRZ6rMNuhbqTaik5h
AcxrZ6o6BmPZ/D0N2mtGrJ2YgbrgyF5v0CBekNA8Dt8JFRBEqBAt/l4KyLMCMn4U
VPkuHRm+Pivir4R0Wlr7xN66m7qGNxelV7Uaw5Ch6x9XiUXQkCkCFL5g+3i0aE0k
Oj41eAfxrqbT9U8Uc6X+1rlDMIBfyZ2jg8xnOq8Z2y1pTwFGcTKQQvFVCt37miT5
um1qloLjl0kqNt46G6r7Pes8A6W08uZgNnzklOVfBSFNIRm4hFl3ymkn6ES5L/PE
9efsnTE10CaB9QXVeOBwbjwp9CNibCuMsmsujAzxEnVoQQcgVFgY7UENVERUByZc
0Bfc3LlHM4xqiHmPR0Lqzrx7ZFRyqhi0eifotO1KJRtGXzR3GL/tvVqbWedx/XA3
qiXJQC95x8qPhGGjOJVlWtqZoxcTsXxiCu2oNnff0ipmkSfdf0S9vhkq28+3Tk40
bktCWsqHq8AheJupCXzaDLiAFOVo9hzbLsj1feZrfEl1uJ44ncQES0neetyrX+fL
CYzXAN13JcUzWFyvEDf5foydnj8gbe0TpyneSyLRX/wO2Gba80DuzTUH2NMf7m4O
4jfa6srTAQRzGEQpH8ne9x4TxAGh5y+Gise1Acsjh2KfAgUurxn2+CYSiblR5llK
9tMbEepFxtUi/38PKwNS9dHcg1HtrgPaoZ9yndp1j1vesGZ5I78hr6CHoeIfWf93
Gjz2/BBHyPpWwYUshc2IqHrMFUvVR4S69/oyQBYYsjVsKHEbzpFkZPZDls8oOHog
/n14uagV6z/D28Qp0u/1/CUwAI1G3c+91uXJBJT5DAMsXZALyAa/tbfXTJvDPtlA
mOz3LBD1GfdrkAWPYYVxqExoEkhSYeJVDj3ez+Nob3msLO98Qqo+l79YGa4KVKq1
YWLobMlXsMNtutTKbMGPm0+vcZ62/qC4f+Zs/Skc0dNvI6ZRD0YcBhojj8X04y0X
5J0Ktvhk/FX3Kqze2BMb/coR8yHx6Lim/tU+mYProDiElmnH++29H8fsrfhm4D8N
A07K8R+rJcMnIlNsboh5YYkarWEOsOZAh8dYrlUZyxhPLZK/VA2X7BHQ7m9fRUtb
3FpfK4kSYiV0UTQq7uhQ97UQc5nyf56W07eBhBoI+1DYIdLZQBQA8tV/PoOWEUt0
/2jgHIDcFYHxkJOBJAJHmeOGNKAxy2I7cEIWxAdf9g3egWxTGzQrOM9R25kYeT2/
i8judK9+He6oyV10CeEgyZu9B8dqsEiTfIS15U3m+QSJJ19NTyandovdc89QQNwk
RIrZvP3B4hAcF0FQmdOk3a2QhsSrxdYaP5I9thoV4++LE3JL+L+Z9nexm2f2Mx01
Pw8VjUIbVBBRF1NmsQL81vpd41kYs11efMHn4vEzyHJJrHd1nzTqpgE1KGSN5WTS
w6er2Qa1wH0n9Y36FLZ5Hy9dTasxb9xUsX7l+ld6JbtbVsTDYgXEOf+cKziz49I6
/+cg1eXcoMtPWuynShRoF/X+wZHoO/oExGlwfYRBY1PmO6XpMFOBkiP9j1wewh9t
8G1TjYpNQUrZffhMtf/99GnRwv9vEL5i910dAdfiws2yfUw3Yd6d1Yq2/PClvn8G
nbFKeHbi/4cfiqUmlnXwXa/lXVShGDiyxPQ+8fdMk0uh0xOtW9kWgIHBWqfR5hfa
32pNNBjqyQu0tlRF9rSvtv7UVmVdkmab+W2F0SPo0fLGktE7wXZlte++9DysfSqF
wu3C35zxLsDdRceCKhuPZFcrLeF2G3rUpMfUxsJjuaLFxrNPX+T/5Ao9yFV/WB9U
DV6BnbdZl73o8wnBalHGBX0yxpttffgdemOF/iCejRGoOlALugCX3zUIA0KoWlFV
944jCda9whGGlpcdu0vqYkwOK4dU8yTzh98vGOI3S3vSfV0VUn6CukQHx9lOtoRq
x/uwn5KA2opmfsVudwCm6uEq9aK0ZIZdswimv/97XolFdHzLDNISaZ63ea1ddVA+
qWjJUZJi3W0yWlAsDLWIat8DCBfXAaPX7csjH9DDTarYmbSKYI8EaCfnJdItbNUm
Gf6VwDPnYMXzC9HWbiK6fOlB1Qu3IKfjzpEpf1mh7EpZUX0R5tSPOtpmWNQ5XDE/
ad8iIZXPmyJGHM0Jj6xgsCaCF32zhot7T+hJc+MP/arS1/Obkv2DtCvwbWh79hs4
xZxhHlX54ye+kUM7ej0CJuhBFR4Aq+SGuL+uNlJhoPu+GjZIhs4xz2KcxfnwWM1M
L5syWrpo/sPUE+jZPzTiGRRFN70JURnk1U/2+TmNIse51pUSIcsS/buqaqwNvl/g
9edpHRsOWWUqnrCAsT8anZrvQC+0Po8tC7L9Ojyr9jJm4FePsJj9gFPt1m/k8L61
HcNOUJAs7LebixutAXHEEuQMrOk9OOGQMB+xq/D/OMt0i9xeGFWRjB7qf7PRaV5O
Tf9m3JZUCLGbpsN9G4+lWzTXWlPibvge6LUP4Ky/cpGshu0cTmE+6kS8k1fKkgvH
i7E56p/ERN6fTMi3weyyjHMbrXZ1zWDbZvQWu7vXkf1LT+OQWvpsKNsPBNQjDObP
wef28FsFfvJ8BYHvUmL48X++c5yliHjuOdqgSSGhezYXayLxZGRnJSikGRAZH3ET
NYm9mxisuGpOUsAOh3Gi/Vy2xNsBns63DRkgi+dlX8bpKmzvI3V/BXMlqrZjEfk8
L0mei81mtffZDvSiRLFFCN+AGMnI/BUMb/KEAVNyhgd8LeIH4QjGpcraruDeo8Qo
3GorL/Z5ebjqfXW9wZbLxcBfhLodG6VHxDL/lb4AOeGZo46obh9GPdq/uGbAhR+d
am2y6GPuo7AZaiM1CblQFb9hiLnc8WW2ZW9NzkWkYxireDk9iB5azJ4JL5boMqQj
L8fSuNCs3+1mwFPRjmP8FEzqXxCiEaSfjThU1ldzP0EO/0bINaQmR0MadrtXP4j1
CSllt/FcTAwxVeH8u2uZIvXcO2rs1rDer8mS//kPoKXbwAUcaaOdOTEw12rbpJ93
4yN7CzpNaqFOR8zXrtQN1bcENSFb47VGlzsQJnqcO8Btm0ZzolrQSOimK2y3SYew
eJRrpqauppplgGgxQWc12Lrdut7HhKKdEFG7htOiNnIufHzpY+G8N4ATOGw2Q24o
CgSqCLfe41bucQ3YM9U86mZBqwBi68mupjVXTub6pwsm6JeZom6Pt83+9FjrjR68
b9ELR7m7UfoDJ+WVPIL91FnlLVmCWU9kllXixj0gjFMHwo9Kl/cx4QcfqjigGjY3
MV1qnQV92omEn+EN5AGFFqpPeKYn0l66dtnMci0/dEioFBXMoi0mZFRyuZHWkC8e
xlkBH25He0/zRg//XmuGFERwweL69SLJe56DbUUV7zgfahB0C7CfkeN27Zjw91DY
JqyNyOMoEnrkYm9TQYO2Ii2BYBw3oNCFKhNNRTEweIWoALAM9kmDat3MDDcoP2HV
nBJN1gx8u4OD1GR+2vLVwI7qCOvT20Osk3n20N4LS+CiuKV39AACDl8r871gYT6W
CWv1Hy8FlmosGKxeP5I45FCBMDb82blEAuRnPyrUiRef7qVAuLS2periOurdQFiD
Z33WL/JNKjcRKYnpL15TgazN165loKb1Ys+wQSgnIZV3uWPIT/tUWdxOXFMIoECd
5UwxVrbrxbYPTYFKK8Gksun2d92rW8YDvQSZ2hRtaPhTHowG27VIxfjNagNpAc3T
Ss9epGa0gJzpLD4rq9/vCrrvxisFWQ2rSBRIIpSHzLh7GccPJIivPTTNaPteuWEN
ixL6i3fgbpabt4GoKC+5bH4jLk1jggH/i9MGQI3k5UXNqcPRbwXxwDwl3dGwhSiH
9scKZApdUrX78ykB0ISm1rQJfalDHPK+0zpnuj+Uc3ntAl9081UJpS7ZGbixbvxW
lh1uZ+02r+5vFK/R+WGLM7+M3NA0/6MxpWt+oHdHTRcrsgXf8eEdK6yJMVeNWGmp
PXVKI1xguYDoods9creKXWUKp0jS/7gphzO71+KdsksgNuIEJPDur2he9tuZBglB
MFHtozEQh5lIpll2v2lgrQA6WeHFQgxvLUg8mt/6kp0ukxc3oU1xgPj1RaxLSpYF
lXEEMtfVFOoHgqFeRUc5p5cXY9EEqWNdUXNmrIqET2sUrqBpyZtEpujzksjKKoZh
DWeoxUtBHWHgv5Dob0ag+u8Hx0IPMyEXQe/bLLMi7Iz7rmxg7o9x9TnX6Ft4o4sq
wOQGqfEZXeZGwaoAqc0A1TYU5sh741hyXdfEziFrxD/q1AA/MF3yXr+bG/YzRvIE
HsqZKxU+uDgwLr8XbSko+3oGtGyoZOf2AvUICo7Tpsx+w/gUPXrWJX4D8AjNM55m
BMIxOUXQcZKdmJ0FWYxWoZo39JNlQyNkg7mzy8P+zcvaDcGKEPUganATuIYbDcLT
HmQOz+0GlWjch6SyYRueqAJoVFIgEKHLHldzHhEWPbww1b4TnthMCI9FtVe+DuUI
AuinjyAvqhvkvq6bdPSNJNwZ/Sv4gK3xsYztJ7kV1WQQ2zxdfxBqZkpco5YABckj
0yexqn7/7qfHvdf31TjjHDdB2CnFxH0iQDfT0p6A9Vcwic9ZYhFBRkkQa+NysESP
7d2WTNZGW+aZ13Mb7xjYlrdLNdwyb/cPscplRLq7mgwFNeEr71FEIjDpJ3vda4x5
X4aDgfzpCmWiJQuM28yT28UNFKSOuTZEvjToBv9kXLV5ldVBB1naomEmhMitLEwQ
Ew2OsWpPl5zEgeYDMFgQMAoj8fnhuy4MHUn2fsfDMJmex4/GJWkl4Z7q5dYSk6q4
f8t6hRCTCOBkf8usnKPkkvB5t2HlLFzocy2NOh6uabJgj70jHqNbiRQYODzr0KR+
5Ee1oDNl2SbS8AeIpjjE2lqGOuh3wCuoZaDCTzVyXAqavxqEB5TcQZR/bcMp+H9C
Rto6h1BD/2jvyERIpUyqJLwl0O3EM3UVEkCgAGT8qyitKs6spGoUvjO65C1TE8m1
TIR5Z3M2pewZtosPmblrB4X5HV/2a2/HNs9jC7kxyYn2CezqWqAOI2xG7BzupuDF
2sQRoHK03tPie8LPKw7gry8weI3QEkep1Flbq510IZ77nVoKv9664fHK3OM+pb0B
r12EmOQBfwhYOHq++RgqIAUw2mWAaCWcKyLx4XytWMBJVDsJRpB22xdw24Rwhyfc
8RZf18xMlAZP5EtQcroraJBDNVHE1v0qvpexNncpvcmZPqkqHzeKBP/SrjrMuwnO
hcdxrpjhVzYZavbORPPaxfD/9fp3ojh8yC8aD21tMbL3X6MK3Ei8mQ7duUyFCGxw
eIZyqVtZYqeIo3yUt765WjAYrcEmirfvvyhb/4cTf3nXkLIXY9Wgk9EeY1vzGynW
O6Gm9SE6lz3dFrAGalyDb4UqtQx8c3uIHieO1uw02YZ5x5KEA88FOkrjqKkpXsf5
WqIuhze2bcotk0tTq77JOkaeThIEPEUTF08+6MItr4mjWgJiWU8GGrHKH1lkO4RZ
X9s7TUuBaQHF0gpRuZW/tIkni112py988Ki6Qdp27HktQ4ZzAbvXLqWFio8qjcak
cb2AQA4b40euHtOGO1fhbGCMa7YGPKUwZRmWlN/zCyFCp/o/bjqWAWj+dd3dBm88
WTxQGSmlg/IajNXYhT2zI/77n2QFEBm8XYLGYbcTHqg6vrJmwR4r4djNXmA/isIo
YsYXYVE1JoReqpHLMnVnHCE9gW2TQQ9BObLXdVe+jwFgiOH+ZfUIc+irLvNkaJxg
EaoAVlMNw1zNJf84Z3ZLjRNboOAemzRddoloZuHzUzjx2qq6Zbyhzkt2RhGV63p2
Xp/+TalWoJZRy4lb3Ty/tyNjHd/J3pJpSKmUn0jg3P3CUpzptGHIpMi69YLslOWm
46jf9rDLAHIPDfkGHzWqnveEGtRO0VPqaY/iyJkS9mhT++uxEpHM+VK/FaoarjVb
WJ3DAo51Rb/owpdMuvW0t5fYFRcPWXkQEyF9yaDOt5qqtJp0Z2POnH0n5C1+7+8O
JJpkdrUF53lzknDTnKvUXo5hphn4uSDzuWutN1HQBxH8l7IeY1XMrkIt0BhLXual
4m3/DBTzqBX8fDM0PadViHS253aW6ZzdLJb0ofETS7rjPJL96erzK4J16YU6J8jP
RYBFZDqNvi6CJKwl7LPaEBGbQgREqgwe/ZX1295Yq//evf1YN5iiH8TiF9c/uxqn
jkxozT/fLfrmVePlNcT/nZY5dzGIkq8ul28PMLnEFao/N+ZKifKKiWJBVlfpIa36
K5KmzVp8DZr/oj/psjlE1rweZ2exJrw6aW+BISXRwv6Pysx4irphMCGejbAWwRxp
ThfBs9JYn0C5KNlgBfdY5Wg6Qoe5eudidoRSmd4MemBSuAV8+JGUqV41Y6JUFSEW
4gfvlQNIp9aKIDmK2OIn6wQ7cghuWnHORDDAoHhCVtnxAsLpc36er16cyGDzV0/J
kJhqOvlKmRCaAnt63YAXZHs+ePG/uAZmelVm7YvFJuTTW/h93dU0MrUd5WECSBh9
Afgmf+JZg+00RA7/P/t8a23YFfvHVSS592VccOYiiOAgdmIIc2Rk4uxlXq4Cc3lT
BSr31+PmXGO4klXsDXqCeT/awPUTH4mQCQ6k87Ia6hluNRqJvsPFe0C7juO9Cy/u
scv/Yyba8jQ5r4lyJCPKak5glJ8B3iOj7OzwZD5pygIsdvgD09Sk8K55AZai18NI
Rz3Vgnw+WmI78WuTAD29RKhuMJn8LrkzUfmU08ZT4esLGoYX6G7pyim7Moy4uhEI
lkmwAyWz3Sq1GHRvN1gvMfp/qut/aazGuSKPvhYusSeZ9HdZHMSMo1mcu8JPQKhf
c8jqRIOnYVRWfPTc1TitGiCZimN5/ScqSc9Rsc0szuqcXiNWjmcLT4G7FS9VIbaO
u/d25jEDsecyOPybp0WqT3xobcXsqBk6i30LG25+rwb6JINqw9Kl7pLJ2cPrJoBE
eZ9dhEvuU/acH8IWv5eR92yNyk/u3S1fO1fOaleiz9NpRm8+Zn0LBnnKuBW0Gb0w
gyixbHze3i47SG0O3uX2dgWGsUUdBTEAR+syT/F08N23gdxw6O8pe5NYpw081VUy
UeORdoZu2z4hL9YeCEwIvxM4kYWTjZQXuj3kKH40WoOmQACb0NQ2/3YdZ3OIKtyz
or3kh58CdQ8uhve5D7E3bKmhhk0XPKusmFwWcyjbXLVgqiVqHZG4YmUbSh+KH1/N
QCBH8EeRo/qThLcLKaJw1+tIYMuJUjzEwBqoHtJ2DPv8bdWEBSkmdkrmZQY1Ra8w
rL23PGK8T8T9nBOZ2Bp5bdAbBxp/Bo5JTBgIwoZ7r1Z44yXNWYxKhcx/NiP/j+7d
CvICcHUVQDIqpNCe1hjzxPr6JVa7g9DMJMiSwt36WRBUZc3+I+CkxLGNZ9fYVe/2
z/YDx0RcVw2puliflhJY44A4biSCHq1gtlChir/TEFCEZzsgtm/WjgugnRTFQbkt
0kQTq5XIdELiHZtYRY9QnbNWTrVSLXxpOE6u1JLpRzu5c22YWZUW8YWihwVWrz94
xuxafmOS5cyWcezHGD63B4Rwmd1BDVinIueA96OAuye66V0dOv4E0r1xys9sMDWV
vEI6scs1wRFOyFNrc3fq8NTLzLwt5Yaydw1jWHQlFnOWHW1NgIA4ekgu7xfdAM9h
iXbYPPthFeRFlHPRWt5vVCprKdc7Pt9NGwJULIeTtp52xDi3oShC6a8Iu3TSyMiI
MsNVZ1nXHS+ThvY2SSWCu63gRNPUcrvihGULHdQzpEnvNubUJDachZtxURw5oXX7
3P0Gg6I/e5k7xhNm1+PaTi7lFyrsVGNOvSsvlvFT08Z5JA5ydS4l868tEgLtGbeN
RzDV7gmu5ufjEpoK2Nv293Xm1YQs7JXyXARlhKZTaRqkRF8ihEFWm5+1BvG9yG1h
aGIPHmGnSdHMYPOFi7ZHInQUS4qSr1Cy1CXxh6509S72+uhiMGULksALZvK8CdX0
9dAaKWKZtm4TDU6y1sMDxBte0VbbSGjqzm0N1Hdj5ORxlieYETNPrs/R9a84H3pA
zZxYaoHxBgWUQVUbvACE9lqJwUqMvHgjNjhRpHFSZpeJ+zRb1+YuKnCB2ikgjN1B
Hl1cdnMrNThmu28MRfhGOaoARFGWqc4ajZt9nc6GTPnoMmTgQH3+eqXhzIXkvbZG
KnaIMcAYlMimcebOCXbTt9wV99eha4IxniwBuKtHM/x6riQf0aGysIkJ0Fi2k7bf
iVgj5AZwpGP/1I/A8zpd4FILZfZQ5CHxR1JsivMVq6WMvnpigmXXtE73b/prYO7l
f/ohJ0GryLZ64G2oLtCy8zgmdFzNGr+aLwbkbd9GxL+Ns+Oe7u17COJnuSHYYBM6
mHvKmgtOBM1h1YHzcZYDO+uup1DMSJsYUVWV6FtsSLgW/2fGUH4yqYZT/5+zgcxp
ytBQBmHRrvez8QpEED6x0rpTx4/lMzVtaiK9FKPV5WMB71QJWEdDnxxvFYWFbo5l
4AEG+zlUlDHdee8i7PyWjqpK/gn6gtVHeSOPqhEgcFezs1bjriYnR/gesqI4Quh8
hhA9luDEUij70bJA9Ydtbtp3OpnXdp6xk0WkDWsCtFAU0QX8kuleZ/Ig01lq+NDc
PV0ioF+MEZ0a5DWQ61pzGoDCseEVYihUYt9rLAZJVNFJp6SdNbwxEQw8ubn6ScTC
VP68fsBfKf66RXgWvuzOo+CxPSzyN8ILugm2W/pKErulHZr8Zi8H44LPkCi0eqYw
oeqNti4oaSqRkiNQtNKh0UDz3wj5obqqjbiSELpeJkmB3ruSDZlsmO6311z0Lttd
RpbtO3xZmRziJBsNiO4IwStwQQre8Qpq18tgaS9is+s+DLxZJuyQJTEmBOOEFQzi
eVHHe5yaooK21KyNG4SQFbKtTpVaS4adFgZaSuvoZpMdnGk74lkfajdguin7a1NR
he1er4DJEi9saUe0QnABXLJs4Hzhu432AkrjCmUgHU9VyyBP4UZ9efnD5EAvIh9L
dopcTJbgER038p4kvcShPj/1FdApWozYnHNC63d6q4HcfZtVdaQ3sJ5y6SioEj57
/a0WclS2RPFaeuL4mFyFnY5lOX5Iz5Jf1HmSzVNPDHyxw/ck4YO169T2w9oVXuB0
JLNNaDcFLwCa4+Anr6OnmmmH68iAGuYaMkeunUqvwtrEMFUd17Bsf/+219nOVFmd
pF6VEV0VX5MyhCRiRLICFKFwVD4u9kEDakbkS+e0hYuZjsVz0V+Q2ZNi93BVMwl+
Pl69TCyuua8xcVVL+r86lgFxca3XR/kQEAQFvfuhnWwfrwRQH1Li/j46b2nTxFpE
Js4MaWpY19EeqMfWcjegeMtR/gllMp7igUv91T4oFWTTssoc2ramA0PwIE+R06bd
UjvZ5OrYmq5vj3aicSWnNqMJe/RwGqg3t1hfd7D1fIIQzSTQLqPmTElJ4Annel1j
U/HnJf6qYP9c8uNkQa4IiYsOwWOaQsCnYerZd+RBQxMV+qP6PCQF+xMHAeXCNWXX
xhU9Qq2Dw7nkP39YqrcTYAGmV0RI2y84RQY/oiY3HkA3CH6jybj901V8cvjkCnxZ
acY8pG/c1sj7JNVe6dEJakgqHwESgx3lH+/Irk7zMq9vcZXRRlDJnF+rWG6P4c7v
uBfKmfDplDCpCC27Qqhq2WQqN2zRz6WMO8SwAuBrO1fM4F1zCspW/rND5KrMRdOl
es0VbQWnaA9DocdJJtJ1/4kijGr8nQ17PMjowP0Z4wcGTPIYaA3jtXVutM3I5YzU
k+zL+dg2NyQnf6NKA3pvX/UY9lSskyxhMaPRY//ybO5xtn39KRk+rdPbxZHVUsN2
ZFymuqluBLPR83tgYE126WArsUdMaufqQZNEwxGUJA/tG8MfyHllxA/tb9c3a080
kKyiHcU5IAqDA5EE1tLUC726q+dJ3yqqChxCnidwm46JcMUVEnmo5XelnzMVYOm0
V0J4wSjk2uS1GV9DpW1WE/4PKDbQrgmaixMF7s62RWosRgku2q6ftX2xwqfam1pP
mAqrfMhqYlb3kgvkerNzVnvHX6aRn4OSBZtfIU07ME/yN6LGfat0EWkMoXSovxnZ
IMTheNGT7As2HnYZIfsTMpOXBLsbkaPBwYyqte+Osy7Osbp08j6I3hTTgwAUixXs
0Min0vCkB1+4dlAeqFiEmoLVchWGy0GPfohIzMMwhnQCEbVSyyJj+vD0f1LMo2yp
PAywhwLG69HY9hEl0D+HFRper4z9EKaYgs4OhZTng1L0+paNG4Id+w1UJcU1hZZr
outPlIrn/SNuqz9WMsYnGklDa4JRUPTL3Zs6ngthOq20Q2g71y6nexjpvgOkBacT
P7YHGDHSn/Xcw8K0nnHiWGVsyLbGT28rocZsDKdExKbGLHQBeldD0NKIL6FJoxUi
ax3dN7iHwufXLKmJTVn2CssRZTsoAHIsvx/D1cK58+75EyW07O7hkGCzcwFpvwTa
st6uN7p0Esbn5VJQOCWcY4HB+16Z8J2/KxmH1YXixslorg6rzstRKfykety+2yn0
//oCEQYfyCdCr8/i79AGlC0jC5UyzQnAsvjABw1KN5KpgP911lWRP/vVU5V50P0T
B7gw/0KxKE88stNYLm6XBvDblVTJvv8nhIHQmvRhLTmU9DpB7fQSS8dWeFkFHRD3
Ybz6GfHanGt+cAYAD6kVOko4Ptc0t7jjh3r1b35wMZr2Gy5qS6qFnhOooBf7Z/SI
PynX0k+/vgiu9PSO1i4ifdVvurcGc1L0uKugf0YOYlOkhLf91aT5j6+3c43xSSkp
OAKSQtQrZcSE6agCbLuiu+Y4O/zXLWzNiQI2mK0OXQMXW7jC75shV2vVmilCyGxR
wnBejUuIEbY8lKAlC5YWHkfHMjGAndxYKRWS4tdAAklRUTK2mtDm8WcVVrZBsCiT
un0WiQ9UDP/MGdYKjYhtDYM0+MOwcvFZpFc9HOGh5hsG8UyMkDl4w+Yh23fRGgrH
xg/dtYGIZ7xyMt6QJcnlKvsrBpcgqj+/tEsKSn4h1OTrJDmMeu0R2ajwWT8jVLDz
hjdOPdsBFyyG/d0OrM+OKIyTQ+U7ZLWxbSWquRi262xwqm/T6wlhGiJVBzE6aKXC
koR0uUm7xrKbPUCckJCabpqnxZzp1p11Xd/H33FSb7h2Bl4BAl47pOJ0q2ZHKEvG
vU0/U+tHKe0C5WaoYS2HSiNEi36P7fMUivctFmtbkv5j5+nvVTZQ2hKCBKIvC63c
+cAEKkZs2KrYMHO9GhYZRAWwcfsVR/n3eqiTuJHATn0qojmo/HW6Fo7+5QDYSs7F
o5Y49d18r5/SPYe5cXheZoXrlwtnS5L8A9heX8015RUgsaYEguX2zTWS5OntSLxE
MdQOfwy01qcZ9I1P92m4iu79mFM7IVzEwudOMO1rGUCf1AIJlWsguL10oMVL/HKM
lP+HLSokzHru8AoCBGONTO/wN6udK4LDqnENU1r5S4aJtk+lYkqd78UTN7w42za8
4CKNKDp1oLwPobVgL4G4Ytlpf4+2gyAJgjyKlaSQzVd7ynL1aNJAnnqu2j+zFTnu
2gPVZdBIQzSAFgzJkz235e1tuhTQUClOps71o8CvJ9U2ArXOsPCDGD8hqD4j+vDW
SSivmVnts9Dg/i2x6EPdTWPGLbVh9RPxjLhCY445VF/t5zwFBM8xxjz9IVrRBt2u
wNLtTBmGNgmk3u3Fhyq/ep7t5rQYF/xiJPzk5NLJpeNuMg/2pUs2W1bGVSaSe27z
nb50bcTyyFa/LZMEHUSJDXTMgeRuyxbEx5G8QhuUjIPen4JEpNaRjmG5GiHJAU6M
114bwuoAFEeQRjBs2wiQY/zV59QlAhaIy/90EUZTilYmFFtkyG63nhCLXNd35j5c
8yFwOplQbOF9EqvtPrTJUVe3kEhoIpWdITgcUbp2qsdNgY831VS3d7lb+0dfYRt5
TRRhgeWOW/aokXWRMD8SUMKRIouXIBPb5ywlOagJrBCB+jXDJ/jcmamCvpc+BpaN
4O/8Vw0igmGPeHjsgw0++0YAGeuZLBQSs078sKMyzH6dDY8y8u8w1UnvyX1QOkVQ
tEvMTN2oqBYWADG3jih+R+8vO5S6cdMLaCCFovCKzBABWA1veO5EPyqMhqLnLqTQ
EzgHhqc0WBLJ4t18BpbqvCGhoBgHN5wYXUjyCxXRs8qE/gZ+XYouIN7vZ7BTmOeP
3F/LhbhottnVxZwjXF8kxhLD7OytCZcOa0v8OXC33Z1RvcxM+ChvZW1FgYr5VZuS
DkHFNLePnzfRuYHOmZI3RRXhKj1NbXl5boI9yQXsQxj5AZBXChrcmBiLujgbi0DH
Sy2vAk3ST2IqRcUWE2VfNaFDaB19do3RBKW5SiwGxp4aLqCHHJv1d+36IJ2nGsEn
SAGBUjFflbQugaQ2FAmtbLNx8SigHtpnUxBdT+7XL807cLCaptSirRd8lzKOtfmM
Nmf1Jr7dv92HpPsG3aM2bqyGllRnDYuMNjTgBCrBqN4pNJAsNAcaGYR2Qp5/+CbA
+ogXqrIFrNNS6EoR0iAaWt9dBZtNPWF/Vbn88m5NhdlhN62WzklGxLXgbtuZje5/
//slK6O/xjjs8ONZwgJgK8c8xU+0uvq/sGSjs6zyn25MMaG89G4/Su8wES63b+QS
UNqjYANgJTGbbi00AYUo4pOpmM0cGrB84YxhzDU2grDIZBKpU5V5IOPrKtcBLrey
Uq/SBx8S/jMDLAdrIPBOFXd7j7rKpN5Q6IYit8OYRjexzFmIIVDUloZnLEv4l2Ph
AjC+Ld1+mJaDSdUjBd4ogdYpbGdu+5UwfcDE/raYPqIuEIO4cvCkMnk76e+AdkaU
zXLIog+NNmO288Ud4nohGKy2vkjFNldBd08656F+XJ/GL+uXMgJ2b5aj/Nk56AT5
iuBdrZKrRFmhea0fs8qqaXdWTFzk5iOlCP2FYsrz1iMuvM7wos9MJ/GElgMQK1mN
Sf2pThDh5N/StEFePENrCirhxum538Pc/SYNJDCBhE7yrQ98TTEMPvsOTZIy+HUx
g7QKmU26Fy+Pa33g5qBgMdPtMRt1cOpmUI/4QxFZQvoYoy6OKA746EboQ6Kddo6l
dhvwwd9nA878ZJD4+is3DXDqGAXoOfHT5qofbkZHQNlwpDON8clI8VhnEhstie+1
r9mGiV1QEgwbGl2F/aenJg2zrO0RZe/PjropyHPZWTheWxdIkEnGBGgvYktVJNCL
VwGwyWDz2KepJ05TgWPpakMyFSyupn2aA6RIUXPPYAlIGdlgsCTXkXhmUcrzBbKb
V9HZOYaCi6dDRKKEnU0Kh0b/2LU7XVR0nmv4c2ibkKKX4FOYtzd9dBQJl/7Ow98D
ZaLfH3gLvEGbqXB6b8pUWjplHpolupNM7IsWQ3tKPj9UablQitLn6FgiRLEZROKn
jhOy45wNQvj4Y5wRjv/m2THruPnq7JRRv0i/s7T5cGp7c5nBBFFKyj6mcUlXaFrr
ZQafhPHZFy4IY/s5yfXNsZ3kg3Kos8mWuQtiGIA5cuHKqXqHy7QtBXZArSkpVGZv
pSQjlzTfexzof9ZPurThciu/6YygT9BJZJEauTrHWyMmUqnKTAt0kqSZCb2ormiv
hwItTa8TqkouQ6UVC7UR+wd5ByUDAp2onRuevDdiDL77OIzZalXPxxpVMUNFnW8V
bnIBKealG1Px35Sg06sVIk5J/cWtvVV27W5DEaV1LayZU7QaDTyzUNw3czF/2Dg9
ti1/7f5vU+ILg7AiLatL2Vfau6GCI58B5iMnF13wmRPT/yd32L0l2h6ASkgmFQYw
KUbs1GfwfVDyyZW4OGljFoDsG7oeQVQhmtyECTldsPTfaE+tAGWfdZORImqzG4gZ
P+wZJx4IQan7MES3O5802k+CPqWeda4Cf9Oxgun0+va9Lcb5U6nh/lhv7iOXSMY0
oXmdeE6UIdBI9qZyC+YRIrrtoRWphssE4838+MckQMzRh8DDH27/fkKyXBB5+/9p
uS7zAg37h8yVQT3OG4KRNAirX3qJ8NekqspM6rfqxvkKy31raKU9KktdaT5qeTqu
XxOu/hbd0XlN2YcLztbIAKjRkWSGFZSIUyjzX0l9FIC8q2r2Mxu2tLFtYJPjOxuV
g+P/M7n8S3+qNdJxzlu39rjd0vx8tGP1luFZA7rQDtWzPh4pNSOZR9tHg4P0lH28
yIYX0FoA5ezs4vsHCLpE1aKyaCB3iq3z8nneiY1EwLEeq1fNqB+9HRJlL7Goz27c
Mz6x70wtKtBBuR5VKJp1JmshuvxqeI/NMzBsbGbizDze2lIAEiqMPKaiAl+jyFPM
S1dQOnTLMVVGekHQADTbH82Z9G5KG3GTS6Uh3oKPi3dmMFn8lFuvZwcpWJ84MwNN
wy0xK9HDDCHkQU7czPJ0vZDogvrlGXuxl77nTPXF3a9RraaHdc/0kv16FkWb1tNi
WomWyeZvsxyyCCTlj9z5FhQKDdYAcGURVXTa7XzYoVHFNqq+6zgaKJqGK+pO0US0
r5iKydoDMJaAaPoQRnZ5VCMhAS8To9TfRLQ5uLsT7trpWWV3iacp5ZsW90QxMaV8
aYCqob44Qn8eQzZQGezldWtUZsrrRG2G06Ts0RiodICgCECZDuN5hT2rw2rbrqrK
M4GMpSfEOIXZkUKIcFmd08RW8/LKf5hBQAtc34lI9Cy8YD5hysMmXiwigt69/1LK
rO4U8SHDVCiFttQGE4tlPno9dpFlqPFW/UKeA9OwmUVkCTLDnukLuZe8VhSFg7m2
XIdYno7lpbLW0PSKgJd8uZhfSwT2mJPPnvk8UvfqDADVApd+oIcsxPkcD/iSsKiL
GisQE3UCvYaI0olESOnKyXrKMqBGcb/WDBoJRyWiYTe5CRWNhBN5W1T1lc8xL6Xm
tMjPI8UO0lRrD26Ch/5DnFLRcD80zQ6PiMxIJ0Tia8nKafqCl6LaYVAI9AmVGW5V
QzbzmGofmNuMLs3Hm284Y5hDXYiAmLDQ3nvrVoSi47nz/iljFBtFPtD2PgAakCvz
Y5QcvJAECEDCqLdQ6INg6rZGjx+FAhoyryafCLoKxf8jsRcSlKFSLozMcfsOATVU
AyebsrKsdBsN/Mu+3d0SRVIMExCxEB8JkLnqbmSaOTULKc/kgtjYLV/GYpd6Thi2
QMqYsh+sIuS/D9K4RxT5NLO4bHupN4u0QMyFdiwN0IdSNN4GnyjF6kIgGRQDovgu
22CjNhSuaCIge1O3O3UeQ8rt4RHFJD6x/q+iiC4tHEIVti1qg68ew2a/dIoBM1xw
7J2pZfdamrQSmDkOamceoH7aADRF5elg/CzEPahNispJ5clrq2CTmPC1ffT8kOia
LkaImKgfkG2ssBxC8cYPHTQbBRKR5cMZtusJ+nCrDqWV47zo/vyF5ojEw58tDBY1
BGYrzIpFtuQdtRQtSW0cl6lRY7JVp9r8RmlmgJ3Of/gehKz1qQUIGSq7gaZP/8Ni
5satNC5ynUjOkh60Ql7TTITfUHHfhyhkwH8AFPE7Nz1VsSsgeXFr9MKD1APXp/LI
vMbfbzerEPdGGe/mn9JqZd/KrvgJlOIjeigzFfCzYN+5w07NFNAJ6QKQxLphI6ib
GkeZXQhHrml0y0w5WccRT1iqAdw/7p8u7NuKzPZaX9BbwPurAVDXqUjepqBYVyFR
3kPq4mNFt4XwVSfjZA9v5c93wi9978YFdOnH9s2YKiSmPXmBvFeZFyXsUVF5dCLp
5F+E4pR+9tZ+iq3XpG+WRxTCGfKpLwudWXCDc9GzhTgKPMcka0lULpDgswv763ZZ
A/jye7EJ/uZkcUCYfxmgJKuOCqh54pKwVgv+7T1rGpmXzSZRBzXZ81d+mU/ZWtJn
icqDKaeEZPlH3VA+dh1KwF1zm4yS5RDNx5yhzzjx8Bzm5Q9ybLUtw8rQJ6IhzjQw
7uH0Omfe1KwK+le+GL8uRG6i4VNhkFy/C7GY2ly5OyEup/POf0GFfOI9ggmBfyCR
zj6BqvEHQCcE+/P04LofQU5kzq7YdFF8N+XL5/EqzVkhHVTMkuEDikweUVE8gOI+
brzaZPQ06EBESBO4FEJaFBYxdgS8FBv2hB0z3GpTrs+tGTXj+R6lqiKV6bbxHdNy
G3yVGPEUdKk+J/kOGq9uzJKy1RezwUC+J9/3A38+wYoakmep4WgiA7XdPGy+w2rD
y7jW9VIzT1gmi4DW+f3VPW2B40jxdvNzofBe3gJ2DZSraOqrammkyaU2x4fRRHYq
/Hnt48moH3/aIpnOuNijJ7VQDOJZXb8pDxvq0fn7fvxtvNH7hhQo4ZV85Wi0VeU1
xsUvmzmcDaZtanLG/FSUT3TxeXCFurnFCkUbCVQjgsHYqZqgW9boqKQBGFjFeKbe
6Y6gzQ3PLaQYfYZqjsCm93sekDy+d+4H2Dz2/BYsP1vHZv+7N0rc5q0FplTdDkg+
lxPM9gEUmZEPpC1CCkeNXjmS/U07Q+efaxhdCdXlDFHhKjkzZuj3CQTQaaauSmxO
eCLcNQqGXtjQhV+IcrbMH+8cbwCJePVdm/F9Qkauf0SqbQHhLDCU9bfnDDHvXkq2
/HKnxoJXFxbxw6tUZy5tpyjCQodJGnSZ4Fz/HdoD+Qv0HG9nFhTdtFUYo/5FVNK5
uBZH48FUSTEFTTVBS3Xg/dSnmH13p5p/HNDfTE95j6OO+fHLmy9uax8sIR9fUCJL
gTNzzzUp8aHx9+ljc2sRI+/V8ydq7cACREP/qESY+zvC+7u24rrTPQDm35WqFNxn
OodvEe/qY54fPsVh2fKuMiomRERbu4ZhBn/WUwYd37o70O7VicCa7w4uKZXWDd6q
7Rzg8tV/dXVNca2+MVwt1sEj19WCQYlT/x/EHPbKtoHorZjwu33xBxYHa7gxMjcY
CWeIYDEpTacUTbpZK50dLVUwRO6xOTBoieD48Hvaezcn2EIq7A9R5L758wrLV1Ra
73y9xCsowJcouTui0vJ2ZvOoc0qebBAscUAJETCAjez1nCsThi8BCJBnoIR8aw8y
qtR54o1wsmFJ2tnsWqoK0HMUc/7OSLhoaB25XlKMzT0JIOhvJn2N2xzdaY7PirLB
0AG+9bTUDI4zSy/TxegW/LBVsvt/sU3CAt6wXXvQeZ2ZgqNJzc3rnsZIO+rWOAA4
fxQqrHJfDpEIpG9oJz3Al+aQswA36qtiUdLR6VdOo9nRQeHCttTca2BYiGRGoGNB
peEQ+H9BFTsIM0dwzkb2X/kEyanpgro4c/C6mDMjAob+rZnrGr1ljzo1wSDH+Kp/
NvROP9gFgWYsOprPLbsPp8wlnNNqLQU61sOfyDQjH/Ikt92RGzZPrkhLXgAwLgUM
J+bcupoy4VfhYrbQT3beK+Yd/zlVG6eT+kTpOfHRgQhyxhJjoLdHqXl9N2hdb9Ji
e00kZkTbqBSJGPRW+UO5Rd/u95ngIbzy6Kh4B029UTDdpe1rjEnGqO2vjgC7Xpjh
EVc0IqXPOc6/o6FFvbjj0mzvnWS5NtOcPcwW0Q08o11Xm4dveCnzud22IdiURdXu
i9Nl7oZEdV5S3x/RndLaqsOWYdjGYflu5eb81QPsYlkzZ/z+j+uv+alovP0I52UU
w2+Dj97zT+BvI/4CAZV1kFo6y14zH/FNmRj07fk/MRJ6rBTNAqYZpnDCOZG+7ocl
H+Y3EjauHQTtWDByCHVRuCbvfPyaqLbuMnNE1l83XiG/OFT28UMJ7gUL7i65PBZ4
nBUPe2C7UpeQkC/wwfkykpN0CBJyDRIVEVRxhegCfKGDmxtpE9JXEHvh+t8nBSKY
NL1Zjg8gMRHMxZpJpq1Z1kTbCVB+vrDEpa4sXoG7SlXfR7YleFFGwOW5Ugpdse36
YrGXlARjqiX9MDvg4ohrwjXZfnUMyFNNxx7hUMfclDSHZLOyeT+mHVNfDgswGmLd
YO6krCF+OTp4/3MChm+3hPSgnZgCsBZ6LKShmIEmVFp9x67dfhfiA2daaBlGQ/dV
TltrbnK41EdSLeVz5cYftgamuGvuva65raOWCR3E8korRa2ZbxZgGixKrnj05PEy
Eobo1HnQn5CSlbomL7et6HMpWEd+uroSKn1dV23fRoUhUcca9hDzdmLmXi0exqMh
Ba0kXSZTe6s0tk9+MQ8b21kle17o/KCOAGIetVPnHKI1CF1VhWVgV7XOG7Uimucy
8KA/KBwrIJmktqyULZVxrHDpIdNtAVae/nsC9gABITwoMetqHVn/hLkM+QoEySyQ
p4RqnT3rz0OUmhw7DfE99gG6TBqJ9dSORbnhSxjPxz10GKZtV5IoapWd4D7f7k5A
NwPYNGbOCHCBXLXj85SQRe7M0BKcy+YESPYNezW/RbIwp9wG4nUHTkode0T9gSLr
QVlhzsZH22Md9lETaGi0ZlLIirmNVY8CaqsVPVDMogzwzSUTbgl1NO6CwaYkUccW
E14K3UvkyyXJByQk0dkjmfzzlTxdogMtN3ZGYXlu2/eqGtD1DfapU0lDyU8Hkivn
LaZOuRi/1ftQRotaxENx+sGeZ1JHBJsnj1VUFr2zopL3mjNhN2mGyhyr/vkqKlzM
CXFuWygqGCZ97as8AKFBVShwR+qMvs9U65NdRb30TphkwqFbqpoS688AMjcw7v3g
DkktWl9nGC3pfSeqgddv2neWW+0c58IQpmT790FdTQd1APSw6x0PXz1njdw2uEQ8
okJVuLAwf3lzTBVu2d3Xry9eGinJRNnJwNDAMqv0O8B0YcVJAS8Rw0B/L1jNmx0b
gvPhiJ80Cdtnc3AY9vtz3DRY8zbRD2FZEM/uQv3KuZ+NRYkl5EeMs9JxpUKUj1VI
pJY6wUwPTVPdyinBBsdy966wZWQt/xKUO5ftd2yvUDRAeNvDAMlNC16ePt8zPgHR
jwLro1lDaeXJzk3JWn7+PUZ2g/8ynQCj5b3AyRN8CVYGULAZNELO47qsES1/5gRM
MTMR/6Tf7w8kKeYtzKqptNPBC/p+CuWxwQDD6iu8x5UZJjC3rYnj8RAX50WkjOeg
zUw/KcvQ5jb6bXQmxGOiH3QAgWgNSCUnxP1vYyl60w/feMKaWvgZU5YdwDsez74E
Uvj92eusF4W8N+BiITz5QwXdGa03WO9sRU2Lgw6Hg4o4Tdpv2i33AGEmKvWFSL+A
Ez8KYIKnMZoVZvbksF9PPccdKbhYegskoYY/YaJtWOu7XNGj59Nx/mDh/4hUMvXf
zB0xqdN0VClOReB8G1IA42B7wTZvFrk6rPW0WcDQDNyjrMYgbpnpfkMzWsrtmFE5
GOeebJNMQhGGeXyKDrNZw+At9LBYFtPaKygPfVOFJv3FPYPlsa7Ym3vVNy5ykqtK
coFd7P9eepF88+ooK7KELXwKFXtiiFXoR8zDD18Lij1XVyfJ4o8EDvUdoIedY5Tp
2HYyQUhz0mGfCj9sJrxIjaZz0eR1ljr9Z140GXMnH+flyiK7WBoTkzy3E2m5D50u
ZwsViOdfPj8WzWtfuitmjK9LmHIwsrYG83JfRbewekDjzrm2TrnCr9dQ18wG91Yk
btrCy1Ww5/Tw4uVJi9W5iuic11vz50pxIB8y3APATaL40stocJkW9/KIQTzGhOET
zf/ehZf03c5VRQ+1D8g0oF4iOvZ8obhRIYf0Ftc3BQ/I6mizZMg3wDa4XgOjoksV
qd7D6dLyAfLAsWy7UJ4gILbdmn6jwWvzUZkRSXaIGLe7zneY34IC/i8mEnyQR0k4
h6ucTF5+Uw48IE8qtrA9jiZXQp5sJzhCfPGn8GDgxyxuQtUpGVNaXgTAfodCIngY
ftAqqmX3X9RVKz+yi03ZShToPBz1RopafxeWQUGL1MoakSLeLmx5Zi7JRjCorVI0
j3tbo/Vtxs3RmXS2acJ88WEWzWTHP9kUZzcZ6f28GJGKzLoYXL7Qh6Y3z2WWT7uq
woo+EiIbDsgF/NOqG+twVwD2TXXuAHPhurAgQOd5T7OFcqA2Bpqbpe2Z/wlXRikL
tW1L9Yto1Cecy13H2qqpLr97yJZkYT3JSmOmkanMDaTlHtDeY3dZM14aG+1LDhWC
Kc1UwDAb93+a+QoOfs63ZY/gBTpWVGClwe2O865Ct0I6neX496Z1EjYlM+wW5g65
VosCnBQuo/u540uJT55jpOrs1pDgxzu49qwZFsXO23sB9w4IOtulnZvVfgSw4ITQ
PjIBhfonkFuqOF7gFm75TH93SHCtru+UcLHZBtsJGEf7tkKb1GdlK/Tu+zw3wmMG
J5CCkTXVjLORAw/F8HD2pQaeH7mtp2yMytszYG0g/0890U8DpPlBcdrjVXJRIQhg
E5RrejRx6exKdfYm5padpHT2vBo0gqSmnre0VMCcZHftR6x6rOqXmj/HRqe7mNOf
wibrBfrwJq2Ef0QUGDUmMBzRpbU9yzpzOsLMuATfI8UDiXCI7X70MXmMzYgHLOkk
1CPzg9dn8xA0pC/mL8erx4jWMz9PVYkItMe7UQAKqoMEJrmTV+WtGNsMkNV5cPzN
RoZQ/S6Bryz/c4z1+jfcbikhysg7jROwJ1DOcdNBku8E64kYKetXHpDgTDb2HMQX
lUZz9N4AFMHrUocqfefM/av5I8zZ7dTZFaFNRlxqiJROEr/G3jM89M6PwajQvMvR
X5bNJoR2k7MyyZucAcVWI5p06xKDDZOSi8xF4oVmJFeE9und9Fyjm1LCPkLT7Ttw
zzcgrE0lVXHTT3jqA+XqnfUITFMFAEYWLdwOoRH69RI2Hqs2TCXCahGjFs8dS7vm
XmGdaKQN3WQPrS+4QHip6Xee5EcV3pnQiwQnTfAvpbKMhoBSKZD3KYSr5JQ3EUDO
i3suQLGWl3Rvr1xLa+g40YgSwm2ZWa6Vcf1j7SFGA8MwjbXdW+uYk0/x3Yjpt6K9
2JL0VpQSNYtsXQt1XFRiRfaA0dmQ8ngoOrctz6klKtPYq6bT6b/BbX7LHgLmp9GA
wdPlnjxaz1pglQNat9BVdVqyYnl+VEJDDF/rUrbpT+8+PECzyj03iUjO24iwoqdl
bt7Yv6GC231jREbbqgJnDtqsATCT8xaS2SDvB64ZJsyJLArF+eiYm4pbMXPuy5z2
gwnRyAZz9GgDA4uBtdySw8YkLHwzDF5xt2mzylh5Tp+GGSKDNsCT47UkG0Kj+PL/
hyrDrJiJSItRxJK5LJrtHUemMMRI+n1Bmy+ArZNiq+L6ZvGtL6B3h3HS7PGV6f1A
fcjAEAhLHzeRF0g9kfWj+kOq7S0uNNr6J3t9RwouHYeB1f2kq3e7vwWRShwy+epg
XhDLdMsKgcrTXpm7RrexOlHO6YfVesTsoAorfQxfiLJ+7DG9JeFfMw7bG8o5k5yx
P68jCPm2FwAnYQY7CJ3bvB4YCKhgv/R3LKwnh3rHkInzTOuJ8MNnSUUJweFX0CYa
9VhkVuLqorQN2dYDeuDt/I2+uBZOMbrC/X9rhwQ5sKPuwPCzP16uFTrDgsNX1zB/
B8n2Z5XPUa77Xa9Zkl+6GqvBrvHayFhZbDnLIvPZGuhxO9JeJp4cgPhHmk96KB7R
s20EQyVpyitlv9xzSbUrh5SNFi/bLCeEPQNfh7hwdhxeb4UarVmXL27Dcu4trAGf
9tckrow22E+PLTXUzrvxSByY90B/LT0HYT7Cqrw1OwhVHOenFB/VrIutbOyylIy7
1RfWiAw5AzW7P4y2aG9U54kn0CTJVLj25CCtuvO333woDx7Q1RhIngI4EDMR+psg
mNLst2bQ8ARLpN2WilxkFLT+X/hw2JjmAfwHYWm0q7OjCopkNivUi1IN5+Tk2wdS
piC63y8Bcdo0xItf61T2d0VXBY1Dvk1GgGXIle58NEDdhvnoUKVDTDdM7ZzdVpbQ
ZMjpfUmF5fhNEV0spgA/IbjMUtZmHfR4i80VsBI1evi/AUCcFCGGbNTw9kNsQFa1
E/kHPl7LThLYlAOlc4TCJ1WkSFzWAaBddSHfxjhPdWEyKG0Gbs3yV9xpQNP6nGJ7
qGo1dsxU8NSdWE/LpnkHlNQwjkvZU7ZrpR1EdxkvHuokkEyQb0IdyKWN1hbigb9U
1w9p7zaVIJlTQ5pHxwwTXuJnhj67J+jc7TScMpJsrO5WUcRjOwA8sv54T2lR3nF2
rIe3uKD2bvJvs947iFBqS+6c5wS+EcC6e2/m7Bk5gXvSEGMYq6+1WnaXVL3gC9DD
riLq7R6e2isf61zGf8L5bG0swv9baUiIzMF9OpeaGHyiwIuKi9Ip4wo5c2hfJxsj
vYS2XsjkSDIcd2+oXx9IXem7tHJKMvFYimow+WT4favW1nUbpSMwdm2cwwjO0ZgG
DQP5sO9A6ozJ6fSlY3/YHZQbnX5Xn8qBj519d5tLzojGXLjPJ2Whn0bhaXOdeRwm
xiuDSANvX/nTTi+GKskI2SvuHM8ORHumem6zU7dNKfpRa/WTaQ/xC1/taV4AlxK4
7zEu0RUfHLA0gsYfdY+q3r55203CX5uuJTWO5C2vFNowKY+6BHZJ3NAsyF5xCRwH
KBkW8aSDXXkj2sCezUiVYGa6d2B0Hr5o1GomqUnAzT3oVft3xvIGv8Pt6vNDvaYf
gui7REWnpRdNmOUvAVlACtC6hGSmOzNZ9/CLNgR1Ih7PsW0BtIl+c1eS5ojg0AXQ
FUmOiItS4Uq2zhPXCkCkUGaTO8N8oFUs4aRP7stVKx5D70S10DPtkLEMonncQ//H
K9c+NHvZ1GQ+wJbDFd+e43q7plZpLvhIErZxoFfdLL/PFSqnq+CnMgwsgOIIVj3t
9hG1EDpWAABjUdF5/gYS9ITyLmVxE4qVAUpo4U3frBaTNBv2lPrD03y0z1Hj8uWQ
rStIhztbDAiYbNCPr3ldnbq/NWQ7kKolyG/qFzzNh78votQ1hkBlbArzDuDs5azY
rWc/uCmmwoOpZqaN6zETc7ZPJkdjfQXXti680XaXrby1NNtq+gnpAM5/coKj4Y6b
4daFgKn7PZcO1MDaEL2C1RVH1MxbnvymeJrUQEQ0SsH2I9g0KrsQXhQlXZknXkSJ
7tM4YCTkY8fjlxfrUQRZ9w9kCvq9Z8mAlGsgYVuQFrZPxcO7GkbD3tlnLFVeruVK
wtZmRP/npxnd4MhrkbgN0D8/e/fSwryeDJ8DENDS+p75aurPwVdiz4eCHtsydjGM
ZVc5Nuf51phK/OJ65n3d26Gc8UGVrt6gO9asqXXehELs9lEgeEiF5DJX1r3Xdec8
sz2n0FdifWe5u7bvgxau2p2i3SZ4Dr9Xm88fwmsFuv5W1CNjEsaZODapT8/z/RNH
EUBkXhIGJ4L4WocJMqAczl5t/NWCRsZ5v8cMNjlSaKKFxXhsw/+R/9unM980FGW7
rUEVpLgZ7sGitiywuczgqam54+RcBPPJpIAxHGua12EcF+2UF3MYtX2Oxzhx1IJT
J9DVflxEcoKZ/nX8SSXANGTghIPcpa9xZ0Xpe2O0zVNLDtm/Y0X5OJMJsPxAMkt/
Fuyuc9ntxUAd2AifHnrm/Z0tEfwmgLrRUo7i/UIm3LIaqFYlMxSKZKhyJnJuRF9T
MiMU8lnysukU6t7y9oFr1UO1JZoddlVaVgFm3VPZ824BfgpHpDFoizyvw0KVIBJR
S73CHjAULAkYuiVF+hgZrORfsXTHH4q7HGaRSe6ZzJSsgWHbsa19YP3j/TR1RMKY
YfWUUNHvm2AiNqbyY0gmnkPAtq+MNV0Udm2P5AfV1K4X8c3NWX5TV0Y0HNV85Adm
f3jPQT0Lmw00LLOMGwvf7u/gdfYheESonDC0z6Ox/yHkR4kKwg/LJK4B4Oj6+tLe
uZGniOXnBZMBLdKkaKLJ9AmJ5QHCbXLpgqeuJnqy3AKsFBw8GdD5DgrjnpuiO/iL
kna9mcyCHwGJR0Lh2ZE5EPCpT14eR89ryFEkVW4uF9o1hdJD2T8axuUZ/oXdUM1w
GtLETGuPXSG1QgK68A7ed6Ie13U49jUrZ3efANUKLHTYs71PlMINaAKJgw2a3VjA
Wt84YpRPS5JtXUOrbjpz4PuM38TBxtnxWHFXXRuX4lnOIwExAgybF6Q79PplUoqu
I7z4ctc/r9e5aZzzhekMYXQ8eZkV4t5MUpzuz+xThFcgcInwDYwONPWGH+bBL93Z
5GNpw0tz/N9Iuv87zvyHkdF7wj6fM7j2jl247M4ygoTjCAvPDHS1EHm9jVLI/nrK
UJgOnyLMS5tjGcwvLJrCsY3F1LPJh2G0DGk1x+Bh13uKikx+dQvdAnhG3Uy5ExoT
aPGVVGa5xFbsc3SLNHS1vhBEZ+DxRRRnxxKmL76QYurMLNZQmp4Ug6U8+7mu/w0N
ewVsy9AJJ+ztE7suhYQHPHBaSGL4PRrLIR+R0z7W9nipXqCcDsPAhltptJibepR/
A2VLkeyuibV2CEkvaxLe3jgm5tZGdvN21PRKvmNYEbNTNW/iQhHCWwMnLTooBAqr
j7B/7cceGdN1SJRRsYn40uMPx1xu+0VJq8rP98/o0OyR3Tc6glvnFBDg2qjm7xRD
6M/3MpS0hK2alB5+A+RCNWQp7mhgTFDbpF3dGwH7we1dZI9eDTYQ2a4nDFu6OzDJ
PGrNi1BPBJiA7oqg1wuX8siZt1vlbCQ+IChHSaQyVWQm4g1yQXyu06ZFIsoxq2Tx
flt6lUcgQ4Jfnzs/5xNPBOZR+miCYaH1hYVbqo3WBANsU12gfhvaY2ov1mq+J0+1
0bSZKsUYJq4nhe49qDgxrDyX85bi9h63Q7KN+GRvbRe0dv5VVaLwW6OhE9xKTjiz
dA6o9A5MMN0EkL/bJMecVTGihjE/9bhDKcHGm/iDTdLEPk8YP+oIDKzqHr62dCOc
9d8PPz5trDMYUK++f0pFhKIToPhvkn5cPdh8eRs2YfEnY1HHrHa/Vc/0qQ3S+Qsq
6ZC7OktAtLc5LzyUugRfmb12XzEuZd+vC1FxiyWwc0iyD+2szpkBLoo0bFN1dWuS
YeeMogN4bXc6wl6Gc3A3VH0JWIuCMX1pLOqe1Z1iiX+TatJTKhYVdDC0ejFvXYQ3
CG2QEte89EWQcMYWJqmBsCWgghkuECv0uptny41Or/qMRiCEXYfI+++Wrqpa7q5w
FYDgesovf0QXSxf6LmMHBtyRoVyFBawi7LnMWEI8naITiy07e6UCAFlHMjrR47N2
ImqevMcC333pTFT3VBblJI8zhJnDAvprMdtl2BykBm+p8g8wsY4+xFeXtEym2yTI
zvgRvwOeyt89jZNYEu5IBS9Sccnqk+Lrc9T22Cu1oA/0zvZ31bItnmJCZQPapUfx
3xr7kaKdRBZswfmYp0+QotKZTvGvnFmlgQp5XEgPQ4JtLAQI7OGww+f7Or3Mg5z4
M5WezZnWkxm5Q8zJOA6OOJOW8F3RWwLtqeia+RXBnRFDlGgo0W/fXUnHwzQ4g8aP
ndPD67WJFddF2QnCkXYMTkhlMSyeG1Za833vFxHYRgVzea7sSfQ85KzJQWNsdf/X
GEUBXzCYycJ8pgx75lapJwQqq5j1eFC2YsycMO23pMxNfTlZIbPZzsJO7qAz4son
CpJn6qs9B7SeBYWOeT2IXg+AKChm0glDaFSz765OUp/Deear0RtQKrlr5+5/eoqc
mbZK7ofB9gx2Pt/M+pLZc+x8JpIgHurE2QBbMtClnzrZ/Gt0vvaLLI7yToZ+OSWq
fapWIkNgS+ocrVamG/nkxw7h5Utw7l6eQIPwdYRv1KninV1Je910XoyCo9guYkUI
dkRq9WbLl+sh7Iz6JxhLKcY7E+ihy1t4HiEO1zNkot0t3XcXm1ERxXn7m698q5mW
Y1xKob+CXUq2v+odYxi/tR/FDxciiMUX/D8NuZb/5aIqZUO4i+HrTrwKohksh8o7
GKYioKZM1lO+UqjCIdzKulvGkqdJvH9UaGKBQbF+lcXhoDX2+KxsRTYWkR4NIG1V
+5Oiq9T3Bmi40t3mYLyzyXP46TyIzpEUT+DVIDv2MyeM0UQoXkoiSe6lw1zOWEF8
nHNZGXngNQGmBODbQ5eBJJZc/6eD13C3uCJQ7YTp8AA+USXbrsUcqo0hFF2KqnqT
DUpQ1TgCft8ns/9Lhj7GlF/Tdzh6LFWh+WqGEkzU9GjzqcjFWcIf2aQciU5CBI4B
x5CHMcI3qxu7jll/4Y77SsANR/mFoXItkMOBjiXhl3vi4uKcDb7UTXgzRCvna0tN
D+kdSEMqwSeRWHCzWY65Sw3zeBaG8h+wY0PLDwDBUvbsKTw3jI5XuwHepqjaP93k
H8ySZxafoqf0Z5U8O3tuJyOVwueiBDc9yDbn1NR26mbzEU6HMJO+HrTHSIv9Tz14
zzahKrs1ui7B9czJ4XBlKBGGujsYA/UDnVX0pyTSw0oXNzUty3GUaxPfkjG33y/p
7HpfhYPAywhk8Hnlm700+01Edn2bX+lqzf8+6ScRsViP67bAY6SbQsfQgMcL+W8U
AgwJZhXATDFXGnYSVEtAZsRNVObCxjuPWQG/1lC4tGP3s+l/2zl08Aw3EkbdfoSO
r+boi8vrwpEnTwj2TB9XQ391vCyuT0IC1ZAvWvERQHB/eNY7+kFm0liQUsD6+A5X
x6DfLIj2aCU7loKX4Sc/IEP3XhepAB+bHMAOD767amxYHvNpqV+8SdxxP2H96Ax4
0qQ0SmtcHuUi5ceYfhTsaOzZqMCp9go1WNJTAmUROxD+J7S0zZqHnRMaEwyg4cCt
iIyTbaDrAxLobI4ydYaMSXRAcm28D3oXjzg58dXzaefCL262d1scLa/I0/PWHWad
7jZB7EKhd4PdF1AUVbsm9157EqkAKvZ/gLCx6MaFezdOllf4OwTqo52+mUfTrV7B
R033oULcAawdHn4NWOd/GYHfQqwBgP6cq3dD3KgsjOAfAjhCr7VlRnmDPmsT0jYN
OrXlmx6tjinxumSvlwgo6pzKKq3iJgWUDhpiwfswClLMzB56ybGkVoD+pUcO1VKF
EJYxcnkFedsZARenM53Km48Z0cQfJbcjP1BiKnSt6U5yE3DoESnfnDZ/QFrViYlj
kkBmkXLldfPYcyxd91xdJSyl7ItfjN7cmxaLsWq7/FI2/ks17IFRL9caT9YpsZRF
ov6phQHrkoIRPwDHen4VUNAky73D6eR++IHYGVZz4hcZT6ypxkuiPEhVM/GRdJBa
H6E4JRU8tVj/Pl7FMcRCe821RWv+8I1Mzl2EBUt6KAJd6gqVvSiFYcSWMVVafTkK
cVTKP17fblDxq+ft5fROJwEVvzx1yCiCKZbkv6TfkOZuaSIohPeox3Rczfq5cZnr
xg5P3+ANk0CAcPO5Xmn/IvBaeEme2RNogKWYKs4NcJ2G99XWIaLk8nsuF2mKLRkJ
uq8vr/7jST0yV1o5l0ogeyoDL7LUzcQPmhraGb3VETz6oaxLxAn8WNvK/JBAa7xF
FXz4St5XmvXuE99Mv8wIjdgVkA0FYLxwEDvo0/s8jRCFGO1ODGQC0CEZ8vI/FuE5
zNEe1MS3j/7PWJyMQLBaqJZnTHcSxc9PmgBFidu3tlMh9nCB08JhEeqsM9axO0KC
AOJthhYkO171wqy/iadxFsLL/eMZ07G9w9lpl+ZAB1+DVOPz6Y2NAEKzascxO/hl
zqxnyxqAh0aAa/c41H+KnQgW79LJ4UN4p9M88uslGkutwR77+2WRFk2PpzHiy+WD
3ub+4Z4T1hNuhoaQQmVjEyswmae50bJJ5VesAl4LLMugaJnDY3+j4MnXidLdXRS1
eA7cVbzP91QG8KABQom1aHIQdII68OcR+H6vHPxDHNUeGq+vGSb/diGUQwWQFRzR
AVWMiWvrc0hQQqzr6dye9VLup6dtNDXaO6ODc3Qsccy0Sb14YweL1p/0BSUnNPrS
/ZZA0OIzU7obE6DMBdAi+IOJ7yJ6mr6wXDDFo21D4BLGr4PNK7yNP1w1EU80dYZd
6k7ZAG3fUZ2s9lRCSjIE3x+Yvp5O/8gIzRBhrIKXsHWK+wTEmsu3mOWP7cy86jBL
+mt6Pw8KhCYO9ufK/ZuiqPrGu1xRrCG7aUHCbfiKUUhLf63cxvsOASW/Bm7xEjrG
hnh3kg8Cw6QGNKj4FWz8+QHWsqjCwP4fzNXKmepJNb6KXOu2QDFJf+V/4e6peoAy
+Hxlz7gj3/kQ5pFeY/A+TkUqCnQ8ww438p7mrfY2d9AWjCxm3ga9vUZzZhj3HHnM
LeUWWVDqalP2GKfGaoMpwQ3kK0XDkhpCVUwTqwTTHksKJwe+7SMKw7IDUniZSAuA
XKEUyeY9Cmq2D4o7febo21ZhIvYThMUUGZvWwxkSwce+nERrymVz5oko3xI5odFt
B32WZXa0PJwYpJzH3SgLob35i/rABeRq57KY6v2UVvZg57VnuT0vH+DfjnKQWpVV
jIOL1XObiscY5GGwUXgNwKYKst43FvD+STgUDMttxf+JbS3aBWRjfxNIbDv0Nhfp
F8FjW+MsltplkdkJfxnMTwEyqYptATk8XCHynm9ybADg1OYWP7ltf0M+Hi0K/bKj
XmgjdrSC4ARGUK3P962Om5BBTULq4vtOmJQY036IIO2laLt9vTab+QqH/czPT1Kf
nNT5iVrbYZXDNLwPB7grCYLjrTwWLnZkjEhdZ/5GWfeiymI1TgCmGlOfsfy1U9GL
VbeAhmyT76BxcEIB0/rDD3Nuxdip1NUwAZtUB1WbQNLprlmcfTv9+J9Lwe5vsFRv
k11QJOYuHcriY88ua7rAcOU2tP1Q8V7oTZNDg0Nyrkevz0s4j49ic3CTPIq8KZH6
JLoKLJkc0dmi2xumVV7NbVsqGK0hNbN44qzCx4lsov64L5DzQQ37LH6i0d0Oq4DX
jL1ijPUR1k8Ko7TtIRcBZJteA8nKUUwwmX/9i1CpSsqbDm+/ZAlRJ2rptGSQeHvw
6YxvBRjUrFvViEv3CrT8EdNRDaZ5WngaiAJv0bPdHxvg/fNAw8qZXM4AgFC6dSG5
V5T6zb2GiGv1mjt2pZ6JTRugUaHyGeGW52OhluHdNDvqW3bdhVPF/MEiBLbi+VCX
epfrysuiAhY/g+laQZgXi3jBqMgcNDj0wMkM5oWwMPx2ggoaoZI9CmVzPuqXn2pL
M2tC5ie0+gk4UI7z/s1k/v1SnCayWU68zSUoBOic7gq52cATp/azkOGkSJCLq0zz
l/CDlR7dYa4QZ2/PQGpxoNeyBJVCjuOQjxO+pA2RNrM5ESVW4VBfsTeapU0h7nFD
ONFhJmNyhz5U5GlI5+D80WbGEVOwS+Y+MFKTKR0a5i7gbCAbPEXh5zrOrY/PnCyj
NPaHXePrEWM2V1oNl5dfXSz0b/JkFMNXeYneut7KTStZT7mwADXmtI/AuV3AXiVq
7wnABoYeA3CdIPPJlRXD3JuYYbR+VdfmjoXxuIEIoaTXDIMrhOvyMVZ0Ba0Ymf18
4SYkiEEGmOFpLJsjo5u5R/E1F6LNTuhHtd6degW/YWUCcO2+7labLaWDzgOlrbY0
cypQ5b5sOc+WDZ4wuL6vtin3iejtmKoEHYHzVa6zZ2LTnzttUZhzo9XUNoLYaS1b
77+wzz0lCHZSNRNWhfaZN5yvtm6Tyq1r3pgUTUXBBRGWBufNYcLut32Ef71wayZA
GYiTWvvxLK6skIsF9Ixm6O3Bdsk+ozoQ6OFkBkaUYF6ZpLbcW50VRWRfkM373DoZ
kpxp8DejS9TXAY+FxM4+Mw3qwOdMvqKlKP9/aWV6TA3VHZSgFLrgPVn4f7vZfK4i
5+1L3e9Z2ZL8PyvMJvGeLi0LiMRmJYHAOSbuUosGChKAhj/7+MV69GJcjx8s8sBR
82REE4M0bUtCPTxPcg/VLtNXQc2kKGAIlNNAX7oxrc9Fd+OaD7KsJwHJiHMJ6WrM
svsAzm/WyIkPmC7ZYFtDSZPhRMR+KT188eNZLvhecalO73qibEteRGGwPf/gqfr9
x6VFXTVRnY2/4Kb901pxMriPaLr2+gsP8kUMuySLwiEdM1wTjwry0xwuKJq4HaJc
EcDZ+qIWDMz4efzAPKEnhKQwPo6v1Vd+mW/zm7tY6IAn2uNkT7VwE7yWYLgAzMWz
LTBWJQIHlOvw4xW9cd7NnhUr98nDF6Tcaf3HfzAvsGeyXYEribv8jKjvQfuZaKNt
cI+hkP2tqFViAeSY9Vk6klkqf24R7oko88L0qKOImDtQyFAQbw4mVj63wfjmHDLL
BAN2rXXIEusBieanUx7mhccaK70pBMKUJ2Y0ZzTevol6eZwmncTXbGUy+prEx+1b
MOuWVtQMJ6c4PMnLVaBlrIA3sW5z5GcAeC/TCd0pAXYsWHj73JwXUstih0dBDrNb
z6FWgpMBr0EE1ch2QItJm2qAiKhZ5w1TlSQ77+/oN8/C7ghCQxODjcujKEjeGBym
yMO5BgxsVKcgEPL4fXdfx2Ppyr/I2YXrN+2BZRcnw6fYWLgRO7rquqRqe4gZw1/J
Ktn48FOS/1aydkA8KYjciAhcWiP2YvQBmYasQ0eopMfBwfT7sPUTz8tjy3bmAz+o
nMYtto9um/L/7RbtQal5kLKFO1OrSVgAjBLZUmxk6bd+atDsjiljBpaRjz7jdQ2h
a6RPkQYpy+pZpnp+oaQVkZa6F8qPp8vMCGGXLB3EJXOjZSQXCxu0VC2zt9JLoHgM
PwykoVk6gkItIaFjR5YZNya4WBnCIXrHQuCROe3izSbueHH3YYDbeCtV7CG90TSM
gFlgkTVpF0/sfMMNWTf/6oOzvNFAiEmw3OKj2pHEpAheRUBvWEP4S4OYqYVwMetr
Cj/0dPKMni3pmupiLNDscDbtFKpETL1AOy08y3FO5p/wmsFitVAKMfmFootR3Eya
sUh9oFx+ryD6h+ZQ2MPbERdcwygamwGO1+gCK5mfV3/nOUSUgTngNeTfZTwYYHnx
9tBLaXkhoSQtP/dbGEhqrC0zu4ssohs3Hf1jPPze2de0zVprlJCsbg5CKM/ys50k
HWt5dLaUpmI9CKbgbvdUpsgD5cFCannmxd2XX0/zrl4rDGybxpBKneSS100GOAx1
XQwdLVyT4GeKbJCpkey2x7dfBlgMc4JUY0Y95GYzhDhneo/U6d2EX94zNSZvG9Tf
iwp77W8zk/tfqF1t8nB6RgaKeXiCoLnMppp5WPKtYuCtaryx5cezBJBHntvdnaFh
t6VP/Qz3GwuPDBc7dvoXCtt2WWs+ZTkigAFzLiKpqDPNk7JWu8blb8cMlQRTVKK4
Z+lH0UKXj003MhkPUhRWhjHD5LOYNhjWcEKbwqLCJtOSJygU/o+TdXjHcg+zH7Dq
s0bKWhUFRqJY9biNoPCUtmFNOahCZZshiHlJCrAH1+QNILBmZ/4m0kPfsD590rBB
mbG/Fahc4tqznR/LhHK1qjNxjqHWkGcpr1taoqJdf7tYKCseNgNNb1fcMm4clF4c
0hd+GoX25PrzUhkbYM8mRqreae7CoGPUv0Yynn5dBWRg6O/yVlCTrVRU0lsKsEZG
FnTV7AriqFS+DYE4GRKFdJhAV3BFI6dWJF0y9+stDmsav+x2ay6BqsxsqeNzUC9S
gz6C0vdPBZRC4Iab1q059OcsRa6aOw6Zjoym1jKLFiY7mdGgp+blIDqa/Qaaup7c
EHUr+w6JBnmd315l1r5s1ANT/nwJORTxOa0QTJ3d6LGp2socgh6YDlCmqJZS2kDM
MVm/vgmJdFbQ0wcfYRUt2+nSnIDv4rAYDiLd3bf4Gcq4Sbj6vTqSavrQLREWlxCo
NgVzP5jf11LCI3EpncddAZWlBh6rq8QbY8Ri4EkOTbocdi6w74McNEhorK1yon4E
LjtGX06CfMBjvazaro/fnuO0t8nTJpxozeW7mVE9eacyEQQDkq2YlZ71vZCXQj4H
pWt8H2zBhDbDrtB4dk0/+zfsRo+qeypa5w9zW51OV+vLnGrcvseSn71fP7ISnQtl
vhYq81L8Om+1wblh6Zww2pONFK4Iqn83ZRgXURJSuGTV+zxr4pQ2ij3YgWXcGH30
ncriCI8tWcKj2YcLnQUHv4gkYesowzXcSui+gKidKANfwU09xWv9ULnY9PBpMbVX
0HrzVv+5A9f0oKypcX8gz8GYQ6fwHrsUo9bGpBwAlazq0jTE7dl7e+Wz9lWu4t2Q
9vM2rMtx6L8Hi+zcg+fqdg4RRyrhBk9PuO8+a0HlerboBMZOd0QMgc1o2IlLQH+w
XwLV1Tdt7d4qvbWmu6UVqboATG06aFI7KlL8eA0Co14eWjlcSQTqW0FXUS5/nilG
V1ApLS4nbgt1FfieQFOx/eIDITQiI2mcvVm0jRpfpW2jUceTMhHxWIoIyFb6vp/j
bh/bhE1c42zLyWpuJMVbk4Z2IYqb00hEhDgQKSNmOIrTxc+T3OSfqa+x4oeNrnh/
8ezy2T1BL+JYvX0+xODLgb6BnfNkBSbgxxagodvhz9M/wt1HKBHhYHa2cJoyZjYs
qhVhpbV/zta417u/rU4YP05Nr+DSBz8CX4HQdz2Ax+tE0zcWaRcmGi/1EBze6MT/
eBwdY7pfpC/6oNZOUMNonVq0jlqS16a7KIB1vGT3SvINO7hr5dCzyFJrchDqcIGx
iFHIXgkZKSCvzDl3CCKF5aE1wbIKKDlk9pK4fp9g+1hqRBe1VKZneLodFZO09L9l
kyw13XgNdDyTnlA3CTYc94yHTSBhEnYKsYSPZDXL87l8QrLu6Rk6MSmkpU4XCiCY
tIQLsVMB18F4rnXEZjeCLJW7Fz6cAfoMRL5lFIUmPwBgwHNYFJWfvKbZzQksceoE
5pKtxGT9fSBqtN5NCkYR0FIwF4EYu87TlDE1ss6kQZx7t1Fo81jczbRgQ5MhMaIz
z9wcQScO3BdqUAoU8uhe6mcDEni+dgOsTFAOoLFYHyyaXCNLsYLdHhv1JhHl3emv
3ti4lMggurZmNohR8s7yrV+vedgb8uACYRmsWttm6PMxudYPqmKHUNC9r4pQyDEY
A16/uJAor6ii3NMpvtr9CvkevBaiiWUU4OlCTdaX8bzuCBe51QhzDPe9ZQYBKfGr
QM2RfpXH2k/ABlpCBqMvIfRFOyxJKMMO+1o6MvE0QJ6BBcyC9efDwoCidOdW10rP
85XdK2u/zNedLD+xw5FlGjiN7hUAWY1GVl26V3RlbCGlPq+dUf6I6Le8lDT2cNnO
26wYH1IWyMIJKkF95uyaFHQOvGGjUn67UpRTEsMQH9No1zOOlG3zgDlT/ADtgK66
4FKyxJDBCNhjdCy5To/64mLV1BtiMmZDq1tMN8+Vfr6Z2fm9fYJJ9Aj3zMYBvErY
i/2xC6hkO0OU3abgWrHXnD/HfMCnMGExTMuawXiznQSyy+UDBT4nEy/levB69p8x
M54rQOMSJxtvg+f1eAwTJatbOSjo3MjxgH6LpJs6TM2Iu/N4uYBclYTd/qhbupfY
JxND2ZbdSdLS+H6lfjXsQ+pkMcui9LxRM5HXURWZ6ZenKta2FPq2piL620IxLSu+
G8mfgGw0PqYz3dz6MU0ayWUQf1OnuHWlhhf7lVq7uHRvQcZQ+97v9F9hgxTL/UWd
nDSpNZkPmO/9/ivK+1NlvqsycXW9lUADQ+jcEjPWwhfR3W9wtVqFiIykrgikhQrZ
U4QABBzxbHMt/HLlJN9QPNbmkyI0K3iaQOHkTj3em9R6QraoZwUaua8kBC0+OjTM
IaGKwnSLndyASj5Ps1ayaNF+CiwaAdMMIyskW7FgRtj0UaQujolayqkzummjGxo/
Rvzj0OTwNny2TvLSVXtYmNTVm1v7Of+Y7s9Kdfjs+oKGDNTF17hhp76WnKiHK/x+
/Fhik6A7WSwsyHXKllwMYMJmEJLkwTojeYx1D3X/uL/ZW1juL56oodUi10jHz4Tz
Dew3NjosdQF79/GfvozQQdVre1BZDMB3GgWzkUwwYdkve5YUSQ6dKdUUXuXyWQLK
DE+ZGr09uhcymjil+m8HCemj6gJoL98vVKHLPMWJDNBKNOsIhYPwEyVr4Kt+bR58
CEfrdQ1XYbTqI9LNDMWkalVapq9Ii6RflpuoUcCy4QeBMr6z1Dvlksp/uRoQqiO2
Kc4To9pkKoT0moqD+nWpgrMyLfbkzjV3zzF2DQrkcclytAFsgnhkj3gsxw0m7TU1
tZ+6p/YVmHCxw/vjf9JPzphlW6VUHI2q8bCD+e75D5sE7oT6nIK8lbf1YUFGOPsD
ETba9mAJOcfuV1BVY9rbRrK5dgKNfEIxMQQwzwAgYaELEXfce+/5iMNQbysrMyMw
mx5dSlHGO9CrtcFS2JZF4+Y7D/k/hIyL1LLsMg1sSWWVUVw4S48F7GnwTHwO+L2i
SJ9f9ox3bshEuxZfxUYFMHO29UiL4aA5Oa/ESnujMKfi2C6t7TA7PXaGXeXSuJWV
IPc/JoEVD4WqcgJVPZEf1p80zoM8X0n1IP0pfXfHYLLLHgWZdTlyKlN1JxKgXUaF
c68HdGMPMs3ZWxtoTJbKzUuUJusMveSwLfo5FRMw81F2WUN0fdmAL77IIlsIMY9h
3Toa1KgnkoNSB3SGtzqFjhYkNLpNxfYFD7f+jVvYwB+VsDtOrocR9YJTNbyXKFr+
HLI410IgvTqPJpsR8Ctzek1S+9nZrmVS/YBlqWLNGFR/P7MzBOIcEpMGl22o7otX
NxJDO2Aowq5DK93Zlk1EaN9NVBZF6PlrkqGaxpD7QHDnvTfJO7dqSb0Y9gb19p4K
SCLcbuINuV8fdcc/+VwQJ2XZWbSVc+5dEPMRWPFLicc5Z76RvEWCvtVoMZe4GurS
KVYMaEU+RI9IL89KZBZ/ifioUbWI/jWixMJ1N6xmi+rR4KoWoQYFnrYAbdTlDtQ/
791NxiTochvpIgC131fZ5ZdR1R8uK2OGKROhbYuapcuL4rRCuyPjxp1BRQfVanDV
oaD8Fq8PAzSHgNB1jhCshH0HF2g1uclBCgHxTzddhK0bKMr3AjczyjeIWGBl+S/Z
S3nWE9FgPnp+sQveuRYpG083v56dxfdrOkM3OXPgcOuGVxzfvjY5i+28RZG2EL6Y
JkOlgqUS2kXVMfWlQDRyrsKMURUCIUHLSSAQkobGH1yzmoWeFPbYB0wKV3rTO46V
i3/SUnz8kJ7/OGoD56h6uoCem/0UAFURdTUHgSYTYEl5uge34CvtzOg0QEEBP2a4
vimyQkUTXfgaYLjCRSyxYwiRkXOKhbKBIbSVYfJw3F+pf7bJj2H0tqurcNzSk9FG
gnGMLVgoYi/YYN8ZtcxqBYbXqTYT2MDHqR6UoLTgskOgCKOYemkn5VuKyurK0aPO
RpPHY2Qqpcl2rdgTrjAaCTTndHmK0bPdNCna8MmFIxtmH0pf3rQt8vYPNflAysZP
ru+S9IhNqor64iKgUZQjxifZ54mY6/R+bFFNrS9hBQNmj9O/cQIjYdJPVc2pdoz0
zuofqmJkdrhMb6qZDv85hkIoCXvUMqlbY2ILL92fwEha/femUjJDEfh/Y5taAprG
U7BdO+CWI62c73hSTjez5cdEgCPO/U9T6InzLi+Foc4LAbhw39DCaamQpuKrrpLr
bFudHTGymd+8MKDDMgPfH3DS/OnBQi5xyOX8A1qNbHwcq7q8JVw7xtciUmdvBnCI
EjscwiREYm1pZBJBz8+XgRy49642/Zp+DZXHilIpcuKdMOYiMRtBj1sELz/r6RDT
ffa0ZwNjcfipi00cmI7nn7sp2BY++C/EOPBfxtTxH56/YOUt3Y2yOzKQk/E2uSFc
+T+eKCGvrVbeuCasq2Wr1JF8cC42bqu4/xIzd6KRVH/hae18aKMIjlDwH8ZrRNcp
NAAfQ8lfxyBL0xIzljj7ilwjcVmibUMpAFuzg2NfUgqVezuTTwb2gE1t8E7UZJ0M
5qm3XdLe5R59WRcisln+SShzp7dociAbfG/DlwzSKlzDgnwpuei7P+3lfTHwa/pN
NXozKthswyeBaS55S5QlWgmaRnqWvdOwkX9aZ86vSJGD6u0t5IWj4xGryj+WSeHf
yui67eDqXiBFXooDhBqk1K49Vk2TmmLHFN1eFeEprPi3j0ZO8qVm9gT9ezekVAwJ
Rey07c6MC6jOmGICoL8SNZKfgBq+JTDLPrViUdxijo2cM3a3W/MeJllbipX9wx/n
Wtr2xUGITTTEOE4P02bmH0ceosMY/q0w3usxu1TeHEJlW/6xE5id4XaAbiEbYdVj
aBjDofumuvOZic4aGL0pWxnagUyPJwDZix3K0hSx95bnyPWtZ5dcrycyblzbCxLv
Vv72POk77gNfPYKUJAHmZWkucUg28ANE9FV3S7ACXR8egfRyHo0eZhPp10ggQazE
35t7tmqJRNzApKmbFJMbgT6KeSRYcnnQGAvxyJb6elpFrYHVqghPFbvbhaH+6n7x
lKT2lpt23FTQHzmwkvfWPbMcbXwl6prADJuTe8C4SUoflzw1IMxMNNw/tU3IAR3D
WMDid+klHxP8Y0CBr0DnKlGkDF7rT0Qd5lpm5rM/CBBBq2w+B4UQ3gtjUmzZQtGQ
ccxVCPQOo/J3aA+Fhcj1eCuVXDg7Uzq9hKnwMBJByCQSFa1P4Ze+Xot7cH4IGJKd
JBtzZpiHhfqY+ZjroM8E+RKjKcOF0quu5GhlH5nox20R038TSDGIgXAoBxPdplMH
qGyoT2GQ/zsVC+Ff4F0l4ZZQ/JkUnB2FNvNEKNooWhk/cXlEzHkV/3HQCIIHq8PZ
1zk/rMkpJXRhvn/N414QZ05i7INj7gCUgltZIwpwElpMPVGGdj3Pi8lBCWyfZ/SU
gYmrq2C90Zuln/d2fVmzha6WWYbrqQr04jdoPJrrun9g34cdUt7uQRUYUiJisLDV
ket1FeCFZiIza9Q+xtRl1TcPXXQA925yI1QZUPDL2Wse+HD8DyRQW+h+lx215aDd
VJgdGc3g9z/NL7PEOl33tEfG2Ziii9A4UNAA71bxYHXvdC5qu+T5YymByPbKffvZ
szt08JPB40L9vpdRiVV9sBOtbCGC4ghPmU0holk5q+BtIDSrCqqNrtOyDVpm3ipS
yfUG+MN9f+W01t+1I5vm5q9k7k11fb/tYW0bKn13bZqexQjkx6aPxoqB09sFL2Jq
a1DDr4AdtXJYsyiE3YbgPE9Si3Mf8qsU/F2CjGOGZ9PkhT8yFkrjYgj1NfpBFlh8
5dwzj3d8MgIfIlzJzaGqFZVT097NpLXhANkf+RgIARzwHPESBeVvrz8JUBrpnJci
guSITRD5beu0PO4QQlJEkAj18FJXAXaVEP4m7eHbR1g711eTR7Sx5568ywVZUivX
AVUeQUp8Zfzvni1uKdL3ppy3aqaRuXjhrvxKUX+Jm5ftNnu6XjbWMbIFBIBgjQ0H
90h3vJF/HsufuVytQZJuinuMgWesmi/41GzoP0gJggcVVlV4nJ4FO3PeMGiZyYTE
ZVX0lW4q83Ug/ffh65hIv41iq851HzeJxfFKScts4q852UsiFngV54sWOm8upQV2
Jomvuo+gdCnyCg9svh4tu7Jdg0F+8j7hZJf8JgwSJjjXEEKUdjXM3Hj2w/ArMank
EszwgPdv7fkf+xVP7cTWQx9kvD5ojLvqXEK1ZowCjNnGo1TJM9LhN6JoUf5lCNx+
srDA5pXuPZGNbZkgmE7Vytb64dzhxbp+eM2cistP/UBLelKvuk1VUYvRDL2A7EvX
HLPc8MG86GmT/3hj4JFRDH1+GdFNu0Fz+JSWHEojZ6wbbNqTTcgAscN3Tp9v7g9b
hZ7XJirhF7953V4huxvgyTLxAgKwi3d69/0UPFJYBdsNLj0O5oSXzC/P+YZ7adj2
Q2yS6IhoIKMIZH+dn6uMzheM/GC5XU3rDuMY1KFuG4JPnzbMHflhz1APgSnRwx7t
Ueqk7pOK7XbHEAx1lTyfVxyUw6vnmhhhfS2kMeGiDY70kN5zV0rhaE+SQvhXjszq
cr6jWscXbkUhhyUU2AL7GDeAYy2MEl7+LNhv2o8RzjxbEVD66bgJRksMHBSYRc/K
1HKf3RJI54S/xICYfYbk6JlZFaY4D48qntMoSpOjSYsWtiYyVDA2ndmf5iE9N/VZ
Y0ruHfno7wz95PDw5ryr2PRHoxUn/SOdjY+IvNaueF5PooAQiSwcmdnl/2lNIPkZ
MfIHpNvWAVXx7mrY+gk8ePLu35/xzIwjXNeKf2+XGLh9sM7ljQkVSPSBsqRO+Xot
Pr/oCAjmIsUEZ1ac43rJDn5wznDOovCiJtBgYSb/lu2AQ5uUyth8Vv6qP3rkrmW5
ryQEnXirnyOasc8g5M4rFwNovFU8/TLXAhSTum1BTsLlknSevbR2z73uMPhUQn0G
RH61UC+esLfbPXDIIPM17UgtUZYgIt7pDYjuzkVRDFCBwGs/367G7mcF2gxZu8dt
GKQP28VGpW7TWd8XPRFf9dLNmS9ugg6oT/0zehY8YBc/pPBD77uRoOSWfQmZWtMJ
Ex2D/mFAltodlbIq/TGaC136HaybYh0ZLZ9h2SCixnckutpc26ozGt2RHjahJdZt
wT8RlSegMgpZqE+AGvnZHNAnBqUCGoX5NIT7wsaGSFAz6lzoDDgs7PXK6lI00wzy
80q6iX1wwCxBN70jiHMXOqRV9gl+N3Bbi/AMBOpgU+q08Td+p+OYeMeZz4kWXqif
Xqba05olvtHUUwky2avhUo8gWMS3qG1T4GfWXJqcdKDtcusGzUi4a5sY5sj4USqo
ugrYUHcCh2BPk9AqIe64PVGUKOKPOWQsxUoK1balFMj/mdQnOHvVpy80FK05+OTS
C5CSgS/xbTQXI1NYEaUHewqSnceoRNB8fIaXfG37n5pxO6IbeFY/1Zw5OwisQi/a
j+CSBdW9RcWukscyofCVKDex8ZE5bkKooDTItiYi/yQ/B7eyTo8FZd0y1cwJCzMS
2zzU6C9wwIy4IAYOF5TeHWzUvlGL/2KAqiru1/CBrIwWa4fWEGzijSRKcvXUWq2R
K8FUWthZLoUbB1SNxhwaht8CvfiE2Q251UdY4KNEitSsJ09pFnB5Rr4hj+5xM5nh
mZuSU9QCDpgIXKCk5zTuwk16y/gjiDCdB1qkMgmgBRYGTpoK/ztIk47qTYLijWeN
LOtpSrxadw7dJLaJL/TAefZUEblORW5Q/AjNcvu7RjYBfinvViMpxbaomTSlsZY0
Ftd5AHrdAdXJ24PoTFOYasLW5wAIf43hCCTAp8I7XNzxx6fLYXlFrcQLxdhxCjaH
vgcz9/T42NqGrp+X3L/DYBzofeKM+ty+pPKebrier+BD0mholOuzfvcq4HI9jst1
qg5Yivd9s7mdWXH+uu0F7b7pCgEIPzSvOAJ7adxM+fCunypKSoGHyuSi+QjgT0ZF
cigFIGFjjzVJf0JUAaaooAG/kn8SpWs3NvamTfq1NFRnH0QalLER+07eZ6VbaQCi
XWq6zXZktKPDJV+yKco6NTnVtrsUoiEetEKl24ewVkKvxDcLMQe32LVO/pI/9upd
cuNYEtkEtVAKfO9jVAFcRodbJiTM9a5JtWF3JmhvoldNZF2mpZcWBviMt9MjYSnN
E8NkuqQNwbfYv0UDRbrw9NptSRRibgGOwv1JRMn9A9GqeL3mbYTfO0C00mG2XcGJ
1q6V/6Nrpi/Yr2exk7X2Dy1WLg8C8FRGih7BBPTxVZziH34xcu89MfvauLW5SA9/
WF694jxOjGSycZyohv7ObbKZL+rCMbIFgUSUzvwAaW0ZAaXMZ9e5FpSvii5y7T/q
BfWzW6WFipjMxfdjFKdeB6UYlAzCiRuYWzg+/sV0vRgDOjue7GRh2uhJWQ/n4TJT
Z1+Sx6xod6mXWUVq3/+bYy+fWc7Gs5Mnxey2tnAqtRuqOzHrngDxWd8isIImQERb
IPfy5IKx/puKpInEoZRSgAhodbnmAAtj4URpkebBV9FnjebM8BNP+UXlOz8QAHB4
pSa6yDsOMsVg5MLlJ4W4bRTvvh/84AHdVv5XNCh8JaGA4h3AD7WuYHdjawb7yCi2
cYOYhtXkaLfIA6TtaFZZCcOgXN2TI0blYAXI2wBf6uOydY23YwR367Jxf22CNX8D
/aupHg1iyf9Hfd5gintUyMv7Gy9vQYgUgFTC3JwxyQ86d9ewbZ6YWCAaq1+5SzMA
miIx3w+rg0tfx94KV3xlRPsIKps/B2Z5I8UyeeK0UvgyWZClMF5dmeHM7xjIS+ya
1JobnDIttM+0g7pMVW80M+LgPynmT7d42Aof2qaHaBoOLTfyZPLDGiplWqvrWZC+
uxQWzVGJ1yaGnpL16TKCUaUmw7GslKTyT0mIyGqkn98xS0dXdaDHKWEXrLS24pJ+
a0mz7mSCJEew/Xa2EetY7wuOMCuSARau3c6ncW8DDv/SkHSjvTrsMX+svZ9nh+gp
5/fyHKqdViiGNgaCmeZwrYvLpUIpjnet8HzLrSKC9Eol0jRlfMvHNwPxWrDGG3Lt
pfmLhoFgWgdHUreVowUAN2vcmVOqzsQGKZAAMlKwoB8ec/PY2yTvJzOjlTLj725p
lfVliX4wpVdtsSoK3KQ7rMrFuLlADjaHyoV0AJUUyztRBH2V8OXDI6ocRF5CwM7D
hNDYCkpnAJC0VMH3kAaMt2SPhQn6K4bgyni2ayUGB5SdcjxsXj4/Vx7Ywzknhg1V
qJsknDEdeIBXbjvHHwVjPS9UZgTtnXxBDdjM59cKhA5jyulu+XO3xAaDg0g6IGDR
7GrY7OZt2Sg+mZ+WmM+8NzeCIyywfGFMY7DwaXvlZ8naoazlteocuVrHga//ZI2j
p0NjdNGKMksU7xTI/SZQ7387RDcqF4Sr8q/QpoTvRC400if5RWbURVh9xLc/lyxy
KGDn1X75fVBmKmRU/MyEhPSe5QPE27bQd6+wxUWmo3d3Jw+dsfFzXSdoZePAa+J3
ZIicboOocrFgulb9NTEzmZE4ToTUa4F3qpoNtdlPyRbksVoARhQQIEY8VSzeZ5UC
yF7Nvs3r/hvOFxxEFZXWfcfkpleVJqlkIsHzJG9CNDClyZ4xpZty5x1t8x5waP+v
+NgjjRcR6/u+XB1wXjNFz0ksmQm+EtMjblw4KZcwWjH4wSApmsWZM9HR+wWAno/x
guprEYFy9rZJ605lRiKBjVPMmuFg+wBzbuLV4Yxmty3CoAcBs+eBECCbSeQJabDh
rt+xA1N8RL+GA1Us5bV1qAluAyf9xXKdUZkSfOMIssiribpkmYoJIheXwl40ZeTi
+Zr0kW5p9Pulq/J2PVNJVp9U5sqBjpZuo6FdhoacZTKEGbySV2FdCqXCxj4H7BXQ
qcf3+TPqhF6yHm9nCzYsShTwFt3x76H3aK3EzL7+Uotcqof1QMDoIM/41+hA4xuW
liJIS2B/+CsVFXpqijByQ8BfdrHCmiTYshllgZ8q8/pkI4TbnspBsQ3c7jJrrEFU
6EULZx7xpuLinuipY8uxB4T8z/7/Aemq+C21pdZt76bz0RCS78/R35J0vX8HUXhw
f3Bv+Gdyi5+KW6uwXaE6yt5OQwSViundNXn8xqQFNfI6zmdALh4j0QnCU9R2h1O+
/4wBBlOndUOrk9xropTtwVntZvx2J3J2mKbGXSmKSn8Z6JosE6FfXzyL8ah2vwSq
SCQATZnqDKjASEZkGoC9Zb3X0oPi9cPP1pOPa/KXYc3GJxxP5UpW5sHtuTbrBJgA
Zyo+uOo+lq5tfcf0vpK8f05flnAMXbvgfxULN0nd1g09+kdmosAp05QC89kbMAOe
2W161zAIg9WP46PXMAT+YWD/ISM+pLm+gNFXbsCsSyXa5G5SYlqa0vNHiJzLjHJL
W1zCi1Z6Sj3+1CMQEP19KahvhU1kbvcLqyByGy3OimlHDGSFJjPm8VJed2MyGCy3
+AtdETPEchg4qCTRi2JG+DmxmLQOCacfw/9OflIDxIWmeergwIz4JXqt1ucqNpHr
Wtb+du6R2E8mpqrX3PTVohnVlL07AkKG3Z4CYSR6Rq2+TvolMojewJNwb8KFZ+fk
oY1/8WcGYjvJqzEJwabMCy3oWaV29SEhpPkugrJuPyvp2MWiE0qKpJ+tcaVrkY6X
l7iwBX+6JBeBl+hW+S40CsxpQSvA0hmJDV/ZCjBhWSZB53TM6zz0Xh2EFqZtBZ3T
+gPhb+A/GMSW0dQGDZWKso/dNKGtcVu3Qz7GIIMwYCeFsVx/bZWohHvnqPejLL30
oosM9LYJ3OcR8NWVMh42fqPIS/Nep+Sec86uf7vH0RwKOD51Z9MEmC2aPd7wmmNN
ASAGTJ6KFZ8ZHNii3vQ+e/koqxprpbOtDwJi8SPve08hRTiq9EjoSSqYQZmdyolt
iHkSt4aBftNaqHzo9T02L0bwAbspX2WfnNSF3aCpJt4xR4vMCAcZ9lUcnGU8UArX
NDfqM4SjfhqBuFJo6oQf/JgbFbAkp1xJrShZo5Fllf6naLT0lN1hRSAMzaL+qiiO
t7FbVBNz5SY6u2dxM6CGxD798AH7GLsn0ieEfXyYAAhXgUCSor9kmCP2Rfy8Zs+n
0K7qPPsmo1gdFKkWQvMAc+gnt59gOPlkiJUdE8rRWlJ4e2E8CBsh6OSYyi4wZ4hl
VPo3cOHBJk+A+RDYHRcuDGiq8MSGRKQQtoAb1bNNQ+LAtQHazNxAIBk3uGh8zyBV
hHWXuQ8BF6Yh1h2IELeTuzXOJa90+lJtOaePuF22yPnerrB/AIuU3JHhMnibWuG/
nmQl+5xyoXVVpM2rVLVfOaVqW5+TjZf4HRzc+ECmRe6LM+o3xH72yjMfit0axMh2
pgB0WbKAD0duGMuH5sKVXiWo0rtF7uv1bqpzhRv8l+TN7oQgzrb3YuKuHN467njY
QkdczYL9TnbAD9/e+Cm70Y2y3n0JbM1OZbFVoonp6izBlF3AxWc7a4z8bNcz1XtB
wLXRInarZHtqUZhuRBiuXJaPZX3C/NyCZHQ+ogvizRG5abMe5Q5p4g67019h/f4C
nscubzSE2KdYU3pwKC3BEQVa9GaNNaqfT7/10TXys2ifNER9OQWTNzuJ+TLO6nop
kv2Q6zvuvT8MeakzuUHhDhdJ6DGPeJ6987b9mFIxgDXMfvtN80kBlTGpv0rQhJty
MUD6bA/f3kzRwbLZx+RmtFVGZzPwpUw7fbJy1yRrY86mie/tDvZPBckSgUnKUlFL
JHUxl6VzCobR5LUHAaBj1pr90IU7EuzZxzJep/ZULyKjKkH5Nd7k9oacuqF/godh
lTWOxLE2NFTWSkCT56BJx1taAtMyB34m2HxBZ8xhY2arMysp5hPo4k/C7DvRMYtJ
Rd9EZM/zxdYXOiwE+DykzFPRG5FOhi5czpiMJi7LVBzbh7aroZXEplHA0BN06sKt
QLqdZ6A9wBnBki4z7S9G6DZjZQSHt+X5CZmfTBKMe6dzHX846iKZJcl/UQll9Tk1
qCRmEInWZTuvhMgA7Q9ep08/gkZP5+3XnXoV3eiRtjvjHo/L5//JqXKax4VyljUb
tKYnEmo2psm4zu8mlD2WP34Jrk6++aggYhnboeb9mwvQNTcsM/aHagXoq7vVOQkg
PmnSjmLTiRI+ICoAn/18JTUW8lM23Gmot8Z6IdhxNTQ0FN9uAjl3lX5V/38RjelK
1cDcwdJFVprDemMG9Fh8lAr51YvnnftypkclN8MHUvP+RjXD5PBVivvSqF2nPcKM
6qdT6kBY0+Fmhhy+Ry8y5xYQA1H2uhwJqQrUzbUclb9E/lRJaXfP+dSQlbDjLRJt
oyXg+efhOoOH0b/6h+kh4gFTSuj0KliaKebx/+PAUo+pfTmZ5wsRo6F2rBURI1nw
gkIkeI4FeQ69m25alWdcGFK7gDBIG27g3Z0J2gHDQSP6UR42bgOXLz5VWjfYiARN
TfKNQUQBNLQm0JsDNw8ml5QkjTGIVIAwzQUID+GpgB1N3GQzthvJd3fq3tY1kJGa
a9hUmufs2hamtVIBSb0Y3ppGhv0NvLWPW+jHzxJJWF9rogdtxI8dyw0AqlW0HBvX
Ayr6QJzaoOrVbC/qqD1ZdFcLb+Mz1zAVLifZzPFF3DFa8IURDwUTV1Yo6NGQ/i87
oyDacXXTSYr15rdLKovosNsx61RgochEpKdT6JwvTkGlZdguv8WwuFv/ORxUbJjx
S1FfhgQzttNZRfYnVIfqtjSq1SEr2n/fiUkf1311VDCri5bQDgFs+X6Ow1pw2ngB
BNmrfvJlAj7lyiivCMHFHoXoeS2ewL7N9uEN9z+D4MwR24N//N6A8etqVkNb+8k9
0cPpCt6E3EJAh7U76Mqq3k0AooY9863LoXuhetgQBKJHin4ki4s1KIMyubeYq9zC
j97df5rW3HWyGGkaw7++hFXquC6GTs6unNQJBhZkmWwNW+FW6qYy1/lKPiv4tRYs
AjvKQfGAudIbhxhk2Gv/ZK/bwC/ORgvX2Xm92iDugwPCdd5p2wgQVHDrJJ0psuWz
vkfiQTj6fcF3MA13iCjCa9oY9g7yatxL80HQD/v61qQBDUlDdDODwp+ObImbMIS2
ncZmzjc/IQejs3sebTVL7tlxAJaoTyED9s5buuTs6NFStM38PfHGUyRu6PxYTdkm
MMsp7rJGoVcYNihUofnvprAN5stxhrcN20EZccaIuMmfvvWDSIiU+/tgh3d3qJfx
Tyd6Bz5sGtbW1B/wc7/h5CQGUkS35y+HRODhS4FRWgtjZdx2bvChI6RWiPoKlYFN
elSjJA65lsLiVzN3y4kBN3QMncaW+MgSBhkIFVZSfA0cfcAAHmozTSWPjKxYRWol
ZnxkfnrfhozZjN5XQ9c2F9M0jxCtpPUcgQQYOKFLCJgFwpoUp5+9lRTO/+SnfaEN
B+RO24SbjSLWP+vu568yqvmTGr4o2RegWrnz3+k+yBer7GMScTaYrw87jL4cQScc
Q+l6DM8THGnorb6Q/DSwNi30Mv6hOsQhafuNvn97GkU8023zUXJYROUEnd8cnhe4
JcRueIDQT7p3Jxu0siPwX4B9GLkRMVY3hWCYZdj2A7LM9QyHE8ztMWXPb8hqLi2e
BQu4esvEKhFT1B3S483XlWi24jZCcXX7a4z3Mu6+meMtiyjbN2aL7jGRpvCiJRKQ
Z7LPqvYX8pfTmmo9yTfi6+LRytmsf4i+ygS9c/OqSNlpUf0sK6FhTE8428fJGwfU
741+hEUWlQ8TFhw4FmJZC4UFztAOjfTVH3AppOrxsdBXs0/vxCsyrVSV6S5sqKyq
ARazrROC5/YsCyWOuBximGLStLKiO9FtekvgnqcIrMZvTudQGnSkVlQVZnV+sBiy
RYO2zfqVkCgmxCrhZbfP//Ir+BOy5xkRjz+9W76xjAjIsRrUrxbBJpuBAaV5IKdR
QmrutnYw9xKR73NQo4f44Ex8thVcv1bFfuiKFZSVsGZ0Lqd/CHTcAjny3jz6Yvby
McANuxGTAH0UBYO830weXVWL+ai+GpGB3YX2yyBnVtt7KSyFeqZuhygGH4gmlq6u
rX3BsGdBfefNdrpJYNyMUQVzB6/m5d1+USD+X6pA2hlNqgwQoh1QM99UATdqQ2Ir
j99quM+0P+BZc4+GUa6f6JnydlTczo4N/yMffWBIzK9O3NncO57EZcslGED/VtXA
B7ykGS1fzSimBbtxpekEY1j2DrFGHxDNsSX9cRAIW/dnc8Xcw6bpeerTs2lxi/EA
ERDs+dAYfJsn/FFlTDlg6r07ZGsRIieaWAsDTTCH4mMPn+ZuNJEDJ5iy3mrlpL/B
q18tl6sldlhxlk1ZqvwJJ9ZVxQelSggdcRutA5XOeAGAvq/27d+NWL3hbZ9gkQvA
87QCR0TvwUEPBJSoH/rgtA8ZgK+pHjOTsWOliMTbEZjwk9GevDEWphr2liREPAJ/
IgXVOyw1xH4yvFlPEbZ1G//aDLiT/kH3A0sdYu+4OwhjNh6vA98ZJBuKrBdSMYfp
gg0Sbr3OWj1F0xbbbMxF05wH74mdiKgQ9GM6SEkSnkrP1LH0Ha60F7bTkYFjlo1O
Bq7GNMetNMozmplh9QbvhdgqtzkVuOnwpIv36Q8jUfqg9/BN8URfAUeH/sBQnNKr
fIEnnQbLpHpgmPAid6FsD7HsXvJD82HkSPFIy+plpqfn7kxYG3noH3Ttbki5rbVd
XJpd8GCGq027vcc8WF/7207gEvLr4eQ5Qi5ALevVoGbYxx5hpl091nggSCY8lb1D
qqWgXCGkJmKZqxTHdECbAg6LcazJ4oI3eTnNCDtcRfX/nTnP0KLcgHlijebspOms
rDB9PhCfPV3zmC1TIpBEW2D5MQQCTr9J+lcaEOHRdl8fGz8/FqqzzMsELzu5BKjo
JFeV/0jAzLy/mMND0JpXndnmcbKd4+e4pILsKcSxyaW6zShfymW9w00vGQmUK7vJ
HaqwWSq3mSSm8KOv8yLBrgqcl9JbqYU3tMXxK5OOr3sjOpg54zneVkneArZFOPXB
sRZmyToPn8cE+6lC4Smy3RRCHWY/68r06JTT+mxSJ+WvyjRDfvfpDOXppo+VndNF
TZ8ryrqIJpM2OPSKYE5T4ONPS8xebu+saxVaBhnmNyM71n9r56OnwzTz1ltkfB+2
K/UJrfqUBeXyzqbPfdZ5H/QwpMDq+zrB2GgegIxiwlfPz/KoyRye7Ah2OHdl2tIy
iAFew+AVyZXlBGDKGyjX++oUCLwhhnT9oTHPsWqDOJAiwNR7itibb1wut4qN2fcK
Qf3T+KsJFM7LbjZHkvMTL7uW+nLRBW+bB8o3Xqyhg3rfnGyXVXHOMpWF0d8T+C6E
iYrxL1tzR8/4NaFkAhgpYOQYub85hBpn6fUMLqDh/6kli2x8fs78KgnmJ2lASqHn
CG9oo0aqu3Tm1HrtOs+49neS/dFggSKO0WiO+ol6GnrgZQeV+ujb6vCk3sm7Hw72
e0OnX4uHYHPG4SPLcSD7UaHxiDbrF0xkh4E9Zeoyxl7PPnrtPAM9/p424EqTvxMk
Jn3jX76WWXOiVsR/7bss6UTgftt3wHZ6WoubNs+qhikQOeVmGldMVw8Rwe1CL3Ni
l+mA+ujnAUF3UvYcKleNYaQlcYe2jeS2YPFnpxCA0A4SdF9PDLw1ZDUyHazpJa4A
5hiZkMTI0UYzj/lC2gBSe7D1UR5Qvr9l8uZjvKvcYrvB1JUpm6QEVwEC+tNpZF1I
oyblFwvju1qHqz5IpSss9P0ipXuAcHDoaNqdqSffWIfI9CcQV9EicWqB96fUoIFC
HHyqw0M0H3f78BYAm/hxoPEGKP1Da9FPk3ELC8QWj9fGoCt85zqAoHKIP9oj6DYt
LwoNJPlNJ3Mb9P1+ovDuUvp0ZW+1wxBy+Z8vQ8a9r5GJrOwkrI+0FKxa7QGP8cDn
Qm5e/Vm0YTMwYM1Lcx6NTod431i/ZOtMaG6zv/5jzYh0WxDRTfk1UjdqhvRrxn91
UukWn0GGgBZSzbhQNW1pYWG9UMoSaq7rcllbu/oqf+rZLSzDfoylAQIHsbu/zt4d
/nIJ38QBnasyB+X36313HTzEOYS0Gev2AbcAoCdKfqHULhS8K9QqkcIyFENBGI9J
w5lekGP2VP+Wg6j3SbrPe79iClV4U4bk3Txl4Ev6yMkC2D5Rd/NSoCkyU55K0Xpp
Txb7dV0M1no2sB4eAzs+r2eE/D0d+59ZchV/rGOiZoXsx12pGioIHck7ymqwzFG1
GWTiGC7ZRmBU7sxYgxoEpOWIF9W9nrlH/AnAhn2mkSk5EvsMSDT0OcYbMqJDy4HT
Aok3AlGN7gmAJZf+RolF45RVVKNbDE8Z4Rw8EbzfcITqbVwDwVSugb8QhrLDyWro
oT9u+BLlLkjrOKYMH1Ki+RTcwr69mAoQjzJ4OVVuP3XFLZDa9Lggz4A3NS+S9NRl
b88+3bT9Ts7ASTHmYo/WVaSwyyN6CJWm7/GQw6loH9Zgu8Z9Ght3i9FMvTHO7mEE
wPpFYf7ML0CvbmYqLixqNQ69CvnqAcJXge6WxsuyFxpYVGxPGcU3PXmzpqyL4yaN
zZKRNuzwR2G23rl4AODI5rW7odEJzf2mtFDCKXd4FI/de8Hp1stxG5CX3Kl6MoSP
C6HKg9/R3Vy799Ump2lwM2+qrkI5VHZHMT75viSXpQPjLWIb20kcr2xibGcfsQWM
oAxp4mjzLXEsi1qtijrc5KtTd4PTSg0oZNxE9aRd0RtFhjnNCRHRqDd7W7L1VbHn
ulgruyqaafs62YWX2fdvEOGdXQV2a4rJCioZ+8ugqPQzY12QgNjYroDnFFHV0KhS
m+SAIA2V/uov5h1TC9Ef/Ee62cZp6bnJqYp3YeRbqIGpaR+lPVCQiaztAX8rbM1s
R9KM9NbH36iCz6UeIWopxJTRLBO5XFfDaFFFVyzOVI9uFfBlpa04cUN7dnxaBhsc
0BFTTCAqtDwWkpm1PY/t0pmSsimByF3/S4UldRxQrrVSXm+19OQDowAY8afIjbBb
y6vLyN//DzlOC62GI94LVc7vij5O0Yeyt/2SwFl/AZLMUK8/d81YOJtHfJdJ26Gp
dLKGdW5c+/gw+RNDTFIRIWu+XkiT4QaH1K4QtV5MQaP9n9e4te3KcdlmT5HLLIB3
8ktnVGVRnMjPhaUjQKyPr6N964TABsdb/upN3L9leD1wUirNrN1G20Iu8AQVmuUQ
LFpOW0wdtlw+dnk3DlNCIgcP3wK52JXbqMJ/JVdWsBpvYzI1LP9afo73UoQwvjh4
DI6zCWBaQUPnq19+JstPfqXmMF4DHuqrayOlOkfbijn6r3eVqT9grIZHQvwx9+f8
XLTEahiBG883R9eZgACUt6KqvUgjYY3BRrz+HlKv5QvLOl8HXhoPcpQjjJ+bPosl
S1bCWkVb+F16tULYrgjkMNn7jaMUBN9UMC7UhD2XEbpe/k+QNPsGt5S3bFBQn3n+
7e0qzsuIeATZcTDL9L26JpoyJcK2ERavAiaqG/IIeV4rDtd85RoyDVM4ASJ5A9Ff
04ddsddEFRMC443v8NoS55xUTDpDFTghioqp+FYLocIEaJKR7FwWA5MTv4PTSG3w
EMaS/yo1jyacoYyBtLjTzaHG+F8AmJF1akdXSzHR/ESqHMXs1MBoss1G2hwBxYNJ
FtWOryo2Sjq/68WVfEHXyJxBRATDgxlEjDuhx6ZDF6ER5n6qykNJr12wF1jeoHr+
hRrsK/aT8/eDtqrxsXQHXO/iFrjSUOCfpOkDcAc9l7s5/JsjcjzJRB+D64X57iUX
8iamOn/Vld3xg7nvO/waaiBtTJTd8xt1Kt7SYFWw3JAQnsWoAOqMmEjjRyDhcFqz
TDZvD+g1fPXEMrafoKS9Esq7RLcXjt8FQDa3Pxi14VZ1rkSqWTyE1zRefuqayHZh
e8rEu+9KoWsMmOJcjWZd14HBLKDRzjqU0wc4WaOAHefAxIDbEezuEECU0bnZ08UC
KmeZ95TtU6Qke/uvIrBC96lSM7UHOp+QcxDLRQTi0IFRlg4U0h1Ex8UOzQJQLjG5
vJi3EyM0PnTFNxQgv4yzhjNfxTnmEA9xfbEqAIrhoF3vWyEXp71Nf+fobtTpiKgw
pIA7tEEU2s7B3jNKshvfoqV22db4A/vl/srb7CzjUx/ua04+DG/6cA+lG+MXeDWl
fsGTZC5amt3aykYKt9QYu+cafvL+W/FGWVY+FRLkn8BD1W4NW+LmiwsYd6P4rOPp
EMk9BjVCjMZQu4yrx8yb2hNSIUE0zXquMbvCBMyEWbnwcIrFNXkObRqQC2C0EIWT
EPVTHPA8zsyRmJ0KcGYBmDaJAXDh4SRQNzTCD5Ves2+SGlIfrrGf+Zs1PCtCo95m
QN07aRt0cHecMDJ0vVJzVuyy1V1T7HFkffmOiSpn4u32g0TJ7wHKyvzqWkYpsC6F
VK9MYmpbNd4Dsys+NLwH67hxQeDQZgSsKEnUdtWbXM8Ri9BnmeDpG9fUZbMRi6LS
Ccz1oJ4vkt2K+YwfYxRGi+UdS5hv0/ulP9OKh5dx1CNhUlD3TGTXMwASokvxlWAB
aSn8uqU188tk541LwIY/bKwXO63rg/pF6VdUxsK1gLJ/uv+CGMngfo7re8mJLueL
ybltSvmVYaFWTu8Ru/JEOBvPreNS+QZNZCBXFyG6/mp9eLyvxVhcPGLGm0MC5mKd
Gw7Dbts81ga7LLcETeRWKgfYw13Fjo1Sb8+VqwntP9o7YKvRDwF1MiY1OcIhKSFr
Lw7EFOd4+/w7XkZx+pSrONMc27ZGYtyFFVEmJu1G2z76gdS2cDC9A6WPa/nDJZ5I
ruVGKCFORNn24GLTKZDnpLTj3DccICaSDo/LZmFCvSC63t1DVJ4eMZYsbEWhdmHp
f4NEn2ziL+prQ4vo93z+lPLnBw+R2vCdQUkvvoX0QUVX5dJA2NXF3MZ7hUKKllFg
llFgNU9wm2hBxYsO2yGEictkZ6FwR0o5+NvJoKKSz+hD5t47UyyE5Jw0FZ+Vu6I1
dlYdxEc50rRIAmOVvi5jVNaS/ZCzQWzkiAFzsZ40sRgpr6wIZuIK+eEjsRAIPImN
nDBO/RZ+lwUatcxB2jks6q6I+61yJCs7Htk4MlvlAhS5RYGqP98abarDJK7x68TF
PHKusQixCd4DWfsqxs1IEaBdwXNuilMe4gxlonbJMP2l+oVW0uRX+tdKqeQW44Tf
r2G7UitplISQjsLHUhQawkpWrkYMZruYDRDHWryiv3f2av5oAJ9mYEkzmYai4UVC
qdtWSg0M6GbnqOERkHFczTJAAfC97g933Pm3EiIKBrI7uxXewXCWT7WWYOQuKgEs
+w0fXLNXhqaH//XumT/JasagL/LDSF94JZB9k8PnWOOAY2xdnaqiF6C+vHXROcGy
qFmyY9i6W9Dble31y0DqBeHxW+9atf1W5CjdKww0VuF8SIdFmm920VuJxtIQ6MVK
HWMICXGSscPiLk5wGoByXz2GKYZT9xq2v3Aam2RF0DCjsAgvbaSEdrMXAm6w607x
3r0DpQo4SBFyx2vF+mUZUtNAiIyMgoU4wtTCfsNdHuC9slEKdCpYfjXkYXpS4g3z
eR0hyF8rwsd34K3O3PobD4a4kBkzy9k1/NNvKdQ1cxjW+5cGyKJTf+0zlJSmS3qb
2NFZ15VNLWqj+W/L6jpnL2ZrjMpayqoqi3+gV2L5kfNLpldde814u1BAh/I5TIw2
4DJrnFCmkNh8Yvhte2VsgT/3CT7IVB30IHegsj3EyOj4UiQHQXGrUh/GDpluAo88
mvMDfCzsIolzfuEPQojCy4GFiRo/AnwrOq1BorrpNncJ2/m1kJ3iPz8VlIT9zF84
3rG9oswjMJFI5KZ9HqM5N4F5WobWh2pBrwRbfMUmp8lzJTUsLemnCNHTwrbNG966
tSw0r3Gv3lWpApVQ0tSocFioolvK8Xaz1sFVxaEk1eSSY84EfooNNj2G/ccOE6eJ
Ilr2FKvH2m1CE3rkGXw+NSilUy/9lQJ3Cje6xhjb0c7IS1jKvO0LG0XzOoBrsJMy
B+6nJukzLYREIM5qtq1qP+pA+GNG2aOnjDGnwixz3wr/2rLzQ5G6fvlgnmS/gBKC
V+F6tYvF/ZzKwH3LmjxptaC6LzAd9nCOxkbEGQYHIJ/Y4J5HH+rgoJXYq7IrnxKk
kpvsdu/XAeWr3UXJtXGqujm37i1cMgtim/zgOQXAdnv4x1cp9oXeke1ePVFXwwg4
lYtnrfVkChNgaH2uT9b7oJIZGJBsuyrsSbRUFqKQB4IwxC80FtQdgPkswHnYWW5k
KQOxInGAz1xao+81FUAKh9v4NIvZHag/6jzK1i5Rfw+KEOb/QjfUNufUXBNwEGcS
zKQYS4p65MmPgaXwL4hSiyDJcWkW3wb4bgLUb9CgAupo9YOh89yWQ87e6wY9shMR
j8OMXCQuhjW3a9rhJ6Sxdj+HUqEln+fXfPRMLKQZ+DlkeRaR8riyRBQmdrnItLap
8gUTlFnEcDXsE4RVXEEkjLYG7TWmimgMSXd8+0E0Uq7tWco9+lEfhemsXr2sObcF
YKY/zUDmuPkejzvujahNJnO94ss9SjO7emhwjJq+95wcI/9O/+P6EpnKfJUoXGLS
DURqb5iUCAx0tSUyi56V3PoowkUQ/hkGhXAL3ZB8WhqwnOHHirYT8H1XEEbjYcIO
f4BrFy8kg/8cd4Lx4km/xNZ1Lx+ybRXcA64VB1lygqPT+JgmYxgC8rcn6PvINyZJ
Q+e2eT7C/QYLfEXt3cWQyMYiT3v6nKGZfBFXQYrahLDmWVqU0k64/2rQJuAnWo1a
UKinJbrN5YA8aSbIqlCA5DX+bUNqdO5s0KPQu3/5W0Gjvjc1k245JecaaI2xtb6Q
2cwu3c+Kez3pl1Bk7mc3TOdHFhaTvUHIO0PO7/KbdaFu3JshzuRLXyuu396RxE//
QUQNuqylZ8mW+rEdNQefsbR13cA+Y5J1VebqfNwVn4fOwwN90YuQz1ZFxjNoTwi6
0l1Cj/jwHoC2reQXtgpZnDlIlR7n57af/0TowcGWKVlhPsEprkbeRgpdalvh0R2S
U+edESdY7tSkbvSVEkj3ip+vmQ8W47G3T6fljS+0my/hMjFPDRBQ585BCT5xOB0Q
120JjViwjIVDDWSlnwA3EiFmsnTA45YGKQb9acivmrJ53pYkRAUEhEWzpwaS2DXf
TFYOzbF5/qZxzotpe0fLgx6nPr3QSzjJkVznIW2LkrRR33sQXQDt5RjFTTzoyhT9
AOREQN2zGIfgUkdvSJMkvSGEzAqYH1jJpelXIiHLxSj/uMEuC1pyfPywMyvMKxkB
S8p2P547zyfhXqARqM60jB3KG4SMo9T1FxoiCd1OB69QvnYPr5QAne969yKPtRji
OcD/b2hdfID36l6uNfesKq4lZ9wGhE5N7ceM45TqpFvTpgrYZZ5J0lmtgkI33qyH
DbGsM1h92eQuEIbwN1jk1jxx98YukZGhPOMOXp9VWrznNewGdcQqlzG9cGxFI46Q
FVGsnDDbBukTQhVOfcuzOwO9Xr+qsbImnQe3SHPmHoPGNvQe4MN2JlPxFRI5B37b
77Bjbrimofk06RMz+e4uBrriS4A7z3uO7bI4515TfcRxY6GbvxgCaJ8FctgQR8Y+
Ex/tArLasZsEChEn8pwFQeZZLEj6Hif2spIHVyYYk4CUWnx4Exx7QCCWPlXSvFQu
iteS5NpRuH9yim2uMc7o5hJWyAju2c9uym45QShzRYgZu7d/r+PWRDXrdLC2ItsO
S0YVoJ9qE5bJM1vBKT134Hem8yOUiJ74FTD6T6F8znay/QDSa9zSuL063vFRkqaj
Rhlws9M9Flv1q5a6hM4TpVStb6mPkXI1hU9skbdYpIQfBxnyzkKzvY3XotOdLW4R
Po+25w4Pzo9nZ3Mn8YGn9irrVHYpVVxAd4BqIaQMCjb39SeN4eZYK+VyAMeGISVd
TMr1nGMxEmGd3dJ0V4CsR4TjGuaWml6nMxh2B908KBcsE+zSoUROSzs7Vos1iNu0
+duQneteo+3bwxhgdzOpDUFvf1/e9b1ixgmvGlG0fqN+8pgg3x31oBWBJzFhjdkx
QB3fPAjW/qzv/SUux/lqR8t0b3AIHDYoqfk2ND64Ev/MJUS0ugar/ggbaQNngIfR
D9iwMwyRzteBTUmxVbWYOsX1j/e5OY9k8HYZdRdn3277XXg1M80ybys8PsLBq4rx
s00LNoWyMkg8vIaU0LYQ2Pi7+kBATiH9QRtcpO8VZ5n+s2OAPrifDCgY+OnP9uy3
Mp5GCiB+Brmm+3WzOUEIJ9OYq7ltctBbUYSLQWdaJ/WsQJcBFIX1Rqnegr+8tw0D
aOOJRk+5EB0N5BOIv21mpQ19bh8mvRHFl531b+UvTmDTcov8ZpeHhWnvAUQPZSTG
/jLV3DKta5OBirPOKRbbpYHXJ1/VgaasDF5fnSiBuNuDRTAfQV2kBPPhhM3j46XL
BRRj44vgJVZmA/2TWf2p1VBE0U4T2mNX1euXJFagDPlGbvKprq9hJ/VjMW+sTv4G
Bzmwud7x4Q59D0S50zF/7KZSAASKuAliweYi256JkmVfh4wT1hyy4xJgXKh56X/r
jU6mlg9mNpe1PozIllm9KqtnU8dHO6ZwemhVGXY/mrJvdIqEoQGVu+eGzBuLb1CX
Z/LBdTUm0c2CVMaz2YcP3Mwpj70zJ7ucF6u0WpYdxaIGtORYd9aI3DSQ0f7AlbJU
62hFvbW/kDidCZwCTnVEfXY9k7AUTzagh3XiEfm/hpodUGUDi7qMZd7Vq/OyrPft
09Urv5BpPbWEIkkzzsKeQiesdZcbfD2x2n6YGnKmEQgdFE/9KDNBCLkzJ+ymiJI7
gWMi62o6Vt1RN/1jGwtFNJIeIJ2ovae5A7EQFJNngBVJNqc5rFh6KWc2fMkiOAS4
gteEbF8d8t1g3VNELZjyNjfjNuEGl9qde5SazrYyEPFx6fuclqEhTt/SqJYy9Jh6
dTEKJ6v0ET9bIehjETmXD4UIeIVdSmnSP4I39mSFbbiEXnTGmkhgrbuIIVugO8vM
6VeNvEHJS7PuXtHVTk5tjt7LSBJZ2s1qElrz2OgA4OZAUuL2g/6vDl9nzTD/DxrI
0ZKergOkXqf3XHXQUdt2PunpjMhk5bZEZrP4wl0eMWDw093rx9W9YTW6u0XIKRrT
GDBgX5IHHn8KgQvdpbmXuao9uOrWb8dZBOzP0eUSyDo06Wz6A22lWKwZ4E/nAocr
on2uZu7NcBMr5h3Mp2djz9MoD5H9/I50Ma5ud61XaCVmtZ8qMLViAWFAHWVfMg06
c8tTD6LgnXY5vJNLKAF+tD6pObMTCjP0CGdduQ76iNRRApu3alEr5/eVprnfU96e
Raofr7beMoUYwocq2EQC5wsn/0hmOPQT1SDP0d3i/bXMthmBr5RJ6fA+mwjxcMzk
6ntmYuiu9lRxG2Wk9dVF/ukom/Pgofv8uaXxEBX5KlklTxVuyZgZH/H9gmD3Fz8H
L6nDwT9+EVDpXKV36LfYoBB/u+zppUC87XMXfVDZTa8b+wwM4o82mO2gypBMqNIv
kF8GvP5Hd8fiqXrqhmOvDw53EBusx0VC9Seja2VsRBDW+ZE1xWeFc2XnJ2WG8qDe
WUgBJWvWSDvuH7tebADvgvqJgSWlTSwuAfOV296EXLe/oyc37ZXD8/LPxXC8Mliv
l/iVieCAss+OE6hU+VsZ2XOzMTgwgfH+pxPitamlGwUshJSCRuzJMHJqiOiPoNeu
NQRajvf8ACfGf3H3MlbAn1EWVGzM3FbWaMJtYD8cwyaNtITfuEXESQW0WBTQ1XCf
gSQp093wbvQ3+NIpZT4d5yEehYvFw1RkATRuOngZiqvir0kFc0UfPr3reDvFg5fW
2b6cYIKBtPeHyfB7a+xro4I9srvAbMmN+5kbrhiBWhA4vQr/ybvq33Gd88zQV5X2
twXyVXA4vqccBaUmmv2K04iAoevy2Ze8wnebeq4DY26cYVKYxOusfiYLiNK3FsNI
DK0AJIODTxKpWQ5c432q6Ioh7yl5/uRA+maSLrl+kxfnkGOpQfyUgEspHl1E/oaE
BWxoszjVBFbGVXxz+6grSF6R8+j2hPZSsLjGjuFuwyRdG4XnEHNCM2lqUzbxApxV
6NkMTPX1SCirQyyDAAVsQL4sccaYKJwBXc429WpQLzJBdEJEmlB5F5TVXfnyyrFO
wpTzxTpQB+3KRIY4l4VbqC/m/trZJv6oBurfCVVfuHvrZaXCRbluwswKWybRZrvd
JkeP9bLb2wjUZHxRr0LsqkONAHYaRxdlFKcrR9ZSVuZ1R/hz+yCsxwz6Ya3EOQHy
RlBQEbCRUx7iJK10t4+XnW82G84vB9wA8i9vRN+NTBU+TgjNwaF+tJ6e6E3YdKrG
wKtpcL5NuP9zqa869iGAMr2AC9fIY1UdBxQX2b0LdCbn7LlqdN/Aeijd3paVOv6r
23iLInOGdqMB5h3wCyEZpcEpd9SsFUa7Taju8sCSCZl/Fpje10BDMy2WyhbtmLHq
K51Iwoc2QDYb2WKVtB0yBWHGddHjs5S5SmF4WxCqJ+KZKqazWRLzngmT+KOSOupE
3LDQg0hc/aRq4zDT+3JQtslKzRoDB2wDpPVQ8yN/mSoDjsAoW97rKPuQ3hZYwuFa
/hhl6ssgNoVd5qIfWWnhFmiQYyIKG8WlRQetTz1T9gZ3ftt6amlnUv3TKQH1IXDL
zA+BR332jEUUPDieYXrEZzVIQSY57GdOFDHq03sqY9GCMEfgMDzxusMd5E6Hyn8X
JBozbtkamM+wWUpFuE2sP4TK9YD8p6TFcdshAufDWGEC5pxHbHyhoISORfkWlYBs
JrhI8CKeX4K9mVUwGaTTQzyKFcBwjMCokcccnwuv8BJ0Aii1pU3bWWpRJY4hkyPC
f7ti6pEPwvIN611FJK1KBgbNU1q6gqtVN1qHP6prDSliXlnpTKf0htIb7vDd2K35
KdaJ+0FbVyYYVQomn7U5alWtJ2dvkw5xgkw30P28T1g0Va3jGhbb8lANGUm6xDTS
U6AJ3JYjd7pPFqwdWmRmpMZ7jzWFaZborPpj940XpZTVH2K2DIjnxDGcc928SmbV
Y1TYxM4NsLQOfmIeah1sYawivtFqGQa4Xd/DWQpNe/dy+Iry/b0/sAnCFnTfZwyL
XI5Cd5F3ApclL6EhPNgwvKgPUvnnR4FJCHKJ0sJbWfplqMbxYJb1S5VrU7uND4Wv
QKeZ7NXUH/DaLtT1J6U8MHZ9Vy93HoUR1FDbLhx/1y6lzdydOrjSdvkjl08gHq8H
AsvckWfyj/sVTY7+RM9/FFbwpj+QVwh30Mcr01nWPXY16vVkH1MfgBTQDHCCV4mH
4JdekoU/o4mpUjYfu/VcCj9iemHSq6VmXRvrdbUuWK/qGpCLjFCUmZzc0sQA69Ov
xYAs9tp/E4jRHpQboo1zBg+fvbtEN+A3M/uCIk8iM+KSYeoQflS0SdjlN5pYgSRT
PMATe8SSbmh+lqn4lJd2bW0V19MVPCL/NZJnKGqnwVQ1ZyicWM3QzwTC6bOaSL/v
m41JHjTVAwp+iY0W3E08zM1VYbdVw8OZ3asiEUYoxPgDmnFA4Jyg5JLvJ1mBY4V/
HuiHOiGP5ndHWpxLVm0jnYWDKOYvZru9jOg2JMipR4otB7r2koJRNxMM6DQYHclX
GiAxsmyCq8+ur0ThJlI67FYlcXpwMJnI9B3Zk9oFsn9jeyebAYRTSjapiKB7LOFw
memlgsMpqrMl8EFsbAFrC5cvYDX+Pi2bE5wRYqn0/NZpaAUkBlx7EZ94J05CK4yA
22bmJ3FcNGZrkpcd5PyVGoUcNT7dIa4xIy6K4q8sz9j42qakeSGYiokgeybQyHhB
ppC4SbaQAfFSlQqIVpJGO1iwrrIgZv9pnbzRJtbEUjpIeohqlfImGBgu4dxXIQek
kGGSptvl5lLieB37mhUEyHxz7353NNB8TiBDTpQcoOVErqlxkW3FlNIBbtAQ9gs7
YSmT9GQDY94fQzIBwptrcOmCqJB14ZeX9EwRhFhAgEvJ0xbp72b2FOakpefgD9NC
wwtX9UXYWsSp+SP3dQaI/pKbQY00zgmQfDflDFsayQNQhMJ1+4K2sbIDJkFKFDvW
wXByf1hK/4RgcdGoPhsmxs5fhxuChEnkK7U6VaAIxqv9Jfl7JusFPlfdKqeTzFm9
cp1H3TDCrZn9unEnUHwyvTkYjy9rxjNzqFTc/yX51q7jLjfA9b9GUai+4w9ntUXk
mYFZZWk0xE5oNwKnDy685irbX6U+1sE3sAQpMteQE8XpFtZB/cchrTIVdNisS+li
lKS+fHKwr8VFeXamE5uJKCY0RE2BNtS92/TNW6VIBZUC8+XtpCfvCBZ+BOiefjtp
YgriXPOLavmsIp7mQxnfSUlzxWGgRFARLuKQIjAh+tY8737PqQuquIt7rKi56u8R
UG6kvPoi8oyyEtHNJ9GMT2V8PyCCgBioA4FJBrlsuXzjOhvbQbIjV9kDi08n9geU
fEKB32cgaC/gItnlJp+LIYYFiHbD8FWvdzRAnfulIP0kahoLZXmOMfGDjxwig+pz
nLdmj6jHT2U7dIKv3lI2bXTkZDH+W2lX62W7U/xQdJDANpH20g66VEK9N8ajEqol
5JZWwizdIsrb2MTiywgQ3+UuO3vSH9/LKL3jipzwrd2RP8LI9/jRwx3wQYpn53HS
fn9TgOAyhn2mpmsoAfdB7WymHjKCGP9OqUIP0lzv7k8oeIrPkAnvLVgYSUQ3syOd
vIPayJAIHugeUYwRkO5E8r+usjqY0QMnUjZCNoi+D7mL1LobXYC/bjEOYUWcMTkc
aT2WeUsbSRrvJjfWDfCv1KzGbVfnwRSLiDKBL1zlavJ1hkwidkpSkWjq2MuomCx4
y6dYCJXPG0nX5hFpiBQcIyrOK6hXpTkx2U8vos4ohPEGA/C9zZ1bbRnxOa9kY1zo
SGNMb87tRjyTLsRdocUwkl++x96hUAeJOSly7WhD3JXu6m2POmnSxCxklfCjBHrr
j4uTU+uAjjWQ+3VylyXoTKEL3L97GHFzzAytc+vFte7ciwLkDqeIVxC2NLjrgYpP
MKhI5dlNKJNBrC7rS77X61I8XTIxtQtjy4qiJ/dQbb1fuu5OOH/wtLmEa5Y+g0C3
dtPsTwKdx/Qq5Puw9xsFpvZKJv74gLsBhGcXC0JVvphR/hzOiqPWohQcr4kPPMlD
ttB/LHUWJ0X0jlK3RlcNYU/BR3savEid3aMqTnxKwYajJPB5cyvJ6FFBOfZ0P5bt
X2jDWHjmepDlnf/WblZoO0Hyrle5p91Or9UadQD9X8TISzkS5n3arvjNqikJC40B
qSYB3T5Kz9TkPpB5LRkQQAnJvKScywHi90qFiL+yzdmE93TLcFGOsVsozOHa0MhE
DQwS34RfZlv8k8gqjuNMx9BUxBKE13t0x3n/SMR1fbpt8FfrOm/3mekQXHHqktH+
ALiVYVkX8wdOJKHYfMAYg4kjsfPI06RbaonnyJXWqERHvMRREjn0/9g6iBvM2i7K
iTJ8eMxK/anEq5F8CrD2Kq8bpDZsvlmpShXOnA2L0JBPSEoihoR3iI14u/kSvydH
TOlMcuh62KF5USk3jYRb1fLHtlXf1eoA1HquZb9ci6UqC86Z40JVBdMldaqVsR6V
8aWt0LHbk15mi86JzeKlHayhQoYtMbJwuWu/SKxhyVkRgZiMa1gonk2L0gPgSNpz
5+DzBIvKMG8BitwdyqEk/TOdRO1NZ4emsGic31W5GOmVHujiuxcSQSK+yM1bbqMC
DuNtTdQjvWyWnCAIMT5adM+tSyYazhUlD1HpXz51eG2QePGsz6eKfrvXDA1Wo1je
YDRnbP5cwp+QvGe6THTsB2lkB3ldxvAb2NohF1UlYWGKCE1B64C82JUaBtorAFVM
wVCFVuec1CXLRQsBW89XzHZ1u1bHuysBmSPa0H3T5S5Mkqqeu/Ui1Z5sXO8YkJKl
y3gSN5wbCnqbmmqZ/938OJpd+sTS4BZ6hqfuJK3io4PU/9NNuMBiz+PY9jrG5Fnc
pWbsBUIJwZB61Dr3Ue+xMzYfGEbESWNBDKAth4C5aC7DIQZs/dszAlN0IaOuLPgA
022m+Ckq0rBLRItqxW45/3GKw+c0nENjkdeQJT2bGoBSxtXh+b1Zei3R+UvkQPOj
pvPr+UerYq4WkUXGKakWHO1aO8kQwrqSXSxm9HxnVDziAUQVIQPwWBqIClTRodAH
T4ACp6J2uOZ4MrpBgaXBiiaOw2GUlfBIHCoPkEiRM2z9EFuYeKZzbzOKKQznP5CF
TN45fSFF+9h3vv06KWpzMCSuQ1rTC+JqFn/QNz4YRgFB/S6FP0F/qpjoauTcMgsV
ioOwua42V0X5WNUygtLTCftXTuuWi8H15P0hw4hm1yVhFrRJS7Q9wG7Ixy0nC4gU
NA/INFVsBswSCuqEZuscqb+XlIJJ3BrxOh7fUvdc8oHF043M0vf/MN15KSYopaj1
Chd0qPWUUv2Ia82mdtEiphBOaghYwdIBZh3ynET08ISnKDyl+qwXV44kyXGDRDdO
y9cxJAFc4NiznOVWsoR4TETIsTwcEmx6IdBhZXlI/wRGYKBaK9deUKUbhfJHzHUn
Vm0S8KxTJliGbTRSL0p7OSsfY8OAJXiYjPVGj0ACvE5bHfQsUPI50ndO/6EuNU+b
sCLhDqBsZpxQwBdAbo+MWz6KPK0+u5dIxKM6ACuU6ODFl6f2KSRxfzN4Af2DYpHJ
RmvzzQjSI038HRT6BHlCyp7mEiVkpuPQO44iQaxkRl09ajUAxAjqnVqUP+yRuGKr
DjOs+ySgZ6KUs9LEDrvV1auvK7QCncFCXtidQspsfzhKN8hhp5VWEQw950k/db+8
ZHCy1825a8XjSQO5XW+NqNntrKpvMa7Q1rcv6uFD9sNyxige6ZQ49sRrAhF9sHmx
y+qDdUpYIA8C5Nv7Zj/yXWfDTgOKDMn6wjcebVe6b8t4bub894C88rrmkpkFsT4i
P89jY9ImfQXJ3GWJR+u3eFKfw/QRvTgfCKekqRoE400seNNsLDH+15pC1LMF/nY3
PLrNlAxDKi6ypKsKJrkyt+S4XU2KyIq7aQMAsg5ZW9WALyi9vaX/QrTSDf4AZp5k
KSu6CrDiKAPnAOgyemj6/KgXcNibx6iMB+FDrTEd9X7wAEgVPx2QK/sCSUBK4RV0
PJs+lYUlP+UT6Zha7dyiYF/F5fbWsMhiNgK6YzgmqyiO7njezhfAOVRv55PsH7rw
hHT4TfnLn37vUN9tIjvuiL6bikzZoglhaIjJlFbaYTjDVfQ4AQpdHBqGTlLDGnaP
oT5X1ksAbWfmo4LP+eBeM2mpwWI6ZW0MdQUkJwegvHmWgSq6hzYnrDT/d885J5UW
Rh4h/zm+AL1ZILn7/K/hiFqFLCXR15mYRtg/Ryl3EbZO0E5rDJkHv4g63gyBrwhE
miVb16DSRfGHGddtCXScOwnZgpdGI5hL6XJNQnfaEtDitir9wEDBArx3+754b6wZ
x6dRBiCoqHAdN93iWOVWQKfx3KJkNh8PavGE4zBMVrwmEj4UP1qaiqw4FFAIesnh
tsaN2BpESFl/5Lb6o+uFiftWXQ6fe49+VZEGXalp/IMKWA1b8nzm3w3AjTuh3l0z
NAqGl8SEwJBzZE8vvSx6TXBoMcbOOjea2LfCsdVFan+T02YFLAG41Vg0vwcfCsaR
yi/zJH0Zj0pgkgpldChLZZclCn4e3r3cVA6cLWemPH3PQWIiD6kzP82zpk9I93GN
1B1dkqUdki00WhIKoRfm4boFKTgkvInEEN8Adyo3JNSJEs37ugO6rOpVA1AFQNke
VmpGhpqbCyMklTF0mHWnTr22r6Zbg6DQbMetUmuxnpR7V44L8AdHiXR6SeX5310h
uWzP0ryy8sWlCPGtpKZ1DCQTes2bIpD27fLUNBDC4HMpG/A9vF2dYv6lK6hwoYPQ
zqDTDFs9HdPz0gpwrZ049tSnP7i5IeUn8QMhz7PWbvgqrrZw9iWVCWk7Lgoi7WY2
DsCY7JEwvM3QgZHPomZAzZrQWP7KwhXnT+O5IEFPUn+YLe2NXyu3r1mzH7PasmCV
MPHIWBwwdO2mokbF/MBr9VZe4qdo3vWi+fAr26dGdgqrFqn3V454WOcaDzEgznNo
C9NnckyoAYnF7Py5ZSMCRNxWkgJSlltAzfO1lFBcV+8xyE5iUPja2GpstzKEOwSj
atzn/GUtutzM8+SsmESwEKtmLrnZwVO/69JkBWhV5An+TFIPCN4r4lIeOklgh++d
qjqeKpxRLJxiSeMcpE+l7MuOLCVma79otgd8gKk63NO1Eg3lP6tXvDFPT7y3u1mq
zUS3/6eQdnWPr4mwNsJpV+fC+TppGHWaNxXpivLlV5AmfTXJNp2iT7K9hYWAoCrA
g1ZZWsrQ+TvZooYPVcS0yR6vrDyriZ+LqZ2AKKj6YjyBdkco/F7rCYnJ7FPfHnY6
4xWU7C3AFo9ZUFFHqT1hr9ytjCURGc0Xba5VShoPUtxCPeArbNPJQMed1ncLieXm
jhnouQ0c9NkzDbSZ1ZkT3NIEaFZYsztKIFIJLcSgLFIURLW9KihT5p9mBJcVQ3cg
bZEJ1H01J673G776xxn7XfJO5BST3fVGquIXUIAM4lCCLB9RxIr7VXhhKDmrMUYN
4Sypuxk2dL4DOlBJ5bpKf0f2rs+psOhb9XIu3Btl4x72/oSUKPnjKn78N5GtC3Wv
5W1wCAfqeUQ/OaaRnF2Fysos6MtrilrFkI9lEiwDldmVrlWPAzgKyKyEhVuTY1ek
bHPFg965BiFGoh02AxYjnh6Bvz17NcT8KHWtkOHEmpFcarUfmDgjUqWW0vEN4zE0
nNiSId/5BA6pcH3qQ9n+4PNStpcObYm57X5PU1oaTGRxGrOJEoB86klvoefiUH4n
8PjqcCHFcunpoBKgUrkomPNmbdnJz9vDxCcPzeUxGRB7F/s3ZidrAcrRgz/mmrLy
lfNQ1Ga3YGM+xaSXdgT2mM7muGJfniay2UylcQdZ82tnC6FcWhGGoZQBgtj45pFm
ferAidexzAgo9wWfDdW4QmpjRInsL2T81386bw/GFx6j+WxZ4qFuWO0FE7KmcG6H
FJjJCcVqekxn2ryd8TIY/uAvJalmI1fNick/VsxNIkui/GfdjO38qK3ibd2nd1gs
2zjmZUEMx+Oa1aqoIEcEwdNwEyAZpB57X4ehPYa+Iwg3VJmij16q+cR1YrJiwp3K
TSiTwmXa3WX2PQLkO041HBWA7HuE+fOD85Fhy9q3V+USTB0+VHCoHgLlgsamcx6Z
SY9R0JdSzMJU1ULIpxbvFi9rF29RVYq9a2eBezm1NX7UrFKiPnLh6qsaUdFJgZGo
ZhRB1EHzePO9XaUK56teyPZOC76Bqddzt3PjFC9JplLqkuMdX8P97g67zqj6C6XM
pYA1XqteE62D51QijocEngBrCgSqrf+sI3nwZSQKxCDChIaWyGFdj4LS5ymDxCg1
Qaxa7JXgCvK7P7LFbx0wdkqsYKtSxN0M57XDoSdypxsv02DSWU/ySDAjkHFmYTfU
P+98Y40c+llE2Y8gEWsBCbwdzaD9bWISRD89vZB3kKIOz5W9pDpoM6gCBK1t10SQ
IpoSTAW3lZxVcNsI5q+HQMt3GNGlAhgDd3wpsCLVYoNV5Y4TsWjgjVJIbY8ivG0K
KQ+AyN9Ey0CLaYldkEJJBfdtXptae89wdyHA0zPqM0EgCko30xWy4hAhxw9HfMcx
fXfyZHgAvfIIbug8aCh5sb9nWExHwedaCSVbweTHmXTQTF9WDUssRai7L/y73yrj
/BaLIzNeU7AbbT8Lenrdzaf1ISZn+TqqFRvkdYUtpzqhhiR/YPaA6NURXIqM4pi/
cK5nmrKQstxkfJrc+5yc7tKi3F9CnbW6bQNZv4pNv++557o8u3KOAgJomw41/R//
udOIc7pt/k5amelmYvQmkFPMDt0irlkxTeAE048QN2PuZk7iyHggLV+ocq0ZTDeo
ZyAFiojO2lQISpqWdmnyYkAkWQfAwVwsc2zaHGVP0hLoNrWxzJQsU1FjzGMFh7HR
KxU2BJmtFe/7WV8isyb60W7C7RiimRDqixEs/NbCJ9sCILDM1BhkTH7Jl26ETbcF
3RbBdh4+zp1XBR2ZfUCfQryEbdE26+x1snT3NxoY5ZPYJQyJbA0VGLePCMQp2mk3
Q+jusSk1UmPB4n8F3JKfWFQX12s7k4DrJQe8drzzZ+DHInlsgrrrUAh0o8BlyM/c
BR1Fc7HFk/Cdf/sCwEAl/cRISlbiU3IUgiEC9qOzubfZKN5UNX/2VkhJ0saahwC2
XMiPPG2zuEF3jB8BSKhFyYjb5sWltwcgqQXEv8pjm5dP0f2G6KxQ4+x/4TMbl1uK
XUxOw3MpWs/O/qkvN4G7BZnRhfBntwWDRdc86fFAJ+2BJ07rJcrZy7nnn4E8CwVw
FOP6BP07EURr0Y++iKqgzDOqVyd3pmvh8+Q7uWVxdLyCptozLvXKH1AT21aJP+5/
KERel07QnKaPHEpIbRLUDdA5b5tSB9qYN5Mp50ArNW/kCqtpTHXDxOxUwv8ZOksd
dlttVkRHw9YKhiAWHMz+kyAYGBxyU0+UhEpzfzJTzR3m9eb7+MllXTF3svXsfWHM
cQoTmOVceJNUQYDUUi4gO8idE1bqEUivCgdmPQS2DUHDA6E2gvBGfgcHkG0/bypg
QoOKWyTwK4WLFurr2ldX3wFa8dx4bSsi/Qw1QWUNUghjSSV4Zv/ArDbaYCNl6XE9
zmj4y9vX69A4PFfHVeDvqwx1LMQbEkghJI4HaBvtQEyKiH3fJNmHkaWFW8FX6pG0
dbaG0rWUOAIr7Of6gsE8XMVpejKlg+aK8TJ2BubH8cfxfsiJ8k3mGLVmW0s9bRwu
ZVt+flj8WGCR7dKg8tUdWq3HCiKgpalAXEQItZrr83lnVJfMkBv/VNkxz7YsOJ15
ZxPbmiB8RdTYvx68rHLPsbuAEKIBrglclASE/rumSN2lFjKtZ5ybdCLnVX1klQmS
pTknsVh9q8Ix7augcTn/f0mXid/MDWrKbrUyZLjOlqU02SgFUh4DvV54cJyUtQe6
jzDbyVnQBrMzXSojX7Qh0S7TnNFWU4YO1ghzhaGZWxVkQDwoba9d+mp1tMubmLZ7
7h1jKQT64+wA1CkXK2K1YEYGY6k0hKGnZ3hKpwRCknRsDz/+8hPdl0G4luyk4mCE
IL+539k/QLRcmub+oV1vStM+xmq/1fSRqFe4FLClFdOdid3jvkVFnFKhesujsrj3
0RHhEW+MdrzmCtHZtCelajmJi0dDz2ESYfkm9IymnKGH8PCI1pUkLlbV1Nu9oW3q
IWLl4hAszYTvrhzB0Te4+6qyuyPOJkJY9LV3z/LNcxoz5+6JCHIKLKqxA96oWMbT
uYF4c3D/gzWj7nH+7Nn2wWiz/3DLMnE+QDr9QngNhIIjChdJkxrRBk/eCLgFNvG1
fwNOvEuW/qcR6UaPcoqZdO+3D8XYJr1OgDWF99C0PGxOZOPuul5xYMW+u/b964Jl
NTJdSeHOQXmA37zOJhkS2My6Rs0oyK3tU5DaL6MjBuMhI8vYaWQf4nUIXQ/ieSJm
4csLY+1j3Jce3Z1VipUe4kt1DCVuroxWoGB3zcYkyMQVe3YWwNG8g3ZZuyRDiJIO
PX097VpYRRLssmfXunLBMu2ZChbWlArF1oKaDdtX0ikZZy5BgRny9jDLbyQufnDR
S+USii6aoZtcqJhxJGkQCmqxZg6Ep8Sih2kz9p3laZt2wWWELQzvd4ehHtCUfSNl
7gWVCL6Wge5hDqT1SxnYMCa54aNbGY7slJ1KSOp7I3+ALkCijpcO4Y5+qjIsh+AU
54hDOwk/WM7wKODjqUDmcad+8/zYLNBdYONPGEvrpJNm8YI8IHluuiQu/W/qGmlh
JO3Bv/KwfuOyaFMzX68KMIcTr+OfeDN3KNyYaO8pyNsjIbA40mxRDBhbgslWPxFg
QKbZFL6oB1eF45aJAzL0Eq61jtjHkr6KYhf6ChHn6MeUKJxs9+spqnnYyZcSchTI
mCVQTITBgkizIzMd8PVYv9XJugYPSjRsfLMNOP/xg5HIiTaviC6lA4qZAyD/KebY
/7Jj0S0WAdWfX/VUVWkvH8J2PWRo1jykQrB3AiYuahfj931nbwrxpk779QiQOgHm
oH7t6OXFRaeDdxzTiKRrpBO6YIrs9ACM8s/FkTu7x+9R3x3a48g2P2EC/aPd/ZUN
CwO/gwdzoNQgB8IQrHPV2VgKeM5w2x7YbzQr0ziZrVCTzeMRwc3Tl89jkZNpBV+v
OSNeOcAULbMANo8S3NH618wNFFL+selR2xo04GyOGVf1g844MzaHAteaPaEm8S3c
QpTVEBfjytFLycRA5Fp1VGFn2M6UFv0lX8XihlxRckfJ5zvUP+g7i5UJaVGy9WBy
hzXHryl8ym5lNXODc+pbMrG5SuYcHVffNdBHdPgU2pFs/huF9oBamYs3i5+I0iz3
Lw4ueiJ8LZ0GNLk2mlpK+f1h+qxHmT3W8c8Ctsbf4d2ptNEwdH2tCIy6p+tli5hl
Sz7JAbI2iOh+Nzfk6KUuWujANfOVgL+y/0SPrNVDSmcbXFQ/z6f+JGmUz7nOa3gp
L5fk3BUw7LCod4tPmyULEvVYQ4mjS95LkW/efpuuCkhiEnVKdGZfplYyyn5x5wFu
D5M3ckvUudH9hKXkXJTEOHk90wKC9RwaKve1P6UK8RXZNBrz27Tt+RYyASLIT1Vp
ON3xpZSHUORTxCfDzY9BfHnYMi4tk+t36is7nN0LQtIhPq7SryPx+O7Mdt5mfBPp
yhNtXCUwBUMJLe2lAA3Xp8WFMG/YFr5/klQCnShiiGTGu8YxhMx0ot3nbZGCOAiW
nMbVpe3pAOwBAAc6/MDYzXRS+LmiW6MBQaWoIGYxoIyHHz3PvA1zm+1ZLYpmi2Nl
8ofHICXgt1p+5kXM5RaT43hCwnAeyRQ6RTlsJtobtO7LY45aZxcL61JceJccGGt4
TqcEs+3TM6SFxqOObtNZXJ7+BMXDAqtqbib7QNVjteXMi8fPHvVpbHPrCHJCYK/d
CCwEC3IntWgzVt7Mg3yZ5Pt5oQNN1ZolijZnc13Ze+e3ygWmv0jnNbvUasDiwUsO
TLE0vOS70m+2nCkCepxg4OsMbpqeA1eM6v4EFXmZaW+2IoujjHJb9Y1YG41FNiu0
3kyhpdkMR4jTEnQxw3QvmvlE0qxVvbT7SFwHrpLTcOwh+QptL3FPDwJHxdX3/VSH
Ew10eW3MM2r8rzj9QCzQD0EX8qAhndMUGDCPV6BfCq/ga/v34GZq/cKYewHSHocd
b7d17SPnDnflzVm85RltXyHtH4kgmMAz9sBOdj9kS7nSo3TVJl9VZFo1pD/ZXJWk
2Cz5UwbqypnLHG2TGlVvUP8391JP2NN3S48GcLpcmjcNu85QNP/nwY1saAMRznRZ
lfAWY871Pg6zHAVSo5fd31aB8ZgVFDg2sBRIHXBSGlSmEp8H5gIPYyxqZGKM5Tve
BhyRlnxV3qXJs0mYHfrMNDUbo/d38V6YpHAzUzgYV9s0cC7Yrw9pKeF66PfBe6Ex
XFMoqYozturhhvQOdkU5KM/b6VccwjgT5ciuLJVpyk4X3uT766M76gB8rAmMwjy4
Fly/PyXxWFiqfG9Vz/epxQ/HFgwo3LS8dpVN50O3UibVrIlChcIr8DjNcPQ/qSr0
70bEn0U+HsOs0ts1vGTtkTEDiFRZcXgFuzTy0FpJlSukOhpc2He2ydHBrlzV7oS8
8Lijjg6St86QBZzUEZvvlHwQI/q2zwf6iUEPvLfBP11w39DqmupeT2uN0viD5vRd
Dab6LTsaTGBW+O4l2boKGcESlIxRgB1ZHHPndesuLAa170dKmpNgJvrcOsuoe0xe
lSz5kMJ0GNZnm9KIbViSlyoqftlXvMa7NEBZqRQeKM/sLoyX2O058OF60BVbEiXA
oK3uM8N9MdJYsgezzusEOLlZUHDJFAOriOTU56vAcil4D9S4iH/EPujO1nL+YNu1
KZ+wQcgSFXz0Ss5a9BnZ0H5UWD/6EU6V3MBnnWo9Gxe9HLc5Zc4DS4TIpI8/OF4m
d+Yfbo/Qson4LJRU1HkbA172uJhKrWFVHJX4VkZdeYqlJtLb0WUjgI7UejwZraCJ
OL/xdsDQsBjUVf5WjmpsFrVZ602m60Q9U0UhKwd4NBUjjv/EvUklOB56zyfY1HwE
QlKpHnhdPOcvIDddTZB2CMc1M1BRiRQbgvxh4xTa48dFSQ9ChDWLj8pFDsuFT/CG
gjutGXpBGp+SieP9mGrIPlNocIGQSKorHzuYUjrJhubpagORmPPGKoZcLDOC6PGV
ttQa7017GMLQJmcJZBM7xMlKrPYRbuKp7a87+LVPPeZu4omL2wuQpXxhhn5c121C
gzqv0T1SFBrnKYk4ipaf7pdpLpBTs2+SI5SDbeY7iMGWHtd7ZQZ5eCEw5zYb+gPE
bCbCVBFVXAcwZTe0suMEx4t+umqZvfCItwLAGqE2lb6Qa0yRCCoEneC7H1r++Sce
bkWuiBUHVdFytXyd6HCsgIjzq71J8WpyrZX5fLAn4G7CrjMaf4DUAIDt+rjSB/zc
HRuMtJrSqXJjAVrGGZv3PMfRqI1EaMb9uhdo3LtupzOOJKLxYEE4Bw1d9ukfCshn
GpdMDmR+rGw68Y316P8duiC+mGqu1mrYeLzv3xFaFiX0D410145XjYyuV5usII0G
7nRV0Yo10Gi6fKH2hkmfhJtjdBH0cvRuEGmnZm80L/G5Bp2G0V3aDO9J8+wgt/cf
//gIb0raNpymX9CLFO0MrwVKKS/hnquxHFgkwl9zpgQTyx00WZHFgzkZv4BQrw5Y
i5E6bdgg4om8dDtJSCZvE4TPBuQ2XYj4SgHtb7lq5WOHsGwEetosKh4J1y4ZpJEM
n2laoVjbyINx/DqQgnSPENKB8sulGMFp+F6mWqEYMUYZTBTc92yNfCHRlkU9t+Uw
pBfCNQWXdmSuEWkHPy0L2xWcshEDPDYVCsu6vXP71C4hTahqODm0DkylNXw8dS8d
cYDaK5ZSb7JkTfWpEhUGzR6Lz5oXY1j9hYGeIvBoMrwzdl0K8KFNDJh9NJv5+OXk
w0pXwO3oE9inwtkGdNgSuxZYvB/MhdcCMYOVjNuzp/wEqD/49VI7zezfkE+RaQ2C
vBrfvEpAKk7AW3YM5IAv9ILhEUrfkEueY/iIm9dqNPoyEvl9L7rxFxQMzPjdA+3o
PyKSsAoi0gmsOkvPqhvQgq6qo0KYiEF2IEuRFdeEFXdTrrnqiQ5VMFGCo9fyvQcb
+ixuYJIMn/SWklqCvX7q6U+Ba6xQG/jdzw394SoTg8wvC5Ck75Qz/HyGqPdnKjkn
w8TwSea5R2D7I4PLx9UUNkAlTZl3+xiQOvX5JmW6AX+Twy5xnGeE3iw7zenO4M68
90/sRBBim148QPLkj1dBpOcXUEL1P8GTBRXzVr4OLXNTjfhEXTXlhRaQgDdsI/wq
hm1+tDFJ76X31nDilMxeUo7oLqq20jWOv7efey31dQPtKm1TXZ6AxLCv7YnbJVXG
JpVmJSUExeocxeTemua2QUVoMfuRU8IOdVnAmrrhxyqSe2slHrf9TnPA0YJa9oRH
V8OjbTFbyyVAFnTCkVnmF93MQMf0ZLZiANVdPmWmB66qHQEEVx5TQqkpZaH6Ep2D
vvUUZz7p6iaSPO8RuQgrt4QRDQhquKY62PxjdcYzSPzQGzyFztxPxvajkjbEJJZe
IZ8tohdtq9MA9aRA+xnmbYHXEYfjduk4hxjZg4bGJaZRwj2IiTjq/GRr9iGbmbbU
xsa9gQ39pjrJZIyfOwL6QD7q0QyuBUDg5G7f7Z9F7BZEC4e6KTBOWr1DNRij7923
8ax8WBN1IZ2BhZoTf/YE/5kRCtEYpZ6XCwv6kuSyczS9TO078IDflNSqLOBDvr4Z
QiDnsjOjDVD0A251eBj7CUjP+GsgjUHY5qD7Nvgpy2tHy7lYibL3z4umfQ+Wrv9E
MuAOSroVxpHMRRi4fnWvQuzX/zssntWRRPz0AeR5FN7ETs13G9b6WKXKb7bMoBBs
j2VI5ZQpRWTEyGzf19aW25aMhdkb5/0PspgahcwJr1gQzBwgY8P7sDqMcGSIEUvf
zNNmnahYgNx7h1gC1HErXRGf5R66a5Ri+imBuewgsnpIo+O6poLak0hge8sBnsIn
BOEsf3EY/kBOxEVxa2mg/9FKlLMuy1ZcXaqj5TDiql3hmAEdG+INe2jqF1qGHo1A
XhgUmviAyUnh+fQeD2DS3jk3AZVMO3HkKuCntnd/D1WOFN/BJwIvkxvJWgyL+TNp
/90J3zWb9rTXvoN1uqy6apoQeNPH1aJbB+ckLsFsbIkKW1+b42ppLmg4E7uRXhc8
EIHb7s/aIYoQ76mANBSXFmxECor2KVPnnCch4bytSfF/aKxgXLLg8KR/UNIBkG9Q
0sPVfSkHxNYQE/ZRGEOOEZcjhgLwylT98jTGa+wsLxd+YPh4HqekNPckfeY1vEBn
hnmjCNP5pa1vHP9mjpL9QD8pgBYmQCoKbacZrIR9earWTpCADM83FcKSrm3+r9RX
/Nb1KmDY3/ONp+zHbZkkpZCdHYBTBtf7It6ZxQ5tXRg237gGmlbB7A81kF+Y9XrK
3cH77ifjjntjhnnOa30JseiHvdvUb392bZLjzodk7qvrlAwFjkbRq80lIA18XKBO
xysrhaTaKxkLSkH//FAELUntPIhv3NSJH6x+IAeAlddTuSPp5Mq89eDckJrYn3Ou
WkCz12ul1o3EmpcesN8jQOKSE9tHoqJD3h/TBTcmrt4vYNFpNoAS5Vnv+ovVbpQU
0WeMfq18GIOKAO+2azrZi5nootoxrRK6sWNMppXQNHNS3dxpm7D7/S3EO+N/qtiB
7CcVvhv4QIf7VoW+9N7q5O6mqlJQb/AhPLpxjU9RVgflUu675nnY5k5ToAbLCQ6n
IK4TzhhRkn66k3XquQPF3K37bTHj17vQTnTRD8GLWHP03IMP2T40kIrPNYseMtrB
SOr8QmQzSkRKv1xXJTzRRQfkKD3871ZaebAwOJEA25cX0oNVjkFTdwyD0fs2VsuZ
HeLAkswEqkIzcyfGw/ISnWR38EyMyWSr/+/WXTM6PoK4ghnsoUUP/mz2FiOsZfXl
nlENAcPVlKV7buqq4vq4s5OT5+YpBeyWoV/9a72qdEEoTiVwwIrCgKpBRDeJY9Wd
fnSQ9eh41hp4mjc745SkUZKqNtFjsXy6Q/d92Pyw1+wS7UPJAp16E5PONVR9o0ab
+P6BgWQ546/J7u4/rRb4xhRV/Yv2vs3KeRUP3lGhpOwS0KK7EwQo6LF9LCa9Gn5m
8U37YJnY/WL35wTZgSr2YjEOKQUnGQMcQjdRQrFuJcFiZHqA1+xNXSIoGvHCbR63
088Bw6Omdwr1fddt7WCfkEZb6j/Rgzvcfv9ejP+acvB9zWUfiJ1pFKH7hu4isSRB
y082Te2tCIYcRDRy3dMfx3DHr30yvvHMNZu26UREpKjb17Wd9SgkopvPVt0t5PvB
NyHabInF0vzJ8H6zexR/3sad6fy8ViWyALQepIbJGZFtAe9Yx3aDmWWqoYZ9vtwN
MSyTmcOYFuvzrmDtNIGZ8f8CNQqdT77jUoUKRCM83Czn3Wae/rarjxS4HrSgAHkP
6L/CaLRuHNyXjRkUwfWSgX4WrleM+3XplBqtiIDrB1SW3chGrQjSVgKiQ9nRyszH
yM0ptz0D4hirLhJBdaMll9NFBy8zHCcgA6SBPNi1kyrXrMr3r8YFwlt2qqsl2gGo
aLSKDtlPKW0ffukk183ddVjl+E+voUY5UAHodT5PF18FPjamDXkuDGLHH6TUMsBZ
6h0PsQxG8f/05iFFVw3nYEwRaI7GARuz4AGRigHzGjvUoYhETh5HjKoJ0gXEdebg
Z895zAm5qOBxe6MmCxTyMmiatWidVv1lsQSiphZF1px8WPPYkTItS0s14mPz+E6A
iBHnQFfYNCfCZsMJSWTCvc+Xb2dpLY4cTTguJOdDAXYAzlm4ku4NzPz3qlzddq7l
FJyVm9SBE3aaZMY4Zv2IchYOtLrOFMAw85vjo56mBbkMWBAm4s4QAq/QNSHETFW/
HuzedpPY4an+LxUvOQMFKkXGfzgpFZF7rs/mrTQXjTa7ZhyIYTnt/e4HH+bZnXDX
eVSMKIW8JjH+m4h5t3a9SJP0P+7NnMaP6UQ62xrjqIx0bqL9LsVPvKiTWOYyTIu2
UR1CzadyG+NqsqvtLQzTxaetQb6q703R3sg0KvhNpJO4ndRzxL2Hp2iEUcybS+AM
zCcmID8coQoLgj3aYmHShiYyVaSy29LZj67E/6mG1yp5t8Vcr6rdIpSZ2KiavjpF
znihYTbe0OcFxZoVVIc6aCEypDYWWmfgLvC3wZj3kewdbS4kqE9/6txnlxdy7Ok9
ByIfeUoh+kSwAWZn8BhOHfS6R7T0k3PwD/agkSRzwQY/61K9bXf6V4O2xHu2snes
xe94nqLRJ+rnI5Z1NG9XWBLO3KGsZE5xblG1xm/4yk324ok3zeeHznnbTqI0NHNE
m1T94U8eZ6t3a5+0Z8PJqC32LHK5qVwu32bPPHdUPKef/avcc79+83r3IcBh0u4T
Y6XybL+UTq+kFgnAOrwoAhl6hit6rjxg14V4/GYvRVpWQm60YZehYmL1U2lLeLO3
mjkg2Wj8Fa9ZAzqBBjnSnmi1dO+pYb8EQWaihZnNq9Ixgn5gOcWPBb6/vi/Q9zbJ
h1EYHmjAwVPGu7NkH6uGSkwhodJLITnZSKPGqPYoKpFAX5tltcQ48IeAAkCeYBt6
FbkQCnpG/c2lPWaUIWn7ipCb6lcQ4N/pVlc8eDaQuxj7MFUrs1VFrk4PdENe6u/Q
fA+GHO+dr90VFBF0/8LigmzPIZ5rTIj4RXmq1ulPMtLLhMwzUx7rE4ZJSXq+x58i
npZcxxcnOay45QarNugRSZvSVznYkR/4fS36ggrAzGk0RAOGaoIUoy1Dx0isrexW
RGDSWaU09Xua4+ofuPSBqONYWXxJ3w8ZqHFiLB+qQ41WdLmaI2sqfQsYy9tu/o6G
164Rx7twU5e1svAXYy9JjDDaUA9fEMOG+/Sb/ZmSe2d48q/1IiKn/mupTV5gbREA
vMB6ptP/mMSzBJB1D58GEsKjJ89fSfAW/jNSmVFoawccrszmSH/EmJ5OmEIJaatO
W/uRkrfk1PM+Sp1OfXuqY6KyaCAwLCOpPkcqF0ajJZXz0y5pLctFc38mXHDv2P+B
SRFrB7HPkdLSu/rhZvBBSFxLcNprB9vfLrjO2lWmRRtEqze0OPmVBU2Kc90DcvAX
l+P2gK3KOOGywQ90bVhfZ50fL4D/2YMe256HNtLSsD/E46VjEeqzQGR659TH26wA
lTETNB9jUwVFhI9vzoglytT8tKdEFFc93ZdIvcpksV/GRIGGZbjH+/16mlUeJT9J
5DqYXjGGCKUZEh35vusuX3hZHdHmHt++Dli7xYwbX/ro0oS9YJeI/RVSPys++rq4
7HKMcpvkR2tcQ3ZGk7IB4pAV4PTzaD/6Jj0V9XgRDGdZKhJuf9Kk0yZ77Z8UPJkC
EvdO91+5QjJyh+twuZDNCtL+zynB6bf7iq4NNHHQekst2TnKIm9bXBWp2T0SAkVn
hlalMiVJ1WAuojfMevq/dIazg1QKL3qq3IZGDkdy9lDke00DDSugO049+r9bMbTw
4FH/5/O4Gu63AoN2uYy2h8jpf1OyuXJLk8b334nYqDJ5pX9rZEeroGCC2VpCvuPb
1Z1B3Ns5d7HUvuguYglsKkfQU4HAz7FfVQrmsNQQN1qE6x4o//eZD8mwz1ZxFkyt
rJgw2rRCklrmw4mnfsDMeyTdBrH8MkCWcbrdhQlTDEls3RGI0hNpCHCCykOETh3I
+0EknusPDFFmwvApDAmEN13nT5F7K2lMhKJ40+Ekfq1QLXI345QoixlcC5nltzqT
6E4aRGkgcfzetDGft7MOZDFD/aq+s3yKP/4gBBlcudbYPohGmrUtkFiNOEvX3aID
8q9CkWyiRVj0bwDJ0Ybjxu1VB1DiJSEvJ5aS8CwS72RcCns2fdxYO+sBBVDJETjQ
UDf/tfRmExDuq8zh5pkAHwKMedbsq8UVruKZlAPpi8qE5orGVq3rEdkjY6TsGDk6
tWIs3zdi0Zki7hw+xAcvDS4/TSRTc3tTBNBBOK5uXb3v4jNjtyVX5pTYX2crlAlK
IlHJCYH+F/wzFTrfmYMCGv0zyqCVunTpX04DgeFrS8P0ES8iJN0mJ9N0SzmNOImc
OZSE6x1X7eemIiWqyK8G4vB9U3qM+MGTtRZyIPGQsnO6/vYkI/I3QRSI3K2X1Ncf
0yeFQOUymtL8ovN7An2Wmy/ek8rSW1TRX90oCClOg0NxRBUiFKt1XlY1A+spN8dz
9Koevrr4KJ4SrbavJh39z3Dod04lf8CKYdTFHLw7r8eim5rvXHNWEvCWewfthH1g
/KThMxPbep8uJroxmJOF5OrXyp7DLV8tnoFibsfGZtpbCyBj0qaRymFMyeExqdjG
M36dohuh+xYpeLdViZmvGD67d26QyRoupKghOJUwWVmhFnRTbOjeG6rbtENcz1p4
Zse/i5DdAbfS6Vmbx1MQ4ymjfmW2AzfcQiIhEdAsB+WJsb19nr783WL2dYpYK4We
wph3ihNOjuhDA6mcL6OySsQpK+GIYOak4tyCmc/f6kncXnuCfXupqWqJrS5iCRoa
4rxK/r1xnSVOLgpYUX9gn0QMEprIVVBouaDaiWtuZ9yYJNqQke7n9QmlpnhiDbQm
4T3PR4b9NVvrU9qVVW8dS5TPK2fbLq9TJlzBw8GqRUPCqGoMEzo3gyXC98sxifZH
U+3KZNusHQAdehFvT9aWo734AuGsST0mjsCHEoqIJQmkJTKzIlFWLki0efr1JbCA
wUUiri4Fs0fdJqrK4TXZ63Te5WDHI53NjFmGGqI3c5hWrKslGLvM9LoNa+I84wIe
p72E263iKLc8kHjpAb+ly3arWJg+ux8sG4+2Li7m76mFqNBOqmIPJPZUztGsw9U5
1901vo+ubWLaG6JZbmEWkh/Z51UgjZhAeqmxpy6u5s8ekB95uir6JSUBACIi8sFU
lES2qD8SiDCJsuFCaNf/7Nfl2geWL8EKnuhAb5dJMarjfZ6sZu8wnmgtROY5pM+Q
zLZ1siemslRCdBiIFQpx8mmJd/hStQRXzGXnV17kvNkNX4ld4axGRTSBO2Wudixa
umuCu0tDD/NMtC7+kAAdL6qIgMJhk0pD15h1I6GdzMfpkH2If8gDFE4NQFrwK567
yu6K37O+ov/WH9cxgVaZDdeE9IXPrPzpuhveCB/hJRxcaWCmeupxfTaBpAKac0zJ
FoFFJxdE0+5fjvR3RDofNiHNREm1sChRdQ5Hgeliu4Vr/viawGp54aPHTu/7VFyr
qWC1vf/OKHpEncRKo9qY3fqp68Fj+4vGm5Xbwpinw9zdxqP6wTD7pmyXIuvCXS3+
Qy7w71ITHQ8ib1M24tWudWHV+tS+YTTXi8bEXBHWvsqtj4osUb1L/4h+AMluZ5bC
twVSs577FhjxFOyuXBgYVwInZv8oU5+U4vb5pDylUgXs0RpSXmfsSw6fG6gbps5K
9efDA2wcBNpEyFEkMO+hXW0F2Kq/LqNnEWEn4evzW9Uiip3IQ4BhqkOqMBB0MRJH
gq9Ier7uOeRt6OvW5WnItLREyn3FmxV1Ahcyw51Fho3gHTbuTgMTrS3HtYvyI/6W
WdmAXMKL9/rrjPEPWi7J8GNDhg94RDM7uDy5septjzoHAOEt3IghBUtA9c2E0EQ6
Wo4QQMTBcLSV1dnqffX/xM+PDh/JMr9CY2Cr4Lwcj2wRdrV4iEaNG1FjeYnTnmYC
qduRto4sfAr0s3NNTnnDNTVnAznExiuyDg4uqOJWAOX1cmYENy8pfyPg7az1+g1K
JgIZCLip2taFy6N58lzeSta1Xpn58hqLB+m1XP1YolLCWv/m/py5IDJVZi4DqFSk
vYuRL6bnqdAbwuU0eG+zqC+2qBMIntbjS8JlsEz8SfvkeigH90gvCckNhfHeZ6p1
5eNimJl/zan2gkiXhISdhc+Rcsr8IBRoQVd6wUB/zLdpZkrvQCm4/dqXwP1o9yas
nDnR20nrsA8cPewI8GdMnBpNw4gm+Mj07KLmU2SeAcN9EFv7G61N0GVLh3f7zYrz
Hf5BpnT/NI4fQwPr5CrOhjIHhh8TwnmOxWXI5v0rd1vcq63bmj52ar/LjOUm5exv
ZJhiXUbprGsQic/fYJkjvhVHidzQlzXjmZp1srK2sOuWqkZs56xaenV2wdwYT4sk
BotB+GxDt2nvAVO8Ekj9itYKv6MdvV3Yc7cCsQxjCOgdPZcBnNNmzlje9U74H4qy
/pQiNHlNqomqbljrNPkRf1ujSitWA9FjD7kHmoNMFX4tfctfybxn+Fn1DimlEPyH
qw0yMv1VsNyFjxvK/ABuxOT6GS4z0gvIn472gdlLSac0ER7VW84VGXvrhJcn8KCW
vVb2Ts/tTuNuGbYQT+xkSe0t4JiUU/fDOoCdUnSSpaLnfMzq81efIJ6CV4Kld4S3
sYlIjn0qA6L3geZEW7h5Qb095GdswzMByLmJNkWmh+0sSCCbOj9WG4DdDiSJvmi0
B1ehvACHDrSjQnAHN8O5ASm91ugge4xW76+QKYFY9LUWOIXUove9hGYIcteLL74n
3KGgnODXtKWlA50U4XdQLGDa8LixmLDMR5ermfaJ7xCkWa1ENq0nCGB6r3Pm4prp
BJUg3QHyq0soPu+Pv+a7pSWm0bOGliYiCa2UuV87aEDDCioeQZhxe9v8QgBJbgjF
iVA2lPXjAYyDeOUD4E50GnZp+KcnocmeJf8q8DZT0BoGIfVSHZjPViD/p8lufJzN
SqthZQdao3wW3336G8RBmx9UV+M94Ut9I6B5MqpL7wXAT9jAyg5GgktAz5oHkBKm
EKwG1Z+Ka/mQQmhkbD54mQ/bV/bbjBf1gQvHn1BizHpw6ySPN2wN46/HFRjhdfCa
4SCG+3yX2hpWd9tzfIQe75NEH314Nup87f8Bp/OuC0zEAWrgYLQ5Pk/IyLzglhvQ
Ul+k0GmVtsm69zozvW+UtDcuFMC+cOfTqKIXPJnCZGZivfKpwI6JVaQ48D5OPv4o
kowSKXNpP2+Zi79RDN6WpK8oZo66V7Hq7eEAxRcqp7JvQ+WeOwVhUMmpF4mEPFCd
NFw4ma7JYAuchaHZ4SCukNxSrOJwkdwE1eCM5NvuHtnIyll/4c6qzZy+44KkhrLC
siH+W3GgGB6Zp6ae/WvAByiT4AXw/1mLbqYOuZiMjOG4MdrRYN5tMT/mRDGAASzH
KSqzH+pZwgCwfjXJWrtub1im6c8e5zln4mj7PeH2inaTbq9klB2ksDe3wovUkhiz
ZzLzFY95fToETpwPP19xbYcfN79DzHJDMftEoHxm8I2KnKf5vWPQ916n4HGfhW1h
317/WRrczC5SAX5sBNbuESfFNzp839VeGYAr26pXkgr8OciqC6WsUcCCMFhfBplz
0bsBWhbnSV8yfeT8qptoaTylLZ9OVdoEPBJ+gsMTocMAFLe/cvc+wsp9NN38CO08
QJpfenHMRMXoGuXRGvNJlGP9bqSQb1iWdxd4x9qgnlp80kEwzxITQQbbMymBGIxc
VAYsZZsDhr0ifopSGdM6C7JBiVYEUFA7mJpKmAEhMa/gB+TFiqf9aIxWB8i6BsyL
vYfGzQ2iRTaBMc+MP1obCuXEG8nNX3J7m9wUX07lgHeExyPBmOIUMPbmmo5RdowV
KLEgKNQq9m+dcKCgZ/eerYlsYpDvIJzH1phfY6TF5L7RuTNRvFvooGcVHQH3fmC9
z3/Q6J66PnfJKGDReWcPq4aN1bP7ICBcGIMb8ed0Pf3xA9cv84WuimTMYBhNV+n4
5iw520UojSPs+6P/Cg839J9WYgZzOAooLah6Mf7llpKGEXs4zGznzlJVYxy4hVrz
8tX8Jr90lbemhc4kYhRn7TE+YtGA9jXJ+PF0HCFpZz+DuuRv9tyX7Evgp6Y+/eiD
9VIO2/zUwRkcdgII53eOLehavmyUfhUya/OcKLdME9yfauZ98GmR3s+pLRFxOkcN
iFEK453tVv6DkK8FhS0ecSPZRmVa/nokmV3lpgPP7kW/ToS0tlG19b6bU8bwMZ76
ysclDRY0evUS8zf+UKkF5kEZorHrV/6djO12bFL0O85CD0CCKKQZmpxsSWndPb7w
UjVUWDEbzFqUj/Zr/+rwhzBZ3fIgN7A2s3ue8sfFt6NrbZkeQiZNZMdkZQrc5WQq
LBBhlZsAOxAH0dfDNMDZh7WxsL9D6TAw+4ZDtS7R2n4RfvCDQJUkm4TCVbn9RFSt
6Z+j/kXfHjqibdiGZEH9BR84Ev8l5sdsi2rY79BuNe3xc/ejOwyr+rNgNflaG4yr
+lWN1mub9A0ln0bKyT6naXlR4yXhMG2ZtvCIPZ3nhAmfObzouuWdv9LGWi3228Zw
b2yXK8ySMgNO16N9kHqI0G86H+agtrPAYXEai9Ji+UeG55RYaSfasiOLiaxBdjv4
oKZJELmtqeOtOr1mx4cSm5GUVgh4Q2EdFj137amHJ/64NEIbSI1y5Bt31SoJAkPv
6htPVkyAkFZ74WAP24EbHwamU58kSj4UdEQtC277LAxUB/uBLzX1iZnmDWay+9Fy
sEyX+Ii7jPsZim0sFpRW/VMNUPWqDbFv4/K8DjylplxofLwlTGPM2YUMHUQRFNRr
rifdtVr9rNpipvl3k3Az8PcBaazXlPyBUgdAtVYnS+L8JJYRLN45eueMJ+nIiSjo
mWVBV6NGcPV6rdlmDZNiPjBuvFt8uNca7v0lJD7nt5pFypkBqaPgVMu2a/CvGV9B
juq2Q6T1iGTdG9RCNuI98hjv1a3V7lmH9d279vUwG4kjAjRbQCmArlcItm6CgWhq
nlQABJF8UCfwzc95F3yed5eU5nf/E42y94uZXv1aEWs8id2rEzcKb+5nwXIa1Z8y
n7iq3/kiS8EdnznqikRGypnDu4jG4x7MqguDZB2CpYyXiMM7VnBexDE/+CblYClq
UMKeqfJQrR0kuTmk/xMPnoj4SmNAfb1IIMvd5LGs3SOyiAQI4lSJnom/nZNQeI/T
kBgPQrRQc9lGx8YGQMuXR8UqbHfbvzcOZZJlJ7w+WonRR2u7hBmxGZC8N/wSj1kE
UvO00ZXnZLXZHJBU3kQupXdhFUhMb6GifdfjlHvOydX7XDwERFg2ixQsZLxQ2dMj
nhGjG6ltdZYmKGepGnLsTYrWdNcdlru6Mei5q7QlHw57vKdICVglakJXjxG9vsfY
h59tjjIwZsMlkEL8etm2QYugtfuOM716exnD42LdWwKfLXq7gOeOxAB1SNT6+cn+
jK7jQ4X3YZCeJnrNuAYufnRVVnOU6mbgN4hIw/N03k9meBxU4KDkELo9cbr3rG0B
0F4PEmL2OFGHh0wsziIJv0+dRaBu/vg29DC85hI9lfKa59Z1zytovcU6Lc+oitTN
zt653LFM+04pD7i1YIdffYn2/eO7ptU5z8SOTt6kzhTTGbI26zLlCdzt5qEUtkIz
SmzAAbblh7+WkpN8LkJHL77H4OoiISVA+kuI6+F0lEj/5jZrHXjBAHX++j5RNJMJ
FtEaXTZpOCLPpiSB6al9kWy9KpOIZ40RxRvyESzhSsHMO8fxu+PI5sWsDdQLteAH
92bhzZRn3bMMPF3XxQ0BlZw/8D+eSORRrJKfkk9L6i4r6gYTU005K6UfXJ/FDwPA
4OXxRsVuE0ZItcl6tnLVrOktV3d1UbzkNKqwAQVBjk7egaQdY920xzLu7Wdv8Hae
x//lqeBn/JC8gJzUtWYJAjENBEcOH4CRkHVBEibcE12+VWTimN+WZIRgjAmQpYRY
xfkUYmynrTI2RyytED8Ak1QY/Oe8gQyyyqOcDfc5wpks0yVzdYf4odunG+f6DdyP
wkuMCKwstmIKTpSySXl355bHSpyGlCx5KcZ5+xfSD2XCm2unWRuRxIb4Fd1Cq3I9
y4XS7TDvJ71LmPYECTo2x2Ow60ZaC9GCiwLg5jVgdhyK+edi+M2+E44P/9pfZc/8
a0K0vIyP/d451fFObT3bpZ7OZc8/xnXvEM29mVFG2/srJL2NpbW5bXnJHpVjUabE
uUw4tvlSZOM7tda/6uWgye9oNR+AiuEk+yDy2Sh2sWzwelpEUOuePCvDxkefAyDp
FS1TbADYTnPsWVD3qDIVA4vbri22m5qBc1vgKdVZZITO59TlvYxwfKBrb0fyu+8c
2u2GyPUaQIBKNptI9vdnVp+GukMM+pZ3uYc2aJFLKvUc7KJyXQCBbeWr8bAIjq65
HLC9/oLcnbFJJWUken2XDyP7OYxDkGrNVuadbLz5oPxUi76wrHILxz8jzzX0crVL
70oSpyvMesvBPoqo8CeYKW9gI8Fy2W4k2wrHlhN92gzGmEiQj9tSjslybjbul+KV
lTivNwzJI7hR41lAVl9U2WJKxLcozTOUDbJ5M2ayRaiK0J1P278Z8RJRzFymtrYV
XLmpvbJAOrP7NCz27bK5sOUqT8Ne8yzYWsWAU+LCTUpcQbmROEIUZVWZakoz/f0e
lC6UXGGnBEWqQF/nFZYR5PuNy17J5wmtUQBmO83Pdeq4BKBPFDo+Ow6KOlQRTNVL
OjgdsU4ft25AgRd3tYAJK/oGZvv8Um37CmN5IGhHWCyr7v6LCdjnSGmbAqGcacjz
lC+cduJvGd1Xvjbj+k1i6eWbj4dEr8gLEPb2RMhpudfQBGWnT68chnPyT3tahTD2
OoEU8MnCVrcMNI2Lr6XIYfKYIR6v9I0pBk5tYWSTS0Z8CNp3SVFcgDRXsz7vTKUW
VOKl16FwyLilJFQa+DGJG9Zyla1pqRPtuCDPaqa9HpKM5RsOWIYWmwOccYMU1u/O
WOiGF/6WysyY2KQHQN7JwPuyFMtqyCYw8UWfnrmIDvXCGUMSfBOkiC06E0ljtFR/
G5eTIDn7gMq6Xnp+GxxEy72T+B5Igi+Rroaiy9WRmJNXzMnrxU8QfxEbQFArjeRq
OnOGexxpci6p+Yj7eNaQR2lcsWHJNX8dGZbXAknsjtO2f8uatRghOKjrmaFh6w97
83r/qPG/cIzm4HGvDTr6Sh2aZ5931+q7WYpWF7V0kvOt8DAJ4nGvK0In7OeqwWC0
tYpJBZeaq8OriPn67zi1z2zfGDXJcwFAHSUiqB6OizolYqRtifskD6tB+GclN/sc
vx56s7n0WmTF9SXn0MrPSt1FcJrc+pWfpYIuQlqCs5660nAIkm+5/EOVY+hIhhBg
rVTkaf4Vke9cukcHT3tXJ6U28WW1q0Rz5MPga/sMRJgGN8ppaLfD8aJIhF4kc0jI
kxmbwz94CPyUfj7ccP+i04K8sUARbrFG2qXMnTO7BphC+eAhKzXDQIxGVMalswYm
TZiMpzw7AdAteeqjWO4te8JHBdQi4YmEEkmKMFBHztYhM1qy6tdCuFi+a5MTo/7v
ZjIyZ4Ocf3QBUtB3HBAHF3Uri6/jAmG50urqbZbDinnNeMYl2dwcM3u0SDK1R+Ny
kD6pJqP7lIUezrQo6ki3zAqtbmFrr1tnzV4PURWcPL/q0CgpLU/DidpBaD+vQzo6
VDRNE37DlSeBAf7bc8uI9mocubRfzKTjsF2ZIw5s1EDsI+I4euak+nIqSgFpt4nI
Iau0rQ4lwex2Tv/XPxS5rehri1QqsM3coSvsFtii2LGgkpHHBtU6i5wA7vDG5XUr
FzNyaZkvsofWQ13MJOon9G+FoIGoSAPsIjIqcCJGjDExyl9DoFmmfE2l2PDhReYe
0hO7qMjVLvUBOsNQpr/xfXKSuvFvs7TCaCqD8knfCRn9+1Z2aUnPS2ywieqhd9JK
hWJnMu2j1A+LX1yLX7yeY3PbFgwLukFr0VeBStKV36SD090GhcvaRxKDexY9gcRM
FwsWk/pxgub+QchAhtGpYOge+m2wii8LCZxJkQq1foydgLiDpJ8ehbR9DweRC9lv
ER4kTbizONpRN/m7ruelmbl4pOq+2d2FI8R481azXTjaahnJiN4GdUH6lCDBwz0b
8yPcngA4paDr9F5UdpQQ5i09ar33eqxrNI7w9kkyfPXsYTF+NOWzQAnPKAPMim9z
Mzf/jPEI3VXEPYZSoBSjFJG0DxDO3UQJW/d74IptYVTe/tLbVOtDu7inNYIc3kCK
OhzclYqcjPeMYUFTvFFLjot4lue7Vn2pB0olIogS7XHbXUoHgmiKZTc0Ot7fo5mj
m6qhD8yj4LSBGn52kw8t+RLiJ1BAGtzq+Fn/kRURuqrM6aOTx2Sb99jBic0zDZb3
BMft9QZ6tW3GfbqiSQH2xLbwKFKA6Sha0iUggD8KtQ7CjiEZfji9XHyudCuUc/Eg
AUavMvFtXY+cg19WQPNguFk6DEdqjctxfAEHoNFTnUCql/Qe16LEW+0HGhpFbuAz
ncpCtNuWgsrqFq73E8bZ6f3M/z1oXWoUOf1UQlsVsrEeeCtTnwJkGHOlDOAkUHyT
dK0sBwxxoz64dnKGrqP9BUDauZhheX37KN0FfTBNdLzw+mYPE/6dhXO7sypV0n3y
Xg/MCdncQnppmUWnmXIXqT+PsccrUvTqZOUqRAgqEkRhmdB/1M6Gfm+CPHlkCRpi
D5uOdm/76dmVrcboxKXpnzpFufHglsfgUplzFq3sWa/qq0nrPv2i6l0ZiGitoCOQ
MpbwcB9TbLa2VPlOblsSHfKneNowuSdLIzb1JPSU5WhEV42HUgFJTpyqyNwuU/fK
jahMdiz5GKEqC7MnhM9OZq20FVcGcSHDaZ22tv3jV4SpbJqwsbWttjyiCTf0HX6P
/QHJIwKwMcAKDmcAGKotcRMnAC9wY+3+FJot2WT9lNNxjrMF4nWi+wcm6w3IImY1
r2FZbufSSYBiRXCQCGEzjRi2RloVaBfRn1vfNI8WQ5nXmHbk3vuQ9fmica/001XH
gnwWIHnM/aYquj4SUK9uUCsO5tKIAyXdGgsU2OMgLTcfa52Pjt3ooC70NSUZEmcW
4L98J9PNMOVit4uLqgFYVW5HVWYgK+TLoU4+NDW+9QeVd0EeNVg1mxd3pElsL9YY
XUWi3RqoaRgTXak1YVRdIIJsHDmBYFnNtjRNg9rga4z5yKbAxUKMWSV53GxBqomf
Nka6o876muvd68vsCZ7Q1InRGBHHdpxu+pHPUtBGYzgnjgXFBPgZVkSz1Ho7LWaG
PrjNBHXSRE2ypN1agAlFer7QamAu67lOYxtBsCFmgMUl9XB6xvPF68eCDT/A5RW6
7qSk1N3KG+f6biTUXFI6DNPmeRrp2gaKd9YSsQU/TFryl9EatF0DmPlJ6ua39Hlm
5HG/B132cFPVgjneCrJNNKY4/CRyLBjlrH8Gy+MhQQeE8Mh0j2jO12UoCxfsgcs8
o8my06yhB0SqCJb2fMmqCkeuL9/2Kd78XxZhHkwAjzSsRVtMdg5VCxUIX2aRXApJ
No1sft4ldqUtYHKkqzOjVO4tzBkdp34jBJw/D6irBqhutYmZnL60dqLLcqQoVCCV
N82bIo7K6VoA6LNdbRrBCY4oTaJi3/idnfmdPAoZINt2Jf9CT3BD1UrBOGydcLav
1TAROy4UJX8UQPdU/6XgDKHbfHU38snVaUhwAgK1d6CoyfTIhcIH98v9srmjWpuG
EuO3Fd90nuG+5LngY1njyVcl4Jbrb4u/yGe2QSWvCR3kFbCXVabnGci8zBAIMQmJ
I1nYBpGgoDvl9l2q7dHoOSBJxWbdKKOyr+SbICPYYev529hnO0XVC/u2hdlssdcV
kRECpH/6EZHr1FHCfmww66KUCAoHLqhgP8eiEMpmln/W4peb+tzYesTDj6ZJThjF
CCqY3DJ1/9D8SwOo/PHEHabXDdu5cYDjg38tIFKWCqTvBrUlFgR2REug09B26ha2
kbmcIm1BIw0UjUkIIuo3YO7SfIhqeMsN8XuPeLQ0qJZbio0e9bTz+Qoc/F4GUBJP
JtmuCL+3D/mCaFKMThGjlhPVWZBXLAM+fBueQicFgSSrGEtEpYvaI3SucI26048C
31DOiWPx6kJhFa9gRYO/sa55xQ/OKCKiPjoqb2Xi1HzyFg4/YkzAcK0FKGYmzcn4
vN0ztNZiUSqMmrjeDaI5HsLr9T23LHexw9cDDu/PVffjcgjFfGNw/nhz6rAi2GZ+
aVfhhh85hCtv3ePBYdsnLBnSIOdNJI8cI/FEwY6UB55uKIi+gCQ5EeLbYOKpSo2S
z3VO/uI3j2StijvlF5B5T6ApKzdEoEIYx7qa517GCopxlNTzZ2LHUShJeFu5Qoo/
HwmuuMaWouOahTFutj1x4749gVOuJkkfv0DfUexsh5Pn7NPjoBn1hnlhpjmoxvLf
8rF+BDgbpI4eeSoH7lGeyoUmgkQNGgZS1FC28Qu2cSgYMwTFX7xVXzyQZXDMkiQm
3iLkMpbq/HMc21d+wadxVlFJTQMrr/ewZ6R7zvdtSPS2qyasmAIg/t+HNYlgRf76
g307/JcWQmBjJEvi1gBsmTPAKcgEU0NqPXw+pDrdycht8q+pJcIWgi7zQZ3rwoK3
MZNcqsZET/0KpU3YfcSkOZeaVK/y+dvkJviLTuK/zHCpd8gMU2tatWnXsYGcoF7Y
28eetxep13WjKA8ERpPodbI8NHv59Ibj56cZdaBxKiALGcBbUOgX1c4tfvAZUuTa
yCHDv9noBxM9A91/gPOPDxqTStj+vDrYYcJnwf41Nrf5QaJ8z5UgwWrfLytK2tOG
jH3+O1AFnVp3kS+a/mZ/+6jhZjv/ziEDgW6UKPGbjyXyjJuWbozxkOSe6KdKlZlv
d4UKTWsudcPuuMFkZ54UhJIvJYPFyI7bIFKbl5EKJwfn89H/2R8DjMdLmHmvVMMQ
UknNWJrzBRgLlD6IVDHkpEFUBhX4lwPxzr7s47OqZ1IuiRzuyBTRuYMqMq9+Z8FC
3MSXHJR6AdlGwpvVKFRWfTqRI4hWSkdA7pHZa+RRCav4gGKxZae/P6ebgHHX2JP2
fFiRru5Tycn4XF86SaeKf5SY/QhFLXMhnZdoee+pSYJ3GoyrLHh606Ks7KEzCAvF
OT5v+uz3oq4EQxxuj3fgGwHolnTTEnEvvbAttfKrAEtfixRTEcvgDg6Y1E/KHys0
mwclJ4nNGXxb3NtMcK8GzQeBjlycBKQaEQfVbQGO+LZyWBl3zltOk8h1GBU66ZmN
IgTOjTKf0vCN4TnQH4dtlpdCtAIGJKvw1/XCSwsp093aRoM8Nc2sHm+UBBo4ABMb
vHoaun6u1v2srEM8MVHz0tl+tshFr39mV4lWdJyu7Vjp1NBk96ZVEnQsGVhc9L6F
yHCDnlgvS8xGmMC4Sd8ACLnG4Lgl9PelieF1LCSa4V/Vxb1AzNYHFTrifi9qqRul
kDG7aa3akC2rcJnJ3o7TtnLFiWQHclZM5ETo8yIKMWp/cDfZofYWg2eZkDUStepJ
oNz4NIW5CUszT15XVclX8vOasjMgeNVBGudJGhDnhojUQYHmkqZYQWnQztg7ah1k
/TyM1nGKscqT2N5BX+/yXy5L1xdp8brbSFfa2H1lmVec/dfVvoRts8QTfCyOfwJu
D9of9liFobuYbyjfQz050XRnwUDOg3wvo21T4CTfV8HffMzdCZhLh6gTHksR3hln
gzDqJnuS4/lnJJ9uUQzSI44iDukaHOO1REd7AJ6p6bslXAZyibSm3w4eSYFUx7Ny
rKLOy9G/J7NWLWu4hKc40sReOQp0m3zWbmKERtSEx2E80SJqBXVoTWrl6KeXDSuZ
0pgvBlKTs/24rEiuDvowDxrUuNhz8Im+m7TxxX1dvXZM2sRKq/EQKZok1waKWfNM
YCgR9sgLgf8ZBqtJsLW+QuB2Dh5fjoedeDyYb5H6YpOEoXUUymhqOU8hq7t9Nuuq
57OQJf+ijm9RLOANieQJ9PwHlsbw4T4UG0L5FU8BfHohiU13tXLy7ZShI47vIJHF
vEAzkEgZa5WrsorDgdFIV0tromsicFedb4mPPocDNptpgR+I1ZnvFsLYpRTBYTZY
dEJowmfvxduR2H06lQykH0LOc3lTgmXWfkoCkgqHoQSSTb+PF8n/tA4uhcGmnUL2
NSY7i38bydhpbT5osr5TJX+M3YDeRPD/SNVDRndXM9xJh5XIdayeuSG+/bxiBL+H
ahd/OeR1oRN0JHd2hpPbpiko8oHaTft6W8Z+y3dtwT8w7eY+ZwvJtGRzi4676R5M
HFAyC3pQ0Ub0gOB9Ww0TXuBF39nbGMrEg4XSBAnUJ0/ddxyNy12LDGq2Oh0Z5+N3
sNSy3R2yxW2lnrXvWycLayFRK0AxfFkF7C9H2igJ6IacBlJmjrQ2G73LC420fALi
RcYT6Hpjc+USQJMVPxDliHOeE1RZO2MbDPxck58t9xITiGWYMU8ciHwbn6eK9FwT
GNzLZEuneCPD+QoHReM+yore79CvQP9WhTZDR8+jvuMc0r5avtsk23mUuOD0CaIZ
DXfBasHj3C4p6tm8W/e8oyfsTESuVWtdQ1Nk+NAl4TN5pN8WvH2MPiAENDC+x63p
Ifk82jlJadC05FeEt7oXpeo3fXV6Hs0mY6HqsIrYXXrfYgTnnlVXXQvlIQK8SlZQ
LJEcahWESD5xtZAFiJ9xbxfTVDUi8kikMjm9g071ywJ4fRsNnfoi/qxfaBD6PSpu
zP7FVxXnwYrcfDO/9uTcLM8QA22j/qMBKu68zyPqXDlbmAlWRWaat4pD1gX11mb4
1PTMnoH4PMrUzXgKDvoKIrhmxr1OvR+7aAwSOG/Baze4K19qJDSjPhi7G8RfnTh1
8/EkVlt/pNDscgXyCognogFULRsP8nwIki4TmUPxaQZd9t5GZotCMWGIlBIF6rHh
r+Yh++5TlddYkR81jVv77UIEM5SgXVZGZg+QTWSDN/k7HsTWEUNMPm9IPrijtEye
Jn81Uc0qYMyVpnZgJgDP/Mg7keLu0zJNG7rJ3XNavLKZrEr3t+D3YIKcxs5phvkI
zrAubiAt02NF52aXsKFpB3HcOeklTDprbPPH/x8j7oc3Ct4A4u2Vu5M+BSzhtBu2
xSmmP13o3mdUAKQFvu6qyUosoYyCer5WJwdQ8yaolL0tmyDZ4NQ0czJs7dQCxk1i
T+9CQziSAo4MTYHaMpqDh/aKFLqZTq8i2AMZ8XZi/zWKhEy44jCA1wKHS3V6Z8Tx
6tcDxkSP5/1rvy7Rk4tlAz7IkrQ9kbdMfHTz65R/8IgTXzA6iC1y5rElJ8mH5ial
Sr1x94UDwpsrbqcmf89leekfcvOZd7NwWyTbm1AKVQcS6Y+x5T+mNQiLvGFyYiJx
mVz2TBI3tKF0b8qmQ4t7Yrv3kgUrXN4FU+lbFGCBiRLUCYpmzxTvCsA+U+uLqfhB
EseVvru6eU+buZFJyVNPt2eHgwBFcBFqHiG6qi23SapLnbdbUsTN+wCq/dxfS2N8
3alu0XbNEjznsMblvzAkBbVyC0dwWQED2dWSCeg1OMFhcOMpmTZD/5ErhlkgUbzO
QOJAbsKlDRZSfFtsn1ppfaaVSz4993B68qyVq5ByFOZSTXg8HUc5P1s8BmFQvzmc
CmX3w+ya+IryWx0cRacS7jDecTzW/Cs4K0jrUvJUjdIu7yVh3Fu6DHscVVWdMZwI
AFTVRCe9o8KtXY9cKw77jgxiBebJC/fT3DH3dyTxcMdpN+lcUJlMQKWddZ2TYMp5
2tjwL6iJAKjMYclAaZ9wCk87VVoPvEyGEQTxAlZ+Y82rzJTB9FCuy8SX+srP+Xj+
TOEk7/VwXheNBiwsoWhj41mBNgFkGREmFbqGmlr+gRlGraxOOjvX40ed8Gb0JNAI
CCwl3alxOMGxEHxmYxcaScH0Qam9TqEroI1Z5JGW9TvM9jUE5+UGM/LRTFBo6URQ
ujuweeNVRlnnRbFSH92UEsc7ICqj0AlibMj8Z5j5sX6OsgEgwR4rF6g9YUfvbLlQ
j4vjSIt/nOjBsT25kWpS+11gh50mQp2sMGi6l01zP9WB7YWl5XxBcvTIJ+KJX9bo
WKXsFW8JEjUYIQKu6aQc/QMu+o9qjZEV2OCqw4Fo7gBui28w4HVucH9k6sgmtf9J
ifx1B2G7VWneXUHBBN7h2YrBrCJbrr/klHqRlQUOrLaoqwQUCEF9V4R+xBLYndts
Eh9YXcMdibazMbOZp+kGAxCnZ0OsKvih/c2S7Ft0FINZhEjUUoJLCn8vJwvdNJ+a
fV7q1hLei+xLx5X3eleq+qrcaC+IR+CU+k7x637jZE+MWxVuVuQuiMkjv4yzuH2l
MO3agAlkvkqh9rozR74NSrR219OGAmKs98sYMLyY8DbpbejCQfMYihFvchW0LgAF
ZIbCwKwGliZhVOwwR5dpHKhYaGMzssGNxqc6cLAfS3pl7ga3A1hfG/XoKkIQvFlB
pwdtqbNT69qznDxrB/KO7MDPh/47xFmlepknw5r2waQUF5a6Se74AMi5p7cFEFI6
dQjkxfmWL0QFAqoEl7VUDSyxfeX/FYPhRS83uKAzoFePl0jnhV+6rQ85qibQQCGA
/Ssz3TcUeRfcla24Sztw6V5NDW2+qTa0q0qcrL1iTH6LLv8qTNfMF33ZAxtP0N5y
FmqaB+AtSyI3AwhWK4Aa5Untv+pCfyH2TWibty9lZM2FJIETuHs1ipNDNfyeyfJV
cyq/wekHJh4kOXzzuMavoXRKmLLl7xINVyLT9/2D/NpoEQxvc2EOcxLvC1Yn/NMR
WuJTzIW6r20zn/FZ00mjG64goI6IY/IIeGrd9fSUxsyokhbYyXtNDsyciPuiGZAP
4VPboM+Ocx0pWKnsFEOKFNRGd+XhRyzn5yxGRETIMKyJtJzk3LHq4huSFq4bP3EI
B7UAdAnCAh4YPW0HhADszZWhUYBPEK14H7aUC48pk+sWspeaUjQwjxKuMhHfl8sH
jMozfdRzNmF4MFKa/9y51mJiSiXiBL17z3M7DZtyEIs7PuWY7lCeILZuwmly7JJo
bQg7QE3k1UA8Hiwd4lAU9bMUCmO3qmXu9ImyW3EWocqG30uWfXLXAYneG4eT7JSr
eUDj9wKSdnag+Yspvw9kb9o1ro7nwhoQXhyKojepuIU6rimRrSI1o/vHnuPlzT+3
4bQtD22qagruJQVG/FMcE2r5jhRnJq8Tcx4kqoxXP8CoGAIBHTMSAzkaKlXnrHRf
QwkuPGRk4RS/gMQGXITx41ufJbquUEpVyfaBwGG9ZgvKVp9GbAKfggen4k1SgYRJ
/srUr1hA2l3b0wed/NKG1XzMDIQBrclFNZZMlfv8SF+G1K2jr8mUg2w34CrVVO6M
KmiKO+huByct5D2owDYbSphDXUX3AOGwbSv2dm2kIuOMPjt/jGPRL8sl4vocO3yr
jciuztlxk+dfXfaIoUJGtUJ5cqLYprWTRhcaxKmcbqn2MDIGatuZf4ikZthRMXWW
WI+CSTgbHnvYvEiVZr11TvfbN0hmOpcwrHh0+lYLon32oi/h1Z7iO+AGE9nivhSu
vqFP8QKX1alVYpN6TB/5jO/u1fSEzxbU18bmmL5pxlo9C+6q3f+uCNCpnch8y20s
CA3gIwqUUSPOkWUQwJxjSHlKT3sCX/SYyd9iIYQg4c+8fYgo5/8dtmZRLjzLdCFz
+iVOl2CDgMjyPzRsxjSyYGbSiQP0Yk1rE38BYRZ3H1XWljjA6cLfzh/tIgcjFtTI
o6UFYTCjgA9qpisZkyC5MEPOcCYZmpw3EJoQdiwE4Jr6LXl0kdjY8idIj0o9PhpN
17UE3gj7J6RvlRMAhmXoCte7/83xsiQkKgy4Gfa/5nzsvQ6O5Fsk6CwCgzVBSbNX
DcGI88yl5l6R0nu0yauYHhegWKUj9w7/R1D+JTmtCdQPdlsToEIoaPw71L15UeyL
ogj+wApDtCjrLNeIsmmwXYczYV/+yzVxoxLo5Qa+tOYDn50MuTNSY/wl64zUrNV7
EcQUtU5vwuYxk4VY/Z9d+UCNTMymbyVpeOEYGagciYI7VeqrSqUGf2ITDv9NFY0/
FXvadK8CvFB5JBIi6Ipz6eZ4cwXmJI4Dx2tncbJy/efUaxAK+qjeohiWXstcCv57
nKUFEtCTlYWUw53CNvdyshAljI9zg7GRoVZeuCdqFtF04prvYnCEp8Sj5dU629Ab
dWlLKzTeEqqvRfvtbRH0uB/LI8Ehu0RVEqsIiuIx/A/ESs+3kzcuYuKg0sjTuklJ
k6pF1jS14BcEI8NPCsLTuKytSkrnoq1uZLGjdfHw62puwSgidT9C4QyQenpT/+ck
1H3tnHbydFfntujv2Wmh15sM9k5HPG1Rxzioq5G7XyOWjTU/2Nzy/OT5oJ3mN1tC
GQ176OfhqrwiyoQj3PvnhrqalqpNdwERtFTVH7457FEtcQI6Hv81W/JfE4rHcQPM
u6miqkKikJM1zwFqI1IVa+al5wRC+szMb2uuJ7d1liSY6O3MJwSgkimXXbowtwxP
hFLwi9IyC4Hs1KoQmlBTjBYZfi2SrhnTUjRINgZ4PMPwDvS4r+OVfwjO837K1T/A
3RnZSdDepNScnNN2qPYHxHSAAskXEGXDXaq8iiEWRmkJ34OjscM7dTM/lkuU8dF0
t+nIXtxwJEJS/m5ZBG52ukhaTQ+pDnK4E2ZVUXr5GwqNIaVqTp03D/lrmg6V5wLu
Ws5bRA+2ZWGqp5IbM3IO70Z7BGfHFfCU3kfk0ww8fyHkJpgeeXQRwipa4eZ440he
7Eu4oOqztN+g6T0oKZAU4jh0aBRgCt3Fo0cOBAR6FQj5m9/byLuvl+AZyhVyAaaP
m+AjK2NKfOcUeXUdPN3ROQIcSkUllhhYfmKdJJfGwR/lDflfcWjfEPSn7wOfoTPg
e3izo1z98/9/ZMO4cKEogjiKfeb8YkVGNSpklRE9UoqqLJB4EI5uU1gYR0dnGbM+
tDaL0HLze/FU7UjdR1rTfxplC5z3V8Nh+lyPdqsaQmMamj4W8LpZ7BEvP4KXlULx
F3NHE2tdbGT7plXYLNglkJLvZ5qquQU/GAVs9jKq1qS69mFelcbGGoXqNNhHIJCU
kUm97RhXBSodDtoZGaDeMUtTOWMgA0+hWXwKcM99VAKYu4BOyt96pUIpeLBweyja
jXGvdlE2zMQuP6hW69FEPM6aU7Ud4LSilqTtt54Is7vcIlfpSUiQX7ehwv2yq1wK
gwLymaSzjm5taHqD2FdCxwnchAyXwtekS+rII0gDLu66EWR4F/aRbqTc9eDlzrYt
2POuQ1jcpDaK9j5b7afB9FGXT4Im4iP1qOA2SoW5Ga8jml3RDR1VLqiQC8CrUZZ9
aPiVc1hvU/YRZmeKSCU88aidhp9WJ8qvUNAY/i1GvCOhvQcOSLduY/A1zqrv/X+t
BA6wD192YG9D14Sn5i9JNXqwbFlVc7sOxC2gMoEzTjH52iaqHExACxND2gBHSeTq
tJOAkMbxaeMAmoOcGaTD1BnoJUao8F+W6kznXMjFrgXK3/EPX+6/9b7sCoLhTloC
r0Xz0XrN+Wu8UTHAYOINP7bUiZtY2/bdF4qfwsYpZnjrUow9sX//3ZWuxpXALZJa
lC2o5ffZ6UO0e9VuNYh4QlsGHcZWxCyR5AurvXT7WQC1c/wfs9Nc+fWsOtRNcqxc
45os/Bw1ObjGEdCWlGLCEKMIaRqhquQaT/DEIzwWVoRW3oxbmCtyusnqvZUEi+kY
N/eQfLUC/5+BucdMU61NbqvjgIcgxWGRCiYgglH2dH/f5m2jJYpBKd/1qEsMNb7J
zf35qSCHBmR/K0Bul9JvoulMAxWgaowf5mwOPBgjIVytguKpDzJqn+15mxJ1PPGX
l+d2mfS595XhIcVLScc6DBgOENwnr8PNg57HT6k7VUwn4VcwxAHkSpG7PV3Cxmls
uXJcaOXN2XbleRTX1BkA8Bljwb5uBFtdzHoKfAN7rJNz76HTJXFZRBvotQxPyb6e
vE7BjhzQkrQdySIkpmWCXkBgr4funAzwoSz2Zomenk8IuC2paJlErZxtXpn6XGJQ
0gHGRowaoZUJM/gwtfO3R7zXkw6UkiMZXUn4FYrNt5/Ny6t1S0NsMEHUxhzzpp/V
hyITmsTwCU+VzTTY45zQMP+64pEJvths+/iZ6LTBum/I1K9GhYGl9a0/s4hLwSi3
8Yl1DhTKSd0QjSzckXRJFkzF5cteEnuHpxcN21t/KMOoREUTn/cPXz+iym+47OGA
rxtELmWrWnk4fnlHNE3Y8LlY/ndMS/NNrsEPLXfgSQfDCdp5DWoTmOJHk+eEjQWu
ES9OlOJV9dhZK8dYQVgkIctu09+AfKTW+RYC53d/7JJPd2yCiDMFXHGMqTxi/3vP
YzBg64dOV4GXtW+Rzooplww/C1I8uUsVnlI27hwbxgkJMkQaXmsLcMaIPQ5ZcdmE
4hOyIC60AgnnXrn9RaQ1yb2TfyeBpeMq+oZQpbM6++MU28I68AeXpm1xhxwy7DrI
YfZUZfL2uoE8w/meFaQAFB20QKmb8T2T8o271jSOvYTRM35I9hFP7OXCjKBqdyY/
VXX0TcvGqP6VI+i+hWBZtmb+uyaXo2tBm3JUdu/r4NvzAI19Mgg1l7Qa1CvjvQLV
qoaQoppWluzitTFchf6ogq0SuxBTKLd935rGg1/BGpghf7dRpWg3XAPOa6SfWD5o
LMlzFuL+ZYkyOfqlG6JYChRz3+tx+kYfbw4k0/jIlcEzJUeRPoxqbaHordc49FkP
zmNHZD1SaKhz56PocilVGYcehqHE1C9C2+zKPg0a1xkQ6xBVEVIa4E/fDIR0yoX7
3h7fA/ugYOiIYgT94JXQCxTMkmG8wCU2YX6xjLI0QPC10E8IQCIoCb8HPQNzIDH+
wAAdrjZ69KFb/u/HgpSQII30nS2meJMOHo9d+OdQ1MxgloDq4097XsACdbCTRHTs
gqGrFHNDl0woxZuoQdoT9G7cWpEIyNttSH+GXlQu/h4EdqrbaxW+IMcUTnOca7Ze
7MSwhZH+56rmnNyHlgP30mUmQaUbHaXjkgjlkvaiM2IhgZ2NTj/E1MVdZ2Vt4+7M
htfclFb/2OdDBEnfy/I9zINvXu5RsZ8V+bXrd2yIo1+YSzPf1AYZmIjPO2pbgSOI
0xBf3J7gDu2hgLvExv1uxfD9RAFkb3QuphsvalOF/omsf5FG91eTE77jFMLr8dJN
he/ZNxWrux58q4/7TDDeyQUA2i1pTSHWBetepMGazisLkWkR4HMQr6ev1bcNpdcA
9m/x8DK7qTYuj724YsknhRC5EWakBekBhS2SZu1P8S43D9qu9rhF+G4D9/eRHJe8
UVZSeSHSIu1onwoefAMheQyjZxhIdAnLDjShp2oo4ElCMXVoigelssQVnEZZw1io
oQ2oGOiifH5LZnUvMlcqEK5amUWLiw/15AwgGYFKHNiYB9IafiqeWrXbDv3C5ihg
k9+qIe1ihbDwrrcGmB3EuC4wDxatuzvm2ITP7PkCKpzqsi4qlIsqUuCumdfghGuw
q6PB3VYxN15Rx+CV4wHLk/RxJmXX8/hfRPxY2bzMe9VP+8ny6v0JvM2ae23kiH7X
xRhpzeyJDt4QPH98sz2z2aYAncInL0JTO2ipYzk3Q9lBFVxcG3LiCNLZxsyD5X0M
qf0ADhyuPKz7GrAra7HjXIRS0YFgpSj9VIUSr6/UEATkJ999rxD+PATTFFG/TABI
xx2XmdhXVlM7ZIdKyrNt9T6LeTDutz5Gctvar19Zoo0BqBTdVVYiAHOdegJIzUNF
6QsF/426sWO97X6HGrrn2bwKJhLeNBWlMl+tZeCoLPxuN6zQgok+1n/MXrF1Kb3l
cBjC4eOdJOY1LjVNQmtJxzOA5zPvwLZdwUNhVyzDFhtY+KWwi02Z98lAsfjABjw0
sekiauo2xbR0MpQ7cRSiEOaFUnEXhgZR38VJusnumzDP49zTc8FpgBP/twxt1x3T
V2rbjjHnyQIPizGOyz7P5/TxbByCrnoPqtdpUolepncij5H9Bz082gsc5Bju4qIH
1vazxDt452VJkql5IJWe1z5BX1ErRMi7HCcgIiuSwIcBI4LAmP+sy3vdx1EYcRA6
AzfXhYXVGmhRwRfoJdhwlMmB+gLgOpTLjBSD/kKstmPGf8Pxq/rMDZV32Qpk246q
OV70sQ8vQJ5p6erH2j8fYtmakUetZh7CreHOiqXgm8eFx/Rqj1bzrp+5d1m8Q+lA
oMkxgImG4XWA3MMKy94mP/45kV2cKvQjl0zw6VJ3guRqWzK+1GH6HfxDASKPr9DQ
6SJp4cBfnoDfAS0HGAqeUaUjKrNproyyHFZvK88kbjS9/oVLQRxC/u/cOJC2QYmJ
0XsMfzOin9DF0fcgTquzS9kumBOpNxYCERPwlOleK+9sBR68HmiN0Mp5iQo4FslL
y5m9HN4ohXxxphUQ4YgzwcnewYsFRyQN3VljQhhsEmGaA7f4SyfFNv3FLyrQwxoi
9HJVsFcPkA9gH9/fgBjtsuEu4xyIkgzqEewsAhRPL42qGVbUyR4gZRCgoR7pLQM5
UT5iJwRSWsDSCKHh+Is22mp+3VL0JG5qNTyWyft8vT0lXQ9mELFSzymF/8w93nia
x6KNv98QC8WIoU1cI3ffLlGADhxEnVK3HbxYkUGQQ45LsRKv8PqOU03hxm/0BVeJ
TWiAn6sYSu0Ae5XFKFfSjzegI8cmEVl1VegpttBxjDh/bYbJx5bteLZGUw7bbuBG
bhZmvWJ/7VnosAKZ7svBaVVwOm66uyErLc0LwJPumZebHpXmA/NSA02nfk+/1aD8
XxvxZ8/80reKb7O4Wmh66goAlsnhXUiVClR0BtNtmpbLjxOO0CUigf63RHxGQ39B
KSG/m1yI9oiSFpCC4/GVoiTWnMCQSm5Uh4GE7dvBDuCKoEzrS7/BDMpVc8YUjZjI
WaCIFA9n4gkjW9E+1TA4A3HG5xX/q/f70kOC+XbggjDA55//NkOvLxK+wfWgMg7S
nZQPAX65jT6q98rcNiOil7uEdlItW+l77rrNNwgbmIIRSbWHRC6drPN3EnKht6KP
oNictnzI1OjXkSIFIxCgiuCkIGUk5jwEwYSAdx9yRGKTQpvRyS7roUA7Gjqzlp0l
WKVdi1gFol9V7KMUwUf8bq379lvw6T8uhgJdqEt8gW3lgV6J6rCK76Ol9ylcfOkb
YK/qCadaxsFarOqwNe2FPgyQCQdXDNUmQ6rG0yorOBnMkDrGVPYNnti0n/ciC+4c
ihZoG/U/kayMe6JUhSsbD/ZWXWyAwNbsyGZ/+hWNmZLnTAyZbYmf/6CdRREOqsZs
kZURUAaNCBhSZBeqH2HdHNDHhyTPS9JZ5OZEdPV7HC/UkUhF3bXZxxkVJwMeDxrD
zrfXlhzX/r8Z91bcqC/1YpB5DpmOw5o+DKRaUChhErCb5FTJxPabHkCmVao1pDfS
BEX+uuYv3x79VjTwpvx+EVbFGTY/FnaBM4yoWOA6Li80bc2FbW6Oxp4a7sCAMnl7
F4ACMx28INtsHf8ChHFIUWbnYfnWwVExB7h2fHTIZj6ss05E5qtnFRiKr4pEb2Zb
gbIIsDpzs93/kG0xGA4KsocFhKUeS7R2Qrdo8hjcHYB71bXAo2baiuPwtSWbyW6N
m6brxeIGr2qNTngBYq2nKVlszkLP9Gemnw0f05pPNKlYkjV8EC92eulNR3eVNtTY
UbcrdawLRNQ7luQ2toADXhV7bIquiTGO2Bpve84ef/LRWnHe/naieyABvMfqN/MF
N3A/i8oMsc5AdEOQZg/DJaYfE4NGRywSYyKjSZHb4XE0a1eXYNP+R0pDQTrQPoHK
E1K5jDXQ3BPez8NPzGQpqB8sH6olSe2stMnnMet8mEusudZGq0xUF3aK8f/kp97H
iNNKaE4Wx7XMQSjyUc/m7cGdWXMFFqra71Y1/wmKrrcwhr/Vo1JJZtOAzI1PURqq
+xfFh7TCQN6Zg4enQv8jkE2vuIr+z6ElhvxPRv4qAxAv5GGtJz78DVKOOXEZBoRF
2fFAp06soElbFxnN93fy75Kii2SyOKBX+aMw6D7CbFjBs90pGD4yzHkj4OXlGsoa
2nK6Wjm5HHEXwSpQeDhzuG9VlWZ7mAQnRtEWgtTN1bSCOKTG3ZVTYdIsyNoThw7+
V1pnYDkYvvJtYW1vBPaef2/TELb+cD/krr6Fp1mv5VBWIdMOPW1U4eAAI5SfWMnk
1qaseuQeXl179pfcR+GijCOtotAZRyyr8MtZwMI0nXyf5SWmjvU+TkgK+dr4F8p6
TuFfwEq9BVK9d+0oYmV4e+hsbV6PKba8+240Q89QPu/5uXZIq+opDLM0THDcIgI5
Drwf29LjQri6dSFWbWUH9BKvhaqS0UQVzx/IVBeL9sdSd2VwoYkpGaNPV6drCUtY
fi71h1lTCz5oWiXTYXOn3qEn8L2w9uA4rmSBvLXXEQJ79WkPBKPzh0ReUu6+YQCH
2caj4RMOwhMiAVTpHNdcPBawADUjxfZjb8P3C1bhuktc6F6hfgC2anGNRfkqhf2+
HXSRwzRdnks8tuEdhgMMGhw1bVW3++uF8BFFm4MuBOP9GydM2/ltHQlCiZ9MC0nl
2ZD5XxzS9BrNnFU4CBgB6dm+GX8pbFOTBqcG4odSTOAmC+7aiBKpB8cEIMeo7rPX
hSFblQuZcB7DB0eunE+JIW+TkQe36yqu7DnQ4lV88Y5c+PxUvWOf9/v7qmAA7c1A
pd0SvV1+DHmqTR9/XhoEPrZxsHnHYeUL8W0Im9k4aH/etXKiOpNcGJS06+thtoag
O1/GFx5BO0FQu6TxbaAFzAtm5Pxmgrr5AI93HjoD0+Ra+JTsXNdXF/O6gYs4f02o
1RiTTTAg2dwUWhWj0xchlsvBlABP1qa3BDK3XAXTeQpUrMH6ylDWud80Fzim4xio
x/UrEEK6We9Hk6P3QPwMoDMFm4V4m7WALxsWRYNf+7ZpkxtMojGYrkHJB9KMR16T
MEHtzab3Fo6oV7jzMSuIvIl37TefhPH6mejDYnH50RjZnkfmm5b7WkCQ3iSkQlOB
yIrYi56YZGdO+mR40J4xpgqTdStn/d2JeR8o/cjeZDoSEG3V9USngSNJoFeYu2hK
iGlI8m6/yqjAEv5ByOiaHvPFpr6VUnFppvZwq0/hQZbyhibcV4KF+dFEKufYudjs
6qRWx1GXXLsrXEHHy/zWDA+kD27i6FX0xZacOtnB89HKo/kfpjweDlkh0ewXE2+Q
G3JzC8aFGdlG0HPHVL0wlgIvOtpeHfWoTleEyro0qNU+5FDeNn7dkfvG27ds8tIx
3oPAvmi2ERenLUFgH03U1w9n7jE1zpFVMc/z+fn0VT0/20q8Xm4FJV1vob2YknPs
1afXU5e97Ej29JlVOMa3EzeyxSyFgh7POEuMaFppK0j3UktwiFWmX4dGYJVDRkQo
42vlwI7JbILkUp1ngXxBZIrUDfDDj/iB2P0EwziEXEYQ0WuLZzd6sQyPtqhebrVR
w2YCYhf+mEBIHvPD2+SxmliV051lMWNmfbfSZJboKk26XAS4hAq6t4NJmicWl5/G
yQPv1SaomRD8lLJDrJkazZ+/WUYQ2DlTkFBdF3rprgKnTw4hlFdC4/IvDnpgOKWt
e8YfHAMf+XZ0pCK2nBH6kQMjNOD7Cl0FORolgVVO3yy67jl9jYXVi7Zm2R60hgCt
EXWceQMNZ0+qTryBhj8in3qk/ylupH1h4CeIPsKMn+dfDM4DET8/A8CvDhzNvgp2
OqUmJWIG6UmmblytCTt7mGs3tngZ4ZIljfPTbBqsnPnCYFVXNUJAB41itVNNN6CI
kV8y3WMLqctpgH88qzQl8FNaD4+RYJ3Bi06ydCxE5IRADk2xZYVPvqahChaRSOli
LlT99T2CGvVNwjJkt8qEge+GOITSTSJ27+iwlSz+ZWl3/11KB4/he9y+cie5YSOm
yTMdJX/3qhXJ0bYKQEshZdmqI+s7dE1SPl/Zn4e5F4garIg+aL0O4sha6PkwJpI8
+xvQ6JEDylDeihAwFzGv36Hk5PzbBYYT7VB7fgxyeRLt4Lt0E+YCJjORRX8KgjYG
YVd4bZ8apIhetsNnM9QjJJw7uncfGLAOp5kZ00JjzlIwoeDaNyIWqQ+Ea4blLRXa
50OSZRqjNZ/GrcuObRdG8yLzPiLXRF+nKaIp6tTZI2fJvZw/TtNsydFokoG+oOBA
LkAqDXME0pzlvmdUtBPpmNIqygEGwLHp+FRcIY/PRgPqW5hwY9BzJNi6ubmRwcje
sxfEM53nYYfg2meDUuyIBvXgNwmoQ/QI/0WTBXA43vKB0UEIsJ5phbn9Ui8UDBt3
QfyeKrrUTx6quXVkKxl4w3jPTKdGmEAScqZZDdKqYQf/3eBtbGWbAP7v0qD7oBDo
U7ws8VuOCQw2A9GQ6DqNYWlbM7PWwcAm0VqoFe1NEDx01KO7soGPEg/Yja4T9Cbb
JjQqhE8AZAT/9FCIecyWVzgUsk1VgPUn8gO7Ln+IX+++B7m0NIgfHkfrD0CcE9DL
cqfrugX1YyxMUDaWVcwTCf2S5gxk+tT0UQ/wfSPwo33DFK/fwfA97aRls206fxLl
UTMsoYoF14lSsT76qzmpSKYb7AzvIYwZAYYQJEp/i8Ac3E1DLZsafWAWChhvi7iu
EYacey5RTvxrdRRmkP9xLp4cPRQw4rL+TLoEjiF4RcxSbNMgdKfJYjTm3UqqXv08
F/fa6ssCVnb9Z9aMBkUKjXpoM1n1mYG9u87upom5GFCQ5tYqOjnbzOLxGexBZyCM
ykbCpzfc2JZz3LBcZzFxpaKvP7aYhOWFRwR5mBtPJrvcRU+njJQhYLUKhxEgEjOl
C8a0HKvCPcfbz2BM3ibcn7t3IBQGQxTQAv5Zsdoyz5dr9inoI3m/d89yPTvWWCmS
KYzZhIlSlLsJg7kchXJpC+jhkdlSS/V2ZaD78fLdwvXq/YIwzIemLVWtf6pBvCC7
fvdZ5vQ+/KEzRpV5agiOOypjwJNYR3pmwcITF7mX1jG14g96OYNTCGhB1ovelXwS
/q9M/e7hVvzli0R+SsWFYtnIBI1Zrvj9tcIW4zOQBaxuCzo/8r+4pNWkPSfdrzDk
AmRALay5hii1daIKu64mctYQZ33aE35jGVMXIhDu37S//EG9Pf+oM0uV9XMcGjzR
+Xn3aWxzcLZBf7CKLGIAyLgpuE/7Rcrg8dbsjbqMeFs9H5D86IeOjVpuADbtPB14
IwZMz0sI5vI9T2jCatKrT20bGjfPut6H1nIP6JUOxeJiAZi+Sel2nlgBCYUFjh5P
P7FfwIefKwEjXjtEITvfa/R46z563JY/ePYHurVbe9adZ7XflrWko+bZ3Uc463Pc
zDiQ+3ckkCbAnNk8ElVjOgS9LabWKpk+/iuCj5KznnRPuNBao0cAtoTqZlUb1V9C
hc2Iwex2eePBNWc54E8MPpP64RHxc0USYZ9xUVLtbU60tFeY40t34QGhezLWt7j1
PhDxk7uyIxdcozIenntYTzB2ljWYtpMmdXtcJfV5EkmARuhbELrnnLogCq3fNqu6
p/MSv/dTxLtivuYPiYMqkmvJSSnIv/vmbIOM8e57j4pd8IP0ceGbSdHN05yQXlan
DoXBwRJYZEQ2LV8pVUquNO1DO25tQgE9sg/UU+0wrkCDdsadRXhFaWP/CYJXuM0N
nOXc+LtDbHP93Z6W4X0717UMoQDN7o2qrjTLNnYXrPYffvN9x0qlV0QMUHmdU2j4
4Z/LGOKoAP7XfJUQUk14JC+SUGCpAVkwPYHrhy2JnelSjQDkf6hQro3P2BC/gcqB
5p+EWJb5MAAblfYv23bhDTvf9QwXPpYlJzBDzYV3b5YefVXYnL8H18t+dpwOYaUP
07I/Aw2fyc6RwycpCD8Xi0KqMFqAh89QThCPjgPo2pXW44AZ/Eb9aMCqGvzzIeQD
sEaJgc9t2AJ1pZM7Zzc/dBt/He1jLObSuWQs++YbvfK6hRQC2xc+rnGl938Tv2H/
J6IbxuQUZKNj9pzPGwXL1lZNJs8qwVHaFbzCsEozSUBEAmIkQYgpL6OK3C4iJvhT
qkpQ9W9OEtV1ISXW4gq5aFBYLNoKL46CIxyyAR/9aUJr+9IG/k9Bg0oq/pRtWgtP
BfBtxx+ZlrzVzvyXhGfaMNKCVFDF+O/Vjq+xd5YB96ll+5U+Joegd8w3O0ePtdFh
50U7jNh3shtBw2WhqxAmidDdlZBJUtbl3C56GHj8Y8BZZlaTdDlxybYwL7g815RL
LclIWiHS9hfGh7BEdi1nw9uidtC1A83jo6NbOwPOLc0YQuv8Ba1q4eKN1Fk+jFGI
O7oS7IteKK5O2wjlTCYfwmRIcO/MiNWlgQqbBk9ijf9yv0QyZ/WRZsdZovKlNwtB
EczX7oYqXWyKwXbwGsvdV+SqjtL0pTHMNn0Mt3TWGKviVcQahPfoMSiP8PDSfFwR
RWHIALdG8S5j5KCIyZ9oA2GMJzpNX6gOgA85sk4tora0cSEoEkiPItSUKr83nQoM
NwbbCepg6YPEzOZ4/2xQRHE5tv8n8vgsKdMt9N1f36u9mfwbRwCVIsm+rl951M87
KVaRkrmGwCaZta3ptJSs7uykIqztC9Ym4UvVd1lbwDza1CS3aRSgDG4Zp9fhrs3G
hNbNaQmJLFrSVln7Uwkg6nwutaYnE7FztLYJwUOjFFj4oZqQK9eyhbjH4lKwwLfO
xIKFDlVMqgz36Em09wRknNPAqWS+6GTA7wVO0EyQ4QgWGkLMTksGnjHQmH9pGNms
1bgplgAfoLJVWQyelA+ZzgA+uVCAUZyzeh8pvUctXGaNkdhjpp4AiYz4FalgRoTh
E3jIF59ZYs0RsxFz5pXJDug6sCpApxUkKElqD8QWFztky7H/CgHNMs8zbDJdEAhh
3KG9IWcZgPPIUZ/urr3M45/PKCYlcDku24xHbBOLkNLSOXy+04vY2rEYY8g3bia5
j1tbtT0eS8vmCvWRaMydThdYyN+lhZgHmrY66GCro3lN8b4/5uoV6uaDPsLnNmzT
yhNxIRMyJ8mP9zStlmSguh9ZooOiAhthERwl/h99RdHA5Js0W4IoLqb8nNlG5ZIC
YpoIJHgZX50zIr+BKP640pwDDN7lnGgzw4OKKdY1Uj41cKeYtx9NQdw3OmEHtPS6
/GMKziVK/Ph1glibABhPSqcfVahDZMjc+4NudMhqcs78ODXmZceR9OlM9ZPEI7TC
OCXIzIARHY2pcKerddoorI+MSF0KKq2HbfDGF1fpO9qGyj+zdPd/hCGvYvx9VZ6M
9Uw25weOFSB0EdsRJdL/peubRqGZOTkY0KoFW1dk3Me7qMvfv/nTjhqhmG52HW3p
cLSDoJQWcIcrFJ0kgAVr/JiDCIfGJZFlXDd8/HMzUrJwTI6o9H7b/OfcOuIZnyXI
QniActaRQeVFi/klMU6fmOlBdX8THZ+iGoHfXMu3YCyD0ZsOfYXW+pkqkl3giRKM
szaT2OpGxVw0UVDyqSXtjzLsCrr53tZI7dKlRqOEsZgStnVyNZDBZE2WwFm1QR4O
xyIBzO/PDEyC11BYOe45bVx3vR03n9994Q15JrB4wlcweeHZ6uA2GreZBteY8YxY
Nhq977Ml1gUsfTJHI8CnLvRXDSwmC9GjTPbmT9rNkbRZlbEyJaNBM9ctK0FdFxN+
Mv9BFJ5IMsMdEyG16sVN9GcOUjLsWufCinocGAd3fuiIEuMf+uoWGmAQPUcOpoCY
3XuH5aqcLeG++jUITk0WFISIqKUkwjtBHu2fpNYKwi3b9uRnIkRDjkRb2lvi4T/q
CQnSKOSbe5YsgdlFg3LHpRrDCCdFHh0hGCqeT5NznHpechkyfwix346SFks93zLk
YzPNfixKmAA/n5wF32lTfdQ89/EvTQyPbqB8sx0jw5QALIrH7pDPXyn4unhe91Tw
W66vZ3K+Sn13/zUYN6YMQ/sT8gGUe9XG0DiBEeJro5A6Fn414F6KZNlp1Cs4d35c
/ExMATkfWCv/d6JdR0xJIS7YCE0BQ0rxUAd1RBfGNBFUN3GtpAyN03P84xGXJyex
r+n8IKMVBVXiR74GaNUFKxEWHcnIIfh2r4uDJcsgEpqvsICdl+yyQqTUqoCTTyJT
jo8RNRPPcrUsacKoD8NnkRnwhxMuwlKRTD3hilxOLoXLRkFRDgD1AAuFcODagOq9
Ri/SXdbr2KOghKHTuDtGSKmpq1sQWI/cDIjZtyeRC03BTzVzHxrwNmVGQjD+03LB
omr/znd6FGjNsI0+m0XTMnFGgNgioNelkg7Pk0D3XU/gBMA/N5JoC3BTVIGQc3Fj
2aJO0KsemT3lZm+ea+IPLJLBtsR3PtmrBaAkU7KGNDlbadBzYja+dK4v+EMT2KhI
1ih8Efja+TsCvu8c05AyXq/reJ1/EM9Rx3v5DCgxVlrCjquMOnWVYyWC8zElp6V5
BbgU+mDoPEYPjkct8/n0bJcs0NL5F1mQaDQi4bA6fQKBRu1Sq++pN9N2KpY+wm9p
G36/sJGA6nZxFHuAmCX5LdLq8Rce3Bklv21hwz/PnTW7xSzxakfHjNILbX2PdoGd
ceGbi48OTWt5tMzHH58QgwGeCYsIR74XsOvTcviJOy+jsdBlGGVnNn5cWNzGZ4ps
DSKyreoyF5vo0+frK99b7MvwuvLabMrEgygOKOCofXmEWkR6eIG5bkvvXsigYr03
fvmabZd3n0XS6QLy/3+fj0z0owgQRH3Edrw29VVhcgk6p/Qy81BO0Fkh0Sjfr2lW
N+jKn1Tjwd73yGxqN6VpylWniulI5kDeA+rEndgUt+J0LSgxorhHHoNXEd+GQrpP
JHSGND/gYj1xcSBGU7I/htL88wYXAyWHyziqvFMnYZSTCgMTOLfsvbqNYrlOjQIa
/OhyVQAJxU1Wr2GTJznwiOdVpzDM+dsfmiuTyp6V95sn4aE2ENEkWN3X9OL56GKQ
SUS2/8ZVXx42+5xNz4XAbPP0qqEAOptm9wmcdPovTQ65wS/udekNY2dm7v7xj/sG
Nk0testd/cHPZ+ixIWkMXPbBwEbdrigB6gFmy6meRhp8eGmoHgufyQR0qPJ/mbGc
v5o9bWKQMxpQ9pM4hZYKZoymiT+aUCSIok8TzwjPMQT53ZfIzKjqI+HcaVdAqWY4
+H58KSdegx0KI9z1hZZVF1dCXxYnfgH50FuP/P2R2MepndIhMqAXhfXqgoEez5RB
aQL1XmNDgsSQ8gxp2fR96JhymWNNrVOf2hBsm9rRHHXCjSjggLSZFQ/x00ZdQJ12
BuNzxcDQWJCJAnNs1SAowxy/+DJimYqfkZH8QrXurGyeNFB5dR1aNWxRfBLd2jZM
LTf1kQ8XQ72ImSDB9dxZm8BQg5fqbDYt3ELdRs8WNjxem1OtDebvxvUCG7znIjbh
3zqwXxFKIX/BmfGchLEyR7HL1hWuvz64sZoir3D1L5heMIFaN+WRCD9V5gHHjAWR
fsNxZvZpWgpA+yJ+ONohzeIe7VD2HDXA+xno8iIzWMHddxB0+HwGlOZUrCh/Zw+3
5CGwCgsuXONrRZQ8O1IBZA/jj3BuYt2VkjsQqWXm3B2GIzCPKZ6XlaqW4oM7nsWY
8TzYeDDgqE+wvaZ64x8CI42yDTNVe9uVnH1uvEipxguSD41rNyljTrjC1U4rZf+p
ZestAgFbZka2MFNb9AVdxVhUPYIJQ+qIROegqhJWBtFyvq96mr/WDiX6cDX3+w02
t2VBhbfNqH0B2sjY0TEe5z5IPC4SETWamCA5kd2yg5jsBdv9R5ZEbDrrBCyRUIFD
L2p6BAGDGfQco+zC4iHWk0Fj8TF3qdZ7tLReWKLwogd+YmvrHctALIH5glqzEXS6
i+TbdYaCceV5EoWQNi8Ln1dS8YHDUZrEqlAYyw8tpk05HBEDH1bisiNbOcdipdVf
k8Fn0pveITg3T+7YF6Dwy/EXX448P4pY2/iBKqOhoXm40Ld4RsrqOp3AaTVChSU4
rIk+keMTJGtt1MRZPFAKlvhtEEmX7LG9mJ/CWL4A3CIVD/ZZFaWIRoTvism6rZEl
/O2nSLdxS1gTtxsEqNBoNMICtB5up1/zs+90ya9tcBUwlI0GgCaXeC2Xu59DJdqw
7YIl1d0pIQHVQSzHofZ40qhsEUj0jMrFfWY7YT5gwYWRYDJoBe50L2icR2RtTZc1
p4r4iarnjDbcJEstJ99M/qW5MyKB5NtjtOZTgC3kisM5ViXzkZtVVK1ST7dosmlf
IRDFolhiBDnbQC0khqtxFDJTlZc2+JJuhmCFce2m7DY6bHJxr4UJcEHoOdku1wWB
cNTSYhsNbisAEDEtXswpijMMr3XZEJgWlHc6CjhJV9ZS2c+a2SfTeeCDoLhh0Rmo
M58ZT/Fgsv4iCFkPH3yUXKW1bAYKVVMNBLV9oU5nebCw0BkM5VsSaetXBr4UQddE
bFkwADuyBMlmqJE9ST628P0wVbQrllVyFXk8IYjlc2XYI2cdetN1/X4Lyg8+ZSUu
gK9DN8rzo/6YeUY1zpHA5ha9FUIrCperoV2TQkEgn5Cd4Oo7rWDkvstwcmPO+B3H
DOzmOVG7omlEIELc00QVlOW8oxQobpz0BNdUQboX4H2y+U4EjYZ31kr0hEzKBKET
m12x3IHpPvqscCWb9XX8ODAYckmlLfxd2FfQ8Spk/vfb5PmEY5qauVAnONFH4gzy
nOyp/q3G3/KYdgvT3xwCiifcEEnjLur5GfHJcHfWlaKN0G6VErAMySMAZtqGfxks
s/LVxtIrxg2AzDvnd6EA0uEQoD/rdeYmUb3VIbKmXCawwB8xs8x+0wEubYGrYKOU
0dSBG5DOaDL1bx2LuR3WBtbUooOOLtSbfm6URPHlYwn2q0N2XPit4VcOuVwITGVv
89SlsKyDFcgxptPphhGF5bP4RptHz2OVOFPVh0rTdGUgZ4cIo0W8xvBMiywRlJJ5
b4ICX1+ZLgLHznWf1dlolVtB+PTWbSFMFl0rrQxEF2rWcBPDf60tVqc761S6Q2Bi
idnF6NZ8+i+z3HbxPKFbtiBUiNjNfThEGKV5LgesZlZnqU6CRs5ZxYM2qujqNAzx
rx4e91+E9pRlpFxhp937gDRFRFyeJ8gVVJeOj04izMMK0KfyL+3A5vbTWX2nsRx0
yAvn5yroC4HK64ZNkAwdSdX2wlbmfuPhBp4wRxyTQrpmfC3CF154ESxBMh/aB3zj
5/NI8gwQD0wIDmHhSFAy9n33zMGMKBiwcAQ7ZvgO3ge/5IYUOpzQ/jS0fmoaGz14
7snkD1iiQbmgdQqMbkcG9tAedxGrme/vPIZZmgrw8IPMgfKyf+sKBF53SFkR2R/M
20rCWvQYCP6njjv35uimPQTS7Q1z/n5prLUYmeLZ4mW5k9WmLdhJHXyGaERPCuHv
0mIKhQQYNb6OTtXWAy6/YUhIWsmvoUkTZkcKgsif9Us4odUCt5XYgwSMLtBdKjnt
QGAuqxiciW3a0wSIaPUzwAn7WTYTu52+GPbLqHiFvSJiBqCcs2QvC6izKszB6aDo
VXRjziSolmy8Qlx5ly1LxpC/RXl9xz+XPBy3YbUuZP4B00J+LUuVLQ7tXOJg/iYW
imAazd7O7LL+ESxMAMY6AY4fIy2XITdRNu1l7X66XckG0ab9OjRd97LJ3AqsucvV
a7u6sgtzBmN+/3VFXy2KAImm/Ol47TRKohY+5PP4TWWKpVeQ2YEZMKuvAIsAjfnq
pY3zUcsy8pAnQvXCZ0uoOQfvHnkZGGHhtkwq/ttM+9xMPSkcKfT3TVBHwPce8Z3t
RcwSiFN9i4of1CZG75uH7zWeyQ7n+ZevOYacCgQylIWHoQRxvNFHTRPoVoUjOuAK
gTa7fT6iTdD51ZB8dyvcgse9sa8WwhUYgS3jhVrmjwTXUOwUGhuk9xA9+w8FPpFk
jM9xBZBxEjxhgDAGxEaDN1XDkLIkcjDQN1frpwSTB18c5kRKqskD2QaftFB7gj63
taABwQmluRVHAzauj9MPi9b2YEkyxTt1gshOk7ky/O3uPPi8musG7FZT6/7u0a8h
gI3LKEhM56a/O4pVG8eBmVvfPLpai9Kjz99cSIjwigprQyta9vSNbQcw6xHiIG4V
AXlXMlUZgdB5fU/tfvgTfV68FmtAyk8voKYuJHAM5M1VXiqRpN0kgphW62w78CtM
xD3D0Djs61qlqz9gHt2ad/5VTwCmdaPtuFUCWBTTp/0Kh2QqP/mr5KVW45CI/zdn
fMywkpAqbj3NCxa8N623lqPXWJMSUPEU9mdZ60HcGuDR49GZlJxG5lwE4GE1YUNl
Nib4lVgcYtWYtT+MhCrhojOYMw9FF/16oyGbOsy4sz2ngG3TCKOCcHDy3EZrXwOK
ZeyB3AYl9Z6FdD3rmgpcn4DPaxPdIzkzYLe7tVEloyXnsB+IU3WnIaDyYFlnFUhK
0c/9gz1vvldeqbGv86jYgBeh0DMqbnbe5pV+VDQCwQrg2l8sIiUL56+8Nx99d0vN
eM4SJH6a+DJnVK+MnK7SgaNng6jerx9I24GI/MWBL/obV5uhM49EU3niWo8arGWz
3X7liEpKYQPjLewibZutWmmeSqobpqclnG59j0vrCoIbXi1fAoBxSCHKMQRjirjN
w3no75t+bNrk1JVX3ZvCKo7XQUCFogXhzE+vYBAY6UiW8ouTFpVyaj4Z/EaxipQW
p/pZn/9hSwraM/p0LLUVXlJwIJ4CspYx6zkiSnkZ6LBNePJEp1cxMe43i7U3gwcg
P7rECKNkSF6OfjzJo76JN5kImZf3xm2XpJqhf61xZ9+l+7Ns4DGeGo3NgX5FUyD5
b3ek1OQ2BzhR7cDF/wY+tx9DGzpnshBdDPyHBpozctAVSFT+szHHTVjjvqviQLu+
bKodi10Jru9gp5XWsQNsPfNednd6TUJiZpuHDJvqd1yRw5SpdY7LlfVVGa+CfRus
Ffb2qX9fREF6yHS9OabvnRsSu9MMJdA2rmPyztqbsLKjDf82NoGapzwe6sUPfGpW
4ZVIrlGsloqgBPI+7MZU7wHnbo1DDdiQs3V/W5jMGgFDAdkqX0P4ST7qbCxqZDSG
1q01ybEhfuHCWUwdpG8X+e36Aecm9WEhLw627KbfP/Tso8eLuMcBP88OzZ4hOn8R
IITkN7Sn69wpqOrEr3fXaVzRlKz7RkH0I2Til75XZT/aF31sG5ZLDoVuF18MXyTS
B/RuIEWtfF+RL6ZKH0a6wktbh5QM0OPhsXiPk+kFkgngjBG+WNSb9sZyWo7yZoqQ
2kKbYTO+fNoEfFvGRyE8sligZTeMrZ9ntICsFmjgIXHjIVWF6+oWAaTSnOpwMXO7
5xcc+qXY03u0VGs7Yh/AluBGI5ipNIq8F8J3ECTac/1NxPlgGN9gkpkmrE7P1fd6
uPtsQc6wCgrzUQnZ0ISyo/W2l2Mvn3WXOsx1NijZKZ4lvHMaxKcMXz+GF/yOe3gQ
JuH96lrOQS5UFxQVD9Xn3LXQ7t7HQSPalv2J8XQ17+9AqN9Fx50xlQBdYTuGwWWE
P9YIFtJmAWduu1FnoR9SfjwMEn8F/qofcRdZHiDpO/FczRv+Zvl/hJtXdiK9ivj4
Ws+Mnba+TUHbyAvTFfN4pH4NswMPQUvjf2iQnCpdkOMjwoKOfWoWzOq4au7QTe8D
xPj9kEG8udan89KKtjw3qOUsBmu5e9UrQ9AmzsCXYbtlL8zRUlf+MnI1XVqY6Yvs
NkrE6kzkURSijncPnG/vuXGx/qVl2gyW4yYvoPuuTNVS+LJOfNd8k3sWp0eT31Tv
A5+lEBT1eOlRxSydL/irQuXw9Fy41xChd+pk5KCvMQwogfRPqeROAu4LrrIP0+ZS
cwk0db/9oET+OeZq36G7l/r+ItZbLOes8x8OYopQGoJZnVMdd6mAwf3ZUFHORivM
M2yGsxbGNPkbYC1x2FYGE0AYhDyriN3u1kUqWRhUqVCAqq3/Za4S/JCP6BjGAfjd
D1kcsQVqmLONC6GhGUhYlgShx3jQ2Norto+XsHusNMd2HsFmT5bGD4Q2Gmbp3qAQ
pdEVMLsgcQr0IIySl52Im8PZh3KrFb321uuOHf7AEOy5y66MO/MURsJDgIq5WmXL
b86RqNvSajSOcwHd/rZPd7pKjLdFKjhSvRn9eVOT1bFiILBwQWbC6KSB8ZT+H2Nv
a/Uh9/HdSOBDaVwYFGR58Ru3G06QwAyw1387vV/hGDI94fU9c8f3mk2ZyFCBLD39
bAFRyhdmvaHpY+Yo1J2E1KZNvgI+FxJMgHFnm776rXCUB/0dQes4S3XIcHDOuO+T
Eq9/AE3/8dXPo5lPaVyOcTAkzcEmtMXZJZcTnz03y/iSCoAMI+kLtJsl8E1+QZ1t
eH2q7es7AgNAYZdCtiuLOGB6ZScya2VE0QcruKOC93i7kC/fLAA47w86GsH6N0rG
1g7a0xGzuR+SQm3DvaY/Zl6EIcPmCV54lh4yBq6H1mRKqSJ0sKEdqGojdTZp4QOe
F9eQMBDGKnLCfVIrv613egZZ5rgzw5rU7cMBrUTPBqRn+FCsNL+cdi8414e5N7xZ
I3ctC8rlbYC/PzDxVqdyisaitgaTHo4SjP/2NK9VC9r6eMMfg+Vud8REJM/iPXvn
mWqO83fDtN1O8IrPPWsfzklh+V4SejD6KQP0greTqlptgesAi6uxn+w3EG6tQL9k
4ipc3kew/WvkI0RF/yUOnKcMiE/sbAgkELZF7+uJxMpZ5ltv19zrQ1wpGgLCSy9h
EVCsues3ZI5E9XyOupMr171s1bbIhejn7HXjlsOQ++jihGIsphNLo/5BdZT3dRnx
PJAgMJqK5YiQcSlVkKvEW8H43pEmrtPfJOlMMKCKgVUztg9T3DJZmI3g3nig5sAC
BYiM5kKtsOxUBYPd2rYaoAJ88fB9zF8tgQXYyglwr0kMVsPxtnnL+sV+ev1srixL
AUpPthYI/BUpOgfyu476P+GRWVsYt/ERc7oeOg8qpWhNcUVSIFmjutiiIvanCS+G
mEodgZ1DlQyBpJ2V9lnzjLtZxFRmyF9fBBaGkTMAoziNKSoO9q/Z8vOzMtbNUDqp
K3v3bEfMjh4xQd0gZI41Rn8uRPuzSRUona2wVtH49ZGI60bXavbxstrcyFFSs8sR
v9vV8boQO8q/2lV472z7Hd3+WaP4s+/OuGkNYzcF2X7w344vYNul9YOODfCJqJbN
GFCbziMDm7TRHwaejs8c11B9M3H8DukPgnpTHXff8jghNCESn35IvYzw6dpuOfnn
p3KbViTaE9bYYdnbEa1StR4q70yzuceDiWgc8ePAuJIwVlkSQXJFKDkld31uIz4H
mQHLFUoryWqqjYNUbjzKQyCFQpuQ8//Ol6NdPonTPea3PXxQqI4ohKl1rmMp7u+P
d4KCn8kBmGnoUTc6aSgw/Gq92LR54lRnhSN+rLxELfOxxRrlge9XtQF+gQHRbe8M
Pajq3/A0xRKIrQq/jlP4kTqCoOJ1ytiGJAma9TM654rXzqcFdHwuECOXaAumI0rl
f7rXyKuqV0+Ie2KSAeGY1nazYijBGAcQoWNcx3CqL82YTpg86zv12uSDh/RQT5Mm
qVROe++Aj0J1c2YTLXG66NAwzY9hYn61SpVQZjxs4hxGqb1lgucXhnlMuVpxE8un
QrP5aPOjNONnsJY1VHN0ft37zjo66vCiNfg5WOPYd4ECOx39o7T7/+LGF5eQ4wu+
iHP+Szty60IjVaWN7PXquxlJyYORns2/cH8jXUh9EahsCgpzjd8ruHdOA9ZvLMP7
wCKnlO1caeUqsuaU2ySdZMBCCm4w9D8JsgzuantCLRwsxvD08+kNJ3yp0rNtgVVK
oSlQ3byFIFnzx8qyjwAQKrd5DNa7lOZSSTiWwP81YismxGTINjcLAlg0MBrEGbEF
qhPW8bwULGugH7Vx8QAKHRTla5ZM+QMCWsW++Y9W2Pb4GkioRyI08kKxOjI0nb3w
pRfQTWfbPBmpLUmTg6HI/0YwcB8cxKpT2qDeZ75DFXDxpnx6bWibRILSpe0VqCEA
FviqfniUX0hjYtOum6T3rgNONr7B1HrBAB5V1KEnPrVe8pzz188qXbs4u+7yT21+
oNrRYhdZbh/HLAqbLL3oA+4rZ+ScALKDZ3Vop+T6k+0czSDC0p59uWxNl8S6F0rh
qeXqCsQIH0tp8vu7JJ8HLaPcYpMFAfQyToBishxYmLSg1G2RfVl9HoXoOsRDWPXp
HZ12/+CEMxBw9rI94za7lyB9zSM36Fi5BtaXNccbQ3jGiN+HYMrfnhgaZNT+Yj5B
gvd2TysajzX33o+ZNWlDQL6feSPNaB0Ch+048kgyOmsMVXP4uUfQ1iiGiHuyAprG
rAWPYGZJahuop4vwwNin+3gZFVeZz8yeHetb7uDw9DtKOkDJVHG61U/SoiEH0z1c
2keIQ5VmM/8Tbx8GCnC/WaJJJgWWKYNn5nFtt4AgYHrAQyk+x3Zd8kCpEk0wNLF+
1/7oD1A/Sy+IJc3VI3bsmEeWdhz6HRfDtp6WntmakqOUIkXJhdZwLywrBUNvxIZI
p3T2SrXFtjP5LuoD3x8JAttP2Hhurlhz2rMfNKYTUd/NW3Tmx95CSrKAqkGPdNDs
OkSgKvUtQ9XQYTsOIoQOZ72ri5uqrG8oKgCLUMZvLs7BozKA4WWYh5l9V4kapHSm
hpjvWT8an1h4XqUr8wI2kV+n1KhsPgQaTsLPbiRJYZ9/3hn06lCbCmlw/+7l/yJy
Zu1IQFNeoxcePcWQ0qnkIL9cCxOCdWl8DXku49X7UtqBPK+B9DSQeBtMrV/4hRsv
TAsZpP1w+qyBwQPcIUELnJP8yuLth9fJROYeySBte5rpCwqhiw8ZPrDlPFZwBylv
n5Tu+EKcDxIkGanYoFBEKR3W4TJIcxVn4K9bVyQ0Vq1Uqfo8w9VtZaBtlE27allm
3f3EXH14JP4VK1BoUaXOpLiJCKBTDEBJzx5Q6dd19j9G3JKnDccaeJf8AtMa3E+A
Zd1o15xA6gt78LBfATJoPJL32ZrsOfXeHZ6G7+RGouqYFMZKZ07icSfoOrOmcUsY
aon/0DXZs+mVVK1WrUGGdsXpB9Ky7U11tj+dLKwmZ+LjYTjLLjXLGNn1nZ4JF6yR
5l0SIjjvp+DmtCtmHwRDlvxKpdIpKiOkZ2xXrdfKmZKlnjHyXWr3O1kdN0XY8eYb
Ycxt5Iqt7SIcak2sP5Oah9oyvABKrFn1DAE/LXs/c6lh+YaL11WxNqulO+2HsUiN
xUHgAEcLiIy/UyN29G9Zr8Qvt27nPT+MPuhOG6lRbyLVKs/k5lDTJSzZy4uMJV5Y
Ji91qh4TY9k8beGwpyVDpFJS2Df5m2SYdI6F9gLHPb476478DK4rwVj8b5CCMR7w
05Qfb0q6abNCXIYkK77BjB3iTLgkx773F3wCDGzCwbvYONo0GqBmUry8+vcG+Z2j
EGIgT5RGXddwT6+KmnoqgoDPvK6KHMQXtGcd5Boi5Z4yLwo3+LhsAKW1l0Ftz4NA
1OUwEBwgUUxbzvwyUKjBNUB5A8nezdkRSDemZ5rnS09qlz890kz0S4Z4jHzuT9+E
FQZ+1ugIbjfShli/eq0BO3JXMJmZAXQaNkozIM5PMeXvUDht4nIFpYqtGigN41xo
rQzOGnIiwAfPP+54UG0/Dtj7oL6Yfzv/tRCWG8SZk5g9IuhMlVIB1dSltPgLNEqw
5+p7zQ/HUOVKUYX5EM/oTy9OGFLKMr1gRgVw7U42q0BkRDnVUJWsXTKMPpbpqYNa
lsRLe4B/jk5aogQnGlc+2gRG1+Ela0wkylS1JFXr0KhSihIVd05Gz+0rR8VnW5Q9
VK8ojf5MRA+u86wfE33autD58qnV8f8WDke4b1DbVKeRkMbKbHQiTdSv4vnxzpvJ
nqmAdxFyWFcLDmAjcYSmicXY7ZaG7lwo4O0iTZelcIsVV0q8BpvjPHiKwHO75es4
4jsjyz70jKQaZJu7/hctFoXQ5C0bQlnezwppqTFg34O4oEd7ytKw5miPlFdK63nD
Ft2jF9TVlpCZXWnJe45FKxtNjvB0NGImBdGe0L+dm9VFJWqql5MRlbCq39H8W+6n
wj2JvILrvdQtTDmtHD5VJPFtiQ6uVBg5d1Wa+ZbcGjGdprYH3/CfW8zmgsFLkD+m
XxmbnkD7Hm+q3e6jxDWjKDMtvkyNnjWLSiLkiUH9ecz0tafczoTaV2aLkmj0YQlJ
4RKh3y7XYJPzG6a0/5bzVPNHVYSanymAc1nEmSh+GyiJhq5BoZ7SsGUFcUe4n1V4
yufEaw/Abe0UrH7TSFD1vFlaVVdD/OjxFCfgmLm79oDjb8KnXZs5Nc5yGmQLktA4
REotUyHUewP6jX1ChLKXxNkUdxz7JIYve9PsF1W88+kxkuyFgdNPnO2qK3arxD7H
poWhax8C8ylo9t2gvPdZUO/+hA3zIlVHTlQl64Ff0eqcTQsOXNFCByYNVV3Q66xI
JtRNw516U0/Z7zyRSZJzfHyfIbeg8WDCRB5BoLqI1VP5pG41RbHigQOhWDc1onM4
AbSqkxDS1TqbJ/dqGSwBg2GK6w6REBwZuGTCZzNAAjEnCVyiHO9ir9PStsL7lmUL
3IeidRitx2LPD5xO1O5E63HJRmslelmznvwEYY2WDR/sMqfbTNwlGTOnTPSevmmw
HgpZV/vkLv0uZJTUYWXclVXngaejFcWNA7J/J5H2dEUaobvsDt5EkFtqT0HP1XY8
v14iKlioht2JY82qNw2lBUW3mo1W0P6uXfE6Oo63oUOnMBAbdi9A35MmAEbQwxs2
RaTVP+UQAvwEggYRewNVMPcb0034TnumaCxjcjx594kadwtoVl4FSPyWO4x++L5w
J6Rs2hqSKQO8S+c+B1fLqmsqt0Ojs6nUWkT29H+wA3aeFuWNCcNDgMTebE84LzPb
xY0BzlkogfSdAnBbyvD60SgmtIe4s4N3Csrkt+Ow9c76xT+esKCgdHY/hAIWx3g2
l+rwrReL/gwH9iD+YgPXJ9n7pqmHzOjYFC3ProGfBmgXjX7qVbdSZ4yaFMgW26Gm
Jy065PPoMMmi7PIdkHFTdTE/EjtlnBvFxk7bSj4YbBhtaiRaqKuMxNZ1cyc2yNUq
aRw1e+EJd+Gz/BPTIzH1Ut2RPi4kXaI2717dHqRTOOnb6iD2+wwXKQ5GX5vfw74i
+qz6UWYYBYXl2RPUNROBxU0ukD3gfMO9vtlMlcK1JkKO1oIdijzSf9Mn9kQqa6T3
9mX2jLc4TOUlE12xYjQfMKrdN6AbgKson/ZVC/mL8PgWtL7Wm1lkGqfPC13YWssr
nel52H7ArEL+kWz8u70MQz04C9poPuMRiT8+CTnU2jv1z4tII+/p5w/pJsQ3Ybuo
/ywHAmznTq2K0AsmVEgG/okCCmvilp2xFRs0tA3rO/VfWaTq5JArJulpMlC9i0J6
zHg0oLfmGDAIGx7DJCSSHgZ183FY9a16ecvJF6+De9CnLoyFMu9GDGlyQgIf+qRh
mQh/Z62qn7ljSDyjsBTuYFcaRSub+Kew+IKaQ2SUDxAgiUOibaGYtFVZZ+Mur6Hu
KIwbcWGTE9xgNCy08FI05kaZxHM96IgS9Vo26kZJCUznrQVeqAtyIFtYT4MNihWD
mSPBYXQs2HytgnBYHYwn0qylko8NZ2RERlGN7Q0zYGKTmV0pc9wCZVXso+NWU9kU
PyLW810uG3mVboNuwEqc+yVA5OGm/k6YntRelhMSBH0AHY/0Z8TBcI8Dw8aNLRBy
pYY6uK/dESm+l9+IF/mkrBarqw7FRz5Uh7C5kGEsdqnMqauXodfnHY7GnJG3Pt2/
q5K8NnXWAdCm3XVmSntazvUa4dtX2ESl+6OfPWdbY59Ita85D6d+kl+BB612+8DK
PfUcTv0p6GMqoaCFkdGMFqwjf5kJy/MpU6TayEPbPOL1O2HZuT5ThFrJAUtiRO+N
FD4LxbLC/ZuF8uQPrgPuU4T+v91ajoUw1reVuteOAsWGuMpb0+Y30XbJprwRbCDv
ETa60hPpMmTgzuOba3ba7lMtMszHCdSxU8xKpA6alF919zw/n3W8zFVNeA8kQwWy
Rsj4BIOHSBQgfPwY8NOceGBFJ+U0lqHYwMZ7KmCqoBwz0MzbLwhT+2AQDt3Iit+H
5jmh02lksOmWyQdnOP3j372pVC9/GFWZjEpK5ArH8zrwBQr3q3nOtJPaxW63Nsbh
eKDtX9rb8h75/D6uO4NV6oejVADXi6mBpotamlG9kd77e5GJ1JL2/Z1zyuwAc9mX
m7a88lJ48EPunIsfwjcY6BrehRcFCfib6ilqJ+73OmDJBEvPblFGRqUhWkpofX1c
EcGY78KOHMkImaNaua9/tu7tu6gkVtXaFLfOPQLqXhSqeDXvVe3twPVIaZxKd1st
LwXPnO9ztZI7aagHPUWD7B4W/xlCv2NC2xt+8mNeBSFOIGc4v09SbpmP5Mk1mDqG
4j7aLWhZey0zKv9l4bRlFqG1MrE+fIB9vpJOCJekxh7+P3yj+/DWnnPg5wSVEwnT
x/Sk4bqJmXrGcst0WyU9Pxdkf99fFS9dL5BUP8Bcx09WB7tXgmM4htecNUI8ROAe
9Ht2T9E2ofrDJQzyXDrmDgfOhfmCikoQKJaLDtwzsgGgC2GGHPQpzf/y7vUcTCQ9
EIp8fibXLhsxOJgG2UTc0/Nkurv4xfQueFFZ7+v4riBI9oWsQlgt2idDdpv5H0BT
1oxAZzDjYX53DZGwUUumGeLiby2wVZLw0nndHN2s7PW8WyC7AjxEL01JL9w48C+u
vY4rKLF5mk8N9WsfwncF/wIRyZf1qX156c/bzqwKKC2j9cyQb7+g6Zpvf63vX17U
nfcBHbrNbk4MM2ft2ScgkSIVEbVPEGQjbDVtr8RHZc8BWG1WhjK43cMOfPfBApG4
aWCX2BR3o5hcI4ln0EawRlzFuhC7q0tL4coyp5zqNCAZxu0TniaJC+nhUehKiXqu
OQCjmHXu0i1EgUXP37fUV+6ZvkT80O1WqtiW3zMZSjwgk0mIt/6sUUD2srHIVM0u
FtZ16Zxru7g08LSqX7tMVTas9tm7G2I1KyJQQ5+WHlgCXnVbYMibO4gZT028OwpI
ErqcRdRcWrbz3fy1kYFyJdApW2zL+EEeeCIrPnkjHm9gkA8oh5/HPED6JuR+q0Ua
LWSEO/Xhiyt8R1MJlsTVp+kJxPfDER4vsrWCxqLt4YWeR8j0zHlWWaOVz4X/ItRn
P3Q0X6wX/kXaMjzeoUvdILCr5auz9+VxQXSkzPZYV7LdTaMWzuJgkBoXe0WpJN+K
EutX6jNjkhzGI7sUi0wCGv5s6+7WCp1gztnCHXlfgjc+R0Mx0EzXF/sOSVsxblvY
qHUsgKEOkyVFmBhsUBkEnMZUHdael/584JNWFCDec0iwwiWd1JlN7WAewv9KIllK
IsRn+UD7T3SvD0v4C4HxwrK0SQpisVrRaUvIlFbUTAdItJq+W+Efhf2/Wv0wYfu4
RLZG8YgnyQxou/VpD2FK+hYiARmLTQDumg+rNe7gYE1OqihZ1OtP9U8WVb5FpVCO
fDKRzoAnugLySyWaPtYsNrB8A7aLjFj3T4qCRDaychFBE5dz5uuMOyeuNin8UIGy
fRWqGqygJ8/99jal4uo35vmNUsqQHIp6CbKfCjx/xryynAqP4w+Fu35N0Po923Cg
KpXIlMvoldNPByc9T6Rp+Av0JnTq5mjv+iXwDmZhUvtPg0H4LFm3QSCqCsQKOsY+
kXSaG3wFkSn4Ckkx7EF8qm4vCP5qn8Y6ozYuI7MJC8e5vIH0rpx5W5jJJHjMhsrF
Tu9J48KHt2C8g3tCQxxTSNiuC6pnVa7RPJ0MK9a5tiHICQvaAXB1pVAOZuxjsBVg
qdfST5Xvs2Z7DndDwOlVl0qmO2/9nu0PrnZCohlgN1SC2M47RBGWcNXV7wcskIln
6LqGmgQlS0q+SOwzGo+cngMsziDGRYDLY7aP9BSMlXKL3A/4w4inOsQbHA+tR2Vl
r4XLyCzB/BdWZ9gBCcyg9YDt/sntfKSH1n1ck3mMBwvn5YKI9ZkwtCKZTF3Kgqoy
tJsgtgEsuvCB0miBKySbWWO9bS/D3JhGjCgqObWW2pQZNiV9A+UV+HqrQEwRzA7d
Tay5X08fYGYdooZLgA0SOM/WJoEdHSNcQjNGZkqa+6nEFFWcIEKI+/yeyngcomX/
HifY/mHY2Y2SHuuwSQisV8aUwwVb5LxSGeD7HUk4eJZbmvyug9mow8nSsiC4A0qj
D7ZhZr/+FO5+G1H9Vvmz3aVOTZlsnPDJUMdPso9K1RAjN6gfINObNdL3UCFxyfOO
56eOoyjhfZzWJ9GZdJzfDTL7wB/RCImGD5OhW+LkrnUG9RQOdEwAFxu2emRH23bc
zgGjTCJqWpZiJug1mNKxIwNZ2K1mb4FACrn1LfGjI5yZTlsbLF9qxphL7Dh2/kT8
kNoaDuwrfovgWHiskA0coK31Zu8MAxQ9Hqh3ebvFaVRg1eG2ULMnIkqvlvZxVea2
Q1AivvbHt2meUnX2HV3+CtNdZVgnX/8sIgkBdHfg73/jJhN3uAldgCuxW1RTZBq9
dDcrqhIGD9giPXRtve5SN3qhuupSHkBv98PS3R0JtyMu3kSt23C9VhvEsSL0PInb
WiKzOT2NtF+qyxIk5vX4o9G0jY71BZss3du/Yge17wFDKX85EVSjh0zvVxlD+53V
ct2Q8w5JpJr22nno6uWVrWPYUjMuBpP3yrPHZjpqmbteMUd3EOyCgT/6M2yqVKcT
5nWYUOokA5iqQSNo8yVfthBB8KhftvYLnxvTqlUrJgJmgtVwwrgQl5cKh9P6vNoy
FAu76jp3ilNZR4d2xuCASRwqyWKD3OYSRPHuozyljXB2s2MJcwlpLhvn2FH+Hvi0
JaJtNBSKamd64iKIkKn9K5RC04cBxaOj9696rI/MhNyL1QISV7gKEttDxssftykV
GkU7hzJaiqOrVNH2XJ1QS5JMSbnd8//29j2YDiKmRxxr7g86GSvnSH/2k3Sd0Lkp
ABkJVtPsTY3iO8T5l8a8509wza0WDrHjrNcVCkvgVNIV3p3sa+N1IuezpfcchNVq
k13aNgRq3o2bfqZch3ShZ3ovt53CuffEWJDGn+1V6BoR38up5wI+V4m69+VbzQZe
S8+mgbXVo0hST7op99gWSfRETszKeKr410W9fvdXruIJiSN3q+ACwpUEq01DtLt9
OCG3sRnkT71pC7e6oP531yDn9KtX+rof+CBtdyv5t6XvqOyXe5gCaE22n+rFtTVK
BbRnJMNbVlZ729uXnKyFEOnOqCReMB312Hh6hOneIYTSFvf9H4xbCFpRV0L1C1oC
OQuB3/K4ajpWTCc4szpbJijoeYuDZzPYNSJ39ySEys3QoK+CtBWcdB0Gb7fUHDws
a81qBSI3V2wG+/NVgux7aO5WB/sAJ+7qcoV8mwnhMTRHW8ypXNa0sor6sHuWAzxy
M7zNy9XaSFJBwuJMzoDcSc6JkHmADGDN1EMVtRRe9Cn7nY+zd027SpjqpNnsb4HG
Wzz8r7OmNnpRQV2/F58GljwC+3OTs62XgJJmj0uzDp0UqMxCIRgaLjLJZsZXP7+7
UEQU71MghyvhCUA2e0TM0MQchqtoLNW+/CHMcDda/QYuTNUUb/FD9cY2Zezj6+4M
hF2O37EYL7xwSLnIbw4r2aXeyYhkBsAM8gY7coHi/cCwqb8M66qp64ELdskeygD0
e9Tq0Dg9bQQuYPnCQYVJ/BMPtgQ1Ubv3wOt5nkqRVOwTOTburXir15uLTob/bmkT
vQ/iWrX304oENRmHStKVeSCBTIJmGLey3HcHGZbLx+rghtThA84kZzs3/Y5wjwfb
Z6sdL0rmCzQVvKd60p553FI3hCkBFlw68QT4gScTIrVdj81zelgIpBOi2kJBDwmD
uTGyMR1PoCDIOugfFXL7I1tGEf7LX5MGAkFAnVxmf+2+MbiEkngcZNwnmb1Bu6AA
0EqQVSx8Pid+5uyGBANaALt+XBGG7hJg3BGRWe4QhvEU506BVhvgFyDPecqXKhSw
MCmqj/Jw4cxHiYgmBOxroaHzt9K35KxKgvW+5wI11vHed55+LgNSfbNDzJ61o1G+
zisV/YsIbQavk2gTmNhpnZ52PfnZmk7DCLmTuE8JM2GtnRartShmsdmeBNiODgQo
Ev4cFEUJtcLPC9h0MKJe7cjBtS3H05lNVFIlpyju2VSUVrfU6zCJh42c81L3ZTip
m+Wlq00d6Zto5rI8lI+qj2JdKJyq8KQ0ek1YcJJeiUYkFSGYyujV8I87W1M2dWC6
KQv4oDRItsuF0mh8hKAyEQpkoWyt4Aj0sIxlzLfdFcbkxIhiA4LQTVoXbrzrFX08
LAbPeOZ1+NoSSUYWZ+rU64isZpvbANRE8FMmk9uFz2YJVbpsbLywyy0JRXYTITH7
kbjPf4MMxJQV6AwN0g7/aolphjOG48vVu5t6uYUHEltdHgm6S5GmG7De25QWvBw0
9kyGtBoceOacbGbC6kl2oKpV1kg02m24X2qK/WPu2XOnvmdcKcv4YWFE8QPVNOXr
APx+OnYhQ9fm3CTjMZzfc+pMzdF7by3TyvYZszJrrMXqX1pS4K+yS9ZK/9hNPN82
NAFi49Pf/qFd3r27n47JfqyRZykRg7W9Qmg/N+IY/F36CR5+VL0Uv6hZFrvHOChv
MpoAI+gxnXIKB5Q1RfZaPe5iGMlLqy0q1kw9SKUgcElZJxgPAaVaN8ngFvLvgvrz
6I1Q+mNOvlBaXGQYyz+Egwyk8/5BpSWIcbRm+xTLNfHQitcuEWeEnn1MpXdL36Sm
y4hrd/WkuYfquwWEdQYpKMW/Ec8ynQF1qzvubXdxw7tjDsKmf/4y10M8zJ4Y4pO2
x2xq5IHep8ZeRJkCaY1pXhEc/reELatmlAvp6tSeKKTRxZH1zdBtTAmlWn+6Yl3/
51dlG7lrdunOugITULEE/MNAoJ1nemGbTSVaVjB7vnzJDHpBi6PXFh7vWOgadJuW
Zy6rimmqm76KyK6AB9K2f4ZUt9gLbxQ/g/KbViSClEEnf8m8QQrcqEKyEwrwDovG
gCeH2aVVN4mkbmaB/BoQyAxuhHg31XBlUI80QMDX82PSJ1ST9d94dUKyZnVAO3Ss
YmFBodbvhlnGda9jms4tPYiapfJJKeGE21XNnugxOoJHgTgYWKnd90k4fV3U1vb5
GVr4xxzZCvBjP8bIg2nlqi6mw+ocInYTpBEYVP0iwxU7N/mmz0LawRc0H23UB+yx
dCdXkHDOe9hPGpJwGy/o3nPwHQ5F7gCcDXYX9VTFjn1t1I4pmNZZ6gz5kzJ0WT0c
qVJOxWkTV2xNSdi6W8GjuEPJOJh7eDDLiY3ZBuFFxi8fyYk4a9ZbTwEf9ka05D9V
rYdMOYA5cG4JnO7g02nub7mmJ5GNxnUKsbDgZxD0Hnl3X/Rk526msMDTOypXEJIW
122zKdCKi4jB2J3kS0PkaafvnIgGW2wasguHfr98OODKUTO8GZJ2KRmtkZ2cif2M
RwpS4G/xKFe7DTEZlmBS8e8nIRTAVhwUSJlluIeSkKndBoZk/H61vX7s22Q/S0+g
WTBhzxud44bNMDe52bwwXplCtqJu2FK2+jbNzUjx+bzxGehZ17Fjjv/WxdHnkT0k
hrNajB2Z3oT9s78aXPneKuqC+mC4QkjzqGrdBkK61ZGgBekCCrI4konIAqPInKkm
0F0EDJK7IbxRBbOv8kK5V43dJmM9H3McpNvbxeZ5AzgU1erxPyvHFQQsk7w19Phv
hb4liBDsCldUir2OXcveNF9apCS+38QZWySv3yutZyXvn+0gJPg6W/YVCerTFrw7
hoAnISexO75M9pIIMHsE0H6oeQgraqlQks6yKVat2XBSw1m17cTEkKzXwtOFUDl9
ptXGPETBQMsp8wMllt+Mak6PIW13W3Sx7W2kBEme+rL4lwJNx5xmx33OvDxRR1w3
EiF/XESUolqv0WOThmY7T4jKC77J1EOphFn+VOAzOfe49rXAIB4MEnMgJ0IBUMnU
ZtU2I9j6IuuINfIR01/g3PtgK+EVXpVlXVRGWGTsv5i7GOhXEI2bBvGFqg42yNtU
MGsiYRtsc+ScaKvBt+Okhi+j8DwPgxXEWsFkggs4w0rS8acS4c5poqPihAv5HAuH
vgTAacetuR4OtXJQWpHlRILxlwxkyMgAooDuSD3e+lRsWXc8VhbYzLLWE348ugfL
WEbuE7A8xXw1KYaRIJSWbdECUxQDVYByQX+clblpOLHrWeT1OT5yJO3nwF1yYVJ+
h/YKmYbPYWMQA+GuONGUZme70yNgZ3FrZAYsLCptmi1xopl7rJFGLqFhx664hChq
p1IOPk5rPvpVB20hNQ0tkkU4rctJ5MI7MbBvzj++WIKlGQrBUB0zU1RMHxszkZ5t
IivWD226W/sFT7jew4H3mxMIypYH4/80Wq6b+FXSjpzvYFm7T0G5TCdYt/H6lwG/
E0mxt3L11Ggv7mugWDpwHNy92xmZPpbMUaIUBrLZSZHu51VSNCh9TJdftFlt0EtP
uglju60rgS0X9LbUL1LlzCVEMhFoTkUvlXct2W+67i16wP61aEFpnZkLep+80QZM
4ERSXzMM6fsE99fkPl0uuqq/trc9Imq5VXHi2LXo/sCxE7D7lm+C5Zn9EH1TYZmU
H8gHmv34El0Qf5GWDcX5fQBTjqd7c0CMFlQOsiYaIu2HgbuYAfADADofcgduUGzo
WQHfDgB5SL2N4DHI96dl+QhZgKvAlgPYLrUcVLwzMxHQxMcRziHMX8JX5QCJNpaL
cH7fxvcFcHeOGFf0ej100Hc4KwClByb0uvPuNNG8LnJ7ZKFsuiQVVdSlSO19x84z
3U7xM5Qjog+WiKCc/VbBv7hR1k8kQl2wipNEkpM+BiS4w5AyOX6JXN9mKuHC3KUz
NQNpoclMXB5ydTZZyTrGi55GyL0MSKd7CZsXJv8caBQI8FIcsmqZEfykS/Fbnrb2
Q+rsfKFkpDBI9ARikBf+vnRXlO+z+AvMACOoH3Onu1OHJZXV/mstieT8GM3E4H1H
q9newUy0Rg/y0nZ3okqcR8RC7s8VYbmxbQNS6Nwyw8RSWPAk+Hoyr80jDS38TMR4
Ag2VnC76p1WGXJuPqXdkGIlpD4uNFaVrySxzh8pP6UDgYx7r/+60T/0BA/vIc/ot
dJtlFr81aik+1QCJh3jDG56ruyj3+E4OKxKzENYL1yfBsBSSn0m7SkDk99b6279/
9JPmxJYIoCOlvNQcpDGHM8DCEvicWbSEoktdaaiKRjfXxB5k31VKwm71skMo/G9e
RSlHBfujvb0pJSzhJGYAo9UMiOz15rIgozgpwsMcALJEbOaWKEROMuMZNc5wRooo
XVBqrcULJ+3OGFGhQjXxYmhco9wQXWzIn6xmGsq+BWrQ/ko//7j3x0qXaJx3kUkE
xrQqvzUBC4Y/ZL6JLztFRPWijlxLEFkGrRoR8QRUfmoVA6LprT+aJ+Odhdzf/8+Z
aE/TTqDQagVxjo4lFVhhIW/XfKdcErkAo1FT3rhKOOS/gmYrHoTwUNS0/LWtoKzA
U+Z2QHIAsos18ljIqxT9BAwGP1E05JCnOMzLe0DbWPJfkC4ChphmLao9/JIOBLPx
8e/e2rnRS4N/Rcw4KrOJIMCDY3fLjkqztjeaeJS80hGK321GzapnH4+qqCD7+uwN
7edoABqxP7gmm46yhVDDGezOgQSuv06Q/NikfcmYD0LUuhKhb1eJ4NSVr1C1UTju
I97mcQ02F9aYJkP/ReBx4upInmWCHh1HAjFu4dM0A9JQB4DId2c/Vqa9rUmFFSbD
UdcuDM9FsZXPNB60Xt+3bZsZShvJbrsA/7s8mYSNEOwRWkfbq1Cvrzd7yXdF37EV
nVcIqLCWKPmUOrgPqG8dpUTaaEZzlvjWLsiO/o4L4l7z4nAtOq2ZwwVf5HF9eitp
depc63TW6AjOLFGYDs91E/pbkus3D99DolXjJ9qgHEFF9UReoqDwtaRUDU71EJ1Y
yLJZWUn0GmHirv0heFbDdZER24/57wLyaK0eWB6AKR2LGSxEPSDTRTdFXztpWBW1
+qzfT+QnsSqFoIMjcbq+avIju1ZU05xSjKvgUzNRHyFE/Wo3EiF0phxH2m8XDHWT
I3D+uDF/7DoxUbG5r3Qfx2efOsee96x5NDjoEjjOWCi0PWzy4OldYdlsKqU3iUUq
aRkB/bRnIoZIpyv1RhpDUL82gKhbfHedbndmolYZS5FvtJOF3brQOA1gauVPmEBR
x0aqVbabgFcdxzxkUJWOx99HYcGC3Gh1+6eg6HCf/o72j6linyc8P6qAPk++4evX
kh9jQCLTCOgmi87g/Vo8oRgZNFE4lhxcSYTHv6nyB971Q0DdwLP7JHS8oUPmF90z
uJHSgheT1Fsq/W6DYDYwvIWJwynpZCbhpoEdnhYVbQV4844oOCJSOCnnsm+h1rqg
DODwbDveKd5sH6ZQG9lZCnAKzYDzA+ifIwqiWRsRjuwMNbxELBnN+XerY1I2ZIXV
EgCzXrgflyklo3ISy4Bb3QJAI1T2TELwlsnPMtIGBPiBFBPaRyF/bcNHvREVSquu
S/uhX1P5NRQce1gxnC15R/8qB084vACx2o5Yu2WAa6YTS0djQGqst7iY5VL3RI/m
IGErM5Xr+Pgf9QTVoYWcaY6+y5RVBO8IfCL83N93FyenDzlPuJR/THY/kD4KZ/wz
3HqTTia/jpQal/s6q78MRIgqk+MTkrjkG3NDCzRg4yW6MYx8HbqY2THEMd0LSNgb
XZebvy++zKA0Nuar+N28pWWR4TSyH3IIxqlImMPIZ1kKrr5/dD5Y8k1P5aSH4i9c
DcNAsf81M9VEdOGu9F5031m6OIzIMxxROy/K9PM48vQQucqk1QEPMEH2iGACMY/q
C4nF8F4KS2nLo0WIcqJL4Hbyid6L8v1CV8mukIRtkMPHVgb+KlCCDfYcnjJRAc3C
/5IVJTGwuiAgBXyrsi4kBcgo25rrOHDXQzIY7R2XJMQCShZYTtq7GmLjBxf/KKDe
luNv44SwZB53JO7mfPyNEKa57tRyCCGvYQSjospJ8hOqD82rYIkI3FU0dtzSN5C/
r066HsusW8dw+jpevfH5pE6eUbtoIVfdi3YT/B1nFejnqz5lxBToqM/V4CFhFKJM
vbQKEMzMMaKNySC/M6dJKsllq8gCRfYiFiJwBgl2PZzSMKPZsLs1fTWUAEMjiFuz
sHMYvxNKkLcswUKl9ZoRd11UVj7711H3qThbLHOPUY8bXoyRymLTVhdvsQVBx6bp
FLIz5MdTU0yGWJXtrqOQweVnIEdulgvDD1uUqceruvjxNVKYjGdmbCgDPh0ZUGY9
wi2I5Xmn1qWZChuJgQwThqsypQNLwGo6sS6sbq9ukZxtFcEtqVV5YQ2rhqS6sBcn
TfpkN26sXcNrXXGpD3W8Fkfkf0DoijQ+8FwfWFuM2u9yxZFdAvCCbrEfjKfHK8ip
b8HFSFhK2oO4kCb7S6nS+qBXKMtuuoVmmqQ3Nkl/ZBKCa+Jlfc6fPJEOIYVKV3ny
8RWzMvi5ElLCyrk8PbdeNA//4zWyYhVxZOO9ExyBOw6LxgYUo2bekFiYudx+vDgN
FwDAQvhCaAzWH8rNO8XRGWI7eSs8kQv/1PTzgu+WMHsjVhE+VKDCttYvJnr3f3PM
fHEI9fCOIvDlzPutmddaYzKsHMF55FliHMuVdWeJ9XOn7GEkOzM1Ays6qUBCEfN6
ej2gXmfCKcUgi56dNaQMl2CogzgtcTJ/+stsIp3DLk/0aYNBXQyTRr8JYbE3QMfn
E9hDo9BFZwVNN3SEICHlQG9jtcZfMyLca934CCWSqQStHdpCU64KlPZm8Lo19a7a
AnZQB9YxV2LOV9pZf9o1EbbOs+L4Blr/cvudzJZSxZhkIZuIUjxCkbbkkKAU6cMc
LCORUe+GEavDd4d2Nc4DXRV+L2Mosiu5w/vMsL9myz4kpV3ABTTDhQXcEWmBnnWp
wjYGzI37JPAGb1ZrA2EDPW95+HvtzMOVJ4AwXkD+pmJ1OocmslzDy21Zeo6xHRJh
mPJHO/VT3dB8VImu+FPtEJN+d2L/JvCFOLx5bd8KHTCX9Wqokj9o97KnMiYTAMLW
K/VZ4hHwcxeKEibbYwinYS7fr68iEK0Z3msQpcGwp1ryQ0UFy/JpFDvY79gu1J2K
V7+PC6cyHc+TDcGWoEkIGzul+aprbx9RzhHQc1reJ3gEFyVMkRvJP43LAvjN1XnK
8jTi+y4cKqZN3jE4CNboFCtrvozoz4bBImjxv0U+dr2Y1m9KS8uHpXLJ5PG0EI1j
Ncg4/w9VULlQ2iu9fL1SstjQkZEfbketkISzN56TU6BMZea6JzCzTs7bFdUStgqR
uNqa2joICS+RJBZAFO3sppwsu/QDp3K/xnRuDB6xeclgjuFTZBruXV0vVEyu0p6v
0aApgxVuVpIbP/3SpEWEome+9eLplwrv/tLa/qIx9ussfJ0XOh21k2VwSWv0AGbL
xCZeGXJOgM+0dKtp1cYRl4vlMbF1v+j59es+zd0rOMkMGYCuAxtWRNV1KRBi3G2r
va8Cijhoh1aH9Q2CD5PfmjZDBk4GxBr5/ekLac/qUpcrXZ7GfTwsUE7z2NzyIxcX
5EMkBIV5nXqe5Oji1lj4Y+23rcIK+J3TLgc/h2p5J1GoigvkTDNYAgMUqLn3rhyz
elHdy7W9UMPrKulm5Lc6ZTi4DtGkUOZazdHCPwkTlJ2yiSRuS4sAGUs7ah8u75Cr
F748DqXsD2K1Y9rJBSuE0P9wGKj3DgJCWQQOOWiy0QvAQwRRDxuqfGQ0PK7kc+TW
G0+QgDaN7cVVRGuTGiCLoUmryt9fUt/tHHTaCclSNOxLnv7RLD9qu9/98sBnHqOs
v1G1YriPer2JM3jCnzAmcw4i3zIWFyW2WaJplgxkffDi7hD1SLhc23LQvs2k6cu6
1B+IOvBYakg9Xm3cc43uewV3oKHNNze3Lu3271MuV6zQ7qS6uUb7Hyxw9MCtMKhH
ZYo78xUgUxg5bwNR/faT/WbVpuqdM/+ySWl6Wqa/9+KlUFhd+qmfVmzsAjVD+b6N
4J69HTHc2cJh5eCS73qQPV50VlP07DFKPxHTEnBRJNM7M6WUk379KUz06wRBtc+q
2X59OkCaAjWZQ0nSrRSVLxGEFgde1uUDqJn1hU6kAe+X1EY4B/UGe+x9+CyQnAG4
NsGW1YCJvKM/sva3zWBmhA0mZ11faZVxjh0puL7UeafOQ3T9XrDW5dVWamerHNtd
hSGSBSa7rN7TUKWvLtrK14DG9K6CKnk4vXjgQv6hr9BBghbcLqWEPEXkbU4V8mCW
K0KdCq6lYBDfY6YdHHUM5CFvDcx8Epn60o57t0QOENPpQTutIGgnAbipzVoRYG4G
6+NJDt5HM/zMCp3jO4AQi4d9uOZLdgvdm2d4o2V5YJbv0UYT48pgPxmfnyzpVOsO
z4OHGCSHURTqIART/jygi4M6p8EMyUCbK7zEfkOBi5Ae42CY2SG5WxFA/vnhGkt/
R1R8D1gqgQJz5hMeyZMIV3rEZWnBs9LTucWnLOHDyscUg/TJuJw9pt3gjhVF/2ir
lUSfS/ERRlWT+CoK6XkSWpxhVlwZEPlhAi1eXzF25Zy93kV9JHFjfhQGbgn8v+JH
83EDZQiWlwl0l40uzLP4esqYKxwK6In/AHf521TCzZjvDDDsFvhnQF+R17avPSO0
yTShp4SIcnfK8NlpSrer0NBbXJSdPkclgJX/jIe2FB2SmhyxRVcfHqstRRBo/NEW
Hitl5FsjjfVuI7Efk+NqRUvcsTY9WAwQ4lGTqPdCvRlahlNdKvFmosOwJtjYnr5G
x72n2WGk0n8T+pT3HtnQ2d3RIAkyw8WSrR9TjZ+UGajeVx4IV6fA+zP1tbBM2yQ2
Om5IAwCEUEHCUkAB9q7mJv8GIf3nKMPB3jfmaD3hh0zJBSdF9f2H7tLRrHiO6vv6
/hyNbXu/aVxPadHb6BHN1DxKoVrsAp7KzSyeLi+cs5LNxDVPrA9dAy3Rw+zPlc7b
+Qxennt5S5DNpgGEwzt0p+66xTjUMtMNtHU6C5JziaBJ4+Ba9nr5w1lNKR3ztceu
IPvvZjAyjD0t7FvHicEgXB0P0G956DWCYlYkdu/htAD7J2zZG2nsGSfim2r/uvGX
cOeAHbHBzFFhBi1hQMh0uYka28sQwOK5SlaFgsj3PXavRsMCxpD0NAEQegcQuyw8
oP5S4jFOQHd8EgP3QVKYo7zewT7ucfI/C4yxvMMb/vW9barM3T0WXhqEa91tgvBa
TQ8cV+WgaFwN/0rSUd9QDPid85za6XAe1MOMh5SXC5VkTvd/GiHDr6r9YaIQF9eP
ty6jQVtW7W1sfBHHaL8R0ux3r3aJ0XJLxI2lA4g30ydwWs7ZZqjLqKysdww5TLSZ
JkCnc0IguI7ipVImDp54u0qpU2kjMkX7GJ+otbHFGcRC1TCu3gQsHyMAv1gWuzla
HBwPQLpfGpfmGmGMnJBf1w/OVyUWt84uX/XKJ86Phh74lc25DFaZmDqIS6whZrtV
pmF/IigMb2ceC7W0nsffgXqJPAN2u5d1iNbv+CeU1LZ8LT+g5vRkpmyBHBle+QzR
1GGE5drGBlvDxagxXDru40k/iUAbmg01WU+VWKPmzy+5RrXREIIuSd/Z3xBLtDMH
bWgl86GKY8xQJEHmZ+g4ra1p5NK0E/lXxrhICRYNOSqDpHcsIz3XEHTecIbAfr4h
YKxwyaNlnoolgeCai7Nf0kYQWMFTUsjuZngLUYXfK8cg2Buvf+cUAgM2vBIjyQoj
41WdXQE9/OsCIV5EFeHN5LtFrThSTWT77+pq9XiQw3YPyAnyR2Ui0tTV1YE/x+MY
5p8GGlUfcr1oh0tu04+JFuvScV90aRSl3zeNk6raZwThwV//PZBixJFzEKXMT+JU
ylA8vpOixX34b0Sk5MucgTWK7WxxLeMq9+cQjDUhx+UgFo/Zy+X6AJp8xqUqRSOu
yBSFDRBrYHssub8rEn8GJ9zOj3Z7m1RSqoHLmDll7Mn3se3ajNJeMl+r8YqXFhfq
c50564BI6zsY5nxVGyyuU5p4aDDguNgfQp5wSLAl2DfFj9SkYxFPQQlJBezZKueZ
jNUreB5fzweRmQDteX1hGmARA5cOU9ApoqLId0h1nFkwjHZ5LvI78myqCvYPdVxf
8rxi0QPnrutniA4z7JuEnbVQkOohXLZvMAsfugNKz5JXoYKES8W2tYunxH2NykEf
kyIh2lqd7Wl+ySLWV2vnbcLjZ5MkPoTHKjE4Ssq0t0ytUM7+n1wS3yF/dG4cBllT
72l7v7iSlg5bFbds7jIWvf2nHMTNOJITjnamcIeSFbq/v44yhlBxbA6ycPzIVkqF
+RmSNRQAw62B567dq/8oYmBrULHjzs+TXPELYdwiTIucPR9WyKBP9RP3cwX2ze+U
TzxNuAXPH6vlUYRMpExqS9FrIl49WN0McrqSvKLAevOs+8OqT0/huuMg0wgXjI+J
6nz0LHLLA2nPoX0yxE+Tucsvv4QFAgtokOMebxWtkCxng00CY7+B/JdgRUn0EJkh
rbvICYRhiHzjqts4S28bYcHBeC+1j3f+V7HIi9s/iv59zIyOybznwvWlvtBIudaV
Tz1OIlSx4LQ4xXNUIg29fsJWU0HAK9nqqdU05Aee/YL+W9F3h/YDLjHOdPzaGQxi
boC6RAbNGIvTSdW2IPNMozLhvas5w73AtZ7tu/TpJjMVsA/M5zDQiqR1hJ3tktez
hEhBDzbs2O2T+O7JdITAGSDU9IfH7f9u3HaRfvG7bvfcUdC91roN/MNHS1vlLP0X
KoxPRAOX1qslOBxzlm6i7OVQBuITeWSer6oAmiR0OB1WuniMPot1FAf9/Dmpqjgu
tAW3OgOqh1ctEx7VCZh2WRj2G/RZbp0Kd9wAOfjFDxrKx61cjapN5xvQ6cuhyW52
WzLVYX6QRsHuTyT8DrDsfqf+j++AqfxQQbyL7f30ATGa/VkLxfSnX86jeAXxiCNY
7p4IAWSBDRi/sqBnv5eF8kiRL/xBhEZfddNNCaEPuoHYi35fm3IU/3n8y+cVTot8
3VqMsmXPettSOUqWt7sOBX3T7P38QlRkA/9ND7/UxPNh5te6teO7JTjZrFQUiXl7
jFOqwlwT8YEbM9T/XJZuZVZg/RQ2v0DXRLgH6PvxqhaAlsLvvYsyqqGJ+/6wyK9y
U7kmkro7SuaVNeP3xdBB3v+6DCEBBvf90Ly9IsT0+Nk/WSbC2hYWpTYeFGo4froq
R3dMfXIIsKirBkVe3Q8v1AeC69WhSqkx0cqKmfSnGPUKSV2KogKUE0qNysvREtcQ
O2vXzxunEUc+EhmvFt/4Qi9iagBNVMZXJ5HguDEyCuOcUR5YmxUi94dlTToTSlDj
P9PMdnWYmTO/lwNmiQur0x702B0CTY6MOWROV5GuVOYw6eiEip8kSwfFxDNO4XvF
ETLZaGJIYN3ppEDKzMlKtb4RdJejzeEYHkpIsQDBeEjS0EvbOGRnG1Wr7TcOsoWq
sfhuezmo8I2Z4BMGQYgqazgW9LbjIhoM2Hc83fevCqPuvTAYCg3Lc57l2DcT8fFl
ism3m4xktQsNwtPR9zqsCMpENgUBoftmQ+0EMsG4Qsokz+6j2GEVAADtNOSIvDom
BxFk938EJAnzAmM78nFyGMuhVQ+A2vSMF9QiPdUAhb3O64rK0wa0sXarwem4cf3X
HgZ7fGvzFo8vzYP8XfCT2ZO2G7O2ZM3fyHDcT9KFz8GReplrvDH+5d/Lbb2hVprR
daCra4eq6ICeJRmhPDR92a1xqUgqFkoKoCU+nJqcps1I1rCOcRjpqlO9NMsNIOUl
adGNPOhk7uaOo5AMpjRE/IMEnuDtX7IxzPMTbkHFm95HLdEoDh0naspTuY1lelUu
GNghTnQSBGfmciyz/dFtR0EbWIqK3JNYH4rfVuDoiM2m5DSn9bCdSPy53a+4ri/z
xq17eLq1WVfKHBBVf1S7qSBUVNWL1Dt1Yg8z8yU0zqRfYrZ7b97sSg+bEvU+OzM1
4OcKDxbWHoFWUMnrAoKfYcKCsldoDGfI/O7SI2xq0dE2V3mzNV4E5f+LhP0fNzd7
dAA36DzJ+rfoJto4DiGSYQmWX+Mj9o1SgjY/EFnghAe9uqIvupCycLHyA/KVA1Gi
HTRZUdks5IJUhfP9lmQQFAs+YNa3eVm9imAU6IywuTI47B34R548mS6ubsm6zV+v
USVtsXOzVj9/jVaJxznIdLOBvsyiTDLGzpbwExu4iQqUv+RFM3HWWyo8FLPwIPnj
F7cCER4ZeEwsKLH8So/mmPSZWfLGKVvRcZjYORTfUIWVH+cs0mk1YkawvNTyXHlX
eUf5ZLqQt+FF0BRyDWK1aBdQG7qSY/jGoWNtLG4p6tdIptS/q0RmbD/71vafPipV
6RqJDnNTGknaUT3eDV+JXO2f25E+M3JeHigWsieDPEm0vvwicQJRa29VudEdocg4
jyoNno+Zgbe0lPgNd7q4Kthcwes1SexIHDefv/z0a/dDIYKzSmlcUChYQMTXQmPl
FiitONyXcq2yH6L5//2A08+zp/G0/9oQ307yicN/9b1DhJcNHjZbwDa6cYIhYBmv
JH3C6G/eP1Y9o8PNfZy8eNfQ2MY8RxQp5+9PaDkcfHWq0P4tajAOJNtEK9rlbqHy
w0TGz1i+UnnAlSuIJqXdcJcVUY/lvznhDorNoU2g5vxibJgi7jGGTDE6kPFu7AL7
J0JUOfzG0teWXT8Z109/ZklAgjLhBQgil7cHocN2F9i/Lk/WxR8YEOMw5NDFiEJX
7H/wPejQloAaesY4tqLNYMIiQN59MMgUYhJ3uXQbQjhkAHnaGhyRnikf9RPkfbDZ
ZPBc1fVDARtvFAR1SXvNrz7NuDB55QvWDKvpdN/EiBlIQvCVHPK7Gw0eAXsGHMuF
kFvK2u1q57fVPixrOG0R7He1YaWCVJI1ajEHitwz+kyf+P1pLbTbqp7ks7tMhNH6
71cGaij+KgEY28a7uf+xt9uYK9Wm2V+LP+1HYbw/6vs9bG1vfwkxqJww0p8+QKUG
hqLkEB36/m9G3tPtEKM5cU9eljjS4q32TInl+696G8qKbH9aHPg3PKgc1zr0DPk0
xHjFmuqjbxp8sjiEkeLYZGisUuqZmfpbEpaDLOABLJPprKxGTvS2Qi5jloLd2TLp
yje8imiwAdDvbvxzLoTfpb9cR/CkrEU7fFY9OMGBi9kxGtmYcoBE8b07Wh2n84ku
blMeYJpCeg7bDy0jYlQ6274P9T6PZY4ewCCrcHz4D08yP8gHEI0EORoYgAPsc4xQ
6qpfuUXTMOR/rWFFR99pwcsveqSXgnEAQHkULMH4PSdWFuYKdoo8cBD2cIX0i2yU
pHDPdssAtnvw0o89cEfJHB1OeApAELt1qgLydzwP50YnhjvR2AGxoUAVBD0ep7C0
cc6dpGU/1oEViIFi14eOAbbxPUvWHZ5I2iZlqyctySXxBatImdf8HZ4rMS4GbpdE
h10qIsEqlUTa6/LaxmZrS7BYdRnWGw11c+cc0fisLh++bAS762ZEYJXIX0npRI3I
2k9aEVGcvl4Rz1dYp3YfrEF5ryDahlKF7/1x2nn6ERS0GJY0/EUwq7DwvRQL1kX3
hnzpfNDiMIuepiRDB83ZRmRoQukdjyi2grJHVDoTvWBRndYp8eXU6c7UBNWPy6XO
I7BXMVA4KlrqYYcD6Xd1ji+NVBLpqqOeRMQ3AqjMk0IztV/KiN0OrV11quXvl7OY
YEBrh59nKqE3PAYSTSJ/aL1KnWx+lJhRnNGOkgAewQFwu5FIAs/puE/m0hOG0YYy
/lMlj+NmZwHr0hJPGufwuK7cpPfAMD04eYo/c/z6130Z2bhLsykjjM5dCAbTQheq
tv0Fn+T+GVva43mZoQSbkKlFfHIEyBFrgq5WsKR136Zo7OWPsFZI2HzJ9T2R0Gfh
m7A4UZ26nECq+0FmnolnDnFjvOEFw4X4JBmZ//nNUue1u0m2Yo4kspIb6JkOfhom
31R3KbSkYIIbY9+sooFd9/X50/QwGhf1NWBWX91ATD0ngf3zCweidjTBxbSJ+8H5
awELnUkCFzhPYN8QKLLEqs4nNHKN7d736N5JlZY5A9IK0kziJWx3SIe5yoaoh0tW
2A9OtgUyjIrPB86ODVBrPT8cnWreebGWtIwAcpv+B+e3zD1Sp92vRXvSOv/4Jp0a
QuZvxjuf6iHi+yp6c6DI3LWEKFNQW3nH+vzUyv/r3Vo73+fRfwnOfzflBcsgqld+
zkcchzXbjpfrksY3GwEZ/yJPBajXPqbSLztaVIUApQ4Qi8hFI+co6ma4Q3UTcSwr
1vQnZs98f6BH8Buf5WyaLCsPqV8V4hkfrnUIkwohDxURyE5hfRAb0ZrxgltOo2q5
dnlYTGrqygYvTaVoGM9qba9eBVkOSBKWWzgONoDt18oaEM2b40yJ9aC13SmqgB2j
GlK54/sjclD4AX2C9qlFV2Ei8an+ak+T/+16K5n22yfxuDxmiWSWVEhCYe0EIicC
z/fSTjukZWgA9TCN8FUeYL2xH75IjBauX932udlWKy2Cy8/58TwaT20PqosgVS53
S/z2+D/S5hGXDnN7N4APm0GMpEhXF9FnKeRmYaktGe9YhbzKEjzonzAZc6aWhTCT
vo1fH5cFIUs/f4UMVAR1I4YzGVAQM+pfjgCnyuzA2EygGRUtJ63XLSKpsntA0TwR
ZF+/4un9Z31Pr2uHGEAWjR/I5YtGG5FrwY7nl+aguMCaj3KRPz2ftXEnlkMOKOv8
wupEuT48sUMaWZSm3l9R14xMU6Jp8vBke499sDGapcsJfmcWus6/YRciUuvJtvWm
z3Q5qCbaujHmxmijlRVh9nqPHkqOFS1BECkTAXd3JG6nVvaXw0A3DNaB/e5sUe4r
tDZb2YRoxf2Q4OGK1TF3P5pzNR7P5Ccze1cCjR900jqn39gR2l41aCFJLRAPBQ5e
VF1SOApY7YVl029Qf+mLs7mzD3Ut2kgU3u6DhYXoI+WfyCnNHaM1ur/kLRzy7e1p
+Fu0dnX5HQxgDje2Py1Q9M0OfE3MN6xWORZTIk+dIhM92hxwcVVCKqls4vBrXVTH
0LxAcujcb07uLsp6ICWjpFQHO72yYEMl9b85OMdNW1s5ojJlsvtZe5/1DwyC6n9T
O3nZntZvXqvP2T+2e29LR8K/LeNleniHeYifj+59Qn8PyLAoSR1LQPpLnO+opxFv
gjw+2cYoGHoagtH9eja3Chdfyn/nI7ADooHAMt4Q51s72yHKoANjm4ICCDvKDJIS
ehlD9n3l+JZeJjkXTRFgia44S9PJ0DlCP2pb4DvJSwYuaBJfmG1btSche8qAvI+H
9t4ru6lLFTw3LG+tkW1SvuqN447vnOiXgQee0Sff/yUgl97hn1vGtojEraXjMe/F
g4VAVyzBp4cmkomoDLom+A8LxhVOcUvBmxi/Yzi4Ukw0/cwHK16FcSl6i7/wbcTq
3Ww1bO8NgCCc5YxdOIXps16W9VihgIaysCLb9gY2xh5wrDvnlOn2nwZdtfMimOW9
75U7Jja7Woa9ZicllpDO8ZplUJe9Es46zzsmTE9HXgNtxxlS9ln6X7Dhqeguh7kX
/udH5XECaV0IsNVmBQ6iMc0Efh87t3s8rbrRs4OeS+3qy7adT42/QQiPwYb+5F87
BRGtf0pnrn5XbEnNFifEfBnB+aupKAWAeYV7pi8E3LeHAMUtGoCwk60LTGOQQ2ku
CGit51yD+PTW0XAZt9V1KeV3zqU7x7MmskiUHSH6In2qXvJa/M9xp85ILzeqGWra
naVLz+VeHK75vzIo+Hlo1vBdwoio2wUOgVoFcSrSDnORo5SPbIXRd/vh74alboKX
uxstQZxqBVvEkWKjhy87zJbd+Cu3am4CQo/wcD0+llFg3Uh50VoCDwaGY5vEiRvx
XBK0etNyynMLYxPAOt80lXaaP5kh6497Njf764KX2lH8ULOvPZDFq3RA42k9PkRL
QpafYYNKAtomi892YCehWAXcQhNRIBpQllHcI1US3+GUvnaxC6rHinqlKv9ZhaDU
TaVWlRjogIesSLhpUDyVARHW8uKGFyikX0+0ddeWZF5jS3pgQwVWXbbt4oEthGXV
qcVnlU6iHIQks4Vprug8UrgpvBmRSnIH4xrzNhHVtaaVblkPuXc/DjgYdU6deLjo
0PloMLz1z+mDFfziKNC82VY4zoVG7Y5phWumXCcnxwHPPK3Bv6AfV+SPz4OdND1a
o8hbucjTv9uvIZmqbfqIkDxomCTymCDEyYvJy8U46oYUaGDdPR5/uRjOC25oMyIW
qR8/nqngaNAUCRiadBUfh+zo1zPXTr6b4hTtMIsRveDOxHHfbjzZ+nBOgxVso1G3
DnAtbPYvpdQqPYFAOeCGIKXAq5B7fxstw+cO0Mh/BgQFn5/6Uxyn9dPGgwoWl2oH
B9SILJQCbtu8fPvTBkwvBOg6PzA/2rVN8WJdlJs89UNH36r+2n+w1ncnDEmN/mWP
oT5vNdbGPNATq32cSz2FCUG9Uac1vjEuNVU92zxXpdaBzNcUzGeetFrNiO8xMU5R
dPBqKH16Hyz2kshDcGqXdkYpWUY28si3DVu548p1HlUEMfxqhOXjOXrSQOYYiuh+
lOEeR/7ZZmOCnWwM/DRh2+O9jy+JNYBGNrg4OT1dR0m1bfg7KIQHz59356n0Lvs4
YsMlDvWk+X6SbQWh6IZJFaykwO0zGQlnm1x5DQQZX7ebjdvJuGw9+yVhT0RtYf/Q
uextbWhYNOMW8j6vpdfCGXPtbnlg/rtoNLf7IaPCUDbuaMFJDmfWaa+F936Sm+EE
Kpm6B9g3Tf7UpHBpVOsYB3+ACTXibkSXDLqvBWndjubXxEhcpQOWywHgZaL68+DW
CsSJsYCXPNkUEkMS/ry6hCDkNESYSdieS1Mx2kP4Vvnq53z4Zwykf3ZysEZ26sFn
2psAO+sJmKvJSpaA4m8d3/AWdYeEwRTSfz5H5WNoPaG13S8g3O8a0N8xh2AE5xId
72C2FU3c32uW7QGVMDTi45yK4rUkcwBtV/8+knqYmWFQRJJrFNGqApff2RWMEgNH
hyFOrL2ejGAUmOZK6PBVjsd0cPGRXVsO9D556oWi9tZ0fXol94WTvefgp3j9GMHc
IXc7U1PKoNkhIeD46w22TnB4QSyFuRh/YZ60Ux3bpYfUXbQUTfZmsE1CGaq+t/+I
ekQYssTtB+L9rgUJBw36yItCscKn8MhXFgkHHb4KnacfpLYP2ARp00hRDVQXZ09c
AYpYZo5RVvP5u8NT1MmVdOU2GymH2Z2DOmvi9MWQ1DDHekjZcWHbAU7XWkMf55Tk
DvrtJheAoPAuRguqr1ewDMTCKBdsIq1TPXGvtIAHsK7/HvFpukSbKd0N9aYZ4Fjv
1jbAErHzaVquTovc4qkueTHfVgUGHpAguDFbXPyuc4Gt66LtKzqUlXopBQg4hZ0b
XX3cr8hoVdxZYWnOV024Is1Ngpax9Av/Ju3dY56Kc3haOPert5vgiGJ0WmQnUiDb
oulJKz3pRVVUiUPn4TXMf91+4guGTqrCRkBRQvzNDyN7CSmfcxxZ7HTjlQjZuyIw
SU/9Dc/1QXuxTJzfGuMGp0gHh8a7H0xOBnZ5PX02ZI4fRVbQSc/gkbNaXEoNvD7/
70c6Bl1vqsgIfbi1sBmK7qzMT7gMKeFhBpK4ZPXGoIyTfTs5a631/6tZztz8Sl58
6Qrvk2IOL8mkJgRXjs6jLZWn6NDvH93puoTY+R1gGcgwqd/VjOLWIDB+uvdRna3j
3TCM0Gxfi61OB9HEFyLkMMmA7c+6h6pyCDAXagrVumCqaDM95CQjBBGhwYR7RMU7
8Au/lm809dQekyF8n8/T+8gsJi6lgDYw5lxwmt5zXX03FbYqWAQgbMUVgbqemH9J
ZG91TWpUOZQZ6geVL044PJ/Udbcs00mBWaXRm39YG3cOKJBnt0tYCQTgi/7diqoT
wz2Ym/cSUdMh284oMAuXzuGUNHefW3fD2/bmy4v1QY9DoBHxi30PfDyxBui8OdaN
UfUWQfQyNSe905vmhetvpNDyVP/w3qs0JiDv0+F3fXFH8SpWxj5Zzl3GDf80YBWy
cquAR8b4AW5alwHy9z32bL0rOQP21G7TFejRtFVd0YHXCMd0aoyJd1ZapN9PFaAI
YgdtTzQyk4wtL6gUJelkcDkQKmY5M/2K36SH6GkSVjKrldvKwW1YBPM8/xTWYun3
H6neG5kpDDi4oNDB8+TFUFdYTWHfqQRjOnbzbXVgLlZvuElD+5tNxazO8n+ceagH
UYHFc/MIzC2Vrs9eeWcnTCiAzWt+a/8zLes9N0hoMbAih4UQyYR+5HJVbIo3lsbN
ErZ9CipV+QIS9IICon8UDYWA+bnnUPplw4rttkFneLJ7+/d+q2kxQMbFGa6ZNsTz
HDtY6AVvQEH7m5p6c1juERN27nynyQJYO0VRDgN5w6oYb8kV/DVpmgIqrb2gnxdM
fmR1Zc+AXJJ8daxgneRrQMUcDzSIS10MSgypPU6xSZ5PCFW+wZvWfZhvqfV6r+wr
tpwn2M9+UpdwGqzZ/yZMTxugUpF4ud7AEse1Zqzg6C0O/PSjMF/lsUlShI2DrTiV
fq0pYGa5+TEtA2YytZyBGDRP4uka3W+rtXduPf8QzXKajSwP5O7VMbvrgDv6M34J
/9jRQeY6LLmBWujUEPbYJe5uyU1Evc1g4cZhpQKupYtyLKEZ9fE1Z6v3+ffVFgB2
LnsKkMvu0qmP8p6nJ9/t7+71P9KKSpzLaA3uc/9jmX27gkJxm0iFj8BlcqyvgShR
lp6cvzx91LJPr8GYBHAeesdWoamyFyjmAyBRhRAYajxcrvgqjd4+CJXJ8v2GyA+K
POgSUstzi89P5TPjikbZTkik0kKtMjGURpvAvhSf/O/fQ7HX7jpOhYNM41jRsyX7
XnRKhAj53qLCwQQj4+4suvUDjVrNPNgjG3Ksg6dUqxGk9JI9qKzdyIN6LDAdJSBR
Kby4EFaerfkg7uvkj2c8VmHvKAd0r/wUODwdrr5C2zA6PQMox3TbcMXcL5AFNJwu
sM6cEmCRhreo27o9FEgm/GoWdqhZY3rzSirTOAIixCscoR5R2y89XU3MzKTh1dQ8
PO36CZ2xBsDOl9QODSN12SR3OfRRdWWNUDHCzS7tpUnT/J/3wBGy2y2caAfFtQIh
5wSlc/iaUIKtNsmM7uPL+WqwjZYmIUHgY2DR2Wwh19yoYuEbErDYdLRvbIUKb21c
1Z01aueh05r1j2xbEKEiSMZOknBUjj7cfnmKvo8v5mDwgx13TiHVMwKn7C0r+Md/
HOIbfIABvx328d67NyQ6xdr2Z4F2OZKXx3w8QPa+KQM0I4Pmwt1nanRLdZR9oi71
3HUgJvgM7EjZWD3S3B6F88/5KqppMbcrYKv0EhfRVICLsquR3rsHPGoGjFij1mkr
HMTU2zKMYYShRdBIHuM7wEGxe41BrlPwC/OiRMSaNzJW/Ki/C7JZqNc3NEA+hsB+
ChMuJ0adHxxVt00HYJ2xbIW7w1lgYTGtns64jFVSt1x4WSWOHkQCrzqy4xeVJtBp
x7cJ/gAaKF34AVGNKFLfw8DBhy2I0BS1JWJ+wzpuOgJRsylttOhaKzyCYZt2j8P0
7B8rlD6NqG1VII5Xu4jslLjQKRve4tRpa0zAMnryWzRwHRg3eIoT4oiu9uOJFXJV
tN6OVv5bVHS+wWyNP/fj+4rnfy3uq6MGFKzc89zHCfHbC1GjhN+hMgfVTHD2oXzq
BlDTvYF7VrCBb9Ol8eILX79gi1tBDk+PS+JAJ/enBh1PEtR/K62ZjBiwfhLBHFFf
FcvYT7gbCxraFvbYE6cZRDyveZ6LtCxbEJJWYJb2WAQz7E/0255dGkrKeP47uqCr
lA2D8e0cBkVNY9J2wqiSAe3sKO9G3nomYQu033OyJstWOj4k/D+LK9XB6AL3zuly
a4KJCL9rprEazYTwC/GTsw4++hgXng3kI4Xs6zOwFtGvL+5eTLyPOp8jGMWf75FE
2CZZp6zypinthKCHkeH+ifFHtsIwlvhO/KKaUSnMH/flNqq3YeLgTqAowsNi/Cp/
Miqh2EtftqtmsBFvlaOFBnfx+s9mlGXanoHI+gdM2haAbhc4O4FFut7OUKoCmInq
9iWD/YJ0dA3euKvs6EiCJnQ/7W4Y0dkA9knwwfR3+cn8XcyldeJ254WFOQ0pue2n
VffGgJ5fL8tX0Bxat3GdI1Opw/OyGwoAIDwR2ufwWxctS7N7dQxEp9fub90nhK/t
jX7/qLF3R6SWlouT8jL5L6Sv0m+PlvNXDYsrd7SNW8koa0gYX7vAQ3bS4SeMtaE7
WN9F8xIJ45Gju2swCAxMO1w7DnuK4k4wvbYFlbqSnj5uq2z+6Jvi2b89z4qnlwGR
m9F3joZN/LTv/CLs22VcRDAtk8vPTf7+5UhUdWD47nh1lBfNn43/boH4nJXPd5et
hKCMh8VZ1VsfDyGGbtPesK2/9lQxAyy69H1RrwMIivNeMJ0sdoxJeygzkT7ZuMVb
esD3/QNeeJOVUc2YHaOrU9Ygl1digU04GWoBZ2opr1HGWpf6hYSzZVcJiYjygHs7
28zlwNU88IUwbM4X74aVL1yyNJMpyk6lI9ybwaDLJBRbPGg/mZjHv4IKGQr/ntMX
rdQ33ubvvPxxb5WmSSY1y7AjR3G4HMnyQDJoMqs7rRm50I3zT5kjZoFhC242RDox
SDR0q4CU1gzb9Yoz+buY0jfq8TXt22LJ3AXDckmobZASciH6IAkkB9dY5ttF7d7X
DieTU3O2OvQ9NpKG/jFAK6oKV/Ce7iKdWPxHoh2kLDRo+z9Fd5QeazKuPdcrt9wF
OSPyhtnVByot6T2HT4z4siAcK4s14boE8VPJmcFXivgO3JeLNnRlYn4ge0RUM5um
V9LxQBNxRXpm5RvUNQU/ScSIdg8qoRUQsUd4OW8z9dYeCqVrMAeCDSa07j2mon41
KwqmiIoz9MAqgUpfK6Rwj2X5u+KgKCv1bcp/dcZwfBZlXE7g4sCWeWDXHjJJOnZC
VBj64GaIXqpYGlQIofYA5wMgbXIvcKR0zI54R2jfQgZMVT9lgJf0HeNXrvDkK8Wn
qU4Md1JtlQ78bGBFq0K5NexpZ2JCoR8Dfu328MAszNDOiFmP7+hUHDC76LuZWFmX
kpLKZoY+X1VpQdgzMEF1w9HfHPAcUSBRqQQMZZkSq7wXQkabY556wwTu6BD6wBhw
QVoJo1Dn/l3tEBAIMSEXfzGJNFy7GYENq+NCLEXOQxYGjtGiisg6azfV+blLp0/v
7mvvsRr7TiqN9RazDoUF6QJ5U6iExiCfiqZEewHSqu2FhrA1jqRh4GnUO91/iJ0D
hVtZ5ctqDLZ0GpbGQt+6eJPQEuLurfjA0TDv2UXa8P64/r0lytHOMpWNVjKJq5ml
3k3wYEVwfV36plZO8eC4WTAT2LQIk4Yg13mPPslj/Q5jl/eoCgY/ohHIDh5sNEI6
R/oXeHuWVpNEnklB5iIMzcLB0LfkLLT2clO/o1avSFV6MW6I4DgU2O6Qpi6vNbSv
soKgT2arZix55DV3sJaWrM1+kJoFvmkSdwSg/dYEXgQpJJsn/uE4dl3ZfyknUqkp
aEJ3jHQD6omMmY5DIM5QtDzv7HNPkX3cIfJmtnaGe55DpJbqC6zIzPec4vqZ0HgP
5zZIfsH9oBtmyDebRTTjafWaxGsqoyTRw2qVqcIAADxasSkLIrGCQm+bnQqhkRyP
OmIhKrcvFAG8dr3tFtvEowRwvJd3+otYTzsc319RlhIsRkMHFprCrvTVFDM1UJzK
omZvkvhfDGwPhZKTIlrqMspUkBUaEccHC4zM4Wo78K9GRb5Nd4B55O4f0aGVYdDd
5inNZRd/7GpWztIccCkQNdKIf+rulXfl+n9mKVq5PL5mewsfY2kprtOZZCuniYD4
1boRfuGWfHj9I5JeGDC4LSVrqlZzjKNrK7PMOUcRzXIZwRL8Qh5jKwbbcT/pZfRf
Kg1otLqMQVfhPlhYFdbXoLVdkLj7MynWS+at84mqmT78hCkBah8eDWxiY9Xwf6L1
c68fE8Kn5Qbb6nnj96F446IeCd9Cm9ydEXYu+s5hKhJiZPsxaBxu6PXHBN1JPElR
TCs+EYoLPKRPaGNoGoZdOyuhR+gHlKuASORL5G4R8kvvItUGepbVcYU/DO/1OOu8
3L+ZJ0OMoAlaopSOE0c+Y3pGWpDZR88b/THEhyFLIkMA3Wiwe3bC/XX/0s/fXLfq
j1UhvASkasG9m8mFUQp8eQyEx/Oy2U2T+ZmzuTFddzNWHJESs0Vl422XWJ3ARKEq
Rx8D0w1XkS9oGEL6kuSkQZp5EOCQsQqULZUaeJPq3oVZ8b3SCHSwfu108egQThGh
L89nJy5ET+GOJZiYx2hOcqFX/xHnMoEaEM7/rakPQnRxSlaqyQx2Rh7eosMauOzi
gcKjwsO1wd8oB3wuCrT/ibSWLycRdRMwevNbJ3p5PxcUqY/BveR3hhxW+K1uNA/P
WKK87GOlHJ3I6p0wnGgwH31LM852XGr7f7UK6NDTQ0KROtFkU6eGJy48HKhJtpde
xaIUj6LwqtPvzv/z2GJE3tdyMTeS6mik0giS9DjFP9HYVm1gcIcYwKKLYK/Yt8mX
5ezLI4x/84nBRdWxRG6Nyfm0BpeAlGsAfAsEj1TO3PkfYZxaLgjp7EktFVun4kp7
ettX9S2yu1RCiYQub4vY7Cizm5VPzJ3HYekdiUh2RRudonAkh2MdJ/fbqKDaL0pk
HJgeKAuECg1ek98q6p4zOmlXbgB+mGArtbKdZIDPZaw8QU7FP/8UwxKsGSfMEAZO
F+F/g5yb/96AxImvDttfMWBQMNq3xBScyvjBokZNyByWBibErW1VwU9xl+fh/8vH
z7PrF9D6qWCBqNis7Q8fvANBz/b23MByhqBCZ0Qt3NIGScoLK6J+gc5CylWcVmja
snTr0/4Ix20Oq0dbiigVXnWNoRYZp6Dad3RskOVAj3p97hUDRQ7+HPnWqK4WP4wZ
J+j2XlDFzTuW+qWOtkkzpF41fguGJn/IUKLwNxCE94KFea3oD4BFtOIcYLW2qW6O
bpzP4ea2WtYFh7y3mn+H0qJdOsOEI4LbMvVEYjIGRYYhbDVB7Yq/2MlhTkv1cbTB
RIroI6pqLVkwy0JhX0UnRIyLTVhXHJSeZ31i7PP1FUT0tLsiJJdGFwQxDMuo/v2U
wiDJcZJnFBLHGpCdMPVaNleKn1x/qNjMfKKMGTbtPoSN5X/c1fsVLzlRxV4hKviB
hxmRLtfPt6+FIgIiFGXzLJkuM9kOjyaCMsg+cGZjjeSRccZ303N+l6bRKIW43pzk
BEfw2WNVH2BxB3NxTU1vX7P94SOSf2OGxbaNcGi6wr9JXhDkphNRt8EGQWNhQNYQ
hRv9km1j1CIg8nVL3/srJdUzzvhSCm3lY0MkW0631damt9bBRRbN8cEL0Fsj/gUi
fHo+sUiB9ZBTDAWyszzeum3USgs5PAisGvJ+Be1E16Sykg67jpOIRqqqgbtJCxs0
l88UuELUoHM9HldiaJPxXPp9L+LU3JOVgmHzHOQdKUc/O3znF07GXc5IA8g5cfkA
+d8eIr2jZaFfhCXOyAxgAQr2ce267FPJ4JiZrpihEKWnV90U8Dx0+JRcaOVifE43
NUhz0tNg2PwD57q3bPbwSO270AhqbindKGjkjDL14IYqeDuG/ngJJt0vPDv/TvuB
ilrzp/zOp+bpvWVIAbzWLPHkkVq2kuFRkbxn3oZchEhFMbxlZ9JOLjyfs12Nt0lt
keVpxf+SApCAlZ27CzcuTmbUJMLC5aq9N49N3I3YsGssgwcGIN/HaC0Sjy4zD07f
imlVeCJ0nMtINQ0rkT5DDXoVs2sHgex8nCOCSF7WYdlYFIUN7B1rNQtYjU8C6r9I
88fSBumGsjjZ/UM+YXyq/0vO2vHn2lOxsv8o1q0pKsQwBx29cM433oPlyaEngKgz
jQNSzznF7IaZ8kxI5ADiJobZplKckdcPc/PM5UrUaJTyUpdX5xqKz7EsugEi6BkO
FkzRurndN38A9aeCkmib47F1eHPChH9DxcCAl92jbhGdWv1msXau3TuMjr6XuG8I
f15sQWDAQakzE/D2mdT9OQfINtajxGXmd/5MXGqVqXa2HJGbnqLai2Lu7BN8s6hE
wYyZHGZ+tkbcqtmBjuR89Jd50wYjVDB9D6hNFOJGBSx8H0/DTYVsl+1hu+5fJPEe
/BKDqAr4H9EqH0g1J/EMXO0t8w/LgLuWdzweAmXHJNMcLZugueSXXNNNG496Ybwx
rggogLEQmAmCSKpVbGLPZ7L0ZPFA5cavc/z6okCE4JQvaylHdh39Zz6Na2neZ5z4
GGcwVsnR80CIQboer9CKKqBJdYoiWrLQo2RNcefbUyZxPcRa+rsfFz1OjZo547ey
T4JmM0Q263+HuXnpHW7rhyL+F2EkPW6pRvoPrs/oIO7T4uuVsd02XQrJEUy9fNUQ
ZDfH9U1PkHfxHLEK1C7QpUBzNT3TsyEM2089P6OeXwRiH4t4h/63GfNYuB/Wt645
ARSQKMQ6h474MpCKRRkJF9vKqhXLv0jwFzV5sA60YKcQ65kdeDWb714eb+PBOOM7
OWk3rzP9juNPhw1efsNH11mJhWMU+ei911n/8gSpsQuiA/bfd6x1evPjDAsnsqMc
YhfkmmL7B2Jy1mUklbAC45OMwSrqSQ+FNHEdPv6iiK9ZgQTxS73KDxnFcz6bqhcQ
y4SN0lg7BWAMxJgoXDVP+XwLFdQ+0kUVH360GdPFiRxgsbitKDk0sGo89nUucHNd
YV+aROwhlkA/kxVW+Ozk9Xp1gnYbTgG4y3aqU5NV/fVeP9QIEJ730R3YNLUer/ZW
Cp41iL2JeqEk25gF3lx35XARON1SWmA5DCxpB+puNUDiXPiAD+FH4xGwU9mKTjk9
Q8B9q7EzNI/kJeJoUXRVVED2TQNx5Mbx4CrRqvzwYV7B6+GoLxUMo3pJ/mQBszwq
AwZpAy82NfVJrw3KY0bjcBDEmWF8iXZ5j0c7YKh5FFMrFxWmv2np7r4ZGSeV6uSs
dPaF3QpdwsYiDIkGQoviTNesdh/COLiP2iDxW8sUzceMk/mCXmdVL3FmGiT+00xC
bkeQ1LD6IJa5X1G/NwwlJzamIWKtEc2jeLjRYin5d7yIha349+xZ23Ojy1XnCGSk
QJ1j9TkvGJ5sHiPU4I0m8eXC8EXuBMWF7H8XhmFzqsaFv3AZkB8lVnMsL82tt0zs
wYCHCEIcN7YRJHVXpF9KpzBXHkU2kbuwhiAbNCq3JyVOcvt/Hs7vd5y7edPvqkRu
yEg29frg+7GjgGdyw7izvXnyi1ShwN1dOvxFb3xSc72K8bZINP5ud/Vywd2Iieav
iMQkJaubBMy429zt8xJuj+2cEQWk4lPXifIsFDYNAUL6gIKScFj+qmsnC0Upulx4
YX5zgPlxHgp+Xnx2emDUyieuMT5qCkPL2kD+Zkk7tg4L/nQx/TAOAgykrA1ABekQ
fSDzAKv4vqCbKQdTAwiaeMp0oaO6J1PM8ZYW9y5ypydpIWMa8+0WP+zBXksRn7m3
IAjREXiJaTfNXc6pmWQqV10XO+qqxM2YHVYMsJ2KggAgTQA0b2ftZjdnU3RmzXQG
HJkW7QDiCkqcntF7g1xRbSs+Z4xC0NwfwNTDMruJErsdBu9Qhu8X77Y9VNiiIsDk
EBnBQHsYVa8GC1aM3XIK+bizEHuuFFCXAZAiWv20wb6jp/x7JtFe11dWJdBd8ZqB
cjqrb1K35KWJOwUkeRH6ewpl/m6DxKkaGYQcCNkVPMHHlCRxu/KtO6/LjEePhr0O
yZVMXrBuiQwWId9W3V+kPHB1ECrJShWJpPO0ZXKiWQaow987p2/Sh0FvuhGDgUpH
RXO+6o8ORK+s5044OomkG9PniJpWnK32dJUZ/A6dZ+xdOS0y87itT33vyNylUe2Z
rzF72HoRpDPg/2OmDC6L9iXdM5Y9iVvZQzLgcqlY4pceVQcRgAmqcM40AUOAsMRA
Fje+WjZDPOcHhEMvzJntt3srvj8N8RWTA9ETd1EnFMiLFi1Ksfv/Lr3bVkA/Hn55
+J0cszjVxbGsJptop8OiYnOO2jK5/qh5AJeTO89+K96tHk9mjbsNo68b91OKJofE
8J/MF7rz9J2NvUIF46aNAnu+M5xv7MGBE0lvu2RFFxoCDvGCUIoPK7asKKzt1qJS
qHy/7uGFaTkHut7AunKn2AMkhBz4zR5YXe+9Blk+yj2i+b4sSFBtz1m/k1RHfg/U
AWU2rGG3XfHccn3qHEZB0RHbsenvfr0uw5J8XpzexFdRkYsgg+B8fOTU+orYxiZj
Q4Hq/+okMj0oSQxDujkPiMcrb9Bf64qMCmYkE5BjqgExxlIlAk6xdWCWohIyTMH4
zfz+07aTkn74FTasHSo1nHCHm/wFPD2KIeM5T90ozKjctvknBZsZnSCAOyeCXNgC
AMlomeuWPLN30S88NDwpOy7DeRQMQfsWKSajFOpByIj644xvqoQ1gNqNBdrpi4NW
Euv8xn4cLsVaRkLe6x2Z48HV6wmSV5PZaWB8JdkwjW5+XSk38cLPlAUMT2ffdDpV
aGuq1e2eH8FqrALiugqDY1GZuUkS8ExuVKRUAyvYahdmlFblGr4dsQaxoNWAxdYE
VTBsvMDL3OjrV/JXBRY5RBMynjj8k6P5BGSKaXbTNH1h1kIYNLS9MmZH0ZLLfg1R
Qt4+dr6MW2Ro0lQxHpkUoMfSSUgIUQbg4qAwf8ZzU2cxyNhK0KKh0G3HA6vlOgeo
lTNS2bIFoarGw7KJe7tRU9PokDVtQyVzID16j4jVDnSwqS/SMDuFqYFuju5FZh0U
Mfk0FacJlhv0KugCzjVZ1IdYo7oVLnTkDqMluLoi6AWwX1HA0qtGT0ga8SNYmNRI
QcKkGPeqBU9LnbdjKsnaHBfJsb0YmNqoKGuGreKuTGoXSeFrIwbFRB3s+kkNX/Q+
0u4bYK6MSRZEyrRdqAQnFf7oiwc0iem95t4NOXgeKyFVmt0IO3L4gXgk1E6nnUw3
4ud3YFoNSAXeAtbu7O4i3yEDF1onnbhweM/sHC7ZgN7O1JDJlqgk8Gr8jNJ4NWKf
ADcarO1RXKMyJ2AQempypEUE7Lf2JvPufkHegsL0/XAzcRKnd10Gy+j0xQxA5HSI
Ax83S0LSoqYNO9cZMnLhfqy8RztMhSyJs7Itpx5hjcv8NIg1/klCc83GvxDN1ZCh
2y4/3CrdKuzkAcpp9E0+PfVZH4dW1WVsJF0wOql8Udns2URYc3Jsx6fu+/sYUxi7
3P/fmOElv6aiDRjXR2oo1w9WfsVTpgppvsexEwTDF5XJ/sZ0KqB2iXOCfMI+3pn/
ozSY7LFvYc14h9YSlk8s+2RlUy4N5GzQ2kVqyBaxVf/fC5nLXpDLHsStDPmB6B39
WQ65t7uz7T9LrjXLmdvwUhjC0lcVjhY3lYvdbNFZsH+dzC9rgE08vWM/jhX+/fcU
mCqRJhKdNUihfkCg1mDTkHhFOy8mm0N0wRw1klnEjH9nf1+5y/vB4TgCIfb8dfAh
fd7KLrS821Sa9jH8CIeQy9N/ch831wx4424roPys7t8xksPn35bfXenRrOe+24kb
CuNJOd70KpHQ/z/o7qmaOCU3SazKyUQ+GEWkucQ0qyx5yxK0RBFwxUzWcth82Wqw
+XBmpqHPFvQzB2AhrbwvTp25w0XpXN/WkL0nRn2hWfvPK3JYfFXUvhWZDkeUXnLo
IuURCIaGltecGTZ9tnYb7Hbo9vNAIlioDZZb31l5iMp5Dlkpit5ISV0XgPJixACP
ATJsn6LLk5rAXqPQX5eXLyALnF/VCGW0+zbBLL6dFHlr+bJwI7LIeTasrKgZVGUx
jQBUBZGkjqigaK5kgKziLS6DPyY+RKR5kr1OmE/wx052p6ucFNBRNmJBx6PcffXr
SLd1TrrekTAXuAqyMFR+PZYR2F8SF9bJrBamPL1Crw7Qg65YgJ5sW/PT/Qhs9UeU
L5GxYVXFsRkCWMqjD2P5sXH9+WYfINL5xJ6/2Ui1W60NKjknTiBeZHUlwr0ngQR2
4aDwhaoqQj7IbUHJKq7ptYxu3KdhWqIh406bzu9TPsJMqXDWN7k5bFWDa2MK066+
75Wknyn/HpqnVtymknZoQh1mPIQMrKbF6vG8Z03alpEnsbOH49UFnPNjyQmdUrjr
PcGpW2+j4Y3f1ZcDEnOXBXAi5Y+l7+mqNAXX4QcBFMA1SnfdDAA/TN0BYANmyfYg
OmRvGVGjfNdXZ9U7AqAT4E3TSM9xQ7Es0m4UZnT9dx6SeGEox7Wb7n5kft8EapCc
snCDl8kwf2fgSIJCB19vuO3EiDb+DyhJAhUsCawzJ24XbFcOL+vP7BlYYQ6FAjwY
X89jy6F6aHoYi1y4ItMY1fwC80A53jSeShFUZfeLHLqkTVhDKGMo14KFvFw5oc63
38xYPYpsC5BzHAmzv+SzIGDFFcKn/GSjpxTUAmhRP57ffxLETP2Sj2GFxY/hhhsU
vvq7N+aw92LSpKEOhTZS0Nh7Cr+EA1ZZunTSmQ0ZgfuYO4fsm1lMAsC2ttR3mJyY
GHfBu8r2adlQMYBONCIwv0Scxr+inAQNqFuJblQtLNa9vZP7kU7DNIpFMQw9do0l
kzHFYGvAdTeaFP4L5NGd4dTR8qulYGSVFJOflAtLYuzePdbHAC+od9QK+q8fYlq4
wmBW+F5YJnipX9rmAfqGA/sbWGD6P+4GFzfz7Q+L4+QfljYH9drI+zsOmLQSl81F
PzvKWRV8kJ8JxesNukmEM/P9Y9bKtsvsqL0BISr9K8UiuME1dnt0jASXpJwI8t9X
ovWOICQVx2cqWvhxhs7Km9/zZlVM/Kob5JQEVcz0mY5KHm7/vizpAEvq/20Ljurc
22iuuQ3xxh7rRFkQXPsGhTjpq5iUeltNRUSai6Ew4mgMGRMy3nFV0zaqhqbLSvIl
DcS861u0IzK2t99IIYxFE5bhskL+EKtSihpSW77Skhfsu0l2pI2rEKMv+zClR3uM
FzREschb0g8LG9n8fcZKiiPfC/bEZsUKxPaPNJs24iCr6CaHiytKuydncIN7T9F6
GgyoPvljFg4tiHRU9AIO0dUHO38cdYbtLBwMdSFJRRkP8dxuZixTReTjS1zWf6UV
x388jXIpRc74QKg8lYygLrZF1jyZWbJfuUecIO4Q+31B9HtmrBCWgJhyPFJGpl6N
31qZy0Qe4/LwM0Dw5sjwv9/uYZqseO79Bu8TA0b90Ulxp5sYkGdfzyI1Ef7aFvjl
Lf/rDtV0AMqA9TWvvRLQBnDiMrME/BZulMogI8DLG3ufCj8wG4PjtyikoNGtMqfq
RCCdRnqMagmKtmFRCaQ0dRKtr3HQFoxDCnKhDdLyIby6jgQp6Or1pBkR71ybj/16
DgNU/F5V0PhHhmh72oqiD6ZCoTyy8Bt88QSV8d+EkHJRA7jZ/ODKP43hX6kaqiGm
OBzgpQrRGRfdi9FClzK6TOSOe3zIu6BblX8SxbrvRTKCTsDhATEzTe9uTso0xFJm
1gV0pe6tlm/PMvLKoBEHimcovhU8AdPkQgkcF/qZcrQa+lrGftgtEf1t3sAeKDqm
j4I5/UeT/56VZkNwJgzjVWVZ8EktLdWthI9eqLCEFm5gD1KyrLEWvkfBtLHnhc5E
Col17JJFC+wdfuHktWtiI1FiZ0PiCnJbT4RVkdr+G4yEAbRB0O5l94cyba/+GWih
whVivdTNvwqvUZho7H0ovMWutRXeCnApLcrWyKe8b2Gtz1on/J4m5m6O5XrxDkbU
hP1BUleIz5P8sDBrKlC9kOEsGs4FUFUkbab/XEtlrPd4T0MCzcuh/P67xMupzdtx
iKtj2wd4PMkpjVZBqppBQj7iIx3pfea9UWFCnBMtYp99U8JayUMzFnuDKBhC8g1I
vChe4sUSnWCuhuRHy/eKw0jDsKMLrV50BLZpddPQSYsiqZjeZbIqMLE/NfwZRmOv
kVKRTUq+pBxFPt+xv7Poh04uo5HnE5UzEzH9m1lsdXcxURY0OZAoR+DOHxnvOXbs
gJgQKoifmNEQ3j9wHM0/73zsi8fKvbRpc1ajBsU4z9boB4jXFjLzfLY3u34ljLb6
//Su8IVpaSEMq9VoxnWV5rhDrxgSOS3gluplTA3UDGgf/KgCtD18WqKTuoAy1fcc
YauOF7RdPEXxP4FFxz6laFOd4sK/kByYF54bT89YhXlBS7GIdF1y3j+l6OV8y1FA
LygHFoAlW/S/gEnXgbLYiGesAZ4YWW29FvlW7axg3b4aTpI+wHNSEdBsjJc9Ua7d
txlWEdpGKY1LbQxj7cbpzcNh0PhxZr4rHzqrgI+vqCTCSKZvBSlHYylCxAjRmRp3
3tNqkHm3z7+BuHBPIp1kI2HaOcPvfkF8ZTFDld1t9eNuslYy7kVtyBpMib7PpAPr
g/129OphgrFL2G33rAuCNRvdt/gK0WP5CRGpXp0Y+DIO+HD2a+s8RNLO6NI7b0Rc
6geT9l+QElBk+WexbXNSJ+SRBKVuWHJQ5I26OHh0zvtG4G67vP76whffQK9/nwUz
bZ2OKHoX96QO+AENwnmcxKSGJwKRsJkLShLjEg31A5qduKpL+zfFqvjbo0dWsXkn
19WZPY2EI4Kb1k4eyYmdYteltgVm8yFAwFfgHmuWpAEt4zqbBeUg/0Q3tPVOPZ8o
60QZwJNwOtPkHVLvTXDRKsorealvZcygEvLb0nZtRANNYVZdHymA/Ll6Hw1I9MQu
/5iucYcyVi9ssRed1GUoEq86qSw1ZWBEy9nB03Tcw9AtkFKWSk5bFtlNXe8oR+KQ
Y9VZspsp+Y6UMb16AB3PePdqiCZznAsG9QDKuUZOQZincXRyny3jIoYR3FxlfTjm
b2D00l/nJ/rgqR68CH9VV0LROR3/M5mTfloCydQgbd8UNVQ6kAwjqFHw+z6pcm1N
suhdRjIlQDrHJOyLoizDlbk2RbdEoNmhsUrv/dgWI3P34noYET7yEaTUSFeQG4Hr
uRDIjj0Zc+K75PpCQast45kn9Qu0XZPp9ntfwZA4Sv6HvuHAp53Q6Pspf4ytJDyi
bNisv+zTmratkyrNv6g2oUUXR+7RIC3Vaqoe10rIKYRoAqi1e87gQ/Dhglv66bUM
rWKhTzwJgZB4NVfUd1IzWjoCvDhQTXAtHrRmD+j3r+a7Om2qMOZpGUhIjP8RPz2A
mcj9KnGiVWZcd+PWE90LaVHPusqvjT+HBewxiG3ATn10oPhYUhEygiI94Ume3Mkl
/k6jLYqbCC40dJRGBUZZU+6QM9JxBRQeLckKNQHxDQ5+Av2PnDr7TSt4+kI/bB0b
6nUaNnnxg4A666zOyvT0hHJUfY1xIizjE6ksdOjJuKZD2BUnXS1sEdwMJqn7vDwH
Ob05nb97/WOEvhxdjqDvxyAYqy3ZzxZa5GzRDRL+OUBgOSG1JXx460n/49bw5nuX
nUrLJMJGOEx4nnvY8GSc8kbzF3R3kFBrYV47YhTazsvPnQtcvq6h+lMkv+PHf2cV
RWQ2WHdwrH2bkpGYBqJmaua2MZpe4rjFDdF9Oie81PBVSGLe5BKTYouXVHOaJ+cO
rZ3fN3uqyR0AyPoi9G42ic0h2KZBXV3XXwc3fwNOikxhnfzmBuvECuIHLn7k1OW2
F5qRiqtybF4qO7AmHRFQLgC6IEP3Jl7XScd4hV/ABl5/9R9yP+SMTwWQdNs1Gf3D
RSSzcO28pHm1GSW6vl4dqT7r6iLcC1mTLADbkaukeOOdnOLegDiks/phxQ8qc/L0
3SdcKU8OCVx/E4G9zMlQpYb5x1QmZMd6m2bnDc3my2QKvOdFVqBiOxIJov0PxmD/
ft3EGBVhMU+KISXADY34gr9YSqn57iDUxWRdmy4Xe3QTJjmzP35nXTchizTww1tm
BjRI77XBMOKhCGIncfdcgFCReac58+vx/scKTddNzT1e8QN67Yc84xWvvnFf1yxj
xdAi+Dmt3L+1DBaUm0wjbgnxCcHqAkhWdAbVnXfLwCStV+GWbf7y40Oj1LVT6hW/
MFOw4XcWuimn4dhgLAH4MVaI0YqvJIdcRNRhsM+QKgo85L6B/cHSI78Pzqd7LnW4
Oc8qe580zE4unkjlFqlY0b0U8Z16byToGvV0xMF9XrIX19ceYJTGmiVqngZZpW0P
EuRiaF1Mk0b+28g+0iBhfch/npTC6L9BU1wqOo9KH/Mb5oG9ofb8yA2DZJ4iaoQr
jCTJt31xZIhZ1pqIKl6pQf7I88slUNInwVtPek1kY8XxBX7BMlXHU/u2u2PoCcNq
RbM8H0J+AwQW0kQAn9kWHkDhqt4ab+nqikGVafBexgWCPVpco94b4Jw1MdCtY0To
ACbKGk7qZgW47LFYBq3tQ9GPRqcQ6CSneCXIih6s/kdVqYTEXmAxlYphW/aQM8HU
WBOosuA8NYcxMi5awVySFJxtXgulDxREyuaDCygTRPwxj1V9uSRvkGNNCx3jXEL9
YCtMEnd7ybrt2cjPGVVil9LEVS4tTy5E6aqHkNMS7TP1Pls7813tb8hMdirFlOuk
kHCf1RuOtppNFOiKJH3KyIHK18T6AmxQtGl2exZ82xf3N0gKymsyqa3HpUK/AGv3
N30vOkxtOq65gYmB4IeBFK/icxDjvuJG3gwyqAEp7OyfbrUOp9u43+zZTX/NZNHV
2meykWhMR+urs/jowqC7HvObAR5fqT197FZ6Mcftb9fbVf81AlEtBrvvD9iti8Mc
+jo4DV+4IxvG8fu7vALxq2F6hsW5Yd7l3tjfmJWZZjO3sn3koV4yDbn1uSZtld7I
x7YG2ZiW1cYc7C2oRdXqy/2Q5eEp2m4nM7K9GIQD8U0sm4ik4VV6xihLd1ztUx0X
K04GsynmdBfEOaEY+SgrBWGEFpW0o80TsPHPu4ikOTnY+uE/yz4K+dVpTovm9a47
ofTcuamLEVHVkm0/ALl7rmMYZno8N8lOBG3f4nMyYJOHhVvPTJ0siMIHePgHIrEs
9ncaAqVxik3rN1OsZKuZc6d5nqUKLckd6lx++s5Swc4FyDFRep8LXGpqHQsnsHkm
ZHHLwxjhTEFlNfr+LRDwa5IMtSGfqpMoaO7+5uFBvW8k9S7eTID0d/ulKVNe8Ngv
LduRPKGEhzvvbohEChDxuEXpJfzQhPRbxI7449A2hRpI+ti3HFxYVFs5Dgp5FjOL
arAPeT8ED2uJhtM+OcFJBjVDxDll0YJcgvo/ezv0WggFmyFoG4LFn1L8IbC5uWC0
2NGC9p35c1sB/qqedm5T75jkG5uasFRNYOgabMdI3+vz+wNJSAyw6W1IvpY6bgkJ
W/b/lJBTur5ymrxl61eY/ze9qskk0pk6AfkqNqRBQkpS5Mv7/pqdkLmnjh8m2laG
p03VBv4LVvAv1pPRPdnKIEi1EPho4lbbeoLKohMClEw2tXil2lehJ9MmlccbFLlM
e/rUvQ8sMXrKv1ZGgISFJpY9obnOiMkB8QLOCd2bzVndoTqePUPI7oW45073AHGW
z2JC2fSPA3/1pgoQ5dLTzuU3PDZuz1b3pdrSiRrn7El/TmwhFYAyEs+BISdPt17C
RGTFkPy81tAUK3RUJA3s22mIgc5gOF8f5qKxqydeP21tfha1Xwqj5NOhcqhW6yrT
zvohW9IkVo+yUcew2B49t85+BsNQggyb0WKDwckTu3IRqkN1GVJWHVR6GELGeO4g
yqc8GBDzrQ+mczidCciMwQRcfbxkzw9GMn1lUt38Iq7qtgbTRYMppknJpXm7Y6zc
Ud6fhbhwvEXSntwroq5p0QNGKkS5C/KUQf0mIpfajlOkOwGLYjcuT3M9svx6ZMZu
nyCVn0Vlmz3xc6fR5OkXuIlX0EaSWdBpRzF/eOkf/ZJmBnblxYUDkAVuKpv6rIKX
WZn+zgMfEVI6+HxAEfFUTKFS81QUltzEVpbu15XSrQh/bjm0Z9HNRqpp1cxLAoSC
zMutlhdW3rU/oLQWlHfBYvCwspD2IrTTz3lQk031FcBKclZO+CHqdurRj8Wi4y0Y
OLxnH/S9sn0I55SBz4SCUqgQKs/W+gzj7wDnm4/ElIlyfk0/eahMozg6Ah1AYNqn
TbSAF3vGKcGbyGiS37mZeznM9PUSuAL5oe6GseyGVVrTOQDchQy9qmJg/7iEQsi/
bqSwn+ore3/XiKYrk5HXIzT4t69bu5o0lJ0jhitwC6VyoQMbVAvEeG7aSHB5CoJS
UUf5J9bTJRaTGJfV1rKPJlUS21DA7H8T07YNLLl/d+VecHlbvF4LbYRLaCONi/EZ
3D5pb0MJXIOcPoiDYC80wtv0RrhpE5b4ZiKV+2N6FxxM1Y7qDyNoMDWhoTL0l26b
+V7/Xcq/QGk6i0KvFYf2f0KUDKYJnCisRu1UVCZrfKUvjC5eHlcPcFzvEq+Ep6o4
u/qCT5BQES3yPbTJ3axSnIz0UkXLIHHfYLd284L5wBLxYQjAv5DM+bP1zC/PqGHe
EPsIGbnv/3wrr3H4sH+DlKS49yxk7UAJZ4xzsln0yunoQWO0YcVzz2I7A+cUWcBV
cRdXB4NF6mABQQVkrHuyIj62JQLg7FGp5ciy+Nhsz9l+7WQsP572S0WFZSJrf0Cm
VYkZS2yP2D+K/2h9bybTeif6rNqnvJgxOfQBWHbmyOhZBtsHW1UhlmMHf9vRee3y
M9nLFcfZGP7GelsCsJXL+mBrGXlUlnrLlfCOzYVHCr4hFHoaaSSmgocFegqRei2g
dNR57EXpUmtVenncyv0LpOB/AMhICEehuSLXYKhAt/CU8fayW4V8lUwfhv07Ii5a
2OFo35XoBKt5DQDH/bVV2nxGV/LLBejnG8ap52hWq0/NpnY858R/gXJoyUOOiUqm
QLImIR/HVuA/eztPU/MistlCvYW3x1CnkDT4ue0H5DKmVbIWLsQOm5FfJ0DeHm3I
AtKr9N+Ga61aPaUKWzwEF9DuzXNC7dYqiu47hPDiX+xjsgONbaUpd9Q+uPc1Nk+P
wC6sgeNYXpDpSNdgoeyT6FpykEcc4Fzp8gZSx27lwkY/K+wU0GcApaiN8uKn0ZDj
Le+3twRftozTy+OxSjrdBJ3wEoTqiNu1rv4TrtX6tIMGIpsGQgUUz2vWF3lQUQ8K
EbWUJmLZ5PsAeN9V1oVW8nSVqMdfN0TviJaf8qtSl03JODX0OSYgiSpe9IcBXbPB
90KnpWb/2jpEfUj0Z2OD1RA1cbngtwo2AErzj9V9/XJPKWC8dU+lYkGeDCIUcU/S
EDFyOCyCxylNtHTpweZJv+euFjhoEkrcZG4BZPHix2q+k9vjF36h5ydjdgROddXB
KFgX6p3zIt5SpdR4c+gTgqNtBw8YtJWrZMSTvaXe4+hR5A9x+pRq1+hhCasCXS9i
4Jqo/buF2wUPY/kES1xjZhGXr1cFKswVtMbP/VX11F5Fn1KVcEuLohwSAPCHBKTz
J7YBBVoNfDYXHfc/vdwemiUlItJT9b5g8Act/MwhLAlr9GBZqWylVUeYtRPxHvPv
WbFEjqhtsBke663/TgNWGlbiDS5BCk/y6fowazrRvbApP7B9+vI9WPbuTPl3NlmX
pglr9l+m7XM7UcFFM2aBnYdq+uurCFUZDTUWq0rdik1+jr/zd6MYAPOqv62t9qli
nJVcCs/mDslBGC2rUu0oaPiVZeXOFE/RHiv1NEV7CtLNr2q1cOGFBC4WkIsm8GvA
5gva7lTDCAAQHS0nHH6YKYW6whvDA3MeuP+aTMPYkp6+xi6e2EWYhUqZ7DxC9Lw4
7n1T6pkja/q9a9eMlt1ReTfhHd3i+i61D0OEUPZBI+29Z6s/zagx99OnvMgCHL+b
vBgFzP5zX7uepP6fFFWQMcAvQrDPfMlras5i+3OtV/HhwGebK+f5K+z0dsvytNJ8
MmDTS+lRjeLaaQQLR9XExhtCLxSaiiPYj/mK8jLMLQYR0tttdfgmWO5bzzf3h8SQ
GzVrLYKQPsiHVEFktV7Bd+Gu34iY+y/8Ov7iJK7Z3GZKo1UrjD/emAAAgGjQlSZt
m6m/26hkxKsgyfcRIEjevjR+vC9k/DfwOcMnq38r7O//nJN/12Ex5/x1IZTxqsHi
rYFGi2aeer2A0oGkEk3QSPaMO8kqtC5VQRDIIxBTcTGQAP6rb9SDxC4YrJ6UebM8
NFAlp6NY4HTVk+uu6vKBN7crjkMxKWpKyzT2jbwm68pllo8XKyO4AhjBTDyL5T0s
42iX/r/o68mb7sR50QeGA1AG17XYjLjDDeDVv4v9oO5FSRB8cZZhgltLHbG+oB8k
Ef/YUMdZt68ETBXWfxcCblsOHGPph1nGUafwDT3nORZAxR4HVhCgzZsgUiApi9xV
e7OegLPIogSFQkDrmRlf59vUtuUgQ4dCgZZoRW2WMeXHZ4ODWPuODSPgH28G9F8j
U1dEVeLZatRupduJCRuOisu9tkQpapIUahl67v/VBJSyganBatZp3jG0C+rb28Ov
1ynrTZg24NyNfGkABs2yF6FYGuovtw27w/NhNXfyTrKb6gY22RdLewTOPyFCOw0R
8d0B9HmpHDThlqdqxSEsILMXkK9VmJOWhVc4wcJvFX2m8X9TyNRm76Y9LwGHp6EA
o+/eXxiN0USO0l2s08RdC5hNkzlCauEVECRZ3Ke4ESZG7Vd1do5hWDA/TBe7O8O0
LlQnbS0BUIYp6VG+t2lehrmsgIm3ROmWoqCtOKNUaR0MzKJzRFTMFspMoa0AGpfb
snOHljELqUziUYuQ8IQD/Lb6ikfa/wRexJ+UA+Exp/J4b/VBtuYzpZ5WIg6ScF2U
W5/o5wpy39WXOL7QqwRyOKNkMXicFsPszwvHt+bBo0+NrCNrAzc89CQDgvl4epct
1bvNu68jiM/Bd5KY4Jd8SulLygZKBQqE/n7TaPJhA99jqIgYu4U4CbObqKAmUY0G
1uqm8ykp+fR6EEacgeA/pktWCntDNoMR9Y9kCIK8m3xLAXIt/CFqRgt7Dle2LEdh
Us/35U9YK7QZx6VwB5qtw4bQZqZqLc9XrA/bfaLkEZX1U/23nbFnC5o2nRTWBNno
Ey8TY9YDY1RrmDJ6RTT6X0xmJUDRSYy8DeCaRdZQd54qx2dc33jierMh2vMqgK14
/MMRebCZ/ysrjwAcCYLtsaE3OGJJzVWXOU9J63jzqciILdWsVt6lzdqHMFlOW2qH
f+Vv3XxXC/+5qjqRFe1y2WPOHIEDvOAkYcCgd9GEAGVRirKlU6+HUZOA5/tPX310
H7woB+RMSR9ASQ9dILpn0cV8WziE0hyQMiL9IBsqTI+10Jux5Pju4Wev6bWrYaoN
NfYNK8vpcRYZqwon0c0s2/KaH6KZycx6q2HNMlZma+gpwhm15jaXNFPmtLq/FWm8
D19ZEPbFXq9oYxNZzVXqRVR6UG1ncV9JCZ67nbMbcOBhFA/BXd53epsKy+f3x6h9
EML6/Hj68jlyKaKS1Siev55dMX5KX0zWBcK/6s42D78neENy8j05lvoOCuRZF5n5
CmwzvdptiFCEiSj4R24eOeFNihd3K8Ei2UeJ0VYjVQHCiXQreaf2HAN2A5fkk+LN
5VMKGEMBaHQC4zTIKKCWqg/Db+5MEIjfZ1/gTcbdjtKp/3uqpHFKhs5YIvKE6koH
KdXeoMjXccCRT+Tu4WQJldFKCB7S5xb58hv8KoKgH7ftLT5AduOfIv4UGzZj+lKG
nCMOzca2C7DkxBf3eGWbYAcz/zjtcm7RMIyNpgILMTuWGLW75yZCBFfTed1EQ1ld
Ub06QPr/2dv08Ot90/h/Ry6ZW20ry+U1ZoOQvg3A32I5Er3NKqKrdbizTdVYTJOe
teZGxIttDWWczjPZE+eneK6GHHz7UM7uTIVjVzLgpVkYJ1srn+dt7zd+vU5W+GaB
BugNaaG+VOu4kfGexLc4lu1aL0vaSi85LSGkZy6vy+XySjiO8a5BOHcdDOvvyWlV
9FByXuXjyhyqVA6jmvkGaksAhdZIyAcsGNQhUPJmb14zUj14io/ZuCbjdnbXic9+
QqB+J53dNMBGS6qlTQoIgVT3c7IHtFCPZTWJ8pRveYEuguTeIcE5OYuK9AAcKOuE
QNKG+7mm326U/a7ULwsYgdl16B2M8j/9jPHjfYoSdZgrhpHTmwxmkkKgZUtag56M
5fDmL9fwed1KswAGhkbDTUhkc1pGwEOt/KQY54gLoX5oWVtSVvAu8RN4nVhLnuIy
za7xhYSEYjT4uBLXF0ouQDgwzkF16Y206NDe+N2+0iumjWUGgfaHJnfRVbcjY+OH
5NNVQqFl8+pVCDJ4IvRRuQDSaMtoHGANkTWmnCfm6RDIS7xp8rsf6XxPeQiDU9fa
6gS1b2fPpTt8rWXoFY6fRPcQxl+vT9Ix2HeqD6GIyYPh8awwQ0aXlm1+hn66EERx
JXb+jYOe4WW9ONBTDjyJTBddpVPrynYq1ikvTfYmjDY/ny4jqY6UAPHmWWP1opka
51Oj4jBSxFT0AnBHOdK4VwlxuJXFOdNtMJnau1wTMRPRARrHB2ydtPggdqEo49Qp
264dTzw1t02jzgV+UurJbw25HomnnMkHYNggOiFM7BMH7P3s4/N+GHMRpEdb3cKp
ZlA50umxl8BaOvCueIYMUqvdWnvWrF7d/fZXhPrQTWSapnS8thyKNWYhEU6ONNM7
G3zzdDkmwx1xCcwNoF7URS5ksCEDCjPhfqVXTrzBlBv+sfUy9XCIEtjGCTBs+gzR
YT6YXT3+UXUvaUVaNaJlLfA0N31rKIxXdTeK/WIzbrh6qYfbjOLSEiilBtxipQAi
8lu0kzi5NTawMUUpkGwZMYzudgLsd6J7aNQQya9ZOW5azhF4fNB6r1WmHz/oNAME
qyac13L2OV2vJ/dKNzd1QjW6WIIdLV6kbuGe7JSqba4JbWeAtaSTjCgFHpOMYPog
KgniWWnKYURUlbEQRnZKJ9CLy9H/jdbUySPsiSV730Kfg4iSED5vkAYnDY12Vs2u
Gpv41ktyD+Oz/KLU5pgiU4VQxEEqEo6djCWws8VqSv2SHbCImr7GyBD6KmWa5fFJ
2SrrkcSJ5s2OvyyYcNqSQXh7jUuFBbk5SWxBoxmHBJpetooTkga6As0AxwIsg06h
C6PBUwjPxj6RlLIiReuZvymYkrLC1zIGXIKSrsHb5nSGllbejWtD78Ff9xtDMN6N
4b5wgowNuSWxhQ0U747kEHgSfmDcuHxr+1s1hjiHOud/g+TMZfOKaG2hBcoB13HL
d9m306Ho0quuD/b8xgWat0dvLWAZjA3sTYyCTH/l+Bn6pPmwQCbXPbCyb64/4pcq
x3eJuq5pBZstan21r1Gs8gydGWuIXZQxoxsTVum0Ij7GEsXaEQxW/FX/Bq2Zqqex
tPwAPZDnauzaPw4/GYci7VRRC7LRY69jvAkpFYPBw2fRBBeDYtZfackrVGfuxBRA
yw5O1Wo1zx+b1mabB6XAE7WXXGrdBii0J513l24NS+aOzXNY2VUafD3Bkxuhbtdz
9LwpH7dMLfvVu/uT4YYr3yJxpDdWqWQr7TC+hLXnQ9SNegR8VAkpcS6WhVNKLCC+
SsoqA3fVe0YtLVEoej2fjRQWi39dOqLo2Ehboy3tJKJMZ51qjMr15grPCsGgzQnk
ZH0pJgdDPrhkSaEzGOGWWyO3pC5P0OAe5RybkH09+CX4KgbVkD6E4aAItYklAnpY
TxHbSaE96vyQJRktAdZfbynyUVQLZ7JsWjCaDTug6F0ds3r9ORYX3tG2fRQGNnLm
bKyz66Jvx8jZuw5szPqDQJjYBhI1ZGqMkOYFUl1SwN4gAgw9F+IqO4oLqljDGp+V
V//mQRVt9Kts123gd448uZGBVfy1kPsreMSC93A9PrgEDuqc2Lv/qe47zMDTFE6p
/7GyHECRNrGj7Udw0jUv+Q7syXhSHsdWTVUBEqN3PPeuNGGbh7tuhzEl5YC+OxuW
gyn60AebThB5wugYBxZvQgJD35fYglf5lql8wHHmitA4pu93bwyYJjPTFW5SDKE7
f3ys07wUYq41F+UtFGUOF6fATfi6cBAN7Lw1MDVz5gGt5a81srG6McBVz+SRoMPI
n6we3bTIBPYs+YqQiefVBV14hC7jwpKIA27p9taVKhJhecJnuByM+it+0UKrY9nv
80wvNfmyy5EF3ZDpl3uG2om39sM2YiJyGtQOvSbyV25L8wsssk3kYbW/sxbZR9e8
R53JzdYVMFKzDvMOBWu3wRUqnhKSZd0oJHpzzmrSzsrQKkhQpHR0P1XOlnUUu4hG
nBngWtadmcLoEsf2GEoy2ZH6TsgKx9nwt2ZOGCACid/XhNpodQjn3QqvtY6hoXYf
4DYsmJ6vm4y4pc2evTu+INCnidjAf7gnr+yTtNCfJVyeK+U2nYc6fYK6ROdShbqb
M7ZpusRR0Jl0O0iaLvkvo3Oo1iVpchafUjwcaSLg0OeSawoeH8b9v7prz2VBpYKB
ovGyH72ciQ6aHcRWkJ9+YQOMeFF44HNqUeSPasvX4PDUBjLa57fqVKl0jjwiZaRG
PMaX/7O0BPSj2FheBVuSDYdtP+32JRYfSu8FLDIthIFMqhbyPUoKJGPMOQeDI/q4
Fz3nuduE4W2vMLOM1mqRPFQ32AIp1//dBaoGQlWGbEw1RI7wKQ9GIAEW3UXxd9Oi
8eFeWJ3Zt1RPMCtyc368jiVCgFYMC1hPYCPb/6etB/Rgo6FvSCN5t4Ir0RPOHcBj
/qSkqekvnFejbyGZRKuBjjx0xC4efcwVmTo5+4CJ2MvdxNcm4fItV0I5RXFaYcQu
xvfCXradXeCWcRc5reNn/kXiyCKT8kdrEyKX4m9i0/kYCyR4YUMjM6Oz0DbHaLXC
CLcaRijtErczTSM4MLgx5MmnhhEuTM+vRDIxQE1I6KmXjTX/O1zWi0h0WKW0dB13
GVb3VO0hbbTaSMBR7fKQSzJokBDJCTz6+F/vILcfWY9Bvp0+iMQ0KtoTBrljgJzd
vJ9Z4QSENezgd08qUUXTez9nPWs+vpeMdJI5szUvyseU6gADd4V8zlQO58Avw68v
wKfLTMGSujYY6o26pPhRHDzAA4MeYKtVlXFW7igaLjEjBDaGakA6TcFW2mJcvSZe
Q+XzQ249x6eSi+6mpwFsKCQcFH1FLkD8WSO/rjMayN+95uLty4DFUGadMQxkOxIp
AiAys/PVqTTtXYQuZkf73UxbzXrSCkPlYyeF07EQk0hfnDC+jrQzjP9KoBIpQ0el
OuQhRWI5YD3uvOBhmWI8Ni/lTIHqSWA5TsKNojb4Vc66DQhbBAJpLfsOZcfb8tjO
H6s91OKD8i3JdIAYL+eVYMDARjI8HgrWc6uSOKrDJHtSPVfYaHM0Q68/DMbdAfy+
3+4h7LnVHEFL2IR0q4V88GpX3DRqM/evYjFSPGGNUiR3eeLHS5o0UMWISW6y0AxM
/bwrTo+A1OtibLZJ1yhdbVSFJH7++fD3j0WcD9bSEIgwPjC9qrI8TybFjiEnpVS0
bAmixbC5WMvJ8SFCHhXM1XFiTReCKdOTk5hnrfth7Hkk85ga+42eJXL7b5r+4D1w
MiaAocen+Thx7/eSvAqj7qJne2aXZCoox5zpzMuPR4WPjuvp1z37oPFCAb5QXwmU
FF3EgXXie9vBimpktUs0GG6dUf4J49LxsV1kuRLpju8zwVSuYKFZzyJty4JSZ6HL
jtWD9oXLJjYa6ZM7FxT3FGBspABJuJQqef0MDIKdammHIuXpn8oGoW7CUUC2hnAn
OYQWYERkrChUC218hkR0PC+n9Fk2HvZlJpvbmJOkxyu2xK4VePbu0sEkgrKVQPDs
gnoC8CEM8107nPr8t8Vm9MrHJsySATWninnHFp+pjOR8/5OY4XhV6v7/86mtV5p9
wpbmTn3jVVW1Ad/IcsFjDHxTp92MEvO7kgifiAZ0zaUMO8/kOf1/bbonEnCoQ+No
01HRvJLxB//RBK5ghnfYATcWMiR9Qlj3/QiWlCstEgRHnxdzFFBkCtgQzjpt7g1g
xAisKrUwrFzGMl1m6C9sKuebaU9ICfsfceezcx069MdH5QIc7g1//aqN06DfdJSs
AuIld+m1LU5w7skrZDTjkVLIoqc610BU7a/gNytTCUN3L6QUC/iVLemuY+cDnGLr
ailctwZFjtIYLr1VEftVAXEY/QsU3A9kWcvwl4e7eFHaYH/GEPnXFB5Dciy7ITL0
rWY/6VX7dPJx/IPW8g+nzyoCNM7hE4hF0VL5mccTPj58Cs2uXbpF3Z1c0yp9PHuN
usMnekU79WEGS+X8ccaY5I7HefeXTOPX4O3+VPq8gPDr6kDZqFFumdI0mThsyMak
zo4fIl5B5lKnnSAporkAVgusCdCSy6mhOpw3aVF3S0dwHVf1FqAe/CSzYv4j8B/6
daFhN5LCLh+8JzXo7G6VRvTjHZZIqbqVY1x1rDwd95zFgdtmWwhVdZ/0WJ2gsMwA
HoiubrLo1bFf2ohjBerlstddXCov2wv3AFKiraHxUND+wROZG70GaGH0g4lDRPq1
Z/8NtEKMlXjxAKF9jd4aljIfKd0+y6zvhkrW2tRoGV7Km6y7eoQ7ZstguoBEWHT+
/fHYOdb6hiV7TUvocSzwO+24W4OXxEr5xJGzfRB2TeKQpUPn9Q5kMRhpqMDEfHyp
wwvhXr2MzSzAuhMwVD3EPEm8TtQkEB1CKD8+WictdsR685paT8O1UIeRx46032SM
xdTMMczICfGA/hadRnBF460N6ve0lcLPupWmp48YueHWdOAfNgET5So6IOyoQR+9
Y8n17ZEBIhMUw4ByiYhwjAmfXnDNjUFW/BtfUbwyJX3rYzDwIEPupDFwEenVAIAd
rfnunSLe2Zsl+5gdojxHMIjws4m2l+PR3P5jb2Fgikg3ntT9Dr4i/cjPDPYGuqSr
qg0ebJB03PSHXLp8iQ9dg5nf4EGqseyyXyjnMYnoTtLW/8LqYriUo5HSFwU2OGiE
JM2UKm4iHDwcNfvM347oshtp4JIsD7WTPpIPeH1vOgzILO9GsQ9gW6q8qEHPSqO9
JZ+2j59GC3qzvPLnZ7y54ooe5HIxiRepZUThjL4/00zOXo9811UWcJT19+E92vZs
GpDUJGSwQi/X9/YTvM/YWBC14StAbF9YsAZgVJ0LUaRL66rkRdageSenE3sVFLtP
4htQXSopl1HKNmhqu7Q6EQBs2HlnQISXqkaikzRuQbHPlYsj3aFHJU+0vW2q5mM8
RIxb78uJ2vPqWln1+WEJl2PgwznoiNa3fE6MSsB+ikcSvooM1gbZc4CMPb72uOAH
59URHVFKFD0FyIcWYyiIloxDQxV2x/gSj4MaVsR8JXp5kmQd2KeZOK0kg+l4cUty
tMvw5DL0ihjpWMpUjSbyIT7qeDh8+w3/RRPAiFgAbYwDDqCYBbQ3rcFP17TLDO8X
Xw8maRLHPS9+GmgcA4rp7q+IVuGEi/GQnCwfcZoYSII9E9zc+oxb5YjK8GYH81+g
IWR53DKgLpe5K0duT1EZ92JWbowD3RnFNDKpArP0hkomC0FN+/lQseQhFMeS6V0V
QR+WUwq2IY67R7fG0NBYl9GLtDBd/BemX/T0VfsUxVbQD/dmqz8uqED1TU99FjMe
9KG/z0G+ryVdDp2FkUS30wugYsAb6uUXDEwdgSVDxBeZ5Cy4x6Yv2rN27yYJo4Ex
xVYe15eHhwjuNitns5fnZZS7hvI+/zMd70u1nM2rWWhlF879/BiDF/zHEmxUTRcF
x0Pj7OlXQyaHmbNq8h+cJYEcgAVVaveokmKnJbNPU//9OAcyoHMwFhTlzCKa6g1e
85RIBnIEuq4YtsBYujj9sze1jS0FbTbdHMfDijor18O1RdU12S3CGY9/2XOhsBdD
tLyRwbpRoa/VezVQOnGagzzuWSGrg95k19y2G9l8X6ariJgyNLh7sDDqaMGV4scZ
Na7i0N/xVfX/+k+ZCk2cjseEOwCyRTyrOOi0B3YetSc71ObD3mgzNc/0mIeOuNGK
0brFwAyYJuRE+R6uCE4aw+q+wSR59JLvYTz7CLbCWGg/nHzIfCAtQVLbW/3Ciqqj
aI9nGdzifShoVhan1UAAJDadsL9FK6z1Da4frH6Bn+uJPoFEbmyTHnfeobWrWoS/
jsfAShooXA4A4exnEU37VqQ3/zo1RKuS9YyCO3ZnwzL0dRmsAJ/wKvyaS5DTY/ns
mLYwFTb+dOmh9C28LLh75Yec5oRF6rVEG1ZZKe/U5zkBHNgkM/d2wbvB0+lAccbU
8q7VNWNddKGE+1eBO+KD4IkYSNhtHbnhl9NgMWSOQhBjdjjNLd3Stw8pyX3fthCR
U33h0KbNuK4nNZcvGQ6vuDzvhMcOjs2FdU0fhUEmt8nb1vtEPLJQ6QwBtGGQD0+N
lWNw9auujTEBsu8KWBAC3inbrthMVCntMWHvQaD72pXx7Q9IpGA6O5RqeuFiQS7K
afhV5FT52jMm9/9tETFxLrL+EMo7Hr5Ui9LPyWgwbh1LzRVFu7skQE8ih2bl+e7W
5Fsrpg0T6TM8UHDNNkL6vO2pBPyMyIMH2ScfD7vZsHEogf7AHN8oU/vs8jKIXDoL
vCISKtC89aQLk5RtM6abYo6nPhnCOeKRsfpFl1cJYNGPw9O0m4lN/GSRAUNCYsjT
SVVn2cpb9P4Az+CO0msoqSvX3YwALWLgep6iqVcvZrZHGJef1MMkFUr5j3JtzVBS
L9tXb2HQL1iBllUglorQ92xLJWp+2doR4gxkPDm6XNIh9hvIw0koEeCpGX+9pSLO
O/tpEkEEk5ngxzEshJe8Yznij6MUAp6W8tTrfTH7r6HBHrcXveE+c6jdqIbTw9u/
o/X5aCoDJzOv1EoyT0o3Lnnfn6GRTtP67RGzjCmtmzfS19VWyN4rIVs0AvGxr2Nk
Zuv+eZFsWYUmXavc1whMJJgS+A3CgX/Hethip/gnFAUHbYe4lqhtZPGLHQGC3Nxg
myXnLELpKHaZv8/qwpFfl2gl3k5IiuCMhFr6jJ50keyPVUnZnue+V6KQvQ/rimqJ
DvWq+mOxxjyA0T0T8JT5xSs+pp7A865RpY17/QA4MH/guYCoZf3ut14N5LnV34Tv
ytmrw+NtOlyUDb7vAVTRSULV9ntxsk1lvrwZ9FRvfAe/bAiiweyiM2/66slGHjon
lYaEV7iGtD9erLNsc6/Fkx+/jK7/vHEsTFbMHag9wlycwcOgLFmZNtfKDmAs0Tqa
HBOJ9EaPuTthJTRWKCl2dlJvZNMQcDADFjt5aQi8tvDCx9n4iQEMHjzTRwwnl0sU
rYeByYs5faZyMKUtrqGwwAduZ7AadgIqOSOWPHbWtyp6DXIdUlbr3q3/sXZyVNI7
OEkwlBazYPjIHmya8nj3E2RXA5HVuTMLVbtrYOzSIbr+tEfSjSJNpfCUmp/9tRad
giHGfZOpDFfKHFZCD8/jHzY27ZbDxXkeDn/KZpmaLnZI4oPL58/y2POgEHOqI4wu
r1hwKrTS7MUW8+MdvgpRqDUWTVMX6ihU1NpSnj6dUPVgF+6MTuJ0Cj0BDS2rwvmI
0bkN90DcmLfjj5HgZSD5RsmYunfJVY1IjeyxQLSfDoGrdtYCKbfn/p9cAoJdz51r
iyRJHalVz0njNUjqoLUWXoJ+agkzJ9m4zKQvmduLeo6LWnlqzFDPKV2v+51uR/wG
dAizfMJuOBw8MF/wlTYyOaEBrGRQT83uYNpGJKZg/lSw//27731L/HfjPc0bw9/e
h8YUTG9AYJmXZN09axJxDtmuwLhv54u/4Dr8kLZ/I63mmeqWOI3+1lIroIw8LWlc
WntRac+idFafZdMzZFjlQz629Y/pdWaz7gZNd6Zbs07GdpOzi4rOUEm+wGqByGT4
oz1K94Yi7Q5yo+8ddFryQ0hZjkyQGaKuEpOkwjC43S7j2zdVLRCu7giMcdAan0DQ
eJhjIdmonuWJLcA7O4YCN+RW21a7QUeysoLG7ueszde6SvM0p2iNoM6UhSeE8ZeS
NlMkgQjWbblT5qzZZEnvxfBugSuqE/p6CdBV5dgQqctmKRk7AG+4gNvY0sbHmycO
BI7Be7QWFEg3OTj+9vV8P0vc7bFi/KZl4u+XABgLep8HaV8dD7TrCzebbmptKRSM
FNFEPABWnD6ONh/Z0a8tLkO6GSxRgKB2FBOYe/B0iXV9OBk36PcYVt7OMBXaV6qD
OfFNqp4MVKL2gzsoK+rR/3Ugipnc4JcpczjW6kjGoG7jGHejFd+Kyz/mRAgLkguC
sFAYy+fiKV3izdNH0cBLnU0S/Qepnn+Z4CB8zs5Tm1IxDtJ9xDIAhYrHed6qNyI1
X1eGvZPCSdU7VNyRZAYKIYZera8MZlcaEcWa8I+Fn2gO8SSI5mM0ymjTWUxNoWan
SGwHts7lHcT6ypUreSDzk2bq09354wnd1bIK6GeYMhPc+FJlorEgl/sehxqGWXc6
Np9U26X0J6tT3sy6pB0/kEt7UuywRFZaRBKdJpnErL8ZOM6eZZxyQad5cF0frFIs
M8yxCwiRPebUDRPn0ZeNxi/Sd60GmLgZmEkZwLD67jaOQCQD8Mbi7og6Dvpg8b79
gKaRN7FWDYObLiRwSYykjbDo8L6b1JLBHzzV9gy5WNmGmsdTKNrClkDYyLs6OSqy
28izcYFoFb3J7bt1m0xl6344IxsKHw3BkQkLFDaEpSqu81Hdz5P8oxrOutn7qVJ/
rL9G8ZD69ygW2D59JU/OPKRKu7bGFJxlu0+tVIW8YCq35/z+S95yhFj/3S0efNPD
4cK/EqUe0P7ccKXSgFwcwR3CJkWkPJr8thtVwAGpg0E0T1UZ/8Q/rAKSjNksaiZ3
slpTktSxsgdcwUyWN0Nxk1KIUwr9ug16YpW6fKnOa9VhuXTVnvGtvpkZnuhlHp8d
Bv8yNLLvr1rjSX8FiDVfG5x/aN7l7RlizprDzHASRoAFIUj+UKwNXiyTCXprudd7
pxxNaWTY8jwRzUio7AOCcw5NuXyKNCwHfdyEubXkbf10EDu2YqnbkMaaZRhEtTS4
a7rjfCSZWYDEXIcpq7n1d+FRyJ8A5Fzmr2asdYhnImA3JVhcI70NCy6E8YF/D4he
vp8s1Sl+7Kfvg4MedKcgFofGl1YAzRfoz2glNSMT+1CWAmwDOA+DEaI9uR1A7RwM
+vAqnW6bTmTAUD/NHko+x8lzXS4ts++DeOzAgT9uAODMYuVlAqr1e1h/7QwKwr4j
n7Y7cPFgJUrkivGeP7ER8JW2dDWI9Bz2qz2ffGoX7GSdheXrz1y/86pcrcJpbPqM
83HHZ4/gd0cucwQ0DgwnYVRn0H8ggHjm7wgfJIYI0ZBhQnNTlp3ZjL4j5JDG2rCe
cxlA/eAL/sYJmmWJF8bBoJ3yLROhACzRalpDzRvYOENJKkJPcnmiklr+F0QhgA3l
m/GD7WHosLwt6wJknWjO8OWV4KBI2hmQkQVX8umihoCI3vIeIvlUYKRlgqFM+QT8
wVVCgR/qRFEykvsMmBZgEDEuZHi1i1KXYjKmlEsOFX6nfVWjiMzBoGIDpVP1l+jc
8iu2NigSWNO3vLksmisHsofEW5QLjvfYL1H9uZWPwvKyWASMNZBATwmFqbkRSqyk
UNpSN5ZpcpxD80FYoHqe+++1WJ3F9qNI8Hk5x4K5e/vZ+bp5NN97VjLLIVZCGXlv
LDYMqohZJvCjwEUb8K2Qn3QB089ubBvUAZD5KNaaAg1FB6o4OcvcOTNujkTn7AI2
mP+FEcs+5nu4L7XA8COnS0wYjEsN6Oigem0NpMcH9Wqp48QD12Ng5EBzUIb8R1Q+
TuCObgggwWW3uiVJqjoj3uQQnQS4dXni9VZFkCLMyBmd4Lqq+uajZvbm8ADHUOGh
BiQKStI9Jb9H2vm6OkFjWzYZNFYpLMGHOMVXIXQEobSL/HBZNl9oCuRc7nhaJik/
0bbbCBjR05ryZPtE8XjyfjcOvBTLMLi6V4L8VFZMXu8Eyh+8P2Deng/EMtVWN6Hr
o5x7F1ThvZiPz5fJ1jR/vosMawVZ9f8Q9XQdeJfxcX9vNVo7t5TRspOn304VJEBI
3bMBrBzaObCfCOoz8wNDQNvMPY0sb/XjlvLsryx5WIV61Rzomt6umt8QlVD2AKtc
jtbkuWyOfhoEowGTjwqAbLdYsXdN9Lnc2OikSDP7E5F/+5176TK+WQbKKrj4raaa
T4PK1MFk4btSSGGDuiPx7WFxgbtq3+p/Oc4/pt2yJOkQPmD4IMKCVX/qca3IzJ5H
0Rc37e/ZdBjy6ro5ETGb39Bn/UPnqe7PGQ+ZODfoZiKdGNO4qW9am9nQrLFzGsRP
p/57ffCoMX7FfuJh/zETqZCZESH7Ls+A9yRHVTAK1v8hR1SXsBDnDtZs9yHTg2cc
M1GjTLXcCmu+0gdEun5XwWnP2rajub6f03QvvcCu94bkZQwNecYT2FsTu32dn8CZ
nwXtH8JvP+hS9AUv4M8cE++KlzSS7ve5joI5fCQc7mRHMKKP0UYV3Z9COofWC+tV
JAgjYP4GLEOakU+a8cADSmPIfu9D37CQjmcOMg76By1o/D2EfnxspGml8LvGKsEv
q9OX5vn4yzHg0OrkXEOhpvB2qKOQxQFlksqhC0akki3yBuIbtiMXgyc0qYcQKnvV
xNE/xpxPARq9MXRSh61aBNsXwRm0YSicb6X7ro/OSAe0NRp+Ow1llsA5YrG+BUnc
oLaeUZuWJSCgo7i+g8wU9k/o0oVCdwFoEHTFh6IKdaYkPsiMWfzGUR8/KgfBCpIh
acO2jPYUT29oGuSqSx2O6OSU9j7KKdfYWFHHEWUlzJRtLiOIR3Do2JFsUrPXivBh
1XmKO+rHDE175A4kIS6+ZCI1Q7jfsj7luFiEPz5eNXxMcbf8OUfsAPrFpF3JlMHm
MBEW2mkV7Cup5ta8OYTT/LQNNPjj6YEim1snjLzF85VEN14BlrTZJ1uV0mTCssLZ
Sze1bdf+u9O0EBLUV3tkt73O+GrD1lYzO37iobX8/VP404WGQF3P5oyJJuZqln4o
bDHt5iXnR6cs3mL687oJfdubMAJfY45ze965b+2U4nZeQxaxB88MXQmbSvkqUNm6
wGTslRQFoOhxA5xZu7zoFaawnm1p+kAvMLEOl2T9gaSWpqqxjzjJri/M2v/hD2cX
m0trOUFCmmFJahXz4lilFXpXlfIuieC/asNfV/LhjUp0bJJSWqmotQ9ITjer0v54
O47F8TY4xrxITBnzMUE3mIRrvo1sLVhnZ4kAMm+A9fp+f3/tElUOpMyC2yyvkEU5
lCsMAIJyiPfQT21E+zwef4kq1U9s0fZsHcQ3fuNb7lWagIbmA8ctjzQd/H80dU05
pcyimsG6E0PXl8OhTcaN+8BlP3qghexRk19+DXIzc5hVYdBpxMizWS/kLFSPb7MV
xpbHa0vY1HLdKcibvVnUWby8Yq24+GMRSSu0iq85P5/qkq5KS6OoCxhvKMoWV4Vf
GVrbZtJfkndr+Z23+M/ZLgeI8IlBFLaRPvL90l4ZM/NACm6edDBOjZFDCvIwsJkP
1FwJBAr7t42JdoqaeOddbU1Lq6s9t7BP27KJSEL5M3fnoh0WZykhnaNxo80bU4bm
grMqZq8gfmrtFgTIyu6XC9z8YjbzWyUPZFqRZhkaMbuQZlij397DB4JQnl02iGoj
g84gS27BdebKEvBQrNtAxFyy+kZjoU2R6aSR7q6aO2wwFhlltCYKlSaiJzcmMiIE
cphAC11dQKvlUlLh7YdCrxm0uTk/q3EN8iGd3DF/t2PqN+2iWDdfnTo5mwfZgI4n
+e52KKiQu0D3eK5OiJHeZHzGxTHUgQLHutIBd5VAqpLUwAWZVyhQgK+V9ip4bmNH
HBI6R9UCbahGDWBivsXamGcHRhWnZC8M2aZTYHPL/Mh6fenUdZWY1HW05T417Yjv
UOKAR4iLOJLtEUSBN41TMdW+WIY6tBvUJKGREt3TxBqn1wRNXay5B7ojHDDN4T6u
+CCdiomHOKMG6X+ZrSP9w9SyrvEnUKBOj2aBV4rDHsl2PeTboeGf9pbENcMWSNtp
cVT97jJqTDExQDfU9Z53COjyp61eDpJkDH54hTitozd/dHK9BaBL4fGOfsTQJcZh
kPCRpFFefrIJzjpyzFFX9TOfoVn/hxl1iWALJxhQWINq44CZp4GOtAvl1sYjbpnJ
dxCslgev4aIwgYAGS7vwwmaRDuj8rFwxD15lGAQ+70ykqq9PbM7jk2jLl0qlrU4j
P8LTSEMpX1hktUVciDZg3jLlFMMRzZPVe/O5rNiyrH/uKTtLvxi2TleS3qZwBz8o
jcXGLhS2/IwTEQrIvXd1itl3Taa5VtqHb1Jokq3La/Yx04eYpPolbmRem4DSdaqL
sZXuHTZZAcmt1W2tLU1BOqQpdMJI0AtYzbPbUfBSKhf2wpmMh2tLeMwPvqF80dTU
Rxd6LI6oQdH/S/6NIA2v+rLefKdEyF0wCPgfokP+5dDu0ZtE8LvzkvZGHa0UoM8b
gaE1P3V4cA9LChtDUAm5ieh616fLQBD1DyS3asRBCgbqs6ZGyi+W6c5+yz4MpRU/
RNF01si/Fp2NmWpR5/Z8t10wxzVCk0ZALaSm9+HWMLHJwKXZDZ2PCBGwM84tV3Ko
1y8VHQKXiU9jOXuyg02NaGY7dHpkWsbqbr+n5j8xFBVRAH2pVJ7Yy1r1trGxXtke
DKcQtk7NsiHi75LVwoHF4F/+FPjFlZj5BiQQEsVb2ei5sWVnEHZR2wb2/sY8Xv3w
c0AZl2zltWWV/YfZ5+cTGo+Xuo0QumsRsqkq1tQOUNC2ok/JaNZQDleVd/qwF4ys
JeBQe1l04JQsGZpPP9LSWfQmHSgsMXvn96E7XUIfZ/wmNI/94FgDAMonO5uNIOhj
P4AVWu5Dq1tTkyDzIzURfaxLov4XXCwTUtkeAULAocL/gAAMa4X2fsO6GL41Vc/Z
GU5SpOrVdiZEim6nf/4JP3B2YuSOhBqltjbjhtlWcQB/8xxGJKD7Er9b3twc1Cc7
3/JzlPwHODonUjAjJCM2ZuwwlQKkZhrUSxkSDzvV9RjgPyoH6OaveFAKTkurR4Z8
lhHxqNps7VSx6kphzQsp0RCZf3HWufBIV0ha7w79HqMn7Pc+M8KfHIj3GqBKsqyl
nDOZ6nT4xnD9fQ8Mi6JZCfA9dlCBsxUwZ6kiBhlZZ2BHlIaNPcBB3CyC+asj3EIR
iiD4d9ufG++Q0F2zZWll1669xd7gVZOKfaLbFDIIEgBikUSsBZmzmYP4EO+xZbvx
7LhQOx/UDXYtXi8asJrfB+xihylNjv7p9UI9NptFccS+WGjAZppqiD8PCCo3txXC
qaqJL9wbcyEfQtKmbC+pEyegLnuEApZWP/P54N/+hOH9j2F3PCWmc65P+a4I7TMd
oPNpjun7hTlvsPB0Dmzd02apNiokmRokC4qsxB19o/ONO8qyXlHvXOgRF9/Q7bZp
5AaCfNAQCAHrfqpmjE/zdzM/sqr2Wg8mfnKc3A3U04YbOJswjiI/LHMLf626VRAp
9VXWnoIylfH3QrVWwYAfW4oFfBc9FZ3wSH7sUTjNXknU8l6t+zw7BC1xFsF0ldSP
PeNzd/7zzUgsVQdrAMCPA/JLGk2sbloEuVoYxYSQvD8vEOMSRlfP3QV7MAJy9w2W
gYAAQC/GEht28yddS6WmCJNIygq9XOIPBCdYdsSQkPcSd6XfkfiwTrYQfCt96BnT
dkMLoeN7I2/2Aj4HN+OdhpkJ1jHGYn253WPaDsfaobM8GohliwBwb9xeD32bg409
81i4fKRdUT0RnLK7KXjz9M5zJmV28cZqfOsO/VNR7IeDXT4LrBH1C8gIk2whRtl8
iB78fS81LCcMiHQKT/jQbVkya8vK6owHagb/Nr3q57l+9NJBVNs6xav58rHHUcbt
5h+43dDWrpbQqcV3C0aGvXcBbewG5DP8xEOdA498MvJexgCwngo35iu0wf/+Wnlt
HQwKVUIdfwqUTea4zBKt8kpBQZf/oPyOm+Z5205I8JFjK1msmBzvNzYzhMeDHK9P
V2Z6viTWUowzhc9ODkrt23Jh8OCog3n80S72Tx5z+4ZMxKx5URMyMZ4NCbML8szP
dEILQcBkD+Wt4SLvQyhngIhHWTJ0j4OrjidLICnFuQPez4+NPO47tMo3c5i4lvAe
cFBJSr5U8eEBHMKlelILPRJjcFLfprMO1pgFWfkeFuUKnvqttNUo/ip/f0DsHfQ/
8PV6qmpooLMBf/kRWTcNUQQu8U4+FoJ0qp7oSHUGGCciHgsgpcrHM5jHKcDotLGo
0zRMOmJYGRA33e6dz4tuT1t9XlR8AvO7jvu07WwmmLfZwk3lPqwzXxZFFLOr0gx5
oW4UJ61zIDqImi8h1EteVbeG8/idQhEVbHtVJ/9v7UsdRgLsUliP/h2a5h9vwLjU
onNAsaky8cHsCpTKRfZd7fVqbKs2+2ghDHbY72plinUOtFBfuKlmwnVg607xTwS4
P8yE70/ePaVMWhsKYKjBinVoWgpxnSc1TBmMKsDHx49WaZ8+4OdpIsgzHbGzMuT7
km28GMn9ECEW+Yy1U4/iORylfTMWOZ5EZ+sJMX7GIrZaA0KnojWt/Work/X61JfP
jrto0LIhPyQrix4wpv2It8H3kwlKOO+u/ulHQS39dfo970W31N9UPQj3ITGnz7mi
/ot8s1J95hi8d5GE+TSGCe7w0cIvOVZWTuWZwL/l1za4vOR5PbtCOfTkpoTQEp82
0JpiJUb2dCRKUXgBnmH+/TAPdmDapeOaSzD2ZrP9GNkQm994DLZGWc8xTB9dGEax
w2rvqfjPcjZXr1pQnmXBn2ziUxjkSBlot7qztAI5w1CdzmM1d+RQ42aTf4BlGJ37
FInK/WN3bMiwWhNEYEPPTdBxW7tkRtwaLoDBn9MPXYRY0l+dZjlXrdpjqZIoOhKP
gqM+LCEZiJ0E1KxwyIBUt2JsKk2S0G7oC3CznepQpVR81iGrkF8tz5O/2f/eaK//
VphmejC39wGZI1ut6QAaNWLIN1gi1SZSVKFN1FcVGm9T56UC6sJIV5W/kF7EIGlm
5N0zRa0qgTYnPZYdfroAfc5y7Z3UCpwrNvUW0U/NBWahHJwMPtASGf/WjjIjdGoo
nKyxOUPi18Y0vZ0nKOJ6TK9Uzmf0m1qzNNjTCaWeRJNrpWTk+4hI0EYcGSevt0dp
6bLpYahpPgY5FdL70AL0TTwfPNjcrnE3n12lMifcW0jgIgbN0R3F2VdskwNxyIQO
0UowMER5bDuULBkLTOh2uriaYWAl+53O9XNa0iaR58DqBFOLks9i9j8RQTpWxH+i
T9nmGUUFX4tSR9sapaqzsC/I/s3smuY1HdU4HrWU0GCu+FLqi31kj/blBWHVrdBy
ehz9S5QPrxxsVPz2LkyNuq+gxic0xXW9lJzLIfOb8S6wKxd095fCnx4OhLRlvjjJ
q8PaHpuaG30YdTdcHwtaxpJtqLhSOlxBtQRxP9SYG4ui93RduMbtOiVEz1HZJfLl
VV5MVZQur/Uq6EuO903X+4lO85gKyK8eWJ/EhRt6jmA4p1GKkZ7YzTTHda/4E3Ey
2cb7g2z+I6aDXq2HhIT6dnDzWpRcNcoxuth/m2LnwnohaQsxHjDb0+l8QETYe1M1
vbkODPEU2aZcLM8+P0XMixqvKzM63+dwTrFf0Bo3s/UiHHBRZC3GhykujTq4Iyzk
Ceb5WOiIsyKoq4XJxM7//fs5HfsbmK8YMqpKPO2yrOgYUYRqXFjlc0QQL5n3CLHE
9iuLsLcFQbObOZrTs46emeGFEk6CBdwMBZf8st1gG31f8u4oz8aJyNB6Y6dJT042
/TJQMIunPHtu6O3LERW3qxh6+qyEBAnCgMDNvwaZ6t8hdZvHeB7kYq8t0ApTgiGx
hQ8neYeTcBJC3llJJ+AxaMjIqMjiaBlkmydUVvdt9tWJuYJ1y+MRzjx6+TkoHMN+
voa5VReqXL3qRqRypQnM9OX6Hpk52TlpIKykAGVBwWbu33SgZU/cpw6sCzF+hu72
Z1v5bnHYO/Krw/QXt3tgRoZAsiVMyBL5H2cnOGkrPzDnAWNsYaHWb9FRgnEYE3y2
lFIYP+hS9Ohkqg42S0H2H1GAKWQbpiTJ0trTqgnqtWDYnhhKLe1jsqIfKD6oXb8C
MEEn9EypXjcTYad33upI+4KPAdwDiDMbWUEa4y1rgwnETwki/TmmuGSn5FLESN+B
Rn9niubJFvO0BW45zT5EU+HYfstfdPYlGIF3qQ6//Ps1G9p3lEnuFziuvPCKVEGJ
cJLPpAFisXUK9qntyIC/pibhFQC3J4D5rDk3IgmO4BSQz9K/99LTAdCsrVC+D/Xq
c+5zz2IrKgNVXUUa02qUPVNR9RIpfT3o/aI/mMpwQ7qziJbzXqqy8Vi6nWjTkYMH
bdyLcSBqaUqHlD+SoC52JgP9Cy5eyLjJ5+Vp6vT3IllF8ben1znmaSuE84YNcmHd
wFVgUjNk7ptpe5Qx8uFuy4ItlL32tcBDiOklSz5Sp6wvDUWK32Sveg63cqFhMbQD
4+WlGx/W003fIMbQ/99A3BSXlxL1dRtDLyQ30sma64xPVCxcV3yGAjL8v9JykNLJ
m06cy0L/XP99I9qTvktCOKoJjw0owJdGEEh3bKmuQ0V9noWMTHU+YHSBq5Is9/ye
G/dCq4MvoGXVllT6NjNW1H0whIDnBDWS3jVw630ZLAM10qflknsfi60GyvkWtJcY
JsvCR00jWfu9ZQVVgLKAF444dSBQukpL5YIdiMRUleOqNks+UxF04PdXJmE0zN/9
vatAdDpnT5ZsSporVa94uKDQtvSitPNr12uA2jaBwQcP+wfx/OLqWiTF5rJLOHCY
4OGwzGHYZWxN4l4e1WNkF6NeteqYjAOn7lt/qwgnP6lsBEb4cRcXTb2x8oSkYj4U
Nlqb5dbC3wb5LRwPXKCviCqMK9n+R32L2lEcqzvGw9Hf7yB8Np+6DNiijA4J7Fxi
5Q6V5zYfROlDMl46ACcuGeKnRNpJowrAh/N4vKFDCz/hvI2GtGVJOfDX4NCQZ03u
pkWdi40V3ikO0sCVHmMGbLtf7qML4Gd9I9JChh5vAfSF9OG5vqG+hOON08UM+Ba5
DZHf6wG/Z1u0Y8NkXREcE3hPYOkp6Ntd8ZagxuuagQRAHb/2lz6CN+AOGwYFLjGp
YeLEEB43cwrqN3lkH4oss+HMf1dPRz01XBnorYtjhk9nIfwKFKohdW7VKZetwc+y
SWYASlrkDFdSTrmrToegQult/wH90FY7rSOQuedGWaSwSIGwSzzgn2wBPomvUry/
hGEzpHRExIkDZpMjQj3s9+swJJHP1oqLljEsY3Tue0keHu0IquKKRaXgNHpohsVa
EfiDCHhDWMcygaly6oypoBv/p6Fs5J8dDCqiYlKPqmN8TQDtj1bRsll2F/B5VObj
3/vNQujKgG9hDyiuURvcwBZCSUjW+IUEh8Q9q/EwKcj4mivLwQq6A2UvT8xN2E6R
s7nyV2Ep0SUBg00Nr20yhP9qYhpDeqsH8CjgsnQAjseRutD6PdgP/A9psS+r4sSc
stRdQsr/Q4rJmhZpBrLcH0no2fVWQ2DNiET+eNKCUPBNSzlmdYYlOU1envouXzbX
suz26YME5MRIzys7zQJoCNdA01+uxyhOmQg2b426Zgh8fCygCrHbxcQxQanJyECK
4jLip3KfiZLMFuVo+uV095oiqCk8UI81T7RJutEuvzOAC+1VxOoUNYBYlRd6KjD7
I6dcBov/QMgX3NMRhYD4ti9Y1xAVRW+rHjEIgVDVFHPd5hOkIn4RkXt5FYA2GoQL
p6XS5UbZRrcQhElCykxygxbecT0ZppPS20CNt+Pnc2vL6QsbZXyDvfUIlZCYHv8c
7yz5JrtKWK0wBvHm3FNbDwTdZ87ZMm/poJ8qfzDJRjHwkRabgipDsB9PSbSt3EqS
qGQLR8bYEV/T3kiznKFJGy60tJfUaKS/Kx2Rj2IwMOrPFOm7liO3q+uy+kosYzeP
R+V4ridIxFQtBFuItXwWkaZXogbpM/rewvfsI7Zhp3VaMFPOa+qR2WFtdYc5ESUn
1oUzOwMVJs14AQr4/sLtmOP+yw7wvPdnm0Ey21CEVM13fByXHJh1Q4r28huMFF9n
lqfZbiQ9A4OBt2XXZBL3ZUrJstNYMbn+LJPT6Uh7I0wrwcUNgzS6Kl68BncZdj2z
onOOrotMEhNbGjajwCA5FluB7OitDUiAELpqaEFhN9/IUeQaJ6lZGoR4mR2rEsAd
ifHIMRCyu/5N6K/WfVd0JhHKMCGN2pKhDKVLrP2GuhjWejbDKY0RUkXTESUBtgNI
j2pNBDEYISTIs4x9t8bmRDidtelnWwZOa01Myx4LoT1N+v6OiC4vtSqaHUinjdKj
7RqJw13hqlhkn4VKsErzbmylFp7R1TmwCvZ6JwuVCECcN07vnuG8c26YFJJ6UwIc
iJGOo4KKuvuZtXnGV1FNsnH2ilw6CfKS51yMcSk2HIu4NSmfLcqivHA7Lff9/F+g
bKu4P0zPJXXcb4EDtutPPSElHRmHJFIUIB2yeiTxueeGJm+K/VrXo+mWQoiK8HZu
IPj6PFM2/KnowjA/Yhf4AwZzFRMJDkzkwxgVpdscm+qK4kMeZoEM2AOH0imf55cZ
Mfk5y6RRNHvmqg8HC19fQ1XHgUs315uMzXqwfwzPROv+dDh60nUeTyv4cUmvw8eQ
C67P57hiYtptxEi9HJVsf8EXcUFwKPfqNuZhZpYAAkGXmADsxhPFTmE+2VE5O1fN
ItzfEV+Koj/l1j19Ml4YUjQvCPgDJb1vcFrVYugqh1zYBroQiFRLyp55YaNU9sGv
pUjVKjkKaa6qnkyZGspIYRs7WGhXEToPRtpVnci2v3n5xPKKU4w29SEn+/riAiyq
xQJz863J3Fn/05JJ1U5Zq1UuSyJeheJG/lKCl8b+mln4lfvlscVkI1lwRoEwfgd7
LanqzO6hZIW8yi+jzPBIbhKG17DL44MIKiOk4cbTUunkrFwchjXB4EBmZIKtHMjP
NRU/XV0oLPoY01ECMZTBps+9jCOk29E4einkW4yLvsSUF3y31LnhJoSZ1Om2VGzU
rjr5ptWqUyn+QYYjq6yV32leNfMH8nA/sT4RumcZ9qtDKm49xKpdM+agELn2Jxt2
zRmfIkCXfCwsR/T7IIgAwEed1lZ3XP33TTgsKmhRVGvlfExlBZ9YYe3w/HxQBokh
bipih23MhMD+5FIyKvS0GV1bCaFcoSmkDPLCs8jNZAC95AESXdCswl2O04R7WEpH
uM1BOM2/TuAPrKqZK5XldLuXy8VoLZI/qU3oIz0mI8mQHIyqx/FUFZ6tFsMYEDYV
xqH2SQ6peDRxNiltoNke+VzYLo5zwZeetDGvdP6LPYZ+2LtLVDdUFQj/1hpbdFeK
n287+3Cumpq7NThRLDm5A8yGFEhJmHO0YkyuA1xGr25o5AJFmKbllyDVZtuoymb3
fG1uhUYBvoxLpLIu8mo4Q6FmzHMmB7nKLJt6wkFeVngzVzcFMxAvRQIyrS3kgDXg
b8L374gRYsgdvXXRfJV7vz01d8GqTADOFkD4ZoTwsCfkQlBikaf8zKMP5EafNykX
MXAxKSDL40FtZG7Vm9GKspZduKETRvRbMv2PIn/CSVe+qqUilQbaApD3dV6a1Utw
gbiFhPJp+74xgURXTUzcaRKrvLxPdeX91KRnRfcobyKuLoQU5vA8f7MYCDGVxlTu
8c2nLorA5MDc0CbE5FF0CJPy8K2eoRvI/40NjVTBxHVguVEXbWsv9LWdMOYGate8
/feQplP6wOScHPiLNVaYXVzxQkte4f4ga1iEniRyd6CsU8NCVOl2BreJ//H6wkx8
jX7pAP30U0Qi9NWfINNshKyJSQ2Dmm/ZbaeS/AFqZzCQPENtnHE4Fnmbm1SWLYTR
fs7jF9blERFlXix9UluZ0O5zwoaAXFUa++se+tidBZ869sF0OjnGKesipzp4rYed
F6utCVRCdt3637IUDWgp1didQYN5gCKnmxO4tH88Kaf1dCREByWT8mm7GoSM3Wxp
yQmbtTsmC9JyXeVuNIY/BuzmOLjuL+Wz/ja2g8SxS0YfEcxr507ZekRy6AWsCe36
oOyRzsouxQIEtth9QQIrq8rnDAuIKeJged9hleFpCbuf/apA00nLrLgWEW5xIA1x
VGJP1P9lUDK1ct735jm+6dfnfRijJypaZvpgKEG7MrdDhstuFCUgiq1lKm7c6A9A
zZgbk2dtADYDUYNfE3aCffoJLKQwMunEJ0LuSO/y49OYKkh4yVQnX/mfdqAnGQcA
LlPZpry+5OAaP7RAW0kUomw4/OB110uYwJK11/21R3Mu1/lbxWzd15eh4LNlfPV2
b0KP+JkqU1B7X7UGBW4aP0P8ojcRU/SqPia2C/fag0KvlbpMfM71RIE8Rz/ik3YA
DUc7tsE4jxRa4La8Hlm96hsczIaQRdXM+oPCTxCWH2ogWkcchJAOO7M8OPLatffp
PYvEqKnspHSBNB2r8eP0SlkZQiFyVY/lCv+R8Ia2KcrHQaRFSt9Hpysvm2GQK1Ys
W7zUhF2KkEuu/JuQVZssJmHhaQS3GdVUa4/sdnMLtlYfBETch3sbCiTz++Lqt+Se
mX08Rz8/0y4Ge6+nnwo0WZ1amTdL3hlut+XYNYnz78YHUByCL8OA7CtBoR2MGbNB
6VP/zo/vi+iO0uUbDIRJ8Jy3qBcRmvu0Mg6FZmua8004cfXmfHC8QghxMPS1szw1
llhFJxz3rXExXtYWRvk+eStQ4olb2E/BpY8AwME5YjWZ9ugYKNoHYwTSubfn+mM7
b7WYHwKlvwi/MB/6nICbT9ipIyo5Knw+eIU4FoN/+bN5y7EDjLJI2vHKkd/71xJM
5nhPw4VnP6J8dPn2QBc4LrW95T2+vkwZS+3dZtiZ3o1JQB138534pdb90empZE3v
lvoQqeCsh3OMq5Syfsu+Vu5aC2eUz2NTujFtls27bdCraD8PilfA6qoWCwt48/Fg
9plb7Q9ja+APydCDfWSUA3JM4qOJhxlHOvbVu99edqy/q5kLwxnzSzZS4JkuvIyZ
CS32v5M4PwT4XDBZ9hjpB8UeJPtd5/rreBq22aPA/83GPY7ginF0xnZLazEZQJyL
WMixRF3vmSswn0POJ8pRICa3fdy0NJ4ZEzsi0WTZ1QI86aLdp4FKeaNAIdl/nKUK
sOSU0XpWMEJKA2HYbNHvIBgPTkReu+V3Kk9dsLpK9mJNnfGsaNh2ImBuX4L+9wOl
ioBFKsYqPu2scrlAyb1ezOyhpf2fTZcoLQ4Ht9K70y8+zdoWrfQsOBz5q6JhcMB/
Z/S65yVDV09Jj7/hULPYcSK3KDa3UEl+japT0UsOXrQODe91lVnlDAa6lP0xplI0
TnV2cPEbQtoGQevtzttyn8pfO2zoFt3sqc84WjE5UgWdoeCCspYYpObYQqvYWHWV
psVy3sEvb1quBAk+W0qCzoo1P5x/4GBKDlFjypoh9qtPsq4r6zGuf7hKhjew4VA5
B8pWkNHnovEezB2xD+9JYHkIuKJHgXqeK0z6Teq6tB/UCdPk0fm3xSeY9jqtfet+
IrnoBSjIBW7jPxWPZV7KDmSYLbwmwv0X5ircMhbZlz++JJTbycAOP3Ybe8Nqv+91
IySw/pPyfqrEyN7p6AejJU2lM6Yye+oMaD1rFU9VOvmbNFRHfddofDZWm6WkvTRJ
bdwhWdX/p9zMOcVKzIJl4Z50RKdvp51ugiohsNxm5KRCjRIXhC2owvnyTOveTBH8
VkaoUZ8mHsZf033+7A+vVqkmRkW3DYcl9OM4ABt3YgTURWggQ1Bl1VuhAGstrKAa
hV55OKeYWQXbOTvqlKhwc306zML4tp66gGG8Kpf8htKniTkbdYDuwOGgit5yRpQf
sWq3KvzOI0WIRa5QVjums/x6PZzVUnE2KWukB8zfdXgRX8Ryh0Fg0NZw60wN/PsC
ppLwh8IWEuGqH7c3yoNiHUiY8kZinZ5vwC6rirPcE19PJ1BBTzv4Ap6y1zke9DXd
yOuDcL9Rdg/GLJwqzAAhXN3lDlk9Ul0Wyq+6VsepWWaJI+RPWUVZkSf0pLCUCy/z
IEgzQ41ZW5mH1/oYVAv8hhdZEVHUronMfVBnYLbTht6toXiLl8kA0NTRBhibopgO
YBDMllPiy0RF73sDxqEfMkZJIDH3/jnn8KCgvJmHjy0cjyJM4mshUYwOokor0S/T
70XtBtpSagdnIOcerejNT2cUEw3YOQl19EXaqyS5+7ipQt1uHMbfLqcMx7U6ikXn
Rbx/dBIA03gnXByR9gU+mQNKmNLy1Xqk4rYRAbVunLcsMDZcq8UIaKUG3ybigcQR
2CB9K3Itxjk/KFzG5zEbWrFY/m93QdXtne+9IX9XSNoViTEp0mGMoyfLUZR0jNiH
4AYVLPpdenBzkOuirL1A0Bbg/KKf1ymJBH/yoZ+6f8NKEsTEeF0lWHH1KVfOx4+K
PtcFjbhnpvuo11OJ8QsAifRN8iGXboSvT1q5NjhN8zNw5EoVe/Z072h2Lx7yHQmY
B4fbUJ+LcdQJR7HVHAx4OqsTYY+rqGC7bPpJASXvFfzQ+4TZ0v+UHUnntgUgcKsb
vjaYKXL+trE9lv6mWuR3pJSHnpUg0ZEKfNDj6caaEHlhFGe3gjOnwBsjcecVM6PN
aqq1iia8ykg0qQAA/l87qaRdT9sxGsm3Fox180dDCjSpsFhHAcqqYHD+XrgOiQXP
iMlW0Kdb1VHit+yNoLnHhaKYuKpyt3DmyRuxrWPQNKe4HhQjo6t5DnQcHM81Z8z9
Gs4O8NMfA5fLlP2/jz6NhwUE6zUTvivfTe9DLm4i8hNw3uQQMsVFtlC857na8Q9H
4BWKc/A/Edvlsq3EPU287y8rc2mykmqPCFAeERhsZpwMIwASOlTvuUImao+PQxzv
nzpMo6nFVp6Pa62MXFLn43u8N2k2DcvHUXJ9dj+cwXitDpNildE9DBXPD2Bd4O9e
qXlBv4JltBMX43gP5KQPVbTjQ59/jEUX+5Cyxc/U7RkaM5vRM9FAXA9H2EdOwEYy
2StFcMizkBBi4aV9JqKqwEZbX3z3XMy4pPAB3kVa5+kSJyJ+59lsAI2VeY6ZkhPw
ikz6FL5md1hM9z+/h4c8BNIRkVzsHf26mDM02vUV9aZnjIDZ1UtZAApM4rcLDgrd
A0MJyHWNjBcSaHV/MXG5GHpjNR1Lve+FVbx1jOs8sHzv4dCh9IqGcI8tVkZQOthz
fTQcHTBSHYrQHPb0v17iXJ6FRIEGKgyOtGWY2YnwRM7vdCahzZHicx1lMrr/rfgQ
i0wqJXlto0JkJiM9rbAdojnlLxuUHnB70OsagQIipHbBtzpqzsY+/nXmnKbigijt
UBYmzkN48WEXoiZtenHtyfCRVNOXdhxfkGwJJO5TiQcsaVmV3h/nsP86No3zfPmF
68tPymLIMtdZ6ZWeFOjkm/J/ud7Yyn7zye5/dxxx9WqrKcEwn/I9jd0jfUlKO2vk
nUcDyjwGl4KWNmQk1YwaDwsjqrkrZq4NQaOnFSsfR1tOcgviHJvnwWEgIshUIs78
kHdwstW3Ny0aEENx7pCKtBeY5SCAg2daYvPB/kU+WPTaWGZGgpycSZ9INqttT4Ol
sWdWTyPFPYeyZs3lpo0Ozvy7/acnSHGfwu05zHQvQgc/qKV2jQu+T961Hbimdfr9
agTTng6DOQ3jYLa7qic0Uqp+N2US3RHmKcJEl6ie1JzZm74mliUPVjxcZ9Xv7BmG
LIxKfLkcfm9gDYKHD6qW4BerWyB1wxHVGHLAwvzJMGVOYU7ksLKKImcE9UrYmbKZ
OtZAzHA7H89DRIgp5gcAlqEBBrrXosWwj7ECjjjtLUBNg0iXxHcnC64tMUA6nl8w
jPbhgPLf7hTCGEF4q+s0ap1Kh4oXtEeAvWT1tRVHp0TUsVKpr84ZK9ohp9K/Lgs5
xgYtWbsoksvVV9a9B64h3VSLNZk2cnJaNUFna3ec0AD1EmovX+LFDfa7cgn+Ai4D
QBfEWnrbvmzKsgJhIaOn5rYVR7QDt6IR2+M/0zRvBsXjJ5usWH1SA2q7NUVZyCQ9
U1x3M3povlYT0ZAP24RYUayF6KqZ4kiFFiEWDcQzmrQU5r9jgbUCgYaWUDVQapXJ
ojGWPjlg0VajnUXOuDt4aHKxWSPrE3WD+7AssePEoZRfUHEMThDM4nSZeaNdp2Yy
By+Qli7E3WVYVewunv6w6p9GX6V/giZKG4hILLt+luzVX+6YRxrUtEYAJ2NQQyJN
hPAjd1o6ND6C6fj066z5Gvl95HQju241lKhTO67OgFDaCQe7RBYRW881H1uH60y7
Wt0q5xJvymYz4Nz1NTzM69mAGo5FnjviIKSXN86tRKlDS1rqYZs/VHL5hfdADwJl
grJ9EfYL0ka4xwxbQq5YBOt6P8j5KF0eXsxDFq6lT44C5PmPH//hFQ4WQ4kzVXzw
WT0ZwiIesPbYgXnXoBMUlVFADgKw+gu0hCF2aGQfbVHb+X+VcxqfyWr2FrTm6Lo5
m+pFiAzO4013/jz6pW2CDWYp9VLvVAWm6cNoPIM63znFB7jxcfTzczi/SElxT25M
mnJeRt0729XWcKkF7skNfHqtEE5FTQ86OznJkYHED6VCfxPXUalAay5E+4IzRF3m
v5HJyZzlBtgFw0uDYa4Z1S0IvPiGoQ0101g1RsLN0uNK9n5GKgl9Jzqt5Y/VnSC1
qkCZkoBrW6OAGUsLisWmjuf0O4Z/2UFQjCNHzA1mnC8GWTGmQIw+eHPUva5iufbO
CbSHPZglhdrdTofXho6RpU4Qv0HXRbBM0EfmbciEEIqqjpsV5XUdJBa9OYdSzLcv
PZHQBevzp0D2Sx9qmPJY5IRUZP9ppuGTHtQL+7GkHP8eFwXjaF6up5AlcqTZiI2e
lggqhyJK53EQtraDuB5IlVLKaoL6E28/JEnAVQOvmyLcJMvaVzz8/bJYvM5Y87Yb
e4KbuvCDRv1pjTyynEu8J6S6LTCSPSP2KoEM2wktb7TB84S5huiF5zAn3OiSpTyZ
Y6VZkBw7ozVoPU7e6N+6+RVACP3gi45aPtQGCDFCYAfzhBMz9aV3Wd/RWQC4NMRM
MxGjHKpUwAUgT9AryfCaGDiRaaMX1UnXpp5wHvrkIWEbv//qGozkydbW8C/HQ5Om
9QGHGNvrmbNbN3ObwoWFfx9lvXPi6KYU4PDJFuzsFp7Bt2xWFKsGxLXqpot0Ojt0
OaO7igKOn1vuKxs3mUTZEEyKbdQY7OHs9zSf1a/U5Wi0LGOyvgQkT3oegOgmeSeq
F+LvkrP5MSHfNytHTBW5nl6f9n6wcU24YsOcUuNl59hbxvJuOjUcjKq7O8WLWDFR
69+8w/j83iS3BW1mpR1lDD2dzM6Th7ag+Apnm92BQKzqKn1fFgFMcQ5ww35QfcIz
2FqrldcijLWYoPwc66b+6P435aOZrUb9pubL5p8jpZQrAojPhFFXlL0FScxbY9MY
S5ZJijmD7QEXwLFR0I7wLdbl3IbSH6Qwnj79S9crkylVlP+1y3lMWIA2vQIvFfFY
zRdUW8JIuV9xADtf92p4hWZ7qI55NiA6//GsU3QQJMKruMDjLor51flFq+qPW50w
y1SZY9Ly8VO2SPlOzCqCfTSBeHG03LZmSJUAIi4Ksf2iWH51bQgJERUlM64OCb7U
QlQZxu+aqNuXrsBpBwAnhxEak144VYjuP1NeglkZPz4rkIKZYNkPIluB53ELGivF
6NyMCmnykb0aojfQi3fOaB9ZrjDPgGay49nWob9rHkY2hJ71F61W9xIRyUWaYwHF
6cg+blrzlJBXi0iRDhixbnPT1Rlg7u7NxNAYwCixgj5XYCkwzjOK/PN95e1pMt3P
q1jqWuHqBxfQ3YWZzwFCTF4cA2F1Hck8ePwrYKwnZhwpC6aMfYUDiyVf9z1HaBPr
PGFWKCNOkNnsXM+aI7LvLr9Qk1QC/9XMY+o8Y0dTMm6GFbBxQrRJJdFg98dRz2+T
sw8fQ+sHsPh243JrdkMYPPyBkFKMfdMGdTwwB6DxFqVjMsE9CCDZUNye4gISnA67
6rsbvecgv0begBqKO+CCGDWDz244mgkEysXbEN0Qj0Rbte/3qn5jjTpHon9SlpHJ
mm4a9wNM61OBr2Hyu6S9xzBG1P2HOiXvVrkk3tGa6f6dycOl4xZ2YADRndCNwYHp
JouIUxS/f9O25xWM9YXXIc7NZc01x7HUI5ZRMhjAAoO5yeaAZdDn4D+i6vQQ/AN6
xoZFOqdZOvLOnFh/XdV7gG3hualccn9OnAks80ioTkBlUKejs0UVlJdMUDNvq92o
GfGN8DAYZDU+HOPyJXY/J5an3+qDL3kBsciniwf2yFrJv2jA1vYfidwQ1SxmoE9S
qyN+obavA9yBoHc3hcaQUuvqBP80a6XSOnwKY+QUd591xOoOK0tRpNhJyJSjMxDM
xcHgaUMln+C+Kjb439k7b3cAkOX6U9+j1bk+kOG9TuexLuVEr/YgWBnJWr8c+s1g
9t584eIUiabDMHyutDy6KUv5KALsifPdVeEzdcH8lhFu+sU8PkoIsXRdnPSBByy+
+aUMgID/7KgLx+foj5D9M8OaYgVaVcHfAHS9xTQbL+OT2vXX5Wur8oStp8rIT4F4
jZEzbx/cwk0Uf9jDfmLUWvok3d9YFmF6vQmQ81stilWjANHDzzogAK74tuQDPAWZ
hB/RR7W1uD/HO9f/f7wIVnsosJUjMJ+KBtfgpv1TD230UgdMqt4UI0dtVlo4hnp9
Or7/nZ0tf5wha6Ofc6DidP430CWXtrgosNfE9qNTjggeTpSYrqVpj1jMQdVz2bgT
DAvjOFx94EP7/elQP1C5wEJ8Pe9Sk86hTL/LpWFk1T8izQkATrhjWTd/02owW9Jq
oE/5gNi2IZTFVdvrNziP/eL+VN7BGjhKgnN0rKxMqQMvccyVR+joOApuw8J5Qs3o
TsqUpRzhNCxA08jvlGswx9wfP0Tpx1YNFXsVVMoi/6NYqHYoadMvNUd4eXJOhD4m
GCBUB9K1Pwwg2Mu60P6LK8aMlyQRANbZ+dyqrIjZkAPROUpjgieFEDetacltR9qr
vBaAsA8RVLjbVL6VnyAjcNHBQKJMbb9m7jtc2ibTLLQoZUi62BZTpvU5GQQwkQ4v
KkigJEaHewKeMvwLHC/9NKI6UYd7cAhk1/josjB89smRjoMXm3HkZgdPCzd6r/kx
K2X1c/U++Hh44uKuQrTBoMuYIMrhgKOtSsu+2SL29Z8audoq54EE+Gu2fuydRCCj
0zGfN/gUFW4lyBDGM8Y8fh3zoX6+Nb1fAjOtpkz6xNCB+l3Or7ktX8K8PcrQQ5k+
P6Fn5ZpCphMAS7PBgfiIzjRJmvBkP4W/M3eKFVZPnPy9DoqG2QLpU0nDXGtFQ3u0
cHjxuApzG7hEm2kbWSPyshe14bl7yd027N+/goJWckBkefXEgaqPRS3FDjT3JPRV
e279t2WcEg8ja/nDjhVNlItfGId3v0jgH7Sjd/NI1wHH+IbOMIKUcgUvxEX5tZh+
C+H6BsjeXFDq3fnxVFdbr8KVQ7/w7vFLhnMFYvU8zq02RUnO2xQI2u4Ix3vpPUP1
A5KZnMUGp+q97t20vRN3YD5JL1lO9Kc7LuhWiarkY46Yotd7SpsKE5XPfCCigKkZ
VsfrFGGz2yZ+dwDJuaUUbNiBxWSPdMNOPEcOFLlPJ0m7tjIEL+yxYuzrRxWn7F6+
1PdcqfErgo+FhN4QvAzBEo8l0oqkNMV8zw39SIQT8fyPsnUekdiozO3RltUcHW+f
qA2WbQ7SlInLjO80/ae/2S42kv/kA364/XnGboobIhJ5UG0SkTAnbvTEsrH9Wwtu
wGWQMCTqI7aOsfSGgzQNdELMtx98RIr6RFgPy0TKn7zX5yzdlzlbqeFnBEUIlHw6
a/ItAq40G1qqxmgnIyU6HhzhrdV4PppAD4vVP7qh2wgdWsnNT6nSbIQ8Jiazu8zj
6QLR5GMCMjff/bz+yWXfYP/sEtQxzOEsXdMRoqJEjpj0CTmCsGXT4o4LqtOAZRSQ
w0Qk0XAx3Tng02DrbbihA3fuIt4BDwoyUXTXMlHBOwR58PAoszl3cXoAZus7yBCZ
pWdLa668IanXuzlAANxf52YYYEkbxAZtetp7zTiPF2dX5nCNUv+65y3dsOgSxZWQ
3ubHddCVxo+JpkJl26Dp0RrLGOran1j8pQDvRttLiBHF93L5iNQPoydqj2XG9NHP
92QyN/Y40AaDByXx2gFbFd8BBJwY07PySs6lsm9u4/XXP0Dje4vmWbzF0qU+ql9L
wUJ9ArfQI6rX1pEdj1C5PzOQTEpx548fva/AJDsWV6X/ats71gNgzqVdlqn6uHoD
37M7BOLe9hhRIR8Yo34ItgROSulg6eZscySADoCx6vFx8ICYnQ3KPoJ238g0GEw1
UQZW+fZ9d3VCubNTudSdQ5Yptu/Esp7nPJ47WrE7PophJzfFgejUe6bwXMWL2W4t
ri7DiCpCLVT32wvkAEjcKR66tZycmKjQ3RW5hwYJGiRBP6aeI04TINIUTZto/S66
91HnL82yPnrmcOApX+G/vjSk7xzGzJZk/lf2t4OB8xnHD1Wx4XB18QmCVFciCNTY
jLtFU/hQ5kh13qeP6WW/QifN2kHpsmGSjQozMFirNWq30fHkOeNJp8zDYBVs4BEF
DAeryowYgA9Vo3SpVa1cF2uU4XTG7+KSkQT4ijG2OWN0kuUCK0A7zJtgA8BAv0Mk
lUdzrKYTwS0tn+/M10vHeF5X+JBbpWCR3WNagWgeMyGoWvOh62uPHHMGCJSLi1XA
039W1oaSWGFJBpnFg/8Hb/ulUS3Z509mZY31lZBQI7jnSph1ad2a6Vkauj0Sj7hv
+cR7ZnLLPolZxK6d714OYVq3BS0LVrv2hQbwptFLz1Aw5pm98qLEVPkjjZtOkEfK
7HHsBAWYdTXGFBn7KTOMh54MPySo31lDs9HnBG4yVvefZjOpAbdNcOF4oEJcfUXD
6hcCpBg7xFZ5gPbrcQIPj7qD/sP/ENPDwBXQ8gwQ5FgvsPwijfkueDXjtlM/AHWj
sMi9+Cuyb+mJOSyM7IrOLiYpbdLKyOGbu74w1toC2HaqNHeUGzlmCkAXzt5v/cSQ
ZzYvFlpanZgjur+lX36xXeZN5A5iwRO7Oox97k9ZZwNOZT2e7+HJlAmbeCklJ/pg
9Gxk8oYKFulNrks5jb4NRQf4zlu0n1EJQjiklFPwUF5TK3LAVrLxm9XHu0B9r8fe
Aagjpl4Bvg6k21ySKvBDvyW1NdqOxOM6Nt1DVJxzVXwKfHiK7/dvxCfnUiTBHXwm
RuuRNpmytvu62hgiw6kKPwINzfwni/2UbS2ly286Twetl7vniKnKwTp1fwYEAz6c
Nr9EWcLApmSRKgLhVrJBD0H/GbLD0U6WHT1MbJiCv/2egvNn6XxzixTQrl7+L73z
hjpddAqCx77vxiFP82rjEBLqPE5/TurAr7JqmAYiIGTSW0GFu79/csxOxnnO19hF
aMSGN9twg6b2v0j10COLrV8EOxREU7GuHpvJwXU/BzDPKPHViWQyhaeVHqAL+f4X
PMN6i61nwJQSO8DolHqZOmOnugd4nM5z7qFk5QiuM6LohmfTOCfeY3hfRGOz6e15
hGkgh2ezOCifavIrzMAw1oCVrOnwZuk0gKBPLEaWIVxiVw6nFTxnniUbuzuBeT0h
N4CVIMarOCwWjBzwaAdCQMT7Nqs90FFXd15PM2LxSz8nlPRIr4sUSDfjK0gKiFZP
uwquKGpt3217LiibDJ1evnDR8+0EkCOoKdIbEleSNUnyT91bzDNi8xkC3wSNaZwg
qIKvIw0+Nyoq31gviSevH2IDbb0JsBgK/7J0Sdd8Hv67w7Cnu1TaOWd6XDe6Ri9+
/gkNhHBDcXBRgdgnGXoddT3Sf6YpIX7Z55RtCjuMqKJz390n6R8ktWIu6RcSCKZG
uU+Hv7pqdSPuhqZ9n+cCPAPByKDADKMtYYm2nlvWS7FhH5R5PqGlFMu/wdoGC97v
DLBJnEfEaFI+C6dFSxul00y6/mHi8ZjbCW/TnnZ+hx/XMFhFsfm2seuY2E3ojj2o
VpwFcdnUUaT8l/VQsnhqn7KZek1zbJi7GccEkd9EnWNRelDQXn5jv6P9l/77NZVm
lIj4vZh7WLWu19EDsj2GpDRadtqzWAkg1nk8BH0b4rSsHYvIVKGf0wFHzyFV/9DH
IPix/8RJXf29eX2GWAko+XpAJo9S/KswZI6aGDdJ1uWYHyZFlVG+6ddz1Zxu+umA
S2eb8MfxTGZDWu/Wbf8WecQ2mEKYZ1LXwl/6nzUNPcO/KniJeYnX8WrsvTIZDYUp
Dc07hYsqVrHe2ja/6NqJ8WlSTeLrj0qYUnnLXXyBjg6NJTtHrmBrNixh2wA47qnT
TUXIKZgXw1YZeCd8eS0X3YR1TJFKSj5F00tPutS/xUETalW5cN0AMHh9t2Z4aBd1
d3tDR+pLS4Dx7hJN5SOJ7uuAQ4yX9gJZxyuFa2pGcClcW6l0vvxwfwBcjBSfHz3Q
6GPpCF4Ws5WimABZogcFQ5tEVSkPiYk7EBtBAmNdkdlFyV/oLwrYcGZE15gsCNrO
T+CI115IDnNzLyKVQAKCI8Hy/Vav4yzRQ+BDVlHIBDyaNmFJHG75kxSJ6+5ifR4Y
RwladNZm1ntLuWUxclWL9RoNauaYmLfZvQbyw2/Rk4VZpPEGeSVE3TTB8XiO6gnG
cG4C1Mahet84LOW70qLKQ6R3W08qPqBa5BzGAJk58cDNGP8PB2+5d4PPGa5knLy1
NSHCL+/ni7rFlYvl/LM9yEi8pzz+1z3JGap5S740toOCUQvk3LDvEKuT+XAUaL7L
4ATGk063BEdm9rxsfcToM4z/Wta26/PCayenWfvvpmkfXgwIu3tA9vWxHNQmqcMA
k7YjmCv83cuCdPd/xco8mQC7h8qi+KACsPjr6MzZVHB3QQx8tEOV75Bgu40Ur+ZB
Ulwtjh+i0pXUMgYSLD4w8xQLXzi224PdUjTaAsbP4Q1YZLaXvg3ItWimdP7L9AjW
56aX9b1kdrNBJXLZMyhTxPim16XPuUIBO0BbbopAfxJJOawpJWLkiTJmN97OgyKY
d5y/TK8b9TDGEVtKhYe3SSfBKeOX9G3dcYVO20wLFNlC4pLhduBbAQcwb4BooatR
xQJhgR5Z4XTOEo15iAB9H8WAwPBtKmqXp4V0EwjYvhue49P/l6LH//gMdWmaf9Ix
Y5kpFTUTckjf6OrNGVeopvIJFIBuAfoqaKVolZMtNDg4I8A/jU5uy4ipPyi+PTXv
7jqbHCeRxxxYAJLybuBn3G/OWT5ydH82XFXGthEmeTeRw/qSK1Q7IkajNfGqtUk5
wRyswJw/e+JyzLolrOmnc/rQsEEbcxVs170jK4AXm7aGHn2tClvYHrMpm66J9ThN
gtT5Of/4ldwbiMZh3hYex+LH8itUBeLKJoZHgMZjPzOkUJdt3h9gUQzzxo8yjj4u
Si9E7rLZi2dsFdDgVDnxD7iBjfLhPwIJAiWHuzheVA+bv205qbISuTMCPasHmwam
duT2sUktC1c+Hi/CLRpO0Y3xzixqhTYEvex1ooHGC7g58QBukk6sdVRMKaC7oIGj
9AhoTfxHvNxbGOEbRPdKAvVS6IzZaEPrt/0AKX4H5p8NPlFVjCl1t7ILwa0df9RH
iw6x2HrNq/uStt+yDUwkKk3D4mEMmARvI2jEVGDIHny8g6TMb14SGy7jVgIN6vcP
72NOdqas4xlUtErgsr+LEMW02+T7nJojt0XJArd1a0gHz8VZsD4nVgAWoTAdLdLo
3K0Ff5avLmwceLEIIdwtUnpPBTlQrvgD+/FYdVWxnudXtGeu5nCMZKtkA1sqgY6J
ssU6bEgYLTeJuSFso1udii/4978pHDA4GEgIqj8I3S2QFwHlnR8/WGgmACX/jijp
29QjDCds9sK3CPWav/ZynbOhbnlxBSoG7WXg1ADZjgK4/5Rs2wHL/3lKTK3vPLcQ
uquz8IYGv+LKyKnpXQHqGLMujsH7sCi3FFwot44pLFFBh/Qo8bwGEaJgbBk6wp0o
pAkynLrZRRGGemYr/SX0ICo73T78mKySqUngqgzTctpDHARI4CgpvvB4Uj/0khP+
Yd1JAeNyjeV9FuZoOuFYjFniIOD5hs27n4FS/r/Jn4duSwq7zwzLFWoyZo/XshNS
ZJJAwNXduxGsuwHSXNzvKqn3kiFDzE+/Biu/H+mCtiNTjvtY7+7cQVX5sDctoKYH
lffJOCA1+MWO0j+siTiUwHIbFzii9ro7wrnEOAAdZt1PbMNBQfPJRhp+etcJw6E4
Xlk0gF+CKY0XfMnCKCdSlRQ5/Hou83LJrqcuumAYIi4AuE2GSxhAWXf56BDncY32
bhp1iEpEXqdzLYCl9s6hrJ1mRKVbMRT7xHx0AnzMLWGIFU/D47sU89YBBCpWC+kk
qEaWnVJReSUNEskYsx86+qJmVpM5UocGzXIfeZhw19Z64UQFQDnuutN6bdzf0aGN
3Z/fefaO4dheyn7rTmLtAHWJaN3NvMNZxLrPxMEnfeUksrnrwOvOHjkSRhqnjiRi
WKPI3ikJBaLf9CaHiZcEb2IKES48/u74zH7WcAktvXAHb1LUYI3zGCylhhoYF4hz
wzsSst5x8Y5ADtwHNNTP0YvAOIoT+mssf6QqtD6YMLiET5q4ONXoV7YSbrS5uGbI
dmw9BQpW6Z7hw0LIsYPMRIGtv1+TxBLiN87kbOTnNeCuTsTkNYYkUo5qbl6Nz1Mm
dTDBRiece0w22+sEPbYryTq8tn632u0vyuD/uHIh7HLi2cb+E9FeVvShPI4viI7O
G3Pbj8CWJ5oiVueAs3KGhQvG6Fmm2yqbE4BId8DgmqmYFYCl/b+aSGh5JPO1kxVf
cwvQiKTuXnH7k57YHzBy7sKv0ulAy5hXkyjCIkVnBpDxI/CbSinwJ/2ymEmH1Q+v
Er7wdKHQYMtBUqC2gAAW+ddOA6QP493jO9cvY1rCAxTcvHtSb09r70JgZJpi0qlD
0aDuQfhEQgu0RlOsRB9QDsJeag2n+9hwpduksSxsIkLlVsGB7W3OuekRNqN/KnQK
BMJrm3Is8NrZ4RiNDgr6sNzlVEwC0nRF0qMagZuvIu+mK1FpiUfpS3kCAnItUwjC
JC2aeHuNz6mA/cDbO3QVWZOEw/8RHmshKYIsUs+WHKWgi9VRLvUy0dVIWyR2M3mu
tDwIUJlF4ZxlQqxsdHp2wSmuL1BiPaDcbQvVGUTACszZcRIicK/u+SkqJNaQC9L8
xi0z2oR0aPFR79cAHgGjMng4y/hcmEvx8EmnvVkf06TgkliEOfGsGJc3JBeHKlFF
WNjxluvPVAUG+ICq1zLY6INIK20THmSVxpFwkTJdpbUPTs1I9sVV/71QuJNpK6Vb
EId3n50c5eWa0Myj8n1JyJteYyXIlyYtBzj/b5hDQoxcnLrDzOXN2Jn9gYzVvHod
8MXpYmf+lHKcBDgOnb5mQbwARHM/uG1Lt1o66RJlzSs6hgK7W/8KZxYRYeFa8hf6
rbq/U6Tru9jnQpRD2F+bDhHepVixVi8uV8NyfNiUuyLQxr2ta6cHFMXRkc1LIFg6
H6ZpKnJ1ZBHsTXnPEYymwZFXpDDO1bdcezDgzJXiSxlY05zKowsPfhEm9eCdC1ri
MzpVHW7epi6NbFt/7oYTmL7Cs+qKD5JYqz3ktT879J1gt6k650NWQbLdr31jPpGO
lGtICHP99F1hlS39M7hdJU05GDxnGdTVyPKQh7dCzTLa3NeU6HITEMbXE9MZl/OO
08ZAa1l4v0kVUgQc9JNBuOXYVnqDeRE3yxYjrD3GS9BNoJIva/rJM7Cs/m0kW7Qj
PGDX9gkptCpJC/o1VzBxRS5rskVlcOu6WL8p+cUsSifDM44DJW/nONpmfGe6MONg
wJiQ75/VFwuO0Ru+brUFacevfY+ueYXiq/C0kfIvkVE+E+XNd2PS5NlFntdEFqRw
hN9h+NhM6Il7IW10AA3YKoX07n6zQ5eUxFbqSPHH/3bxxyWWF+6nx9gkOSFkRrWr
kogEVAkT5rDzX+ZtGa/PoUPPnyp0Fe7JcB2tucOocexav2l/aAj8I0orNJDbaipy
rGZdeqYkv0nWfODM9tMustX35tTgSyPdhEFxJXoIhaLQyG/l943dcz9BiZCkfIrA
2DR+K7rA7OtyJovSOrGcGSwP/LUgW4xwSNVT3peFseGFIdwQVSpcDBKhhJKhuwfQ
N52A5JKpGQjlF6pDbyPchQfE07wfEOxjuPr05dM9pwQZn62Sxxq6ipHiHAYbN1v6
AzE9VS2+cxgJThkaX/A9z7nFSK2rVfWHHwjtGy07AYKC+wd0/rCXPfATsQP2NEcm
tsfKl10Hr+YgrRZmQYDYqogbp11/mKlp62dmrqdturHteAySBZlXFEimlDen0227
4ZPyMHS1T6yl2nqJm0/PS0Vk9aEg1kX9RRKisF9m/urOW4j5hsugWikCW2FGie9K
/FIgXIeuEQ+sYdwLfrxUGaoiwcA13C+VfP5zX2PIdM28iBg9Lg6PMwAPlyprF8yu
4PxtTdkxX6okIF1xhvamuShnswL8FCX1/gx7zSS7UVSQVV1HHz3NbghO2rmQ4MzD
j+SMhugyF82NJJXfuMr4g8SJu6McLdTwqv8h8nL5viROsLiZwaS8YH6TBdkvnQkX
ft+j/+n8nxFFayrpQhS+tglwJ2rsZCji9zbYkZQa9pLnBs6hUgU7sXVlLKLkUyoY
kGskGwXJ3L/zIYWcGmldWqN2uTkGrpb52blVoX3CXFGSvzJkGaSqHq6Zool+QUQd
o6uLnzHC3L5gk7Iptu+YLRYElqE/SC6WQO9YopWPLYZf7hNR9Q/Pd8APqlpl6Q1Z
UXjPj2ut33Sj9qhrweMR+YCKMqGskXQyc2bxeaVeZ9CQjC/bn+mRyv7IUsBf9HAV
Ld+Maqv9K8pNfdu/D1gfH3ljMrVVnF09f4hvoISlvHQ5eHqyNoIP859D5RSuyPV9
824tgIQDRfW95jfEm1pce5uAY7AA7fFJNJs1EX1awMxCc3HBZZjgi7BcN0xkSgh8
V92j6wMMRojDqKkRoupOtIpq2KJMkQDNiYH3kLUfXBYOjrBa/5tZx0JoGjiXL+9d
3a+i/Fu2jjIeg5VU6qq4yl2SSyqLBaztyKMDLpksf6LML/poz/Xa8hezWdO+2yAk
9mOjjJO0SGc+BcWgleGvdZHMylnLAyMIQ583hfxvZU5SDLusQWPdjmIRJvYdt+Xd
hjbsfAuyOgqNnZn7UBNiE5IFkx0rP4/PPuH0j2OfmXaYV7d1xPFuiUc/03SdgAly
OWRTS0Lx8JDZdr4UdhFsvEoSA2dBV7vaTgVKegUOdsMC67ZCeZfMhgKq3GSziH9w
qAo/M2j+sbpcM94ybl1OLutOhvIaPNq7N2iDYSY1XHQOPybGto6kXF8V22a/X0HQ
UfxTuRFjHaOUTrVlp+dcbJgDUppwznZ0ECbp+o6f23mTEEGvDfdpPvjY+iSboXvj
NME3j6lFaD4YVMzBeP4kHLJrKeFcv4TgcEoweziWVxxMwbWIaZWwWQUVcYOBJl5g
178fKLcypc6vyIG8yO7Qr1BuplASWXpzu7iccYzogXztoPzjjQb+kDtdb+ENW89i
aj4C1XSoMX/cTCWXlKc1H/EvqzyxsES5cXOk3hB4eXqMe9N/htS4Hmo54BnK4co3
lWe5f+1qgscD1yXhyu1+PISIEgjhvUOxDfmYN+ufUYZMFuTYXGatNwbky+Kt+QHO
p2czobmf1cBnMlkkyo/ZvpHMQw2V+PtSv9ZwRl3erjkPB7u0Kiocehbb33zTtIrV
ckApoAw/ZLW0sKdhHqv0WAV9fuZhojYTBm02hURxiZcr7wHAKJ9DutMNlaFW6ivf
ZqiMFWf669Qze/j6KEIcFVM7I/9Frt5oCQNocoOIhlsewM+O8KYztGdXgAxSn1tf
BmE1ts0OKnUibucQzQg8hh2OP4+dlDg0KdA5xUw6Cu/IR2z/WhTD7t0WakbS72by
qULoaeZyV1mCFMlK0dFsaoasJb6O/919bAa8txUo9s0Kr0C0ZNmX5ouuyEI4mWgG
JiHWlhAqL86g4obJHHyaCrW9DgDWJlpFuUP1Gq/gt/EQCGLSu6sVnxf4UtW6rJDX
R9F1hndBe/Z3N84mKCbXvQ6NQl3NyqLokkzMD6yBKEFGUKPG1G5rFiHrIH0I4T4U
XHioR/Bu4mNmjZ8DM3Fng1L8hsrfFHJX8kLYNY8xFtoRBOoxfQaEHFb3sHY1hvxa
gzwFQJShU+B4deYBuuIbFocgh7PiDlqFCYfsa893OP5KQhVKSQDTRRt3uBQJ1G2J
C+WbGQDfXFe0qOqZYopFb6nYmtLtjNp3JgmCUmsZO9uPl4R3QMqthsDoBgjqZRuQ
SVhYy6tNEKbjtOgHiFTSJ6hswc5+P6RPnEeV1aKMPofwYEudNk/2Eaj0cgewYF4C
3/PxyOQq3h56cy9xs06oTo9SkQQ3ukXBuPdxdk1A/val2DRVHoS1jT6kja96FKGG
ZLl/zWplxEf2T/AwX7o1jnvcUG5a12vyOydbzlHniqwVbcH66fOaiOQzM9hHgTC0
lm57q7gTfzR6KukKnIMU/laiY1TO4jsXFmQEgAL7N5Mzqhbgj/Y4wrFcn/VOkhgE
EZC29RD/Dx+Vls11gN+z5OjHKJ6A8InYN1MB1tgbNqxddmTZva1Jhk4o/+cuWao+
uGeHYnAzVlZ4j13rCeYp62LJ3U2oaLiwbM5YU3KFJztMsWVcmCxKaEL2y64sohOw
rYLw1oq4u7s8wHXj2E3Z+Okeu+y9ecYr660+3z+ylr5xKZb4+/lg/JhkbJnHmM0M
VykD9iZshDhuZtW9qkBXdNZctbJgNwUoxs8PiLXdHyffknTxpJbZC0EuvQQJaJKn
RgktlGhmcMVJGd5JSngTPB0lAKl4Kl8Ryz8+WP103Kztn9gVEQOmITP68lLaERji
xy07w5Wo11q8kdpfTXKm3Ga+o7b/SuvYA5yJeZcZrDWAexkbSIstb0/5+VlgKAaO
193O/XH6Q5CNm17vVtNqBy2pE149dYxzrX0aA3hGBB9mh9Vx4CTeTPAcL87gUzK7
CNK9/fdVlX0dTEBc2NWsluFSd8yXytPMZIQoyxJupMP+TXM4tG1swoHAHsaxpiGv
7hCtTRC5uy1IiBxUSdeyXKK827U9vkvb7vF9y5P/+Hf4V3cFJkT0zyhGpOz52i3z
c9/sNnwHiSLVPWgvccUrogmdfsVitpg3E6GLJUlywNsU0MYp46hDliojMZYQ4/L3
1ANpoJiKD+39vE3iC401WDtRcH4H/6xeeZIo3pYbwk+/7qqzyd03GQFDIaulXLQb
2X37uslettItaEYGTEiuBpRDszloFaCITkLC2jVj+xuog1QNWP73kQvOnJXDmz1D
ZQwbl2n0gUH8fu0cs4sfvq45CuV1JR8tpso81+7iRxDcyvos01Ejj5ZuzsluMrt4
jDzW0m51Wf392maXrTVIqLWJgZpsf3VRs5Ni3kH4XyX4adrBbD0sQFlk/5k8+nJf
h3uLcXCg5l6cZ/bAz6KmLrh9AO3kp2lis2rdAy5geLoGGlnbgr6PQNEiJ+vXR2P6
ykpbDhapqTNcq7fG3H3S8U6/mPQiGcd/+xigaGhZ5X4VN8S+B8BuMtNX+cVe4r6N
ZGkhvDzq2v3SGNjGO7XBSWzfBT7oivNgaA4EinZI94ya3yAgEdfcw2RZ5IoMN6NM
ACKVOjUw1jmBGdfRLrPSPrUk9ivtTjhdnOXLE/0uv3STBB+7dGnA8TKWmV+8TGBY
prYu2LL+owp+pnRXyWd05ij+ATdTBQ6sxYPNP9XRVWr0ogIS+0v/dNv0kFF5qYXm
Q2iLLOrdEtid0Log0CF8GMyhQfm1lI3e8OzJgyGuVfUbqTewJKsV38kJk7mxvOm1
iQ86KWBtHZDlp0DlGkP/m5hXZkDL3FUx0zxx9OVSFB5l6eHnNOSoytpztl9gpMw3
l2M2NJ11ZRnG4rIkAFdhnc/f+5yhTz+yAkHws8CUNIJI7HSfBL9aVDB1ptS9+piP
h5IrrGGIqWNoGhtb9XFv0YXunrpbWsBWxFD8+oEdSR06Y0BAkq08aieYDQ7Wo8P5
xTo8Dfc/7XCA6JGMrc/rM5iHMDCpX+V4IGavWroBfuvyNNrWur8546V6cYmGU2Ab
mhqOW9unimxzvzkmLrt4faIrZ2YhH7XK8V4NtJiYtDR/fhE8N3dIPvocdkI5n5tg
fyyNI7+DQ1Y4dwQl3LN4xtr7SIPLxfbq72V3KRS/3q2SxSkojWTCV3t1TDBQu0vW
ynqT88STDxDOvdvjvADVgGoT3YaXCfHi8GDa0VEYbd8YgGZ7xfUfODubizz9bOOr
26ECkWnkHGhoBjDv4flQT6gMaKBJwWg3htilgrnk+3hFFnXWQvC4xyXwWJuTnbyG
NBD2mu1nQB7Tj6SRwmWrZ6193cBYwp6RWSSyQ5cITytdaDTqXyKPyfAT8wdRN2gm
v2ykzxUXN/4rYFOtFg9DCm1/26noDMT6qWiVrXjq1aR15KEo/T5tiDRGKbHXB6mt
pxCQDzkFpEkvOrwIP4OSlpl9UU9jOh9NvthpApegcMgOQfaNNsHXWFMdKQUXchrW
tTNuyuvJJlpgzfJRwStNBVrsJV1XHIyjcs9FcSln2oY3fTSEpGz0r4GcrG8Cd0eB
weLH3NRr8gFVreLIzKTbeXwYszA6qAihMrlJv0g49py4aiDL+MmBTXiUbhChT8YU
4h1gPEJEC53htOI5HSJw6ctUX9+a1XlK4BlaCH7xkQisE/A30bt5bRKocV3JzxmU
24RsxWCSF8/JRLdCvMIx9/tK93oO/ehil2t5a2ixBL4c/tPBCWFbYC5Pi1PN73uj
fZv7dbuYmuRbBYztPcOnYDladXnoiEU1CHouCYyj15K242tu53B3D+3qexyeN7ye
ozlVeja0OwL13xpl9Fuzeqp6EqN2eqrOPcP3B6Bsfxsq97V4QlocYwH78uJE/PYy
Eb+Xvn7mswkHB61NETVvPIlwWO2rCAF/BWJ3UpB/HgYYxNpteIY4KZqHBHp8L4tZ
kIKd4GwOqHkrWQIRkVrTY930udAHSpY34tmenVbGcn/z9m6tplZkwJ1REmoSA+1k
V5xDJLb4CECZdZ2frpeGn66H2j0hVugr4Wa1ocObXkE4UL+qPAGppAwNMeUepHdO
+qolEMykYa/IOZC5Wdb96XCLTWpmcSCs3+k21gs5QVqwJ63TAdf0r09jfFww1rNK
drum/x9qKDSktd1i2vS3U8a8aLYvxmlox23z1bHkf5BXuPU03nj/h42WYTdfFIqE
yLl1hz7RN0zPSuFyWcALKcWI3rJHlVIVhn2KXWLEflf0lOawgwBQ4tBvZLBGe8/R
gelWwfVYQYSm1qVqQomw7LkwdiPSlBaxgSTlq8efSsGbTqt5bl12ox0kAdVrCxje
7VyoeBCTiSwrnKlDRYQwDXlq39hmJOpriB8aFEYp3ft70mL4Eln/sQkvZrzsUW1b
vj8YpaV12EOp6B87xTJyIJX39fg1Vv5kHAd0LL2Ea5yAZqvQeKaKjM3Gi2vykkVd
UPRYApW5WAKJ3X/xVVnKIWyZYTo4LuXlVCx6Bbh5dsDsOuYx6WLnosMwaA8YJ3Gg
WaCSgSz1kHGqm4CNmNDaxBr7+T+iGp1EhLx1BWVQdStHOvhmqrBCqdZu363HXBh+
SYNOq2vZDu6GiUbeQGbZ41SOF0oQFhfFq3YgxtBfTFU7UKMXVuL/CPHcfoNoWPYv
IoUX2dm0/fOWkQQ8OAMmwimoe+GoxMzCYeBi33Yxrfk2Kg4XQ2VF5ChL/HF3L5Qd
VkQQu2Icofw6rdreC7c/O9gGid9AwCoZXil/1QbeQp3iB4s0+cD+CWV+0buwHpta
7Pw/J1YJyUIgQicpHS82amcOrSt4Xa35q4ptTzxDLNaHLrwnxWHp/29UseRPZ4Eq
Flpn6XQTx+x7VhLvQnFvSGOYPPdqVrMh/NAR4CQTDd3M+/OAG4bZwH18Ikjk6YIO
qB9PIs8862BJyY0aAD0zGivyVxu+fMqrZOrZUdbOOVPTrvKa/veQ30b30KJojWWd
3BJ/QKns0P/SF46i63n9HMnAMpYNYm4ohGtrZTuUDu+GBEJkM29ApuGQFoCLIsD3
P4zwwBm6jrodLNLo3cTSPA/IpjCS8hMHAjsMMz30ajWNNIIOq8mIRHQBItVmU2xM
Kr4R9W3pHXMlXxRPAgJnk0R5O2bUjTn4mzbKIINC8LStALlVlNgQaT9h7JGEW3xf
sCUj4KFdb/N2s5tE405uyMTR5ku29lCp+Tfo/U2JxirJ7vPF8QFBRPTReBEQQ868
tfOvjuxQvGCbzrWD2Ja/XT5uBawZ98EJUzb/Am/vB7pTy0EFwKKtvc/oKZLBCzxq
i2oZCxuBhoTD0yxBHSAvzQEA2K3DohEcFURfKCKXkLfoXakAIcOANobKoRZsYDeo
YDxnFJXVexuZ0FmbhAqoRpBzGODYw9qRnHpAsA1i6cEbWud1puoFTaek7bH+ikhl
LN91rQEJadJoVl/Bk6nZm6KF8qHUd1Snr5E798R55rhYVUxL0POx083fm+xLPiYC
pHJfHai1+LYuhHsIjINvP59Mflno186VIYQKE5bVnLOrGX0G2BUzvkntSPAdqMr1
cEob96UVUIPHCSKgYGFx/JVFzwtwpez6b3/d9OAL7WUOu+JwAsYbgXaEYtcZvuPH
utQymmAvLC/0+Yc2m7ZPvwRr7jyw/uEx0n1IpKCaScHcaj68QlfxtHMCdEq2ThP0
FmZ/b2iBeTeaQzpcTyJ5w0T5oJ4dLWyxgoyRY63NO8KgHfWG2it6TYjTmRuWVH91
uIWuHMI7xyXVzMuhVPXt4ABNMkh8fNi6HcCHaBaU4saw7eo59C2fvUgT2A9BfHUT
Vbbli9xnpvxe0JT9Nez7dg/76ScSY1mPxYr/mxRHG0dp5zdZo9xftB1qFU3+cC3m
JxG13SQdr1kS52xcd1H/ekRkCwejEL/dW0QoeJ7YeCuDqnOAByf2YjXSB3/ImUoE
AHnQBO5LDoih9hXk2m1SokZSJH25yDZ3X4hwl41Ud7Wy6pbwhu7uqVihCMu3R5Tw
WOZ4xqI9iYaMFB6jCxVpF+FKMXvk16jH00R4CooMNLuvr6L8VpDnONtOf8wuavzP
2B9vtQa+wbGw7Q9UwW1EvbpMpYjW//5UGN9t12Ili+V6StCtgPKZGf5bj6VXCmQS
BmQZddOKFtmDT53Bx6NWPFbP2X5Dkb+V8bUXDQ9/h2QbWSyyNi9YY2oNj40q2zJ4
A2Tm7ZOOfuFEkxebjJ9MzeW+G43sej0PN7L1el5xEgo5Hg/AAsib4K4CvpBKUCr8
KObTnFpQkHTQQL2zDof1vTJYJ2dbFFG8niG70QoU/rPC57+Y62XxDfvjeyA7sZnZ
nCeL1NP2dVbKW2SSmio8nA53R2KzlT8UeeLTYbiiwQyA6ZHDv231nvLzMACl9yHz
rTVT0EceSerbir9edP//493C0uJXd++VUJSllpXyC0PYFo0/+61KZB0qHgtFXLzd
FupJrjQbwaHeLdKKKYcxv0Td8oGDWN/dhsDQlFp5vii/5Iv0WwU/sdCDcdl8Io9d
ATUaV7TuJQAsbWdjfYwv2r37+sAdhhgfFDSBAgbL3lzyIO96YGxgKl7Phk2fDD9E
EltiJyb4rhJtU/D5/V8aV+Mm+TXMaPllPGxUWk07FwGwNs9y7ZJWhfO2poQgEe3G
npcsNqM+L94Lc0aMznDq3VSzLYJPQ8OJq9XxDDVjMrUXOgT/TdZ7Nf2MR4GFZqiM
e7yj3GX/TDXnZpWwqdg6BbGxVbkG3bRm8MZaxS7xByuaquNTTorlI5ELnBvqrS+X
PureOASJebVYSAi3dciQHZQDNwge1yrB8wezXPadO76wBuAXOeD8KFC1L5axggX5
Dd1foKnDmg1yhGzfpZ1/bNvfheeYK3ICvXBNbDb4VxURAiXQmgEvJCQ+ZVtFHWjo
GmEKfRtYmzxVeopqBUJD/uPLMRRLlPLUpUtWX9A0C+y9KrEIbEiFdLq2lYUWJf5F
Kf+MXP8OvKQlGK/WIfBbRIcKFOamh1EcNTuNqNKEoII7DFvVdBhkCXuKUD/mbgzz
nUxeD1HPTmxCAEQXj0w+Z1tp3WGT1aYiDWb1We/jecp533k1ehaAcDgbp/4fO1v+
VGzIIJoPsdeKuBtUCdHHpEklcfEWSHiMkvule8sYrJ5ZBgBHHHogm/CgEQGksmr8
8C9/AhU117myiOel497IqGTUQfE+WvHQzBRsAPBWQAsEm5/S9bi8AudtYly4cLRC
R6OWlNpQgqokQSCb2ixOPAJZmHvfmpeybvbmBbNL9Mz4RAq3hJrD1FbBnpVePrKN
uGAJPOmMjE7T4HlC4K+tKQNlRdZMcoD9QOoI+HvWLeTM7sYdIEWluuioQj9DrQmI
GGP+I82aFAsbs9zoLeLmBSRiYtSZUvQI2EvnONi5JS6tMJICoUnAoKEaGy0V+HOH
yxdKmKasFg6fzMG0NYHQNh4Yw7eAldLE6aLXh4davlE72C5Gm9j9qkwZO56z8UBZ
IugEiTV+IryzhpdGbcZ4d9ZPuUfUAuGak+A3l3cLODNuZOqvQxCzxPMAl5R221Fh
pXqQg2MOGDuaSt9wJJbhU3iTi5/8N4bkjzmBM4ApTsby+oHsgzHBfj+zeKgglF/b
pCDI0MCDSpTH1CZ2O7fV2yq+6dCJQqogVgz7nzJ7UnEzBU6GKl8OtTJ3Em6VS7/f
Sv7kShsfaU0xzpqYVB1NWaTKaQRHa502VD/mTnmRv9dz3rYOvHTbD1d1SvTL4s6I
LiVBqg+opD5UT2mqeeVzj+fCzMxVxzSb2uRW4feMYth2yQGIGZGK9fvB2nu9YpQQ
NgA3paxuAuVn8Pf+tjL+WMhzHyMw8Nf0rsO3Ac82TqLYzYadc3+LViE3Ql+15PKg
99GXybkhVWDQJcJOxNWZwt9ZsstfzMRiimTlPXCH59uwlvZg48sPb1Rtkd4+eF8S
A74MXMF3zKAafe1hAv4RNrQmFt6GHDyBA+6CyRAWdTzWWnjiF0ZeJ5xs4zMYYX6R
/m85ivX2QmiwLhckvNmFZVHMUb/FBb1FgwIgW3N6REsRCDoqqyECUI3nHa+LvOsf
fQVcQxTSdOz0D3Ygkj9lVEU2u2A4B0ItOsAmwkPpyLMCQS96dZEE96KGGFZbBp/p
+Aj6Qpe7gfPl/tO2cOpAIf38BKD8i8mvFFw2EKmYi+Mk9QAi/DPgzhPXtmiRvIWf
t4MHluv8rkWc0MOIHSR6kcsIcbVz2VPVMSVpGHsR8SgYmWHtq33RU9vD4xCFUzNW
FX6EFrkjvMoshyaEfZxxvjdbNLAMEwNA3t+2CQBZvjhZer/RuLuIhLsSsMOKFR/r
G//5UFg+t2Tvyp/qUaliSEkN+xbBCWOQWS9yxhK56nB7uERUVo3FucK6eXeT9Q9g
LGWq332+MdjA3JBKdNcVXYUaoqcCIQpKHgYsFOuxEuuDhoUmv/t6Rl7fekikA5PD
bDLOYvaFG+RCTQmE0QBcLS/t87yqytYl2/H3I9z1J7ykwUsUChSGw6jjUPDW0lq2
MjiG0B1tcDlgtw8ppLRxPw3ARiLIeJyspcGCjVn03BUzEiyav1d97EYqAQZc8iAw
61YgjIudIn1w1XYi+MwV+nbEyB+j02H5MyBvgMssYCf+YHCEL55fZow76MRR/BuS
bmWGMMZgdcwwpfbikJ6NcjfRHYlsSqrJaoMF+8chf4XN4aHgdCL4na2OEaOXl8Yi
YCw3XFAGHiJHEffn055CQoEmZ21RG6vCXCH1ZWhY12ISJjbtRPeSEgTAx0A8l0Lx
N6CTC4IQApA239i9XZOqZHOMAGIsVJKZcfruci76WgKJDNwHBXY3dHW0q1beVwc9
bXujLMeGAPsrwOEn04exvuWtEk1Gu5Fs7sX24DDyzSGDJ8MB21xGuIqBX3fEQfKl
0fivmTsSPTd3A9VLzSxiy99KM3gPWqr6xSN228eJTkM/vpK3UzaEVEyWk49H8EAl
/O+y5Tex2bFVzSE7v/mwn5dzkZiO8cz6IJO/sKbC08CrQLvCDhkDh5VX0hjSv3CV
/gZgyRMWH+dRO3E7CZJI/WkNGzcTMuBbrjAskN+rmtdLL/buZEJABSQIYcm+2Emp
fV9wvo20Ge5+GvAiPq87wCITJCWMRhSi0GmD7on4z+9PiehmZgA3RU6REQQVizXA
fKiDCQqkhSAGTAXNfZsJkj3BVcX+ui3y5kgv/gGnEYVBbv+mzdCKMeR3a050m9Or
q7FoUcrbskgBbUTx/68GZTLqsKuIJRDmE+G2I/VdiKmQs8a0hoHvX3bQuCiwk/2F
kJ6ATnoxy4wRDuvV4WWm9F9Ja+I5STzR2ThB+GFu2bDU658Z0N46fg9jqMyMqKRN
OISq9v4201SzRaQDBEsfIKCKLoLTrkTgNxlQJKODsTx3926Zw0tt7iJzOdJUdzdy
3lSji03cqB3+WkOvm1gixrGLm9osz36il1DnrpkDSv2YJ3fFesiAjqZ0CNXMAzht
8cyRFGvkdVn3zrVh9CNmsC4QANMEBm9HFk+lJYfTQo5XNOTG+r6d4bE+YiBE2ac7
u/dszktIce/ZAEMWOCCgYckQEphrDCrZeM5zilq3G6Dn5W55kFF4TjqZ3HVGT6qO
RfeyvSRWudVWpnoip4isLHu7BmPIGmhYNh1WqZNuFn1OotL157YWW+j5YdQcu3kp
hkU3J+TctUY0/5/83Iz1nPFNVsHADl5vafVTb61j89n0N3QYWAwJ3tqnEYpiYelA
7aNjKiF6z7Kfo8aFeHkYjIQ/VXWeM7S766PJ7xc5Ko5SiFxvHX/cNjbYkeT99S9D
i4Ve03nS6sUo1my+LALAiHIoHuLEwJrRBKeIlLtVz3if+kIYkBVgzKCiQLGnEiJ9
XQBcXMUb12ZAxk8qq4DJarUaCXWk932mbtm2hVbGyHipPCLGpovJ8EtmNH0HILRI
8vAIdcwE6MU6Ek4IYaJM8T1ciyucMS20PavwKCbch807Y3eqDJqdQqYtP5L/AHY4
6Xxzl6S6wmo8q+UcbALlY9ZPMPl7sFOH5OZbCoiNjoPA3RCfPNTZUxGbuQn9Oy0d
O+d6XxTfUV0eVoc02cE9FQkFbcAlt0iF29v86POtLcRLmXmt3Ko5aBtlJNA2paWt
BArmqqXOihxHlEUKbl/A0xZPaRb0o6OMWeANoq+gThR/GVQLVsTnrCNgMsbFcXxP
WmNtmiOLUrsyZzNoHRAFOyjocx97Zn1MFE/8lQbsBlaYTZIeRXxqWJ5BUb+5c5ga
5iIEy3Kgnc4bg6PYBvnsJQIojbar/5rP8gLs0k3Kud7vMXodvWgTQXh6si28NB5F
jVcr9slay9haCNIWBaAeeA8YXa+rBtUuj+ojgQBd8drWJS4+bcW1lY3mWxFZkgRu
600QRKeefOxcyhaB2sv3nF9t+swG37JVaN3NUG56EAfIRazrV13YzSUkzr2rVKLD
3ri9bCDDbjrmW39yPpBoW2WNMGqfBNmg6kaI7qEL3z01vjC+pgcqIKGlE+jvomPV
stRyUZzr2RamBj8zgXJa8FXgBFwcZupBVbsh8yYXQwq/EFy/MSM7Ikhe3W58VNYG
0XZkpXzAisFL6OpbxyEE8pw2pMF6y0DEkSehV4P3dlG43gERzqDo1x/mHKlz8I3U
CLvkksv5ZgwEiCvY1dq0QwLbnEVIEGJUPROAsLp8t7fxCvLjaZL+dNW6ZYj722ma
6cxh8ZdfdXnG7SK4uEj5D/a6KtneAggWVGjxJiIXRjNcy3YGH5fE9sJ3xFVs8G9t
eASKhgJ5QgCpzwjY8g4XQqL8+thF+4WA0QP1MBP37y5hPDqR0O1wf8UdOcv09/1F
KcGnQVvjpna2e6LpVMV7MPQqfCJCa3eK39YuLyGod1g2mOwczidKya4KTdWbvhn3
qxmsK3rTW0SrrtVsBeTCPfFEuWinlY1nDVfq+lFwZJidjtFitYNNbSUB7w5Xjs+F
UHZmpqu/6hwwB/kknWjCSeqNnZlMXkb8b1t7N1TXRD2lfctqWgCo1HXKxTxC8xdl
BRAQ0uSFv07LN3K7AmMJwVFvuuuT7U35WtpNsB3PI4x4DvQFt55YFfw9b5X1/yVQ
t3tDxkSov1+L14TmSXJTnHkEw1NJCf+tQnVlTvopdTsAVk7dNe5CZDJKEedE2fhT
XrhCLcS+xRcvWpGGFMn0vK/FiULg3uco8JxSHvSnajK6SSSmfJXRXqfi95DeoCEF
fmNtbSwo1JxMYdkrcoscr+NKDT7hzayKM9VcAuq2FXK6Co3qu+2JkpRD0wukBZ5l
NCvXggUH89dRJKEzvRltSAYLwf9n3g9FnwkqSlVZqZo2rmtDsHpKQXsisHzA5OOW
nWnVgNbefclmsoFYOdYQcSnLEbRwlH14i0spGzwni1UxKVTXDujL5zTlnGedbGNR
PECDSoY8i3AgFq2cdSENGVUF4+tq64rrhxxsumNsg1CyK/RylhN6VJwhu2aIDtGS
giugKsdYO2B9HUFF9HiBtwpXHBCUVYN0HeBp5dH+PbNyjJ8BtIR1/uINzNzr+DCN
OHJwSYog/ibiQn6RPgpG+xW/F+fxe7CfUdsMkLWL6/AdssJR+3PT69I4AD6dgdZi
olWkCdcaCNC0nlDwej15RdNxIQNG/cvhqdNwjgSrWHy0WzTmikPOEl+SIiXCom7/
Dcssd7rFWoptEiUfXfPj9trWXqJB5l5VBNigPDP/DoXasbDfi53GExCDNuAgxDMK
Vz2CS1oX7ehxK8frEkHYZ/o/JFqeHwilS7wbVdE9D6sIydsBnHO+WDXuBFDkV3Zh
efByPdKrGdawqVi8V4CeGWitdkarVhQ0m9Phj4jaHJfW0aiBBVfuSlvP3A3OXZVn
10hs2Yhu83g5dNpBGNtd5+2cjjc1mUaOCcVz33k2UISukY7n9J8bIHJs7fCFIJEy
KuC124PSYEGumiLnweakk/klVZFDIZcgpTfzhYd3xNQu7BijEcIzJIE50f97lNDM
7PKjaY3XSnV1KlvSN4z6TNcuoAIRNL/gCfEAYGKf+FVnDoFuFzJjGzu7OOEh3Hd1
SDoi9NMpWyuLEnqKiD1YzFpU4N2qnyjRYtZ4BdAwK7HgQenHe4paAc4byPhACHZ/
chRhggdm6AmuFZQNS5lpnXTVdSecKKkn8pat63N30RDm2xqhSO6jmZ4dgZZg2Sng
ppuCScTGFRmwszq97r1LlH7ATji0/3HIYc28hcbe6P0yvVY8SWR75khBs6L9lcdQ
Q1jhjO6Qh0qrG7P83EEaCXlNRMx8Mfaa0abnb+qdsuCrbiGVfbvdav5w5UqPvpTm
207QLJh3rBF6QRWf6/Eyt0lMCWCLvdfx+tEDHYFwx06Q3C6TsWfk2lKNEaJ7i1wc
H6A0LvKx+2iE9XrNQp4ri4wkPdnwVft/OroC0t97jORH/ZuE+npC72IHy9R1NDyr
SKfqZ8WIRLHNmonpk+f9x7yoAFGZhdVHuBU6C8uOollDEk6Th/tlDpk3c+NTZ9oh
sOeby8e4hGABTajh9UHTidZvNuCLCW2UEG73XZvvElxdsFPs6EulWSANeqAl4Xqq
KoGhVzXhH38lU9wNr2KqSw7PcA7q/UB4wK3lX55pUF5Eev87NKkyKVpGoVhjxUUP
DRXnuHqm31HOMLG99z+pT4xzA1P3WkQ+bAWEdl2nJW+9yYpOIQUPcMm6DWScrKNR
9QDSAPIjJDlyG3+0H2mhLsnsdBkVjOKld/2GrCBM9Qay39M+x6uUscr+B/Gx91ir
iEOBTguM1klY2XiEaokQt6ZQ9XHgxzE5vfDykBHl+uRRg/ogsG4aLv3+ZrYIxGKi
sVrPFOwiEHZTZK3SYI0XWhKHPmLF/fkS8Oi/GjjgQOj5oxMHNCwTsNZYaRvQ06jk
yVxFd6552TiIdOBfN2w9xM8uQHnZX95BB+a4xv/w25Am794HE2yDUP7+1eTZGNZR
/LBF1i1wPN7Wu/b77T18tXvAFDJqHP2JEwP+kOIlAmMEzBaKsc0WEw1Utl07XNJg
O6NhtCjw2sZeB8H5i0JhpT39VNwFwBhFah3nwn5i9lSo3V6fFIeG6UfYyg6RHdLw
t6VKISLLYcV8XwktRELWr26PErGuk+iYjwV8zmDiTBSqM9qStcXBFnYqmNnuWGcF
/Qe/Mzu503uRxEkxn2xjus4UZwmVj64Z1y5tvhq7OSafo8E/eiGII/lceLGZt0nP
1L8MHa7WvZb2n5hxJb3j7F0KseglW90lYZrZTuJiei8fznVb7j0hOLmBjg/hi4wC
OgCqUmEYPe5XA9OhvFGCryK8OKpcfKwyLMrI8wtwEuPOAJm6O/dMCIrrbXUQvt7w
yml8TPF/pvs9dHYUQF2Q7wz5xayFg2PpqxnO6EmAQYujziHQljNtbpJBurzyEaNZ
0f9swpIhfWvIBQZbCAcFVuP90unJECjypXvZP4x4Jo9zl1Tl+qpI+SRw3ehjPTV6
QRagimnZUIpgheLmO+z3bXuEMdEVgzJWJTxTKrQdYkn2vU8e4GIj1y40bzX/aBx0
ZWFFBED7p8o5uaaVkBFvPPKdaaMOkyaBh/kDcTTiVWMcoQVRhkeha7KdW+HF9eh+
cnnySPBdp7PPX5QgzNwV4Xc8A9MNEIF07LfSI4rA9EWf0/qlazJcEgYW0mZ0Oq4M
WSNZr9n1cR5NXlciLccp69nlJ4waeK5WhP7oaZEvEQpJ7kPpp0JZVJAfoXoPTbse
W/s5NQ7m7bHDVCFOa4Dsusk+8ywvaKJwKSAMSpFLTxChhlqZS6JW2k5TylxmIyCN
vlrURCoYxqfcdhH8QyYrmiNpQ9Y0ML8zWFSLWOGh2QDrfETDCiiQDC/bHSFJCa/Y
8f4OXalJi6ck3OlI6jLPFc42TLUnVM1a2nbicPrTdIkQIpOTxZ5H1ch192wZ82ky
/Yn1lqUFnQFKUI7SdIoaTQPwmRFxKjEiZOYpquHWI9AWsUSjrvOBeqjVRC+KwCZW
V1sNlPXKn65I6YqDUygXoggIUk2f0h1eMVjXEjUT5YrqzCOx54LNmSxK1W+W5OMn
qbkO0CRFHzPO+WVPMbLw1rZbQfkWdR4PfmuZqyX8Fr7ZUs2lQ/7Mlb3Dv4v++XBx
cnL7FHi6rxcA/yvnTwHIT4T/dCo9gOTaeYZMBmVQ5fjMIqNUpL7SNzpfqe4xLjtS
PR5htxStH+onxgcJkKIZNu8npxindPdCWvEnVpyimDt6EViVqHRxdLBNN2C+4q/p
B+r0t56eAVpjXQmYpvvei/KOfFKIGqea3Ron01h34BgrVaIVuV6tEr3ygs0VmATt
GHLzGh1H+ZMBZLTmcxSXBYcUz9rgR7FKnogSwoekiN904pMbPQFMS15y9feNvszP
APKzy8eeziSiKXvlRwDJeByGf5f3MR9Ou6s7LVcxM0Qz2QLLr0wyUm8Wxhk8VKZ8
jb4hWmzIphq0mI8Gi6OF5lWt/NcQ5GeH/sIqMuKnrGttb+pwOAMpc4w9fmADJKw2
RZ82QdxYtbNCdtuhayOYdRGNfBUUHSJ9DYezckPDVDu12orQqtWyJmQNrdJFUnX0
awRtrrNbfJZ8C+WhkFeZiI9aobijavtZ3Dbds1wxzWHUWHU3MGe4XiLqWCZHut53
FSBqrR7XeT2HBlDqXdcXv9afw5qVmy7rEaIMAjkdpTfshyISgzMXi4J2t66yHEI8
1xPZ1X3Q2WGdMpKF/I+hBxYaIFBlhREh5lB8dZtlEI+h0BQ/AUKO3FFl89mjYdib
0AcY9fAHz13L9A36sAz3V1Z0mZMb3w+RZObILZzlnaUg9QPB7Gbut/j0isN5yNO5
YPCTAigziWoBLzkXdcMLXpQ5/K8lOIHL2P/jmb+hMVUahvbLWhEWwdAQs9eQWAyd
lWfuv6Nd2+MZ4XY+oYk0CkjK8JFGORlXa2bVQVqmCEM1vm61X9JGlrSsX/S5AcHs
fxo7B+ZvfOidFvwJwNdGWmzH3O+rNOyVmuhaRCq2GDbn2G9U2bJyaw6xm6rUFHvz
WwRvz5bts4dmVD8Etseb1R2Smn8kcwt49vmEkUdfSspv6Yi6Wl5hZiWRO9LY+xWx
eOJMh2aTCrGOw4KBorf8Dspvx4YGqD7bhuZqmbn1zXUYmNNz1/lQy+d+eLvVz1iN
9jJQQhufL3DJVvBhaHAtInCw8qMGH+7ctTmRxUgsFX2m6aukEZMJTVYlRJr/U5Vh
d2ktATHOCbNkK3HzZsn0HoTsaiKPN9jjDyXg8Uj3yxO0+J4qxsesVJIakTK7tLY8
rEHaeST4DbLFeRTO2M4ruNufAnoiXQ0yByEstlzSIreEViQtx/0vs6Ef1XYntrU3
slBu7k2Cp974DLOiPtAQWVjxFbqwgfjC6hYHMXBmYzAiQMREO2yjIsEkKA2tqdub
3Nh0/IsNOM/fKFFlOrdWPGF3ASsiWZ7qzT+Fbz0TsV5bsW4U6VI9LFNg2ZZ4cMvv
Ykm3A2Km8AbgNXNyxdgcKl+gBCfN88YAQ2uDxk2j3iOoY9FkyTdyls44cwcf7SMX
eKeZVsGtBsQ11phgqugdmIzY33mEo0/ypoY5pVT88hXC+hKS+Ihkko4QmiPSxzKC
vppPKm2hApGjCivjWk1mp2JRD6BdYMevY2mCJOpMSyeblqm8831V4zKybMxitFeI
4BtwS1EXlCd9UYfZeePC/48/eJNgvNDRtUHF6gyXj7Ep9Y6oZgkY/BlbvCVL3N86
J486+VKFp3oIyOOvKcoZotylplwIJ6miIbixELcEqBbBy7qBYSvrV+/bqGuv24pb
kZHGYkcRcYIkzLwAXbLsaPEchcIy0eGHg2BjoTHX3sKdj0YToarTXp5jGV+ttQbp
3qn/kTcjaWWlVVtTwyUb/owSoNnSKaoUBHtIj7SkouvWWYwphlTJPvpt+YU0AxV1
G+odsaPugHsJLkQvtfgup9o9Y0Q53PUDpsN4bvzDjltq4DTykVsSRo5WJUO2AdAp
QW4t0Axk9pwBKWdxLriFaD2wrwQZY8DZDlQcBiVJgg6mA1WJ1ScTVA1kIglqLIcF
x6ILc3fjws2baClbisLDcKCj4Cu4HZ6NNgEsjE+9LrRKw2OTgbXrUkBUHNmJk5pU
DGYKDXVrQ34fi63e/J46ckGwEdZurBvBTbP1GHKaPPE+02/aXShKGyPGGLABWID8
MVRfHnHkAK6ziP5vD5aiWTyC+PZxY2YO/Co47m+v0/alfbpws/KCIVChWw2AnxUZ
HIxKH8roH/k82i7LKZzDvL7Xs/4TBD9lIn9aNkf3EDbpCr4ZmfLigN8WwyDseND+
CkWyaz/ixcaeb6NW0dUWpjUv/MG0Vm4Sh32BwvAVW8O1TA+rXl6tGOD5sx4y1g9P
qiGRqT9Apy5mDZIVVHo0X/TgAVCiIHegzaEBBoOvjMiKfP+6NAZFLU2N+fz6tg51
TfEocdX/sBfSUMEAYVgdxzgULaU35xX8pnWCdW34erdVC8KSVxv2nBn6F1BXpaCB
Ck1IvtjZlnArsY2uZ8K6j0NrOUkJSuhhMT3TF6oszZ0QpdNO/nXuqtJfr5LOtVgD
6H8b7QIFnow7iV2OHeXrEceaAFWl7PRnU+qmZYfNkTOweBnVEeP9L8JKvei7yE1O
qjMoTSlTCuo9S9+jhInu4efpxiZvwKIf23KKyRVVI1m2P4jkkErz8JsQKZqXEP9t
DWxxoiC5ugF9yOTnxaROjn/7e2ztviDcAh8OAHF+ourCO82DtTwMQWRNaB6juXKT
QPPNKhnKRZ8tTWykd3BwbpAMUpaXhiDpMuq4xfneMN8599/aI6ILsxidwi9Qk6IH
ZpgRZTg7bLPFBd+OxY+OVK6Lmzg7vO9K3Zc+1SSPMEbdirNj9yYvcAslgHe9PKBZ
c7c0fe3DFu6bDR0NQgRjFQSxtuoSkxsM08XlJ97ymiIPyCJG8x4jTQuY30e1voKo
6gJDhKXeTtHPgoK5m4JqvDB/EIyjmElBfIO9wJ7O7u2UMZ3eB/2hrHeKBUCY90Mu
jC30G2h+7R6BvnDcYTMF6ecYjTz5wQoc/V5sM75IHv6oPTmJhoEsezcNS7RBF4Dx
OvsqjcAdgZfWeSo+0GcyNRvxK6x910itGQ7CwfvXzWmsOt9TrCfwn774hTOOb/I0
gHg/qVXVR/ktu7bNsjkD0w7mLFqKeWFuTDtSQGkowmzm0E0Ba3GrNVnUlGwCIiRI
ikB/PCrSZXms3+Cj8aSIJoXMrMGuNEiGIm203VPGlzQf1kYGur2CSQCblxENYzJy
jB421QEv7aFvEmEuAczRSwnxUnWFz6g3DcAWOyx+gFOcJz2p0wxVlycoir7+0NhU
rfw5RkfyMDWfLlWDdNgltnGdCH6J861m/XyiUgzv8UNvRQsj8ghJed46H35ayE0A
C/hpUR4zIRCfS1g5SuQk2+ZrLauFjijWieqo48l6QxK8gEPDA03MywziPYL8BDVt
1nhLDuKYnxCFJpEmliYFmMdujZ8XgDCa7zwq2RNibi1ZGcnAuaJShstzOb4cqMXG
r45R9Zd+88Mtbx04oDh3mM1xhaoEnC1eIgpTRf/OAYn3MghqzbZDAClHlXbNyHKH
A9/9wCyDoUXazQT27/1axDLh4uUn4FHR8E7z/DWK/65cto4gWDJVmzHxJaRl4vFK
/mRktdi+fMlfS/+EzPUtYzOeEuONvRppBwpNC6fC2IgR9bhGdRTCqflS8uslOqo3
b+m99zgNJn3qnrqTOGTgUVZ/x/bOFRNrj79okXXYTvSw+XmaMqiqOPftZQcpEKb0
K76UOFuUtOziDFxZTeK9H/6PIi8IHIX3AmLLymz9lLmHRjqAGoYfsKKEnx+BBmcP
Np6xUl09ZImfHaoZE5o/BgxKiRpyIdk9x7TxJ2VDdWxtZR78jh+Zk950ZKUDJ9Rb
KxueIsiiyj0CIznJochY/UzvQjyGPqGObi06YMHM1nRcJxMZ+XeiGZ2GCVLmE3BC
2cwUKR9/jkRUeYaj7O5AclnXnQGLsnARtO18fjn9jO+OCHRadD1Z1T1/yri0udrC
MQwjbvHYrWBeikn741qYbdhUjGJ9Flv8h9QZxh0scm456FUvCimGg2hAZx8iDBe5
0KwPSXlwef8ctjE1P1Fxw98eKTda5FkMXUd2cINIY16tOtpthIvf6CeRhrjT/4DE
xq+UhTqsKvWWYrrDByC7tiwU71to8Qd/ObOEZihSDiVeG8nyonkGu3yD04VeXuBR
7xa7Dk13C98ENuxnl9UG5BSAZJWXkwVAIcRBeRnuJUtcd9qRfaLdLk1Z5Hn75T5e
7DQsJMtP9zAcfce0fZeYmhVu4cT7kJjszg6MayRX/PfOaOzXyuW68LR4kLS9/s2b
Q9b/sT3i9fGUp+gLYaiCclhd9ukzskzpkJZDWRbBSK5ajEsxE5O2JSIx/cDzT92z
0QBHZ+po7s8IYnVlvmwIsn9I7qJ8vkbQ4sdsz4AZ1kgHFYBtzVH17q383WF8jl92
EbqV2YbFI/ZtJ3D4quegpwvyBvG6imTKCB/Uh90dMLdzjzU0ASWvExEULVRKhsGR
IGkL9KO5CmOZR3iQPae/ZB94EUZAb08BqglcYV0SgmKTPlFh5FciCc3yBT/Pim8S
GfFW+glTa0cbmpJcTm5u1j+u6NZj6Wj9RSNbiy7YCZA1aeUdD/pm82Rtm6DjU+3y
VsKpHGIdS10s6VGnl0g+H2rgjNNYSXsXPnjgXqNVTCg7sOrH03h1GWTIk+NgUo43
8DqBRHFRFAfJ6rgFn34jyXEYaWgILHTGHkN+rqDf5BSpmccpk58Y/Emdk+CJHqP3
vV7fulZsRcMb/tz9efncarsgGsl7hCPMTrDrditLwuGMT6B5OcToTx8icGPBjvFi
LCHkwLFLzO1is10ETi/O9NrXJN43VAsyAcsuKsyE6GsuCf/o/5m8Ax7WVvqIVbhA
q/lGDKSCwW29JA2ihu0UKCXJNei+bSoWdphSgRIfdX3ShUXPPWr3PRMFPVcyqIpl
zdHoK+al+UYlIi9h5yVTDD2iaiu7k/H7jiEjA6sb0sJYmKQQjIpbduGK6H3AAFMx
4k7vlrZX+PMotPw/m+IIaqhhmDejur8p6gx6Xhb6zWc1aSTbleiw2p/2Z3Y9+ga0
kHUJPJXawXIb25c/owEJh+Fn+pHsA3ZN8SENljAbYRGue7LZxy+Dln7TLNHrGmw1
82oqVYqWvZg4oosh6cSNOsrj8SFFIZJ8M2rrzJcg1zvUdfsAS2Gnr1pCfN++1B5b
O1XolGqFX4e7xktjTaJFUyP1v9JlzPrzW8mGWNBGDCqahbCnSu/cpR1A1a8LOpbN
QXbS4zC7//b/1MEk1h6ZFNqXqYQ29D80i2Y2ltildjRX8TSjCHFixHSmb52ZZvlm
XuxTvfkeLhzs3IQgVEw9ZsodZi8zW8FuLSFpJGYr3WW99TfBxjAHGxgBEUD9blPL
taHXzB1MJXUnKvVGjn+/cmdff9/M2kSAoVGWc8s+01C8TXAEMhWVP/cfVycRwXer
cHFhQ5dx2dH9dChM1/d0/8aJY1UehyQGC6naCtCDkOBJtXt0eV0yB6dEBj6kGb9y
IoqEdHVJQnBRmRKvSsIYdJf9Y+uKSYVV9JaQm7hksMZjWkZfdFv0Vd13ML812ZoN
qfXTvcmUTcL74Y2RBFXgHFEOthfZFVrMcG0rNkoS4C9Mz2yPXpefz+6yWAhb/aWn
+BR3HlWojU4hzLPWJt5bWPe23WRNPVYF1UYQ/X+M13M0x+LkDD4ugjIxMx5lfHGn
gWyYpWNjXrOQ9pSwhchYXoilgm8HkThFdbV7GT2YaaVV3l3V+P26CJZTr2G/hWy1
MU/1oIysm98gbeVpdwWB/Bi/DttOyfVWFMsRjredboFaucKyHKRgVD/IlJ+f0x/F
7NkHYh3BiW8J9PTkDycrcSaJst9KK5M3evki+uLXWicQMu/STxdxL4LbmLfwAWXF
UBejUfeIR6wfCck3JU9sBVKaaHmDfj9fjI09Jjgliy/dfjxQAB0ijp602WUbAXc5
SbUidXa+QEtoWUcjtM2RBKnrHQBeytKGNo8c1QE8huoV3m0PMgSAF8ZH+d5EwQ8q
sPU6BU4r0kAPVNnYdRRYLjA7/LlcCTPqGKJIfqw6hOlOfBe1ijL/rkO3S3GWtOrO
MVm7Xbf/NGvnqnMf6Hglut8cCy7Bcg1eadGT3ine48gSghR9LW0VabarhBEVKRTK
DhUMM5UNKTcW7LaEYaOy6teRJxZGm4l7kjv4AbDuf+s3Mus4nGgxDH9gYuiroKlA
G2oxGUX4cfRd5/4yrSYg5PeU31v9cdVB+g997O835KRmYxmNaFYrvLxqNKyQcYAJ
M4CqC7Wu91YlA0Mb/063moGh7KZRcUHy8Ir3ZW23jZuwaOvWepxZSVkDbbgEVvnT
m6PyREPVEPAx6Tk6fRH8p6WBjOgdnCWJRP6a3gOElxDL+MntwxNYwjh5Wdr2pmN9
BQ7nv4vZcRPGx5T111MmVAFnNnVyfKfNJJi/HCdkyJ8xo7mUwApTFvRMmpbbkq7E
TA3sA7Gvhf1FOmQR9rhJnpjKRaTB0wt4zYJZLCxJ7pxet9eeAnKdV6/0DbaXsXaP
CL4s0KCSfa24AS6l+WBBPf7iML9JcUIBHp9Tk7kFNqPS27k8YVTjxzmCzsDeheuB
GhYWxh1R6tEXQDSP5npdI3mAvcxQ4rJvhceCZQyvGUrUw9pRShCxJ++FOWgMirfP
1YjIv52k8mMXZGVyioQvkrZkAxeGYRrPA8BaF91g0P0ys1LvB5jM/Sy6iomrcJzm
ks5qj4QYwhH5qZynj+6F843XAlJCa7qAUg2IID2b2OvrHZTpxRldIW5c52f752+a
fiqPtu64oLIi8v5Xy1cLHICfqiLCplnjONI1J4799g9pMh4RaXCBnqWAXG+YTtbJ
duZ1CfuySwGDIS05Xqvd542eHOECVyMkIr/ZfKrQiaizz6ysYHiccHh8sIKppXaf
MxKs6fAW/z+QddwjExf1MamDQ7b27vhn8Cd0RkUlLHXF/jD1v2oYgaiGoqB+aM9c
Ppw6MjHpqE1rsNwKygMQXs2pDpYF7nfzmbUgFGYHBCgzeW+7/R0Ghk+3Iu/Q2ndK
YJrt7D9+ekgYFeNN4FN1x5lzABe6TjfzLG9jTu5yeNr3nnu/shHW28mPr6F3amzS
DYUPQzgLhkAmehigFLEzvn0eLu4nV3hTf0xjiA7rfspp89EWSv1TmrTwkei0IDbq
bMSt0QrHmr18Usd5nRtnePpoVMmE5V9rsjGNtrwPdDLi+XaW9nwykCRk08nJ4hX+
0oR0nH4Bz0xDuQzPmSsK5FAJDv3+QFlCH5hBeCCTjlkwnf2p3MiBbseLearcBWv3
MZWe51xB8yJI7UOCah0X192exIL8sOL3YUugWjRWQdHvoRYKgPobHOTElt+/sSrb
wBmdppm0yD8M3JVTL6L83FDismPdFfCz4fvuz5PvpjpRXQWWTeUavVwgdqCE0hV3
veC7tIHVC37WDI+o1HYCMev6D2EQ6wyExZNBZMGxwQsdRZG8NeWbzCW6Adym9VT5
q86MTIIOaXyLwkKVdOUxDWuYhrDs//JsDeO9HgjWSFnYyA3mrm6l2YNMHtu7T9lS
WmZsBsc68fRyNdHcraHQKHeDxeAqOp8+Td97F7GOOZKazxLjh3q4Ni22IsUBfXp/
5YX5xjALAiexjRH4EeXu9K0aptfRTBj/C2V+Prg0Ry93+D0IIAKE4bOOlLfd/8mc
Sg3snlqFewh2/gdtxmogJgFUBiI/RB3Yn1kY/meqlCmmlv0+UlAovQaJV2e4u2YA
hNT4X+Meehpqns8hrklPhgiOE/LR9QKtD5jHx3YP/oJ+r2awqXaWCpGsM2MuL5AW
qbJykY4cpeQA49QgNXk3dapieICXkjGhTOa+eV7aFiX9+gVle1KsKnZJbHX9nJnz
+y/C0rERic6Rf8rVLL1dRfrfgaNFR7fc+KZUIKEz4qPjSl+lQ6xR5oTXH1ypef5d
07vCrq7fXrVqOoeNMScFcVV0zo3Q9yhoTEryC00zs5oq9lespc+c+/Gi8TGTqf2j
Y5GaWR3qhAGnVLWvd2u7AGNuS9EtavEqkMPDJ24KywbzFEzhzeO8wA66Zn6rZ32w
cO0/qe55F25uS4oYrDuiLbjNgdpBRFTrMW/VDLoC1U+o2EuFXD6mGfMt/4DBF75x
QxnxD6tM/xNVNYk6LvuRUV07J2gsVmNaO+mR+goQyV/+syrUOUw6uPcV5epq0D+h
e3HGa+9JyGtTB8aX71HztYWZGV+SKkBFMcWbKHIMib6op2xaUhFDb6pgf8668F69
X51LriB8XsOlahpHkBb/5KXj/G8IoFmUgoPXINiWILk32aLmYjxZO15Y8RtYNo9X
if7hrTbjlgY5QS6oD4tZ82vEMqVBPlxhcNdPNkpLjUW4quiFIDdm9tX5CnstvFh/
q+hNmhBeQPkeeCZRjgxaBgv/Pcyb73c25SZduY0tmpliDbb7OYrzb3NDEETpay/W
p9xS3FjXH8xg6BPM9fC4P+SdLPvD+S2Dj3XNrWnpRWq4yEMfQHjlHy+/OpRuvSeh
LV0oIw9zIWOvO/2QF6HeltkXzCJBxLY0etg1HI0425RBjwqZLcqFT3jlL4mE7oNQ
5oBu8NtEmLBfWxv4z4usAzFcUMRAmWeuDxCzYGhgtwP/zJmOwkY2HROfV4nauskI
DNeOuydWPR0w08WvRhBr9eeqgX2ywnnIcuUen62YfT37fLMn/v8AgHcjv+uM3b2U
kP+Ghf7QoZwYllXQqhjaIyLV6eyVV0I5weNKw18z6yWnnfKwPiM58yaXc6fzX1Dm
QjIysZtsZDHoBXwCa/NH+MBJ1IBR9VAarfT7ORjEDhnY9t5zeLffurpKsYu1LZ0j
rZOi/1eOKFXf0DI4EgTP6efWGqRiRExCpe+JSayzloAb3QSei1Vz7cpwYDP5GwSh
EwHQPyte2jfW5MZau1kjGmNz/G/1BuzzG75X/Q+MIvbvgmqPdATh4mShjwEw/MBt
Y49t/uIwriU91fTRlfb8FdWZQayYzE4zVzqAiPfwlH8sgREfoSuVC6vrv+oa25g+
rbN67jYWabtYOUdzipbIHxNf6oYoliX7gsE5HZ2t7FxOnrRdWIfPlrj6aBvGQsQJ
rqax1OGp9KgH7uE40Ysnoi1K8uLPOYf3kaQGs9+fHAQ9F59cvQogXcWTWqq6N0/d
GkS1JDICHFIVsVFCEyIBHMJ764KZ43EH4zfhE5exWgiuAkwKp6EZE+EO4K1fg9zv
Fbl6D28VvpuiuKQHwnEbPl6LWXrWoNUiVhZSFEk0cUN+D3u1Qkeue/i8/HfQO7yw
B/TYDAbMz9iYAuUhY8aK4BXRK5SZGTSZo25Mc13MyTy7V8D/5QcknR+psZLs5xYR
v9HRUyzO8QpH0xp/WWAwxKxFbfRtAuo+L0ZRrTF0htrWHq6nTXI1eRfzgS95rUOP
4vecFrQfEHBAS8xsZKZc1ZA7i7jvQspYB4rVtC5q5HZfue5XyS4UcgJY1aG4jDpp
JZaJB9ArBNad/IvwzGXfza+RkfYEMB9hJ/7p3BwS5TdQcbv/RTKl9CHopgjXvDN8
UOYbLoyOC9kd1ln7JMJEeUW6ZR9wU3mrNjm4T+XYHrfCNAdnTCDaG/9QJMRGQI3Z
KNHWV9G2INeftDLE6tztTRDsXLm6S96u4qSLD7xiOnWSrztSxpOpvASP+AlxqtF0
ISKIkZuGFJVOB7qm3Mo6ZlKXEcjY375dXvsMHAgCthYuxIyKPTJNvKYZDyqJjg0N
MbgQFKnODcOdhXqMPXhVwmVq/5c2y4i35ICewRGpqtqlfvtnmsv4UKbunuumUotV
BoZxuW7XnTUi4c9jml18+xksLCIMH6g4kadKoAYVY8HtSe8AXEdKZIvXJY0FJJD7
uwC7aLGCGd5vMa/pbsV/MWe7HS/SOQQODP0dofpGXX38MO5gTKArf4RpTnLlO36p
8hEOsr5FPnxwyB+0ADChYdI5wZHh436iHB57pESDals8A5zYRVbnfN6B9cxRmszN
oOJQo4FVnXIrBoBoinpaxW2YXtxg2LJOLMYNqYpuiXRRvHfKPNTzollOLXXwLO20
Arb9zXiIVmB+fUa9qgt38kRC4w7ngRyf1MVodEmE6N8+HHSrbVTyQzvFzxG2wT+j
JZyKpvjImOXUi671vjJydXV8BbaPN3UePHFpdKuEfe6kxX3uHN2enqnAgC3JKKs3
jFUynmezS1X8SAGyG2ru7CSv4Z9kHh3ZYW8ERmviqvuwuZUwRinBGt+I8ARrSB6l
LrmI3pOmL05zzT3ph6mioqf7oiMzqyeJzLCgECHsMxYieFGZ/AFNuArZo/H+YKjX
LKuZg74Xaunxh5cYFq+kHQiY6A6UWVa0EOeAqSf8MBbxThFqaoETZ7+4QNecZUza
8Um6kaWjZIGmjsORTJ5G/Baqm/wDpzZn3kU1l9qAW8Z5R6x6XXttJISPSdPiSb6v
n3WGR9dWBkrutrcGEOtvWObXnjP2LPey7J5t9uGPGyk32ONtk9Ud9NZfpCixYhe/
w+yGg8nK75FAxgjqSyE0mfRLXSIeCSh9pmSkxBztklh1+PMTMetWfTdQKkTqedfK
uEcqJ1+TLppKQr7BDlpfYTIkgEj45npg/r7MqGnWG2Dm1FQUkRhnqNDU5LP31Kb9
dbiOU42jebZhAJdqG/CmvsfLd9Bsuys+IQmOt3ihalTiRJsRT/cx4fp44zZFWMPA
CC396GveH5Xldwo4kjaDLJhW7TAgqdigVP1uMdLT82nJ/sIg4CXPTZ3CCwkpFC6H
j0xUJvuIjXAzwc/+Fz9KJwoW9EaQ0Zc3AGwxNZG9OFesFPuCP65XK/iaPQa+pFiO
uADkmtBep91ZXUe4J1i3lmQRzND8TCC2Txh41RKFURLxxfqLLgbpIs+Hm8m6Tn4j
MSx+iFpXTALS/jFxdEznC+HhQxtv2V8nC0kuJxa80p/BrUGup/guR54hAfLn6nHh
FfRsqq8q8Av32YIOpGXk2DsBIizuEjj9YQpw3LptpbBp9ykYt22fEYcVpYX1/Msz
L0p24M9MD7jtoWqGddpvghPX5GoqEzhqhVobcfF0woRjUVbPDdlzQFEM7cAMuTSU
RFcmAyE6otLCn3eQM+1T6PxYZX5tQkDFf9B75eqVF68RWXibmdpHrdcAmvSg7uCB
LAlQFXSy2qSx+t5xjGkH5j6acdqFlfhdWGeYit2nGJ1XVgnhcwiYX7L/qmDjk8Fm
TctoeaiXEmnwm3wRozo26rYNDkUQOZsRAIV0y8wC+Xy4J7eGWA79qS9jGvYS68rH
5976FpG651D/uU8HmP9nSU7LQryNgI/Uw4z/e7mCizh7//xOr7az4ghAd8T3Do5e
Djob8G6MzBggmf3EI58RODCT0pbR9lm9zGPuR70Xd1vBldhjPYfjC1Lvy0waTGM8
abhCjZmdUuGZZ0q8eCrkdsiXQQS3ihmqVOTiU04izHOqUsLvUEMgBhK5w2mXgghy
wx6h/ssN98Nc1okUreW+q7g5shVhPe5gE+HnnmNHOAISv9rto2GVq1x9nO+aLvuT
isToikvQmJjxBLBlkog1OTQ66DqY8z4qUw0msc+d5FH6ZumQAAG0L38EEOBsmzdY
6pX+V0Fb2tHM0bqBZugfBcOGdQzJF++Nn/etEKFw5uw/TpWQ+zZvaJLes3tCFZau
lG5Isl8V3M8GK3Y5hdbGXfPSzym9+RL/e+vddTlIM6C1Z8QEpAmWsxGdf/D/uz/N
tRCqP3+2xFr5pUAVpdlDKiIz1V1dv97PVqlnYzsrAuxHSuL9qMCz8Y0JjNtkNA4d
OslPbVI4uVSXdPWcutnOq35GqQxX6XqxNHJuQsqTTwdvDVygqDCKSGBdokxI1/r4
F+lbGxQr8ICwRtOY0J2krmxWq5gp4u3Uf5ZxlOPqYs9V2s6HRgDfNCy/D8gfy/dF
H0xgwmAsdAgJgRehK8Xnj9dOm7oxmQEwY6cc7uHE6SPWN0l+BWhcROSBJbRBM/Cq
gZpB0F3ISXdD5cncayoQFEr1MDfTFSJBq5n49q43lsCEWGOcigZGTE20L0EdILy7
F4NwP/rq/wCM9L4tDRznobQ6Xcv3ePOlmMqYrcJJYF6fUBhKQ8u4184CmYz5zLMU
rIn2hX0DYg4UkoEnfipy9rRqEyRfrwhG0Zm/AfKCPy20zgOIN8R8gW7RJka/jyH0
3pywOeqdNrPiiMicvywwRBp4GSV4iJTlYzR1M0u57ArJ8haX+Pp51BIkAN/GgKW3
yzUgM3kTjvnlcKoglhXxtuT/3pE+kj1Evl8xLvzQUZvOUUXPP/qYDirvJb2zP9xA
S7dameN6Yygkx2kEkCySb1xE7s237ju7truQQpgcNygzbMN78mpl93VkuP4FDD2s
AFZccDJa9DF4KIwJK9JJo1GDBOky3X/V3Fe1L/s6DtYNkl/cLhHrE2eKk/ICb5R3
uEd4QGMr/BwslOe/Nua3bA4DfzIW2TNear1B/hYPw8Y06k2rJBH8DHzOHOfJtueR
1ZUpu1IytVWkRR86KYGK3IvQVQE+eyrVkAhMu9uKM2GisX0jYIyUuIoiSybXQaQL
G0vjpyRMENOqIPLZoG9hhD0s1V7UPQG1OLYlkZX90mFfxIvpAQBeSGq1N6j5VTZy
1V2pywIjHHfZ90esJy8PtM+9zZXDze18Nl6snAXzcoTSDh5Kl/di60H2ksj9Fzwi
2Vs58nglkbATQCOu6ff2jPQ/+5XpQjTx5JUHGPpmaT14WGiPi9ZQTZS9Mgon0YkZ
ccmBE8U3nhOijGwZfxTBs0jAgF2ohZYp09mmWv29JXEpYVxvJqcTTo7LaaOkEXV/
2kiBQp+VZD8AKa7m1AKFNZfXfE7uq5W2/ErdlhZ9uowYn+oXECNXN1iAekG1UmRm
zDuVCDahKvxAcwt7dlDlbTVIzxM/E8qurLWJLnYccCiRh0bORY1XCbzK+S5AVeXt
EScM9XVnB4ZZnTDXDKEwejou4AiF/nUxGlT4P94KMy2Ql09/bqSiUq7VIGc/TF2+
KiY4dM9tG9GJrYwI+rzAZX1qMRznoRJAYVrK03TOAL/mtUiZGei4HilYixQ28bxc
+6Ui668HFLx3/H0KLeE59mXLT4+tmofvOIwv2AbwRDYDwx0EpmCBRaZjlD0BhsrN
yCREgsrMBnwkLy+zesxUhBtmE8eY/nVBqZslJawJzkw/7yY0obTawUh5nOr68xTe
N+GK49PDgRvUgU8wZYbzt/xRWxXXZvpp6QTXefIrjt2srbffEeUI/bWzQFCKszk3
MyFDJgJSAW1xnTdamOl8jOduQXWZCBI3UAV6y9+rlMtudvehW+/EGRwosCmTjptN
KUju7I6MHuLH0+NGCwpaXcJFzLXD7sxz+ktXnp8sOuwFhnE6cz+W/B4u3dS9rJ6r
I46vmbaAzR8PLIo1CLBBIGYKRo+hCa2tA3V4Jhtt2AovfxjGwm8HVm2O+mouv1dE
db0r8SSe6svtdMkZuX/L3OEukeJDtabo7ZYq51Qa/r5O+2nssXer8gbSjBkdsm6Y
BaZaMzd9d5peTljxg3VR3k/UTnH1ricZ9MpyAb3tmYh8n+v4H3UvChTL3XoxORUE
43TuflcCY2A6x0ccmGa/oC48hwIn2MUUgI3GK6suP9PmILsOP62TpxFlps3Gvv/B
GO50YLoR6YgPp9CiJMkSs5tBsHwLZTDzPG04+CtyyidiZreyJYT+zW9tfzGpgOxz
0Efed9f62Og/qmokISfcUzlCDqIPXvjIiLc64kz+GbSkoS9Hh8SmWo7v2J79n47u
DASFz8dnYarD/FWUdhe2lStKqOaY3GJi2YtEF2WokXIb0sh/FeftW1F3v1SsBuH7
nWBg6zIT+Z6Uh6Z9V7pQ2ZltmbXHXwHm2nm118RRAbiOBYB7c+QTEGsk/VBb1Lxe
2odsZRJ8ctSjRUstybbngKtxKuFvm+lJu6Z7vNkPvOSxiQoIz3ELGffld3SmZGqv
jkdXFeKrSSNQdpgwvVQMVmfodTXTt8+muY4ueqoZcMKWLiJ2mDo6Q/FmI8Pc39Xe
ZKZwR9yW1/sGxl5XJTMiQG2SS6nJqnLQQ4dhhk5dDar09lVI0uGfsl9Lg1iwp0IP
zFN2v19GDehHqP/nUz6V3kczsMXsZZJEIthcnUdRJZgUlrcRFrBz7J37qFIxAUtE
uEoK9PJNK2149jWls+9eLb52N8iSPWv3WIpPOd+SBz+SYkoOeOGy2Cn0rHaX6qz+
HpqQIcvDPqL3WfxemU4Pzr/L5Zu+1GqQqtQIjeY1aCnJcOy3d4imagxE3QtpnFUQ
Ubx1LeAPKqU8kpKujGFlnIvSRgebeknN7v2Atyy8GbGXVkDhMEFrLChUgxcztISD
ldcFPa1axj1w/W7e7Ebs4Pv6JOWLHDcD3EDXY1rA26vxgkRRk7617bMEZFe1w9CY
HGjn7OC6+bR2s5nXbA28Mxa+dsDbELm9OMogg7bBM1Kv33791mjRJab3LDvACL+3
sPgIxR/sWaTrE+vbYHdPPbR+4byQiRtirHMo252xucxne7sCFBGpKxF9h9bGAMek
Ix6TKjh5CkKhISPD+OuSJH5KeD5f7eDaH5DC2j/wACOVtz8kcnCwZAPqEc1saKhq
bsoP8i57laLRzIAKp5RtnmZpX9YoNFTCiwlgpMugErfEkBV/I327kSZSaXizT03k
2eLLMA5tDFhFdRBps/KF3YCeo6cUrQU2bBBd/QmPYK2AM1c/tc8mEz2J9EitJgpK
4YDUrJobfZfGKto4WCltjQF6xhw7ASFMqmdqk5YDQ9QO74vE8g3lUgNKfy+OXM85
7qS+Mn2qKdfR2Fpq9t4zXGwMjOocf92eX580zv1RZkYG6EcJLNRlmNSExx0iXdXd
KwFeaLz+B2H1nUuW9UqOWXuEXB6fsl1xBgJKfixJJRxqKkjapN0l92EkKLAZnMlG
kAEYsaR8rkKM1cvVs6SGy0GM4Srgo/ip/ZwA9QVtzLSi8VI+c9JQoVWZuxXx4NWT
r+E+ZSkhQiu7WZ2DFjvjdJa3e0+5sxEJynY7BvNTEV388FI3OruPVb/Z5GkWXQSS
qtZXLOLCbHYSzyq3Jatm9TzOFS7PtIcEBt07picDyfxkH4Ad8VQptj2uJcMYxO4T
VQFcJ65V2iDwUzoNkj+3PtF6fO/Shh0ocDFWgWY+YJCLpHrxC68ZUvswKTcqCgMe
XX9GH2h+SM7BUidYp2hzEdn5LVVaMewpYJNU7Fjri0GyLjfX/qZI62RZOn2ZQ5Vv
gtO/dg+Kqvcax+hym3BNpxyftz6LxIeufRcessfC7q+DmaL9zNTTN4A/yqwUqE4J
XDICANh6vognUmGcKt06Yed5L1omyZd++f9bJY983FN07LNO8OPHnEslKpGLNt3n
z0F+/KTVVoTba8/5qLZ20CkV2xwByKF0TTlXoksad+OabGyQ7F67B2FYqDXCmJpa
SODNDRUOVBlFpUbWXfXlYImx9ph0cSpu2V5THoz+IFVBxedh5lCffDjQmJxFkQvL
nUTQDmdwQ0teYKuuCqsl4hxMs36Dr38hasfaSPpQ8XVrKF1NgN+EGzs/Y40G1ZQS
FKr5aD9+MIdOCw/rjTPDKr+aY/mOBzui9YpNdUHXlz4RphS37hwwQOR9K6Ptn1Tr
BNZP87QaPoK2WOJS/3Njhl+DvLFYLVaY+UGtJv/quKNU7iprWxMPC11WEUjFn0x1
67KIUiLo1zwtGf58CkFfX8v5u8Kq6clzsGaw7Cs7iaeiXbQKGX+zxkbTmfxcQvpQ
FsN8S3ZPPEBJyuiE68jSNxHo93ttXcZ+KbcFsFOFLLeSkAwsJquidIGvUX0Sj7y6
oSCPK6wszAeXBKQfPovfHM7z9RWB9xPVWYtjpuogo9iG7RiVW30+9ikv3BhS38m+
/L8W+GFMpOyTCsZCuT47alQNBtDmpGIlu32rmP1HBp21376ICfS3iYg8zGOWhE4Z
0Y+x4lpyVCNK835n2qn+ywD37QW3Qj6hXrt33ZWuI1uC2AH+RM9WAOqjQCU13+7B
qb6hO6ULqmYqWsqZb4kVE92xFUR4rgoEAMV4Ftckp90kLZ7pe3f2f1HP4DyV7WtG
7ejsslrfuleU9R1ryGBd6B7qvdZZmZ0waYIU2ASTg3058nwM3b7HvW1opqNrrQfo
kKabxOinWvrCkjPoJq+Hbzdc56pozJfxF0CQDdVqN1vPOKrseIrhAYWccmq5ZZb/
lsgqy/exWEQjQbFBSjJv5YMaxUZe+3WBfadvdGnCB5E07CDhsqnBVFuQqiyAsaLX
Xf9S3LXd+kQlDXfeL8LlmHyKpg5bFl5BanS1KNrMPjCi3GPjbfPX/gPBE8W3wRrH
I7Q6Q5IRKjcggCSM6CMMCqSOuHWpoBMbyaq4WDf4NNZv3/JnR/Hz09x2oiUA+iWO
7mYMAo5nRVsabW/TRVEvruaRDO8qmR+B/A2yG2BLk98NQnxlz4cZiUXSspWssGez
NUHwAtLIr8ihw6lzhk/szCPZ40cru2cj51DV6j7pFe0MHd8ueCNWyrGbWlL/5BnM
xY1dnl/0gyUg2h0MXnCGKUgYPG4GBs0fyrHN+PTEqanKx0j7CAVTL/CGr/GQzdwz
prMRv4zorpWePz+6NYtu4J0V9S/soQZqIzmI4EadU53r7FAltYrxGSj13jIsevVV
kq0JEZQtRM4sXHl9Cv7HstmLV4hzfeEA+CcaKZbOGMVaKs6cMiwg75Pz1EG7P51X
ZV2xMBijnGmOyxlVKfWFsbo9foLp0KvyRc2XgTX7nym2cruzLoQV2fU9LaIIiYaa
5aKLIIZr3DHn44DdjR18HyFG+lypOFLb4VIThUFN1HR1C/Azls2N6Q9HDqQ2jNar
44rT7UM9PyaRsDLjzVPxjEGCGNViNgeBPnijplARBnS82QSH9fatIxfFtkGnU1Tb
cp9ScaYkGrahDlhpaBacfmDfdqcurdI3OuH4kkujDsulY3P140Qpqoac5tUIbBLZ
C3qlPF90GEJ2QLBi9EhDmmO4vtzo5kJ7w++QGIHUGZZUgWAGbxtlvv1xcsIYP0H9
oteHhk6IsmRq+f9cCHtm6Q3azhEoZedufu4Ekn6we50ZQNkOwsHVeAX81dIfhcWm
enZQLLa/lgj03CH7j03CUFlXYhHihwWCzW8O0wrO1zB8ZzhYIgBbYHR6NUjm1uzi
kW11N5Cz7RoJ092RPs4iF/0p8FIrE2gVNe4bq6x5/2a/aH5ZCD7o2y/IVXOGy3uH
s5vMAGPmJoD12pFHg2LHFD6Ic25jmh8RGs8Lz2wfEEZSAPmMrZwDozUklTgU//kz
jSYD/2Vw+7dunMQ3ovj9q4YBe3AH/C+TS5Yp6yH/beqPDU8YUNgM0A3ZdN8mKXMg
33ax5saZOhFHi9adNgszfN9bbttARBhhYSjmp8pO+ILXnnvNOJhLHBPeOBNBmJ8m
UUahxg5jVLyUFG9psCUEHpWOjJv3TIgd9yD1amh0lqOCB6Sw7UUiR75TnB+kxAvB
qai1i6GDHRNvpq5co01W9vqYBChYL6b0tfq3f8TzW+qmOjvau/38U24HJGZL889f
98nHtAKWigAqAhumm3mxj4WbLYxbYga9x3m+gPeMM2Gcn2ck/8U0fkUJ0Hdvwg9l
qQQMgeaWGe8Cm6C2Cx4sGtWGEQYjaUs5OzutDEf0gl0B/EWQPpbphuRGHiWHEwAQ
eBlyM3eNiMXlhor87JExx+KcFu8zL7Hm46Je3AQQ/aSvFi/yAdk1JEJWY9/lrDX3
iMGn9wP9j/ZVE7KYH/QFnphS9DIqD9V4JLyOFV6aanVKj+kH8QqPnZ949E+44dWU
ALVpQ8uzsd9HNwPK4uRMKlUTZfLxMFndto2T79Y5MEIoRCV8SwSkY80ZYLxutTgU
nrnKd3TyV4I734rDAJCZ7VzbcKL51uFaRNb+T4KgvxSYKXl3KiGlnww/yMcJe0hZ
Gmv8f1S4cTWKipwjp+ImBqlvyPazKcRCs7xhk5CG63qZI40bcxBHCxLoc7lr7RE/
Z9dJdthjUlnhOyCVrXQBuD5k3bxwfN9E8E6x0aEuV1X7CKSmMHCWhCrFsJ1Is9iV
y58aC+jyrT0TLYheDXOOtTtgZFTV4klq6wQTS747mgW+sqE/TwueYzj9vJi+FuCK
+f8mcabPonEFFU5eVRQtbt7A/jHK3lSkQ1Aib5QwhhH5+1Y7mj8FkLoRZBXyb5of
msfTgUj0T98FbwMFfsmxGjG66zsTok/b2olo18Aq5MJwJcaIRvF1Aadx6j0imzrx
/kEcxODxZosOMRkoMQpxlfLFq4rb1azd4Xu1IwSoZG3Fm2SDcIPp09g6l5MOS9EB
GVLKgnIV0Bm2De7WlZ/YWvad0wkXPzaxNOFQyyzo9AZbvcWEvaGBCZdJoAN8TvaN
DACdDdR0hV1Zd7GDbudXWNv5owzskq71DQ/fhUsnsEb4g4/WMKfK40bRbPMPrqL/
7qEtd52hUMk7gHlZSfs2saH0gyrUILJkOSD8fnXq4BffBn0O603cbbJ614iR6nOv
MFUQzAsEqzrocbiUQmw2w+e2iHUe3jKtHjnCXZ1tnaRFfUVQdAk/LWiJKlsKdm3P
YWo0tiGsii5kER/WSJMPW4G6Os8CV/5Wf0YsfWi0r1zrQU7yYoQ5tOjI3Jh5fI+2
gCglscUaIkBaPNq6Eqel9JG+z4//ZOlF7EPlhVeRWeyKakeGFdt5SD3Klbkifh8H
Y5ej9gpnPpQ/D2jFka+aJzjZ++pe+jWy1edvTAqQIUi7LKARIDc9ZWeIz67ItT7s
Tyr7TVpnvpfPNe+MJJ543CG30KrFja4Vvcwbae7hX56ytHzi1ecV0xGyoPScsO0/
F5GH1T//wi1gg76vVSmBIL+RR3mRZwgA6MIWp/tbIWe5O4HW9rj7MQ25EQ53AlCT
4xUFpTjCKd6Gl8MXQ21pJ9zd38nsItYzQ9hvwe2Lz5qbgqeVK475dbcElNTX+HKj
2J/fx14bvnfM3jPURN1r/XgSbYvc0kKXRWljX8vQGxwk2B6cDfPiCbNnN0N27rnC
7BQG3A81QuKsNbK16R8jQem3Xi9D7mXBXS+7texjgp+1yyAmcHP5Z47Sc/GoWVHk
f0wz+WDwOUNSdBRaU5BSPfUJfWg5wr4yctmlf4BTr95v0Ya8mZPLd3tevtGOKYfS
073CDU3I0fA8kpv5bBBYUU6IuDSOmAhSl176JDmH+1HqOyYFmKx6Lu3F/ld4r3Xm
JEEhHxIOuvydvvWz2PeYHGKF673Out4Anmi1U7V1k65IqatiViC2IFbFV5aBaijl
DdZdwis9xlnI2EH9LRfRBn4E8UUT503dTazOA2Pfr9DY8sS/qomzKUCwE0dEWj2M
nthF9RIFmEmW5t+i2afJKLdeRgT8KeG3yUDpWhjykry+/LHX3JzlT3OiaCTt/7vU
Sh4u9cDMR1gaEc8RLDD3lf6/YKgYDeDHIEfDaEli5v3KwPtrsC+zAe0u8g1Mblz+
tcthA5FIui1WmOvq55oamCndfNqGNBQWSF/F+38bxdugOiV66RjPliwBwz9J1/ny
MXl++KyxkQxMB5xU3a2N2Rjhl0B5o+Pu02qhBJwPMjozB7E/3mFuc+GwmztVOj8M
U1t7dHUBGl4wJ5n37/CyRwwI3Nnr1A4gPc5fU8ZVwnVXXXSiiDsiqlGqVSNUn9iF
mQ86AURUP4Im8WfIx6X1sHh+fjRQwoAqtBYhuv7H4GTFMQNEQk07jSB0N5Xq+j6W
iuUxSKD3+PI0xNtW4cVUVymvrj4NHIUG3OA7t+DuhsPr6Gy84MmNl3CpLNHcIEPw
TMMswdePGzkCQ9PVTDDzBEevJja9mblidJ4wvmgs2gq/wL+/eTkKFgshrDRwxRSA
nS5gnPVTfBwm9BS34RpocIYfjTYaTYuvLR3Jljle9vNF+fzcouajBdQtT5bKkzo8
vplG9dVBDXUly+poNvCsHmFiL13vHN3cVEWiFXLcM/F7EYn7SCisW5HXfPJ7BdTi
JH8CX8K7g09D+Cw4cx2o0N9Cg9bAiLhi4xVmwukbNcVBS9aLK/AC2cGiNjWkCexS
E3GFTkO82fxJdjI7XuNpV0Q8/20nnt/1A1tANzDid4oBPPLr3cTtmIu2/e9EeDJT
LWP0KDaKE7ruWaGnmQJW9KJVm0CHFFAl4FUERXj5tKIY3bKf5+vJVATvrqgyWDJH
YZqc/zSga/rvDEs4iv3c3Y0P1Ut2YBjW1GgV++hHOIlDWL0pZkXY1qohEa3cDYJ7
04p6421+m3grsP0ecMpH2+zpA/l4b/olbT+XleLeGf7SkTfMh0m5j2y5SlESkDXP
XTwiYryTQNYymoq28oGSBN6aDK/jy6llFYph9cl9aImoBhhYIMsSejQDe5ii3uwe
3OIRshoz++9GL/DFyM5HELPC5bwEcZagjvI1+F+3+dtdz7dSsaRGlLSDUKMVxxX3
yxQgeMoVV/D+aiH4Ge+ckvELNpFfVzTznwE+uaP4zW5sHTE6p/3+jRZz0eJ5cQXK
f9ZPzI5QS29YbCPcqOjHTHb64V/MHMYcvn8WB+Ll6/SYLo2z6Qathwr9iucOBplA
rmZN1jIl7CENy0PNiQFTWqzO5YZZbghCJjF76Z2K6Zfg7w+z9UiY4xG9P3ZG/4y3
y6QEg/24jBEPE1eT5xoO0txnccowE4k7lFr4UxOpiMbs08mVO0Cf/IPIqmrLvJPH
ix0kOr69TEUhXj+rflBCazmB7Dw8LENhRky+m7cmlY0B1Z4GOl6PYUaRaBsgrzdg
ouA2KFK1pBeh5L3llxwDxvre8u7PfGW2Fh2zVmZQCfWvFcl6OWI5Ai9ogPXItOrv
vl/OumVhS3vM2PfdKuDpz5foU9Q3+7EVHDSA2kK3XwSRI/ucNLvxqj+OYFE/TBSY
rz3fAk/ipZtl2bo06/tH97kbynLGPhViaOulsZI3UqpwtG/4Fkx0sWS7R1Voa1ei
oOPIwVQr1HjzG1Zw+TuevAFxNKR6kuBsqoms7UflxPChcO/ADy21q4uLFvFxOYD9
ZMUJB3Eo643pDIpAP9uV45+Ad85KTA5FSops5NvkhT47nfqxv6vml2CWUvPkxGvQ
/YpP4qZVkpscQNz1t9e/RvJQeOn5MB9kaVMuD78Ry+pHIdNdb3qm8njb79heU+KT
smbowNr6uiAVU8q6UpEkGf63VIhHkapX5d6Aowx8bh9uUtHcb9T4V5I8jYgbcKnO
oyTcWGHIReQIVpFWemRifa1EyJJ5C7gISi1jGDRDndSsg/y6AHQ9UHDmRQSodzJP
Qh73oW+eSpM/ee1Orf5UpsNKNU9mZtb9zlcdL+xKtSPwseyHtGoGNVVzfnBBjpOo
Z9v2kY2yXBYwzAdxJ8t1Kb8SWjaZBEoIp31tnkuHx/GJxBnfjOTzZlG4lzG+SeUR
edc2oEEtsyau6aCciBUPrl+dXS0DiFpPQtNWZtorYigk/uj1YclFL9RtnlUovqEY
V8Nb8WNwZj4S5izorW4jG7OB5O9zeKJLSOVE/gCqSgT5Ds8z+pPwBEyOxR9ze97g
Sov2q3GKuauQD+7kbtL97nD2lghxSzQm3pBjh1qHBSm/p2cKC9MoqSxfTPhLjsOI
ECsxkhvlN5gjGbJ0AyOsqSOGBF4vRS02hB96+b/nSD1mpgE1kbLQJd9J6G+1zu0V
P31+0w9ESBk3uHoayPi++J1XdMs0T2cCi+6zIDLupS9isQosZkMsncmFlubN+DNZ
Ys9dJDufdba5JILmSCf3566SSaDO7Wwj6+oOyDwQMSG0wtGgSVEobMIwUZraTzZp
pzl+qEQ+79SGt5bYfUtijTsjw9/flu5R2D9ZyrforATeFJrG4y4oYwMr1IEAKsrS
hVeVG5BlM/TQEwYbd9wXydNJ+MXVC7YxINCLPYsMR/osLN990YSV6doI8A8at0ZP
fN2zAdyXoDvDmScC8LBlA+AdY6MXTWR8D/SH4s7CVCqyO96Ro1CwG1FqJ0w0LMyX
u1JCWEKmmaqWrNIn7ppNt/ltQbrnoJScDaagkK4v0Z39ZkPke+Qzkq2DAViMsUFA
2jKfgSdgt966AQmS3zZVI/geP7VMopJwoC7CAkG0oroZo7uCupULKn2ws2J/Kjnw
Sr86n98Czyd8b4KrJrMj5onRs2c9To19/a2rr68kBT+tVs8MWNJ/dOP4lS0jgKWP
We/L0IZ3mliOyB+38zo6fUFtxWQE0nfD3BU1HIIF4Pzg/eV24x28ou0ZkvupA2Fr
aqHl8q0PL86OdafnFx5JCgKOmD5I1HHPFIYq630ohS/N32G40FKG7LiL4BXGePpo
GB8KZfZF+AZY+LwEvq0HLApokc4aoLIP3+QsijQC8Lr0gcXs5DK5R1QWxPPLy94Z
tRHFGhbrKKw4hzWGLHGl7utYyZVcWb3ElBij1NPq3CMmbwSh7HdpnJsmLXOaV3rc
Y4yGLP7FH+ZCalDEB64vhVxJ7s0iHLCgunBYNazCzwSRxH8cyTZeMOmK4GRCb10C
w+/qxUVmo7XwH+s2MK4bSK0DbWaEEjA4xFXi3c1GqehrsdFWvl3kClN8rH5b8b9k
jk80trkXDzb1JS2biMYEpsdwnZj+W09hRx18Rb6EriuLce2dzU//mBq5ulWTfKDa
1eS7n0g9jzp+g+mfNaji4exRzPeL/YcoZGWY9ZYwhMsbAh/CKkLgwAj5e9Yja4z+
KTBps7xwVS0BS33f455Oo6DP6vmOGEdNF7rDR/NHFAXl2iUZ8VrpM1I2a+QKFtRP
Wv5zszU2JbRvHr5JLmEJwYcdOKsANrdDXeaIa6fI8mg4f4DlR30ROgG8u8NQ7H5l
O//9obaVv6BF9WlSLdfyO+pgJ99wo33nAzlZQhT7bzTuRNxzrmXwKku6oGr4lpxL
vKP4IZZLDp1YlLEhxdL5Kap+stE85+WSN9OHPOn9kbwSvxX0HUzvYIJ+/CmnB0gS
KTN94bluHa+rKfbq3dpPKMJE0ay4fuErenqBYN/LOHskeFCdkVYFdB2SRU7wcROx
g/2copouDRFqP6j3ttamo8dyQaHphcs82HKkLv2RGXhhPQTA0Ip2qX6WsMwCFiBq
sl2ksdWPBfzxy5cKFSpeSSRM3cY5+HINz8YtgvEobJP0v5AqxXCKq3TAbtpk4/DD
m7aiP6BmZzWlrEY6w0wRSAx5gvnctErI7800Efe0RKL7CQs8tEj4DUvnRDqgGhr1
ww31EYx+VymNSlEnNzJl3ydQAs6OlpWq733jXqzV0dtG3shtusl901b5uw7rUs8T
urJQqnZjSnz3yGf7ntixPIvpDPjP2f/qK4a9TqCR+smQ2Fut/GOvFhepKXVAP9Q9
lPW8RGYJEWPnW8PYQ2bupkxG3SZvs5V2G4L2OdpWL6gVbRTfAHlzz2SRkOBGOADd
xrz+otQSSWrHVM2vJPuNTS7oCAliWJcXqheifb0YnVwkcCdV3lWlmaEB1prfTz75
1DzuF9v6bNPbeF0Nx84TDaBJ2qx/M4LlEDT0QWsgm5XKvBa3nouSYpejj2oHg49G
/zzOBomP+QnsQw/qk8ngyVOvpkKm2gf19DsxljyVDZA+ezLZa94pLlRZpXOG+pSL
Dg6c1gaIlcOpGsv6+KNhIZmZ4K3ol74PgScCuVvE/G+rDIU0iflawBB1fj9eibE0
5cRRXxGSL9lZhKhoTgB/cqgIB5GgR3NoBt1tnnp/MsubqYJS7UrH6yOEjZV27o9d
QOXHUXiehrzSeXxp1uOKoMBFQVHlIzRnudyBHISNjF+Rcpl+f6/1JA2KMnECoFpq
m8P19Ezhz4UUNhCwaBXHkl1eAyHXPZ6hxOwnblsByCjG4OEbzmWMumK/U6Zj20Cg
74iXlK4BoupyexRsOYQ3cKheZfJSBPqG7Rz/w9juyz3GiOiPakxkQ7zRiZEZZzWq
G/y5oiow+xEewkXi8KGZZkBVcY+W4YZ4y5rMnuu8Edtp1elk5Sf9wksOW1UgIQkD
O0WPIWj8detviqMf8LN1eJ2isb+248X9Hn5P1S7EvN3mZQoMRG5zrig0bQs8AZkR
yg6Yq/l8P/PCoFtHDt0lTMlk01aNTWmKPJqZlye/hg1Mvg1DTaeTZ/hEJCbhjy9Q
lFSicFxYm9lzBdwbfXZJWV32WdA7Ck05bbO5CM9LRNwV6/xo9VvbdkXg2irOdKcM
+m3eZg47+j6qFbEem1DufcWUF8l5FnOpdLNoEzA78nzJvKl/9E/6Y7HfIKhWv/DR
z5jDqLrdXwd7u2PuMttHpQjy+LcxSvKRQCQuvGNwjVqORsHR2/n64cbxV6f4I7Nk
pzW2k1L3ABGqZDfOyxTGxlCIrm3IeIL7jD8XmJ1CesKat9ENiMU80+li3iIBiBkn
3Kp5rcR5nRn/AXAYbgSAKfF7JHu5+k2c+JUIBXa+/iyZ1vfqrCVgNKR5Yi5SOokD
waiJ2myqxzNeWtlRUQlJnpWOfpm364jqVYR2Nlvvg1ZNNeHeQf4UF+TY5GoeOl4h
ltI+LvA2O74qkPzrebJbfhI4avEkKJUysI2yNfC6NUXkisitvtW3is+tyP+zsN6G
PZo48ug8wiTw9rq1V39aZ2BFC33Howdo7RyO1OHVehGPi+go/MJXVzY0IyFEaT1y
7lgqm0lJa/MaaPJAwbhUUvey48z+TInjen4cind+NdNNGRf61Cw0EBKli8BfjLv2
C8le8RYSEMRM9ifDS40afKQcsw3Eexhuyd+8cmoFh03K4ZqVQwcNd4l73GLH734i
1fSZRoHf7BIrBTF9bofjjJLQBQm52yM+foHurx0cA/S+ZQMv2pCFr6qUpr1M0qpx
tbIehFDO06DgQ+4+AqYHJdErnjL13o3NYsbTjCanNcINGji8ml2qpXYsBwiwR6FB
gfKMZx7tUmkqyVXi7T7D+TSJrO/+Koi09ll0Qg79u80T72b6vx2pJKtSCq3tgiF1
Ho6NyxQb22XB9k9AqT3qPNoHOEUrqNQ8o583rqiG2t2NngtM+qrt7WP7InZvlHh5
vPlMhFGq6/hAT3RQ4FAZuA4Rd3rKu48OWZp6a5p0XiAkLJrOM4ImrNcYDEVEzESv
fye3NBfaTkEzenjpnvON95gtQwAVCi15YGQJ3Jif9MEoJiG4is/QPqsy4BLcHSdz
VlDikaJd9HKDkwstJI3BoNsTjjUHiNWzUhHaB1t3LaxxJ+JuV3/Cpa6EooFED0HA
yhysMhmtxXBZudRGdpruf+2RIlXKTXR7FEAJxDm2LGBslKTrM5W1xxNJwBgPUlgW
85tGNjNW84KXEZkJYr47RzpFtotsrH93ozHudZ1TfGGywAsqsmQ1EfNajhT9dgDu
NH/9b4PSbygtCTgkK3jqsDkEhisYve7Lx/Xa5g8IJPXxKTsuJsiN0Oj0B3hFLyN1
q1sBeL5MhF+vWCHqn2k2CPlKxfQaUzGbRghPHRx2CxexkvHY4nmk2vkIPsgyjWxN
oENePk3lQgsISHg5bbGh+WCjmeiL7GCXpzbx6ZZGkureLrUJlDN1rmp6beZPisKP
dqzg4L2GJpugDAN9dxuKQNhpCsjx4AX9+tKNsfybGAiGHVrkp2OhMm9JG6aEg2aP
FzOfqWT61A4aslNGQ+nYAROuWD7X2dBXOG1sZBp0/CImgeJDJ4fzt5X2xhknF9d+
ptEJIVZiOFdR9EVrrmu6EKFynCwM3sXVmqk/QW7LCeCJpX0vzTezz8PQEzVv6btq
gP4DeQdTcdq5PUUupoYAtlfKKa2tnprGys04RtJCh9+RpM0gOZ94PajfJl2Nsyxb
yE5x1KIu9RL3DfcItWFKsff2MS5rjS/jB38VTcTV36KeMyliO4BJaoT97Izw0vqx
Vp2IjX1bsWf1WUt2Pp4F0zjWIAUKnkqnh2lu2z5MainvoPDIDWfJpwjLufujSD1s
S6j8uiUg49TQcnN+RLq8hXTkbtzzgqogC4XhZuSYJBncttccYrdoS8xiY2vjhG/d
W90td3cq81kc7KQSWsaawB5PqHAQltCYQNAMdbMjPR1vHPWCi+unFwFOuQ8jiErN
RNWl3ZfqfiXJMXEKXZQdLOY5zURjt7kJ47PQI9x/epfxmhQYG8cTL9St0q2Lsjtx
TTHtw9EvU2QgRJoJgzNR64CYpahG/JI87hm1z9I0LyTw/vPo8zC5vVU42xAl1QSl
AXIE+mCPfwltn4rVtsiYT+qSyFrlDZa2Ese2o0j3aztTL/R+4838xIBBmHxCxQs4
8hoVlUM1XDT3hSPmffqfrU+JA6SG3Oi2SO149CT8Vy6pfQgqNxL5H+xuCu5wufQD
MYcaH17my/bH6mt01lWe4MEC2PcYqSb5eCTVznWQD3H+wVQmgIqfhFrLjL112YF3
SEuCFy+QTn7PctHlprA4swGUww2r6nOhaHrtTHdb+/v/Gg5NzdrQJUsM+1aoXzwN
9sZ/FkKy4u4rdvWSiK0c0eJu3bEE86k0u0k9A9tD5rFUyHbNhjr5waf4LRgvc23C
Uu0V4UYUDYQ6gu8YD8Jv+5S03lq2VlSc5lKR4zN7cKd44A/t7cZTWZzTSV7eJG77
j5FB94DLWbm7cd9CqhL0Y2dbI8zhfBg1XzHA8gCRjRIOpVHy4UcVO28A6nlgTSZP
HB+wsj4rBEfU/PZ7hTjnbF4ytbJIzK9DrLPub+PSJCT8IQuL66rIj1GGtFh7wzUg
7k+qrwH/I05eFeUNutVVw9D/eG2apK3Sw58bKu8j19JPvuXTHKBkGQLkgykM3baN
0s/xE8o0RqOBZ0yqG24EZqREuVV/a5xPAq6+Jg0ffhot6PR5K+SKI76lhWhl1y+s
AUIdLvovhWkqkhJGkZqQlMK9kzRjBBrdpUm4YNK3KPrmTDjd8KaWKPO6s80u8tbx
XGjWNFipAtUI2PcDM1IMgYZlJW4JBHtLKv0/sPn/aWFvnSH357GcvfP5VjbyX3IQ
Eii149VngfFqFg0/5wGn5A5u7Yj4h64AzLdCx4vTcVrlMB++v5cSqT7UdfDRAD09
oYmhIRkc1ekBObSwLUsXybJ2frBdhuWipAolwi9+0ZOI5+GlpH6lML0/5a200OV0
mLmUhvOThN2dm5YBsQxO71CsQ/etXRcUxwyrdS40wQj27anxJ3HIbvgOFd4Aa9Oe
VSurP3KOmwn9kM1v2PXXoV/KKRndxh/S3EBj/i86LXjqChOM3aqB/Z5di9wrlz9I
BEDZRohvHM3ckZSvd1C88PXRLF+o0L1lnfubEbIXuq3tfTRnNJcwYHbDGzKxFHoH
xVYPSL5mFXVsIrjDktlZ3ri8rrQSsbn4474fJaopM5OVu8nCd45CeET+l8HitiJG
bcCyR3WYpJTasvQMAbyW0mywoZxpm7IQEMYgd3mBvR5kR0tgyhG2QnmZJLtTIpxT
nGA0uOc8D+5n5f/kAjLMwXlaCql2EPQ5z6vBiS2/hx8BEQ4f7axCvZT2se2iT4Cb
3cjRUZShfbkC6vb8HDvW4z6hoiPHJz/FPQDvhHfi6Y5P2X6DwM2md+XgX4Qyw8gb
FO4NscJ5cDnj2RXvH5bo9FD5VQx/YuxQ+aw8o7rEMOMPIcbnsncvINitSNL04J/H
0tyTzBc3R39RuaQdPV057+whpZ//xW9lNiHhrwDJE4xFoCYouXPKm/savWRO3lp9
yzZuy27+4yqX2BKFzvE5cSWl4wrvkMsRSaAGTIveU5m0gpSF3WPosrGDWdyUypfA
rDz5ojP+VcWfVhDsTF1iFQAOJiyhr51VRXvHzMxJUDglCeGH831jpQyPTuUC8I1Q
m+Fxpj/gwSvBCbtonYWkvBrYEZRYzMelM1x7k79npjdrp3ORUYtvzMRHauiZ+/dp
EPl/G+v/2UOISe5Xk+VPNG4N8BB6A1y8KL8gaxQGcNQ/NlHOUnT5dAyIBOaiE1oh
3It6qsqeh94/AIwJVLR4s107lJgMDxhBh2e3san0SJM5HE5j2RvssoBT5kuSx/nO
yWMOWI1FVoAQKPN/Wd3CNNGieQYKoPNduPUGcHseQemmGDs8UW9Og35+7LWImAvE
EAjzFlaZrpKDPZeUZQCBu+ursfu28j7tG80pWZyj9LMu9wwr8xt/dbAetdT740cu
sr6HZzDgJ5qIbFwLOhySZTgGRMaXL0CtvAI+9NJMdRyV6e4lTdnWQCphrcZRv/QC
vvfHSNqL3Ua093B4IdgHUDUJhcMqqjBvfWc5xT6KFcMSA1halq1Uj7NG67KYhZ0R
YOOOEPVJwXnarTn87gkhII3yZu62vz4OkiDUm9xTdWa9ZGe8iDDV0vr4/jiS2WzO
u3alAA6FaP1vCBrYxwaogIdSZqoi++CRMuLn/pD/WYSOZOdo6iYo45k4Vk+jsuLW
ub1ZoBYOnRi8Cj2kGyW2cr6ck3NIb1y366inN7YL6Lc+FAhrGYQkLbj4WCUWf5Kn
pf4zQ4kG1z8B0BQQFdE7ZrIDROO0GydMTLbN93E72tacIw0voQV3W5s8DYRQ8nrL
dJwLcLvWK6SsFq9QR5Y6Io8zkwaBRzuzmnHyFMaRE+5eOySL7qOtmAVLfpI03muf
v1YcZ8ytwqZqyePO7oqFC8yGuHUUJm0+sHoeLp+zFdbeXTl0agRyOnqgJJQS2t4f
iRU1PFXJbMo4ZYDMjj1wriZS2543a9LwD0tEAv/t8X+FAYnb3T5GQS1TuZCaiPZu
Aecr25UTv8uRYpTO1TlJt8958nAlsm5rnuXwbfVmAerNugy93tGAY4IF5iEwfIfr
FvLe7VQTguSwsQQXX6OZvbZszZCG5/26JNw9ZivxOhl0IjE0a0HPlUGK7bynmWD+
FD2tW0EzBeubktj9LFNwu+fqefie9p1xUGlGI2T+dAYWvwZGZXhxzGm/u7oUwCbw
YIAIJ7+Di84e6MXK9/diSGiDHuSvHwRHSntZByLajcDcK20F/DrQf7qREgNdbUO2
pUiOaoihpog/UimktmJN2PnNuoCFODjp2N67sZYE11N7zGx6BW+dS+caqqYMA3/H
YCwNVbKC6XuEPnye524nbTm0d1MGrb8CtR1GR/JdbTRxkCeqhhEQptQFK29j7FED
djWX3u3rWCtq3xG+yOj27yam2v8OseoZFrOYfTt1UJux1EJ08EcIl+7jGhLHyCCk
oZ9hBaUKEr3TTyP+6VHHAovpR3K/ega0DzcfXpbkGVpVXciVkMtledSZrwpaLS6r
Y3fYnOKOV6Eu+g3peOvDDnYtMLZZnOvDD2VImwINRrgZElXxJT24TfWgRNqyrGPO
qH7YpkRqNUIO92nT2aasvO4TjwCq1L/d8e/5Lu5mQNo//b7vehmIz+d/A2n/7ECI
WuKczdts84oqaB5bkpSLBOrsTHQViJP7y9A4hy8M80/mJQPKuLaOeVuYhGEjw1xk
e1DbVKFBKJwRewZmTcCkpnz5429ZKEFoMIDqnY311UbmfHOiBC/sEtIU2C43g4Vw
zQ5Zzu2hXafzn6LJT6ZvPjpVDtyts+2tzbWEr1/AeB7Z/j4Yb58Gw+cyhc4BpBFv
PhU1ecKAHM2IHxfdMvj5ng5V3QtGZY4cJB8erUZzfYEAdcqdk1Z3A1DZ8ByFIZ/U
WkZ135N3EQYDTUzBN+vJmRwZ8ADdWV6DOqrkzmI0Ozzz4DUwgGi55MJGprCSdqOX
f2jlI93BVYrRFSiAZ89GhpQqOF+exxH9vL6OQWjy1nRNpDuyxCfRhm9OFogi0Xjy
pFHsAZxcSYDvytMoDrIQa0ltl+BwO33NkBAtXXCwqLDV0EOw3RoCns48x3nC2YkY
698fx748jKs2xcp5NmYmhEe4oVQYVOIjxIuLHWb7f6P0z7EcV3wIs9SSHGpWkC7i
mWT6oVkA/D1sTllzfkO1kuoD7u31plCUS5KQy9jofBD3yQ/bJTgLmWkuH+CZzyd2
qZkz0oZkhGCNCdlSAsOnYo4CvPac55Zb4HeWMUgJsPivWmID2FaRh4GYPLHpZKqV
fUz6m+F1G0FJjaytVbkactseMkpr49I7qEiYT1s3fWv5fV2tgi/B5wi9cPyvuwWd
HUUvcIssqcjFNFnhZ0BmqgbGaZuadyQLYZqS5jmRC9CCg0v8gb8xiBNsyesEfxPA
wx7wqvueNkwLjdiPGA/VbFsLsCfg09K5MDOVw2PI5S4jfoka/I6oJ/vM+QdRmYhJ
y/bEWHin9zKSRQwXfRCF4J4c5p233gTChB5tUUuQTd5V/0HwLp1zH+bawsYO8O9M
Xghx1GrTKs0+VkgvohzGva4pGU9aid1njJf+FTkipz80LGsbs3+zpivmbq+bSWoR
kxO7nI4TxCRVKS+7pi0eNrnSfvlK/3VkTKVsXSWX9W9CbqyA7oXaIJNH8L/WbXDQ
3usR5EnQU9yNEl9BvsuW7YHva6olzBXMU9f8UNxeUVE/RQ43t64Fk/3uHjNQWhQ/
t3sIQt0WMT5o0ORCN8kk6KJRg7KUuuKsas+FoR8CXjhpATJqezIRAFkCEfX4VJ7l
+gU1bLEKM5OOpbPEPgklDoihFJEwHIAn5WUtm6l4L4olWwjgFD8gKxVYVn22AVXn
HSL773WYDabNxQF9gv6YLmLEmSlZuN1qjmuXBR0mjJf33oRav3hQxK5hd4zRU7RY
9mwEfwKz11rt5XMZ1dFITJ21URPfPk0Yt9vZWt2g92qZox1DT54Nj+AWawNMG0Yy
KmOSJTfEKcFPTkWS3uWyYEybd4IDAdHtLDCfayPRKFA9oycc0ewp5SutfrW9Etp5
RJLZumx9zfjzO5TXtQtYZErVXMxNp8NHmTXnLH8DNBEwEPhi43TbFvF1X1NTPJ7y
3bVZPkudZMv+uu3cMok9rZ49ZqqLqwBFqSBWaYorm4cJQS8QFGqCFWewSXNMaK3l
CpRz48B1NqZl16xdZdDDTkd9q9xkmFxf8/2SrPjaJj7/+rD5mJUnwExt1atxxHSs
8DftlP4Z34xbjP5FGPrrPOR1+l5dx83jAMGVK3WJe08GzEfEHs6Nj5isem4+vKCA
lopUOYRejWwCY/qbY8frFLGbodlsgduQ7ODWpqx4T9BrvKG2IjPl/luuuVs9vLHy
EZ3BiudWNF4QhMsTXcQrQeu6tAO9/wsnVvEuyRpnJr+T2f6q0osSRkDI0BdmWmBw
Tga9Ld+0loJqV9i96hnUPYJJR8huIwk6VDbVeQZqQUZnwnti7zyaZ8UG0ODFlJmg
QQJ7YGMKxlzSeyXn69yxcD/Wb6s+5Uqvk9tFsqomowKztZ+dEXQs5LdrnE6TQNz7
5nTfreMV3CzBSr5PvgeKH7FSaDajAIOUWaJCzIqSxbakHucvOAqvOG92uOQAUDPp
+I2rkw7a/ZrZUYer/MBWrc8oSNsT0q5Ml6blkAHrah4Nk3MmGRrbTJkhwxGMxsow
PYg2BPuXtAkRt1C2MIEDu6N21IfY7MPLPL0TphYoY7NISLQSZ8SzzJZRESEles2X
6TVQ1rx4nh8J79Nk5jr88wuQZe+Hk9/0tgtQd26KLh1ngyCWv2ZAlhYcRvIW7NqI
pcHfsiSOTdi7YMSIG546PfUDDDtVnuh33tH2jtVAnAHdNAN885uQsnUdYXhcHMgO
DUnhan337xMfQ7EUM/+vsSAM68IASacVWnM/WALZkuxtzrbVHFoZQmCr2llOjmt8
cB20IBRUsh1g5MKIVbs7QzjSry3aU7dMaBvrqYaiMdAOGqsW4lipKdufJu286gOS
suvoM92N1XaoAveuw7tWrIkUQSrFimbeZRKtq2ZQU9HT5YbZEVSut3AepJ5Z+eIv
I/U6O8y2wFVKxI3qdt11XKvSRrlqUL6FWbmYJYLIKrN/dGTAtCK9gC5NzWIXPKx/
01HzgD49Gd0PZjaRfzHaRnmnFFzLd/FbAwIqZzKDQ6MKqek8YmRbs9Xx8Ki6O3+b
foiiI3/5vmqozCZxw3Aq0TprXSD9t1xUY9ECVTP9eCHoaw3EJXft5vOGhN3+dLKj
PZTtsjHa+zKOO8LYd+o/BCFvBmCirNOnKh6pH5tw5vUFdlpCz9pbfsIoir01SfgA
N7vXMER2C5puNiGuocUwh+5FKA5lOF6oCPLaZPAMa/JRZ3R8KLsca3wENKnO//qW
eXlkgsdZDBREXPZbHREpmP9jkR1itxCR4MQHbEESgYatkH/fTqTbjpDeMc0rTryX
4Y9VklOMprr6YLi1x5XAgLwf8hQlOTF3213UYZ+qcT2tGtFePg11+Ay+mL/KNnGW
qoN7nKYx/4pdoNXDOsjedtAvAi6reo8cqHnBx+65Upm7uB9B/3G7zUnksxzyRVjN
n0pN6MU2qtbhn49hPXNsNjZwpfCo7DIswAZXzROYue6/RG0equw21sHmarebgbYQ
0ygYUCsIADvxNbHAmoAD+IAlJ4XLzaRRRrPDsgfsnogwLzLQY9+ufKOqOKoWzd8X
hxWGvU7XilYWpXBSOkAXTDor7HQc4JX9qEj6XcEcAvChK/WPNWcK3M+zM+ZELToJ
nyn/AkLtTchReZS5ZukcAH/5B/Cke6P9WmihSHFyiLKO9+d6YsW4pjP83ANi0qh8
PNWekKwGhL4XJOm9F3MsGhB5WjeAalOzxdUzar+A9thL4hLP/HFyHrBMSe3/XfrJ
m1BQ5jDT5dvrjKRp2iqQc+hZ3JyMcgBwpyAJ/XHByYfyhowH/3/k2yV2UvP1xNRN
IeAiCArhz1ZYv+OWtnxvCakuUJxBkeDFP4adk+YLJb+9u9gUoW81bQBgh0cZvVQT
p8n3alZv+2cEU13p5v3oaJPlKRDNS2QWWo68lSatD8cQBN77Qn4SEfbOBIkgZOqu
PrLM7/RDyFL7Fyaxx73GQv1lJ4Ry/kguHBt4OTZbzhwbtsDnrbhyuvyfyTKcjrWi
tS4hqkir8Pp21nqLPiQpuFdjWyrNM8MZU6TvAkP8LhdPTze0Zu3kvKFmvxviNOXJ
wpR6SV81vWRRhHT+6H4xC5m3+T+vjrX5SYYzvpEkl04fnvrRBa3KhThPS9R+lEgC
s4TevhqMChQFGbznVhngggPV721L3W2cJuEFHYmQ81ZkdC/A6nkgUA1COYl/HOn5
L5maGM28mTd/CSnNquoNOnQ/a/rcqU/ODpSA2UwMt6fnAoRNluBo9RAn83qim9KF
HKce8xm8U+TwTyrM6moxe6Ih0cR5d7H0dxwM2CnD3R2pkkRd1LXWTbQBEvhNdSw+
R90vD9VF5MQNk9l6F6nLJzz9KBbh5YHvxnVmHRYTNgtShM9Tz1SXZXe7D3pDkbay
FG3CsLoCqpe2uyyi8mwKWm3uyIDzJGlV4Vtp78xfx+17iQAnYL2fIatU2hcBYtu8
0yPXuhmupKyGcwLcrkfFbKpUwhXgJS3vFXfuPcLCfKDxktC7P54VWrNf2kdMro4U
Fo1H3Uf6/vRtIvfe1bAa7xGr43p4Xhwj5mZkGbiCg8ZGRxxClZ98R0sQ/7eElq+h
n8Opj0keDC0ZG2PJHoFL1YwH4DDZrq9tOh6qH3syw7pmYi57kHTriik1R8iP4Aq4
vrmK0bzX9RuAuwPNFnCuSW4uI6W3sOfOFWHKGvBtmWdZR7Ps7TPx62V6Ny1OCRGh
dhgljVbprJuURTHzTOYgKo75QivJ1VanFFycYBh949dOtWQs46WkT76f0UTqiVRf
MKfwEB9F8UEr0JMUI66F6Kb1o2fRCDWxWw8XTf4iRztDdS8PgTpEPhoF3ukmAT67
U6E49yzwRLv9eaqE2688icObJEZys9osMV72bAlisrLwSMZRxodR6giG+ykwzmM0
uvXp+uEMTwFKrkIBgUSTc5lM+wS4iFxFI+TFE8Imxceb3WdBU5EkNpsH5Juu0DrA
n2IvAJtELS33f4M1g5UMeBrGz1IVdc4L8VkAtc3b7G7QOxoS+Z/RT5biHzBVSaKC
5UFrptdKM5JFFKwd/vqenweABFr1QsfKgh5qOZPBHCM1hYYxO2fTJYR7O/dAQGV3
BllrCaS87y8qMd72789Y89/Odf7gi6bAtQQ45KqCWLbY9KVOrq8Uy3vah13f+bcs
EoLXb9qOcjWez43/tZAhnmxDFfoN6Y3rl8kU6dvYOLu6wcARv69A+y/OIQhIbCu2
k0FGk0O1cdN5cEK7ez1UUZNNqu0up5OjSawhtLI5ieWtm7KNSwFnxe2ZxaqT8W/V
iy7uHtQ1ieQnzUTs9mrWYIiZjAIdOAuxbO0kW2bvW+3XJkbdoA9giTixOkCfOzWA
IccoCeZok7Tnprv48S/AVlCSaSHPb1JMJNG+m9Sq2Y9embBRWARd4uBDh17Ghc19
YKcr8EDwYs+3u9NfoPklVHqkI3QSXH5JGdqT2uXhNY8kvSJcwH3aZ77s0CSpqTiH
nSQbMvVZI1si01ZqkArYjb8MQP5s1DH4kElXGSBKZr1fpayk2hJWoHPTIqA/iXCT
csNh6YVVMXw9vGlaKOV5fJ8ob9KU2RZRabt2V+FSJrTKb+IZww/9zEkT9QWJJVDs
ion4gvy/0mTtYYcD5iBLrv/Hwv9BPq6Xns/4WCv5AAJhjxHl3v7Kg1uilFPK4HXl
8HOzPedr3Iys4zp/k1aSfs39zsAX+A7IajSePfFf/OmoQd3yvv6Gx7OB94vW6jCq
2NSSPLyxvB6HGZ7zHJU3VyiOhRDb5cTveHlRPIqX+OXWl2kGU8M6jjAh/qKJe3Qc
WBL2oKNAKD6zOtEX/on3UHXKE2ucVzpySarOTngNi/S9OUcR98fWf9ObLoe3cOsJ
IrUFrJlwkHQP2mQQKgf5xdyYL48IxkE/8BXx+ZTZTSEQPhq+j8VzXBwRpMo2/SR2
qp5WqNLqhgHMVPBHD+/T5SbdT+G+KRVnL8Iul01yfVAQ/CZ8jFOoDkwmfiIOaxi6
ZAC9PnUguxdKSTS/bFW28F3I0DWvq0jVO/lEUaSGwL7ybZjbs5A/E4S8wYeaLaEe
Yuty7ZmqVj+Kbhkw0ryoO3wuT2c1jSzaVMbkUVpQhsWxrItmiVU+XNTgAOjYpMcM
KjWrzDC0WQhh7AtYJ1do73QTGFL0swuF5i9KsH7kGDpxmDkU1F7gQF/oxttRFDwX
TxQ+ZpzIfR9sN/8hZeV1Mp1ppJ/ol+Y917Zv+tfsYccs7o0ipWp5Zia0nQF/IYa3
P1X9dvTYaMbWuzSawi4kJmTPchLCJVa/iGS83XRSIRsXthwQIhwTPmo2EC5Q5CJc
LTO31GHESCQTqu3YE5PELd14ZB+cjLOPadLaVS5jhMsCCZnXv874LTAoO+ZH/MnD
nu0YNvrPHIvE73nkPkc7dmdb+0ixAmA6nqaQWeCSz2DGRCf1FHbCNnHllDAyolfZ
Q+e3ML/BqTtULvsSzmjWfxt8n2daJM61Br5fQIH3CTqIi+n/G4Z9qE0vDJ8RzaIT
zACLeiuUWLUUJWoirXSDjE12wU/XLVJCmFkm4+v1NzUaG8RpYMiE0ot6/bp95Evk
y7ycnUpbbtcXk1ZvtVchwhL5Y0YEdt1x0br3Dh4nrImwKErJWOUOWl9dPm79tufF
4cmg6n8OsM6dc3vJTDE19PwGCbcplfaXQ9rCW8TrjvKZ3SWqCzZXFc2HIreR38Pn
svENgW+9X9LvNo+Dp3oZyMBiojURDIVtgpTH+cVi1TAV38Qvf/X6okgyWQCNmH93
L9fVuIpzAZzJO1yKxo7uaStLwjHmIblDuXpmok2VwB4qgOuMH8HpIj3iOk1l9CQH
3bCCLOziG6NEzCepNcbn4B2C0xGR5Flvf3jdYqCz6dGhDFPPt8tD1CyxDr2szRmK
z+bg+b2iw1s3HXWAoX9jybQkapewXt1hxPawe+g5ZzC0zZers0psvb70b0PyKzlq
Sy8IacNtzjKSyOuLl7vC8speb4P8k8hLXyeEQVLGeeBZxluGyJ4GIFfYy8TJxT5Q
jxEF0pFXjFQu5YhDkTdTESO10IBBfMtbegx9K7tkCn46fRCTpN+dTueK1HJCSzeH
4f6X74QlWTDazus/OpTphCGo5lqFaIz0xzCCmtxs4PgnhYCnqua1nI9gTwY8tHqA
xrO6+9Ho4yDUzX1+Q+n6JjijvlDQQLicLb0sktTgHzYtBiUwsx/OTj1C/jONQ+8L
hUEqBLYZiMU0rsGwodWEANELZ4kFAzhg/CK4r0srYQfhVZZvxFahBGKG5CoyRkI+
qg5dOXzMgke234XKNK3brA5PfuWwP6+3g8O4aYG5q9EMreBOiiklVNBpsbqPEKBI
Onu4ENYiRKkz6U8ME3z+OE/eDQfbS9H3egizo6bQ+gYqurgcFcsky72/aAT9ObVF
5NX4BD5dwNQ1Rqi3FgbugsfICMfD4ya/rq2KlCO1P8US0iu4XH3gTfOuBRot8wG6
xwLpYMN6M9EXLsDhkA8SHc+UkESK27pIEULdZf6IfyYTK8PtHLBSwLT//bmmPRo+
Fi1gwKoYtiTziPOk1zjZVPY9vOcIbDvALPePZk+qoLrV13blzpWFZQi4B1+wK0ry
eecTXqkLJ0RjPjMkbgmHKSMYeiI+JF5sO9a/Q5O9pBlq6rwdaOVN+haVfZsFRK0A
ofFQ9Wtwme8ukQqYnymjhmJa9GVjlU5Ukc/ZKHkRGeFgQCbYOei02P9objoUlBG8
+/m24xfUlvRatgFi1ayEJ4kAt5UjOOmR/JSSZtYEcIbAPFdtf2cZER2ZH68CJMZq
T1mbKjH4GKMU8TKDK3Eff/SYyNthmKlZWLfz5CycVtAo5WOUJmaJ7wDbhdvdq7Ro
ZYazgcRl14vSyU9PDfGo5QBYWUxM3CxoqoxIjdfx1D1Uknr39HYyFgWmbxcMt47Z
hPI58+8GmyxvtQQpYj1s/QHBJfhSlvu1fDPgA63HOHWUHrcVsKAizVJj2nfMuIIu
59J/H9vcC0++9TkNikKSpXGMN7N7WiCZdVnlSuGrlPH7jfhl3n3a8u6lDhctA8s9
jOFdkwpo+D0JyM1YAp58ejRcVkgFNiqOHOYgS4boJ8+T19AwIhfS6POtcJeKmmYd
7fx79zf0h4znbGsvUcT5RNKR9CuJHraeQEBT6Nl4u3HvoeRES6IARKBXPE8nEqFY
JiregWh+EGEmDUK6rz6fb6hKLel68/VzqXaMbLH0YlLvUiRjaZtuNnsrFVCVvAuX
eQVNXQi+dehtlvPHoNnrWLyy8CdhMEuOl2zsAGoECmLZDlZcDPRjSyFxPtFl1PUF
g+4cUwkSAuc850fzodV99ZQzUhCudEX4zopTQRkF96zajzfqc1dnK+0HvNSz+QWJ
nIo2/J0gA8zdYmrVTNlsZzQRyvbMnBtYfWVP/AoE1P3Xafrd0op4nW43mAeWQ7qa
MZGRsZdq/9N1qvKzOhQI8rbrFu6yUej/mumbBNw6cgJOOdDffmMsTSMCZGm6GCVR
IlyqTrmGUBSuMEmxTcWSHutC5KVPErBzVzHL7ot5xYG/7m9qU6kvjCKeW/Ctx0dQ
uFwpl8vYJwVAUdrl5U8GUe6Sqy87kNcYMcgC9xM8baZcAy3DezZUcVhZy0iOovJm
UHf0oiBjmkFlzJQTcP9UQq+d715LJJ3sMaWMfyGTQywFcLAg8ArkMcAtNGz4PgRq
WkW3ljlb7R96AMIAKsC8d3kmw0HM3rY7ZXnaNfJoUtKelSRL6L6hHR8QNIMDRZqA
x34xe0UDHxpxtLc0spKF/vvdYCT0STh622hDEjk4g99ttUZX+QKKKx3JlDS57J1H
QwZ5gLhkkOit1v03QYm8se9pOZVXa/YaRnQ+i8sOqG0J39eTey+8P8PGHURuqG5t
FqcWggyXXhtwTHCNKTp9T6P0Ukyu7bScQtZIgbdbeK6bR8/QMtzKuCvKaMasKLRA
kZS5WbBu3q7+7++YtqkbuHJEEedyVZVyqheuQIDRhh/9ByZx5FfarjcHo+AHyC7Q
gYlZ+zNw1bq+bzp4F1G88rvgsR1rsbiq3BaIOeh2I+QcOYy7Qd8snH3Dpqd06Qm4
9T8BPJhLMDA5OGWOE44y1fNvM/P6qq9rhzyJSRyTOiwyqcjSBkA4B3uySqK2/Dkr
RVYvpuGrQf14/+PHUaSvtCeyxspDqr8TvnjRXUZ+zGp8N5GFbCaZ9nbJnC8j0zXi
m3oQJruBYe6gly/hmel/ZwNPEtuBzI+hXiFe6qNPa1tpJzrPgeWt5tp5ezwflqIY
S434gycFm4oJZZZ6FVzWeLbXKNMQpgCx5vobT0E9M2XlhZ5LnJYm4Opj64KAFVwq
wH6Cm/xgZWJTHWTgT3x83Svmlmxwysy8jgxrBCIl5zp52WkeCDmzkoCNraqf+CTY
/QW80Flo5wTSe9bk42FXd1sWsuWK2PRzDXVBk3s0tAzc8ZA1R/D+FcKIzBl8M30e
UexKFR49xhNSuXVM1MP6CaqffksrNfGGRgYM/dl88M85pfJOcoHNp5lf7Tm7lvPN
3TpCWNJBPX4908PJ3WFEafhAdV6lvbd6viMXW32AJs7dp7mAp9mpEMx3+pYTxJyH
UmOV1xNcpwuymzzRSsxknlGbtWL+P6OZftn7+zmPIu9mj+Bf4bl70K60tQ0ZyPgH
aJlvJnucS1peilsEg+2K2XiCYzLHdU8AaGdb2zn8G64+x6q7BM/lR0Ip4hzj77Zu
cXDTB1uzm+2yp5cwQPLA7sDyZSWTmEdhPNndWZgwHSIcjKqysCq3nAhFRmYWP2nq
Gb+PFekpa3qN7Iu/o9mX+wHet6LKN/qowZpTL2NfPJdLIrIYDhsfkpyjMRvLqpAN
vCHc1fJVV8pUpFcFlgqyjlWw4NHwPN++tC/n03ojPe6zuwLvQpqKRJ+oElf3V+Fg
iWmvcAU11BBPPzv5hAQabu8iLnPklKG77ZRv+FGV1B++L7WvscD0fdlXmmyKZmO7
1j3wFdSiULXLOgnA4jjPLh0jZJb6xmd3Yo7x7LPbF0z5BQl82jZH3WmgyTg/4dZG
rtdVE1CUaTCaBQ9x5Wp3ZTK/CkEDAMDoGzSPHvWZPIbYe8wNQvoW9znvSOsQGc/w
2tKGhTYxVQEb2+uwvZ4m0ozqwvb1SZCvqfutqYTCFwowevxQNeJzEVrA5JOdQjoC
JHUoU27OhEfK1DBBepO0mjxBGyscb1ybzS8+0zns69SmwGNW7zpO2W7zNSjUjA/8
V3cGkZ/5SQhu88XnBUJqazQN55baEWljQbaSjpbWrGFH/17E+PUMCtGxGOAZBmIW
yPWxl7Jo+fBYxmUU04xEh2J9J8fCnHIfoI2A3jeM8TdkTWuXXC403gKvjVgn0B0V
oiZ1j7e9IaylgWlPR/20uTa1iZdTSZW6P8gfW/svKJRgM8gdJp7JsXjmSPgMYwOO
IcnFCU0jhib22z0iN56tDRXv3kAvJzzfCpcQOh58Kl/fleWJG4Y6b8OTiaUAubm0
uiLWXEEnODejap1Dss8d7gYAFysIJaL6oFvVE47CiuA++v4zL39yIkP0bKgVQdDx
8tdPb4Ya4cg7jOWsz9FWy4kq8QDgbR8uf9CGd0XmtfTFUO3H02HnyMMRgfxz2fDn
gUcZq3j7NhK1QITl8ZFrzv9PziMGeIc568O78DRBAgXE5M9ymF7mKVMoiK52JMvD
itPx/ydweSGTGVp2cKonSUkTHfONFgTSrgNoB4xgfxhO3eR3O/PLRRDPoaQW8ZAx
R9K77yzmjDcccMc/n8fx1P7gJD/4Jcfvirwys8phC+Jb//1jSU5loQjY0Y6FRpPL
+gpMZAlgaKvzoHuqYMglXNTmLduGgLgw6gHM5+x8JNF9LFZls8cXYBcWSAN6Z/tN
KFs0BFcZO+JrfvWIY2nwSBJHZevl8rQcdgLNNK7WpkIGo1VUwYksbLWy2I+0Uvlm
OOiOlK6wd215piJ0GYcPMzW0sXQxDbXJbDMttE8cs2sQSGhVGo+BzRU1yq+zkvat
sX9obJ25w3NlnCJmp/bkNictToVYR+ULv2NDPwMv/QQ1hDj4gVu9bRkwA781phOP
54s8QwT8fwS/G9gQXMZAX9cr0aMnyY/96sjHmrT9pqYnkxlAIc05AFR7j43Cj5xh
sF6okBkxjgPH6fr/8BIgIwrhZT1aSKaSP1qIXP0kRblhGsbBLqzba1r8QSLN6sln
M2W073PzjWIHJ0b3/u3Wm9uvmAs3Nu1p/YSmjxccj4Wvq78Y1C+uElQhjMSZBA1R
uXqRJqhAAm5DdlMFNBBH7ILbciep7FhXbBQv0Xx8xfaIMD9qs0iWbBNveOC14Wof
QF/eJIEMME/gWjhDi7vhu0rZr+mBlOm82jqDp97cJAul8JgVDFgbmDeym065Nw5p
si1SpLE2baeMJlqm7s+6nSkaH3Qhcb1bR7R6MRes8fiin/lVtBQVg1EGNaQJoo5Y
nkh5xgFlsdGl+OuTqtD2XsXdY5SIsaV5+XIb8F92mgkL3M9j/Ee4yM1zyseXt/va
tJ07rayXUvDmvkz+SkphNBLZWQ+SV3Kf60kQ+HefmTXvLZP1/KhszXws5L8LH7/O
GdlixJesk0b4gCDq3+y19ITEbLy7Gloyk4sJuxde5WgnrSjORsvbEQhKeESgfYPZ
y56vzYMeMlQMZUGTYy8nmPjszVkb3uxHBPTVf3FHz+yA37di6driXW0HzmZrQRuu
wk8rlrJKQgxUyO6YiJFDaOgj9vttzvsXC9NnV3vZpryeIt4QW/30LQC9dV5nH3k6
qClkP8r+CltXmYkO4DVgWHh6KrFtKdGNftyJjPvX4WafaoxhJKzYU2SGCN7gDaTl
NWP3tVs6wIB7uy1uJXFEHsuMr4qa0wbZiq3Oe3XHXJ6ICDLPwT9aj4v8xTZlcK4C
91IwPF2R6Drs1MBjv/+SrTi4rwxx96/7/gtXP2V7fCrqaorWrZg/HOx15xo9Stfu
qJ4YML2nM/EJHhNSceeI6FKVSQ3ySOnIrzSBiiOFNiqXMhke/Nj8AvIP1whda1mt
ltYNupvTKuuQtbOpLcanAeLwW6WZvE21DtffRK6ytQhLJaeAJ5U8NJxt5qcuT9Km
IMm5jep6JiFmhn5FafGYJWCt/KlnKq/a3GZu3tV9ZJpBBKHlSnZPvzHSWORYuhGz
OfQ6GjY1oSyRkzYz07A+kmLJdbj016920E9R6iGCNaGnKUukTWngWudsV8VJoLbq
k5hjbesevUWvfiqlTXVLZbxQjYFDDo6kG2v0byVjBzN0WW7M/ANPqD8rfdFb9nFo
EzBnF5zRVQdF/W22ZoZKYIEMA1+yDqnHonNb0TOnmFuygWl8x5ZTjGCjXfJK1tg3
iTv47ogItcrLclnGVh/iitOFUdyblyF2v9jdbgCE2X3sBlZ6H/Xsr8uCaNpEJQNF
sHJmeCa20WMsrraaQzUCLWWwr7aRx7lFhBF805lDqE1+G2bk/vQYT/mdrKCQUMqZ
/lsR3DxqhGPeMtzt2rmFw3NafyqyxO9Zn61ZjKqHGWsMxYFD+nJc+AWLbCYRjnqs
SZC1asnB7lMGwXAI8viJii70MfC0BCq0OeCHWBpHwPqmkgvbBCOHaWFqUkorg0Q7
X2yWLLpMHwPIv4AuB0qNfS6ayXiqpI62sGrH3wdl3XQQ/FNI9X2NVlezkDKv5xcq
V7V4He+2szmaV5n9A/jl1wMT0X+fiif1LK8+VWXxc3YRhfI4VYdrIDnAOGlcOLJu
pnGtK0VokEkKTCg2G4vUQdibN/tC8d7T3l2U9T3KdQnpy9AyHNLdkPjzyz0JRZSw
DvBy/pd+jtRi3RImtbR8IDlbvCi0BCbNnGlPmhEc5rz8c0Cwyl7zZH8vhp7MS3yF
d2aItAO/WzavR0iZktaeDFYK9enHxPtw23x3a+DXpYzk0fhsMhV9CLGkYJHf43Ih
jjB428Zy6P1ocYrJgmYqBzFGSmPcXHQlBDj/sU4V60kRuTIftQETELr+GVOW31rG
uU0A7njoy6h+Q00vDxvX+ybdPP6YxbQBn8Qii7CB/h2CoOVau0hXuYohAVLIXi+Y
GVIt607C+hMEppqVBWBSriXnqox6DfwgOTLXaqyz1hkQTCGCy6cr/ds7Arb0jhqP
xgrHT7WdOpTAGV7QcaUfw4tkVtNNpSUCbL2i4FtuhSw3ZKWrqTcIhAsE8EDchx3h
3bgEi7cgriRj6ibQ27H2pr5lFiC5i+nsB4jU8IDOT2R4ADMpGfW12iRug/UjB26m
+y6HZ4nLRED08d+fiBLWBODCqcHDDdXStVm/kJXKzp0MfvwJ6IfaI4fToZQVB5aW
TG9iIJHKiXzzbo3gBRgGfx+Nx5jV7+ktxGiNSjus1d/wmVVS0rhl4d50AQPPDW7A
2tDO58o2VfBPyooBBUjrv5ZcohOAyKLu6AlxZpZlTrzWn0eLIOunE60pNijID5rh
gNA0yQYM0HzboYNkSz2x1hb76i9u+q4KykdpiDb/xNjeD/p2hyp5cNys56j3f3OM
lO4JDLCEQMzqtiZYN7DKIh96gg5C3xZ1A6fu6ucVZ4+Rt5ELp8+3L8YeG/1imYEL
iFzbRGYU+NBd5eMdCcGPesB6bv8yAt54mR5THhtpC5UGL0kjV1QIPDENHuKE2BHu
HmJtsAiE6ukqPuOuHM3ZBGy1YOZLx25XiFNUl4w0qx1l+EAyCN1of1Tfpo8J+cnc
Ld7b9DkXv5GxAhcH2wwFT12V+57YHyNSE0tW5vmcyk60F8JTu0TGPUGds+tOJCgg
XL07ws/6aSrBbwzJ3AHQNOq7UfJCgqsPcNeWXcaZ0DfJD1BtV3oRoBciQVL8Q+7a
BPo94yRXQKbuCOudoSmpbjpE7P5m5iFnE3ZHSSeLBBhH0ghqm8T9nMNjWeWFfKPv
nP4y2v++mk3n+ua6nfxEAHhbt+3if3IB1pq7AYAE+Jt5SWtigxMp39KaYqdoX5qJ
3APYcEIiTXuViPDj3WJ2d4B1W9480Db+e6HjMCVEao9jooGW9BwBQ2ycJLfjGXwA
gAJzkTLWCeMdFO+zcWnAfFzjE7jdAFOUraGj78utzjUJhWfDo8EFh//tXD2fVbsn
1GHNCvp117cuz2xTzWZ3cSTgrT7D40sjux8N7EehtTRE0hrWu+VJBEchbgzOYh2b
sR91dX0lsIooKrPeQYybfaufEmBRCPW2uMlfXc0roLSjoT86ffhQ4KIRydpGl0sh
9BMK98qVTtEw11G1ya9roRmU2NoqW/s088rV7uBRbqnoVcXjYCccNT+WuwWtQKfm
soScWHN1O51PUWzgv93OVNcOMCOpWvX3Vuv9cTDhdgXvOaw1RIET8esg9EnYDsCb
J0KOB7JB6Fh5LsDmoeT/+X1RieKFCSIUoDC4D3FBFRw78ZXUQQUMZPPOoGX/3Tnt
fVKZQuNoMz4hmbPWPtTFyphJjobFj62Soiy8kgM0eBA6GKQq42nqjMkfYstIDZuQ
VtG0+SCJFGgLGzlSGgZO7PI5t+QCXsyDZwX63ptcvZlVvpkPn87Oanyr7u1vnG5v
HX+b/oELXjKPqZ5YdTtLMNf7WADw2YHIrTYV5Tfs+THOimkGUs6usC/TmmZaXIxm
EmTZyLj5a4zt81ZYimClxx3vh8Iu64cK8Hgbb1RkoFugZ5svJetus8nQaoyY+GYI
GUSfrDsi30htTvdfkg5Y3IRyRTRnWVHuHSuk6ZvxW3I9qSJ9OXI/M8kwT6hy7pnL
RA3tisiBwqkzsJoiM+09LBFSjTGofLogDQqsXx6SBSoNBxwrZw4fX5n2ojnVMZhi
O+ioBjGroKKTC+DqgP8jVVnr26UTWjbkF1tKuGlLjmwwuS7PsjtblIzvwnWxP0Fq
RNP12xQWTYXYSjUtwvtezhISFiP+MQMsirEb8jOrkiwszRcH9zGGAfyBrkybASEz
YQf1n8/cbD0BWU94A8IWFloDKsHSzsKPWXdpvSL6zbTAcNhJ4oiR2deGeDaYKFgg
iGNAKJBtsFe2gpCueZ3VCVHHa7GnGzYcm4QwmsOixznC4PkGVEXZTaKpJp626fTy
qBz3sd+dazgqEoJdqcbqMoW1ZByJ2oE+ewD8B/5nbirrftKGkIC5F7h+Zcaql1Ar
n46ofg5zeDuGwKDaBagP5pg13BktNAM+At1/dQD/QqI8Fb+8tMA10l1tHeTiaB8z
OR7sgcGHuM3fVpPNYLdpmaRCOM+u2daezOoxN/MgcjWxx075xy+imjpxVuNjXvFv
BlISZ5o4BbeZOP0nEu9xPGSK64HzjSEegDK0wlQUyTKM6MUwH8dD/quoBQgstrDR
lqJOpXkCpquSlalrAQfYCp0Mh1ObW5K9VvLD/77XMVg2wVcZ33St0Q3EmrHt8iAQ
AqelYVJ4kVq6qwvG4Ne97jfFZWEnE2VuuvqDiUR/DKUvbzTzfyJgEL0XkwzPqm3n
xiVqrW+yrNaw8Uf7VRSsCyrBwdgPvFR7dFKhVGyVTpFWIxIwzJIyE7GB2Hjg9nRe
FUMjLdNC6FtfJqaSx5x1mmMvGk5HRtJmw5ouP14d4AibMbjdVqJ+E8yVYS/SNfck
zXgxJRmVNhuLS4Hc/noEun0lM5RMFYGmz0AEuHqBOz2q6Gyj0E1hUTj7e8DsRTjy
nF37NaY/VPKHphilsVfpOkj/nuLoyvQL14zZH2dtW8ksxH1/P3fq094CgHBlOwbO
9lpbAzzFNKwbspX8O6LPBvDV1BHLRofYd4L7QqHW9mR7tg6gYS9pmEqhCZGJfr6Z
9VFumRx08S8Bwmx2YQ6mVxmDy2QlgsIHY0faqpaAib5wy2hz1uBCxVHDXUUOqcFd
OORCnJ7UioWgZO7vvguZUwf8EXWfeEPaz3m2BS4UJ6Ho8tETqGsAy7kN44oMkQPh
o/XWCMfj8EchMGnEFFxNn5kjhWB6peDDF2KsVZA9nJWNNBTSOVcHfe9bsVNsuS5T
771ZzXwxU9AAkatLA51xtUx3xEXapHyR73xUV+htzYmlW/IuSqooj/detgsDFc2e
IXUa+2WguCl3RTic74/2RS3JLk7VaSfou7H6iGt4j6aKoaMu6uhN1zLqnBGEq44i
XVpi0abiECHZo/rIu5FXMPQSBkBUNhUQduVvj1JSf1E7mFCiubvQNnU0rMatRRKF
UWw6jcBXBcxPW2HVsHjt740gQrCSmYoWWpfwOKHRgFB5VyLogHIu6iv/PQ4MFOKA
MYDcn8qwzQrLyLitqasvG/akC0+EbURaHgApkiUW0ImVebbpLUrpOgfRwoVfXqKn
UGQeFNzfDyFFn/Ezv4lfKOoJdIyKNcPAb2VEpoGaoydhD6WNsCiB5vrQLtyokivw
cujsas3ozzdfoi8seFolUrnRFK5ZFEN1B0wGogZp8ceZDQNnszbsmKA5LU5hLsEA
WUwNIxuXkTvoP4yU914kiXO+XqGBu9ownbfWujCvWBTw7vb8y2UkE1Tj5YqGqg5+
RUYoECDpwGx/8vOkB1wdhP+NBYekwRwWF8g2pP82UPODMu3j7zDoEOJEW44D0B3K
okFsr1PZw+W/xju1gWbPS1WOuvGlt/5E0PAxCtL0rO+tij1Iq8SS8SR/AUnxwjil
uQVBNLhdgWE75CiJUWoMjK1/8ULs3ZcLrDYBrPlSwR+9Yd6zR8qsF33mqLlVss7F
mhZIY1J2b4kSmQtrAVkJ1wPP1M9VPaZxz4BJGywOL9Y7nneishW7pbx81o7rrFCg
ICeFrDAHUMc/5FcsBQNW+vqxBP2GRGBx6alQU1d0jrSmLqXPNUL3JmHKPwSotgDB
99cLX/4R6m/hMGwJ823Ashv9crZeaIfjl8yyKbA6ynYUE8aXSksdt02fmFgjehGL
tPUu9z72pg5ThxZh1CvPCMhE9Cbt6A9jy3EuTbRoWAI2tw5CJAt7IDevHXHCyAy0
tneuuUyqlyFq7oxAt3XcAEIFLNDCllLzhcT3r/QWn7SetLWip6mIqkkiuYdYFqfF
gXOmOX1IFObSjk9bRkDxDbi64TJETaCGCaYGfeNDdE6Q3Fij4YX+1flBDHUgfKuq
2oxO1MUmmmhUI8/Tt8c90vvdYhLT9T38yIZqv+fHz463FqQCjfQQM/OZdJhHPDCc
2L11EjKvJdjGnME++FzN//Q3j4KKgpcqERN0M3NMuwnY9I9ydquFmUVQXaQZEUmF
MMGRjRpLn5aq/V2l20g47R3WI6It53ZRIGomMoqZXeZ4aArW2YEE2ZSQIkkC1ZNU
MXr7kCdHsKGK5BO27aKYvZydMGloHzg4FHKqPHVL9KMuvuZaGobYBCjnlmbWw7pH
Eb2KniEOIpu3zoZWltJD+B+24C72gyWOG+OqvHIxayizDkXX5PPj005iFAxvEofp
f4j/UITQ2Eh85XlUtgNDuEs9bQ77MMzd1MjVfxYS2KVa2K1dixdaaKSEr2/xsHns
f53qPiYNJuqR88IhJuBkhUXh3U6U5NUweEvCCgALf1uluZR9Aa8b10hf5//btTN2
f+FUmCWQZjtYjFtwl3nKgh+rGv85NRCllFhlv/gAbK8mzfdxYOTt5UhPWfc1PWjD
rdXq1Y3j0mpAHveME6qV1QtGGQ3J/mMdxJspepY/LsfPhjA4ch84KLt+VZC5KFuS
tekjPaGXzy2Z/4nrTLpQCpzs+jiXvxH/WXJiCKq5Y808BYwmF2m3Bl9rWob6JcPY
uLXioOY9voCWusMDU03inEg9u2ZoMhKE4piwRsI0G3MxNdUK/K7hem3tt9xLGYL/
qawsKXLymem+0jL2JSwgB/C55+EW91sCByCeItyN2tjfu2QbK/jk9879lYCvsNnO
UD6a2EcxvGN6e4yFq3Kd/Pzfg3xN2yFtRkMVcGQUwqF5tW2RTY7QgrI/F5vPbWpg
e+n9+m1ZeQ7OjGNZ4qsZLi/+UedfHWTm/EWL3jM5Xnb2MLuJ4zX542t6exUMPgW7
nPaev8aLSfKluH2b9V0N++s28YfLLfs7GSA2pe/0ZJzi7DQ9f8bJce+yV0BUJGOF
NS8DVMiCXUUc7YIRvt/q15zFtRXmA+ttkDelSpA9E+jJmfTA+2xLwSdC5wJ3EuSB
NJqaIqSUH0VPTSNOt6UK9rCWfwxiGMHHE4j7ZndNviMZfmDAkoKtvwIU4o81taE8
B7JNHRvl9NH/yjStyYoCMvuHyc0Q6E4sxDkRyNhoM7h4iXf+Ce7TLUoyRdl2aH5C
vYllHv+1+cWe8TAqx+x9+JP1Fw5g5yHxapDQ2ToiWsa4bk3qlW4Pdt3h0/0KJCOi
odNS4aKD/xL4pZUFg1tp0O+IP3Ap9NClmeQoZ4IwjgVd9k9Bpt48Y8m4EDbGXbdx
6zSQ+5yBUOzTY7C0W+KH/YfXrUtsTJNhAva9bFTYZ313vi7pbZyDSlJX/IWuLEIy
5vWWRsDIO8qfa5S13xkNFHtG86ec1cekfehSwnRhTp/Taz8UdQyuwQTN9BG57CDD
AsZ5yhyss/laEjkVJiv4uBq+/hZW2GrpeS7qxn/Z7E7C27tyaAhYa6d1VhAtVknq
6o2xdqVt7hVps98CHHD1wMPflgChhtjBA4UNY+HfLveayInLX2mTv6Cp31fjOGLT
dUoSop/lsz7eNEQaImhpIiGBpuYrPRVPFeFFyNYuWixE6O2Db8Z3Y/FI5DLL2t9r
h+Q1c5XIH7EYmzOLN1t/OvRLpzELxHw8rcaLgKw+k54NTMw02K5Rc4QZfFKm2ulp
6t3bHY3A5MU6HtElmuNlRzEbVuRotRqOy4xtRoZl/1o7Uz6T1Xz1Ni2PdAnAoWBv
q0bdRp+HdltBx1kWZvvOfJzW9BljkDItRU4W4L5KJTUDIe87R3QQZ/HU9/RqbxPc
fZeftBunZg/VvIYuw2PxkCP3sGdb+TRDv0SZXybqr3ROzZqwkIUOP6hXOppv9cuA
T2jAwfzdgLMjQImQejhoUNOm2Ox0YfYjE412OQx30yjG+qxT/F3p4Dc9cUpG5fj1
MHgXafttdxLcseI2hszcncNGJL5LvQU9qEHp/CglCc5jPbEFEpK0i4R3BA/0WAlf
5plBK5w3nUCvzSC8GSNte1pSegnv2dllR7T/MhTTJXx/6HXanLGVfZjIvLW/dIGr
jdmmVJ/dbQOC59ZpDmjMkF/+7XNnU6bzCa4ItmG9VHEwLEhKScAwP4XAqZp/hgrD
FlueMOfIMCmZEBERbv6+4Co5z4KVC8rlVszggnPlCYmqe2b3LRfApwhDvOnwAi1T
taIw4Q02erknAZLI3xImF6xEH1cQtRzPnOEGUgLjFG79PmOeKOJVy4iRdKTOcYtw
0SxYu4rOyJP+R67Q/Ew3LKZI3taGlFSsE9BqqmeqjguHJn5o6/jGsA9jJ2ftaUiQ
rfNBEbZK4llWOJxO4kttt+ADUgRIaeeWgAeJNGb0escjwqUDCOHQd0Z+7qH4Y8ex
I8t4pjE1pSZykiLqAz3fekheEqisl/qoGJfFplwec2oZFMWuxzfqpg0oxf6MM/bP
li2qNh/Fqrp0na//q9HQbIJ8qQddpkBTNSHpjh1R7MfvAjG9NghndPlQ00xRpBhi
xZChAgzBfLtpmWjx3VCMgSopOUvHVasTvvoSg8Ci0Bf+tGqMqTlTk7zHl6/5/LIH
6kSCNHNd1CFIGoAzWwyM4+mLLCTAQhJOJEFhFQe48xaWrpdliovyZpH3idMkXcTA
lxsqhz15tdnm2aYo2PsZKysE0UziB5i8tBHqJNPCfNk3YVnr74LmXHYsaePQ62Um
L2q0+5VpaOoyrManK7/CYVDYl+sJigDZIkB9ncdb6kikhkls4lEyAmb82YAlF5pW
K01SIHiVn44XJGUBulQUYZzY9jL+0Sp+ra7cCuWArR5zCx+hjaX4iQikvZEmJyQa
xx/sdnbp4YkcQIKzP9axHGJQj0dGViyGw7sCCQC3wsyvEOBUjpnWRq/r5zg/fold
AGbbIcv5UxnP3BLHrPctYU5K+HozaekEdkkF6Xds/DdghQGzUr/jiNZunkQ2/NYO
dz89GnQFh6ZVizMtXMrGBsVyQLpqqPrwFKUinHt1IKHIwTfQLeW00oIZtnfmHsf4
VHUj0Fyup1yA5+HV6lgF4Ueks2E72Q5tkFyoAP2a2tAjfI1CchFLTnfXaeYNP8ti
qswBNVMQ6RGl6cBoqPiRphK8/0ntHC9do+sw/HotIGWF42/YPR/W/dqEnzxjvqJg
cGuiDhTSPumPoiZUT6+7OLmDl69shNwEDs+EU70JroUCVV/f5jX5uLNzJf2VuXfB
2zAZ7Cp3hl3ynRI8/WRBrRVTXSn7x9ZyMxkC72JT57cZNSOMiZGR/fYhmxiIjR2H
/kOV05RUQazAyvmJ5Zrh93zmLXiUluLnGT/rWYUMHeTaI0Uo2ylI6vX7JMR2uRUm
DTyuNr+589PwgNp0gzL5WrslaxdASap/9ymtquDJTiNEKOAL989tun9vVQRvvFhl
KY5Nz2T5yOz4MbhuDeMtEvX+4vyj6WfubzhvB9r479Dx+40NQbc4OdBLQcK3PPjO
LKEaQYYjAKqlMBt7C8DxZaEkq8F8vj1tugf3ajrYXjPpw3ZgIV4tIEJmALEFjWJS
fC4EHy0vRDAj6fTNgcBDahQOW3VtoMy70+RBiWQrib15wIxzgivkaA3TufPE3svo
2BasvifspZhRFVAkljTj5M+wTugjkdTIwyo7SbAoUC64P4IA5PeGSNxYFsFHyYVv
7EywlDDIVgB149DAo7WB2ub7O6bldWXfh4fGtTEB1JZfs+EPqhc/znVCsOUVMO27
Vy/Ks1mFt4pXaiA4UkeB09LvKvYKPRPlV6X/qePCV8ttlZzIKP9rf9Xk1Xrqd3U4
C1C1YEAOzsrdR5oGoGyi/XxjDrEHP1Iv4+Ewiln2SVZ9FLLNA2BiehoHD4FppMVC
Xtn6nKFON8eIdsQjEHeq+UzcXnWGJsF/3C/8RFzqUsCgQkMgjST4xuSiu81FYhCh
AryypeiAm1+5NjBcVsX7FHV3+1UakwbRIvmTqqekiRNPTUWmmuIYQJ/JmOJa4JyB
vfKwOWHVWq8CMLriPdQdPeCqZJCIxqLhMLXnMkJnXVVxYUiVW6oO4d/VJDzB5f7e
ptTTPBUD2uy0ZglV0ASM69inez6QhnI5dAj5msYaQ9UEQE5RSQ3T3Rr9nQsxlzjW
248PkLukljHSXUTHSyD2C5J1lNgd1tr8g4jP3UX9w2e1pRBiNIBU0MqJYxfxHr03
zDefRBxQlsjYbFKttPUNkAA8tG6oE0Luz+R2op51Tpq/zG7JnLf8C3LasKvydb75
ayIsripHvkbSVW2sPM/SW+n2lnoL9j2lPNsWTuYeRQS17RF2i8JB9LDuk/TlbM/v
qdYRepRIBe0wZ89+ydYlamq0bFNpkPG887LxMT6bm7sPT360ymk+RromuRzdREsT
kYE75nyV/w+ur6QjRaH2n12zJ90rCAjQllFz3ZvlRGmXauOcQPk43hg/HCv0A3Fn
aaJ3Rcer9uDlMDM8fI+JX2rDLKbz1BKZo/Z1aVV8YGkhSapmL1Bxm297NE+I1Vfy
T9xJOfsLOjNljg/1MKJanmX8DCIQJts6XkEaDCT+vAeeP4Qx3C2gUfpAGRTHWk2H
IWFMryiYtBv6CPf0pAvYn9vRGJt3bJafBihpcI92NZKrkn6mXEmiufSQKufGIOMj
FKcCuUVxV1572cqCPPVkPCcEF2jq8uXPLVbanxqDMo+gBXkxq6Ce7mvpy1DVcMxV
xJccIhDsDH3u3v/0sJn1mpMtkPXtR5UB4a6IdJ1DTFbj1Q5ngtll9HcRkKQc0L4x
I0F0a9NPQDwXp1RYVWd/pbhQre274NYz/TWIn9dE1ESlg9Rdghl81cBiB+Y0/K73
48gLIlSlH3Go8w5QQwUDsXXfR3tmMik2k7aaq0A79IBSGE7siKwil9PvdU5McRXc
Cmplfv4cPe23y7eryYED7AShUhDiUSOexIV6RWt+xa3BRaN7xJiNZaUQfrQws3bD
PcMiSvrjthTRSjCwwqZcSfGklzjWAgtytOvDujKEvFzH9C3fs8YPvmxOyJPOocgi
xM6/LQe06LB+ZalIpuKtAfF5sIWeKAOfMvSTYc1Tp857dV3w5HetmdepLungOquA
criXzCfQDifEUyVJqPpF+qqXYvj5jx2ELc/dE7kRpYGZuV1CsUGs/K7V2pZj9eTw
ghZS33h0occNxzq5YoFM0o6TYKMZKG7mBSKHPZUEQvG4KdO/LYY1h/1iXg8AqTe4
FG6xV+740tXukJPXYnmnEnSA+VK6DVSSHkpsGYIxAbyLqWN360UvPAZ4/YI2TBK1
aNWY6cw0jRuYnnoUt2t3dmzfj4XTThEGZOJg7vZEyGcHAQxMhmTyKP7S92t/KQB0
aWFZ6bMkzJawI16+hhxWu9IBMljnaEVyztoD6kJrxrYYO2lt6R2HF83YSL0ydMKm
a82jL94kCfS8Szcdp2ssVOdLMVrsfi20t+VsQid8Z6MtyCAwec/Zlaoy7uqmk/O/
yhj1yH+vFKZ1fX3NRbAxBKHWgGW36H+AwVUjOQlSH53R5JKTIjZG5NEpDTNiEQnT
rGtAvbhKm34Buik93o3KXuTJh8iYodBEeacgij24H1CNzyiNclUpAvhZ4z0jN5uo
mW7/EOLY+oUz9HSNjzCZHVk2zJsjLIp7D8Q4J37busSV3HqqeXuCwY7e8VUCdbiM
a6hmsOwhy959864kL5tDzIqngQ2PC8PCMwKy9iDW/g2ckQTABRA/uAANoFfpLodV
kg5M80kxY7TXwD0r4olnJDHXX9hIdCiDvwrG3Ef0L9VbQREj3Dejqwo6AOpVmJxs
4VxOYO9fVIoEAdyEZw4CzOfx34LJP6sEmpMkzTpXPT2MNWm+a2NVQyCQ74PKFBDK
k3jpw/dGRzMb1cHMInoLbiWahb3mUHitKw9EiN2PCqZMUjblLgjFzk0cCF4OGIoL
70tML1wtOhOzrgjrGZZ9vhyyYSHSp3McXf4flmgNa7BGjYpqEmtSOiZBQEVc9K/e
usunmWTIOSUBMw6DC0kw0DQ9XdvE9X2/6YWQS9qMPRVNFItTqpv7Yhf17Li2reEw
UOg/YxLcSn/keCeHZdpzEjCJFqwY3AgkVzAGzP36oWVFRDXBGIhsNAy37Mty7ES6
T0nyJnTDj8l3ZvNbCykKryjPtyu67jnzYBLvKqAg4GttqyDpIhbjdWkAW4Pl4P2g
Q3ThvouBimklwE0WU6xXunwIPiTalx8Aorqsv4l+aqQLBXLZ4mXgSK+z7gnot5Ct
ENpfkJR5cd68CXOWr6/qt9E4b0uVBqjEr/sylOP2Q+eXTshcrEOFt2Z3oCzmzgiS
g0Z1HMn9TB4N3eqYaywHPBztut/zzfArKKKq6JhU7CHRiJvSjZVfB0/H++/qqGJ+
lh8yyD4i8/LfHAYpkOfxBR/bi/v5OQ95D1xmOHoxegbEJaSO7L3hxiFX4LvFeusP
wW9bqJrzsLmNynHRi5IgSxeYA5ZIOlxPYh8U1KvUTWo7EsSuHqBaLEGLRae/r1QU
X3Ew0o/NGV3o9xgSvEJuH5dlR/bPbPmlCbU6GS/mhx7Rvsgp/bavUyPIUqagsLNm
5Gk106/ZzMwVGj1q2UJyRohKr1Z+l9aFYLBMnjaNgTSrm0UkvYk6AQvB/+PmHRWF
aaPKuSi7nY4bqxKYd5nUwNHpBghY/E9M4UoiTYjsdkjhckGSZ4hw0Z/bEYWNFiwf
LOq2IJxX5cS9JfRqeyISXltqsyWoGDGZA0H6q1oh5NL0OSNZKW/yJoW+2eYobDcT
AcIOfwaqCGQrImWzlSOVW/a1VFye0NmvG9la4CXmciQL2X9YUHBWRBupL7Hq+haD
3aEMijWaOaH5E7EVlEQWmAbcEXotJ/nzbFXCs0mLoKnNIAkW/rVvQR50ot1hIfmM
zg86Kx5bMlIU58EUsH5ycyoCaKIO8DZScXX8VpL3ItQD6AYCL3+kcq0sPV9O73WZ
plICwAxMVhA2Ix35ZNReiFaLmQMy4n6BXOPtOaluHXXpcLUSu3qnWQfLBToK24bd
2A84YcUaNBcFUIgJepIRpyJgVO3UytnE37BDbXu3le29IWAPjni0BjiyvaP0IYk8
Qz7dYmQ/2L+cicOynmLi9HKHuG4fAyd27VOcdloIKK0w+iFfeE4WXQp/nBA4S847
c5yC+aczq+aiBtwv7ntgiTY+Ikdm3HSBsGY6QUfoc5VpSibtq5cd/WIWtAIAONFW
jmNIY2aeFoeZ6lZ48H1uo7Tbs9cfX91oA690uVtx1RFuP7WdzAsonuo2RncUbMKs
uSANFidz9oJyGxX5wgHrpvHSr//f/v217teVJwk7XpOayeIlNNVPpBm5rZHyiP5Y
EPVzrPf0H2JywnlKelyxVuU3ZBjWa53JTxAT0kmMSeqZTt3r8XB4YGFymXIUOLF9
A+pgojw5v0IlSWfIZTP2ddgHg9+APg+7jEXQ+UDhV87vrHCddVo4Pz1hTryni4LZ
aen32uhCD/T8/gd9Hu6ftHCTS8saFvI3l/aDcVBkTT48YMtkqSN9NBCZnSeLc0NV
fQsI2OSalXiqmkBf+Lp4Fminv2bD/+Z3wmhj5FbX4svADbvsrMlYAHv75tTZwuuK
Cp/XdxM8lFnAytpBnxYZOWVI2REzhsAYiKexpm9Vxl8lNDdTVfGs2Htrr3yxQbHK
5I7FNMhnGZvF54XcAjJikWxXkI+EbQrkSWtV8OVzBddPg306vyio0TMG9f2UU/II
gMCtTcn5Fe7ep0tjjaFG+XaUeKcITRJbBis5wgQReHBIOlgXR3t5UyWI0IKlD6UZ
UGivyCik0jOmQS0QfkljEH1lehkYIjY63FnGZ2z23x9wFqYR6HOllZ/YzO39gapm
JZzD+WreyXL0LlVH0epxPDNFhkvJvhOopwve97c2afmvMVKuEEJ6g8vQdeAD9I1P
PRtVEi7lsb3qylnOBPjqImxBAYk/8SZixCbHTUetek2Xfg2+w6nKhNIVxjxwoY+h
jLPP0r+U1rK6J9AbiVtJAfRfs90Fo/m78hDeWz62wFXxJWXKOehnGK1fEsQPVLfu
/G0bgAMzKZDcMk8Flof2O4x1zhfkTkhYjioWfYo+URlyckjtHVQyQZfe3KT1YQmJ
s3pH6kl9paLXEpSp+W2ekPmxqd6maHqOE2MVukCMwH9vKoU6PUkKC4jgCddSFfKF
pOvG2XR1kuO+D21CbNAhTTLgwCqkkbq8id5q6ZTOkaRXT3E65NX1xF6sVtgpa+/0
Js4MYPvyW+sIspXRIwXkGAtYoD/geDjpjhYzKqv5dTcsWTnzWId8eQTMEWTGXlDa
Nd8s30q1TYpii7e0Z3InRn0EsfcxOIKympakRoR7DU8zzggbH90Gyg4qbrSAwAgW
REqoVrmiiYnsdqy+ROKJi3JMOCGQ7lFW9lh/To5p105qaIYPgTDCem3Z6Dyb2aNq
KVYfAoGXP3aCvgWPZEOBQA7hQmTqaoYdfrSZGdUFBmL+gC0uoQnK02WRUEt+hRn8
ku5j+aoEZTKOGOSxR+rDlVgr37SK+z3CuoSPbhNWm3ve7VZnhieAyCHCxzhWRSGR
11ZT9copJ57/HTUcCup5Hf8cpm8fp2iTBf4pmmoOwnKxnyrqpPiNSErci/yQnfny
KrNkCoSiFBprfu/gGf3/Mx3tjEfoQRP1+6mdsVwjHJkbsVvqrVU9FbhSQoSz8sZK
23ui/v5gn4Cysu6OmX3CYS5MrxsP4AR9g5la7ieH9yrx8tTu82UV2sm3tOo0W6ma
kbZ3Xu28UpBFPcGvqbnvNpqz4d56k+nWwO+r4agolBpXwJUk1H2cI752X4lJbcJA
Hg9nKTyxxjSmW4H/qeuBNu3HGCHxjJJJ2v5hgkAdr2QZI/60D5xqgqEsYKUhxc/9
e/WsVbjTPX0ScE16+sOa2XW+jFw1IEB85eaIotLq36MUHwdhDrKd2OhHSG5S+EVf
5+NCz3N26tNPbeCzcByOPC1xErqjGNDZWO2LVkKi1p56FRP/UaNY+4LKXJMPd5LR
leP1X3fEqdhaNH699lAbqJAwU1bY9JlUgn9SCHy1VMIyc18IiGJz+4HLwFqgpHRf
2TcDeLRnyUvuX+pSMd0iuIRzpTDTPIVrJ/bdtVU9X9Vj51v9WY9pQLrUl/9X2Lhj
0aJZKe1l9wXJxmqvkmsmm1Ph/ej5uegq/iYEU/p/mmro01Q6G+mCh8RMgVhhVwfe
h9KQQq/2U/Sw4Bl6/iw/60qyJzlJvboWoUbsoHilDxB7cACZDAozJKfBY4xniKGs
RRuHtomiEhjiMMxHm02mQyT4R2LhMcaoTr9MqHZ0ci2uZEpIzrGNidoU7FyO3SI9
6BAF8NdV0ze42pDu6bn16DTyhftPuq9a5xRhbyLF6GdwfyW+XMQociTVlYqpeJ03
Rb8LRMJFzXefbPJvbRXl10iOM7aoSTHXUpZb8xjJmoLPl9UnG/qGwMOcDtJ+6n+f
cwL6dx9ixVDJ19VCuXY7rvX/Eoo9PmoT9Ekok1VGXOMIfobZtjsY57aS9pizZ5ct
r1bbOlpnTflAWbO89L/c7qhgERR6ez7GlmdOyVDj1myw3mliaLiu9IY3EcMp7btb
TTczaTuXgAUw3nKsev0mOMvun+/VKcrUrgwgHi5h8EhbAC3tIvtw6ctDlgbrqt/a
AYhUdEPmOthnynU+yZh17Oq2XT5Yys1pja8STCsmQzeyg4WZU+nCWaCTzIDlj+fe
Orik56WwZwarGi9/w4FtBR5hmLnya7YP2TdT77xQn5FYuzkA4gl1M2NgcZ4ILe+T
7twdWVv0CcMgmQcFgDLT5pBgBIdiygBkr6gcmidYq6kSRd2rP4sgumGABCEU6rqD
YqcHfQVFRiB/rSsR6RNOiKt3UrT3tIOD0vLzWgiUPn4BSvJuslq3xpxXc4hwpYJz
YZeG3cqD5UQ5r8U+1jDIrEi/gwzD5X7/lmj/MP9Pf8KSSNH67eiDHm76D1YePmm7
RshqUeswkxQegmSNyRkdfLb7AjFeQFRxou+DsCdTxcgC/1q8fuGGkTW3B4tidEBg
LljCspWWn3hx6zIrDyymSW9sKoSbt+nfM034vk23UNRRooNLIlbnw1p3WePB6Odq
uF9kk904miQcfQoJWgd/yp2Vs+vNQHVSRrxgzc3b8R4EN/Qwg3ABdSMDJwiv1rhj
8zIDwCgUIOmoq/HIxFYF+AjUW7BcZUmQ4ILZCIM07Fp9lrzbIQOfJcOUAvKtpLoq
rDgYRYKF9H5Uf6UeVONJwSROoOwpWTfvSnNY8GQUF4KnUmZDqKiCFefgsISi7KMs
esjIl6gUc4FPkdVOZ+BVhVoVh+tXuJq/T/DLv9BKPWbxNroDwZ9ILE9qR+pmqHjk
KssdpCwQXxKucFFCG+7Ry71GthmtovumELJ9lKvuOZJkjvqcTsjHLmfipP30Jk6+
iYTwffWrS8bnjdDhqV74GJwBihkCTGnIR45s1o3LHHWsClU9qxdMHWAT6BGf9yz9
6tZKrxBa0KMZ5SfQ0+zXZMgBPYZnjnlS7/PJilM+kRbdoD2p1RgsT9mbC7CUuRCz
HypYSHjxB1Q4+7nKBvfPMOMoWwxKCKXW3dQznDiyZYdnOq+n08p3Mqv8sM/4atU0
GOgCqQWl1XIH0TOdoVmfUvXcwOE7sPj4adMfq/qyJlI7kiQOjNuW7rxuwW9ykJaV
bx4JnPu5B7PikcS6DqgpCU4ZO3US4GA+bahVvLxbeG4VTBLRUnMH9X6GSEae8Dwd
zKZgWSlltwIwnRQPxGHVgHiCCgsMKayOUr4fEHzAs7t2SZTOqIFfnkcqXeA3Jq5F
axVlwte170Qz+3BLg226Wla68LlZvXZXBAg4bw9XDBg4DIIKCzm9xy8uOpAjRIa+
6ele8uPwu6qCVyjBWPGKJ9rwgmKhN9ky0YuPBGW4w4VeuWDq+4BwtgjBB6wlKtVn
7NMfJFzXDuT91gLY4q4KGX0tfdcYp4DO6/9wlFqZW6ZoQlbOXuXluctWk+EbSmgp
Qiz/6wP6kLOlpSIKh0fukW3mF2qBm6IuXHTIKERYVGj/Ga5/nIgIhmQgKXBx+oAC
h1fHa7HL5Z377aRSFVPO/l9G227gNveXYTMhTOqKYRklTZ6JYf/kTNcLOE4pnzAF
5zIknKCbFdv+NlaoTWlvRftp+Es3ujJZbP1QIGzzk3UghAtcIrbZF9sWXkkN2w5e
WWbsrsI/ProG2mmM7imak4UoPwj1EH8L9LRwLeg3VYwSrDqm6UQgbiA52g16T0fi
wn+kU5A1NrKqrI/ivHX+8bxCqVOlrox7nOqE1Pf7xbn4qzS7uErO174CwIIMg2FP
VjQSw3CU3H/yZMJIoSSKYZc0gKGVuDW6LRHMpA75JYuD3p7dvFjf0CcGYSwwsC8A
kPS5Y38XfyOvjWvk33GMhLFSV5/hv0F89YY/HrrWwX55VpaIFi0lJ8fP/oVnyon5
9rzlWuDqPTVxMQsw+XaMItV8owkE88OZuXTcdHv5L8Y6uatqnfnb3t34W7S5k+8P
moTh58v2GSvwPjXjePcAOxjyItKjPJr2KhW+gq4OvzoxlPhykmB2ebnzhnG5bQ2c
/YThZtzxq+YV4lsAZ+qiqQ84RWIJIqvfaMrhT0x+CWNU2yPiEk1lnbptUt57fhVF
hH6GoBzldSEVp89p8vN37LJwcWu00p7kCz92ZdJaHWWxrLAEJ2dj3ToXZIeluvzh
XbAFTi/l5mygE7gX8ApkU1D5ulVmy6xeqKV8vY6ms4Ro489kqlKTsRBQeojhv6Yy
/ii5scwgIxah1E1mV9wGZhiBpqxfaPfgcsAt0oRQPXz531u40KqQfeX3xrZlK+gZ
DkbL43A4RbQc3DKIENPQpo2muHIa4akHIv4Nacx28kNStcZZrzh25/3dmyfA4s14
SaZCQ5KB0S2t5v7Otvqcr0hzf0UGcjQMTKeZDfmaQgmlq33Sh3pXmAF3BVW1LbAY
c7mL7tMUZvxgKFrOAWyFeX1OsU5nb26eVT22sqSeCyezYJ5jsVbiNOsGp1hWqawb
6ZsfrMMBtuJsWXG1hP06mjRdYjB8HBg4e7YZIt7q2HZh4ntr13mL7f3XGfITzkeK
XZgWcVH3UTzGC2fEGVQ8ISeKZ8p/GvE/t4CAqdJhbTysv0A/r9N7M71kxYZjZCsy
JcB2cRjzU2ZJEguQz1r6huWQj5TQS/nhu/7qOntQlqNaYUsNkTzleO6EB2UhX06Y
Chhj0M2DQWaHe/d9++c4OSzd/R6JiaxCmHWDOSXzwPakwnA6zLpiR2ZCDc6bM2YJ
fMBGSl4kWRhdXPN4+k0rV4A9F1+fvSd7EdmE0y+NewkV/9oYqGABeSYD7qIvw4Vw
Tb6Njw7PJxotgnVkHv46sTG0M9DUdICsdjXI83+RLMEDlx3+6sH/G4uYFH+aw6DF
qDsb99o6WMjvoZezW3IoajYM8qJvmVB6dP+dbYcDJK6Kq7emqKxcVFNCjmboSc+I
nuCAWxQSyF3teKhOWZ13N+Z88yktiBwA/1rrdtP44Bjd6rt8slHGk2lhn9ghaNp8
rWRGW+DyONEE9DptysxDPpOFoCbuawijcG7bEk+HHyaWr28r+ayJLbBOc32pf2ol
x18fnLMqXzBoUEkryhXNLPJ3hpkhjS/NTiD2rVmGIBG6HzPNdJRTtkJcE3Nwom+B
EoLlNG0jm45vJ75z9jHFdIO1NMrZTk1AetbEFR/HR+aY3V9yqL2gZhQt3+lXhyJJ
l4JYVDAalD+7+0b+jSUyspe0efi1V4Jf2rlGISrECKiFfyfrv4PwQj8kUStgM+N/
EtDBbyegbQh7H2EjoDnrE+QqkTj/eXmd0uEZ05bFrCQQTCrCe14++uF2nF7S3n5j
D/UFUDcqTp/SDZFxTzuhpx9GaLqAeNFsPg3637pp2XwjVTBcUtaqQkRqYDEIsrMe
B0FQG3+sluZx/VJY8RBn6oC+4At/upG2APR889TdqQgkEiTmDAkC0XJgw/9zL8dD
rOh0Yv+45c08KahS4Sq3JAShjLel3CO+/fgSpdgqgNfj/PH6Z1CBSJgST53wB0fh
PJnnqNJG25k4V/SHYj7kt6wt7R91VrekeVNveohxBWMsOk2FNDtNDWMJqiJN9T6S
wQIJjZ/H3CI2MKa0M+LBq6hJXpeuoGwu5L49aPpe4Zuk5ggQ2ZYaTHbyYh+GHqDN
+5oSVYftzGeGo/hIvKDxusSvyOJX7e2EK/9ns8YVeDJOyfn9ND5PssazjdOjkbpJ
Hw2Y3sKuXxgbYgmSh1alv3Wo22bli7kCo1f8uOe7YGZzyowh+1yB53y/InciEcdl
b5HCyl6qiRO6DRQFLKi/ZjoFivro7zzGFPIWxw/AtlxB6NbBr219vQ5m/Y6h5Ahy
ESsLpKjda+bCAxndAzHGdX2v0C/9oeYlDBENYLMbcaB2z9FEqC/kCq5hpjtRp7PQ
X7wCfMo6kXpqeMHfxFkFfyqemoHYRpW/j6b9OQ7OJYcrAwxnuLsR8GVneN6hsAB+
ympPq8ZAJ6lffhUsmd0fwK/CNP8xMzKXJm/WEvdem2v82SpaMuhOStUGvrHBow5g
MDMWgGbwTiXhmXsIH7xxb6rlyiHiLS0oAdKFRXg1d4Zf8hp1brI3Ppw+HluZ/R9F
nVmvOtQNVt69qbe5XUlQ0j0mmArmRxGtP9paiHnUnt6ZkwI5C2G+gVsq5B9sb9We
8xRYriZA2JWDK7ha+Kno97Y+koJBvOjT7al2brVPE2t93quuvVZrkfWDcA0m7Z63
maY2EONuc4ia3lHTx8oEIB/u99C/59QAhqkbLAPonuoVFzYOpur9R34Vwq2RXsx8
TDp9H/81PUY3qnTbod5059FykT/mSxFw8y2gBPeDOJnlnN7JJA2NsMcMSCTV6xHO
JiyIFB8FMst9JSkIFFfwgaEC71AMrmkaJqU3eKU7a812O4yK5Gu9z5i+yYc3OSdd
1Zq6VJU7OWcNujHASqfacnXQ+4yPm+loHJp73UVgVRT0rFhz3dTfKulwmjWg0hxw
FpxELryM7Fbulw71isqejWncHOiEcMAnB+9csqfDhh5YtUOOyjiWhezMM64gLwyf
F3UIQ/CCqpa4ZDmU7PtCIqtJvKXujkk+la3xWm3u3iJ4ZwmIU3OlCzCF4d/0Zxmh
zfjpsiqHfHH9qrUujkq9ek6da3Yp/36FldgLLsUACjjU3flfkTBsi0tdoin4Xno6
/69Hb1ERmtldsDJB+MrjDKreIU1VSmwSdb7i5pwrYFGewlF/354QomgjulqXvbnY
asq0estD3bA1f3ZjgVWK+tSTa1DrTLK6kOmAQcqQ0u8pkKJxxD9O5lrO4fMmRf4C
xHdSFgXgNLOO/d9uI6fwn7LzMzUdeDGKUb2BcJQ+WpcHH8H2XOonXd+THZVUvStj
GYWKujX6mDHDtf4CVmFyqeALE95LeSZLu0FGjzzWkcimR9kcJnReclD8KHS7Simk
5LV0BPA8AnGRQj/GjynMevzzdZzak70QozpYxtyamftFQaai2Kg+pWjrfy+nTOOl
yfJZNe/zaLUJ0hjaDF/c7vs6z2MnfnvA7ins74yg03neYH2rTdCous92x9SBbQH8
5pWprp1Fwhfvni9C05ViJbYpbcBEcL9QLmjsNz1CYfVej0ZDcx33k7FOtsk42gIO
MsMhzJJzYxDGHRKqQzXNmp9mRd2QGWdWA/ODIst0Trjcv/BMnv3k8tsAOA9Jznxl
M4og/ifTLd/FPJqcjicvP9YHeB40/tZK7bBEMx5IvmV1IKiaL663TFs+1QK4YfV/
tcBs30FkDrkCH/FoeNyCKfpzqNlVBKvl23s/TSn4pvmrm2pce6y4/6tyr3xpqrly
AXyB3wBQhS6TDzYWfbx99CGbyT7cwcG1OOnne/XWlZiokwDHcFQeortR6pcGfy8W
eeXKq6azEgocADPJkDFiXDi2Uy9JIybRDe9Sl3XCUdlN8u2It92pWY1lJj2mgyy2
TB90cBIWXWVrWrHpOay4xAXyBGP873ZfQTFezzDK1y+2EeB2HP4TueB1Il9o32Mc
477MzVUgt0wF/cPKFsS2VZMtPdqJYcEoJoqx68Zu1+wkRHNucuXIVhImIMADvgoX
SYoKwgF6DUYTEkXUZCyqwYY2HvPVO6wQ99UJbK92vK0i0ePYmAyUaHPsREcTUizf
Anfhk17OZIWdpuBB9oVNJqKLqjZZ1kxxwh9kyVlCeVvQAjlGhXAJUAES3HNfQUxi
h0E/R8PR5s2aoiqFFtxdYW43zNYu3UZbicwO4r9WLO2AFfIrnWDyxPhlyU2lDP9t
flQrqau0OfwHEFsrrqknSpKAkRBq+uIhl83jK7g2JvK2tyX67rU+kcgq7C5JaCmV
+MLoB6tskHK7i6zVJtRRRfb1L+lej5Si0TNHNmj0PBxdTGnz5x+RK5G1iJWZKouk
oPjioErhm8Z4TFHpnA6xHbeAj9Exbl3cA9Z/wjxXYkLODhl7MWBiqTCLqUMNS0dz
3439tAtq/EI5ML8iaI55ysVwEXQ/uPb1/+jXFQ6yw360dqUT3Fd+e7VtPZuv6Fr/
OuDi4gY8hZ9mfWCOsXW7PV8+W87PxbUfXk9pQ/RCvGMP5kBMlzhhPbFJ1qfFPReQ
6q/Sq+8ksNJjANmZcQBqb9ThzRccL6F/fYFkbHHk016HdaEA5vrn7XYT/J8FLBXk
F1her52VKXTQOBXuNYCvDDgman6H5UYPg0HsL5w99vrlEjT62OX/mVjpDORQyAOu
BO3K2TEdETkrJdbOY2ixTq+TH1d6h32GQ+2kKI696+RbM6FI9aBmLJ4wlIF6MXEp
naLaSMzOi392rYn8NCFRNxptupWTM2k515wz94r/u+T+h8Kbzn/YEbuDDoIsOFcx
yeNVp/L7fXybFjUp7xjS4/IhcXhRP9dZjjppZ+ZmF834HJ6XIwgFPSXSuhuZmzn5
MtQ7rxTjDM1RB/hJI+FMXIkAoM765O7IDm9M9i2Y22HY+UV1x/1EyckVEvAVdkfh
NNDnJB94DIqxLZXuZt1JjvzO6EzUVtiSsQTtpXQxN1872bwjJfA7sVgohMMcf002
kI50IdPIdsq/T/5rBkcGCmUScrSY5jjzpeyfqrGgTLJ3j/5+ElV7pAa2AQq9q2/E
SrKG4TFB3M05lsiw0Mcz49/AnQ+LOmgpv/j+YxJbCPOA2siVQ2eB1871SnO/PeeR
cUMqnlvtGs2MXVW/amyzoodCAe2U4rNYuxLmocpaRhgoRJD0Hi/tJHLWar1oMtD7
Jqf2a8/6Fyej7VEEtKIucKUF7BAVFowzIoyfLQ1Z86sd2zULjNDgEAPL8oIw+hfh
czuNz5acb4/rh4KQ1Qty9QCzNFvH3lFu4anlzQuoq07vyRucW6D3PZajITdzJwyb
SSQneb0rLmX7IpNWYunAW8E7JW81fMJ5dMnM6TT4ozxcwaREBXaAFEML+qEisU+Q
zGWUU9YGyoiom7q7l5KV4JbHtSPbg7plyo9FdDWMAoErLfMONB/LX8rnPLlxXT99
a0hW0VBP7YJZ6PkVVSjl0xSUvwcJvAHRKsM7ec2mAaS9z58fpKJAbx8uUMoogmqj
KcNY2Q1yCD8ZmN4PBHqo4/HzEQiCZ7wgnItoOozEuUQBf/I1sL0deXQwoOFkwMgN
i6uz33kR3528zYy75QJO/5D+rXJRGOqxfGwUSSgCn2cX632zQlJ2IW/Mwg4PGJCT
03+bdgIkSddBsfaktJ55i5nUnxTCxDI/KS2chwX7kF+nY6cG5XmPXabCtAxG/8LA
WkLivjQ4mCUKs3gAAL0pAOrkL2Ym74yQ5HygIGJj7HSX4xtZnHNBJsudjXaui62R
zpRk7CqKF9QoYt+vieEV9qNn5bHeWopYNxZ5P1XE1FrYJLykVkPnu0XqCtiqcyaI
lQpvJkLxOPYdjyBZYQ+9vhpf7zON9yAPXVgNfMlA00Lb/oKMAAh8L2YSUEk0WQoO
lMt4Kqf7pwxnG05K6RKsxfgWPirtcKF3gpKwjQJd7NEXH3AxeELHU+8e9wqa1liG
hEGRbA9CuR4JCHD/Uld5wFxWH00S5iKkyHEjBZd2CI1MnoI11EBQ99U92uyr7EtI
RbVusDH/7S+Zrh/VgEdyszkDTi22XkT5nDO1kZ1H05tzk/J6BTUqtR17BycWnQid
8Mhfhys7GmWJXOwNfs/M/q9DnHWvnpoEMqX+UImA0uDmc4Y9nWVk3sksCCUgLN9u
uwt1hnbbZYAfjYRe5II2r9qZv1A/BFzar6HnMj/up5/YCYNMeozxdK0sWN3eKuwv
TxXxS3E9nJsK4AMRTCH2pqyIlZHru1Cf0Ng+J0wl0HZNzpcN/gSHw09Bh9OHzxb8
MPyTDcYCIpjErZuNI+gQH6D9M18f3tPbvmMK0a6AP1fuM4Z28tBNXrjX7TvvCbLW
oinb3C0kcJoLH73iBdV8PnN0xWRYTFwF852oNqLJ8+L9c0tMCJ5RX5ExdPmUi/C2
igjIRH41T8Z5t3nV45pzP7smIKUGj/HnpRu0E9bU9CpPvXeYQKQ4IuLRQhKLJfSP
0ZMlt8hqzfQtwzyQDSxzDNJY5jk9gHYZ/YyvphVjAsyD4HEacTew9FHyEXs5c+1f
rRleT+xXjxXsybrPn0af14hrXsyN4eBoqymgmwRdic9jrLFhsZfUHk4G5qNurSAx
0KfECDcL+7O4P7QMY6TNOqFVXvjLBPfG/dhJ/J85HsOW1LX7l3JrBwxLwBp414EU
8zGjv6PKLdaZWX+UihbyATNhHcK3aWBDK8zQpHw8TpVrjOB4XsEitNyhuIdTG9g7
HY6M7HB1HrG97HMi1pCV9QDJ8vW5Lu0Tqu41MqE8HxBcIZ4YtoYljweOKDeH7djn
2m8SrL98+iYydxczcbrStuyE3GTL7efSp2hjhapOkh0eHgoPYYwyv4TCeo31tuCI
vUkRE/6Er4c7zhOVBbkoFYiTDv/iw4mUrwlEoXDUjPYhV8keCq9xChOTXLxVeqxL
P9WTf9rdsz1KWcOYEWvxSYJpwOegPEl9pxUD6cbJzC8RTHjNqiRr12qANuQln+6Y
dauPDyASKCMB2sQYl4FoPlLvp8RAcIHlZFGm/dfYKuDHAm92LNc3vQ+R0ddYWujr
rPU2XGp177AWg6AvegSmVkDGsG/tCM9QIrkRm9NXz9y1gu31rXJgfE02tOrTGxWi
weVoOuPuc3cse+kR4CBqbliIfC8v/EKh4hBNG3+cinVcvMDcGEc9APfyHU2SFPXK
1G+4vngmMmlo2LgY4RdTkWgX53Hyuf8ENhayU8hYZIuptxNapk2UYKeVmRlhDDCq
8YUoryMPztVlbQeYdJqyolmiqLwGh2AdcWfY+E9vwgDGQZFRGQYQyL45u4/g1UZW
rj9S/6CqG40rjUVVYwiFYgunoTNRwdlMg6UVt87v4E365QH4ae2cNlJF3NlLlCuD
ebCZsQPYGmmxAzLdW9yOJnNTZafO4x2AsAudNUqwQiq9aN/b5u+ZeuW08kAqlRI1
PpSiSLxwnqPVAChwyoc5Hhd2CJyjGZcxYMTLvSUEL44npRnoTOknHZrPuxEDbV3B
oDJ+UbWQkq0r7tCSYGA3v2B+fnUy48zo3KDQiLAtUsfU9h9Vhx47DaD/WAFwxVGD
ZOWUu6oGsF8C53GfcnYbP8pf8jKRfF9ZTCoJjXIfj63bHHaGGkaaS/NnMQlyGyXE
GgJC277KF1EHxYVhg1WiccVpHbtCdWn5W20TxTC6cgyChv+Crg8hVpvLigQY595g
wjnVL8TUVbAGr6E+MtzLq+hl1nrJL6HRbQmY3MrrTZ70YAVvrw0A1jZIuPJgLkdd
Q2id/XN6NKyr9CkeiN7uWafBAX6Q/Nw1ZkiDqak/ZZokEaOIOcHlFqq/Og7NXg2Q
bu4h1LsicxizmYpEQ4ss3OP+JKiBpdTIq6nMjtDdepuUMzRoq1vZGZ1diEYRDe5j
snfWZwMa511VnaDZy8+ehTxw36q6Sr4m+g39LsjAqy/iPTIoSekXmvpIuBJK+84O
PEhnO3hoc3gS7PPo5tpLa8LI48EJpm5nXtjGpJPgNKIgSCc5Opfkc4/eiW6/zkC9
7dmmFhLWyHwIyqwy3EFlayrNeHCllRGr5PZDUnl0ZVGBRuIzPyhWeS1C95sgI2UA
9OfQZgOGcE8EyOE4kQQmpHCNNL7PKZasKzaFqxd3s+ngnWgY4acQ4uphcKM0xadY
9mBOD5gsWyGDCvDcIgIBrWyIZKLe8KYYdsmUL0ovx/V7zo1TeB7x22MImxa5WPpV
CSIFORKxSA3A8G8zvR1afRK3nl1yxWyNDrbr7/M+cAYD5jX07O2J3HyRDnpN4H/T
4zUlS1FGPeHP1XkD67jOPG845KTKPkiG5u0rqaPwSFP3xSP2jmNerHrpDurthD7f
wVf127kTk15APQ5ZsdYCVlqym48slJhFyywO4i9VrZ39bF91GzFyrilNP54SnQU1
RHHj1CrF61SOg3V0z3wuN0F8r1tVP6y2l2Nf/skEd7XQ8cw2tMpyoYy0U8KbC4c/
bsA5oP4uRwD5FLw9DIrECAWwFxjc7XAtocBRrCIoG/KHtA5QfBZ+Y9Tcgugv1Cp+
Cc/yWfWoJ+KuqL8Wv1oD9hBN7Y4i40pX8CFrgD/FrHuMaFg4a/wmbmXJN/dRsSkL
4WUfni/TQe0cQ9CnWg5npqV1QM0z9at+xYKnaOHz5WYXnpvc6T6rTWiR/Pbo8SfY
JdTFQ17ZQ776d1C8IMEyVnAsejVu8fPMHnFjbzSVa6yHrzBVcIJG6SKuSJF0OYUy
/ylR5mV9S/T3sDcnJQ4tBG15D38+EeVuolEpRR+hdmIaz6bV9Bk8SIwgqTysiIva
SRz7FM/7zwci//XAlBbuqTFX/V97rlbmE5lQ30xoMJsEZnPYE24WmCdK3GeuXWe4
rhMaXxLaNM2Poqq4ijIquGYuAl1DX6SRA1XVXu4l/T0TDfZ5mbn6KM+lCNVYEIsB
dDEYIXvZcXUddLa3/sywmdhzlXq44UtPZZ7LqSc9znT0fcRoitEUZopE/mPvP0Gt
kNUwQwvRmRd7ar5WW/kQalgZq6GLjoSupSRIf9P6/T4aKN+IaNtuKyU3wvawsMFi
govZH99Wz0RVePxMyumkNlgozFSRypqtwZF5PIlm3kQGJmgC8RWBzUp3kZrynEK4
Og3ISKJvtRNeEecBXyKVLWjc7xg846va3Qe14Zt0OJeMNpMJTHltXgJuIiNEcbG+
YTbxMbJAoZ7381eLSpmyUhNiAIMIacXDebfbe6UwfdZNdNRWgHxlcH1fQLNVn0HR
Se9gVt8MSU0dzSUWw/+q48qIPzhQVGbipe0sdZhjC8I56XB95EUmWo6UXAoGrRn+
JRgEnKCB/QUlvVfUaNQPs2f2g5wTNcRyliy5XgmsE2w8eRL37XYew7YCTyr3GU6j
Zvk57FrP42aWuIAUOvAqMsNc21gm+TRKgvtDW3iXwB/Ik2vJENYrf90SpNQDuVXQ
dsXPsiT5n0RwCJOT257j2Y7cQWvfk/qXudrehKFhZ2UctMhRXoMdZBuXpp+kzHrP
Hwtrj621KhJUR0ikS+TBoqtMhE/wRrQihDRZt63/K9+6845IImsSn4xqn1u277gR
CLV9vIgAgMggohAEHfQE0/jepsvNF2r2L8zxnKDWa7SuPfJ4EQQqZZlVVvRfRbkS
uP+1TWFLibBJxwRhzFiEhmxCVJK68TbxvEWLxphJc507qUgECudmHpNpEut6h5VC
GPOasHJ6SrDgfdRZXrTXlfEvTtNmuo8Io5lMqr1ZVm1hlCOSl4NEn+Z510nGx+1s
1xWTflKXvSmKQXMCqpyyPiCZJH7qoMIEGxnZtqBJFdwm5Ogs6FSTD2czIKQv6uBp
tampvCSnxr8sVTArnCUK+o82PluybwmodznjWKWIMwLW28N4m5GtBGNEuwlH+4AB
tiq2A9qkXnTfCWsi0gyfDC+cXO4offwj3jjeI+95dkLJYGJOIx99ilkTwV5gZjAu
rkgtN7Q/CbeYtlHLMP54e6vHoOwNqcUqgpWqr0zAmW66Es70Yp8m1k+5n4zocrxh
vLZzSKskwmggMxnanU64tT9qAOelGWU7LLxdxPejxkVdwknAEc1kHP4xfc9OOb9o
MBcTnwfdLyBCZ1sKSNMnCVzIjOOmwWdjmKzwW1q6sJik38aPV7Md6C4F3tR491gk
97bPIsWCg9CyoR2+GR0ph+pVnEqrZpMqHmiMuFNxCt11ipRH+hiKeXgCH1/kElCj
0M5h+PftZaoZdkl+R/fMG+gjhfB6GqH7fLeiu+5i2B3wjiXy9Zhk08Sck+dqEvb+
U70jyOEvCX+1f1TRQ5q2Uo2pEJVwr3QrDzo8fBZle5qzvX9/uUUYBcKoTqfaW8Sp
gA0ZJ2v/XBGAiVWXIW5e4FOJPmWSYiKpqJ2lzoPmO9yk2fooHP+pKxI9R6dYZXBv
/hIOpDWGZFymJFqWJGuwnTSEwgbnCPJNc3qXJ+OoQnIGiIsRxtq6uzX2TSEAY4tB
MzLRcPlRV77ZK+BAtJrx+jY1YAfYg2iM2fO9CeEov/SbRloRkFxVMazuQ+tpNLvx
LTEAFCTMPrzb3VH/PSTpq8M6k9z6PS8+i8W6+WuvkLCUm1dF6bv8zxFZniEzGQsO
vccsEPHcw0vLLBVyzYNc/xtKomG15MVRaFI/tlxQ0Ues61ZeQ12Zal5fVt7fk+g3
WJSTr3O4LJlKlhFNPpUcl3s+Z789Kvr8w6pG/fZprvGrR3LsiIxDIWiWttuDcls3
p5h/AFdNblWiL26MF/bub1hxBFiWKEe07r5eHuHw2qL9VPoZn9HLOLMPRA2MSiau
nrrWvtnMkQ6OZ8VD3+kOHPzTkV5T8s1XUz8wtV4aWYYcujuqkwVFntWfZMmRwRZU
r77otoAQKtKdHCTvPnfNcTKHyL/5DV6oNlk6or1ZlEIFvzVqeGLhEhjCBuj0NAFw
TCUDI23IMTc69gdLrWuLvMxnnTOWgj7h+hHPH+PPlqbfWy7HS7zcTljdgcKPoKBB
BNXHgVSaw0P+kokZ1p65rZDlE/PT0MPewHIwm11+RDsb56izDKa7hH2ANJJkNqkS
m9nLd6WCqY9XuR11xAaMOWVzB2IjTVeUt4Okt/OWyUl4A+YuOxgMP0o0U5pgjmvj
aqrXOA8VRQMIXP9Nm1qdaJdJjjqmJCPXr81wyCM7s7pOaBuRwcRgVG+ZPexoW7EU
JMYQw9WfmPwM/AvT/RhhAJlruX2sKyxNksEsUT94OO3ANaBXdviPc78K8RiDzvWL
APXAptLGlWh3Lpi5inF7Y8ir0A1fdi+fEnRTreMbegEjo9cvM89dVfJdUX4aj+NO
7guvV0/NbLsNlTGVbz0i8NYaJBkbRHSuOnntSLT9wXkHE9kOz7oSqDvTEz3YLm0w
XScOwiq3IX6BI/pJ3t659s4O0I8thfZmXY+vO5SSDU3AfoD8QsIRT2IjcDrFSoYj
fYzLfFTIhV0RxNtjQDJhyijifwF4ErqomS7NJTfZcw0GjIww6zVihVT51sJ5mNbO
g1LH/MR8MZq5Q+ybC6YYcesp80wIM6WzwUeJb14dM0KnVBjeIA+2oFKJlVP1IgBd
SS8ziXmkrcqmNeKvLX83LNnrlRrkVSRBX1E/c/I8bjatpgY0Sj/FZdpb1llB4UBj
n0FaR2O1gaDFDTclOzUb7rJHyx2ncWDY/XMx9A58I+ttBGDGSoBg8GEW5ofBymCS
piMzDgBRLApqZp58tzplTWm/o8OMusWVJY651Eo1zHnuAvMVpK4lkRF3K8cEnH/H
Gy09Hs8YJMnHDraSofMZBmLlu7hIxWeM/vdfKa7Ah9UlAjY7805xkL0WueQpd3gD
ABJSFhYCLIe83YVmFmv4YSISi22vGsO6o7ZauHmB1Y0x+u9aGoNlKgiqzKxvD84z
+GaaYMPkc7ZdMLetiRgfQxRQFz56vhxqw+kclwCfRm78xdjjavpLKmpwfBNj9lAC
vZ2dPefy4GjRzMWLlRSC6L9FvPWtiQpA7aDGzx3ugBx4Xl1UHk5/RLliC0uezBWX
CZ5KF59FsvKd4AV2SPeyrgWIDKR6BaJsOwl0aD6YJfOhhQYKULxLBlMIH5/U2LOz
d1MI8ucpj3+lY/qWt2HbroNYCvchN9AEl+W8wf7CGUotOknZ01TNm3yx5RwqNs/D
jg0mdiRIyg7T6CsEVwEoChjztYH1UdOpwJFGy4GaDyBuRH0ERuFWFXK8ZkNTKY1f
RugNp1F2HXQHo8PKW1ZFRTqUNouzgV8rzHBvHpPdxWAF/di5ToVYE8S/VcD89PBM
FAfhF8XK+4dhkJfpH0ubkpMwW8oPNSTvFwKIOBNawdOlBoqZ1KnrA7wMGEeGeQm7
qi2Wj6GQjtLKN4z37S9dvJFQAWyvSepz3BO1knrMTWDiRbGF2k6VKDqzp43lDEA0
TVxxreh2B1+ktZLZOiKw2slW2lsawGQcog9j1gHis5ishqYoS8dbQzrYiycAtAxc
j6Av00s7HnaMHsyxhm7RUK5dd2szXN3YlPOD5wMzMfsT6+NpkA19oPDjFxo+HWqv
fkf3M6VG42mEpIhlKEhzwxqTSa8sjW8k96Y8w+l5ypsT+PQ8SrYJxyefOMZ+lZNU
kLCbSin9KnTYMRr3teK1pYvuFRkWo743+wjC0YwT7WQoTSrg+jP7Yhqk7KxKVFdT
rJx0r9le/Fb/N/oUNlEqh74HNO2zwspo+j6Dz8jf/26XonM607cnyvdW7Ihhn3aD
LaLh6cH/32+mqknXmdIkYkIjsOWMzUoyvXn6/hOwdglDz52LiFAObJVWe01RuEFT
RUDFODR9qcIPwd8cLMBaVhhiL8EBzPlMW4g2DDAjmbVfSFpTNG4rMtRLmLkxU9Tg
FmCYo1jOaKTzQhVp3HfWMWhE5D7q4GUTR4yTWP1YaETV8gyO1AmpSf7FgrSXBq44
PkGDmtehK1sxFCxnS2IHKQmbQnOlMoJVjRv7owUGKVv6Gr7CoVw2JFpnCVlzQ485
oJeETKs0yxiVZ4WZBU4J2xAqaMY3lbwJ3RNR+lFO6RY2VdKrBH9n+QocPNdJ8ZAj
IJHtMHHuPSogNLtRdFUdPbnZa5A1zXe9Ek2JEsFEm6FYSDVVQlvoyvw5fiIQ58rf
AICQmBsHbA88DU82NSAYq31tNkWqF6ajYEZiGK5LIkT2l3WxoRZRGukM6y5rO+y6
sgLEQycLx7vxSIoVj5jA01RAmcXSx+6R6ja1lQ/5/zLJWAIKh/qcfs8xH2joN1po
Cmsl3cwScRqNPm1kLB7UowE41oFUPGeM0iEZE1MY6nZATmzb7uOIuUhrZSb/EObW
MHo0gnuOvA5Q+kfM2yKXO4WxBc8Rs0yRZXd/cFtbMv0GmXAURYc78omtrG2kEt1m
dQfNRiDZgH2usYI+xlUCbarmg5PctzK40M8CruKDakDXRkmq1s+ATqAqE+yJdpP2
4xOZ8QL5mRyay7rtsk8nOlRaO+kQf6bLVVYsXW97YXy8myJaNm3yYO0nhMZqeQXh
8dZsMfV2/tgRpTgEGRvrW6GgULd0Ep79eAp632oGYAzahk4ykwNU+WvjEKoAyeRm
5w5cj4EY11SOWEQfE0GKJ/nLtQorTV8Jja6gkBTrWyzlauKCg6tC5r6AESrFNyXe
/jdDngfBW2lDfzhvllAioQZ+ugXbaSiMjjGrafbmXChxBJUt1H7sApkZsa9Rn9OJ
AZ/eyw0SEIg27bFEzJJUFWJAMq8XRbkko43S43GX2sYEMmWFF0yolZzE8efuHElt
aas5y8Z5lFSZzf6liL51OMuBkJri3RSm2HPiCd/7gPvdO0grkhcWPMhPul2WwgJN
tiUR+BdSJvnVVN+1+JlmsQjdItb+QvGFx0VldO39g21kcbmbN5Xhht+liQtcIqGZ
QEmFNClHFh6DUITmWmYMuCV+uh3c5VcFGLxD36UHyrVOXiAHMSe2wccmzd2B7I54
CQAKDbRbeOfm8L3SDl/ZE62aSSPLPPMj8zeBqeVFcIfCTbH+XnMwNL/vfqqoe9NG
yp+FXX7Yu18566dPv8UTjcCO08rC/BrQ+dfxrCt1UBQABm+jC4DQoSN6Msv3vsrA
spap+CURbQ2eyLNkyCUoHdCMsMeG1aLEsJyJrv25LEZaJag9qzexUMQnc83/f29t
hEc0XnkuaAm6K/VYddxGriQkPVOVxY5bkFJnueIEVdUyA09hZ5p+i41r8R92/GcB
4D70vYogO1zt6myPv8GG2+Lt4e4BbDuPUIAVyAGjVByBNAquioXy8CVkcwfFEbD3
y6raaCg2SNtRCh3GZF471W3pxbKG12h0jgVD4bQ6Nt2GGJZUnwU6IcnXKStLimQr
hL0as9DymreDBldXWdaoX8yA3anui8FFZIzd6Y1o9ivb5v6671gCc1sA3/uREQW9
fYAlLNjAkaDQqhKlbBqO7ppgbOHOXKO+1yCt8OlfvgSt8CQRBuNQva2A/2ECpOBW
vlu45gTGj/EbfGNDJCjGrX9pvK/vbnZpXXP9CFWmN3GAnzRn4Z1NLY4Muz3d6pIk
tP5jCk8MQavMCHdXPP4GslOfY2zZ9NFa3US629BeEhBBNkzga8pZK5C5V5225uob
MrqWyORPJhkVK/E75nYhfP/lUqO0lTuOb/9epw1mnzvZbiydOqtxb1J6eCUvJ88h
5Lo4FJTNfoVgEcA5ggGljKtL5TxZySA7PvVBc6w5+LpIfUFAhqpu1YleBQBHIUMo
Nsxj9xct+m4DXe7qyJa1fEJkgZydAGyGk4DN8bEukouH/89i0+rUvcAoC/068qfS
mGk5EqTZtXQmaU4BGP6JKFCDzKMrwIU/cyxD3jcxrulhTmWCNF1t9lXz+zljPgUs
63+ORcyZ7cv8yrRobmiTZ/dWMd2tDVlLeuJ6fcTvDouT4YyiMyrwPB4XAs55BM0C
S49YtvF+Pban/9AH1p0TZw/8A1PdMvJ7FRzmhJIJ9Az8PkEd0kd2l0ckr5hbqvSb
zK7pBNXTJU1Ir15u9AHaSSMVZxXtwramPIJe7bYYWpk4QnF9dS37/+UHGuW1YSI4
Yt5e5T2GkjkltsyqPU1u6ZHA8z9j7FLQod6/ULe6g2T07Mg3wl1kahCNfz/cAOGY
B3M8woWgt5RffGko8pwWXneH+t1iBiDx7MeKy8Wz6inlcNDD3RUn7nkf7j3aTbkx
RXsRFNAJ7TAfSD7vhT4ImQ/ReBuDze4q2hRtZ6ZAqTfZZj5cgKjwzz4Me2f9yEaJ
yuDeCKY3jHuSeATr7UCDeS14323IZAYraj1kP5TFrwEmWTq312qC6I1b3EHA12Bk
ukLV0ncsj590j/OeR/z9SBH6BhUwxNJ1tZIdyxQXVrxOqJHsletX8txwlmpRm8Se
BRKhQHE27iZDNWhb9xEnObzUyBXqxVOojNlta99JufP34frroWJIY7px+4RyA8he
ofx0Hp6lZtOje0ovrixj7myhlvHyaxh+Ts3bt2n3s9SS2wtPRUzWfcIp5NyHbRcK
afcwZywjXXbEWDhU3jyyju9E7I/n0Bz2jMJSSFyX0o+23wzm0aCNFyzQBsE4MLKg
5Nmfbs7tHJiO58LNKO2kCNM6vMy93WLGb/n5hNTbxmn8RM3L0h/M8HF+FEw+qnGX
N75O9xjXaNiHm3DjYk4SJrrQ5Sb76P0XwQLFL5RtvTpMUhJdOQ/V4CPlczMETAvj
amK30BsJKWFI0dUbIR3ycNWqBrOYyd4IKWjVEk8VhJVo1RiTkAppxbZMmGldALA0
oGLC5wJ5MHLZLIqUb3fiREa4Dwdb6PFtUTHo8jc0vcuj6iFnpfuhK5aOdHxy541d
pX96wg7MagaEk1XWEP6dUqFv9sgC9mh+fVrVXYxocfuQWAiVE2JpDt/7pkE3j9op
uwazTiSfV6XTzQkyyj4VOzMCAVLP8gGamTKCUpbK8LPp3P8LH7xI7yhhwkI/NdaB
ErsIYP8n9i7A7mQRY1LGbEffg68vw+ggY+9JbaG/4g6OPqKcHHlpcf3TIl+jU6Uq
ho/2yNs+JIm7jj2MBgBMiOEm8waRrUMLckpMVokWvoaNDy4+Kww47zfsSMPSDVZd
xPhFCrTsD5ulcEof6iuS8UPfzQhaVc4/gogy1aewC7bMrJ9RamDXW+2sGG+vzCKP
dUITbl38bI28ILKCuDOPVwoJ/4v+qedEuY/xuVTk6MKMasXtn5HHBeMdudldi6OH
iNg+OwRUR1t9MmErqH8izJX8+K5sLjxhAh9GsNpGxwSb5w5XH3CkJiwYjpWce/27
6qH741loPsP/ePEtUdgDoBIGEOWzmGJzVYzt/8XD9hVgxqav2Nyi8niynEkh6JaK
kylHfN7ugP0SDAwr99F0Jv8BQu5ZrERlcUQKgiLVx3rT9r8Cs9MUNsA056c/zfGS
x13lr2VTcPrp1fjGE6rnvhYk12wva8dyggQD35O9fLDfTZFGkA8smHs7wmuX+MyP
WmpONBzeW9I98fI+b9P6dA2Kr3zNa0AKIpfdzVTR64JVzJq+M3xblY3c2dze695Q
ejIDb5HZeu4tAJjrn6oPWITmNQy6chhViJHfQnTAfsLKdX6fVihIaw4/FkxLoulT
SSjkVkHi0qQvrfTJbHan6VB2GA8aihkCvJ6VAoqbCYcd5dih4T2XV5QzDGOmxZgO
rvZ1sGjnZ0qFi1aLaIAJi0bypQOF6orw/Ti64o2peKwUaWbDBe9xaTortiMt3g69
rHnbg8X48b14oVCQNUZ8h+ziOC/MIKve/t0NLtoTqefCfXlYmg0TahWDq/8VM2lt
xr0pNSr1wzHkS8zGKfzH9nXxpFQ1tTNQmf+UvdQj5vbwUzTJ+ZUTaYUKWnAaGOqd
bOz6nZYIZTGofbJtatgk9tu2vAFZYXhEDa2A/PbmtBh2H6CfRJzUJO08iHNPBuHV
nz24Jrrrf+9X0sCxZoMGFjrrFwXPRmOlEJLYDmfeL0YMuiRDNJ37viSARTpueQTz
/2MQp6lpFEtQGWvZMHbMjbNPaC4BWEBrjVkIk/buPxnaAy0bl0uo0QfZ7DPhCtMt
QoKqYRsgFY+jiv1puqOuo+uofMGMWXRlrARinPKQQ+jVaypkNHSvoGE3er/dFb5P
bIuhJ6dTM5QDzUfvgBr/C3bxXIJKfqHt3w6jpsspfOw5Mv2IGyGdJD9TuGytpmN2
lZNZDQleVIDy0/fVLuyquIy4wDHnnsnqdwd8MynvxZhnBV0g/oVXQZ3JjSiF+E9M
OkDAvbrVvMkOtpmG/+jon8pr+20010T3ZH3sAuy89RVKPfMoxKkGC/RRAw8y9C1D
wWemq5i+KXcP2l/dc1lw9TKFdsyuUu8iULCqAwS77HHNmVi14HIS/1iuRurgJsjP
ZpjMoPi4L7b+30Z2CZU5yY/sNdhzzrnb7AVJtD6aJpOVYNkFHUv9kD6I+0bPp406
m62Fnzd3z0zKTXOHjOVy6dU4rCQ7/AOvdZUTqwdFQ3InKVFdKmt/tDzaWTzlZJgU
9DfmFIkyVLepaLcMNAfBBhCV48HS1D6xuzpTfQ4OlX6pWwCIZZs1uDCsgNN0L0kA
VrbrIUc+piRJlXLnp3seG2/ynt+xgTJj6955B/9yeuKum5pq9ll15+Q1hOoZOLYJ
h0lRdKpMZ++btDcSUVTGCeWd9fyFCRD/+Z5JNGsaMdQs77g9qENke7ba3XHhAd+G
80qN4AUIwQzGN86DwQml+E6GwYHh4PAeEfg4WzPut+rLPETzWoAKNQP2wna1Q3p9
uHKaFN9W/rgKZRXJuO6F7bMn3aUvzCik5G/D3nxpTQpZ89YCZ9sLioHTfpDrmjQF
kxRJDx9KBQb2jQQ42z/iWogGBAcrMn02m9Dr8X4SABP/F5AjnQjiG/rQNHk9W9Sz
nwoYUTZK/wWI4Eag4+fdEafykVVqWN5pSqjO+OINjTnJs4oDLW+288iuPhM9PhtU
ILWrJuK/uubQjWXs+jJre5rivZnkPWaWX6AG1B3pqDMlTLDqBkE3ORwOQ7hUsGH+
P5Xt3deoE9r6lVRjoNxpiPCQ6/vSlK1JanZ91KEnJvs6GgQpg4f1rKynBwkAnRJm
atOC8pXZYRDcv9WxwA2DRc3R1JawilI/leCd90Kih83nwBWStudshOvLS52jO5U7
zV/opQ/mcL4aSe6xHSAUUgHTWbCBAF76EBAbRy3MzVwvlGufwZi+6CZCQCMpr0Yz
lEGNi505aIQ/X5XDxY15bvjJC6+YhaZytTgm4H2msCVpC/hbvC90KK8tjyp3uUrN
E6U1YhabU36bNcJKnNZeoRAU4egURKPrHFsSeLnlqGk/kb6NA4Zq4KO84GwBXqmS
02C17cbtn7efrLy4g5TFc+5XYyRmPj0ydtvNPgcjNwODhE9hMJ6uvBDkLMlZFmPU
Xpj6fvFuEtjGTyojmQX+yb+khhdqMVzJtKrJ7PTUMcmDPp2tzz340Gk8NW4M2Qwy
LllC0crYZdUPKtArOUPY4bEw6y4F0DYP4IzCqZI+ZvhyY2U0DvZWYCh8pEFzCbp6
Fzx+ZfCe19l+iRibI+jcNSGZ4Qcnn1dGkJmHrZFQ7oZ2JL3Nff7GG2vgGlH8ORyg
BRDBaDwjOPLTnjEdvaPgZDSThANu0wUV/n40qQSf9yHK5ECdbZcj5P7CT7dzo9VZ
kud3WyGaO7Hpa8oRgrV9GeAL2PBL08E+iIWFRquh2kg/oNZxj/sYY/xeTD+MWdRA
JfQCg5fRLIPuJeUZ8zGB9mgZBkwv4coXWpLKsohYKU4HozaqVPYsxRZE8LKcCTxy
8KDu6yOdHwftBbDlicDdNaM9SYiGc1KN3CMfWqzhD8gbIzrR3fZfcVc4DdAsNurj
N8P9t+wZ1QbNMPjZfWEdlCf8/KIBe+JU4lE6JzCb4ju6OLP6bIgZaM//A+f2+tTD
VHCZE+aOvt0LPHuBFDf9y2ZWHnNzJ+Uo9qyayq4+YmFGSea9YGWCKd60lmcZk9vR
H3ZZ/nPk31sQYleIPhMTiT6Rho6Cu9MeijoBxNWFQEVUY0KLqxqNSbjuaczX40ap
c+IhOrG+lzWbpXQNduel4Yc0IotptT7yXYgMkZBEurNqA43YOMw3+NEwI/KnWfEy
SA1q0zXFzwzULpuLaFmwdZKrJDcPks4Lp4WCm+05sLIttgCA9zhbkaxz0Jtgo9f1
A46vTOnEYr0ejn9eWFTNG4ITtVQhBn0IYchWUKPdLoLgr8SOJVvn8LSvw+esaWtG
oL4iPerbkehYWHkTk87ckPGObS6C9+jQbPP7BsdO1i1JtxOJzqeeW0SpogIhQPqp
uQpyphcu+9yZHe9hUSay5W543Ab63hDQU6HtVtkJnt/ofXvRC3aUd/tqs1s33oJz
dKwwwc0GguZKWzdZezf93LPJEaBqtlyVdkrG5/Eh1Tjbb629KaXISvEM69esqnyr
W8I2VbTANJl0tZz6ZPgrKcH0YdYK3ieNalt+ja3PC9WPUBV63HclLfFimWV+VYNw
c8wAXFe1H1uzGosx3YkxxQrPymdDe/VtEnGg4ShkyjwV+ucE9GPnIKr3HOpzzD4T
8j++pfMBcuXETvBGFZ/SJp34SU8mymFkkl7aKIfKCDXPU0+n+5+LUTmGzBcQccQe
XnqDIeqEwafGobDW5uo0jYo9YarUYYE7/wD5c8UVfQ+p77ZH9u75fja/h1rXd43W
fdV2DbtULduZHbdkLp8O2qkZtyV73voAhEMRT3gWcc6bcy1GpTgbvOa0WSunr+qD
tGt8q2xlktRj7M+mGO4F09qgBHquuqaNjo2jQoZ5684eGP5OQxQ8s9Zx+8Kkbg5h
uFNbyb+AMY1ErHI5bwPrg5S8V1EZumGMElBYFgMFowocm0SK9U0dKY++8ZbvKF2V
HDqZMc8nJSE22UrY4so7WpEfS/WPRQEgazKLUrok8qmDKDyngoH0wYQcY1M2Bdhu
KM3Znx3AreR1SqXVmh1j3oO+4b0rdE2xwUhhMb9SrS/e1Ex5vN3AmuOk1EhJm2w1
oLtTWAMEcV+jEzmNzNLWAiDjrIAXoqc4z5v9F+pO5deaedl60Ki7vEBxtIqSEivH
GOELdzuLrXWyIPQXrfRaqVfcfhnFDiZpEtLSxizzCIbiinOI4dTnOMLz7kpjdA8s
jEfLxNCG+FTwCRZiPvuu4gytjfeJwo/AbxSrupb5HhPRmNhvSQ5rgh/uMju2Tc7U
fScp+LBDkuePKE1O0hbmF+Wr1C4N9mNwMTo1736eUaRRXE4n9PpWKG9BWLz2jpb3
a/WbDlTTw6fY93r1jnuvzzi3y8ywr6aBvfQ/Qu/XHVVc7Dca+PuZWVeWo4EGys9k
fAkqj7XFZvpBX7qJ72Wn/AZG9SxthrJNoTp2ylDCEvkVfccKDm8qKiVpGJMYl67o
CMeh1MStq7UeKjXl1KQkOZxk9wh7VI2Zczi2HNzCk84ELIfj50ohA4yrNrgt9f2Z
F6oxTxqtxRhW9X+m4O1t9fLexa+eBJL6YPMFsRfUvC3Xjxh1j8RPAmoNkF4fSb/P
QYbABfZF5DwUX33kUzB0cRauJTBYysiTttPFuXYKEQMGghFOf8bJ9WRvOIcPqkTd
uYFXHJWQW5Q+uoIWlcjaQH+8bMNxbVlLkfFQ/Ny58UERRWTNphvsvbw6BubIOGtm
cWAytWIWAnaGvsz4bnN39GJvawS6r48VBJJ07Nx3Y6BEjvIB51OPua+IbI6h65vq
+egnmfZ+upCljv+y8iAE3U/kxS2CsuXUpVE0qfHEfoUnycVEoagBl2CSuwVTRM5u
8GzPf1CITz3cBXIdYrdj+E/Sv2SGrFZp/5KddqeWbBhoZaYFWYnrbYkiE0wbbEaw
X3b+0RyDPvzm7vKQTpShh9ZQWr8txSVBTOIeOIDQrx1fTN0GdZkX2IBdLfkbDgoF
kJSMi7c8Lz4xFv7c/RYHuzc/nY+DfYJR4QESBXJE1Jl8jIK3AC1KY8oqpgaYTXTz
c2LiIC9kaFmZ1JcGb6/c/k3zVLml3ztRHnqJDUFcM/4j63e8AUWGTK0wKHBAkpDF
vjg8oJQHS0/TKG6o2wTI+s75KCGfSZ7Rosue3MqQ8Rv1CYFkxw8t0OimxEOcUn7t
MLcM5aCeWS+yLEZokN+pUmFRsB2MIkGTMIsq1MVGa43trWKiP1M7sahlCOQwmxCz
O9rucrZn/DWOelOU28b30/3eBUmiTqGoY16uHC3R7En3ShvA1gzuSqf/GK7qd0qd
Ex/WRxE1OPx98XRy9VXc8KSslMcVrpagd6saYglNY/U30Cpq8zShdS+C/lwOhNyf
07iQ2PA2FVLIJxgvDav5cntKFQ/yiaQlZQBKqkob55cPznM/2vUVLYukc2R/Oz8V
nC5cN+EELJBLCBs//cGvA39WW87ekKFmcNKiqlNXqn7RaJKnPDc8iPgBfjKeju8K
pWtYZZ4J5ljUn4bS8EUiCOyOJpnEhv0DpLgm8fBFEhqjo7TEBdXhkKLgMzNaKGJA
hFNNyEzD0PflXtm+cfydPpLtYH5dLdUlVX0ozx6PWvcqHegyoF212OPbu50E5OQD
yNwDYx/Orun3v1lXuRYJp25MElLc3i+MNC8VstcPAjpFlckWa3/ezDAH5IJes/zn
dKnNaBL4qXtN6kpvUMSIheMYX+GrEx+vNrH2JjXkuTDSGzM/C60E+U8tlje56qdc
NViJg63AVPw+xffy24ZGYADMWQqG/EwtZ35t0ljcbdpjfuh8Qhje8ULoQV7237lW
nUoiAIr1gaTZ6eka1bGzjvVWV3k+rlJMIC2VJznMWtNirQ8OprDf083l61Rd7I3j
cFpTcYbllb8zQd1BogodCO/EHQM22Z94H/uK2wRP6hN1ZEYnGIT2Cxt/0jihc2fj
EWyv4dBKf+z1/RKJWZcbmdzbgQwKQas67csnErMUjvBRDAJbWxEMwQ7gWrn8ovhI
3BVssrTCXVWPcpU612Anc9/VB8IOIj8crjA/DEjjhTKmXwy3Pk4NKp36UcU51Ja6
1e7I+D29Z2qD/eue8xkveIduGs4skOS1qT2z7lAKo1pfzqJB8A+r6jsu+fSccf0W
201OgKfsBdXS36KTDNZg8zykJUeg+lz/PdopxkKc9F056R7UIHwEWuDZix4gKLG3
5ZqPCOlvITqb2hHffUcIc9yFS+uIpi/OhX0PmELH5xQRPxp8wBg2Csysr6/PAs8M
f2zknnSiRV8C5w6Rfyn+SwZmxbCKYZNkMs8p30VQF0J0MMO4Yc49i/+7UzzezDoo
Y8dOtxPwt6yRxVel6ujA1CKQqKLXZ64o22jadaxZVHpInjV3Vgj/sZMTCTGjyjDg
dmvmHs/i2ARLEBad5FMa8exzm5T5cm4EQbIDEVE8sSmnhOH9B5Yes5hRevLQiWnu
TdMIzQqKNVUKm6pqEQ9xaZCdBOsKXJcFqmEIGewCtkuAxvEHr+pAZ2f2MNmkvF9u
jzUw5FUEDC3dkm4O8Y2w6nv5qSK7MLaQiENtCUdWltBoY0iAbz1JqWvYfbkS2JfN
uO8Dt4wE6ZBQQCG/P0Ji936wQkgt7LL5USafK5raoARseN6Gr5ZWghTsBWlHsHxj
/xtNCMjmjT6ydg+5k/TQzTN4EzAVxstxDLTq1FIq3UyaLAK6RjtSdFsOKnPQfEz0
ZwKxfl+wiYaGrBWfs7eoFOKj9CfBH6btF3oM8ELDKmgllyUmAAzr9yfANPhMUSW9
HY8u6V7kNBdFUM40cM3fwjxt45I7ElJ4ONS1aQQcX8RfYsphfs93SN7Q1lc5n9pk
8xHdF6xyEz0zQlmfd6KllD7xE6xJ+4mKeb5ir7LrHekP2gUXBQRw7f9DGikxgwWh
IEopVJQisT8INKcYg0OgVPr7mLaxj1bHCV7RmAz9tZar7pB1iXrTBx2OxTgninoq
6VKZOvnPy3+68OWqCIDWO7c1eUaCdTeLpswXlRkk0xzLLuj5LsaNRPxGAnGPxhQC
zfDEZR9ALUoiMzgUrWTuR0V1M3JWcWxwQ1hqsMtgjqv9KETCJcF/yA32SFfu1qMk
qgykBVX7XILQH+CnraPuG3gmysC3pekc0o3hBdPYCQ4UmiEC38v6w1FwaOmroWrg
SLIB8gk1/eq5ci23qS3n20M3ZpOJypm8kzv/kf4YVpuSTbBdfT83VGbXEIKQXj8n
aNTPQRnKFgXPEcdL6ZSOd353RC6XunsXwnpxeZ4IkL1avotwz2W+u5nuctLwyuw7
xCFhB80YVSn5I+2H4js8pWxXAhlU1ku3zbJaYald/QSMUR6lG73DBDd/byKticV0
I15Co/lQshjBrasrDgo139e3LqYzkGhveW7o2xmIzveVmgeILQZbyykSL9TBHsnh
gSIcZ2NObM5vnTbXTOGtstYxIKs/shwdZC7xJjK+Ho5cDssFiuWU0HZpYbm82Kg7
k66A0n3Lej+cmXPbHfOgu76bavrQnZp8XZgFjzAp42IzMmaSWSXkAocf2aq74TBT
7yW0nxxwmzmZBgirmMLPmQq6TamzkTsZKJWMiFiioO788F6Y3IEH12OEjWLfZ1R+
BR9YncBQHfrkYwaXCR7xg/0cHbqhUa/MX6m8q8dww7tw+lwyBWNDPoGjjLFIDMdv
CVYjEdFCBk8jLMU2aBB+CNqyMhDYQ5/gBdE0EyqCgptHisFVzDNEMutCfiVZ1dve
hCX5YXjruF6tzbdeT12vpGBlTQ4Y3i7FLXWQoLQ0OKp0+AGIfW4jCGB+HwCsJck4
xj2nIMF6KWZnAD4fXCVNHSvtx/+bQfvivHO2oUbS94OVQqUthqTHIitHC6w/dlZI
4ALCTJV2l3PPYJPf7/YJMzlyvhZm3zGgSFqBOoU5iQoFi6qCqaWhC2+aC1YuJr6j
0GPZKTyiADhf+jUUyDGikkBDJx+S+1lr7W3Z73KXzdq12Pi9afxkmXQ2SpxKenIq
VOTPXpo3MQgR3AGjyZ0EbX1Oe9f7t//3JwIoxPt9E3R2RLq1Ze900D2mIup3IZco
bpJOI1Y/2UkCrxfWaBEI/c8cG1veQtFFzJAAmPVm78UFGueszSuhIwZ6r7Dg6Y1p
FnWXB2B04Zi8jjy42JilwMyVmM3g058cANdKiycSalrbaZWLHSed/QjaZXJl/aVC
FjATnIWx1R90O+OMrLIi2uZD6drYWU/3Vwc41E1HEYsS4sbvFTAeP35s72yKxSzj
T+rxHvrUnVIZOQGE7gv547WRsmfQ8rwvwc9hP4+yraJoZgmYJYqxmEDJdSTb/PN5
QejZ/LFVmPJQ2f+6E3mS5OYlGxf8y15gpd4QUBjPPHu5WqhMFsIDrxMehFaczkzP
0iZk0m5qa6bnEkmR30tDO1nyLePeOLT0QtNk/L0S9WShG5HbJ0otKw73dqgLQRcG
DsDh/c8fffKw93crBr1d6lBIESyGRD9r0IbKEPBsehrJFvsZAHQ2+9+0++huWN0a
61dFglULVU51K+A0NTmf2CY6nm8PlxApNMtcUBimGjz8qx9PigQRwHc6LWQfAYzs
4esSrC9WZC7dGkqd5kL8KqxQN7VCD3pG2BjXyT0K5ROb7bbNUN83KOPRLxfl3Fpr
V5etPPtz1LnUnjcma7DfrKh3oMUPmdUweJ+BABwjjTxq/w4So4EcASX0jgrXnPHl
+4L6oVeQHQVIy6k7zVcadqfA3mqDFgn2Q08uwc/5MupcX4f8qQa4h+yqNw/4ZAzj
TiIrMeFBipQNToFf/nC6uE7qUSs7aLbeZw/3s0oj2yxmiDiuDI6nr3Klki0y9nuO
K2hgt2/9kaW9TQZyXeGLAUWOJ1EKYl1MAbce5J/bMmbje3BngCIwuDSA+T+2tUm/
jdciEyp/7v2N1B6K6MCWKXSa8MxvSvkNWTHPH/mV2UCvQ/p3ufJ6PbUekPQlcNid
T1CrAIShGUXlArASLOyEh+HUJpp2OrLXZbhbwd/7E8hy1nOKOaXhxSLGy7JGJX+V
0gHYjJkQe0HkqbCkzO/zSwimqUSrHzgF2E+yORhsxX/o9vBX4KuWDjCi/0VpIaHN
fxqm9PQhNQK7u31o06k0c5BmNcQw+hVMRp3xfdC8/ujcFxDUxqdELxsByZf92yQp
ecQ8DGxmrfzO8YudR3NGCEupiKON97Hzz9EVygdH4b7+j5DjDAwjrquwAmrQOKJT
L7Zn0vJatgmIBaG3Rgvc/kqt+BoapG75GCgUrxw4A+Ij7RhBM5dz1i0WL79H8Quk
3STOhhtN8Dio4jRT9Hw/q/T2HXy920XZaZ/mU1KKfUjDOCX/dSy1SFlVqKWpbm40
t/7m78EygSQBGee8IglmNYLirnT0mQDXe+K7hwE/f4n3KqT34MVEVnpOykr28h7h
wIWMMnbWtOOhCprCmBuFKWLa63LpojHCXcimPIgtlfi/JdGJ4X2IlU+DHpoSpEht
pOs7F0c7nq9kbmi9IoEgogj4bYV90/zb/VApU8K2Z2lpO8DltxrL5MLkNSnxMlUt
wsTH7CwTFB3YHxrO3coAWqiCQbBgDJDAGdZhnVXnAS/IlWonMsVzeFBD3AcbbA+Y
C8lZ1DLu4ERsC2ytfafZkNdI02xVF+3Ea5G21CZNb4NJv7UioUvWvbXPofMF6a/4
mJTpg36KKziZiXXLu3FZgvT7n5/9NiMhPmpF6eUpeI2sY5tP6zDqFIdE8at7cj80
931iiqai1XitEe1SexwCLzwU0P0GebL81zk8OYOxxJgyMyfOzRuyimnAKOSWCAkY
IuzfGpOjZFmVasJBycowuILzR/xUpGr734Rp5K9inpyqgkkEQLl1wVQTprwCHAGd
8aAqoqj7BmgcZqbZyAHBARguANhfx17/SGM/pKKJQbL2dEgoUxoqhTCmuwdPzH0T
b2W1/FB6B48M6z49DMUMM33OO20DRu5FKVECNbCUvIVyX2D3HVGd8Pa+qXV10jDq
LAO1aUXBZCovi/kX/VzXIQLRuANIQN0j9HrNiNWfTH8ct86m5T3bXPdHXwjH/ydk
I09IibfnmvxA9WnE0pKvJgri6wFpPwyjK0hntqnRe6h8q1WNYrqbzFQwn/KB4b+J
95avBKYWWkcwM9bVF2Z8PJBpZJkZxl8Cp9X5b6rvriB0kUwOnkWNYIu+PSOlBBdW
DLnC1rpjabl1WPYXn7XAqMOxxurWj5P8qwOXok7k3mC7dTRbGsyFfldTDYopV60V
Z3Sp/LKlJhgMLyZUu3uZttuWAWdL7ZHpQljpAoOWnjleymbVWm72DpMMuu51VRlz
Q9q+pj1wCTBYp9H3/z7zQ7wGkKvc/m4eTAR4Qfs2DSSjPr8Dka0qWkdQiv04QG/X
fuwX9Y822D2kRbikfWf0BqkGM6qoKfCc1r4Mtyz9lwRHpJV92GZ+ldcT44Oc1LcH
zPHK81pbbHVSz28wL0oRkV5eRcil6iBBLxmLtPrKBqLvRNn7ZRsZKBGLeVQUQP7f
dPdbF9CqFYW4o12GKgv9plfE3ofzU97pGtDOtUuYp4/0xCyAlrls2UeKIqov7R1i
F12NeJeXx9yxYWPSRRjknXDyW8TdZnFf7hvZoxwmmUveTJMfUSfonhdS4uCm5537
GjpwSRfvyZvRso69L4CQUPCyDCyupFiCDa+l2Y82KMKe6QXwW4QTB1mwDVhULMMl
4lNerkbAlvEozaDzqX0hfs0ugISyIWrV/UaGN60zZd63MIhUSpP/m2mcWXOjSQTM
o9tnnNTilEfpabHprObVaGXVwCEnL1KTSJr784ZczKkPyt/1PJmCeBX7EMZsL/FS
NW2T86F/J+GBfHjadxqsN5bAL5v1R3YDPmu9IRfhHRhNRDNPG06/Wrnw6q8XwIV0
JWnRIktztJO9dpT8BMrJ6DEbhV3Mzfrj9ZBsfEJPGbSdGxhD3dmrXkJq2CzPM/5o
CqzstHyw/DPXsBE/Oy3l2M1QwpiiVIHD5n9EJy1Q3FnsYJ6y59E3qIHAuJyZm+eF
iN5cQg+2+bZpmpRpQTtTzhgXXVaPDp2IgGgqRRFVhbZgVk9zdtPsAJhkZCSBA2G3
cXayay+bb4t4m+B8J3vWR3rZua2dTDuat8OWCh9Mm26WNDa5Q75ERwnGNwKl6xOw
BmPgSkZlowypLdPTLPfHUI6347BA+FnrlgrqkeCt1P0GgYzeTX9vMdG/e/w2efWU
Y+CAUr3YIAV6msq76zeXfE9T/p7hhZJKMLtKxA++5zUNxHLstS0m+dSkO7Ox4Sbs
QtOVMYqVlONFLxT7ZFpSftmBTQ7h1JXTdpkH05hwHdEhT0hHGbmXXb/fGOPKcjiB
8r+Ad1bjSjZsVCAGKmyTmWuuLtdxI3wDxJpGJI9Eg+4gqBnyGA+K5nbf2TFbOb3U
h6SY/XEN1CWiuonpCBAtw2ydEYZY59gTNraQuhc2E0/6APZOl3ZoW4OhGHuOBk9i
WGBejbRMaaqXXa4Ntzqz6UDU0V6pksDlyzbxdvsHN/gA3YDUlLvzYPMAb4rjCQ5C
CLO9oJpHcd7kOqLZsmw98X1PgBV27PAdMbknIwwTu6wGn1TiY8Lke0UHquPGFQsb
Icx4sg4+dMb6T+SVAriUKpHAHtgayC3D3lpWemRnNtkuqec9JHLMCXlFOG8ckt1A
SWGloHc6OBy9RXuhVkwAgQwZAmjNEW/3HhW/pKFi1LMffMiWLFJJC1+e6Wtt2LpQ
1amZaTQCZwBIbi2EkschV0tYYt2brUAG18tDDDJ8pBfXdnKj0V1we8wnAlZMDI6G
V5OdC1vaT6H7R7hO6qJKdNBHTg1hWyAPBQaM4ff8AnngT+ws9HDFTSG/QK63vqJm
23ArV1x6cnHdU08xMTNtqCXzn1zLCmyvrOJZWeOoIH9siklyhSLNGaZ+3ZIUb4GD
CcpOU/HjSh1U7ssJC9wq8/B1oUWjPXqYtWsuetVnzo9SJde7Ps2uCE5NbsFPKQQ+
gIbJ5Pjt/HhMcgkFdLM3dQYucZN/yIavEXgu5i7Q9558u4liFGVoMMBI/ceYf8oh
zVdjTmJQXksDyP4yZSKKPVPVFuGZXaKtA2WsI61qcS+CV5/u7lSajD0pY8c6N+qp
oQHMi3fWLHsc0+5gRcvzYTCebS6sTH+s/CztJPLIcRWwxpcwCE5Rl+ZDpcXHjHV3
t6qudvQgTlQRA4/Vxgna8ELyu+vMCr5UntOC7NsKHkEK276YUixwRfSGuFtveWFp
AmHRH5RFpZqh3sk5I1+YHboTb+otNhAXCsGOnEBjreBqv9cuDqofcwqbKHwymPqT
pSh+ZfR9XBMt7xRYmws3TN/i/9hx5Vf6V8yRZiyc0ojd6fdC+gX4btRYbWGquE7v
Q4yITgtiDhBfzMnT5l4jtp29bOPgu2Icps7eArQwDnAyHn9r76erbS7jNzenrWWK
s5an2BSNMHqCuRaUh8PjDbgM3qjWaR4Nb++WLOhkKeohQeb/fd9KYtfdXfy8fMlk
/6+LoTzK+KzUs/A8y4Gm3Hg2LgZV7UJWdCg/rpCxldz+3LI2qMWZj6l9IVzrpttI
bq+QwR4sunorobFQNX6MIWMF1LR8a9hHY5v+f0Xm+eQPYJQXnnHYdxTWSgrLjjR5
u7O9c76CqjUEW7M/+sEIHLCuNfWC2YCP8WJp6DxQOVa8SOEvRwEmDq/7IuqXk46u
ET40jD/CMg1rVBcbamnVkyju9jtSQp+1iY3KEnS3u6BUAhJAFQq+Ov3sLm/y2Szz
nvJu06PU5qpnGOwhTNPA1PxkvN+d5hlKpMfueFtxJ5SFLj7i3q2jVq8GckFN9KQJ
V+YbZ1PSKCVhU+8nLO9Ks7L5GAhHptOuXTR5KybGIDcmNUs8t1HSAhCg0EAOGWvE
QBgMQ9NoHpjBpuJ69U4bxxgC3Yt8yGVFMTMXP6fSws5JiSjBjcjgQEdpldJjR+UO
TiElA4SAwqyDaXV4pfIu9Yqqg8PrwsgjuEeZ+jobp/OeiyxuIVuPRxdUQYu+l3s/
zsniWdJ2XBwrNgQcr8gYqSVfUZL52a0w5P+1ny1C6dO1V8FJ5yvH+pqSzIXP17w+
IYq3tEOQBi7gWzIYLvC43Hf10PHVl8tuVc87XCtClSbiFnmsPWGlONmOpYs0MWxj
NFMk9t60MJRR5kS/mljJ9vhBTQzNdTYqIcS3HiWTPAtp321tNUCaz8vKUlp5hEcA
G7iGc3mhAPxUPoFBMtnbw+0VCK2u5W4Xeh9/xM4rHcjxnk3DVcwZi+AA5wbkWHfm
URQPy7VWn/w3EBhsUZ6NrTaWKZUYws86/80MhBrWGjsYdXf3A7Ms0t3UzAF2RhPO
SYPYJutDIE9p2Y1yDx3kz704UoOKTMkHsxZLGQ5/ws+RN9NakK8kEKOYwjx/h0Tu
Tq4N0cEcycI95gCFf73LCYZH86pJzYTUF65f+14LVIBbS7cjByxP3fqufWjLdi3V
LIhC5jmbUxfD+N2GnBJIG+fmDVUwwbVWVSAx2Onym4Qclg2twtI6fmT9clRxlWci
Dd0SBSkUicxukny9hwBDKO+Q/B12+fhvkkFBwXwoNaFRHI5O4mKGlJwNnQcF+LgV
V+0tCg9x6E0pPAALH0ehPx0wTB3wsBkkx/SFkvDewTA2/CQkA6aw56LiUExCga+y
HHOjXlWnjGzoGqpBrnVmpAQLX3pDbT/LxYFGZA4h0VFrPKvD2XnS/DTDZoaJWuX1
ubWWMuZQ3ka6KJXf2HjtBsfKKoC1oSgmRjcU2771gYEnskHWhNQlljhbn3D/cRdf
1La7zg4+ktegYFEL1i01zu4dfdV1bTFK41Jm/1wg6U9oXAe0dR+O5BHN3ay68qmN
8XUJtx01+5oKoFZ/AtZPSIZS++2bU415tcEk3pWXY5UWYwqTzioLOmlhECbEALgG
mERgLU+w4F6EriCwAko+nfWyLgPNZ8MqOvE4H6xW8K8dughVVT7jmEiAr35/pCg6
lIrcQOJApr95uUn4JvsKQDFRqraSwTI0DWDj2MF9CU8/qV4zeUGaHKVFwHxrvrS7
i5zByaU3WWyJJ4TdnD84G8Yv5x00bZU8yjM5O4GvDIUPkbY4d98pKJO2yAnM9ZT+
xr3eQgiplXzbE/YD63dQ9hBF1lUmyH59DUJIh/ycolGyxhABpck7A9LHGoP1aNSC
qQkXtC1DKRqHpVV7tG9EDsPwkrxxTd/N5G0B2C7Cy9yV29LND7YHDlW3gOy8Hakj
gwvmyZ0wzUWM6aN0x/Sa7Kp5hqwsIRHTfjNd7KPDyqYrCNReYv71ndKcCVwtQuuk
Qyu1TogNhY6WpNZ2Ul9KN1TqgjNUSHwtsdSv5CMdb+9r7210QCdb/vOdtoq3DHCZ
xBxD/pNKmLs/J0RvdNEtiw2JlLGGTOtgMTEXy3GtOeORQXPTMjeXdx+Hh9ZQz+8C
DHLcJ3zm07QQ0iz0Z4Asan5fkhlpQxrbN6Ube0WQSSokGBsMceIs3eOTq9R7gdwx
X/eKwyhmnIy8Txse6OUAvC4KVj0EjA3NTfhupnOwxM/3U5cQqGB3JpBd2V2Sd2Un
BFSvpUAroyjCZIW/cSr+VOwegpalnKl/RNjlUR8lsyhzOGQWZ6XQ3uEg4iySs+8J
DEqu9Ji9cUKtEKSrnTaDfa5reC/iOuI86/fFDfE2gLBztu1WsAWe0aIOW4L6mcyN
cFN7dM49TrAqkXp2gGHfniPKiDWbxCtiSLr+d3ly+ZUcdq93X1xH2WDJR2b/s8jx
E4veXNIWud+ixSxM5UrKGONI2NF0fdOA06VjAFOQGdkBvm6b6IfdH9Ji1bvkDAbG
TRPEQXqQ5bOoT2kncahkgnNf6et2SQ/VhMUnGEFYf6bKQFsC2Z+1nCZEDrDUCOJW
2pKMFT/um6Iebu2/okJ8rs6QnsMPOkMgGcABrYQCpeaItOxhEamcWqFqbhBaitJy
nmaJ/si47KfXfj2U2dJ8ZgJLaoyMRg3Gyg3qyHtk3rRzp/WvOLSHoevQAnjs2Iev
6r4xQ1JIckdVod/wWnxGkOB8qXl3g4CRDnggIAqPqkEhU6aCuK0v+fWr0+CCdSw9
ILJUaouPsMMKPvA5RCy3NMKw0u5ogL61dFH9fFGwO7ZvJ0KMV6ZL9CJADVUL1eyd
AMf/TL9ubBvpreR94WwLMS3B64SXi3890nwgeZ4a6mgWPs54S5MfP279laEE1xdZ
VvKfNhZPzZujZCXzE0NlKKxgMVoivXz+1F78L6Ia01tCH0SzRs7G0W6+0zCoIwi2
dMQgn7VIbmnjTDsUDLhFV6NUyg4U/GvMaf1+tZeUALSKzoaA3i5oYSd5On5dQIYa
Hn4duJ38Dde6PIJVrX2uL5KcFTj6tBJX6LYvkb+rBoWvCrC+z9nnL2WAwFF/oyCr
xTzvIIlRnofcxjy8/Or26sjWuV4da+m/homVQHytB039F3t/nW0/OvW7ROhxgkSQ
RW5AsmJUErkVfcySV+mFtueyaaRmVyzbtmIk2fyEjOe0ovzer+bqvFAs8ivOTZ92
uU87pokkP6OGeMBgmTYmQatZrO9Z+bVnLLq8GGrePiWkXAoBQxcrtQTlDYvQMPcR
QmNL1X4XurstKHcsERTvbQbWdlsoxcPvyj8EqeSg6PRXp7OtY1Pm1FlVOEfDicMV
ea1YSpskzOZA3VjtoQyVi53EKTQgxUgR9vC3ClKWutu7GFu3hYfCApsbb4DNqVQ+
VoG5N5/iHWmZ3ykd9nHBn3uhViqAhklVm+yhN+64IbIJzyvlgYTTNl0Bgj2WU6us
yBqNf/p8fv6pSq4OxaKlT5xG7twB8ctlu4rdHvy6wC7X12Pu5JnF2koNl4CCoSqf
PSr40mVm4riQhqfSM8bzdlx3/Kqi9XiyOB9xorxTNxT8W0vJtdcoIJq5VxdhxQCG
cxywPwYl4qwt7q7bEBUvb7EydePA7tGE34POFXxgXXsnl9SGzI+t0j9Jb5+QAie1
LM+m9sujf5N2tlxSv/fDVtUr77Y6+rTQY2ayGf/xjSsys+Id9d4m4vLSupWOvCi2
ldI4SqFKbX9CZwGw5NV6Oxp3xpZooVmfZkljjMK9ZXzq9wmlErr++LEB8BzIu35i
Fa+ZxMrGOxhJf8HIqJnRIiY9J2kVvO+tAeKAdqe4dzq/Nb3UpyMO0fkr/8LixZGD
76wJo4doZtlLYaNUDGQX4yG/sBVYmz4sjFE8KyO86Cc7WMrxLWqzd/ikGqyWONtt
l7dwXChnRbA/uRzaglWmnioqr5ygBiFLoK3BKR9kVGncA1SesR/CZwbA4mcIuXmo
HGfJN3yyipku3uGvZBKewxe+HSAY6c165yaLz8Y7oA5y1S8oi8E6oTWFDxAsoL5A
dSF6As6ZFtkBcv6jy+MYRED/ikIPrpkkrmMLKVN+1SN4hhnRyTWWb/SsS6aDDR8w
m6peL5dEKqAlD/zzhzhq/hoXTLRaawxR+A7dLEjmr8lI5WbNCHPa7zZNOX+beTk5
b0aE9b0fy/JkcnDAxCZRnKU09ZqrdeIfn6jOu1qUUVmE4L22UA1AzNUDFC/i13jt
XxLFodYj5zzdK1c7P1YtMIWsdNyMT+GL03yi1C60xXA5yKp1oq0XvGNcR3jdLpFl
9Wg+60XP7ODPa28GMWMPE9FBxtBQpp+RkU/RKG0aThY50Xl4asawgjd1B6Fpf4TL
2/9G081Pt9gZ34TXMjH4U1Cnp3AyjSrG0OjiTOFJGaM5E5WTAr3NfmR9b27G2NTh
cUx/EENsDe2QObbsY0aAxI48VGGEm61/erstDmSiyIMwOBRuSyGh4+ngBRn5e+Fo
RWpq/pAFqPaZkfa8YmvZVY/bSie5XbakZjSGnlhi4oGcsp4swSL9sAwKfeyEFTlY
zMhKxTPPE74txmb/mnaTi2dOiisPZFj+pyYiEfJPAfa9v9lYavTm4Es2Fdfmfflo
AKhACqNa5xYO5gbvHag2C7MgMe2KVp48pOPCfAOU04BQM4yQKjLWFyckl3hKL91d
lkuWH7nv+OZyy/8GY9WQU8sRjxSiA7tx9KoLpGUlgAN2dtDlhOeinZVLNkeMcfOB
qOJfzGWs0GjzVa1F2VM7UfvDkQDRH6QfzPmOSpj8PXmrAY5PxyGfuRrxJBVJDg3i
K6IKFBkLjNqi8KwOP4/1zIddQC1orCk82LnE4IitzQorsheJaxbigDLC8RxLESWd
3Uq43PiEAwmNCRAw1YgJFU6msjZwEp2Pu945rj/XFphjGQH+j5uxmKOAjlYc2yQi
xctpvQBDWwasJuGSwBO/c9sf7pyfX2GPUUe+vrARuVrcbQZMlp9/QAQrqWvZwcO3
Jf7GU8tkCtqnjnJ22n2esommZs3dITwShzEh9SFb4B5iRTWYbhrFUCaE6M4nijTv
guOxyhGbA6dtGRbrLnc06x3V6YddRQO/+WaLlg8fL66sP1kfhFN4734dWGlX5Apf
1pj+3/+77IsgkY3JCoQy7RQTKhjdHQOGnqYUx1tQvXhpm07m0RSRwAd3QEVK3Xyt
lMevJpNnbpwU7oSIW2+XS1bP8Cu0AFcBJJTPdAU+eJ+pMwclB8WcUGN/UcRDcbRP
gFMlwwwxQdjsBEa+SNs3vR11jrETWR5bGkJv1GR5kucMQOZqi+6AF7dwE4/ayDXb
lbLQhV5F8YhucVWG+U6PjJL0M3P+2iFO+FChA7MYoUwyGjlA2YnHRfMZ9ZUhu2z1
zyxNGFx8hl27Er68QSgKvLy9XbCD3S0I2eRaOtMM6LIZNnB+H9jF6IeopITjLySU
wy4/7c4+KkImFUZPGqXr3Ng1LG7FkinftDkKMueT8FI+/2+FPH+K52G6b4NVB5iR
p4BODImy1Xvxdz7PpHMdgiXJ6ODCu9rXq4HLwVj6Wa9YD9x4Fp6eEq/SKRSGlR4q
ymxEn3iCYZ5w5ehC6XO6GfK6ZU4F5RNdwLoCpmitYpuAd4OgvNmdr/u1QTSrYGeT
JybOBuPnFsIZc8qYm+hobGICh/bzjvR7sKCQWAARUViikZoGYBbwU+S+fxOOMuLF
H+uXuN28EaoQCYXAqCDGrWWSFLKxDlfTFdhAkapdY8tzEvd619QMNaOMNmD/MJwB
d9VYXaDnpKYb/OP+XOey0+DA2IUFUBUGqbDBpyO1Z70qcdDJMi6/457eUwKhJcGJ
VQMGc5w9M7itEJfRk3DnzEEQqU2ZgNXgxg6JLcm9VbFNB2UAghcVuI0NerBtDuaH
5QNs65XqPHZjHo7L8i6PrgnWPGqEV9YhlKB3NzNDnnebb/nQZUJ69gUyqLx+R4EQ
sSoihUWE6be/xOUTzBPjthe5HPDPdmWMkyE9m/KuUduW3zDxNrUEC7CvYpi7Fl9o
ekWBZjsSzAues7lJQsbutlwyevDdDvy2nIOTSepwiXNtwdaA/IxA6oRLepOG/6b2
pgJ9CFut+PjKi4M9l2Mav/++SqoPzZbjCjOcSSOzY7Qewv+Aun9FtFNayhKXKNAq
YPntxINLUppmQ6hyOSSzIMKWZbdDqqGqW7g2kKRvBRBPKF6zS7ztHz80ryDVPXoi
xM21gK19177u+gI7teUi+PvnSnNuwGxXYX77/cViRlP3MAOpmT8ozuoTkKEeO4hk
5nFiuyJ96+n/yI5dmU5zNwjOQPDJ/cE6o5Zo8e9sZPjWddawErjAJnLii2YOKncX
uyKNBLPwcfJ2hQXnbJy/RCyq725CERIOQM41hLARUfxhyUC0eXDL0UMHyY4VDUzc
BGNlO4Atb2y63KdjaKvTf+3WoFOg0Mn2LPUpP/WBYs2b0LdftT7N8OLGyEAiUn/8
a+ukU7YkTahO/KL5NJmIz76H2pWc1Y31UZ/DqxCOLCJx3owC4hSc2XSx7wqWY169
8uhO+XGp4uN1MRk9Eb9+7p3cZqi4r0tOTpVX7ttw6qEo5J+tf4hoCuHYVRvWmFOP
X5ibjYWptQ3PLJ6NsO2wvqGlZAna6D6MNKASbKZn40fU3SmGBjXGZoLl4QE+G7bg
OEA0MpgNTM3b80ALsE3xkydU1Gq06BSqczebPSrOm3d1JhpjGiso9uuBtR/T+rwV
FP9plpBiTbsLuaaauY54y848npDVL7rIX/EDwcOmipFbvZUQ+nK+Y2KqPwpHpTel
uj3Rg/ASSh0PG3JLGyZ16CDEyy2MjDg41CeEsH7eJ9E1FNFHN1Mrj8jnSSj9gRqk
/1OJms8F+m2WaysSIz34b7wgS+8fDcgnmb4832z3m1muLXQUvgDWmNjLTPEtjSA9
RpHYXpS3DJU2w8i3YSciMecAOahQ5vKOhyLS2XUGlRHGGroQeVeTdJoCptT+QiVE
64kmFilGAJf/d/tflruJHAd+D6yPCqDGrL/0vVddy39548IIs1AzIbjY+5+6wu8G
AKJOat1PUGjluN5aMbVk8+3iCYXONsfHzArT7S/8wT/Hm2lWMZ4k2sDLNVB0y4mZ
3oZ6vA3W26OPH1SisIVzRAX1+794xF8LECc+mqHV0SFHIFEKqVtPMkg0pr67hBTg
ZrYa8vOYFb9yfa1OBM9JehoP5QXIefIzhdHQOFBMHb+EYrImEx6HI7cn/fEenmao
3k6k5ZEu9JoX+ObphzXMKnJD1CEATrsXtkupBb/4gjqpr6zij7AGCKvsLzb5oWlj
eNNeSDu4HxBDiJV3uT+CudDpgTCkpk6ZxppB2laS/Oad0INDXTxdXcfT4SNzvcAL
aM9jx8pSKrJIOeDlF1T7QDnppmcW9CLX9tS7OtUhP/UYKF+1yUaLgl/GSY7sCfYi
ADkPyM806I42qZAxSmMnXmcDRASXJhLQt7T6CpMQYAh9bRjyvpznoTLFtwYjCzfN
AODoYo5dqlprv20oWHLn8FG/7mTF/r8Ph/YH3SrFKiEop2xaduvlqh/3ivwoC7PS
YRSwhvXliMMh2YDXOSF08o3xWzS6BNq9yikBQA4yYaTOc7Os5IJQlZmyTWniQJ9I
bVcpbBWyWE7u4RRvOe+i1vXFFqa8Q8se5rzg/t2BVQxfJpPgvB6ojcL0Gv4S1TJM
frf1kRT2zzscmhvSCpBfCn3H4U6XVBIQQ3USBlsgTdTjdE4CuVN+FEkkKxpbkI3A
UYAV+JYZUi2vEQRGSoGG0fDiSoa1SwZER5TY1Ks4WO0Ad1xI8ll/iq03gEV+i+2H
fM0iZy+Fgudgzt8kcIK+5OFAz1AXGlbmHcMjakHrWdORL8kPs2yjMzf1yxZicjj1
CqyrEjv0sCoPa7zF5GAHhGodvpe0eVqhYZXV5zzPfu4dmCfZSbd821Lf/OuFKt4g
JysN/Hnekyw3vAdmc9DHhG2E4EDnF88gPmPeexD5D610AgvDaTgAnLBtu8kXjaGE
dot+/UwqhjAtybW9lq7fSsSjn9hEgdAqt3x39XPHP8BmboUjtmOeDG/9w8rglJWB
/IDQ50yZl3wTKj7vfNG/z55cqFbBrE/tA2bGMTjqfuf7o1Hco8jVUUnM1uDNNMHN
7WyXqILYr5egdNKd0+/WAo/Boi5kaIoF0ZHi4715aqLVjqDvX9l1YzqXqcDs39/P
Ob28Tlj4ke5cCq3P8PElGf46ArsOLWjYrTPtuvog13lRkOgY45k7Mfupo6ZNEagU
S+SalGmOvLNMpY7EH9biK9jpN5DdOfsgkm8Qw1XEWXCvMK1UkZyizivh39bq5Sz2
8YkF6+3U7iKNzs2a/Tv/VWiA1/4eaXZZjDGwVDka1df+wWuMLeKsiU12o92F37IX
TzD4LxijZ3DmVHaGSVANpdry0aQUDmK6cGKZP10f8/Q05oO7NK4AB3BdlcJ3orRN
cAraG6JvfSVwqxe9MiAuqf83qVaQLdAsvIElArqdrGkjHIKvwLMp77uZk/MSGIdv
Ki9jHBrBxOnpcC4DbMqIXF8b63Enrn39mlthAK7coS/m2eMnoWs8dUI6Zn0LfAEg
GNZ2nlaT3R+b/cZINbVyV91D+RvA1gtuSYZ4BDoz8Po7V+zQczeo1bQxEQRWzjIz
fa0vjt5KZeFc4e8kdHEnu4OYVPIbwjd9VWtj4fgYivdmD3pLCSrUudq2SoxUpfGP
YGwRHXVz3ndqmhhDqqCFH3gYbwljF4IhGLI+skoRFYH/RYR67SJ+CYbtLVGIfTqt
HbyEsxGzNyHhywcCY1pG01s/71FPfQOqS0hh9rCLjgB3RcMdOzw7+++PmkOBzRGV
/FGtuTGOsxw7XTzaXreld/eP7knG9NfZs6cgHs0RClFE/KVBMUSArQ1OM9up4VLW
6EEeXIRgE2EFbdmjA3NWBYh/KQa6GwwM33JV3TRbxELmNGwNNZHqcd3dlg1eoMef
HAj83qAPscoUkqNvbG3gnDNbJhzcn9cjgzE6x2Dqz7AGE84nCNt9ReNaqzEzxYWc
L9p+M5HTHS8GzfzK8RlGubicMbMkGjE2dH2Z7j4OhDhMrOj+kc6UaGc8OnupZom0
0f4ZKw/aM+CmOqY77NWlKF8qQHjw6/8s6q2yuBUPkXoh/EaoIfitx65/KCx2WV6/
OJxkDcOCCVMuiLM/Jtr/K1TZrvgy0SX9vYTMey4DLQTPfMBT22sCPX3Dg+mfTO9o
1yMb5iO5U1UJzIX1fCPEjnsWNUz9Myu6WsW5YdNhtI9XW2re4Dv+0TJDRVC6fe9U
3Po+xDoWpJ+B3NiH5Ocl/UfxFnwqdqbXvN/URFctcDqhsQE7t0P9Tk1mZb9fD+XR
FN4PmKZRHrofe58aWFCXeG3Bui1RvUfoiWbPQiM3UkukUGCofBLo7+dNuaXcvnaD
y8szxdnJr1+nw5BLLPXmEAZlViPtrjAe2l12IPFVxneju9KWegiT74zAFGLwIjLP
9nP3VYhB/fwQM5vuIVJRU6tZTcN1W6PyfG+RVYEflOjKpqLrX1sdR2cKsKaXB/7C
WqGxFuwnkIzc/ddaPC+3XsU78kFfVe2O9ZFXC019vgDR+xrfNriZd+aNQj/DzQvt
HF5HiGfxtPcZAOYJHHlSItrbVkz0LPfS9tIdeleeBafAyD2aSI5Fqn5rYnXd1aAI
1JH2CgufI98k3IwdDXcyyHwljdgpMwmnj+PhGOX/HKQoGkA65kPxfjdp0K8E9H4n
NyHJxFMjYoHvMyHUQK2C5DwnGx/BmvtX/V0cHnf2sEGycRNfJAb+OhDypwnLHuib
fj4tw26KvHGHun6zR/kH+nej4HKAzHl8t3UnRuxMn7PzvvL4QA02qr/WiZGheVo0
UOnSoYPhNOfv6fE8bmRQ9l8XAWcQxjAw3Dt6QIeOGdoFFkv1BvRDjLPLqyI9McGj
sRVQQFfAeQMaMHUoINDa1KZQDpcpQ5fm25+gwVF/A2LgbeMECMh4MKXAFbqX4+39
o7LDyc7VM0skD59FhO9vF2n5HAuVAgPFYcGV6cPkp7GLQIVsfNj+fqKA0/Fgx7bG
16NTjUallurijsjz9y395pMuKBHU2MnMw01odirQfpC3Syvv56O6VLjnhEz+w88M
80lKrVAuOhD8CZBaveqbEaHLv1oeA2kO9LfTpn3mOE6aTbK61N8DkMzSbhh/Yqmc
xYY6xPkguZDYtzWGULu+WMUeAh7sC52FtTwgVJnU35Ohy8VkFreXoiyaGqfDTDA5
KwYI++TsWfz5Cc7lh0VESvUQ3XZd3YF/agQcnUE02F0czJNKx59BFDR1aWu9fKqa
jh2zjz/xjYQvMizP/w6vhsGghmFT/zwj6fRm6E9HAA56oFUGi2YhfHdRr5+CwAW5
SkM069m1+V7ALoeBN02xQ+uG4WOGRA0ZzrSTMfryAQFkGRdv4XXJip6cuTv3dvvg
otax1KNBXHwuL68kaVsTWQB35YLYEE4bwbjUzpDG+iggzvD+EcTVn39ROO7CYDcx
6nGFjikmq3xpdM5dZUnAaGWGsC26sFLaAF65XoRjUzirxlVm5EFddv44jIRyETNL
gjOlDLA3iBLB7x4R/2pSjoTOhFDwyEea2Ztw2dkSpDcZmRuM5ZgB3ueJ419DID8+
NyeCXBMFJE9/zR/shTF4XDaJ0JlRp73vGQXfxKrAVmW4IJV2dgqz0IgSfTbCxBhR
NdIGTadJOBaH0Hr/NRRxcjyQMd8OHRv3g237/Bv9613zmqyRGeKTIbQvAtEyZ7pg
HnfLsqNWZksToNB52MQIJJsRE7Zi3FDqb+trQRE8J/wE6M0+7zw3KArKkG/MkUBV
O4TJzvgGIYYzjvXzGTllbLeOlEwwRECgqE+0Mpc1TOw1sVGwBrr4u9QiGdjd3CdE
Ks8Pa8m5ArVNPlotYei+PVI7mH3CBYjROp3cL1gaFwpv43GQ8GeJku1YPBb2ThVx
1qrOHVhVCCwwLzrE03kPKZR99TcWn56BWDyIkVKss+EkZaxRnyCjczdHFGf5Th82
peHHJqKpWDRWA9gYwY4KasrL2zqJeOqYeEQ5xM3BjDP3gPn0nfUNCngeRu30NE62
2LIEouzFn6+/ouF1jo9bROQU4OtxpwI8NanrmI6AFsqOftT534vp1CmdF1R2uhWe
AhcjuxUllRCKmB7IKOnPTIClLpbgH/LKUp6hMRKNphDg76wa+1qtvwzNmqIECaxO
rW0LgSSOtZoWbSgkGj6FR1Eh3UOaQacigymXHVzR1ojEMYLhh0yrJR6ri0munDxc
xgmIzR9J0k97Rm75IK6v+ocNoBa9iqMT8H1YnCN7Bk3dfpXfDJiFL8xkvoroej9o
MeM1Ir87jGeKi3umddllMpZBiJ3f4W+FSyIb3ZNXVs5/7omHo3UouBS+tWtljQAR
zsw3Jw4aA/a3XjU6FN/MP+sFA9YUvtvl8UqRA+UgwEp4w90IsdVYIxMcZfJ+1Dv+
NnA0tT+bzWFdS5q2Dqfo01bP4+1OpnCWf69aVHxHiQyX8xzmvgcy5GJMifYTWH++
XU4H6m4Teeee+bQs9Y5UGLGVT365CNxhbM13cCz/Gi+9hAVmI+fQOgCgEs+U8jLz
owmSQbdzst+NrV5YQJse6LsRmnwY2SyQih2DiA9VoSQUD0tKC6qE5sWxnG7PAlI9
EtLOKPuDkMDms5qLjI9tvBZrrwdSbhMIkmncWQNMHUJz+2W2f21vJLQAlFdViCoR
J8AbtuwvTS3QT34Vu9hxipi7sFicaCp4zd/5G+xerMptwRyIPSlGnQuVDCBw+ruY
oOqnKp39j310wyTPUclMsYknFZ0QFy8SJJ+Uuvi+h4jyFexauqyAK1G3/vZ7ipkv
sTdHyaph/yeHSn188KBQt8h1coUgKttyEtBRDEoCsOnmrr4NXY6I9XqShmdLjb4K
1Zy6XLv5wRvcUxDhZ/T5b1JBohImjPTgN2d2opCtF9RaUioZJnBn7cjKqYecGmu9
42j0G6EBOiDqrG54y1Be8e9CNGvpfccRYlntzKpVAi2M0BbluRtwjyYfgqH8YeyI
WhST3cbWCNUif9OcH8W1NSvFVaQb2IOr7c4busxN+xm5uRcrk/rf1QXVs8LHSAHP
5vjqOy/v7vFqKzZgYZixhY3h+CrxT3oWi7SMe9Q8etFWuZ5HMCJvnu+zwZdH8l+j
thNyZJIicqaTteOcU0kx+kT/urY1Z6sQ3EJgJr4uS2jdNUaSV0vReC0Ul8wc3QfS
8cNYR5y2K5vy1VE7ply5STMW7+5AzAcwVUmUXSx6ipDZFvNKTswyczCwtLIs203J
A4JGsFXVKaHk+jS1aIIUwEkwVpR3mOJyHbrOqxGzhMz/H2VYio32J21CB2IJXp54
Cr7J6psqXq0CJghR+Fgs7Ubp+CYY0oLno88g6Af+bMnRyLzkhAZwN3+uxwwGamcV
O4dcviS2viwJ4LZjZXMySRrlvKzz76v8V2SQiXL2Lv9kL12morI3/75y6wVfPAkV
jUYmPddG20KW8xiW9EfqqmXvfwo/OEvAZ/IWrxfeJkwg/8MW353e+OQr68dcKa83
k6nTbmiyKoDEn5fWUqx0UkfRFVdTcYbBtwxouXQBp1Yot4Fs3WMN8SjjYunkdaFK
kFGGmhJVGgs0LUYON2Avm+80s1Nn+VJSb9k3lkS29Pog+AxwaDE6YLsd0kebtEWJ
P52YmxP2hEhP9fxN6vKumjW5XkuW5FXQsNAmX4PB4FeAMC5ZXIkLqUYV5bVJAf3L
e53RpQkpUZj61MRXyYpzpk7N4mcNZB4eb0CBqlMAkpn7if/rOKyE0Rs66A2xa1ct
ebgjBbYNtMyagRMRRjWmNzJeT/zf2JTaD7kl+WbINbNPCJUQ2zchVEOOTtti7Wuo
RHCB2WTj2v2EbWiGyUemC+xvSf0/XeMSQu/2CUHRiGbePhgNp0GVrLCiGXz5QDS7
8dC5lTGINGWtRuvwSMg1/tDsxApNMB/jufbKRnliB2IGT7cL4ht4ldyNk5OZrdmN
B58foaBSVFZ3XYxgEiHqlWjfbaWBMpRMbPtDStACkHAoU6BVndiZONKhtjaR2ooo
wbR4YHShzE9TUC1SjVKPCvndRIhuwIgiS7qEPQdMGS4X7L3mEGyLwdqYmFGxygAX
ybsEjv1MURQpTf62fh8c70mLSESr/d5C/LjtUJ8aNTx6a/Nc4xKtXdcrfB+lWrNZ
ZLZJbbAm7LjTtPiwf0S3Q+nBrJJMjUqy7ZLa5HKo/maKB1ALRCEFI6JMqewG6CPS
n3Rtb1ZwMDEY2S2rxaZ3jy3HhvdBi4edVjq5O+cKCel42rgKlFcIxR5LQubyW2uX
NwXiOu23Gx4243TjZXLi3Y5GkStPQfdiDXsV2GDu81UWg8qOFyITHCwpo2S2zS8M
pWUuysNMZVpi3Z5l0XdqkzWJ0EcsJWlZPt9juoXnVhIwFXd5qDcZm6cuJrBEGyAz
6VZ0+SCtBkEVDJMPKVFlIii1Qx9igz0Vgpcl5uhxxdhNylZrEI/BOQZhVnAVrtnb
hf8EGyb+mEUIKx4gtKGU6+OreZHwubF1y5dS5qSw8w5DNz7YVB+D6D7PUNOGTv2B
4opQtsw6tJgi7dssmR2zOljPj6EvsNgDubk6h+r0iNpL5o2S2iLD5OsTaaUUrn/G
T+BL72UCrNPsDSKzgzSuZB1SfYRUvgBkqsgaVCRC3aHVvPBFpkbN0+KQSXpjufF6
2yHQ4gcruK/NDGsVRrCdWkOJCNwzelvr6kDbwga1zn+BTd7vSEMfZ0mkxnx5kuW5
BqXEqvzS1/yEAOt5T43FPfF5Yqe0K2dUFaiCPC9FAuLQZ0bMOBJocge+H/yAUnDv
0N0r/vpY4sUI2shtmGdXus3mRuo356Levd/3b+p+jLPvNIlWBWRVBs+3U7dtRtyO
ETad+X+T0svnovw09AkYkFIlyZJ1r7yW9OPpaR92Md+m+OPfNc0jxOyrvjZxXc4k
fE0koGHAktf6TpHTL51P93Nbcpa/R0lp7EvXLOPxk4O7ftHC9nqoVLc6oEOlyn1G
6rittj0dJqR+ktwWa5XzswGeF/IEEiEEReXdW/5GZr+7BSHYNrScR2tPxpPL9Etb
vqXFJZX3MBX04FiNAS8F69NHdf2m4KYuvnWrem6MazogMgazbNJX2dFXRQ9d9cQn
6j+fyms+JpxD+6CMyu5sfzrIAB3VP4jo/9/N9lcTptf8dmttpuycixCO4oZNOb7N
M0WGWWF7UYUq+E2nwjufwRh9ZCLXnNlcZHnOWlLsgqak29QREcUKle0GaF2u0/1c
r/EjmpTjyI8Z/Dm/lhvZauw/6dw5QxabiM4QB1CpNfJdWTHBlczKi9ZzYNuMHYry
q1r/tht0gFRjPNGolbJlexG3mRq3ZUJe0ArWghl9ppEVvmUf3qUSIKMBhJNwqVf3
KNtWDAEMvmTCEoPO7s8qazyTQnUi+t2VnyD9Qy2IYeGutuLyOM8ujfa6gwCm5tkR
9+ZXSgefCf2BTlvKzR7LeBMzv+XkctPXd5DexFNMFSnaWYPw4yiHGlSbFRoV1Qmt
f29Sq6L1/U1UOj4HUU5RTfqb8qd3JO7KwIUOj3CMggK0m3+BgI1NnL1+OJQUeaf5
JgzrCqQ2ER8llZM8QITytqtFz7gEW27owxYe3GLrHLF1zMILCy/dvVZkwh5VGVq2
kXZpqSaJBBmZ9NNGK8pq3RhIQ4dlkTkQHEIMQu777j61biAd9YAPpemtqU390vsb
WCHfsJK8G29DJVSUOECx/tDp8jedgNUD66IuHg58P5m0PNTyxz+Yyh/H3ub7yaRI
CjRsb47310JnthAyPR1ykcaVf/p92qUWGYLxfCJ9hu9bGENpPUEd+rvlByfU+dX0
K1PC1ez/iZraUdAoGncwJha64OF3W09bOoKrwWAADg5kUSLDnLCno+BoHyFaubwK
llMEN05veCc4HVHOCOOenXbb/Ak4GGSh0CV8bM3vPx11qEmRi79ZuW4kLpudY7g0
ngMeyNc8Bv09ntLiztigAicIqp/QYGbb35Wj2q7dN3vYLtwF5Mjv3aDtP576Esy5
nx6qtcE6srCg0zHEoICCqQ+n8KQoo6GHr6QPO3n4XqzT3VRCFId7gWBWPmWvT7Hs
cJdbAfgnb76kvnUUTtaik2q1sSoY4duj3imikS5DUXy8V6aaUa/7fh3wq+HGujZA
Z0FZm3iwnN19b8eX4j3LlykY/UKZrJlqJU+kMz76jBaKafYr4Hb3puRvEDfbKzty
p+liWvgQRaIOt0BccUkuSD64+Kbm9eyET+rC4nsw0RSW4UwBttW8AxVh0T32XOcF
tnQfQbBQ7sBUOCFeMF4e1LBaIVuIIrTkD6e5wDfBilnBVRJK496//dZZx5uNGXJh
F6DUymAYDmxEWYxRvADpstdVTgQAV22N0pQc003KocdiNtHE21aUkaKb29X68Ujj
P6KJoDfK32Xg2dCTwK1zzd2bu0+CSu+NH/M7txn6IGlbdT9BDZf8dnBs2CDvORo9
dxC4gCJnNbFQBdDOvCecO7AyCIDaWURgRrOJV3TcLZWdXCQ5sA4lf3BDMzeJ9k6G
aUw1cIXIcOWggAjORWFaIz6SUKpAwDX4D5Vg1DSrygJQ5htynienpJ9f+IY+jqxn
OpOZy2mxYgQwd7J4yRSu27y+ln6+yA04HpwyRcxeui6vg8thmwe9DWcnyyeybwLw
QxRmuzL4J8Vf3BU2I2PE2oYR1VmNaWRkWZjiJJfclg/vtWMS6gn1v8kSA3/4+bY6
VK6/HGmIO0dSrXegxKs/JdVVVWRV7kHDmKOFNwACyIXmh3NsUv1TSVFWU4xPbBND
9ZmFoclPjsyZvsY7DAo0+k1IResiLNI+FzLGz0qeV6PyLv6zN7SJ3Li2EQyFB1FB
5YsISBp331lsv/P48XqZblpKorY/9ZRxAe+9YLWgSyhKcihRt6VRSnn9bKjUTWxh
UYyWn04ctVZHaI+PprJi+Wz+6VZJyRfbMgeu3ySUq79r0MW1kHlDnxslzshMZp1A
+Vtd7+AREM3K5cwBjhYU3v1uYwFYmYXfypBQ+gsZT6r1ID1Z1s25v/Hyzy8xnexS
G7AQpzDkoGlnyS3VjWk0M8YnblN3eOXUB5Fg7/sdy483hNbmSzv7fSvsEJ3DmLex
SUBHVloJNsuZcpUdoneEOWES47ZAi14P73hctTGW1rnVxvGdJob01q1B+nqliUwL
w+9HCAAIo6T/ymkUQ0Wn1Rf19Lnzajrng+zrrTIi0KoLdaKNjnzrqD0kp063+71r
kIV23L3gO1UG5Ta4CKkLm5FW8lQUggXhpan7NCj3HkyITPjNdlnZ1j+phoBDMPow
f8VkizwfgwOz11HHN+AhL912wnZ2ndlXjsGas1xyQSxE8TS3qVjzuD+cKoGpsdcN
k89+AhWcup/Ndl2srJFRbkIZfMsLdOBkGMJumOLYoN63TYQEaCDbdLCbWkGVcROx
Oq9BLqtPzs9Gg/MuFeIKdtwJDo7+CSxLFpQ//LAnazJ7DzhXihk5QUBlzv2Yh9FN
92a6RR8rx/riwWUSqjL9oFxD8zvs7e4U05YjTB1SyZQEtA39fwNQw0Yd/h8ZXWfx
6AtM35bdCtXKKYickD9mIobsBv/q3eo/6w869f3t4+XqL+ZIjQM39DcsQ4Akyn5v
CifzjeOwhSHaZTKv2IUycXqTEIITUIcGTNzZtQa8xWAXWu8zYBprf7SqyYNblVXJ
4jj+OcFYOnnRWo+joqAtkpifGZ/29I3URKKVa3lIN4DDOZCUhqrsCoTHTVRlq3bt
xbWVmy9Ox8EdXf6/3JGjpLm2Xadqp6AqDcLhjortqc0MdJunWQAwu2kTZSj54Kl8
r3r7bbMovXIz6r/VLuHCACNXWZ1Hq7hgP9tDDfxQlwSqC8Hcvp6Ol9NVdY/fiUEM
JjXVuBDnyMO8b8A6XD7DE1vmca1k+SFOWvz/IECVVdnFdTH3p7K1THt87BESy6FK
Hu+qHSshrbbV9B+pbsDLsUN7PjR3VQ9BBthhtkQJdP5vRFjxMG28QtTyGf3XWPf7
pmaeGZXc5kqy8Yxw53PA8h4SyxnbZPo/QcQ5hSlkhmf4BPqzz6I950VBko5RoDKz
atJ2jMi4gDEKux0rxcwobPb9WJN9PSIGDauy5n14Zn3z2q1kshMZ382QDs4wUpBf
Eg/bIOsvlvTtJe7FK5+AqC1rogchAbcty/8HEDphH759eutJVOxeBGgMMTfktoMV
Vq7vdfhYeQd1pxytvLLAaTyRAPxP8jUscfiP4mJFlgR/lFkCMBYQ4tomvRy8IPaH
bA6e1j/7v5NNtgirHrjyG1LaTUC5ZLYQjcM1AMgJiklpLFDrWB+5wJdi5J+Q3kni
V6l5Y+hfuAN6EXh/Syh/ERp1ALPHUhMUzX9BMncUvp5xHoI1lmS1llbA1UERyvww
IH4OOep9jpfEJzYJHqg/hgYRy3h73FdEE/HwRy+ojs951OZlVj+TQwlMypuj4Od2
d/2H8M9LnK5NrXM6cEQMRXPoQseYnsLlp93N3k3pbN+c6BF7tnSZkP6Vn/KuWcaw
b6v0bDnBl82rZ2Huuacx5nsNCUDbqqxLphnsjgeFAoGDigHmTuYqE1oneh9Kk/FA
deEH1rnr5fm3LxwWoKXEkJZIWdfArBc37mW+cPQ84GWv/js6mFTwoDx3Rb7ulqu6
O+p/IrzcvrViGjCg8bpb7XpZK74iJa4w/yq7ABhcSxh/09jTXBwZojgx53KDQaIp
xfv1Ct0RC2ej/m+J9SX3KdAHOcJPs3iLvLW5enXlNZ0JN8/+RFZ5aDDh9Z89Kv0r
r90RoDxijK+0OL+/RksDzYlF24Xs80ewE6M83uUsexGNrPDpPP+pqcUsAeFL7o9w
/mCNlhJwmMkRzNLNR5sA0GDqjiIzbliU51fiGvEqob6+zAT1BkMbrb87oxqtO37S
Jm4ZRxzFViu0jM/9baftOHhaK2UHg9cwq2cqIcivJlbO5E3vWBwBf9DAQ9jgZbJD
R/5x4VZ5DGMLm9YSTuG5uenT6K+JqZoY+388sQM8Sgy0BQod/EgvWVaHmQ2u80up
/q8p6741c7PohWLEZ5hHOsm8BxlLAZEAZDdc5Zd7y0H+Kqp5TC8jm3TUbDTNPk6O
qlbCBzC+bCtJYLdt4rXGJG1cCYO9U9QHN6CvTE9zlkK+DfqCxzDYgifeFwBnsYsj
So0o4PZG0AZLc/Vnw3x3SC7y9l4D91Rj2j9B9In8V6in6pvmovgClKYkLhKOPN/d
pxqYryjRRcRz1I0z7XLxWbP1s2OhEks8Cpy5tHLBzKUoYDH+VzmO0VWXJcsW4Po1
RnP3hV4tBRccJAtmz3XDVRidhVnT5GaFsRmosWTKD4BDOvQRO6+rFFpMNCLwboOq
Y73tc8GN65Lq4H1kbepJs2a8XKeDoI5fSPKK+RmB2xChj93g5mhFgf4WR4KWjH3u
uEkUFoQT9yAZhuZIu65B45o00p3Qv2r+iVcc2ZiiocXcCpnT4LloXzmLyOnoTO/X
WODJ9ytZFR4NWG4G+7yHjd+wc1eZjgii7aUj65AGVr4IRWiaI0aHNBkqzDtfpTEV
u4C9Lgrz8NzQVVZs5o1sbyEYKDbHe8FtHRv6llFyZObeEVOv2mVCiOSKuaGj/2+A
w3H/r9MCHREF4E0Vkey7gKRGmP+RXu4UEYAmA0QsT0s/XuiAY4vxowbTUd57Jd+b
GZhtoeS18ipW8uhI3mnUz+tHlGkEXVSVztvT9ir0VCLayHOq6miPbJKwDQN4BUNE
84pXNUk83eMC7lzsHxuleY6o5rmk3z7BWNEt+NNCFxkjPCIidbBSgR9zbGs9B7W5
L8wdNknWrURMlDdOFi3ynmxdtVNLb3425YwALpW96O77k97u4NgYun8RbHtG8xdQ
46sgdUIhExaQzetz1b5qtyoZpsXQU+MsygY4+ueMDpW3i/EB0LcnIPT/QqIReCak
DMY9uTxKpUpLvs71BsOLOXq3IYpFWwGXasY5tjOdw5yGoWNrde45JTZLNYMv2Ciu
fwaV/LXcgS/3rcOn/xqazUAXNDDVkt8lTAdNzdRyUUDgXf+L+LY8SrijbVqpWbXb
8xnvkbxYkRTBJVDvgFk7gdi3rGFdj4mgwWgmE0GrMz9hmUlnB7scNnwGh+YgS7vD
GaBpqCTDP5uz9VKMXeV0riyM7stQv1Uypajxb0hpZXSBrefH5p+FBYkm8GzsAcrx
INUi3q4SXo5Dfr32sSm8fgJyKJu9MBjzEHapm7zDNr5zfDB1QGA5y1tBHzL44tok
U06vwxCpdEzNAkEsiq9OESn91s2JPrT0us9+XntbMcT+zPgisHCf2HZYKaWbeasW
hOOUpwlYmP0RSY9w8ikrJs+mPsmO7Hh+kJ6tJh6qYmc2mW+lCKxheKU7D2tp12x4
+t840ET+E92ZVK/I/1SBo5nu7C2McMFzAR7CMMSzqetvXKJC7NhNgqDuhJVmezKf
Z3lGdhase4LP1iK1A5qzBukreQr16Qr+dLnF+MGDRiLhcsFP0/lW7KDmV7QamICS
yJ9xjUyxu2JPBaSdxmjKa4u238QP9ufzgWeleW33Bg4vg2+0oNjeDt2Tp0KZTw3J
xOY8pqUDF09XnxN522OXei2YhqgCON4FjQiB+oF9xZoSMKxtBo9zWgiXvJXC+VWv
PQcF49a4cDM0XsTpamDuYtc/I/SoVU3PC46Zabtnq+MWW8em+nPby4H/9wEWAZhx
fPklXj6JnrADp83yygmdEeZBpNMKEDoa627Q1Gd7MqE8AB1JCLRQ4zubKZzdDBEi
XEylqI0Nr9p71lVcAcSQPPGmC2lDd+mWhFm0bMQQaqFZxJNx0eyhCooJUfDj50Hi
l0c2uv5SHNcgV4kPqG6P1YzAop/29kf4A30zl3wZKScQ/NxhzI/99j/rBKhXJFOP
t+Ncj/hZICKBxUVHIJ9Q7pIVnaHXq5peBytM+gYHL9xo/v0wOM5MzNKyNGkSBUK8
zq18pqyp5fiS4K0n44oVGgHnILr6mE0gR4FzhsJbv+Q8CsBJRpd/23rsQKajRqv5
oxYd9PiD1tFf4G0f4JWUrvS6Z2/M9RKFWQgEv76J4djvoLP10MIFQ3Whv1ZcGkkh
It7WD8Np+0fUT0FVRxxYwZnxlAmiD1Bu2pE6DZSa7ZEavckJL/n2God7CEcPdBAR
/FLe5axzMepl02ltXnNpDOnRjUyiRVWa7IlU15ddSZ/yHWW+VtbtqtPcQBXhr1qj
C4RAfH1j4FcQ4ysNO1eU3BsQvjmZM7CdYTMzo2g+qZXAMjWM+mWs+48new9NI9yZ
SDXRRfUs0CEaPwq9C6mRQTVo7+0CWju27ABQ9nxHb1NTkINCbcaXu2nOz2fsPtMS
7wX1KntbghPvA0wT1K5sqALOvSrlmj2vnHxKJJwQ4q8xNrhxhlhnBjgAW18+ssK5
MvH+jbflK7AVla3Q4Gwk11GvnB+x8MK1PWjoqprMScktXpxn6F+sr18HUKnOlGqv
C4z+pbT3dp5uI00BATdSXSMcydAEkCUJpQ0QGNQyumzogOHfTrpH9xjNN3loLX6w
hCbC7klZ8j+c4Wfavr78nfJCqdt1554pBIZV3YtRtHkvf9Z/yE4BlYmhphz0y+xJ
BKgbPGn5IYtI2I+OEehoXYUYK1GQy0WK4CQHGeXvc3q7ZNdBTmU62YkRO47mBR1Q
OVsXmTmZDWqVP+DOjbm90lot1M1NL5yoduO26h9ER35toFKmjNRSkTGeJxX74pM8
eJXOqjGzKfx/vc5EucqHRvLbi/qhQ+21iy4Y79Ts33DwOgRlM0Y07p9X0GNaHp7y
3BbzLZRfN0KQAgTvb3U0TB8sNZfVHA4kpmoDRPPXlQ3nU5EPoep0GJp6/NjGbBfw
d0kj/mbybu/D5UFluFwNNsUn7MNNoglHpyYYD7C2Q2rB+oo13GOkxo3PHt+HzswV
qR98NFRD70w+BNem+3CWksJYxERNWs9yCwKTzKZ9XQdttzeUoL/nsCojJ9lZqV+F
OA+zEUkH2pS1r6+aFV6uy2bs+OJdO1fbsHEvVPQ2rwaQ8PpUgWydbqMbt+pSvbHK
jLuMU+gGEn8CxJ14nYLeGLzCGGYhipUeyf6Vk7Ov12CJ4+R2Ca4abWaF26opb48H
/To6Z90Xr69VYjAUnw3OD+Dvd777G9mzJkuZYas9DSkAYEXk2wdBTrEYYi1DNDs2
HN2wAliIboCpucfXB5MjlyIKVTPQ8xMJ+JlaXfr34gitNPh43B6bE1W59Mzt86cH
ARQdl26xcc/J3RiSA5yakFIkKy9q1jMPBq8fdq2bmyJpszLMkojuh7cCGGfkz2i9
r8+Gfonyh9qu3x4Z6lEeC8PqUG8bZBwh0bFh9vQlVF0Mxtlh61T0YLizhkkCeZly
GsyZp1ZtIrZU2YU/h30XsqKqzfFXalwCGyf5GUzhfYxRV67pE03UsQbPtnQmjqqM
XtH3yRYwq82QzASCVK+odjct9aeOAvBVi5S5mCW/CF0DLAyiBGcsDSSn+XiKXiQL
IEHfCrtmTLKdvhCvFpaz/I4qE7pv/E08bWUlUDhrFaaaa4f+euAshKv/hnOBPRaq
ZRAOqvaKpAnY0bDMd0/x50zzDORE6W9NwyYFdC9XjpKQ6FImFwfWIVBxBoow4GAo
0tuPypIcEz2jzYwGGA7mO4dOLNwoCVG5XhtoV1a3zgveQWTx+puPX/SgsArBiDuF
0DRUPab4VvinOck5GHkxJ1CX7N+P443O9cK8u5W3C8ayesh9M3bWBW/kDB7Mqbig
HGrvJ7rKAxs1rIBO3ZyUYFZrc0Cr2RWtvpVninI5ZW4Y8vECI9K7b1cWubs3XbfZ
gQFVUm+Ku0d49cF0PfK5KGWBy0PiQjb3FrQY1QdAVTzepD461HB7oG5GMfmZpI2M
+BsZFM0cHI/zdmgvbRa+gnzRJu37ugY1FF8i1/8VKH7GAA0T9yP3F+/4VWSIUECA
c6EUJfT0uxFponMNc/W6iHU9r8ah4PfGsGzHQGnjfgmXi7rd4LSJgtCSBOq0Jrro
qIx6rl/W/Dg+A3ob7YdBS2ZDjhfBQ4B/1d1X0/tj/N05BLXbMmp5W8D9zablKEt/
WcKO82UANQ4enF7DWADGcAksYIWNEELBFR3xGB6z5PeqOhcCNXyY9ETyda1enwpF
2R6HNaYuPGQ0TpbdrmY8uqfHOHx4oy0cDSmv6xli91PXTF7rtPWBSl25uFLVhTJJ
B0SUVTtrLgyOy8v+r3Fg6JVPG4qcYlUxhbChSlNJ8Od7EmksSV9mGFb0lLmCRVG6
nHtYGSjPPe5eP+v5r2FJaWJVxjUAt53v2VQPVq6LJmyvSMVUQHlbdECPbaPHAtYm
gvwIacGHkwxAZ0upGCt2V+yJSXuJhqKc43DDc3DsOLGltKGFR13Z6Zu/n+Px92Nl
GlkMuiLpzWx4wRfVKUHbDJZx71Ryu6st533v7l96yblv9w7RhVKTI0zOPMDtMR/w
2k8nCPt5iABhnRR0ZkXJE5oTJjeLd/WfKULOINDMjHy0XZ3OHJgEeHv/tvaNNs3W
CP9bem37Qk8oOh/VR3NrODTdP/DjHLSNrXOPpuE8HVItzuAn0YIS35rPPUYr7fFj
yWgpgsTsirHJXCJ7+AaVmMX8aild8foV7X+WVpN8T0cRlyVCgDI/HN8h0iHzudDu
LMazfm4roPz6rRwL9ba7MBylTk5puis71wHtm3MO+ZKOKvNYCnNexUuLpuJ8NKpV
eWEK5vce86svgv8ikV6XQzzbTrthA/8lPqHYTBjQj/m1uN8dzjU5VOYGQKOt6G9T
Qa7JrzT20deAvMmqCS2oB9CyEoUfQuPwQYClySc0WuyqiMQWz5ho8REb/k9y871v
M2/7g2OC36SmqyCNYX4x5N3HkcqI3eVUj/DerMmqlbpCqskZrF0YeWFiWO+R0m7v
6AVihB+ZJ6zXM2Cfkj//tiZBkRrdt7RWAqwBJpoq1EElbDN8T2mA2tfzTK6xl5dt
wg2Ek/vGpIitka+VYWw7RrfEr/DAGk3eB5lgEXampBAWFS67rVQil+dfJTFuhBvr
0SwR8XmIsGR75jdLAQOrYCRr1Sy/CHrsy5V22hFzv1Y4YWU2kgMkC3ABm1G8m/ei
YwnkhpH1kymzgstSUG/ic2/x/0vX5R49BhdFPXQWf8R1hKKZbo7zkcFAFhez/H4w
CzkwggpbblcpwopzEgwopmrXv9KZMh10eXio2VhlsL7iOXRzCLaFWTcZnLRYn5KV
pE8Na5xjwtuh1wYxkCnsvMP+PukrAvJ5aMYqAg7HR6Tiq0gtdQOQvGHxu33e0HEe
+Cyu144wQl1lpmHg1FZyDO+szlbMoggB61alUYfGNQOcJtUNF6Jsswl6jeRiyOxG
mgs6u9ZU40hdyuxfLxBDtT9Jm+TfIIH0ygx/pquzTjLfj273icp/fTdH/skI1ixX
WPlIG6pJzE27fyQF7jYGlizS0K5J7Le9pfHKTqLyJUITo0znT72PJEBtybjOWEs8
E5sD1AGpiMtpycQKg15ofqO0+grkg1R5DqlglhtPFCJhvijq5FTwLvOdbWDmlhXF
jYtzv700tkz+PZJ327KTC3j68LGU2JiZTbxjdaxJwyvcR2Dpl0faKV0jwVKQOUjr
s8IjPtZ3PaupLVSrNdUPyVtRVsDIyt/evTpXJNzdkSqZiD/vPW5MPl8yFruszA32
9ZZAkpX+KVWj/Y9xXtEDzBhtaB4XqoWFTicUOm3y1Pqi49VuDHUyaWanf80acCKz
ne2Nj2G6uJtijNHtBtPo9l3kGbfuz9BZmxbzNDKjmXba4s5tSPCzThrxdOAK1A3B
uwkU8Vc5P6kP+juEy7Q0vSR/t1NcWVzAddA7dhl/+tgoNqZZPyljYT1yXAdMgcaG
/ILFImaS/SvZBkVvlVNggGHLP1hlr5hO9VVGvgGSDex7E5qGxZvDEfSsA3Kaaqgo
rtrZ49B6b9jtW6mPXmB2+Jolh5Sv6K30uwHOM7JOvx93oOx9AJmAT+Lb//NdzGfL
n7afwW3NxfY7+fexDbUjUlnvxiLzQPL7wk1eYdf1eOWYBC9xKDwwS7ug/V2uySvn
N2LXxaRURGCKQlZCSzqojvhoBwNZAotfB+TCpnwCwHGwVYflvQL349RXwcilXNVa
/srPMAC/0wtRv9XY64d46xibQVOIqK5QALoSXxhn+cytsMB1Mj8dlaC5sv5bD37N
HPdJQKb0w9PQE/M4fYpzDHQhH27tElWed9P8ONfZOh8cey/qnnQMaPyIlDg6zvMl
NVf0PreMStx7W0pm8r5eY9PlRlOdxCsu98LLUCmuZJq2pjwb61KKvKo3bZTBVauT
2/ZcPuJm3cm0LO8GNDIKJBu7axM1SjD+0PhM3LnTSPARjtKB+FCZQJck8sCxGDaP
qIQ26yY04x5VATRoq1rIEurCAmKvCOEyd+MvQA2JgVIM4qpCHQDR5G5T1CbAbpYE
4V1FEGGeDqDR0Fv8SLSni+ueTNByxda0w4taEcxSDWm0lFA2Msk8Rv5k+mitf3LL
SCcDxQQvIu7BT/0zzAdaO10Eq3MSNQfbOnMtt1+7BmnAglM6C90zlsJeyfbjL2s6
POE35uD5LMmC5nq8+t0qoaEG5MhH+uYrbhBhDII2fhluN9qN6uHDoK6v3vaohMW4
zJWYA87P4YpM6TRBGYG9yKn4PaJYrJvXqNIlwSS9grVaKQQ1k8X9rngocXOrQLwK
P8IcRSfhsnJydX1MunL/q9eSBMLomy+XWIXxS6i4ncx1oF9RzYxtPQMa472XAAmh
AwFoxTU1MwSpjCZJ9Kf2umBeEeNchITH2DByNejwwL5+2TAE2mVp32y0QSqSVk9G
fRaj121hynFBnrr8PkdWnGLnN4EW7h9DlzMzLMiey74WyBDj5r8WnUgLx3URybfv
2UXNgee9dvh9Tqj2VK7hrUki2COZMG7Sfz+RHV55WrwsiT+n+kiHd5AihC5dYNWc
u46MZVvGxCXGmPIJ86V0eQ0H6dvPu1fADJpnMyEv2/Lk94yCWRHgUsuMCzhDu3K8
3cSke/R33D+I4U0zYEf5oJka1/w/gEK0OaTV1craMfBXRCqkmkNyEwzRVS1yiuGY
yxSg0H076cxoRYcy3s4xwf3RgYEYZwSu6WtJpG/yPkwgsPp01uHcJmIXIbQL8UUB
vQ6aNzr4eyO0URg+HPtj1BjIaaC7EafYdBYO7IZixYfDziizu05r8B2BuSjRpJq8
O+9tmkA8eXbq9oBxfAxeKhBcRwrVd5+tjZqkfYLBGahOA3kb9jNpEnnHl3H/vn5x
N8C0SlHG1AJ5sWDUtwjHorV+4BEaRz7qdYiImJ+iSjAWEbzP4BHSsLev/NEoR4QC
EgM4ijHrxUc47pZkqZ2ErmrtjENJYnaStB2Zo21NtdXMJWIOVSy5/0xceRlRU7Q6
CACSxLVnPDQngNqb17siwyugZEsj4lNyIX3VhIwYBtf9JCEHFR599JBn/39RDC7I
HVv71nOmj2R/4OcfRXJrPh9kVvYJ/aKlb4EEOHRZpBdkn3XQOe2Bsolxlfz5+u1s
+yd2OQP7+OMaPIx80o+Zp7ZafDDQIwHqh4jKjWYhIifx6ggjTRuZC47cmzdCnhSD
IoE/hZN+IUO4/n+LXjw0CF5oCK2UA2oB0Y+8re1NCKgk2O9gXz/q7AHhxddUJg9u
qjAmemhuUHnPjs7Jpymp+t59LYDqzxavrloHrZRsr/QSU107ivB/EbAuXXj+84oC
k4kt5FLjQ4JrCp9hls21j/hYKjkBQqUzVaHoFRhEbc2QKy/m01/jg//LC8MubtOK
V6l4nEf77HRfDgn+iA56f/6P6gU5CcSj4qgtbjrfjv+2KX5gmUufDH8kXOjZmeT3
B60bC0hU4afS0ZeVub5k6nhV0G1Q89h53nVn0d9kCRXtzNvmPNN82r/F1VJbaYBr
uKZIolfWjoEG9+C9vXVkKqlYaJZBAavP9t63zAhcP1Q5kqIhAvsBvCx7JuOFVLys
YXo4kjQsCmR7XXeBHUfuSIPOjpnzAQeWcLLmfUgeY5JsDX7q1tiN6Eqn3Ng6UvqK
YF0ZZnzB9rT3RGEuDjlsVjpXwSo1Kl7THGdYhWVrwZK1BSwR4+dgMeu7wKMxm75+
senP32BK4xhtG88yvweyAcsfUvEIIbX+btqWHex6kw5cyTrTOcaWVH6xyMs7+NU9
kXHjIweSA5roaUcT5I31j/uFpg8impdvdBKsJxvIa1rXA64QMrjt0XXv2qlrj/ZC
2oqxHE/d/5GGwDsL5LXXwBvNl7c+shU5Q+RI8hMbdeEKbMEaXgKs6EnXRq436jg9
2U60qmWWf6fj/SgbXOSKzCDJE2UIIW2Rncb0xsDpK6dBzJaoVUY2yVIMQiQ13Uum
FlWy3n8kiBKcaiwKNINeOuquRT0XIIl+oNz3HIA0kwAQkwC6oo589YcGm+gwxg7V
ttIV4uLkY4chvaq88JVmkSR8Ob0nNT6/e6ZfTl8V5T2RbvMZHDJbZrUwsDn3j1e7
tMn31xcMOJPW/aiXc52tFWb7S9cDkdwc7YtQiMiqkym6qnV3I9JBE1S/MDyAftyo
/5Lq5GECBNTjXsi0In6SeT8F+z2TjM/vYYs8l9dh+OjNtviqt/aHGvbfNA6vaUxQ
c2M8TJR5I2mra1pVfOU/q0ACslNFUpZGFM+gjpx1qWs5ai3lfKBed0aT7esuN7kN
V0rMxvt01FlLbr2T6P4Us+Au+YuqsVgXryWGwLK+UR00ROndzJ0FrHKr6Q/Fel4C
0FXtxUun9sNxAGp5fbk/WV/0OUobB9gQvNsgpyAzUs+mcmBMyQPWu1rIhQ+LCUI1
EgRW1DeioMkBJ5i52Of68I3w7FKzwttFvNeoch1MNaO3imUdJ+powbs0k77DI+pF
bcD3ND3B9VLRiL2DMI6wko3dzsJDCdplxHdecDa2XYw51yaBe3RcGUMLtZ8JM+IQ
wMGiTniinayA+WUbKNSuw4fVN/E6UXZjT5yqPnb41HUjw70YRUTejvAsTMmDX4K1
iOPOeoVKpWYEnn1/xjIHL0VZW9HtHdm2lXtWPCjnalNNcYIzoRhHHctRRSmO0vZQ
uMnqk1mykgy2R35LcSd7HrkxnfSIg5RDZt6noZPI1ZPS9uy+6wsvuvORcLj2Ozeg
zAgst9pkUiQ9tJ1BLFrVz9MpSE2McdWyZ80dyhxpsQIIgBdUr44m+V/co4Ol5JVF
GLSrL8uDT8QS7NQtGnQARD3ojI1JKMT828gwaGWaz2wJhpNaXAfF8y0/2KrwViBb
IqnGImLl8Vow053Zvx2QWmsJYv/huKOmAhQ4PabNQB1blJjCkv62J5lP68UUiuF8
kIxH2lFk5l9QHU12iLn4LEV9cnGx5biNQ3/uGEmqZ3Zhx/TdIibrGYrELaAET/LM
20iZyXWXPLZ3tjxEA0B2qk3LFv8cG3fLOSKP8Rs4NPxFJH62c8sFvhj1cWYrbvsI
jH1DHQd7JcVmwUcm/MYxxoAw5YyK7PieOT9chtWz53Nlq6CdsC8RXNNPP0Tzhx+A
rACowsYuRtsiUJgb6qHCjVsOjc9n8GK7q9h/iVZpo0hCJRGAPF6tG63iiAgW0o8c
lxKJ0wyi0gEohPAFlL1NkFBMfSZ6Rfc2quAdwmSXSgQIaKUHoRcO2riJbyXgZNEU
Kl9KOX5BY8XsS+LRDXHuj+VfGBupIJJIaWBLWrnPCunCWwGvA0FD7PKoiYlX4nA/
SIGuNDDvyQy2T4moWgF86C62t7EnzECtTT4E3yZzIFGWz7CeXbZRz7t5YziW5d5L
MRxmaYa/hp2d4wRJcUMe9thL4vqcgkWJ9vHtajRMlaDpjCL1CszUuLlinRZnGpvF
5u+rVNzXPD/xJGCSDhzjaU5oFIM3zKjDCAkGXTrG1dZeZ7iHkmJrm96LfjruBucD
8/SrFrDv0srA04BKjKvwtFylBT8d6kqZGBon/Fqj7vMoloDZyNX9HGzzTOzK9qUI
bdJMgMzyxav3myoQKKlAO5AbRg1O2mCLm5fhsAJXVvY/tbwOgcqxE2SbUJZdQdTJ
xtvNHUr0c85gl8MpYSFX92zoj2hNXyOW/fBRo4KfB7yWNOBIL3H4nq8TPAwus08f
DPF5He1cPiZVr5SuaNEWNGAQPDM3cQ8XpxbeGyri2TV/C9OFEjWoDqNstuE9dmbo
oWvN+Q8qvnspm+wzl/HhxDrn5zvAvDS/EeU7AAlvlQJ7/TT9IL0jWJH4nCXrzWNa
hOr+NpQlQjuFJeByCTTgeyT+fWN+rP137JZEjaULnrQrR6jTeq97uefbBo2PNYDZ
Rga8nq5+04uNswXgxj5k8hXAOzKxhq6Th5hxLYsuCnmwxnxDqtG6ag7ywQkXE8KW
bdinxXLA/yqM6lu2Qm601PUCzxKJ6/OV4NWTA38G4If4oLv/tLKUUxRDcWYr3Tpz
BO++xTK0t3FqyIgxqYaLSPZpbnNvxfDTSRhA6R5twNAbOLCMWUNOkwx5qAEEkC2c
jmKt6a1UafSJQxee7bN3Kw7hESSgAmMaVkEPSj32CDZqbHPdlezjXWYnq0EL6QAc
daoTF/JzXYTHjicgiZbG4mOG8s/9ibSECe9C7UxZ3NBBKs4hhlBX+fsgsLcdWBc0
l5XaK8upDi3JdoHeT8/ziOa71BegM43VJ709GMHFoYCM52YgvnPZrt0V0M09NMw9
LBPpalVD84JQhntjbB20Kj+J/hqlRKh4UV5TneH2m2A11wBAtROTyFsB9N++Q4Rj
ISKfjzUkR8q5pBob6mX+Qn7evTt0UkijB20HYgRcCrunDDEAsWNOFiB+0pgpgTzo
r7SSXWzKFFq+pcKOze26EXLZNbfh4W89xpWDHT79mXGnPjk1ChSmGOGgWJo0vTqJ
htfRTvvIRkWgL/76ZKOYTs3DssyMqQc/sKKkXZ82MAwrCFEFWrb6r10UcWO5kjnj
WXCnGWeENgRDPd5tWyDKJmHfRBZGuAL3/c4muOBXYsfsFbuB2GKidBODtALAfE8F
tl+s7p1M7x+dxdLQxIjFKLdczvr+cfssNHoAIsQUAhE7vEWd2CkVg/9ntn8ODrKd
qwI17lUGzSpxnqL1SCMPVk1wMutFO9xAYhOIPo7eEJDzECRumBc7tCWYM/CXlEn1
a0+BxlAcNlcJMeddZd9ymB3eSqhIbuy6xQiH+x3zAh+VzgX00moy4DHSYdPivURg
/WqXemvXILqcGcbRPC3g75Mbf1Gg5DbGSpO6NkTkTSRN1+VMOtxYLkTYgwZsU4Ce
odszCOXCp1ajC4caeRXnCgq3BNHMpscOTIvcGTYjaBTOBsbgM4ecoIoc9CC6rdJH
wSCB4mzrbkGxSbIbjSVYbMVJqqneSjNQS2lFWecNRs+dT8NFBXmrmRAztef5sC9h
M7REyXl4DOoChhr1gK6L8PcwOYWNJiiCV1oIWaNGp1P5HupCuQ85QY+PgLl7K5Fw
cWiROszItO8ngVCcK3lyrN42k52WZ1O5xCCejfijtaWev1pjHK6M8ejdwAdJZzzy
ZzrczS+HyiEgzDUFneMrcRJjoVfUbY2EFvA3yMpY9nZgQ7BOphWiQhAiNcNs6U1t
XmI/ZkTL9KE9d7vkl8VviZ8DHdslOH4jRGTiISFRcrXtUzBRz7xBlvOWeUSpucNf
i4FA5Hp+dOZi9QZkbwwSGz2m9y+L3f9cSIX4IFabSywp4g0Z0cTA14kMLAKqp4VI
4jcFyscMsEVfqZOz3gV+DSpFIvCQ1IuVmBTOW5tTRMwIK3G8erfiAswj7mOB7Fwu
X5sE0hrkjYdJnWuINiDpGdqQxEDXTm1UncbXYsdLr+oSmDPmvigTxpZTzmZGtWTF
btdAx2kC8KfQTkHjtnptPmjAauFMVZAe3VGySuRxa2bhggIYCj2rAXOAgnN0Xhlc
eUfkDclAPReEctqKpBr0bnxEHD1JlGGZUiZFg2BipzsajyPJ0hDoE50VaTmR8rBS
Fcbk6BVPU8FL5P8RbAxXatEWI2Zm5RCONkSfAm2Yk8UQHkpVlxltfOBgyxZB1gvE
eDH1Fb5ClbMiCOiBYJQ7XLmma+BSZLx/li6MK7aVW701gZvfyXe9w7cj4A5tAoWK
9YctDifw823lQD/bYVwDpmXi3P0H8eSzm60B04CM/kd+YE1sP1mkjZYK7jXus4RO
MzuyJQR0cGVlQcNoadpx22wPRKPMjghswaTZ5thPoPv/+gQAj1SWEbo9Ocr9fijh
nn+NuOjCpW7y5CV3MirMgf0PcZtR1Vhw60uILUt9zlr9lQA/VZZEQuHYZuT4CXQ8
VnMxJqVztxDGKyIkLoBzl6M0k84HWdnazdqwg7cDioHRpUZjAz4ou5U43KDTKzBt
OgFd4sFQg6rU9lJQAbzUI9cKVfAJC7xOyw1xRXweYTf78CIcMqNbgIISiT1eiLNm
Vt1LrQXaPQDJnSy54PMyzSO4JFt8mIyWxnEI1sVgdL0UjKWeLksGGOTn8czFH4n2
5JBMeleP5NbTaoAygem+U5Dznh2xyzLCROY3535fEEERBqoYOZ05/d2KLMmwTWzl
zFtvykQg08eFApYh+0N9ZdSc/6I5f/GD+bUpnWUzg4nh+GsEeh/I9AB4WezTHFZI
EUqbVYRb8zZopu1o/fyd6UWzLP6slPo5je5lkzMxYNhKwOmo673Prqx11gHWEpzQ
8Y6osBjtALaJFeRXdrFGKgQ4CMxiU7HCKrVyeOmsR4psKF7bD5nqbCVV2uNtGjrp
B4xWvGT51lD6jdEQez9FIYDPb6YnNO8ZRtMsfSg73GckoILAMVCIlNmh67i6AhYr
9SWRMU28fM8o/UcIeEjxUFusI2LXOUvtlfnMXSR6hiVmwy/m7hsKXCItqLGIHWc6
7SG0XsBn0ZgrKgFi8D04peDUMKgSV4bplSyaArj70yiOqR7hAu7CzeByJJMPQd6n
3UifSOUAyr5pxeavfzUZeKjc82zmY2HBAMUo9czfMB3XQBBUvUv6Xk9K+NgN0upG
ZAn4dZb9SZq4wD05wg0Bghrk5KjpWF1xVDgr04GYBUSVZ4uEQQOWp537YYZ6vTQa
mN2nyb1oWCVkQIT63N4I4+jnOf5sLR8h+oX3gjakKwHKUnMSRmVAP7BrDgVoErvO
u4SBLz56H3SaTQAcM3q4U0uBGF25Qae6q8/iDTR21SzRCGu77rhUwXb9EO55kVbi
hr+pfcN6WDi9zCcpskQt0Svkc+kVgB4F6+QgZ/begvhrDtgeaI3TF58LiCfGf895
NMFJ3c+Un+gxW9F7RF32gP2cTk98sr7LytOLqG7thMKwyWHVmHG7wVq/D34e/Vii
sK6ELiGuCWFUv6sk7gPcRAf+Jj8g6G5Z38Bw6GdaO+L+QozWAwcqQsK2oxBpuXS4
gIIP5F+DVBK0BOo56QQsLUYL5o9DR5kz3dQ8p3pSzUXVuvQD0kLsfY4wDGzsYn8c
FFLt4ocHE82cO8hPxeEesyNeWQLj3gCHUJXHjdi8/vrY9arIMz1Fi0xcriDB91vR
A+cYo0tji4M3zB0l+19JSTHgtdOEvZiKbzrPbxmL4mdrTJBDg+NZdijnNb02mYMD
42XF4jH6f+q7UBkhaWWO57v/jn9ce4zE6jMZ6SbnB3NRaikUjJspRw3/7daGXaDE
/MjfocXoX2nUlTfmKZHr47TfZpkeIY+PbnxPTaSUTFiPsJ88VEnuVkmihd3DbW6G
BYbsoTUwMF3KrwfWkb3xJwXSWdN8XGAK8flb/JbXKKqtYg0DPWbTnd/Z/sF9C3/z
p25sWzFvjd+TRwjJAswC0aPMGgbIXNi3WVw34NJ+ZtUtfOsbjeRkpHcwODjejUY7
6889INCYEzR7axSTuiwsYY8q1mWDzo6bCe6SV4LcsBDmZ6H8PfbF1IOunhA7Oplj
Ucp/Z0O6MWDFj7Z/NL1KhII+gouu1/+y92fPwvoudyfV3Ejpgs6IYpK47o8zgJCX
GrW3ztvL5rlI/8wrESPfpmkC+E6odrB7Kkx1GF29OOhjlV/Xif1yPVyg/CUWIYWT
yDDbDpw/Nr9SGsZrksrrSqd4HQOjc4sgspLo0+A1zyhFu5c/pobfQ+urgGAcO+i8
QrBrfFRuzpJZfBJF7WPk4gx0O30KKKWlR20ykp0H63T5gjIheHvosyIpLpYd9zMq
K0EiWvCMMuzL99if/gzOUQTI3G8KApuP5T98mGN7rNi0FKHvDWUEnq/xaF50MrFU
9e9oxXq93d6T7VMvFzWJiddwT6ZKN0Luud8ZyeH5xQjxBgXBSyN4rg+WbQyAIY0W
JQCIx+YLDaQjBuj1Lzn6MhTZYIY5mJ70shR3eBigHLT1Lu+1surgzJ7BOUQkQ7Nn
W1961LKUeDGLp2XKPss5fbmYx+BskxcfjYAsuELbjYpyHpbk0SCjrqvKYKFUxxTW
a5JJJ4eEf+n2OI6B6nxV6ox0vtq/vGUoIkktm5nnUVNgivXfrCXdJXCQBCDIthOm
xS7SsNLGwU6onySKhhrQq3X79mSbj1KKCo2uUgRsNil9hC3b/TqLBVjDzB7p/8Qn
B+wmj1TDD/Dt1/BPfHsUAATIZiz0zWxA0FSz7NYdoGxNquVlTwg2DAR4w6gYiAcc
zDFBvE+Om2b/a0sqdexq8wAT2wJOE7PnxARzoJkugUkFYm0xOrJPW7cFk5o0ULxl
fXstbkCyAXBC2P8Lw/pFBwN6rRv/OZyMdPb86R7W91GVVPL7CVuBJt8Lwek+kPSH
Zis46Yd1UxcjADytIIdbHkchRrf0MYH8/JhQzSOM3iqVPnsCKWzUHAdUhbnj/04p
1BZVCSX0Icevu/ZpBgkNQ/CW41oe2a/MISLVbtmUUBHJr8XSkQ/Pwn2cLgzeXvd0
Ym0y4U+MEu3aJAUoK35cXZlDLR++6/cBh9V4Gs1l6ASCPPmpH2iUuQIWYotm9vst
yzBszgGuWYftGjVA8yLsYLt2VIWR8FumJUGhxZi83qEXCIaIPBPcNEPglJlpyqE8
WJvXWgGF0JHP33dyINLDfIWMYZuNO0/3va8XBry3a0ijGq6l9nG2PL8hypH8tqZ9
g38zlgcw6wWrUBKGL57glivqRvQ4naj42jsLtOPVTI+S3S5r91ZYFwJgew7+lonH
X+Xhy16k+bYLvequFV8kTTKxg5WLt1cv5QvZZuXIWFsr5JIu5JyJnxJdpdiUapeU
ZXTlHPgzCiymm+NQ/KB9PsOtRYhYbtj9SScQFwZ/I9k9nptE7QK3Io14cRhEfPl7
rY/agNfkkQeG01SIDxH1uFJ0Zj8hyCViT6szO/Hiabuw4LqDrJQkiZ4/jXFV6SW1
reBK7ZA0YGX37NYPvMxJ3K97bXTOYxYXEUXftnrbdi/4gtDJyPmEH7oJCggktkUL
0PTHzRL08hUeHBC9nOGbIGXEhoApeqN8ZoywMBiYYM0GgUXAlc3V1M6NHczFwnIH
tK2gKvNLvKbd1veEJS30KpY56cJqeAegniHpWc+xYQbvZhOsHN1g3OHoaVshevf+
DG7GcTLaVXd0FJL19hd3ex2aDcs+TeqSKrtH8m+wqh3Yg3YYL0CCVOrF9vMbeKOe
3qVWtyyM3nC/tH4/6jGn7J2pULrTQ9BE9uLQgmyGrcvc6vLBAzeZnha8hRPVQoz5
IJe+XP4UrPAKIpzFJ8NEoMWRFom0NyOfYuS8Rhs+s7ZY9nSjRnMUiSZWGjXxDVMh
6JbgOGNFF2AyvtY79/QZ2ZHdzctrOKk2fTdQUAaL+i6tBNgrViAWWsQqcbisE7jR
itQy7VeLvoOTFVnwfQ9q/lLYLumzby/Dfhq9g1gfwgD51WCAhIL28XmFs2ctj1Ku
E8mS1wcZhV7zXi1AsrvF7gOp2+i4wYAsIu//vUoJJEb8ySv8SpPY2zsqMSjNLvvC
FL7DbpOk9zLiOt/ZSfeo6AGsDIe2TFYfYHuYIWwCa7XYfTT4HI2A1ShrPvtRV6Iu
ZDCXwBF+Q00vknvOAuLPOWpCSC53a8xtwnIebiT++C63eLoJB1t5eYzDfmYDx2vB
PbDmKyDFd801MhYVGvjNGMPNlcx6g2xsO+3rISi5L18Vt894c+cijAF3NrfO++9W
oKrf/HLJP77Z3+0G9nlZDk4KmPzJg7YQTWmLjMiY1h4W4yen9wswjeU4cxjDeLMa
DiY+soeUabfNi+ee8+VPCryaIUFi7w/XnMm5vgcs+S1COMCfNcesRiHCmadlHdaJ
9hKvVBP/uqHF8UpfqCaObBRZ/xGafbGeYSPbnegRR4VotyO6qdppylbwGbjuZZfZ
mnWQRNkxxJrNXAcB2DkpTRTqb4yqChpmEV5PcD3orbmyJ/BtY5I/BOBja71vJJDU
Li9I1C1HWQ9TdDs1oEitGySEt57wnEnt0IWElXhnKf8Dm1xIn8CUDyWu8WdM2cft
DIFxWnBy0Qp+gT5T9/66Qd5jJy4cscb0j+s7BTqkRjRi2h6fillySzIjfkWnIHq8
OOjjoxwCKZ9AoazgIVwI8HwCH88AVVMi0jPFtzW8bsP6NwADKexJMbYXeMMw/0kf
3/4HlBWVmRgDokNvsHvwBOGGMqLiqeWum1KnF0u/Odj6ZSAH+YdEhGWnHmvlnC/x
dNs/a6rKWpKuG5h0vtUkEBBnS2VKr6bb68wkAEBP+JDyT7hiqiXI1TSoOjdH49rW
D5kTMAqJqoTWNYu6Z5LWi04wyrYizB0pxjAv6Yk4ebaIMj+8tLsPe+9Ese+uoThA
EN3NJnkshK3ICNj4ro6EQEf2aS87KaIRu+NaCbRCPu3Js+zH79ME8NqbLrKSxNDy
ilBytrbwWRXQIGr9F+KNm2Bnz65RXCSEob4cD2B8QOUIhWgMuQZGEkBw4rSaYaKv
In1uv5d7jW6RsnY9wrvYQmnMKzUuXfsirdFfvCCKHePqZAxJAnvxGg7ghq0AHxYv
akrvmEEYD6+oe+/JJTJ4fQkz4hYFtgDDQn71IX9D6XGunEyIoxxJE9g6KCl4lLPD
CMvyxTvWIICFnDi/RbVUW1VhxPkKamK489Fqz3SmpZCxucLmBYY+zMlXB6K2pi8K
d7CPym/x4ie6QusldWlyD7pUObe55RhQcIqGX4TN7bM5NMpNqB6kY8vSKxxEVdKb
xL/IZ6Aty4OediOhp99TCyfSjluEZLAGtArx3J6yKy0zopYWSrpfP/14XCMZ2dDr
iqEnxPmPJfoHVgrxKSv0WJ03TA76Pav6U7Gd16a2Q1ZqCj6gsd2cmgxyCHpxl+bE
51MFm/2i3gmhJ6aI6KtehbS3GDB9wzdZYgpxbl+oCN+tege5Ws0Y7mmE22SXdyN/
HeN+ve6gdKHfoQHBPCaM5oC6Itwdyt+FmvrEgeKdrW5Jf/GrvQw49tLu9HNfpkup
kzkV950k9LwtWI/yA3Q1PJEMXqA3gwh8iTgpg5ykxaF+Mt6gszy3FLBlTraPVKyP
7+SWyx5nxfym+JVEHVT8Y+4EoqkXDt8InvjfzIBGAPuaTqt9O1cvVdWQTwZ58+NO
OgdYYjd0w+nAmW7iEW66Ip4Wh7cfJqbSqv6l1I55EYzGM3jjDCJG5xdclKGZRc5q
igak2dOS1iF4GBvFBnaBbEfHTMyRsXtmJu5XtbnfP7HsNPjTQDLOhuIRqvPlfXyv
QSK00+pUXIUh5zr4ucYM2klvlQIMQ0p3npGuQCftFRS4kY9AVtoomq7aEBUrlypc
wUCcyLq8n2Ze4XDiiLcwfsym7jEwRwYp9WZQG8SZ+WZG94qFxj6myIZG9BUruMiB
b2DRJx9cp08y0+SYS63KGRzVtRHFYkKVj345RSWCDea56XHQMFGmqj3aWhSfswG0
Rwo8KiDR5JuLcKcK2CAnh9LxYPGAsDl0fXkohdBVy4NM3jOAZ/ssoG+Fys4/eAQY
qmz82i5A3ChjmDcTB8qJ3qeAYRXKiP+bjef35x1Q3cZYiT4I+ayHM+IHlSVtTImn
+Qg7IWyZmMc6kCqckZ6n8308Dc65d0t1FN/rJ7bV56UwoMKh6MhOlC08bsPgsnkQ
jDMIiJKMisdUOZV2tzt8IPjrGZSTiiazJHDlVAHANSGIc/54B5oN5BSEdk1RImN5
Kmnrmohl5aTHZJTm5OU/4AoPPakfelAYFT5LC+jwOcO2y2zsKPwZZyZTgn6dP2YL
z6HeTAy1kEAqpHKZxJodtUzqb31Yj+iUsr17YxZg3dXsl1scha4iOdn7TV+7OOUI
8C6B/tPz3cwwNmc5O/L0L+ef/1EeXKJvHCYPAZ9WOSFIxULBDCotttVbyp6n9/5p
Zt+Q3NIjZqcnR7ZNRPysGEz4Kk4f1UgKivNt65L1IMTXmJrGvBONfs7A1JqK4HH7
4yvs/UdHwy2BUeIocJynIK/lvbxgdmUFYxn4WudTfNWhxTnit4FEeaMb99f85FyZ
AD6nN+nGCt10R3dA+VfFg22Dx9706gRq3eABPsILcYGKfCvtEBkij9li/7/wSWGm
9XLD4lHFNTebT2rwBaI5Eaxi5jSmoOcFgsYv0L6NScGLmGzkrmEXS2cWl39rT8Do
+VXAuyp030+B4dvPv9CNRZrz0exQPy8HKpbFRTScZ3w0y95WuM0oSdFhkDr2FCWf
BbhfEDYe8zJ9o6oI5IJxIsQnRPi28Hfkof2cPgavyJbkE/5rAJz2rx9XQQr62mSN
zWGpw6dwMlXmGHao9ufHoP0goNhGM5drx2KnHaDBCvUXmsIN3Kod59h8pk6QEill
WNAEECcU71t+5ey0JERH0Ze0DaIKqCKeYjxpl2ieaAuxlgqcLWz41pyJwW9EGjsJ
7FfxyfvPmxHjzi2G41M/OhyRh1xKZs9eABn2xKSLvyWV8fx4Fn2/6VocrqFw/y2A
oKdjNsidMrmvswiFXUjGhC9YfbRlQZVMjOz7DzRWNrVsTomq2i3zwctHgO7IYWAO
3bVKSHKM5AyhBzw5MbIITv730ftoOTUG/sB9x85eu8oBSLGhn13H+Z3NicfrG7Fr
09A2pDwdupKm6C+5xqoXtwuhNOaAWN1WKcawaQXR6ArxRuBBtL6g5RkJ0KRylewm
lflaHvI/LBukll13bpO6lMekhgBn0aI3RJqk0vf0w2t/XX6EH5096/jedStn6vUl
WBDQhEjKsSD++QJ+I0tHm7lGNcsdzQaeJUgtVNIP69n8WDthUi45RjWDV/HSh5MU
9pSUs7QrMRzQ7hv+Dk2z3dRNaiaF37ztYCMLz9XPeAAo78qHJdiaRTB8DlcwejCs
R/3gjZzxZsw1As6Nt/jbs7pB4lW4N38TPRXGIUXpqi8F+LKtf0BbkAFDGXXmJ398
n1tt/z03OMguVKFG93KyrjTtcb86UJ3ADVTx1wlXIbt8iUpzy2223l13nEjIe/8z
2vEFVhsL/REeYh3wt/CXqU66YKtXH2GZyV0T2SeyS8RuZG25bvsBswDMdMqZEo6E
b4uojfM2GgayZdD8uKSm3qHyG7IrgBFQJ1RDw9cJGU5sHXoaw+FYpYfTuWj1hKxB
pRsj6tHVEpSPv9nOtFVNv7Nsf+pFWKuyxOASFkxlVjlC6y/MtvhZqz2iPmJHggjW
bLIZnkDniCHS8zS/r8V40925nEdb2DLOUA/LfyHuqmVWZTqRklfshLnoI6p7K0sA
kqSE+d31wcLyahcpeDu5iGCRNWTCfCVe6/2r03R+lQYYQfXAnuUU2iBBCTdJ/2G2
n3/OwAjqBjg9HuT5heduwvWwm+05xCpoIV0sMtPGDFv042Nf7t+FE2RPi3UrJpB+
r2uKHgNDUNwMrdCK7O8+zc27jqvu13n5CsgSCExlUfzlKMEteDw8ePGtmnjFw91M
HTmiHBdZkD50owDxGxGh6R6NUjcsb2HQY6qUoO37I2gpzsmlnOUnNEGz6BMUuU63
KEmFeBj0ZPtvJelkyFNB5fM/lITQNgUhTwIfl5TMus6xZ1sd0obAmxpPhxxgCkes
dpEopK/8dL93a2nxPqowLdcbbeJpqOalwNji2nLgGfsTe7m1LUa9h8tgaGG2JCCG
VKpJUlRfNC/MC2MblmJBvUYsoUMX1IIgFqLQdMfXQwGQgBleo4RBMBKwg66VN8Lk
ONBlDQky87pb1+sT2tdnEmRm7YqEwbcOmoiAfSsUgbvyjpnqopZWJ62Zdn+x5nI7
UKo7ZMFi12UONm/kl7bT/4MpudFOMEVOMn6hSrQGEameqmPc9bYSjpaNtHMMiOkJ
jnU+f6U9O8ZwolmNghZ7pV+QJ1CnV5RVyixmKZTjS5zxtM+zEC8bRUkZCtf4bI7Z
OGith8bcBj601+DrkQalDkNaHw5Wk5lMeyHnAvWXLmBkwh6SYeE03IOLn3V0bptM
evFG3Ik2CnUMDaeJuSAQapcBQj3RlPidVNtCVZZk4juQtpnRKsPvRWpFj1Mu7hQX
d3PM3ACGlKNLLXskzibI3584NrcYeHc7mbZtrE1xWCmbSieFgeWq10+RLFaZ7Gay
InzT7PAt054Py7/aeAwP2L5RGLdwZ8zetxClfG2KSEs2BtHW8ZFSnLP0722i3Wy0
7T52Bk25hp4ZQEQmggn9/KAU8lluZZwfvlnbM1Y+vZmVIpQ1t/xVql0EB1Xn6pxu
tNXLVSGaKsTCnFJn7BhlOcb6lWiX5M9ku1pFbsgP1ZW3sK9siqspa9a6lsebroWo
m4dHdBaQUNVbyVaTCsLfCSIta8zBDnO45ek3Ppvg9SDpHcy6YmYUnmNlVxpj+o/8
z0kFpaiYsQI0GNxOxLM5APc7r0PZ56uXfiUy59uF2yB9XyniJRYkb3QRJ61sO6NJ
ClU9OEtgEglMG8Z11eyvrgJa/AW+Tgv7iFuD0Cu2qXXPtdtJ9pYWTSITUQrGht2I
oOFE8HjZ9Gclvuwbi9s1PJyNExxskWQiP0WRDhowBuo0m/9y+bEV/AVZVDkrd9t8
lD8+dzYHc3ZrA3L3O7FM74yq+0LdYwdeDEyBRAK+BwW5fYcSeIUKxlpGGCtwYTnM
0T0KNtcyLvf7mLDeC5kkPXuaf0PR2Tot/qLiHxhXoQcQF6NXIEU9vK4AWdS1LK9P
hUdLGGCwf/+Rk42wMX+2n8Wtk/RhuEp521PK7jQO/F1ejZ9Fk4ny29yCxYb92n+2
nYcX00ISRtxnon003AKuURuJcdQzPb7TYHfcayLoexddzFju3OVUg0Qo78LSU0r1
t8blliWtrji94msmfszeny3+RN29jHcQkc//1TJ42OWlcr1cVoyPcqiEOL89Hr+H
kRYQkMQS5c9nb9thhQ3wTX2qRPpE0v2/9xJX3HGT/UQbjP10DhTolE1C1Sf7+byY
9GVcPlRo9O+mdKDaVXYpq38HmnF0Hyz2w/lcBqoCmSgsKB3Kdz3AWFKLTWghtoe2
rZdlKirlaEnjzu3JeWgRAIJhh8vjwU503ndbRhhHt5S/Gtq6/twnaNagAqzJmdix
FaI99JQU9PK7sQJCN/c88119neDayO0QmhWLbTiZbgdQVFHfyjFmcexwqicYaA1r
J6l6RWlCXGfMbqgSMY9zJXuvWAljNuJRgUEUi3BvIxelnpLhn05Qe8iloWLcJthd
rzX3cAMYjIONdiIyTUMok8VuWfPyjxQKDj6lEqAsxwPax3G0TCkeEVEQ3dXt3YTC
Z0YtMtWj9Z/+6LcCEwjOr9X6SWIB0gzYtfyIzocuM06CIF6wZnU8qqVWEzOLHpSt
kOBZoH8pveBa+e1XNbSc/AvdksgQLji8uxVnX55zLnZ1PNUvZaXqkoyfHTa8V5XM
XbHtGv7TbhZOEBrPEYFWG0XhoTkI5mQgTSKhKuyaNrOLfgjqbkHaxtlmOY0Uoyda
J//0WeKkO7irsV2i35aCrvtOqyTUiV9lKhttu5D9bMLRFjMwVv4S1RBVOFToU8Z+
09TGwnSTSWrBbrRuUtI8X0Wm/VU2W3+IWfZsHy4+CLaYaVYBv4iujYKxMCzklLwi
41Y2L9VQSHLy5uk6LSmQtNnVC8i/DF2avT3t/J1FohXoHN2/jvLj1H8KsQPEsT+z
RmLlsEmMvgH/e5z/z7GqaiQ9nEu8ef/9Ybj3y9HKoQ7LUIfrfWfuznCGHVC/yQQP
DMfrL6/j3/aGqCCeclKF4wlDKmGy/45TG7e5F7hCsP6EFJmLh48sdNvv+orS37Rd
VYOyUz3fKQJ7zTDczRhlkXFY8XYzO0jtCFU1jb6uaON3XivX+QVoaTsyup2E4QHI
j+lWbOgkpr6Ul/+fVR3BKOF2Cg1D8XroEl7nOARmdJTXN7baPzZt/3WBBtLSAMK2
551uI+zV9WSXQP3PsUnBRUcThdTkBR7O8PoZ4XOr2C5vkpfJTnrGSE3V4r3PLThD
kMxRgiCCAMbS8K0RkVHcb/90b/hTctaQM2jasl0LJFF08s4ypPBcMyJ9bNXoqc5S
N1UDTR7Tc+IkrO4u+sdIT8OfTUe5Ue0KWraxZzI2xtIhAwsKhwMEAObq7vaZpz3T
CeTwurOPrWQKAUsYe+bsFytr3bWkyC2v9yX4Kl+HZrOwhRJ165uYGQv4YItIhHL3
pfTwUDem4v6trfSB3uFsrawJb4ffcuTbpbKg5uR2KQxSpd+NzUrD7rcoKMbLpoTq
gVxlz3E8pURCsU3v/bDsbgmylMVVU/jqWmcSMx+o+8cGpIkYJHluudBLNv//E+07
tk3xcsTmdteiVgSrOe8NQd+7idtS4a5WGxwve+s5+YhziCS5lit4gWaJmtBszxM7
ZNe99jnbgo85AE9O5MS2k7cVuCESre0lr1+4+WQtNNLlmxM18SFoDbLvGM+Lod4D
v3i4SDB4Zd0vXDINGqAh5ryNWtvB2R2fbnEvSXgutuNWhsfdH/7gOnid0XNeLtqr
Ko+VLYPl6VT1BxWhBUePI1TcS/xROVa7RjlIpEPqH5MrXkIJO4yFrgBpzGBnxDZ6
7BJ4J3bXLwqKj0linWW00baZwQXj4slxiy1RTrL72t3QbZdMw9SqxczXnDbZFvU3
vozB6zfZE4g74f9LGZvh4hnvnJ1pSrundP2h/Q0Zb21DAC51Oz5aGsTmKL17NFhz
Hs0D19Y/PMQ9EX6VRSZAIJ/jhv6s/8SI2SarvtDnM9w2LsOB4OmtK6yI8XA4sgyu
NwX+mOC9bORTiVruEujmuL1YwgrFCrqI4zRfvDjtpjFUJ7WAqJ6pQ1ZLJQbBaLKk
OBUZNaHuYhJd8eYEOPzS9CsgHF9m/c/ore/RJZaqm7f7SgZGFAenChOZgnIaRAkv
hB+Le3EfpLQ0gg9XNg+WEM59ij5fV6GL4fobrIHUwnjUDkHov0lzbGPNygUsFp5T
fyvBWA0Kqtrl15qvRX9N3uixNiPWvG0uWqKlwu3eMH4eozycMgz8ObjrL+cExZL0
uU3pHdsrWPfbsg9HpqEXc4OsHRnrt2p9iflDpAS+PmEess4fFhxnX+GBwLMQHLz1
J+80VnWbU1nx4R0ALKrUa3Y8sUKkaokbMy8YpNlNRLUl9xhGcLnRUvkrmfZhCRTi
4f0bvkP0d/roezjDlR3Vz7eaDi+FgVS29lAlqfkjdprOlLvDF7+Uv8tFZIvRkpoH
XM9wXZNg9vVP7CkzterL8ZL+seKSJq01pY6eOJESVG89n7G+gVMeRKDAyf9sUfB8
BIpKD9Elwrd1YssWJ/cOxoBwJ7qEAxvzud0gX3l91Vfr3is6G8GH+AhH7QfGf6X7
iNTQCdte0Qz/vayiRLKAIdDbU431dAdsq2QZP8wjqevSZ3d4eLxZeq4MazbgoAla
bGqbtmjMoxE5PclWtL19oXr6sfcz658lnmxFtgrIlvWv9YTp1HhrH41EZZX8iJpp
PbxKpkSr2dmmukEUpzKGq9zvEK5c+vhENWjv1b/PjoAuZPhFIyhxxkxuMvmgGOR6
Za282PHwgzqgTO8pCXy6LsOKHIMg7Rz1OV3OLjR7RY8ABbYzl3qLUi4D+mY8tHOB
wAf/wcw65OrNiH+Wt3am13O4dO0mrEYUhiGby+PwnMyfeGFkeDkoDkG68U2Ew2Bd
IGcTh6ckTjgFYOkRzHTSc72iJNpbQKZm6JaA4pA01mbv/MBm1hi1tK6zI5jjL2hp
npJPQjRgHgCrBEftIPBa8ZTHClLjT/fur4PorlqPuujtXlwfOeSPAEbkqqz/FqBO
Aykr+UV7IYXdPx0wwRPFMt1A0wYnpzv8A/W4yhbWinErALHRc2L4l3qviRpitV6t
S3oxVRRoQBnUXvfYGoW1xYglCSVFLgA/IDaV8XkOwaOEAd7uOV2+O15j2aKVjewl
Q2Wym2vID2ZYJX1d8SA/GdhwE8zI9YtF7JBJ1WVAqVIpQZImitLqrCsTh+ViHlxs
G6NdZWaN2bPsnYzNBNqsjZMaCcBrHc0Ocs2xK4KZQgM8V+66mJieOT3g9aCyt+jd
okppuw+l7ssmSvKYa7NCgM0wyQ6OT/7Oj/SJS1Sl9pOLEcohne57ZnMohJ7cYLzR
mXF+tIIhtwbjyMjkCt9KdeoDxAwnPACds2JdjXHHdf+S62e3CPnbaavGCru8h/2d
Q1NP32yeiEFDe0aOoLJG7U1VD7vcBSPheSO7yjtZiexkksubbeb8ofwqe4FHrRzC
IjbvVxAbkPV1yA4SHH6nMAhQ+vtSaSJJH3I4f4e+wdPTNMdK+3jU1184Fwk/VIVD
1CebQoJtxGBdbW4/wp1skgg4OplNnTHyFUOpWf4aQ7w0RcPH48atPWNrip3/9R3u
05R1tOXDlXouZ26RlRb6th5YbqntCtLOHIO+y9R6lHvHRF23gW7nagXwOhLKXBnG
/D5znTJq1+6kZ/DSkv1XYNBf/TGtizfrfZec9tlYJEHfR5QZjgj0eW2aMkTn5iuK
1SsuzZH7X5WuG/uApd37hdw2r7XLoTTpbkYRST1dGD8xUUSR+r4twvFcE9XA0cWY
1sQMLpIwnjUZpmH8NHaU8f3dBYpHib+oZgSRjJzfA7X3AB7BQ3cMwElaDSIAQATQ
TFDneh47IL3zeKtVEcPowGBihKZBLY/M39I2nEOj5WOJMTf3PfFo9vRQk0LRiflH
S+l5S80UT4qrdhsCBSnci/vBABGGmcd3vkbe24kMtxFJW/4lnwJHbc8p5voMGwdA
34S1GH7B0uBUTvvOIwRsfUjVcygDNpl/Etq/09pymCkcRf1INXODzkZSla1U2aal
WPk45LcZFnM47Drh4//+wLQKXs9YhyChoo1TIzWvQMwdB1vA1Z6SrtTkqFOCMfu8
fu6Lew6lQlk0Rb0nOmWHV91qxa5JySD1dM7avpCDHc3XXZa68icXzGxZNjndpXHS
NWLbh7nwxtxf+M1NOrVciKbrE/u2evlqS+SQZj0wPrPAtkm2ZPgniNTvnpawSJ5o
zI3D5igISnhPLdpy1svxBCknarQMRjVczrhBm4tKH3vXgijOveADEcqI2MER+kFK
GSmezLfgKpmmGvB/tncfhe5ZPRnWKX6D2BavnMltGEUcPEzWwqyz5QGuTuEpQrG3
+Sar270VIOr7msL9UANTXmYstfFWIKSxyT43EXY4hPo4yKLDcHKuJWF6Yjl4AQmP
8FU6zk1O9CWxQOT/RPAq2vtndo1nvZvXCie+GRyAWRrXnrHkkitWaysdbwcTAZQ3
5qp7y9PzkdPTCCMve6y1fNtSX+jmqSiwG8AODOgD40GxfhtIvdPpb1FaK+UHYNjx
HVE0+Sl6waLHUdgAFQU/Mazl21De/okCwXH92QU2yQvt/zq/3MLQYG71yuMWux/t
mlOmOvS4a18t4R9+DgDZkG9N6s2HbBBx4J9Keh+XVDtJfh8zROvJpOE59+HJs4Pv
i5vw2zIs+kvPk7Pc4OAaIDZoAdMnwS1mosKYgObwMeXTO+zuawKD+gcxMPGJ4WLO
i0GBNMf0c2xZzWEMNyj42GR5MLbhctlfwjal27OvQtyeRSuwL7cZ12M8KTtuC56G
ulAx1/ollRezP8q31JegUbToiyc2Mwsrt3kO9IHc4a+CjWqdUlKkvUD1TvqnyHF4
VcvjLlJ4LcnXqrfzZkRVq5yLQ0Bp8l0cjEl3cBa2RYp2h1Omj8g4iO0BMppC2SpJ
scSXl91Oefl3PHL3l0s515QI1ENHst4nz4q4sgYoxAhnFgkT6JsqTr3A9KYwMEG/
7Ji227WQBYvCBtr2BFdvcGg8sWwS8Opt/h9cUxGu1B8PymCkqbUQ9UNR+Xo3lCxK
XuE2HAFThjl+thvpEtBbYbWkYc3ZkNIIqmYSiJRlrH7pXC7lvuUhdW4FL5265sPJ
VPYCAZHEig8XAnW1A7vnYx2p/xJlW3RqLoaCVIchgSH39SiVl4FNevyE5AC9oAp5
frU5f/GT5R4JdA6jOhxu97Zs75wC4qRrMYEz3qxKpG4F9+TQYCyPFS2HKL3K5k41
qJ/ViDtfDvS7enidzluHO/OBrjw7UP0NzZtUgVp5P4sjZPaOlfiLtZyniTzkFO3o
48ffrCdu1neD4XO4+dW/5dEzNYRUFCXe2DaUS82jTqI+DO22KGXqJr/ydKIXiWVz
ZWoo+vgv469ukFfrE9BwOVkDdzCTIDjGRPrnEuJ847EpvrQ0qv4q777BcojSjfdW
FKNCeyYqjebjTtTbfNExt0nAebQMczov81Jqm7qRUlWjnMjd8/DxChwoO9sYLLEP
KOFyXH3VN8rNv8BltfMYOTbLmnIf9K1robXecbSiG9AnLWmNXGTW1RUFxt0QHa8T
IorHs3DPUH+1yWjXKxF8UnTsnIfRitD8qKhdFS5CPUEDScZDToFVyMwCEJfvI1FK
ifaTA5EOV6IkNXJWBEdi+gA1T6666jt6SKbSrlWSPw8xCOmsRfyDX6X7fR5p68pC
8F4rVnRKREqCmsvuvCpT9EqZA24cJamSL24rZWxWqvR5H8PmLqr3SiNOcn/VAysN
GRLIH277X77lbStMDQP2eJn7LhOJdKG5ZsbxFNJIn7VtbiRm9Im+WyPRv9D6URxp
uso1dX70/aMT+/SD3S5z2URi3PAu/9fKZ9C60Sg4KYmkam/Ji7DNVOhzldr4Pqqp
1NZtPCeqBkdjdCKnzZG0CAZ6oYmfuP1vOoKAryKe8oQd6zl2exzpaGcB+KkrKyIl
wt03/DGrIEcEniELEfjHtHGtYqlP5yr8RMQv3lusi2kwfMRa00cFzh3hgHkc6DOm
qxdMMthxlYBBVLkJn8aUZMEwu0cUKCTpNcfoyQr2opWZDeJioa5xAQSOfPlixBGE
eikbalxrrLzNmU29LFibJcvXDOzJFaJWljc0qk7hPCgPN1l2gFBcsbVRKAFW5ixi
Krx3V/EWgDmEYSbFHNjadTLnkr1kWT0e6xFpzh/DhqaZ+qHN5vfFcwP2Ir6mXUah
qZMIvxbYONusKcBLtP2UnSHFsvOMjsfMySxfsjr/uhFDQn4IAsvpynYVeWAzg4zg
RFnl4A8Eoo8dKjeEuxMnwOYn4i4oqmEw7UQzlaiIvdeElhCbA3vSeKKP660I0yR7
SD8+QvwW/D07rf06bseSaAan4EozfuG5RUiYNHrChnzQwY3wA94J+UCWqNLexmo3
8QanGlPyDNHoY5nueV9RTGYzktGQV0w2Nvp7bCeR3+d/t79Ma086zltYO6s9R3IQ
sI+uGbz1z3L2ZA6EcVQf7lIRjQ0llHbFJhc6sRBVCnmXbwGK/CCQE6Z4KdCValq0
qXSSx2kLYrZiC74tFyAznGn+AMQb+eaUnwYnB/MpppRINaVNRi/isDJ0e30ea/pX
1ixusxmKGCSG87/IWmpjaTKJpSvQXw1Y1WDcDfwkUJUn9b/DiFxNbAeBqwurTcw9
f0wmq+5VymwIkec1PzpQGhCNr+b8ta4SP19HOs+kcOM42W2BoirfOass19zKWQFl
UtPxdYcejCvr/XVckrhHBAeR7vB6Qxu/P7nG0WzMfkcmakIcv2OukKmnH6XWkjUh
B968M9qlU0EnNmowevsu/pVRLwMGLOh6Q+Jrvs4S/s1QhZGyFzLRBHvwm3c0Ypcf
3unlHHHvAZYqsp5URtC5qIgMODn7wUqcUL8+bs4yHMkz6f7O7Q3MjWso226Y2rJi
8TnxjNXIRdHgM+uMpo6AsRhSTEvwmrPMXzmPfPBuMI6WI3QMzBLrAdzCH2jtV8Wo
zmw3gveXdR6ABWrks1ZmESyHk/2LH+xCIw4p8HDaBPbq8Jczg1/A9fZMGJ5fhPxY
msCXUDG9IGfOj50oKS3XnIM8oe6/NWWN1ISleufNq0lpNdupFIu2E+miMID4Xd/y
ve9Rr6pz+v+jwL5OBHdINYdD606HWIzF5TIPUc8e3SuePYpVLOkPh40tmwIbSMVf
gfMqwHPLlpyONUWb5fUltTxsbt1Z0cbaU5jirjY/ax2E1WewoWny/bky/CSA7Mls
rhTh5JgWWnUONjCj4bvcMzZBOXubo9vgwS2Xe4Hd/cZA4JcUBQoyO+tGe0iFVG05
wZP6OcCeMxax8NPQFPW08AW+Z7+wR9EC7mx66gyUskzUqUM9m9XDSMK/PC/0WVuM
KkDj9waypn1jvt+cxX3tKlR5z4poy2k/d87uMebEuA+FCigpiRbGZWTcnw1RNpUt
2bPRk+n+ENm0NtzW31Xd2wGOuYTx5aEUjzTADSkInNuhdn7po+3lMTdID7ZKb+eJ
Hh20L06oCy11Wq4peSF/bqVmSJR9lgcl/19LicWjyNGqb7Nw3FI3OvmG1ofZxdUz
EXoJxxNkrU/aDvb02tnBK7FZmfs+E61t/Hif5Z/TwZM+cqCWZbrL/bclSoBkV2jE
HSU/CpOKfYFvrzP4oVkL8EwyiSjWPWIQe2PYmAEcUT3KeD0zqbuLM4SK86i8O6Iq
6qtcVTPEwv4HbaiJbwbwYDeWRYd/OAer7lcPKJLP0d283sDLr/SjwO5DQ8VhoOP/
xq/HBQA/3EIdggPn9YibUJFJ2NUkbbT6FbPZ9mSVt09O31t73Lu/kSn28wGNKq/O
VvRs4b9MRBDCn3ib2TFKw0kZMcuxGElJCGlh90qrP4KoMPGo49HQ1uZHvMck3fyz
fi2QCvF5mMfSI1lBnqC2HEDq1w+h9gZSCs7debZLlm5QqXWOo+6PYMqUZwCzevvu
0vuP9yAKacdEvbnRt+PlwY9HCqCarPdEhOe6N8VdSMynV4t3iC4pz9A7E1BUou/O
4mJpfr21pStR51XRuXRY1c3/MePp/Lv4jgu8BhRU72FBxfFT8lT1KDwwOx6lcHZw
2JU/Pi76RYcR5KIPpiFslkRVm5ERUS3jbDUb5hcDKyfcB8mM2vdBex8HczAP1J3a
gwRxp9g7hJHFqcb6fgO4hxugqMngvhIO2ry0YbRPVMSGCY9lzsHp3otGZPWfPtUF
HR/Il/Kdcr1zcq5pASFb6SomlpO6f+rSahuw1krV08QUZ72lDtemxjCyu8Xrk0aw
U4gEE1HysIUPVQmpQKYyW+xhubYc569x0PnvxdjaTaUlb32i9qBlal+rKDjYdIEx
14zFrzk2upQvarEScU9/SvlJCMBkcB8Pa9GQZbBeVzU4QmAY/He1eAwmjdb+iWM6
JtNdita3dNbc8lU3kURutcDy1FjYiIL5EbRjXNLPFw9U8kMCej0QMTPoMIA7bhE+
pWKw1HPq+kIx1DHpWpHcGjbF0Vjv4pal0GFjYkCG32e+OTyYi1Y8JUGhUcLP54UK
6SgkDpPK0te9Iff0TuiMYsj7QWVc+lyFgQkQP8fdA0Xvyo6X9iYSiMCTlnPRyMNL
DJ6Wky79CIfzblLPrCCxN4krTnSqTrRP5TwN4PZJPNsYqSJT10xNnW+Gy/UFtB28
DA/YZ7BmVW61n0/y/aD2OsRAvuqFhRea4ZcUuPNTUazntns8I93X1MWw1bTt+W5g
uFsY1TX6iNiaXkbt/QVLFJQ/tVe9TFhR6Ae2ptKpdcbvBucMe0ChBkYaDbE41alb
iDsSo0CUTiNK+1+G6cbx0Bgj1ftHJgAaomDP+/t+vhZO84ws5eVna70gOqRnFwgU
8kDUTzRHe4cBN3kNkyi9nXdGhtkU3r07pyO6W0jusgPU6TleKUUaIq6HPNOtNzsu
b4T7ksCjiz/9Jqh2973vedkjXv/dGAOYBOq3Ei5TAK9j9jZLJo41b0l/P2BN6fbO
7DLCB8DVQgqVKqKzR/qHVrlBT+6AJ8MMvJKPQ1i9e4DALUdl4Of5PH180fn3gxx6
Pi/N1jWhp17qKul4eWnRpdz7gI2ur7kvlA1Z/cvu+Ppvy76myGW3rKr/0kXbtmBT
5mtLuDMmOdIZJznbIMTTibhXIwreCHub72VXknZY+jiSyxt+pWNIXv7tlWt9qP9P
U348fMqG6aHXvVY2AaOBJ6TUNhjGwp420Ixiym8H/d+CgXcykbcn5hAkcYMUkYH6
8PURP0DJrxR/v4Cs2qb89UuiORnnXSaVAXscD1nAdq5t/LOsL1E8vyce6/ZQccE5
ctvlL06pKEllbVTYcf2TgXr88Xfum3J6MwvkM3gcgP/YDsWRnLhl9rnQbmTdI36w
/dV2sKIXDud5siJkXpAcF2ucslaSN27gEUEiJbbNK0b4SYqWzVhYGGRB4mM0slzN
y9+O917Yyb+38JbVhtY/KtLzm9GM0UXqVvHLAOmr+F8yX+O+No+DnphTxXoPQxdF
XG6vhe2ft0Gn63CTMOsOSrMg9xwXk6qTtvyvYyVOKSvae1zKmWcD/dH1sIavUlSt
jNs3gBxeaF49xinfgQORz7FlYI1mdwDBLwgdG/C7RbTrSRBW4WV8pfWeQPI2Pk7t
c/bu0VyvOB9jhkKeiWSg/wXRuAJPRfigHtC12ZONN98jH1n23TxKL8ODcsSfuv/6
IzeGncffNDeUbFvzh84kMvyhbNZea6IzSmKFOT/+g5RQxamEmmWZiCOpu5yze44A
75ME4lviYo/f8AMENwU2loxu0sOIm9OCuT69Oz6eyOxw+y8EH0ZRsQM+mxxT/FCI
/S3hD97npvfJigBTaPEkgYhA2tQfHLhBwXSk8tLzQmtUEhQRHVxc1QBQd5g6JLU5
SgLML97kZySgTe/6CXyvhAY4ofGUn0uacOJ+KdfMP3mU4LPln2PdmKSJy+FZJzNE
LlygppeJrnJQ9JH7CGyMfcjlBQBcAG9gDnI2IGfLHlq3dYOaHvOVMi0FPv66nz3s
clI7xmCLrJuVtLy6th0KUmS/8HZRcci/R7MzLeDroFqMet2OfI5sEIHXQX/l+5Vd
zovhSHWYz83qPTUiYgIlts1CIKtIrJ2A0eqQ0ULbygCeqUzX//VDwlyMgOgDQkHl
Ktrusbg8nbe5ozA4se3vg58yhlQNPdzfLD4lsPDjVJVHsoQk2AI2acIIU63OEgxV
sGlMRUAkscf5277NfwtpmPUjdQ9hpCYta7zoYKfP8C4I3WBUo6Z1v4Kcib2IOTpE
0O+odKprzhcwjW6hXaU29mfvi+1Z9dRqGsWzQ/He66DUl5RddG8Aoz1tGMEsRoxl
dI0KcmmBR8aHI4riht0h1/ZoqXjU2BPeQ5m5/PxUGxQ6AEURtOTaUpQ0hmGcZFse
iGitKQTf1ObYchQIH3vATcqnU/em0xaPprm23AwdlwwqDTs6fbjOBjnwpm15nRm8
+MUbXslQZbGuU/Bmx1ecwSSW2sfUjH42x8cOLa3etZclxED5HjnFhZ0mLt1hkJIa
8OCNyIGKs2e+7wec8npaM/68OfxHwH+7zEWTpXg8QVTxVB7ocNlI59ybIoQZsKqu
I6rc9UtB1yCKtBfqIatv/Q4ExPUubGXn9/RgNM5eH+bWfNdCK0ZboN1Gz6ucZ5Qf
U55tFi7MyMxPsJZgktxzIjf7n1cUJpfKNHhJALXMdznrfWmDFPDNAh9spGv74rOI
5T1VjLY81i46mIrQu9vYTu8x/qV6Ot44gK/+flBUGnf/czFOY1g6i8QMjMXJc3jb
pRjjEDCJWY/xuhJzbyTsvg/eZucWSv/rtNk8m8zRHOEHlcZAmHzCa/POnGMYjT/+
rsGS9ctEYz0JA2YgPRyRpdf0yev0PI/3onUWDkii4RveIijaXn+eeeVDoqwUyD48
ABKEMT7g7r83vnwvIBm7uWiaSQCWXqpTprGz4m4xkDpKr5X8ZliZopzhlu40b81n
d9GD9IGJrBKBNCVhgokeM7w8rQpE6hLq5OtGQRA/Xu+PuOTJzBLkXKbtw/yNlR4U
+PQ24NpjKpTXxY9mrG4lO7roRFQsUpZatv1Tm8/ybx7Z532xd6ILHhwoJ9aGsZ3F
m+GqbGUvBCM2AS2kqrntfKknFeeduPgTpdBtItbeiaePhvhqteseiykzEsPAAJgz
ETtYAaNDEE3bzOymuZVMHZODvskRF96MeA+o7+jegle1EdsKZ0oUuKQlmYZTlKlT
E7pTclRy5oHOYb8VKgdB7kQeNOUpOi6CcdPPCMov8tUDhudS6vaAgazu5zUyTrRb
1nKd64Dy8rLNhCi6SNgYDTvSFE/Qt0/D0MFv71cdvywR0hldqxlv9UAQOsvBkSE5
qru8YvIeOhoyFLa+JPCw5hHvbVsz8+rJZmcGFXwKxVNrIQdrX9BAurppNb4B70ix
UQCVlXygdL5a9ZbgsDaJKVXFTOdOb4NDH6uQDbR6C5VE/VoUff1vxZ4baSE4lKhM
1vqv4v81LDuyD4e39Ob0P8slv6XYEkqoXw9jkHUwZ6/4LXbR49xuoB2AcX5OlIuI
l760Himd7/seOpLJqFBB+J/yPfB6ayYcmx9i3UB2lmcrMJGZy7yqa4VcHK7bTWV9
qpWntrD1dylI90ui/ODCQj0B3vC97RKnu1Vq3Ai5wpCv4UVsynPbhiRPvULGlxyn
MlbzMQddJUOU91J9jkL7j/S9KdbvzRkEFO9+vwVui/2zyWGYq15yu+fxtd9MBjNb
illVuPue+gq+YlQBqAA5e1yTEvetrSSii2SxnHzpwkoGVf4uvw1dsR0MuCx0mTqi
VuPi9V1fk3ebOCKaPhwKqNsQuLTtXsW9tvR8kLsVrhHYw5Ic2EBCKS98JLNBwNc/
1Y5aELNkzWjiLagV7yCR8dWLc3yHBGxFfYVPVvEaja18SVVW45aql3vMVUTSVK/e
jOTBF+0F5AvHxQNcRFu2zWLbZluCBtVRUDkHOgN1G/MYCzrTxf0j+KgFwDz6RPf6
GnJdfIB8N7uWaT6jh1I8I0UvDVVYnGLpCA+dNkOp8syXeq2hXnaeXgkX6C23LWtl
UHkVXXKkG21CuIuZndqOvt0mdjihGMv8aVwlS+VtahtGwXDbl4TguK6ftcI7t2M8
FTsNWPQAK3WgTAz5HhVGm8sc8rCqYrOxy+A5yG2nIFLPjRY2GojOGirFRCdsFzI4
34SoPNzc25JskThPaVNzm4eRe0AL4xhXSvv/pA6SvIhowKaqOsngx4l/ZIUDnjqk
OyKxxx9ruTDETbmMf8rgBgS9W8mlzDaPiSLHqEHL6OJyGVdb9Cry9zyyrlQ0my6r
VokRodmPe/1hVK13l8LqvcDzJhLEXT8XASrehhIh/uiZMJVgjOI/spGuuuTlPjyL
Di7TFvNWkUNC+94cF/t7/hKzb4LVQsMr2KBAH7uWYmD+bIdvyPXy1t8kQx4xMtok
VJIP+mYxEsMD1WLd3K9Lr59OVSkOesSjuXO8HS0j03dSDQQBiqhMWqDcdYvyZMKA
3H0+EJDOIumbaRYyPppFHJE8HTwNQuKRu9A72Cd05IlcD0bStK8h+lYrQamJBrM6
XrAu7sO4cibY5NKWaasP9L+E9SOk41Y6OaEZ7c6Cq9k2tE3jNkfd8+qxmAQovDZk
0dtiSp0bH4B91IT0FCUJz4UN8mAp1wRBgsBe9fl+cCLGt0pDsMm0OQw/0NVvkd4u
phzjIlw09B2Jjc+mXqXsI5dLhzvyqQ6XfKxMF8QtIHJM/34VyLRqRZlsEMDM9XrW
qx0Sk8VicpPSWN5g2uBVmSrtV0ppRlyRbmpR1s/2wUa07ersKHiwJCiXBxGRybls
J5DOGSpXGIbL/2D6zRlQC5d4r8k+QpTO4ypU9DwkgtjLoxjTSc7rYkf5xVJ0/mjK
xoaz28rCl56fSyfWjLqDCwq2HRAmM2vOLzXFmNduOusy+qV2dr8uAxb5cix3V8OX
9jB7JGk6pEAEaNfMNJxSExQyPET8xfBklD4hin5vReLLt7cHEa/8hKHwz8+dnaHL
QBnD1GVvs+FKgMRw+xqKSHiZ1yFeBqzQyQOstvm5yI86EtjBKt7Lvz+WTnTJgYtV
P7jCaNAUEM4lbhrvSx3Q8G8/Pw69u7KXLoqlLRYaDvh6QW18WSoE2R5eiLcYhUBA
Z6ApD6AqTKt6e0s5GdoSewPEwNOY8NXMtaIEEGkDye/A9s/sH0nOL/YedjrN3tHJ
slu5boa8kNSBLV5CQ/os552qOK6xDaES6a+xaHwI1b7YSnez7IdeV3YcJ7x7BLJX
b+QO1M60ek7s8I2wPLyOf+fYLf1mx7DqA8aNAf/5sruBVDAoXDljXXkoTURThMRe
lhu6h+UJTJOck0Ky3Gc3iG/AvYSSr7DcMOiVK3wkyRE1W/D4LkaUh3pbtZgUQIB2
A153+bDGgh5rLZjdiVxc7FuJGYQTzW2c6DMACS4D3A0aTNerGbGLiaeqd4JgZ1fr
iuw1RRRiFgP3XGmHYW8EYrdlAdFJ2fHRlbzWIZul5Duo/I/jdIBx1ANkMj7YbTtR
W958RSzZ3l7Xm4qrJxnuX4Y2YX/8BxUzC5WlRMVE8I84h12TyFf3tWzi97ntFVzY
MwIsjHsxt5UFTQ5hQvRltLy4nPPIZCcTrMUElu2ZI5qGUA1HMqSha9+/4nCJyzjZ
gkoY+S4y+VJvxQHVprvlra84+5pJui9nXqfjP4ALICnXlCLR/n5zFv9Q6WHpdHV6
Hh3rYqi37LDwvbEMZwoOPm/Q6wZJZ8Ca5a8zt4Lu64DjsW3jRnuRS+P7jJFym4im
qf5jjRuIng8Xi4T/xGdZ88aIXq4kA463PdjtPo5oclGbjXAEHEmvaM5l/hD9l9Ty
wZskmBtk7CSE88dUqyKiPCnxdGZwjUzXeit8DXjanH9MkiwrchKFQ6kl/JDx+zEy
e9COVjyfwXseewpfgx2sFnjcu+0ERWXXnnYI6+7lgwHgbiTukFFso7+Zvd8Zr4+j
DintGqfUfnBNuIqnPu/Oa2rFV2j8QML3hRqZgYdSiMApOdX0mtoWXFHFoUjOe87X
Xp1rKl82uRFJuGuS6TWAM3IgJAjLd3i/h8d0/yPeyKzxvo9nW/Djx2bM8NhfVw7c
3TixWaDRrgy3vK4bL+ous7JH5jySQ2LQDTUsnBJUzcUCCXr3L9CU16XFjszqtSbM
H77osJiriDTya3qKlRKXpjcsjSz+Guk6TbjfMTQ/Pt8EiNvb6h43kDBOu0OR2tXy
+6i5LW+M2pWqc5Mk6iMiWBubjS0wv0tYY2Tp+cTvfmGf4EyvP7knJas38Rv+9dR8
hAPm1MZHt2fmym1xoM1TlBySQK/od3o5r8DQ5GP96BEr4B1wfDrUSoO6nH5Ck+KS
1U/VmqM7+eFlB0hTFL4iOQXx8K99QnwhXF7Dl6xsBmE1TazMwx9sv0yg8aVVaNXx
qtkq9zAydqR+PK3BIqu7pszXCdM6SiFPH/3CNj7vScXcbPdQ8r+wkmwDkywyOFBV
Fp7KZzKHe2p5iP3hdoadtQGFZBOK1azjxFOojwhWvou8JvZu7NuFQPFBz0Bu3rTf
qAUebOtrQxyiC3BYjD+HAbyXiBA454Q2jMUuJZad9F+tsPe+kd3JNqiyKdMtH+Gj
QJdRfzWRRr2NryQ+gc+hL0JYNKYhMKyMGw54p7d4SfB6FJa+GHBuC4MPPinlMoAD
HfegvC1MXAfrtWheIMez1AG5ibOeyrFR6ltea3SUYS8GySLVQipYOh60yRY8reAU
gNe0IcQ9pBxNZPKmcPs4YnCPhPv116i7dfZnFa0EWcZXinz1UiWUV/3DF+G73V1M
ofsaiClgS19rNFzkstttKg+/q//9/V3OdCRZtycwFuHoQMBzKnMoBQm2uBMxQiYQ
epNHh5NIpBPC0ENFFQ/xFBnp9iwATq5AwBGBtlidjMhdRhPl5pmwhVa/N40XVpM1
7RHn8vzgMp3cLgwQ3KbRelx0eAE/sBX/+6dGTZIxOJO+ab4j/krkhskfG9K5w2F3
rEkrZPaHV8NZa1gDNx1Vv/n2fGXEH3WTM4KLYWmWoJxJ31i2jKzqHMoKESzgq7lN
Tmr1u5De0Qdl787CNYdGJN7Ft0fMgt48UdecQpzHaxufOSrYAcSxzDDOxql0KpNf
Ui4Laht59lK0FQAhyhBLKNSDstS8cej4RlXT0znNVnGXJoFf8d3+Ovjrkebb+Qx+
HyRstHf845wvYnnQt0fvPpnuDDgZLzfp/Ad8ZNYbY2S66xhGeU7Dj/xtTyW03KRz
ob81mF46djnLg6NfDV6tgaGI1gTAJCIvK8VJ7Qxf8yuK/mpeJhb4oIF/JqczEBRD
ele9Ni5cAQ+nD0VPs5a01NGtUIMX/Spl/Cq1SrEOH/yrgYREUAmjXtev6b6xhsZn
PTA277d3misdCtNTs4xQ6kYALskINUXM891i+iccQsLqmgf8Vx4vWSKrEgNaRD5E
prAFHq3e9bpkwSq6PAf6rS+dLcqfhhTHyUo56uq7Hll3Xl+lcbS+E9hyRT4ewZXX
NQ09RUW2PJBeBB3ZlKgpSWE+IitcV1Q0y1OEbvKP+OzNdC13gTPiWLgPSfhvD2nd
gGnZoKmtnP8Bg0ypvHOXMnPwbcl55sAFoNn4dnqfPqfvTXpYYRZmtOWnuXiACsKM
bJEDres7XS52OCsOM3xAiLJlILaXX1i28rDoFafeJKHLXNFsJwHY+EInLSFVtsT6
Wb2a2za26JMO0TND2r/8yDhJJOFzpzN6i6oB9/CsJbmX24anMBqfGo58ggI9rQuI
yNWj+p+2JFpw6RefQRkymLJzMbRqIcHJlnSPJG+WV+sLDNHH3TbICXWFv74FJwsR
JG/4uzXxmp/E/9guZ9zA+z7ucPibWhFpPKco7nxbigsGOH5548nFpwipXzqMjDVr
wdFXrPXSZmMBfOXuj2849wvAOC1V8R3frGwQ1AL2SgHfNTslMEtY0ctc1pLj95+k
mZByM15LLPkelq+FQYBHZPF0n6rtVbAn66ROR+z85moYyIb4PNroVVvp+Srh2uIN
7JnbQJcSp0YP+cqNB6S6ZnAkfXLtb7v33J1htCY8AQplmzASbJ+rTknBHkhlEBa+
3gjoHBAzsV3zkgpQoYyMk2EgWhO031KJEJNwXcmiJJIV+BOY/MSmD7HMXVJIhjK7
GEWHp/zxjxoTVdK8cgYKPH+KYwIgdwKxt9q1z9yoCEWJ4aUx0YgqXtJpmc24Nn4U
j9ioQkHhJ9Al+2CxItRkYGNvyWJjMc59BPNr9U0d/dd7gABcIa0kt545zEFrTuYC
wjG6nCTXS6PurCNq5zt92eeMZ+aIBpBffZTfEfPWj8MAa3Tv+JpFwNRoMLl8IZIS
2wVcxsQXe1uJ93G8p27sEAlq9s3f3UnOU+bZPMs+5Nix372/PBOYivWARFawlUlD
FD9cNe1IjDKmy2VBdYGiIlhHh1G8wyOI5kpG7fFWSkESmkVEhDC5XjHiKrW/Fakk
RKGAjpOBIXNmN/VovAk1kYfBYBkahKJkbOvn7fh+M6iWv9PeEqQSuxpsxhjmEhBS
dkBan+MYaYLp+Fl4drkg+UjobetUduJOrZcnB4Mzr+nC7hTSXZoQHddWZRJJFCXI
PXhw931BJUi/LhvTNb9FBJHZMf5sSpSK+KGkBXaJFzYqYh74EKXwzh1+JlNQyWBK
nVsLnlnlG5HdPicoWea8TF04bJW3mNTG0ApEO3Xe/LFKYtA7go+SCMZEak/4yRxr
ucZWaUovtbkXFDKK5BHI/UFnOcnA3dx8DocKWdtOdxsxo5nN5kMsWabqURcHM90Y
bk07hvlNbJMKdC+M/tgeF5tKrIgFdnVz6mzhtxei62hE4AyGxytRB2TPwXEwdixD
0tCDe5/hnmWzIBugyEE/5H7thO05M36E3eec07sQbkZdYptaiSazZlaNYihPHcGN
fYMzr5LG55ipOInrlfYX/j4IaVWlB3/3YXFs+50zfrhyzBp+TI+dXKs8sAcIUSsf
FVUm7WMIWik0tmKXOuouvRaHnVsNhEpYTi1IVcXwoNs1MuUR4+ulnYvUk6+oDXZy
ziWvxiYBIER9EQuCldSnT2AaGdd36YoOvtPlVsglWIWQWGCM8d8AoCKUhJI3PKPo
70mL84YewIWhaTaWwU4VGshRPEIdYObLsdMWWm+K0Y8p9Mc1dlQl7DvW/LmvHL6x
tWtziHo73tDt+vIzp929XmoYvxaCvzyy1aDUaRLW1TW47wxUU8G4nIq/yfU2mboX
Hwl2JpcZ8QIZcy/opnYlHuhHpaphA8dSj0e76beksZPkqBOOFRsLGZix7aFJMrHJ
hsW2l+J5/bseIyTM1ZwHAuAmCoDgtEZsAkBmPZKM7hHsITwn63J/vgS6ifoo/eF0
jvSoD6XIoEagERr1GcuCwcvEtKv3SAAeFkOvUtWxbKmz1Zr6WgEVCkKszH6qPL0v
URM3dAQQ5TSD9gZ4TD+MNcbcL9bZOYGQw9fiwRijbgm4NKphMeYzCDAskDev/1VS
efjP8C0UL/Cu11VN8yiseEHnSl1J/zpFcWQKzdhrIIp9619fGUVy+OpvYpClA3Ni
sspOmP6ClUUoCQXUowY1RjRM2hTC85X4+eSCEr0iWjv8ez00mPj60mhJVXyhe1Zq
c2QtJUccNTCMDHdjEzrh1cWN022zY1MVi/2bjW8nqfsP76ddPJaWVtadjEnN8uNT
LxxqRVVxjiG0fQIb86uFUoZvBH9stzNoEewooXTglntXvgymanj47ya408eaDlY2
O1KzVifxo6EZUjC1gS1eXgzs4UcNNYfOQQNOsoaCMQ9GbJoa711GxnPvecYG4iuY
+CXH6KudcZFo8JPGNiE7YJnCk67lPnH55dD1U6F/nzz4BE3lFG0Jpw0AhqjpFP5p
EoQMjyaOPbq2QQcrHxhC1kQGsVp+e7PQHqD/vKPN79IHFXzwM2XgGf8gWla4at5r
zOXDk+FMYzUne5mpAzwgmMr7n/Uinb40X6SaGBRqbQ/e3JAnooCNLe15Og8oGf+k
eyiwI7X0XgyeGhgNc8hRkBAKQOcN48pFwuXC16R/E6iRHt0ezLNLTI1pBbHkCo0y
ptBztWeZl7xfoHlcC9hTKr9e7sRpXbHcTC7Kh78NP+r84XT/QWc176yUphnUKY0g
Ox+KmQZzLOFM0zWvraQN7s2pXziunWahe6CL+g0ny84ul7WzZmlku1BJdsN9GOhc
JIZ5Xc3QAAjnAIN78BX72VHX6dFsgl3RLg4YpOr99gLn5odY1tPlDskNoVP8vAtG
jlAxrEeAB/ouEFTPy7BVYSI1FBmchkrVgynVQn5gWG//FX4I/OjS5YqzPB2DFIBC
yNjDUA54bhNpN3jkHf/G4zDRwTFN5OHeCmoV6KissIBppW6dksI63F3e4uz4KGHM
i74M4j6QBP5wE3PrCrfSuchf6/4jHSsJdqwzNyHJBbVG5t8rtIz4fNrwaRZmCn4c
692tf13zrgdXE8xA9xwUfSmpJUkemBK+GwoI76zhVEnXQ0zTJmEma+mDweklyGxd
Xt4oYOtBr1ZEm1hQWRx8iL+Jl1Rakps0vqIvbKZVE4Kd2OAoQmHxHlTyCfZ3W909
IGOkkzz+2Ns9cPAJyGho+YzMCvQNJX3/IS8cBcKZZSF9/PH5+q/URc0O5o+/LHxk
HbpFRbF3Qv8K7lR+B5l17M72WyrQ/EJ1H9PfH0NbgAa4Sm7b8rbztnsSF/7e6TbO
eeb1MnUXZ4eHYXCZJUgqLyQL4abFA9aAAykzVP05OvtvvrX4jr821OlIQ6QKQJDN
aWiU1IrW/lE+Iq6orjNVm8kdJOl+2ix4BHEVpv4qe1/C93pQAb5qrsPu/fy4xi4e
4P3avrRgMe7SDXPmXACwqQt8t/bVwkmjGBjIt89DtLAjlWJwLG/4VqhZJ6jbC6Ji
jJU+s7vtE+8p51qdXqtqdtiClP/NjnWU9BdEMWqeLBWgM/LriNU3tcdGMDUwO/3R
SdyhlT55z87S82cEPItUQVYSDsVPKx3f4KenYHNyeHRz9D3KHdN/ZKYviQASNwpO
nwoF1DxOL6Enxgrn2T7nT9vdpj85t/c1rzc64kfINAVA9qMSH/derbcbdiLaDaZx
Y/BGqmXJzsInZkfUb8k9sxfnWRq+MD8yzgJPAbvD1JjuAHlA4jN7FrKQ4M9yUWiW
BBdvswjHyYlen7fFH+zRuKMzW3Aaahz3wFPKNSR3xRVbPE739IJluNuxijlaAdAo
0VhgyGVX6ARm6j1VUvZzs/zTsS19a02qRT1VA4QBAIcyQFkJI8//9G/pfb0OD8En
9a6tYp5Th7UlOm0/6V9HCxTlEVxC3NrdttQPaEShTBf9gcv8M8b+8yHLtDCQI/Xl
k8Y53Goe4CC4CNVFERJ+bA9VtdC7JjnyMNYtatRR+X+nv4VNEgtCo/die1iimX2N
oUjuZEohlKVy/+53b6hds5Hxp/Q/NMr7UaSspHMh07jY1zgUuLT4aZrwmzO9/rsX
r1z2Mo9ScRwCe4xcfw2QH7S4xncnMSFV2Wsa7r/zTM/w1UFVfMXqxmt7460HZweP
weWUobq2p/YUcIN+2ZicZ9q1pkUyp3LjIsZP3JHWPB8PCftHHBjH85WQFg0t6ZoE
j5/dtmt2DNOuQTqjH7ofXtbO3uqu/sYZZ4FDl+d6FkPp9PhUpBUegUAh9L9dVCmp
N/4IyBQilyKx9GsREe/VZK1zaiAJ3c3EK23jpI3O2rrIhiw+0PCQ3TW83XGnkKcT
ER3f4xPX5yoroJKBF3yx7Of+ynILuJaHklIXTLkSQ/loL7LQo7NtS/az68lvbZAK
rTylKRPEdpEFGg7tW+LzksSWGVcM4VZJDpKrKh3vRHKA2NhG80EAkyQKzfoy0oZB
SJ+vSePtLGNWJPkVB4h8XLIQ6PMPo2eO62chnx6cAw1V2XhPbU0etrsDIS0zFtVK
s5kKa8uhyQXXs2T4z/kizRxSx1uxCNuyHE74ipHHLdhosjHytEKH7z/PGaIR2djn
YHE8oGx2SsQCeuApK9/1bN73qOuBORJtGc+pyj1LGdxw8UXu4tkmHvG9TRpK2QwB
hfsu5DYvz6a4qa1u04Nik4AKMa+JgxIiI+tgz0AcPpeYrjYTH9wlaBmzHQ4+AD/m
ONH/1bJI/kZ9JJQvjucdBH+DuxznLt+sOhE8MLo673m2zUMUIUQfA3S2usvnBqar
atRt/igSRfvwOB3dpvNN4oSgvUCxh+mTy1A6UQUpz0El+5XR0b0aCH6tONXS5jiU
dpZtAU0+/M1Fwr4OVQclykfHf9iiZsm1vhvsxosyEy7d67+NElsnkslw6kFe65M+
4U6SutjV4cq+klx5r6xQwUeg8mojVAPp7MI6BA4Ol8SCA6Eg8ToUKPBp+3G1Ufw4
iXEUJD63NSw+NcJKyoOzzH52ifVrsmzFhvxOdigtXN8rZsJQuueJOP526GEE0Nj0
AQ8Wf730Uqnk2O92cJdIWBNKMBLUi0Ig7Cl7CuY+qxnb+CnLDzlrplGGsAxiPmmQ
QUfsOZbvywgiTOy+84l+qTDqug9Z1tQVjQwS8PVuCZjsyX5l/7C/A6rb6nrTkv94
unvzNlsB8rqV68n0HT7QaxBJ5beT805vIVa+ORRJB2KNyXC1wQlelxSxR6gEwkyw
gTaC9xKerv5I2AoNtL58z7pMiTD9rr0sBUjh9XFgtjlqJJ/zPayyzK84lEX4Zj5M
d1De14grzn6RBFSNkrHYkFXyYVRTJyoF4GBSj5ijk6MpdBjPGOrB5zel+JpChpih
IfzN7+lrM+IOZKuJPMjQiajKXsPzpwJcMWxuXkQLWjFiySOUW2FpArX7BaonIXN9
cMqjYG+S73qamOHXJTKQoofp+gZqeyrXyY6O4WfN2TlyXk/7Sb57JDTAz5ow8uBW
Lx2GOPmHTpL6YzS38IVDNaF3WSrgaGGeR4MxfwSXlneokvkkbtvOyq4sPPRglxpC
sutBCdCzZZDEPw1PozdtvC0X0tBEEyEhrBuZnseysXb4cNqz6/ccHIrd6hJoUrPV
zA28tKx0ZmaLXOKN4v42Yl/101XE4fbYYOerPovFR5GzQRaOOQx0FFaFoVdjoOiC
aXBmotNBWkGrRg7ZHNrzJ/zqv/8MsUAOd2wBXIcXF3332DtElV8pml2M/qbyz4Il
bQyET0XnblhEd8hMhfQjRHBaVnixuicUg1y3ycj8THF7T9Nfn/LI4BtCm/gZjGuk
JywkZ/AeKtknZXU7oX0rBjEwbyr53b0YedwUZyqkk7kZQNbd9vNsONf0Ddxs9BvZ
fXyRaQCGOmX+iHE4GPef2NwFDIFwZXYCSjpk95F8IB2Cezt4ayBCFOSWF067jWDn
xiYbiU2CmvnSiL67G4npvm7Nbl9STOsBVDH6ZyW2qCg6wByh6on2yI9sZIH2eaMm
oyb0XkPTodlhAXCqcCGuaLp62CzyWSVc4GfewHD3YSMjey3WRvwByHOvHtPvW7sa
pjmJGo4lfoqIsa8dOAL41TO0AEye/IzJjBCBvgwfpIPN2ei8I4rwE7CkmJDHsmJo
YEhoGCbaC2Zd8jQ0m1uQkKSbDpEh6wDa3+6cfpyQ9oAXHPus+27y0skF/xXxevzZ
RayPjsRUyW/+s3+tdgx7puvLx7+aEtlKrvRDiCb+uvBj1icwFbVWwYGOTFu3pquL
+dYl7S370e1p9mu0uWk2cWvD+Fn+FNrRMWS2mfHXGNqATTnCapgD/5McWNZmOkKW
0uGOjWONh+p7rjrZxuUfT5zdpAx8RVDncjPNWA7df4ZdO7jQvo7X6Z0pF4qD9Coj
6TOiGb6tbtZpyUquZARGQm+oX4jkxVPt+ZYf2gINXs96YrcMbF+U3Mg6VgA5gP42
2RYf3JUYs3TFd0wGwJ0nZ3JncY2zOJZhp20ZIlRCo/6MdB3Orve2PRJCHqowbCyq
JAl0P+5E5ZbmIDmib8jujzZE9blm2i50lmoVNtF8IgQsbYpk4c8P0/OwYkDaoNAC
jIkjZ8RDRJaqSXA93jihxLh3jzpxxxuPvGJzp1MSmN7AZVFx2agNi+Ti1tgo5ARW
k4cAR4WwScV7wqjdz9TBEkbMh+71BEdQDhxfyWmvqYORRNUkJPf2BOP50DtqiLkt
B6Tkuo8OSqRadfvbtimqtWSFdzHs7mgYXVbqgzt3mFMCm6D7HcKCbWMW2ChjKWZR
Xeto71IZK3v4qbTthbkHv0Gcwe6hJ0mK0oldq4saZ75Yn86xOe968nmco0MaSzXg
8eNENnA2plD6QpmgmdAEIxTdm5Q/3TzNt0jGkGuWTEdJGhtyuppJHj83mwefDRnn
7j3XsVXdwARfXqCNRFJGLGSEAU9iN81HDGLmr4jSKjoic1b2P/6gm5PtyFWxkZ0J
Ss5UcbdY607gzMuXk8tauvyy+U6UX75tG86A7uEBNjmmKd/A92Fopl5/2uJ/4Xvs
keSlj5NMAlvuIPxpEDOQGsf+mOZwFc3TktkSov6bL6AwnCTshTNXCwx+I6WZjpKd
e3hTfUhQwFMZ7Ey7buFZ03bbnIY6DiZ3bhgAbuiTLxuXokpf4GWlSTEyhuAeP/Wp
RncQf3mUDZRKfA8oEUdwfu1pZFfnr+DWEPGXjO1WTf4xoIODjo8ldU1q2Lici+an
CJ/FueCX3RYC4o/hOeVhwmfQIugbZ/OaQj5q1D2kefm5OdBO5L5W1Lk5wwIwGjPW
jgvhZEVS4UlScWCaEZzJBW9cKF4SNkGdJzpWTFrWQwuwYtu1m+8p3E+hD0kn0hpt
fm4TuiCMvbzZaI34vIo8ytn2WOemUYeskxtIV1rLPKdqxqkXXuOjpN4SDEf/UzGy
AdDxokvfF167KJekUyG3zumetc+vBq6uilNBUW0/SQA1nC6CxzW6V4bbT11gxbTB
jWVNu9cSJGQsbGmKjZHGdQELP5jonx4sYPqXK2uowvtycTQl6EU4alJoosARyFqB
3vxBHzzfS6abQfUDymMsy4b2MgRCYFkIrKbFmrohEmio/wKhEqPaA7Y/q853RMOi
KagvxA+Qfm9R00E18pwPaAfzh8RNwh+AIwWUNT1Q8u5CfprtFNHob/wzPyJDHyyI
ohzs8J/robiSAy7Bcp6Co6X9yITkk6pOm7Ob5pACs7ixfu7Raw6FMQNCplnFP3TD
KAQNj2W9FyB04bgGcDWmCWNqC+usQylZheG3OY/4StZA4A06aysChZmzcEyyTibe
cAX0LFyKIGZdHCEN3U2keEaBT7nvXAUqKs2bjTfQgv1zsqV8yRM6WLYqqvOu0SUL
N38owT5nu8WkHfm2ZqarXwv1Jcb+HjY7T3VvmEmWuDk8wAdtwK38soWkXTT8Sgnm
tqPloeLU+UcHovE6fByR5VHDhGEk1oAslK3CUj7ixwmVb1Db9XQXBZ4a+on8Y5eS
QSXo9YASwb7O8To6mwGJhkLjARnu1PVlnzidRnrP18eqEFYvfnBiYn3b+qotFzhm
ISMyT80cIFNUrxi9EV/uHh/RqnPgP62wxyfB4TdB8hPcNIjXuBbBcu8h2tgwlKAL
Beo3BkkrHillHpw25g4oj2xyGzN4rgg4DUt1fEVqJkXhn089RwBzzqdcjKxJT9WQ
S/C3YTQ58uq7eCzV4ZtUNOHjOypg1byd8EHO4184I6B0pl4Idu1tRHk2csiuFPdH
2VSGOBawN+pwo0xNOlZG2US372mQH0T9el0k9lnIJKWFneTNyK4o7BQ+b9jbivfJ
RnqpLPrM431Y/hQ/s/pzfXH1xJNpPhKzBfK01boISZ0nmmqeBVdAmCsU+pwI9bBu
GrUiNbVZADU8xLGYFyqqdHELTOTDRn9u09GFDfBXIWT4SbBJt7pevWEfqEttyO0p
pV437flLVnT7BOTilebTcyPjm0v+UerYsRPUXRCT5riPq58WBI+a4h2lAGgktb/1
jVH3t3QpGgErI1fuwq6bdqmoSMEvGD9+fxX2QSrEFD4CHr7yg7X3opVNlPS17QZp
77jDyoyG2tFHNhamDm4XuDhX3hJISF2815s7eSLiOdfDWythF2T7tPYQiq5Ypitf
kQnBe2+m7NAeUk8tfWLyEaLE5cNf7uj1Dr9fla3BVLFsp7qbD3ZesA6DnAStP7vm
9U1W/+S38WBLsH47/QnHInEHBmiNgQi4P9h4GgKzpAcaceGdhlsmPC4F01G1CioV
7dCrjEdA1doxwH39qhQxcVcyRuWn9MN8A2uapKFSv9Q/IB4bbogWN5Z0/EwGUQg/
HbKe/m0B//LcKCikHNvt5tgNAqstXjt7fNsZGm3xwPHMAj8qu5Pm3uELV/BM/24U
IWGr9/VKlUZF7xVRYSnoXs5orRZeudn56VzYvH3EbK7lX0xdSCUi1i+chJR7RVp6
e9pqbpXf08Ck3Bm6CPQ4qe8Y0Sth2sKz9+MdSV23V48YuqwiGwA2zObhH6rEP8M4
Pa0wOYtM7kLCmSxCQgX1M6kOv1ZzBVtD9rpSFAiDSWkutMWl7P0/S+nLJxEL/Lf5
AqJMj1nW80qvNRiTAe+NKTR+EtepIPUMtsP+u/crVkSJWpUdBp1qULDpg0psSo/2
v9NpyEIra8llnfDyPnmca+I2GoTwm4U1sIAOw8a9hLNtsgwucdD4oOQCnz7OjV5G
o5C2TgmeHe5NGD6aSiHeErhphhzIymTdjJU/FbhcL9z7pRvY5tYcXk4DBY1lIAdT
AUHBwKDOBDHxZV+3grIhHSkV5j6C77HUjMU8FL6OxuuJmWranTo6dqLP9Z+qy+7e
ZzNFghWuGz8xAllkut/fhqL+vY/7wi2X+MPn/sJLR56MOEblrSuE+pVUvtPodF3F
ExsFEHHt8XXAecQVq2VOui+7fh3fxVCzyzkhqIwRDqf6EBPrrpQbE+SXZu1z1jY4
PZWWb28OZnoSOEt7BTUB6uhLs1ReO0QQhtwEeyFYiIpZ9MltCtkkilkEoSEdXMjG
AemH7/TJCauhhGiXBmvO8QPD0iy8f7zCXEqzLzLLSBjA1rLkVzsoAa8MlqXejtWu
ywP28bJsNE2gpM+6CMZw+kGe/fHTd8g+tGahxydugg96tRP2MwdpOB7lbyYVreSA
n2G4sYbibQ83fBDTWHZsA9XL9Xzx4ROVuB0qEXHj+MaIlKIIa86iM9Iw5wiNdvM5
8JjZlFFwKT84Tf2nhH3ctp6Nj6VpqVVopBXkSXDT7RoFjkaAmQSk6+EIe9jk5iJm
nGQpZqcewF1XIm+nwvWHncMPevFEKZ3E7Qmgh9ahfVu2Afy2wz3sZ9MdlvPuO1XT
vjmf7jz91s+jUg1/m3BzAm/PIB1184T9R3BU8UJOhp2C3jxW1h6wz6C4bH94ZntV
nUrXUa/4fYGmHmv/75DKyas+icJ14gpWZhaY76n4zBQ0PPTGvCoCo23tDUlF/DEE
+l8P3TdxJJovBPYjqnLdJMrc2L2YRzEcRW6NEkIO4G68/XP0lT9IJ5tj+cYqcmTM
7wx3L0beiHkqxXHmw3V3mVqS8abdzPPL75LubQh85GrVXMQ5sIuH7/WyVaRY3r6b
elyFCG9t1wFobqrjcesw822EyjgHJtrvI8uSpzQ1z1MO6jZvpGdBCnB4xPqhcvSx
EZCtHLh628ie7gysuLwWvoPR3RRH03Xe4Du8o5hrxx6ZOUY+hwHmSMi34iH5tlBl
GNm41dcqjZ+KOQLZcMEkkJXpy4XqmoxbCBZmxcBEVqv2hXbOKcnp9RmXnOotCtPz
bxwQNjbEaBDP0niQaMIfd76HD41NvWx17wYSftt4tDBwBojR1brrEE1cXmW4HVQQ
NUEr7ZE0ReIk5csn2eVufO34GELtDHXIHNlEL9FRmkFJDXX4ZuAkn5FpgEnhabqJ
I5YdkGtQfdKICzvu/Vz95j6eZTLU/PX84TQqj3wu5wi2LGEFl4YSSlC+DmHOmIyk
VxUnw/wf1651s0NtMYTnS/XC5Wd7qIVKZz/JQk4IZFy5JBFGyKFVHJLIhHnYaiqM
tjPonLi+ZvzA8IYCKVs3jYB0fh6APpoKJ6dJpv6IFCJfk9eEqNj0nj+hgvZaekq9
YmH2wjVfj82VdrO7w0iwHXgZVm/9Z/tnjdRaqhkSDCKbB4hNrFznusrfFkasySVC
m/+p26dx1mm0PdBUR1WxNE7d2/9BMCO4ow7M+wj1lYf9Du/VqJ171Ru3KLG36ka9
0B7hNIuAckeHXoDGAuz6nT2oJkgmA/e9N8NKM9p/YS/VZ7P+CmAUEKJcZ+skN1Aw
RbY+oIm6Swu+O9NKDDhRPfHK2ZMNuRCEual9MNrBYQB7HQ5PT8kp/eYiy2Hi9dAR
Zwz6eMrt0b2vL8lCvO3381/0BV7MW+Xs9H3IC3lOViJv0o7uj8JpCBZmSadC4evj
0f7FUxLq9C6c27kAwONNRBpoPIE51nFB2xzSaUQkql2B7+gmYdnOJJlURXjGqU1G
m9xj8HlUwTlQrNEbhie5KbXceAwQmyS8mnImCIn6tJA+gwfkS56QjVn6YGnRu65D
VoH/ZSdAS2x7CrwWL6mdEg3k8XoRZ47VmihOmzGGYI6ELpOEKtmQAT4w8GGybWvW
cbTvZgfUIZBtupBc27StkYFawIWdLjcHwS6YmCnpN8NVZwBlkLNdZEM+sgD4Px8/
aKFAWDW+wZRS6Nr/vDJaKTb7icnsrvaW5uQUMiG0yOMF2TL0V3UVagmF9VRFE8x1
Fs++n7cAd7qCxdpPgP5V7H0IPZ3j1cKLVWFw2KMdyJ4Dq5kxuVDnjlqQxLsKEWnd
0yeiSWTw8OJBu8OITTDy1Cd6MHRhGV+eKVIkDToTNze0H7/hw+gox//LKJy8JAy6
oc5QttK0gpJFO24YxB4PjS8IcDsfmdhxcR0Or33xS41ljFIP4dtoLxtiY1MKn5WA
8Qw9dFeWTI3cIXtGxpqwQgBQAynVEn63nmlblcnrZL0ju/mZZgQvJaCNb8J+sEkY
0DqcG6Y3gy3MaQTWIMxu9m8Yg77DJu6Uym3KgEwqCmRdntfHxHTu8UVartf/rQjV
UoFTzYAPk8puaO09BVBw4Y8LG7xUa2AlOjXJCd/M+F5uCaS8LAqIvV23UP047SlY
54WH7sCI6vgS46xLluKmD9sg5OAzyrZR8kJUTw41/sinjMn6iv/KNU2nuiXiNxyZ
B8l3QFf6exYwk/0ey5Vo4Vhexkm5OJOu7MCVQBU6DFctqq0tYvO8bCliks0cXIdi
u5o4MusdVpKnWNb1vZCuWLUJwvvjgHueN7T+uN4rsOZG8LeRvAq/Eq7MoDonfxa1
/bKvs6fLImF3OR4hxriJ6k2xr3kwnln/l+GBuGxvwb82k6GcKa1WIX+keLrrUS4O
/x/SK8s4Hgz+0bEBeh32kKt+xROZSb2iJor8esi3WYuh1t14jMzK+s/fl+YCvh3p
fwqkVtExaOYd2R+QwcmnIJquCbTXrdydswmVgpBFVU+OLemQ8X5A/0CXx9oo4erF
QoVBFQ7i3rl99dVvLBE8tWOlqotQM4/Ac9r6qGJ8UEElMAtMRHR33vgXAFvDtaYy
1Y+Gu+D6zXR2nRwA7FRgX+2oNpUaF2h3cm+tEL0o2xR1I2jrL19FuNoTsR+z4fwZ
xEqDFgu0Q9KGTDBpRxE0BoDE0xtumiOOVscVW176P6TIsXo/X5ET0SDSa3NeJjpu
/gzQOVrDdHy6pz7E6DIXwCa0ciYbxR4fv5CbjO8IxUPGETBz6O68Xzba/Rci7C95
0gvIvxpCzHlMYwjAy+DjECX2k6weNZjR02R6zxdh1MinnProCPGCKzWmvVXO6iq+
k+jYb0EGP/RNsh2frMvTX7KrtLUeWEb6FDnoNsLH9LgDRcR+Oz3CJs5/08lyl8G/
94u87bUJ6LZEKoGP/OR1cL6DruOBsVTqwxVV6SF/c6oEFaP0au4GbvrLMOOJqQT6
s9irv70ZUOnzKJiFnwRWKutyLsaWN5AhNFx71WeBEJPE+rXdKZdwGD/L8k/F8e/2
ardfkFAYijm+7+tC9wllVmFZj3OL+X4ebCANzGctnP0W4h7N4tmasDctzxMG9BhM
hpo5vf5inQWc3coM83Rzl8I90SUTe2sTbp+6U80/w8n10zboGbRMK+bHzg5qpdt0
N3eZaxAhxyfd6PSBv0W3Q/NhEw1yKlA2nfaaI8sRIGwygWH38Y3A9DnmTakrNKE8
Rz0CddH/UvTfZAmR+w8HmFLraIvXFHQWI/Pi+dWySjC91Oc91Qp05L6KII3ek4oe
xCFW7zZ1TwwoIYOUbpr0j+xnmMWY2am2kntoBpaiXBkoOGUC/+Jo6ocp7C3Xl97Z
+iLtJfmVq5X5YJcyCOY/DKRfTPxGwnqjaX79pY6HtXa67odeputZgbRrjHAM3PFZ
aRij6Z38UUdqGwmRACBOM9+XO3gxfDJQlAhWrucH/o5BEfqghw/Z7NnoRIdT+BUO
7TaV+Nb2IHIs+5fgIQhvbQh06pHvaTykHAPdIfVxoZKSsppvH/8eMeskeOigISgO
k5sa7X6W4OXGXZ+QdXfZVs1P4XBbfZCmnqpqEsi5YzxcRKMM6WqmLsXVlAp9wdwC
fOQegWeB3Lk5ZEiuBdksbdbSxifQMt+WYQLcQqi7Bdg5ktUD1oRg5ewFrsoDp9Np
B6SmhGhcAnF5uA0ZS/FQRJST3iosjmnxdkz/YILLdn9WfyPibEl108Kmk1+jyQv4
SiZmmpccA2EYzkiJyTZloMEKdSXf2llnKvZYvAQqrRXJHZlGB1wjOF305yoAl4hI
qQnrKdgHpFwSwCK0xhiwEqbH3HL98mpUSk0pu7rGbkp/PoLT5Kfz9QbgAAZiK8mZ
Qbawvl80rW73MnZj0RBwCPIvCKk5ByY78y/28gQ3YadJhLVCsL2eWT5pjfjsqTKe
jOWRw2VOtci2H/zTEoYTeD6IslvsfbnllQZjEwIkk6KeNvhG43v4IJjWT71E4Non
POym5lgcTZ9AQcyrwUAptL/3L0brxlo7cOUrLfQp0haozX/1nmw5SAck8cyQggxw
6NdJnyQNH72erMrVJbCaQyc2+r6pQZFMTrIsecURt6a1pJPGLKBNWxfQlKsVNW79
eK3zPTY7R2pQUXQV+RFieCLgwEmmJwZTb+9D2IFOfcmBizLpIrSgi6KY/YioUBwe
cS2ELP1u9fgcMM0efNqSSLbVOzfz9hnZRZJSmp5DfxXbz9k7Yx54ygfkyacnbcXT
IhBx9yaKeeEsu5vVcLE3CozLBfSb57GPkedli+7hX+rLPyF2v8ws1rPDTZuQg34W
Lc9vU05kimM4c0iAoLfKt8Oqeaw5+9VsGzOM1yOx7Nscf/o5/X+8/tl1umdBQWjW
N/cnoqU9V68N30nIw9xWKusEgsWMWuSlkyiZKTGG0v0tk8ZTqNXYZaUIRYgR4WRY
mup7s3/bZ/bCW3SDXaBfr/yAr9jZmXnKCDP5X6ihNKwQ0cn+dl1jV1OBjGwHaN1T
ZBtZg4HsrpIjlreJgYoI2ijJ3XwL5iRTJXiFIaPIkouksnzRlGzXGlycQmzDKdJ8
IKwVEwcWU6XfEVvxeLkTFXuno7xKtcZjs7JgSOMulQfFSAe0XbE7+zPL/WwIsYxO
RY2nx/ig1hBOb88Ht1Tzsbq3bANUJoxUFluLzBlgH8pr9Iyl1EfFBGYM4zYNbzEe
UR/nGQoSsRec+OUjzmvkqGYwy5+V7pt56Vm41ONl01yt/rjd5faDe8A711X/zfBs
/SoVdFo6JFFz/hRnsLsFuCNNQl85RVIh/DxWnxG2PIS/MBvKItdIeqjNd9DbdSqe
tmnrtdy6IE+sfG2axQ8WE40UU7iGjB1W0Fq/BVYQZuxKuXO2RUYSkWtpIdpI1p/H
j8YBkx2dCGyS3uhRK3k/FJppwt3Hs5uGImmmDep1TiN0vCQmZCHRNGJ05f3DgUao
x51iqxmLghGlRf0Jw9k1KRTKnk2ep/Es0AZoX77kf70Lc1Yk+zR45h4tM0aRO0RY
Y5s+mgldvx7ixL6hgT87rP0+7/o/yoV0CFst6o/Jh1cacgqQncXahZvS+o4eOQFC
gjEzgJP0EJWSd8yO7j5gBy1px4HQ3M1KoUZvbC6Q2auppNV77N9emuk1WB+ozP7G
KEC7USwWCFrars6VWDxCZXIfm/xOD+A9noJOuOLCxw/1yLswZjQamrXL9Umywy49
/SF4wLqoL7tePrgZRTOXvgMzoQvUrnUQ2q8r53J42MOrozzc9wAUhFxB0yW6CGRr
D4hj/OYWZ7OosaT2zDhmmxMxCggcSoAwD738lsDwmddpqtpavAGzR6e2a7XaJnN1
yBkZzFlQZ2j3UC2M0YYIFiFIViKEcEhpGtoTajdBNsSwA7qjPQPo5mP9WNGb9fQL
Jc+9F6RfKdP8MquK0Iir/wqiTWqjemyfW+dKlZ474SKHqAD5akRnK/ExPWq+kWZW
zuYkV1A6MEKoQcDFerWIsF6GAiNAgx7zeDdSskZ9p0nbZuFTk8cSbUUSE/r0V90N
ndYdWNrwS5iYZ34+z5IAE6TeuahG7jIktm23p/56twWt4bnBIm+31h+zujLbOEqn
Aip2r9EPBJGUMsPB2uXWbnEUy/vggPCZTopiWA22GuniSDAdVipmgfu994MxjHXt
45cb2ECkjxP6TU5Zn5SQSZPZ38cVqxL+/7QMC4q1IYyG+KpdKqxoJlMjlpz85eQ9
FZp5z436SBhFeF05HD/syi4hEMpwh+e0Rp9szM7bG3MnCKiHZPtp5oW0CWDsS8ed
r/+gSMsSC+AtxstJ37FAMkGnqWbnh5cgJjzLx7W5Ij5BAhMug+V3QJEKNV5W8+up
1LxWi0UKjRsv0B4zKObIMko7W/ksJGB4JOf7b7eVIngz4HKtdUe20BKGDWBJ3GND
ylTd+ykml5W5OCx0bQNn9FIYgCMYMfn2Kqw8mLMnq287FDxdaftrk38Ghzukm03r
8aHTu1bFKXalE0+qJa9IxgGq/CRHa/psYPHNZSchavxv2f6Sg8tV0+PtlIJ0/J/S
VQD3af251VMgxsCAI6nK0u6+qno07ZtDY9QBQMVL7VRxEbUTiuTk/Y55IjhgE4ZO
rnwwgdj73c5Y5L6XSa2fVGRT3oQEf3EceLdoMFQakNHA6Y52xk4KBtqJmOww+Nsj
0tlJKqGk5Pjvxb46wOE50nyx6OtGAwdEbuRyeciVxHxMU8DFjQBL7uEWDMWYLA63
p8eS395hNGQJsk8UJZVucXDWPvLsACmbEgQVl+X+9OLAiwXnLwiubOyFtLb84qEZ
sS7iLU0voowU1S3TmsCGnWftTwuSekRLyyxsn745o1fkYE+IHStI9+C/ldP3Nq80
Se88WZALrGWEk3MkblCiR5/juOGo8ofrTLvV1aXmrz8pqwKnKTo0NrV0AFgvLtJN
/9T/pJKC08nZOeUQxj85HsMSOOE+5NxoFOVy3vkayB5yL5ZgN6HRcUQ344Kc2CBd
UcqRBQo5HFpNkF5LrXrF/AsqcDPBxeUrAnMZycMyUQYQ0nQn6UMtyMd465TI0X44
4ZtHF0NzoVxO0922TL4UlQB4Lqbz4L8ZskJbZJxtrmPIR07J0hWZOpkAXDY3/7o5
R+Y8k+bCjwLMiXvaBe30WA0CLWymO5Y2n5yay6pyhLqTFIQNeTuB7Pq/t0Yov4bP
vaJqulj03pAdx1qFSEYTbg8r1YA3+w/WeY7CzV2vB5NOgIsyVKo/BZaZcGkh/NOD
P3y4K80HqrHXVdCadiXPfaXINpJYewPbL3pEGE/O8zg1k1IYEB/HAXmIU8ANlBMt
RbJR2toWKqd32KaSkb+SupwcMH2dVe212Urz3ikKt581L0RMu0XM5WQ0taw9KHdF
NpSrXkTUAiFHQkQK4Z1vcxs7AOSE8RIW93k+KiSWSpI7pH77BrJ4vwiiOdh2Sg67
DIv/pCfpu/q6b7n+7OWS83uJ6Bhw7qFFWmMOw6dS+CKtbY6VXGFDY9Jt6fPsPf38
D2gJmrxFB3nYV/HyfTeb0R1H/b/q1l58uNndVXoJPvq1o3gfaGeHwwXrYD192e9V
KNKuoAVPHncJqZorQ+5K2KJsXzFLm1stCbL5RBTuAG6VhQHXZi3SqVRtr2FRGJda
9zCc2pu50+U1CCkVBlIPSNVG29Eim2h2dTb1epdN6b9+865itfJbyT9zotNf/mXE
T+dYROv+Ph8iKAiQQyND0zqxG1Q21q9HdqpvEXa/mPrSgoAQC1z0xd95+wnhMl3v
0fB4w1gCSFyiBZ820H8HUYBqfnh5xQ5XRUmt+HyxqOKM7U2KOGGziK9w06aL9UPn
wtqMJ0YN8HFhZdAej0l05MuG1ta32qQHbR3WCHofOgBe7YDTvU5delVnwjIy6pYU
2H1lk5uixZfEBibeSXPYpchZVR2ReQpIg7okYQLa09F+SKc8tP0avL0iPpEvc2zi
cQbdSLw+Zkpi+3zLUBGYYkbhY7Ia8AUnVXHJGnbqu+Kp67EgsXUbT7cM/ho15cEd
b+iXpkh+05VrvbcHHcG7sMNakre/y4/NxzWkQdykOR+S7VPdsPhSTIbsNubLifMZ
Ohaa4vsDKD8p5j9xQQg71n9k/DPqqRX1NUVc86Ko3fCdYR8llV0z4/jm2yvaTy09
XlC+i+WoQ0M0tl8QtUOOTZpNYAvu6/b8q2KGzTOvC6dLKQD31Y0v9l3WwEYQVi0J
lQD6THa2ja8VGm6QSGhMxQV4c9c3ZyoTBVyrSr8/kjwUeyUkN49DPFBHj2hO74hj
02gFC+W3USOfplcnN1Np5TMPRvM7zm2XgjhqVTQ7+N52PyFGtQfaLG6iU01QC+EX
604I6bxvXqj92K+evwEhwbDuE9rf5wvDLdSoE8Efmdp36LSOL7YEHS8VcbVifC2A
GvymFlN0ch1QkiO5GfLgRaA06tERHzubOihMBtVGvE0+hM52e2FDeP7aZ6TwGUQl
Q97vWEdZLepRz5mqCmVf/SSG/+c6DQIYYHqNT9CU6tNbCwk/W9Nlu6+CVlE67jKm
VzjEqO5wnCmW0ogNXbqWPgHzPe3bJSZscTzD+TqnLKidGwsJ01VJeo6X+9xq1cyn
cm5KaWGLmhzeB5usBr1EwoUuiRoSXgtIUQ6jJgkC+AARPUGA5cIHe7nDfFr/IWxq
5kz16X2FN7dmiaE1XLppM3nf5VkU/d+3YexZ/IhwWSwG5tU+v2hr175yX2YPjww/
iAArdRAtAxxEEAjAjYmz+5LCx6YjvU3oGL8iC0UdRySKVldNXY/48+35bpnlEDJr
8KLIL6Er5Br/GkB1txDgJ3t6BW7Ef5tQ3b6wzDQnf5DKVVkpRtlMBB5Ab+rG9fE+
3PBgU/CtENL1TUb+Oix14t52lbtl5k0qJWgT2gZggvvqQn7LX0EOflHiCGsyRo/T
XoMRYdypcWRg/XwMBG+gwYvRBwcsIUuoVKwUU+dVNa+Vb6LbFKIsncV4eFORsRlw
Y4nhxMdLNymNRtcnavgQZeCqlU+G96fUMRcGi1+eouAKOmvep/cnwpM4DaBLWYoo
vlabXTem80aglLUGEAhbV8TIpnATStxDVR79KuZemC6XfX4YAAdUn7U0Bsigghsa
7rB6cX0hwMRwprwOPGchLabcrJVdFiKgFxgRbqXaBZtix0I90zfIu7TD4L1aliko
wslsngypWCkVfYYuQdF4q9chdGagVSo0A2H9hcI98IVk6DVbJOMpVGB0PFlWPcuK
yN42uSY10R9o9Kfi3DtBJY61L1I7194nz7yBo7lEjBi89wODB8qVzWONlXY6qGjQ
W03KS0xCak4oqBFLq6qkfIDjEwrp2lqw5qfVi9gjGwGGpVFvsv4j9qReRtHpAIXQ
uc4QtGvrzzPem1T7u8Cgr2Lp1AZ8GLwkz8ZwIHonMzFfSOZPtSrnIso1/cEYSGk/
FusNDRtAnieRygAGJtBJGMa1I7j49yoB8z373o+/krExs+4bdkYHNb6wVTHcf8p5
jsOrOMrebXMKxxKjMdcsSLvVLHXb+hEwGoNslPQD/87ZA+GUq+xvPk7YG8CW34v9
//dmr3L9mIBUmJapNLvACg/DxMGZceIGylt7bFLLL7YW8qlmqgVzJj7urpFEmg8O
bBDGBJP65ArghsRsWzBA9nInr609+Dk2SBnYWT9LQAR4JHaLPQWZHvcH9HPnjBU7
XJwQ9DOKmN/IdZjR2beCA6yPUDFsMPwa8jvkxKCJQTFdO7YCqbU6BDIWeIjoZ+UD
ZU7saVlkxUreHBJff1Hs33ITwdGu5f8XOTXFwN+zvRCWOf3Plzzja9OZXYxFgrJL
dhFxnubo6dTbllRsDMCTfmjTXI/JIUTJmlqzTkE2U7S4XMfpcdkWevTxOm9PagWw
Ey1nyUpe8AIu5kquG2Ecyo9da8KBhhZdiLfR+wY7CA/PFmVC3BNLZ6BAoSSeIyDQ
Jw5tqr4muakzg3c6G/L0hzrjIFpb/1ADKEwiGRzKv/iP975ePNrNynLXyqCfzdwA
lcP6C6VFdJwX+ek1qHH89kS8QFdAli1P0bivlwf88s3cZSG27oV8E+RiJHo2PqbV
djB2g//ATAwZDqJzC3GvgbvSAUBBt3HY+DwK/sjCvmdlLLdRfR3Z2r4cK0mKQpU8
pvLxaL7PK6S/Z0QlifO/vqRnnMf/aN73Jqz+cUVlKXEoN0nGwfe5M68ITlVKcpG9
ze06oCCKaPAUtVTlkOwiSQMhIe8iRnrUb3w+lg2NgFBPNOsn7rQ4b4jg8T0iLRG6
Udf5qMZsnPa1l2O54IZf2+Sx4+NqV2sm2elgkiomNgjZ8vlOOdQH5f+V74c8yv//
fsjrS25yd0UU8qvhynR0KePNh6Zxf0ST2E9Tlmn0b2/6EF7JcQ5i3jzk1sr0NUWo
FbMBbn0LjZFlTD95VC0UXgDrMv8aVQuVzS+mGYtTehMCb04x7hE2vVxN9ZqlHxkG
3pVmFvkwKtNXVoAPRM4hk+sxrkwNyotpg9OhPsCT6kfLj3Yz6koKu8IXSE/ySHQ3
FKVZp9JpLSfr4kB9SOLq7Ux+pXsMdQiW5WaE1bJg9ut6DpXDp/K9W3C+mJfQe8tq
MUYTtRBNiGFLg6PDnCwuKydEqt+gkC5OLhhV51pjhkUxxh9la5oReJku4FY08V/Y
NXZR3aOCXxh2OMsYQprV32hA6dch/Qq7gD/tVs2BL+7rZbUfv5YZ0XoRv7lbX9e7
zsWUIUMYA2b/88XVr3RVKRGKFDNuZ+Bn/rbnCfaldwKMF/+WrTl4PaU206YLm7vw
YbosqzrQQSXhK/I9AIKAqWqkEWtnZJm7f5mPP6rR4yhQly0ugdhUcDVsWtERrnun
0pZWQ3Zhvde+N+hQ/DaPtDIOaFKjvXaVnMG/2DTVazQAhiuOQp77TNBMLI8/SgeW
VNMIQhuzOfwS4Z5SWmZQDVVv+Mkn+PldK+oK6/XkCluZBi6DXi7MV2JuGebzC4Hv
QlmAbnu4A8rmTKMRIBJGY9Z7wiPkR9+Sc+4ha3as/834D+8uV98m0Yw+lfTwZ3G+
qKIPgJoy9TZumoj8dpWvcobihcqKbMhycqsu1XnNQ5qWnbpgl6oWKBwk/AVfZ1Gu
HDD6h1iD5u69i/YVRyC593Z0FBp4SHnCLBG+uoggsEQUCUBHv5uLzp4k+DRXkP+S
uS4oRpnHdWshv9RWhJTewD4u+gJ2m3xPR+RpuPOgie5jiYAGVAtozvzBqlRSRPUY
L2pGTlt9YVgnqVpDK7Tegi8DuQaTXhDZb47kNNxg8Sw/jOZ3AkaOcavE3gOzC6E5
NSh+7RGs3ZQGVTnpTdFAu3rxLoBq3Ih3VOXhLz411S/R/y0100caSUo2jZIC1T1x
e10JEasezFgk8dCzM1V0qmwpD/waL0rnIkYjOiM+d9h67DfINKKZOWUAIG9L5VFs
qlQvZzqrBRIrBWg6ZXWirlQ1uaxsgiERiIrRT5FNIn20dIImnp1dLSrEljAZf6eE
neNB8QtfpGbEfG3Dta+4Y/+QbgOyEZqshNLGFAmpEgjMZ25jHJlJk1A0xrBF+Jj4
3+T9bRIHptBnVLnG5VEA2eivXj6d+SZ9x7tgVIBbpz3sFO/x1wXd53/6hjWtwQBH
R3CN4xcZQyM6Kpp+cOmhWI6phH96EdmEW7xTYyfWnSMI0gdvEob1GFy+1qTH1O4V
8J2vcEYtx7I817PA67nGDAEizlhIioOSMettRn3XW9y+4qTCfId2xGKI+Hjvx0rM
D5nnNj0oojwU9FPQNQXQ81HKRK9lKDWmv6MoXkhvnL/4VETH+UT3lDNG7hDvqW0+
nstxnWVGD1P+QP635hspoACfQIR0VuBvNOl/+n0RpGUVpqG5M2A575OviqBDRu80
vd2kfQktPuE2vpfI6PvEaxIDSMysojgelDheLptSzgyeZjoOUg34C9VzMcxfQxSY
SQ9XOt55ZJDsZ2VFzb0pSCsxL2cu437eWAZ9JoH5ho6+nCFrY2nkGCBlr5foDgbd
KqISTMeTbL8dORHGFwXC/xtXupuxBNv6RUwQ81ODsMO39P0PnzDC+7Pm5uuY5UcM
B7MoiMkFYp5dpkoM9XITTh6mduwl3Yt9Af2Y/7bZEhajUi60FP0bQcGUb83Ol3Z4
+OrrTc2/Pz4UHop2PsXaGY2LUJpfV1xxClY3A1eaj2+3P5eUv0SdloPtoxZBl44u
BbS42OOuasQtjm+HjzMRcdID6XYdHJ2npM3Srw0JfCiEWrToAd7Woz/Ej2AmlAvj
p151t5kW8k2yfD6Hzatnh+TaqkjPWaStZ95WkD97oJjeZJHs8wLp1by77EYBnxlE
dq3WCYpqrGNXZ4ivRWqXBUQwUrnbmSc9Sb2GSyEK6ZXPjnV1QDk1o9pp5tGp73v4
5fuIH5/Yk4RXyw76yvFcD7GwL10bhQ/uMGMB5l1WgsAStKxEviXFrBMMtKWuMFbb
3uKeViXZ0F4rWNmRWiBmGFpJwRIzdpi6OBwxnnhuoxzyJodQ3YE+6tCpQ3M4aipE
5z2yYtnn31A7/BuVTAeQc5lrPqNPsVCAOXhlvPdUu6ugsOoEuTRj3ZN77bWKAbWG
QTrrS6JRAZ7HVPtCnOlwuqy+F0KOL4aPMg5TheMHYI40t3lFxYvmVewW5Q2q617K
Djn2peFP2cpemgwyXnjcjbG83L88vHgFyP6iiLLyQOSV9+oYL51sg9jnoQpH2yY0
MXwtVs7Of1tbfrNTaa/l8mzRtWl6yi5sfgGtVwkoVCeBAU+/3emUJnDyiboF5Obw
FvJGzLjTjv6pcM2ihP4763jpe7zNjkQbuK96+OsOJ3+AvICOjT76e4UD+DncnRoA
kbT4czvk+scfYxdiT158GRzhXRqlylOeldQ8oEG2OepmXu5FXMRZ2eXKgza4tKyA
Mkh1VsceczDzbzMxKTp/VX76KDcgYb71uUI8to6skLaksDqWISJV+aRDREG9w9fl
naANbdBFUa0OwdoXuccOJQ2bwsSYa4HJZl+ZYSuN1nekBBtA6AMEMV2FgmENHecZ
ry5PoUkHSszzAWCMGkI3Tpu9q8bKnbQBhp0quD4oKGu1/O8a2FUn51/8g+NNGQCL
sPFPAcWDmZhb7zC4e0REAtAzxDYSYddgKeF3PXfMlg4ROETQoKaJ7HfhgEsASvS5
DP4bj1UARMypAebKmIeFpgvgmsmgmaKFi/qXGXmJ8rQG7PocSHI6+W4JtkRa03me
ZDk/lkIKOEnFDzBDDrS3e38yGXgFjmYwz3/urKA/2jkw8EvFEnFgR02KdGDYsxJC
ILfMnumM2CTc4ZQiKpSBgOQNli0zBVBbWszKZzrdo9FV0Yw0iNGzFOYo378ZKpER
vR1FgARMp4Ub17xQdkh59c5/zrWJ4xNF/XgAGWS8lX+fGyygb8Ce9Qd+uk1fab0R
nt9C6Z9HmELpWI+kgkUKMQ1LR4Bs125RJeuzOIUR0WLCmj53VWsgPnxPCIYcb3ua
mzfhf6aXdF5rOlJotDytMzT7RELLlzTcKZeQ4zDALx0dc4I/cwKHFor7hLptHeK2
+oKykfDhtVbe0HtuwJGaKBrYh5mNMh2+RSR6Vf/7yyvxPHns4o0X+TNs05luxTCd
RhuDJn+sKZdumbUHJQPos6CsGjhZYUHi9V/xYyV4cmeMrgLaT4qCT03tN6d5yYd+
0Jf/UHBE132z4Z+ygl5nvo3Z93zE6cjzEkbS9phAEyQkWN2ythdZk06lBlJYEYCa
D5j2emDXe3o3fzMsw5fEJIWayxtu3gaUPWqyuC1pQ2beHGfcTwMvmvoaVQSxUoV7
LaZ9eY6wzz9Ui50CXd6r60HWqGa9345SqItRmCzRyUg2o8RuKFAgCxysjlfNoUu5
xoT72r/FjPYtFbLkaNmK830NcvhxLXwRXM5YvuOTPQ9jbC6gJgcZ7yOXHFpNQXp2
91g45nNoQWJh/lualFDGH/VN3XlXTvXT6VrPeHuBGaqZ5TcOtTfaqDZ8LbA80qsI
5tMTl7aEtyO8tjg6hVUgn2PX4uXdePOhtjcei39cyLlbjSOtQJ4zR9rguVe/LNqz
B7mPn4aNef0qEH2dObCQu0SBbnjZZmxizl1oz1n9xpT7YLqr0s5peGG77irrOj8m
sjkt3G2TUCNRYJYOTFDgqXJkT6ey4J+hmBizQEVWfu+7pdAzHa7nPriJnFbk5JkO
ao04sZ+RG5Py2BXgM+sWg27LA45AB82InY9HXjEUHHkF1PXSlsQhIkRLqhp5bCSG
aoZryHn/oNzYcn8e4eSR9rvIgDp4pmuVmh54xaDmVz8mkbCuva6+dbQ16zS3XBJN
1wsPQksHvAYelUrrHmxRqxXqvdmF1qYfXlelhXehrvE+OWuvzm3w0u+z/RbawpVx
Lo/7pbP0hAZge5wim4mvMUFSFHYWapCzf8zMJw0mjp7ig5ccFgzPxu4gPx1cZYLQ
39jNf57iC63u38txm+AKQGMzdPJwxc50oAXa70dnOLBDOjTCkjQ3tdbl88uCZeSd
rwfZlwtODLy0yXX3qtdsQsUgfBZaKSAya3CArsI1OSfq0nFPil1HeHq2oHQxmtoO
8bWGI1bAWaK6bc3al04i6g+8etMEmuIGXDBN20x8evtcjC+ipAJz9KoeiP3RAU5N
7uGoHb0pjTIQuIgHoXVgBBQVf/r9y4imvf/B3cBGsNKQ/moFn9BGxxz9dm8Nb6J3
/BV9VgBtmx83lUzVlRO8Asis3BrXsOOCTOobiAMopRdvepogBtCjRV5T3wITcRCo
2rZexBmLkd0SzgnbefzfXwfk1ElBsHn8QKkiJ/3PPpcBSX9usbUvTKnF2n1s+UlR
GNrq3atBf7ieL6YFSDgfPVoYyrhsnLAMRIog716QJR/jAa0dXFGbd927uhBZZA/c
q/DAW5AztTtGmyan7leixP+l7usBQ1dDZuZ8hfHwvl1NcY7gvnQTeaV+nzu5v7jy
VJIDQ4PJVMaY1ld6TEaIf/3/A5zoZomeTC3gtlNQL2tHHEcHAVdhjoM92ti9PvRK
iRFn7vrRUaDitE72qk+bXfVbJP3JBxEP/4m+0Jqr3pT/FYqzVWFl/BA9X76CAYux
1DIQtOtC+0BFgNXS4tSxpYDkvBAsJvRWfBpc63o3u1cCfguXLppen0/EhPLL5Djt
XseKGBv7zK+PJzZGy2gQiwo1AzObFoMaUu1KeS1mwmJ9CTR2gFUkxRidpNy0pFJe
PKDiuq+Y5V+0ujPBYQY8VTX3mfuxyyAr4sw/uWKZUq3kUVsPXYgT+TKL9Y57Pm0Q
7GJDohwvsWI92lCqEemLVdGF1bNgvr0Z/cQMybgz0c7hRDP4CA6dae8xXrUAMNM8
SjUdnEKKXEutdjKk7BiEVjtbOhD633japdieyymDNVd0VENUfEa59F3IkTP0TnOf
ZN3nZFZOpu9OQ/0CZGXusN7LZL7Mh6XpYKqEvGlYJsEWe2wrn478BTkhnP+N8IPp
L/txiUaKXiX1vrwV6hu8z/6LdKoWrkB8+Cx/LggfvhyEiXhYueweBDl/tHe5xprJ
wn7J8TOzcXGO2gGu2wzYt4K5bYowRPLHN1CD081fcTj4tQlgtp80wa6G3gFu3uWG
rDqkhyNqIj7RRoVreqY2RY0fFsq+9ia38i+inxZ8OHdjW4CERFLJHm+ZN3k9gnuw
IHi+fvh2Cf01zDAgLU1CM6qcFGaWKqxVL4y8MXHeQ9OInj0nyIiPYZLqNLUNX9RZ
Bl/y6+TMlxprjGSL3ijz0bZmj964Sb+NcspEAz0rOmhsxlI0VKiONL9HsG5zOvJ7
z4SZucWZe1+1Y+mEKU9ON/g1f8UHsxAIsl6UrjubuRJOuLgx0dDTfQhMyAi1MDrS
M/OjmTaAyyopaDJbZ58+Ek+28MoE+WxVpqIVlCTssBhUgrv2hfKKgzqc/76XsIrC
f/nOsFzWaDeofEPa1LbyTox6OA7Hy3hWHzq1tuOWHF1ri8YLM9tQnhHaLRNOa1Jm
p1pBmqiQpC60UrgG6bSacHcUjby6BO4WZkMnO1kstj//BhrTqwN3gn+E6U3Eaw1g
Tr+cl4du6HO38Fr6V+6bpbK4lgfP/KNgnMg7o8haJaBdJ0b6hXEF3KMPaS+UA/VU
U7FnoZ7VnQCYAKFtTfvrqwmlQwv0ZrlSVtXrE1P06E0VEU5hUvcxUEKfDyZXexRo
1jUbGOuQbDsX+04MM7pjJZJmA1KFqmHWQJNLl1Xeyl71QaQC2D4FXYoMvrTXZ/kh
DNK9BKjCkJtamk5fehBcfFuKLFhBU+2KUw5EWxYdbXq/fivdBMgDh/ppQj9QONf1
vP3E+UxTdNzG56a8adV1Co4TbWVqhHkMvGEbkEJMeBoJ8YqCg9YW2wLgPggMiL/U
i/zN/3qo1pFj2yDhMPYcaM6REmufRVNLAD84RoU3ibmBqr3QSCU+m8czXdRMj6x7
8B/PwaoUV17O1OXooILn+yNKFghpU9t6w8BkUYaQZzqYnpayU9QFoflQ34oQHYZW
2tOOuBhdeErWFPY2tnjdgRY51KCIobkKl5v/AVdEo2+xNklIxxJCMjyybYBm5vLD
qzkqXORlK6jbU3V9Aznqnirzk9auiXO4tmorHWQ8oIaOy+Wn+OmcqAbSxHQhoo/2
WwuF9qbASpy3lpFQ863CWudTZ/98/sEPdPQgiuh3RM6sRWIMnBfXouIbDKdZu2oU
gysaJ/4ugr7Y1GbMKyZijQEXo3YgPhQ8EYPLHzfwRBR4FxorDGnNHu63vHCOn/Vn
UxOsiaVtd1ZlMOLD9xlpccop6ZMkbjUgdpiTZPC5wUU1VV4U0NkH0ZdWe+8jw0kP
3hodKm50RvId3A/Z3gUG2csDR1fIy2u9foNBUESCCVJ8DgSFwqSyYYNuPXl27zhQ
HIkOyBsx3z3UIp7A4Z8USePcGT8y+kNdiPBhl09RROmwO1rGfMyWZahN+TvmuF4h
6l74AbsStBIhP7anVQUbl7pBnPMRGuNJeQ8ECZswE6QWQplHBAlB5Pkrb8MPt4pE
tjGp5sFaMV8Z9RhWoMZfuYW7EGEKfV4El2qTg2S66g0upze07wDK5Gs1wzr5/EjW
sZM6+tnSLhlwE3cvbdP44+T+/Sjz4d812EtFG4oLs2CXfiD4pbN/vIzjoqCT4II4
UndF2aDlvaCAXy8R7Nq9xSP3oNCTnwBrILIq962j0oIOnW1nS27Xq79kkrbbMbpF
/TKRxWi3OF0W1iFMFY/qKIZsIqRnkb/lDUXBfFEsMVBnh0vlJ2C97WXTw1hZUEx2
jgjKCrnvk54CGqGtav04wFPEKMqHRJetYeRKGFh1+LOqotXgTVKB7EPgSyCJH7xi
sIR7FKd8dCVWsqWHmgVWUPoe7GwttMM1jgh1CiG2UrodF6kWWhp7KE02oHlUsSzf
HLdpjS33az+reP6Nf/bm0OPXpP3YLaETC9pw8PpY7+p/6pjX3vhgLuCB/23T66dj
SCT73oa/vAiO/piKG/e4fj3+5LilhsK7tfFh8aIttS6piNZfPJpYhk66il+48RlN
PzUc6WUwcB7r2kFj9tZY/WtmDcOoSeL5A1cgb6Pl/Pwf/Iq03vJjxhQ0xhvCI2sm
2Wui9QBWnOZ/gYDZJj6LZUyPpZ19LdsN4Zmf90xxi/e70Ax8WqxjJAVHyF10Vy2+
hZPvC04sxPB39olPQBhYtqGaSwN34XZdbxttiF8hkhiUgM/IUODonCfu9gaRCD1/
kJ8B6jOsngSXyL3YrbNkwi2lnUh2uaDIBDQpl9S6nmcgALwiyza6Qgtk/+PrzgCC
zjTSzoxUMp5m1DWMBWYBS/mxf5p7u4xfxvJbMn64KOFAVuqT0xdgavsTeaPLqoji
hjFJO4OrgC+xKCv3TY8nKpK1hjOaXK1CG2FeFNldtchjlEhyTcwEnxzP9V03/W8m
nxMmiSZJ8P2HtKNA9qCJjukwrOQWJu/pGKBIjrz0hHBxwByDHYTNn24k3tecLF+0
bCN1FVzL5GPe4C794rc8evoEwrvZdjz9FYntq574ChFiOcrhJ+Wixrm1L/xrDk4S
OvlWBEmkEzy/KB74/7PafpwAxE7Eg06IuMSPW2UHK9dPvHxf5cJyj0nB8L4+pwOE
XtM6AtQIsarjjLmmFHIx2cWQjhwZP/DdJrI188lofr6dE0d1P2vcycLyn36/gpbU
mM6Hh/6aNh8VSFYhAjoBB7Cx4t3SMnp3wJ75P1ZdgDUhwiq9SOgAinGjDQlRl/o8
5U8AT3mkNwwxcjIDrDconch5ImuiinASPI7T1GwJqq0sGZfwre6NHiWio4LQRaoY
p3B50te17Qb9t7tC6DnHReFqhq9wGcw0xvwBUx+3SG+pnMBudXsRcqnNBRLHhmP8
4CchGuHw2xg52KhbKuIFJjS71rIxjSwQcsd4ZyR+bRnSXYj7LFuCif15Iq7xRlYb
EE6Jcds3P+Xomc/52KT8tvbm3esBtawYE7CMYfae85o5HldcTMnp0+m0mKj6L2NA
wmudeneS7x5vaYTVZwWzD8Af05ILbb1xgwmLgP+OCxiuBF42NMHELgZod6gbPo8X
32L6+nxrkB4C7bJzjCdNzmrqcy3y/1w6HXVqO+amsPik/rgDUr1cjGea5vqX/yza
LpRp9CA721XKT8YE2z3rf+LxbccKaZ/IB/InOFE9W8t6jlAjefkK/u9qRp6avt2F
M/FMN/UH4SbeDpbAaY9//SzQcifoqHiY7Q47ExiVqJ7t2rULwxNAYsc1PfSdWAP9
kcbhi5IFl/+oKZbxjaTJ8d7PQK4DME8esvk0Qt0zHcWwVvEdVtowPGGzMA8OvxVd
/Y7C44hTdknQn7/mn0bP4WcHeyPTdysDuRfNCoe9vHy7nVAueFrXwA61eDhViTqE
kK66Nml+38KcLqEg1ySngDFzRvKsQYyQwKwIJDTbmn6MpGL70XcM5L3xlfhngW5T
j71VmNFfdEr9efmJcvjlsGV+yGaQDlys9sO9QlS39PBPohN7dH0ZHpTDyxSWrZOl
JXcKys6KCIg1OTY3WVUyt1sI5HCcHQ8uX7g35rJmQ9I4se4n5/+bkxq2OjCYZuxy
QPkaoGyV42+wWxrm0oKq3gtEDYivsazl/MYIRI2K9C6xrQa4n72a1QMXR/vJgH3R
F6gQ4KuHjNyh2dOtYiyQ64/6U4lUmf1T5uW/G1h+pneVJSC+XCAD7gLQ2u0a/Ffp
E4MnNK5LxkogSWWjcUn4jsCt1rGtFz723ugURzeW4UvmMXg3aQJ0bdqtYSg1mHz/
Qx35t73PDHeY3qWbghovWjojlq/ZAa0Z1d/67n5kOmKjK2066uuOJXCM6gERrKrd
AxkLFn8E49ObRJhpyxY+YK351pI8SQrfzNMUPFTbLaP0KATw4v5lFG6UE5cJCmpV
1zFmBhihWT9q1ssu7SVkYRvw+4SFgyD/9iwB96Z4dBpxUDwPa5hqeUVeucuM/NK2
o1j0ablIQNhfIoYlux44nU5Tw01L/DzPGbp2dsZgcx5CuQsraeq1tOYeNp3YlvA2
sZHI/y1aeRKV7T/fFoCTKHcaGo48S7Q4fSWeS82494WQLabjeVvy/eEq4o53tlf2
VJd3D61nEoIW+6So3uyBkNR9h/+FqaZd0reLssEgS+BLpPHqjO3nnp8j5/PgVcKg
+0suaWxUmaMXOcdXFQIh7IVwPSx9GPD+qoRREUHCkvN+Nz+X5RXemJMPD1xDMnAK
UO2/KWONE5xpDzz834EZ6GjaRCNu+jFPp6LEC4XzG854W38s0c/mqfX4o0dcS0rw
Iz9VsEC13QqaGNgHdJ8BnhzobcbteG0k0ivTWnlqfpSPMitn7RlWz5oULDl8Z/3e
IkbfERR0bnhKythZSsvoo7AI9cBj+ioEqaVWtroQoYqZbb+n3GdGojue6oPtbfUM
H2gyNN6gUcKCmUGimEK67i7zmU+jgwdnHGPVNq31OoXesG97UW2AbUrMJHZw3w/u
x4XQA5OCI7SrRPy6TN8L3AqjV9PlEmfwAcku3Be/rP47qXBiKGbzo4DkgQkiyRdA
cND9is5Pb+r44StP7vZfcV+P+Y9PSgFvH6zbDosLHF3u+SHwxaZ4y2pBlrHCsmg2
YHOG2imLOKGlRNcr7xmqlrsAaHxWyqYYagg/ZyCmV3MDGhnMHai6Z3oxWbi1tEjt
ZyAUKEAdt5WS/Bo1RNLP4Db14cnyDk/Hi/37VH21jQ1WgTJPkd1KPgzWU1I3yTzg
85ry1CWZFmXexL4uNzQbD8W651PodgWlI2rhft/YIAG+ATzV3+G86vU7YmZArfZ2
DzbdCOUHy2t2KKy9xz+O5vjB/73GRZKL7Lrk1468j6BK8WaU56zegYq/ckPHUPIa
Lr5Je1xmkZA+pi1Jp8SOOM7V6W9eHh0LMrk2nPMQYSlzGn6tNxxXGCN0oS5D0KeM
jz7JatKjkSYF/ga6hlwX/m+9mmD0jxppO+kg12f6hLVqoJbEnoORzfnhf7hMF0Ha
S1YDS6SJdTfjZ2H2T7EUfXOg6cvozuEW71PYq7EPycmqjAhL/fHUl2YuEd2K1Uin
aDPSRrW3pW85WZrZXvwLQMhkflsRrTDt+PWjYf+TKLOzybPUTMTqqkloWT9sm/Yg
GwidJNyDmMu9IDyttrnApJsDnz7+2KTnxX02iYPZzIxCWF/bVMWbEIZBZPCby1Ai
oHhPmFbA7Nunw5YDxPU3jAo75OjZZJLpLYSZQSUP44OGqLZ+CtPT2+ZQ1G1BZRMl
jELM/L+JyoMGjo2T8u1I1i+Z1cZCS2HCVRoCnmIabnp6laK6Dkj2tNHYmlxsx+go
vl37zQKxngCudJn5xRoiLWRh/drR5TtujHP62g8Vq7/btYnhDBtqdN1R9Aiy8qS8
fFwObFJQ+Mjy2q++pFFlSt9C8e5ASI5xNNVBxyxFNbAn/UfWSLvk8tNHgDtNn3u3
cXkxl+/uGaxHXoad8VcAQBctW6lVNbAu26ztUjE7OOOg5tcUFp9ZD8FUUt/0SxTp
vQ6OlXX3vZQ3KD4lcqvY8TVc128R6dCTFIAjsdbCiM5ubg6c68GaOWKjwhAP9akK
BcRD2MunARW1dvcAGGjXc11oA0zodJKNubxwym8Q+cdzaTz80KE21taI0dz/iCmV
MMOk0WT4/OvM0+4LSvfluMxecf2JvXdjIzO52rmsnEqV3LX0giHgt2pDqzJahcDn
ZlNcNbgHyIJerx9wZHtr8FEoKCCBLXGCnarnLh/rgIsOZFOZFdWkithN3ZCucO9G
TRNgkAFu1IVBT8GNpUBhjDXGpXlz9ExEF5Tr6KmdHQTI5muUdTQVa9+Jg0w7nSBX
4rs2j+REqwRyNjya5/DNo+VZ5CL5R91s4QjnYh2pbgnJbj7ekFxOB4QSgEYpyhL6
Ey6v1zZ861afOVYRUjPY8yzkJHRyLXTPbPPGIfTNTcgJ7Mn+5c4M9CiWv9/GmOwl
o3B5IEFbKFoVUuMWvhw9PGrBQYi44Vig5aEo87qtNT5JpNlGV7FARXftqnVaJJ3H
UN7U3QNtA9aC1JMb9znds7N07TF5VlOxhNHrbLeyAHHJwrBa+bnlMjwflhV7v9iJ
NnwGOivkjiux02X9ogFUORa9Sa2wFRO++3YNYbkqrFA5onvLh1Fdvfjz3HTpRL1p
ITrFqwQZidBy+IFm9NaGeII4Z86qgPoI0RY131Q4jg30U6FUbgUNaX01h4Z6ddRL
q6lJzCrYZDhkMGzgjwHMrjdPSpHxBku2+js8HDe5m4XKMM1L3A48j0PV/hhOFXvw
I0o3n4CfBMKkmmgWEGRNVCvxo466fKxw4SVbr3Z710iRJb6WHoebW46eohhJSumk
yJlU+suYrLuotCfGOXRwWz91exn1mwpg/Uh3cPfeZ2rQxdOwKImYUNs2xOkPKwPU
AWNWVxOUJ+6Itujej5O+hXh1UndbWK+umEROUDM1XjMh/Xzi5xTLcP+VaFDw4xy/
+SO+5A/UIPi/pvxtQhp7eKsi7dCNXQBxWD5eO9sjZRcVsoqCuFYA+VOZ1NmuOQ23
KgHObR0PuU0qbvTy4Cfe9IWVCsEZgX4UAcnArbMm55PDNMVgrO/mWW2Ca2uJOdA9
v3vR7oPjNrYJJxC8t5zS6OUDpSpEajXwuv3D6UrZlx/uukEgPsNvj8bYcOTAssSm
PTe0dzz5phi6o8+3+gMSWSpW4jlTKQvckMBTK0fMBw0YM/N4CJvmC6JzmAS4GsN0
kt90t2qUbomPRZ6tiZixAogxDk6j81XYpNMmxP/HhTxnAtwBMkbBje4tj/O0y1ia
tvWAwFWGM9Nfr1lPtRPSxVGenRh+lGdXd61Scyv8wJbyeweLH8vN3cenf3kHS3dt
Fhr4bPYRrwi9DQa1o5D74vNCZTezBeb1nLPqZazvjMIFf3kKEMksUINhyOVLelTg
WoUhAADI3i3YCLzM1eRUlWFFseqUH9ifne9BZqo02NPbxj7hfZyCmrhSAmWjMZtH
unR6fVuzqtShVbGJ5YBuRyRk4Xdfjlrs4YhoqCwRD87fGtPh03OS78yZgI25ooW0
e9niXS/jz6IM3gi6YNZ+coEJjWmwJBT4pMOZuPd371R4Nql8WtxgAqULb2MCZ4ok
KyP+yvmKXwq+UTLDtsyTsH8xJPLGPfxbq7tJ7SFohVfrD1fiQfXtMkjxLjBwUOF4
HNJJR2cUjXSwda4myOsUjZQs/3qOZByNQvwZznK64eGhZilQnvNYfyWMnHyBAxFn
EzitYP3kpKtpWa5Ew+qBbxLHJ8CHnkEFuxojELyrgX/E82zsXwFH+yGaMwzk7uxe
gZcejpbcMv2t8XWq/7pODrLd21j6MEXMr/ODSzDYmwdl9T3jYarOWEK2mfhNjMun
CtPM92+05FCj7lluH7iHacb4Qfl6M07H9lsXoREWxT24qK04xUaCGBHM8OifenGt
yp+sp0zSppdEJIzfVLqZKc3odL2CmDdJOcF+3iQhd9+JE9EFcVZbVUD+vPHyuXMf
o+Glq2GM6axCiXi/40B8uP7k9uXTPW70lU5+ZraDW7BIcId06YItYNviPOf9G4aQ
sn4YOuvx8D40Jtc0BvD8w9eQ3/5+pa8XI4yTBo+M5KpgyC8A7jVnUgXfX/m4yHS0
rIeSIGbZCUF93Ql9hUUymRDkqWhOFE/FNb6ACw+OE2jXFzjJYa6Rrw68iB8QHNP1
8YDkzY8kp4twaQC3dc+ZNBJgInNoQ1EgdyxjqpEZNwOwGz5cQ7PjgYdXW3B0T54X
mAkBXG4mdX51YdN6nXZwg0NznuVHqIADnuxTYPZO90JhBi9V3z4JQdYgI7+J0stC
0W/OmmL7xv2FYLfTDOSEY0wFXjVUoog4KrzYW/PDyKz9yaqzUiw4i9xLgDf+sgoy
29BuytS5F+Bdj5mHIzfY9M3Mr2i+Gv2rE/wU3JmhKE/zebMBFkH/2V9cUazXb9ro
+uTlU0G5Gb8aAQY6jr8Ewo6u98zNc07tWv0IHGlCHL0c6sRC04671P4a6McPjkxu
olp6YGWhwmv9eRVKUrlWriB/NOtiKzKsYFCUK7KGzo5VQDJ6IgmAH99EjJTYLgrN
9H/efyQjL/+E26yanL8+9zgNp3YQTY8Rzr7m8B34mX5O3wTikRhP40C8ER8A3+LH
nktujFA0vv6GHtoVRnVMLcjR8pFO9P+kdBRGROWybulo5kjR/GKv+XywoNL7OnyX
kTbRy4xq5FnxyaXK4Wh2XPQprMJdeNzxIcFrR7evNWddS9S1G4xK+ujcg+67fsfC
r+Kl6Wxiw8cIz7M54LOHu0yn8Rh/owfofqO3KS5A9PVqcOgiJxxkYJxun12YaBW+
hHet6AFJK0Ea8G7RjGXB12dndFeNtyd5PqtD9YpAkp+FmO44iT+9dtufKsLPmjZ9
nPzpDTeKyZOw00FHA0EinWNeKMbMTsFrJkHUERRiUeNn6Qkq97ShinkgpV+SpFz/
61sZBjJZS7BKXEihxkIWukdL+sR16vkcaBPOD0SAElm/73sPWNeHromAMYTd8TTW
l2eV0CDqyGUMxNLfa72dt/dqtk1YpZuo4oPhSSXtVmhqBP9guK9b1cUuNnd0MHkB
qZSn2c44CYUeQNbzvyjMsOecxLTRdCfyRj9O/b3ECa1XCxyplgnvppN0EwuhR5t4
oY2MxjmOGqegCmef5Hsk7gmoB2HSLoJovxhay/P75LJg0v9w6sUDD2KtIPuYuNfk
HKDm9XnYfeIKrMhP8gyDFb+92ivQVJCeXL6z6v1eLBF1dSb8PJwAv5S6l+kIbiK9
sCPOD7CRRgFJgHvwwOOfdrWtqnW0uPdxx8TJonj53Tu9hZezWHWVsdick5q98AoF
ghZBvOBVGRuEsLq62gV32uAsynZcvN1WWDJCz3gsudca7BqWC7BAqWmKzYnRZFIt
8yZ11Lvp/le5+qSnRkAmBRuQivz4vAqdbcB8T0ByZOrQ4aIAW8VHJWphmeR7Xkw7
VJ5j9lv5HGXFyFD6xYCLVCmg3sdkYUNXR8CVJYmzEOYpMdEORmitUern2eZdok2Q
QonaYE6gwoHoDBec8zyxgENQVPn0VarVnHlqrVFdcCZ2Vzhlfy3y9v6T82IFZ/L3
yRWXXGdHPjP/T2aalQ/qrjQfaIj1Wwqzwl3BVqj9vr25U4Rp2Anm+CMMnRgvPE53
bHBKFFA2FrvAvTK/wO9zKSGhDVRRiTzNkBxGN5UrwdQNdfi1o8GmAYmhMxj2A1kJ
p0pJKlSJciBwTMH4peHJEW+aIc/LwfSWiUOSk4r1yWyk71V+11yDSgmcTe4ZmjlN
e2fL2SoAYaV5qNzQ8QsKNv4Jbsn8J16YpxFfpmyievWwYMMkrKyzTb4WFASSe76t
rcZXDPIn2vaycn17lWav2RYTK0MMdwe1hy9n+ZVaIk4OKEoqvdytviTseUbxPcQJ
mTjtnvuOMpIRfD8cSzISkVH8yKw+bzzRjd4h2La/Ufxuxrmug02Pvc2X5HS1gtoT
f6FGh/w7HBUxWaN3Qd52qRo9yJpBWqyUU83B5bh7g2ZqYgvfm65xk3Dx4uR0BHVz
lb9OP4ZLz6MEki5eVKdJXIMzIA9hMkGcZHj6zwDvEOnms2FhHqYolVQNdChvfNKK
taht9YIQ3Zka16jV2m6XKoHi3SXXdntfxwTcBS8QdiLwm82JFP1zkv7JQYKFIctI
m9XlLPVTOZV4I05YkSosLMwS+1BNvNaDsgUjW1CUkJXrUfBILbi3AiztTMDkuyPb
VY27fGnrBkW278Hl8Ag8l7olprPEJdUdahPFlv6HmG5NMgS+Eh3SH13byLFuYfjQ
7/j4CcpwNBEDe+qXjm/3V6eSv0f9Ua3XsbLtvs1lJwqmkWsYi8auOwFGf2pZJEXZ
mFBfzw3JKmiBsBPlO1HKrMW4ZC84SKv0sYwlaWieXQ+0umf/q9ZTpNDAyHZe2bsY
+f4Ar9QfWNyOJuPZoRa5JNw9bl6YE9bgsBFZwKwKzSmZulIz5tM+O5ehTjo0k+VG
Tc0I3sXro9HgCw9ig6yigz3rqmeqDwZq7pBZ1yLCPWXV9w/uP6Q2ZC7budYDVbSg
vUt3cd7/ePZViXc84iYgcaZ7kn1VPUQVW0YpjAHyS1TJVieUisBb3llm30k0n1EV
w5TYvyDyBbVlTkw0yh5RycqJkLJWlFo8CHQuFjlBu3oV15mQD4kQ08qMfbXt1WC5
oZgZsRyQ/WPVEeAvvS3q2+F0zR8lr2BYgromDRUrJUy7DL9KzUtJ+mWhAjdwSknT
vKd358hM2HCDQRGpwY+onB6HlH4ElGLU1lkgGt0mbrV0euJE4dADP3CSIytZIU7k
lF66ISXnxisGsEysrp6tngPOV1YZLi0TGj2u0CnMdYNT0DDZb1/vZDz6IogByaVu
VxCThZYFiwj33UMbDHrQbS2DehamO6Jvyant0fwP4NKJ60IwS6NHRlPD77CeOVfc
IJranirxjsWpPPuHnJlDoDRLRxjv3x86vsroG0CyEWcS2uEMgJy/NV1SL3kquNbg
6DlQCKan6Wq+r6hbGvY3qsJyxO6r+cKXYFHQfK/FPMnDcAj4BCApdDsAKlacyOHF
mnBiA0Z/cBbHmLjXvBa5XdOkg6skdQWg/HmoAwGmZPS/6Vz2+3gWOazrGYDY5v/D
AO22A6vNjXkQ0FoV6qfFih7soywp4Kw+Zf6lzcF8Gyna1q09HG2hUratRKcTx5oH
M/ubedPZtuL1QRReonJx5RVMIGWs6zhM/NCtg+KVsJETWFP+PgQHhJLsMYAgEGzp
iihsCo5VIN3iIxLq8eAT8qJ/F8jrYVTEtyZLOISkSNHIkw4UmbfSjcaRoWZnQruG
S3NZyviEW31UWcOOuA7LRRkFzAZZB8iZ/0en4n2dUpnxxob2OYjPl6Nlq1Pt9U5Y
sJ7AuD4l/tr1vrs5KSV59ersYT+STLLI1WOFvnj5rhhTF1dTutCs/ng/elYneDrt
/gFeJYBsM969fJOJE3o84EA4dfgSY1J8CvGyTUvtwIo3ZavONhtraZAo49RQUOFD
zlr31eS6K8PS2dOzmdRb9YEMe2dCAHUSUEj9jjFwzUyJlA6qCCvXUlZWt65fCbgK
toSZHC49d0K5qCgBjdJ0G8x4/iyvXlJvK1Hw8z9TPf2bOMlHVsDNFbfEmV+MIo67
HxXBbJiZbFPCoI8Y6W+XtR+2WuZC7ezbPw36wKdN3+ahDDOc1487He/7Sei5kMLD
+XC/fKRNVVBAIJTpPaowuCTf2I1jcrHa8kzxo43ngYximSCBn+anU7bRkMSDFF0b
mlMROKAQpIlb431y9Pf6YqyoLML9BX/4Gcylo062QTwmDfCZhs6oFF0J4YIdjtbp
kUhKNVMgyTCmI9V5O91aYbYe4ppo23JrHrj7Ybnebpky4JF8+qbS6/JgcEXfSHzX
QtjdEGl18NO3kmp6u5LrYa2aoma6XJYvS/uj+e+7VsrL95kZ7gQZbP6j3wBQho/m
LCgT7709s5I9iJyTnIcYswbdutbjl6X51UmPwwlHu4zLNCxrquDD4Nwq2QqFBcfx
xAym1FWuGlYbACWrVEirfEIFJfb2cOyrl3MNHHLA88rl1CryPMp3NE8xUnDue2ZE
hGt1tnl4YmgyCyrAWFUZT7sySYc1jFyB41OghzEGe3mKPL5j7pBpS510uLzDozAh
vhk9qDqKJ2enlUdq0I/RJ1lxmdX81W3OGVRZ9MmNE4kgqHrJNglodizXz8vWnzYG
wDHpNlKI8uWR0/Fjzz5f4fNzciyNvMVNI6pe2WYRYQJyBWFM0mZikO6+h71GIRVV
5ZwcBlFtvemM2NShdBLYEizZREPZ+RcDNesseErmwnpjx0M1weubFraB/BLmOHNP
NOHT34hP8A0SNZhcKrFOsEIduQCGlCcTaLCGREDVhLK7KOR9jxLy3KvBymcKfYXp
OPJHe+C4ryRqIZL9ap2JsImzMPZzMP2wFUaMz1vx1y+WEFnX9ukpVkS9XoaGjtNy
cbZ/iM3jPfI/Yxz4cj1hlUE8eIth9TlXkTwCp/jP4fYlGdG47qMPX2CUc7rZTK6/
24Ke1GZKw8C5VKhNBpX7gTyevdDlpHXvyvDPtmLQHq43QA2vBvSnnj7gBavld4Aj
X3sFmIwbNCdyrHBTZMsBPFIhtd5MM+774VZbarUQdwqrI0YKFynZDbIPj233RDtf
h2FEWzzgXdicayAaqsmILT0ldXLGe6hV1t2kJlKDV0C1bwU4c7RucS3sbgjTkYyt
VRFVjGOb32Kutq7Yl++KTtFdRaqmd4A2IzWfBKHLtIlMqCCF4N/87c39crTuXGRR
fGBhCFx1NtMTjlaewOI354nHz7eLfZOvBRZn/ipZMQIM/jdz27/Sx+e89cS+eD5M
cdpEtJq6JOhAN1x8lrZRSkaCsQ9/7NNgb4eq0s1MQOso5YHXTJz/ulMJVEq2CUyB
A3piMW0gLVQOnoXuMlYBZ1AVt7u0Y+/NPeqpoVDVHi7+5oPrE/JwfOGo21AXT6lZ
DMyRdvLXTPfclyVUoJv1eWVcpYc8umi1fNrZ3+U4bOirsjPb/GJXf73xSaQYEsu0
Hxs64PYKLkVEp6WVbkVzjDi8xDJM3SoxoTj0Wx4/XjrOx58wL2kKF8DcW/TQB6r3
padyJxNQCw3pB9DPe5npEyKQkUiAunK/qF1tR7KVi/XUR1XVL13zS7BHTzvuR1M8
SvNz4UsMOHZdqvZSsXAXOiKx3X3nB/8sMcOJo3T5lB42FUZwvDFK+yMLRaf80bNK
YeYkTRDpkjgyAk/5xCS7rhJnOS11VXOW0ghuG6NoY1QIXyN0ncwbo5O5lHIvMqxx
T5d2EvblmhL70sl3GssxcHFDkVFrZ3HIYnV0LHiZFa7A5+nPCXeEEgISY3iQFX11
gOpGd9QjMgLMTl+euLdI9HoE21HwvMfAkrmsquZXmxoUlNWEwNbMaYNdh14a4Anm
ann8ArwgFwF3B9hJCasGKfZwo1zliiV0ewGmiDBwODP1CLk5/VbZAEdFRocyuXRQ
axIsW5zVtN3KDQa2dkmND1gZJGT22jgoXSMejTpy2nNk+IdEraH2A7Y0bo0i/Trh
AiDLebk94uYfNGYXQX953c72GJwqzRuLLtKq0CRAdCZEj3TCJOhx+Nlch6C9Cuug
ecF+CsEPiueYMeQ84hoHKm3n2W7qow79USrIYLL8Pno74P8UkfPnxsSPQV5qO27Q
x5+l5oOq7P2Kx2PXvP0b3wOIrNLjE7FSA9hGqT1STg12PcV4iWjLy9w6IodkIxOV
JAZ8yWKYp6fbvmfgzs5ocavabPfANYb1VAvG01U7QVhFPPPAMLIAlJipDleiEIwA
GIGsqPykDsO8jXfxPJbu2URqbw5T72afMOH9rtYk/LHrDwcekRGxO++soHKrpmVg
wPOJXAi+XmODmv4Dy74/XpXSPctgGeDdKv9oIuDenqqtOcVKbKW0ywAIO/Hf52f0
WrsStTmew+pjd1MM9U9w2sKibwgMhwqR9N2qz6bdj2IbSFj0j93HuSKJmgP5TknW
q+SJAUjlC/gRKtj4n6Pr8CRUOTZM/wyeGfMNv+198RLVnB0SD99Ru1K5zfHGYAq/
mfGfQ6wOf9Ydtzg4IiT8jOkAantdjlsp0gAllNwkFkV62eBdZHCnz5J9ZRiSOlTb
pQIYYZtFELQnYHBiktzuKjcgO0Ch8xR6eWqe14OabaJujmvMV+dPA5iYhjhhsuQi
VmtPxHGuqgsMxxDh3jwpY5/draKHSPfWKgc1zU0VxkAGk0xecN5CvkB4jB/oKiwC
IOre3SY7rjOlf2uKg5OrNc3T0ADbOzufrT1DLqnpo3kqPZXlusVQlZZuHKfR2WDG
7VHmGLQ+E/xXV7Vm/R5BXeYb3kXfz4Kuf5tjJlSgWM/YnU5PLlW82tuYwHMWRKqy
GPBNGNENmP0hWXBsPRQXHAuLPicIGVBeCYv5dHtXQJT5lvZMpqkRmRkGUQ+zwBuz
iNDlcpYCsX4UJwLPf6ghcF3+IQ8jqXfRX+Y8McVUS8b9zAFrFWjmQwf3mxqQhUZD
yx6L64q5T8RLgIb9amgCG38wx+O14Uy6ujx2ceb3FjImxgUVKtqrE/DYzn94IwTk
xvOf5seHU1b0RQsaT4nE8b07nEu0zEXkSNmH5bX/v1IYe6m5yfiCLU8vUltf2Oxc
iL6csO+itGDUBOywJBmhTzrg+wqe4FNzQJLDGGUK7hO9xnDdJV6Mj6eFbjfZOZLA
fxgUMUAI6YmjzCPLdHK5eQQ+AgCu3qk8Z1a9RFDVMxWLQ1HLXFfIvEInYeeBOppe
cc7Scy66PKpwgJt/h8xMW/O4l8csZbCUJZEWcNK4TlZL/j3R2zBB+6e1zTDos70i
C8bujpg5LDdX38VYYuI7hMupZkBe+Gym2WnA13kIKjg0NNupIv9EXdWg2Q6p/COh
+KxAmb2e7lzzs9Kd2phQl9kIH3I3+HsoVsmXNa35Xi+pNituauYNd24bqMBhNr7M
4LRc5/GmEvN8/MltaLhLpoX6bLLus0/5MIqC9i5Cz9q7AKzgK/dZXx9E0PDKhJWa
b56A0DKglluKpKIcy1dGk0QDvfA0jg4P3NGG5ZcovJpr49cqOWBxUSOAWmFHPH14
gZSH2t1HNnTpU4Cb6eYMMjdow+7ioBt4fQAZS8Wz9hcFA/tlz9UzXiG79ol+fNLs
QeP+Nevw6mjGSUaLkYnmUZVMu6k8wSWCHzTg4BSkZFFTfFOVDP6jeWV41KWit3nQ
1BBlDUdoc27M0aTRtGKn1uW4qW74shf88vk6TQvF5CX6V843kEbnI8+YFHwEKgr0
R8zTzWVMH+fjSvROKEf3nAtIEDRkWY+AHIGpoyhLd0QMCzDlh7q+O3l7kDVyI+hP
/+HF9DUelNJxPCvWLLD8uU6ikPvkN8T3V2IRafz28RmzJw6j8QhnM8tvn6gYhuIy
t27945zoksnZTsR5k1wnfodXkeVYL82UMuIGlN0yAccM8mYJzHto3zNW1um2lZWr
NeuZZ373C4jA5z0PKAGSA+7S/YVu2BUQur+UIHvD4BY7KzhF8DppllANpRu27fKa
pQDwJX8MJX3dJl/J2Gjb8XtBw+MHCufRCUzMwQ8NVeFU2NR+C6Bp3qBlC7kNMxNz
CKwtn9XIJDbWRnKez0fF15A+dPkpW3RXR84VgVuUEPYg+1AqxTBK/9pWj/FYWlsr
FFWsGZtvle2rrfEWFOkJNCES2PVEgiWB0V3QslPoXjyNTXiyrqs8u82r8N0NBDJJ
OsCi0OR871ST38eDXqo68cEIMw3FZeX+x6uVOrIPmaasHTDJWv3TgeISiq1ky5X3
d7vA8gsABsx3ZcWFGIlS+xl7rPhXejk0jidWKBjvIrh3WNnpp8+Ed+T/Zs8y3g+7
jO42mSptikCqgFlUV5OheaoZircldU4OrPYbe3keD8T3R3R9qxoBnYN2acH+9NjI
QkdDtRATpxd6CEHudsHb6/9rQAxzMCkH4JO0k+2Y0yy8/+QZulP7T4SI24KIZ4g8
3zUyMxyICWv6LgSPuZSE2GNbxJZYh6WQ/4PhUgOL6uEUOo3PLHMgzqGgA+S3Zcrz
DsnQnn8hiH+PpENKdEn6mULCo4cRrexwUs1azAmXT0Pys2ZklZMvExxYBA25yFOk
OawUO+o38+5sVoZ7qZ9VV20p7CURQCIoV3XMUjeVfg9BszI1GD5XKNEvYOaK7L/E
7YVjuUCdk6l5Tz3sKt2vclSp429q6yP9fNYsIp2BshJTSr1yHZ8j0b+iaGH2cKsO
ckv8caNOFdXRMVoqxHIx/e/NGFuqIDY0SrsOymNYJLJ3WxzudTWq1eDbsJALUVhv
+CnKy3FwqZk1l/dfhPjvhH6fVQZp4TmA2eTCbw9B7eZ176B8iVcep36ljY9msPuT
wWI1rr253zJNtEn0GK6I6h2mCFR205Ny4KI4MGUu8Le/R6/WApbEkUkUOtimw7NE
EN71EX2dAh+yOmoqz1eSpakPDmZYE+uCUngzAmf7laY4O+8q+UG0dvRr2s1rndi1
KoPq71oBUGDyClPoEtIxsqx6eVjKTE1m1rsJsniuxp9qS4YgtBwWlL73TW9UQGEf
Mhm0auN4Z30KBQ/GYd42O3POr3zr+5uI0xXGGS/XOvVxNitzMhI/5GiaNs7xD9Xz
+NbnWKcVttJNot764xYZHNyDDRBhzNQxWJ6ejpxbNfjBKrC6fwIyGkEsZWUTa/eh
Y4NGvzbfv0RMw2iTLjIg2F1Wafh+jD5JgwLmafaSqq872KEPJ+32iL8Znrx3mSso
2d6GbLduJ/kQF0Ky7V9iRDsENbU0MopaglaA1ZFq274BV321offO5Q0Tr/liDaod
a/MXm9QGFe+CmRXDOybHxqQmXI9Sy16Uoxir1aCX+yCMOtLhInvdNwURoIj/KyYP
6CGx0+z6ic1bL4Ljq1xMXti4BHQN+KQU47MpRNj7RISb11VbizPX8ZrcBQfKIqIT
vXOC3G84Eer7CoAEQl0HhWk7cekApOe9DSM+htVxT5HtBkDtzEqOiAW1Mw4tGtyZ
/jrtp/ect7KZLSmFpgBUoMn1SfBlMTno2Q8+wIn04gEcN4yDy0eTD/L0wSX8XrU2
mJxGVpDL6rgG0w6jXMVkGS88v3uCcabaVtp0Zct7qO5bmqhM2unf+83RXfQHRayU
H9B2a4TIA2GwYXVXCe2UVNUJkql87PUxiHULtgyyCKLWR1Fno7Wf9P2iBjxYh7O2
u7syVBi+g9Vrj3EB3yof3l868cTojJsUyhRfJ0CE+He/3FkINLkOSjXJgGs/e/Rm
0VyERHve/aNJSzgVbV3fz64Lm9Af9QxO5LSI2H3HatV9wHkQG+EVC4W8mZ2zASq6
t6R/GaOyVMtY3ENjJ05r3550e4wxrhF2XwafaK/2egHqfis5MvQcyaJbu4W+IubC
KX/Bsycz8x8rMJBxtNWc/X7rPrgFTFlFDKtkkgosP+PMlXipd0frfDYWCaccrVWY
JEapc3dKcJAhLQR8LS+qPdTY9CTbSzWDRF/Fpvip3+pgjDF7pb/+d0KtG73TLHOV
Nk/QyZho7+LaeAAayuvm3T6QhQQLufEJmSVz3OoiVO7DKOLj6mh0+YjR4cwaWuH3
LgIm8u8qVY6ekFHxeMC53r8J3755TxWrdHJCyYxcOc/RJzxLdCXEDWaXdWCDWC+m
INvtW1p9sL43h1PhTlHK2zDDB2PbQ6x/Ff6dWOv5loQWUaWPzi2m6MZsbd5M6CbD
LcHdoKAFPUkMlefn2eH6XrEcIIHg2h8qQsY0tWdfeRJsQtGR+HbveKXR98LVpQiV
GDdBxLubedwKFGgw711qxx6ZwqdnlM+Ew2hvyXbLP4Fbm96M/Oyzx/FR9k43ooHA
ZqscCohBd7OfOcKPTaKBM6HR+TcA6RQF0NFGtXunt4veEhur/WT8H/TEY71lrfwN
rpfkKcX8Rp4ERZRH/PJGpZ3jeky0VPtyVceUoXxYRDwus3pJD6/JglL3dOU3CIRw
wWHsr3irtBbD7Nl10EufckKogRZXTCxUpoIKNmV9YgJlrEEwwpZ+xH8OkAaF9RQo
047OZkfdeqfQzeg8lip8MO1rI35PmkeWqDgn+q6oH+Ref49GRFyDOVa9u+TPDlVK
ltmzqyrBs573l97ULpRufP/kdL2LauIOdwVBTohWNO6SSXz45t0l+MgUpRcqacnR
SKGpvKv5kRYo/FDGWd856SlIm84VuF9lKygh6aRvAqDs7qsBMC8MgMPj8T+MDzDd
i55TXorRo+TyGoXLrgeIO+J33VH62qAShNMl+i1P8gbYFa+p+if41fY2JlStBrwR
krOmR0SIwpjeVji/Iin9H4E352cEu38CKujFkCjZsEovkjYc3hMiV7lfU3IijaOf
2OFhrJPb1Ke5Bea5jZb3gqBC7GwdpkwDEVMzyl1cf14D8QYuQ3RreeNgNGzWg0rz
l2p/H+UwJ3tYLSEIckke67MWy6U3d5tVOZ4ZXKGWTPdc5mqYIxS0ZmFeJzCGdLmP
8uPK+bD98aSv62sphZHLpgwDk1QTjdr8KYDFKHMXivDIPRsAhuYYQNVS02nVtKPx
jqFnpFp4vefkBqKdd1WBpnVoSE2r9k723XaN/4y8o7zv4428qVa76L1o127mriKs
y0sSLe2UCThxpHjPPKlzywntLF5LpYxgAa4ZJNJv581iHvpcUHnqGKru5IH+4Bfg
3DMgQIfgONNrnrMjuFMdUxLBC+AWL95vE+qta9VbXH6cOdjiJrQwjHWgvGivqSoz
vWBmOOGaPporiupaG5Q77rQuOnPm09tf4N22VO1PwaMbYG6Ix4NO6A5wPWuC8K4P
XJ4aZuW7MO0GL3ITX3ZbteZIDnkjbXlpG5WHG2vNSZrMtiOiuAb0PWRrA07IlU5n
BYn78SWXd5kL2YZ+ROf2dEI0aMt5a6Uj84l3Guc+vYchuJetMpAbu+H30+DNLxNh
lz1whyUphp2ZsUtrqg7COCBxi01gv5DDqCtc/KL8+odyXVlpt+APba5L7l2oUYvJ
jDpd7cFlGf4aMX+UYVHPtJHnEvBgs8yUHZQLMLIC7d4zSJDmMZ/jv81YpNBdkUYs
fvq7fcWu5yPf3F9JkbrkZGHqm2IuCIQs48kNJYXIC2Mu9ZPnJy4GDxay3L036YVY
TQNWAwIChotrGvKRnvjuRcmZ8BgaYaxXnxLEdeWRgeowhwD/JMVOdQG2w7OiMnyd
l/lBnkn2GZx8ScS4a7zcCPhUY2oJkxeP7Zo/VoliNhv9yGv1wfL/YeebR63ZxV25
ieQdQBCipnLviTUaJBhAteRRELZzxv4JQ3asTXG8QBMi2JigoRAGSgv5tG0zmyPg
edBmvuWSv9FXigVsVTk/LRFJKClQMhnCME475sPO7yqD7bYsvDJZLzCkB8XZC6ia
9lSGm94uKmDGOEkhGLFtb2I2rnrdhusCRc5c3zz07VfGkQIYN9WQa8TxhmZfWREg
uGHQDE2kzlfaDK9+6Ot0UnNgkIaBl18ZVqqIF+bch0XkGL5/+jXmNoGNgMQvk4Qy
vQqalYLKEGg62ElwYG4UCs3TjwIECVFaUlrxuDIiDkFTdc17LPv4CdkxfW5yJZZN
RDwhZFas2TRVnyJu2TRO6VCe6tGBSVBQ2oiuJzxMUNV1PlfplicdaczXQDtMrWQ7
XEIvEC4pT4DmRVoaDCW/A0VAQTSeEficIwNc78UZBU5bvsmh+U4yL61xHr5m7lYE
LIp/fziC6x0OmqZzX8uzf0Gf9c+r1TDHJTiU29pDFE9u6e8a48lKenVFaBWr3goy
Bibe/McHN6XJPnAAuoXGmqO+ouV2QvdjVRpGBw1HD0UnloN+nQkgbUyeMWrNqDrE
MpxwFQAqSBs7jODoD4RdBaSf64tPavPTntXq6HKS6BfFNuGREvI/lVqqJ2qqVjfH
2/YjAugGpucrLQoWEzs9ifASs9Sr6dT/KRiS75iNXDif394rUqg2ebcdRXWTWYVq
pM/Ed3ChN31be/CFenB1Cd7FcIMao4ZAVhfceAiiQmcCnjVw4gQb6JRu85UJrST5
FqwDVeIuMSrB9q0znewtJikec4jrNY8MGzPrwSfq6G8VyfCgXo/tPXnXHlp307yx
AIFldZvfqm4utikFGldw4G+zb61ExoiIO/HUtiFNxRSxQEziBS3oCDCF6pj442MW
cpRzp+vnejHfwB28nZvShwuVtJ1ycqmtYe1/zwlk/c5UZgVHWH3GyMAuNvFlIkPh
R0h2lMZXfbyQT2rKHL1XIEKoGBD+qOGyQur4FjNQSl5xqi5hmErVbxavvISXomRI
z24tC52bXikF2fACmpm4sRTpZ3THHiaMoDzNhQxFq8ku2a9MHQBfsO74fTYw798g
fYaz9xeiRhZrzjQQgjm8E9KKgEhY2l6zaKjlZIztpcJXUxqstVmj6JpUO6oaEU4z
41pfFWmvmQR1hPayrwUBguI3yJKVLlpgtPPuaEcqTvU3x3PxYl2W8n+eBt3GfqTZ
k2CRKw5ECJE+NszY4PDwRxD+yk4bPiFlASQvydq3JkDKjGYy3G4rGyM9zeA+FA3e
XSs48ISK+V93e4U2Was1J013Nb8p7rHc9KTDNXY3AxPuz1EPdLdpb9CWsfDZe+QS
Z6cSAzoSmF/Z5hUB9BEBYryjQMzRKBIRpZAjHt9P+PuHP94LR5x3r8Pb0wagOEyn
vexWkb1OXtef9q3+4K0RUs4Q6gP/991kjugSQsKKWvpbQryTCyKHJhSeA0v54/6v
fMvzyhC8vyKI0pQiKoPsKs5x/6oRyKa52irTq6kSGGZPrD35Q//xrUzWm3A0CkMO
0cu/L0hENXHykNNqmRfDjHt9QKiYku/FScyyM1e+4in89ZhO3g/KLhYo250VoTB8
vibStrgSnTKc9cxpQzRbhCJuycL2e+/qM/6WwOh8gabKSquVAFnQwvPN6Tm4acEj
HgV4bBD51oBbWt07sgnM3tYoTniXn5GJ1bPo3FQ6BJdkpy456oIuN5PqVOAqfReZ
1GNEu0quRtBYWaxiQr7k2fTV2UpDG1MTvN5XANAVyEtdR72gVQvENcxnSI4Jzo/+
Bhe8nvKK4acuOLYtJ7hPdmGhet3J4NN9f8IH5suXkXS//9ZHZiQUqkNOGyPkM7kI
btsE5IHFyion4HIa2kpJfSNlrjOu4TXNvP3Ptr6JTtX6GHaKlqT4jiZ+UcCOPP7t
8iTxoNXZ9OZ4lvh6uxvLlvQfjm2LcqnO3Xq5ycTJSeUfjyO1kF/38FMmEBBDT1Nj
cEwbgkNcHG2W3rtxGdZKJKG0b4tDawhaKzS7WilkddpZgEZz0pxrRfXr2FB53tBO
kcpyhYX7h8rTqEadMNGIdFsbWCMDZ5PffCaYInNunl1lkyBZXSm/NCy9kXTBU2at
0EFdtVFrrhak9zLeFPJZ6gboWViPwe9MuJ3sTPdhbW9EVPKdFNWnsHXbbSVwHRSD
/YbSUCMAiIYjrc824QBmvfhWF2kewPEqVcjkEEUhr9KZ19l+n8y8lTVdmZMXmQqO
3fAUxGXeUgq9Pvj16xMswmW1bYahOiyu+qghwrc9uypLVH+R7PEgEzgzlDW7VW80
NzFDSgU7zM3jnMsplKACp6JpxMxVo4/Z+Q4WzSrbYuuAEfzV4QZumMYMd0FxOeb2
NHjgQfcOEX7zbPqte3fokcUdnOIaRk2immGZl0DyQqqlQNrF2kjU6fC6oubJeSKm
xXe529yzpv9BNCYiMcgimFULyADzGjeTy2lPkMmDD2vRUC1f57ESg17RJ+Uxe2hq
02Wj2woXJV1lzcE+xUW/lNq91MbBIoDSxQbMViujLjXJy1BqgROHxCkGHkUEK4O3
w7iR9qcrjPsrJNqt3bdTwZkdsHVv3A0EcvAC8pzsHKVqIck0gyhiLvbA3+o2a0jZ
sYbaI8GNcyQEltD3mQhr6h05S/pzpXhhcbBVqdEGOYN6nEb4VsQOdfbE5QIkj8Xn
Ts3eunrb80Ek0sj2kF8YWIGz/wdaaZ6mc0Izhh/Uz8zUqXMxkWw7Eww8yuxq+dfF
uygEWYBUfZE7GTTJezS3sZPcQZ8qI4ndD8lXWQ6NT0oUKqjcfJ7ntZQG1CM8oPVQ
SOLjf63MuLnJuRk5ImVTYaX/7mENTzE/zleijAVqFSRY3RaMRmKOFkNmJ/nzIsio
UfXwGSex8aFOk1fDE7JhKjgj4yIQ9eixehzZGYtlLm2Xq0lDiSjef33FRXY9dgaB
NyoX+htMT3RJ5CF9jCijE+lLf36efI64Edp43FskIc7NopzaRXIZvF+zMtpbzMqI
mJHl2fY6iq8QF64luIO6YCT5UiOuvtgDNQu1TEqEEZHhBigeZIpKa/PvXOBNCU1z
orc3+Z+PzM+QK7bgoRy//+ig8envE7GkBkjFUoGZF3Dc5XQRCZF/p7J9yw8b0iWE
HFmFLbbPuoUPGMjpLgxIlGxjrlZMO3AAGTlkEK9enHx6WylRv0Dt9RW08ulFQWjF
CSyeCqCN8GwgQLA6wkfHuheYKh2JG6fInUo4RlJpP2msfng5WCgwvNAy9a8gISCT
cgBMfiPb8O+fsgNiDktZyzm3xXFhnsDjViWfb3XEeUyGQqCKJCmgZQoRQ2I6XRji
9nS5qiJXcxo1a7zR7+kQSMzX5u16ZgfRZw0wWYPwJtGBNvnL8qHHI1Er8P+lZUYp
YlxTr87fHtKdXGDcVcahHQMgWDYKcGpSsy9N+mPtpEVZ4AADES356AD6kL81Xv16
JLMbOxgRfo+H66g/VFRjFWCFq+xjkZHRXsuwFpYrOjZMabQh1toXwIxBVkc7hckg
1UkAiYhbjJjS+Gxg2JO/FEj4RCovM+D/Tjbhpjsjp5M3KVebHWmC3hUkCzqO3Zyd
wkcb8Hba+KmQtti4KzsC/oMZLnwDRm+pv8wk4CGnAv3nMjzlcDkh1g7QggxKT3wj
gov3d+tKMXlkaeL4z5BGt8N3bphXdTk1S6eM2lFDD9zwt1jRKME8WyyOcTOP/Dtg
lvl6E9na+IbmwXHfU6J8HKkW7RcUiWR5GaxmUBk/2Z4PEx1byLPaXLjoTJxDsJox
VZHWJZWYbPbJhiOU5O+ymVFsDbPXiTEMRjUKVdtSgdY4mhkFBa/wt1GyqPrLUGc0
02SX4hFj4k60GaTBIm/E4VMFkeVvVGB7WD8rJLvQAb3rGS4a95QLyc8A6aiFPdv1
fxiHLtQDquj9T34Xu4ANPrq+OM7vGIZl9g7Yev4yN1aJauA2km50mkx4VH20wOUa
CjhksLb6CdNsWPU8VWUXmzQwS5OZH/SQl7gV2EcHeTeTVwHGOZvy2woX/HR/4k2X
7BUnn1TjLO6GOHKLggNZvEYksmIl+E4qSQQuhYfjBmowbkJdoEKuaDgXHTEhZq8k
nyvD6k2n4jTVoyF3cTLcMWc1t+oXu2qXwBDXrWpAPiZ8T/5SoBSvBMRLoaTxo80f
GMfGz7ZFBqzeRmIMieKVOvuYavoS8G472sdZhia+NZjNbrFATgRJokxvABLTql4z
7090SIfduRI8rdCUssXrP4eLE1we1D4lt8dnEAoh1NByybJQ2WfipIuV2cYjD64u
jK5eThBKSRXyBzINeShcbeSJMHM6kL56Ccnrlc9WRM80oaAljV2YKgSjMfj83inX
DApvIIbRGzriZaWrgR0EXpH1edycsdPMQPVJP26YfG9o3d86/W5SsduVhtP1pEXB
NQBtCKSeGmElqqWaUrVcBLi0kXz1Vsp6KQ/A3rlMUnuX6wac72aHoFwm9VmYl5n1
4XydHctHc9/Y5xQe0HpOeaTZ0v/83N9QoCxpAWF2kAD/1AT8wVczI2KRqUrvgWoX
9PzVHSnKn9Dgkz+vl6BaqDHmJcoSGeJERj6XnKuuDxczpBcVK+xWGR3zMTdM53LL
5gOKnVAS+oLOMMkU5c1H/+/c3rrn4Ty0S6Fda0UW9cWSST6xZNYKKefNH0aEeu7l
JSzdiDVIzo/UWG+FoVIYnu4ob1EmV7vDwMoLfjVd0VDkhQt2tVgHIwB2D/OR7I8Z
vOMLTtVZqEbPdLqHD3G4Vvxyz6DLA2G3EMZnFkfbx298sMG2nOWbAJ3dkONTZ0BT
/MxrpUjAPgdGKQFSyGKy1RTqM3d9FCXUl2IXblJ6mDcFCaxocYJ1PbDmFD9ia9Cb
UAbC+JltjuiiypNpHk7QtuAF98Rk91t4CeEBTtN3ttpp4npE49GYn2ebM7YwKGdG
AzMV6tPA64Mu7szI1D1GBw5Xn4JdoH8ZYtxIUaWPU7f5bZ2WnGt26vy9c3PV5bbz
QJtTDzf17vrqqEuBWDZuF0pKmniTCnwdQDwUEgSZKQPjg7e+cMGL1WI57blVNViV
fa87Hc4QcX+4jAZRR3L4v6lpuHqayae2Qzwqc/cpVlmo2xSZWaxF/1Cql3jiuCIr
RUesLb8GUrfF9LFhgHk+DjXTcEADyW4JiWxPv4Sqt2orJSlgYIB1iPEtG78xFF/9
HhRjpTlZ+AlLbD4wJfoiOrY82Yy4XUrv1azAhfTiucmp6ZrNzmtsfF1IZ3BpC9pD
qvfpzyASHwCRFenKvytzXhIBEe8ccjlEehkC/9W8BsBnkMYcPgcywUtlZeoWQYT+
BOLUm20lZZvz8Qc7VliLzmMM+AEBP2FAoSK2dvgNeqHCBXiC7hvRqTIZaHkx13tU
prz8z+v8i2VhdjTyfdGl9r7BktuepUXHJ724/WLnK8p6lM56AX/oyTWUybdxmDf4
w+ZfR7hG9iKAu4YSkGXMSyeqYfqzplTNG8EtTiZpFQ47rVvfy5TxRSQRz4jUmXUt
FHGzE/VJ7mXxF1GH4ZnpXzPKThAQm/fVUudDQ9pD9sobn7qsMk0rxZoh7mfRcmff
EsVw3n8kAtPSre6tWFHb/U7z4QdXQGZ6tKEL1uIdgJwHNC4Z/Qbp6D4FvMRgG4Pd
vSta1lq/Gkw6NSn5xNqaHlBN17HgZn8acpqNR6quNOpfrWFQ2HyRF720ZG9tRv5b
CVjUoG74tCJz3p506PJyw33oIgY+B6KC2FhQWit3L6unmcCHOeKhbky2uIDt5IP0
H1LOpXR4mA7pskhX2ekMwZa4bAPcUtu+xZfhw4HY/b86isias9qsLwEGqB13hiiE
2L2s0DHjjPZrIgL4p4gnZ3vQUmAtzSbBB+3uSoIDve8P/sS57vAngPECMKcWLI4x
nOfa9nTH6CNEVkBpg4jFCOrByshPnY9gxZJ78LXduk59ll12voihr7xsTqOEbgbr
bkGFfB0NMZEEyfAT1tgt8JYEd2ccmYxkjuuoFPylBS4twP1dhDBXEyL2+rJ4K82M
2ZoBwj33TEU/d92mSAyf1qVRTthW+9t2DOJQ0HxXeam/Zme1Kji53MA0dKIvM/6R
ql9vo8HSHBiopzHGrPYjW/tlgjsBBbeyABF3ulkwqtPZ0MmlxOSdHcOP1KRBUZxu
w4ADu6ew42HLFldP7eSHGPx9dDsIkHdA8mQdpkuWerZG7oBwom1upcw67xbfOfUW
JeymiEz3sjQIL0AHUWquR1v4A310VQ7J3eq2k3onQxWJiL0hb9iPW7j1Oq7nyua+
6O5vx6EAnErk8dBaYFhlJ4VrqGq/vXFtYMaqn/GNzN/GVawJvPZ2NY/6TEygM9wQ
osJ5rwW/y7YLa+TwpiKiaT32iQ4F5IJN5VwHVlYZz6foNd0uPJ9kBEJxemLStkPD
0K6wibW+NfU/OFPCfnjwC+nR27s3LzvVIbqfQz8V/QME72SmpTVtPiYTk9zPxTp7
81NMoqJTWI6UpV+N+0Bq1solL0DY+gqYjYn/ZRwarIZRM3g6VvCdrBRxwpLOORh0
Ff6D0k4m8DyynP1ubpBcckx0da0+EOiPCfjUm22uVKdJ+00I37HwE3j3YyUdTaAP
2LOmwAiR5xv94TrnphIaykwCxxreWCriMj1LtOYtWqw8IT3o383RfsZa5My9Cqty
yLD60ow6/qvSFUTiR7dlfVewjQQInf2eX3igx6SF+BlwrZyMLz9O/pRqRpk8s2tq
fPPssa47bPRbMwaaFn/j6/j1kPv817qjAS7KUfKbYogHnNQqCu3AlM66OTBfidjg
7i4t85KNBj2QwdJEY1V7MAWh70f3mtPk0sts97/4giyJ6Jzi2FAxtZJGeozGURMR
daqhxC+kkSaMuq2/NT4nM9mWA0Ay5SyTCD3S+nlpx14RUwsv0J+I7uTe3ttu0fwU
bdbBARi6kokYTOu5u4aOf7Gqi0P5pNfN/unar4zBlMXd1tiH8F/bUxPCOgMN2anp
maPsEcRE0Fzd5tafuFWwtmyh8SYOyd8wuagPmGNywoZJaWrzsIo5HtWBnqRwgh2q
YKjTnE/LPJ4pxopUAR2jkMLtrusTcAEgpQheY6wROg0smzR8p2Y/Pd7eltS74nVq
WONqtH5yfd5xYqIxIf6Cd1ldbpj7dFZGR3wYRhoRCTh/yJXVAAAKWSbpLTGOrrH/
7JyNEIqtvxOM/nDhSqmP93H8R4uT1jmCEM+5wVKX0/XZBk0HjeK1DhOotBUjTvgQ
tDtQiNBOoU9NvGiZkXinzBQCpRfVJSBMyGInMRJFGlrrCZE7ZKtEI5i700mtStAN
wfy74GFc4dEZbteQaceh0iuxdu7POrxq/U7ogvim/B3hV5C9DwAc0B6KjJTdFDVK
rRgZyrn3tsZ6SuNJF9Xu9XzOOV4+S2PiJAw6SoZLNuCWySWBP8xu/stKihaUhK5E
QeiNjR15sjD9jym8O1mg8xtX1BYXNMEg7J8KwGQzH7SJYt9PIIo5vrvxS9rrRv7s
2fLlgV2qhTxsMInNazTd5ZXf20CKpPBERUvhVAFBdV/MdqJpVSk8FA2qFhnmNFQG
U8qJ5x34oZRG2ekfCh9I7aDtLgeTgvruNQyXcqQlTcSH68td2T9W/PYhN8gheNdI
HbzZzX7FI7JvWVr94V6JLV4QbaKc6GoRv9DqZWgtD4XgBiFBdnqu3I3CyRFQrDRC
eQKCtc7KHo4HEU/4y13rb6xzFXx0D9/ygw4i9BIOTk2g2MUgNW0KkimgJhaiAKmu
kPj5oTX4RY6eouv89XXWhw0g87B+lQY37AD9G4Sqy3d5BCPYFbDXG1z7yFSJIawj
srxrhkTtjOWkmaVzxDZvAC2AneWgDhIoc/8P8VjB6kPlguoRzRWRFCuca5hElfaU
GmNo7y9eBYToI5SoNK7wIETxOB/JFe1IO9dw0UEYeZwlcmLKWmmXltW4aYLCIkU+
DEperN00XbjLHgnXiUScF8hXD7QfJtqaxh8Mr5UbMd134auvArXgrzPemovdjWfE
zKGplV3jFs4Zhqg8XRCtsJLDacZP1/kRSxllVQItAlDQzwMmjE1jx8ZEsEWimULG
hZxQcex6G4UYRYCGD68bn4ddlw+IvllxvWcqQCACZjRWjMYwluPEiZxx5ad7Epk4
ghiBjaQ5OTiEs3PaiquEsnAZgF+VIZnd9k5Xku4TB3M0wOs57trVKj2jIX+CIppy
AZw2pcm8mPtPnnI/f6In1YlYESbExdPXeI24ciR+VBS15U4ydQjDcipS24r1NM/t
1L/qQIVipgnHjb4PGpPESccsGL7yIfHNx/yWwxzSVw3WM8bLesNaylzBa3dcGtjF
qEje9kXrEcWCr9FZ5ri9f8m71sdzIqGakzzNkh/tiVPZxlQRrqgd3k2oOLRQ9kS4
OkQ74UyeKkmR0wW2qwwxGim9/eroDu2mG+qYi7xWamnwO2Ahw+U2Ov1Z+qFFRxxe
tw9V9LJz+dgBviRoS4YUxwRkekGOskDFyOX1l4epCcpGda0+KU418JyK+gc6DSfx
utp0cXnrmvCHvoIyRKTaxvHyHlw5Fs+ecYm0VdCL2CYRTKkVBkI6itqy58F3B0vm
ksSJvPa+v8sXDaH4clmovxhnn2itchSWMPwHffI5qG+QeqgEk6YbFoeQq64LsVDv
lK0Q2Z3gV0Q7y+ZZVKKz/ynMf22uVipQB7maBbJAqHTBlDuvlgAfjQSXc7zmdxS8
Kf4P90CUIDvx7nY7LvVJBotR6LKL8ucjts/220hokf+Y2ZiAnBDaNHBUDLz7mRad
YNH4R7dQ5K6No0Ly5dZr/EGwMbhVTJmTQA90P/qO0Pg44wjnNOQMgV/6aRzI/2+4
L9romSD2wiB5N/9JRCFYhM6qJWkzxCJe3xhm0S3cyBPR9Qu0e87pUJG5k2bw/7w7
xssuGZ8BW557yEmJ05bGhhsJNQKoOOOegzu7qVXlvaKOBaQxA26wJx4Q3ohwjx2b
65eCe0nIStS02ZbBtSEjROcKkyVSWl256mEVcvnp4Os1gR/X3D/qQP11W4atMBn4
gsYwxTo5FF/d5F9fLMQjQHtZx9M5bxqnbVZ52msrirYcjEBXZHZ9TxdEz8QJA8oc
DKhBI35hIk2WLEYf02F8S4rY4Tx80P7Ko4b6dTZL3Qfgia5VEq9u1TMfMroBtTv4
38wK0FRtazFkBbakNX6Ree3keYr/vxJhttcn8Q3V8Gy6Kdp1bnri9IcDTk4ekpq1
JlNSIWdEV2G2bRqlDQ/623IYQpk2Z8zaWYbpNjG0O8WMbmuulof/+Jgi/EokGVhY
Qsoz4uQqPNQTP7ce49hn8B2AzItVOcIcQjHObDI1FBJxb+UhB92Y/uXE6Uvey+5V
8H4+am1Tgj9oM8MWtR9t/z6T9DVg7UowZm8K4EaAEnIuMQLFOwjmjkPcjfncsJnw
sacE5OH0bB8AaFFvx87lFmlGe4ixbopKFSdD1R/9IOOc+SMrvxlHQkx1uXwnmtpm
rL5Va+lr9ces+QEQW1Ikmyz6aCPanhWSr09tDXqM+Cz/zoAlqB4asOhqb/40fhRV
Zxxmqi1b3M/WFV6qu6n4Wu+EUQkGD2FpP+jTOo0ueLcRBGNJdQ3rAa+8CkSxb6C9
W5h7kmHJuSx/7PnSqA2LJn7TBHivR2Rr9iIxrZEOBteMWhBBUemiNmQG/Mq9El5P
/GVpo9BV6rEOe/395vLdNeOQCIuk/X/VrNdy3VafFwVHdNnrIwB2phBNrkfxK8XC
E1oBOUyDAeWcx2UwnMJetv6/elbYM4amUsZmuqBei5KgsWVnoEO5Yr9W1oXXalv9
e3tH6FlOJ8TFbmun2tAKT65ClwYtM0LCQ9mQovx0yZrKKI5vhrzNrFNOj8J1wPun
BwlJwrGAtCMCclmwugnG/TccsCIpT+OvfXVG4ovDTF7KM/C8xNUT1OyjYfIxE011
EXHBv8M2hR+FezziaHJfK6qnFtgrSYymHVrmMxXKDikWdAR94FPxpIPAkS8I+q+T
kF+/S1iE3Er60U7GgEk2a+S9M6cGcxojo6GkCmm3QDAYQCGXXrSUqsBTbt+pURDU
r4GglIMOhMW37ISVGQiHJHUCychoau9pvoBqdYd8mWOLLl7QTHGmyfeJiFv1w+Lb
TeFwiRgW8uZ35ljvizNeojQ8sDq1pqFlls9qujleMteA7nLzXZfz/LLaKTkYhaUT
8z9M6IWwlGuHHpcQ0RD0P8wxGuhDIB8e4PA0vBwGob0AauYg8xipIf2TDI5/0p0f
QwuBFZHUPraG0nQXzQST4M2/zQ2tTx+53Ux1ChOBnUvgV0tjE1Pm/qzjqkkc6oCX
9i1a0fh3L/MbXu49EH9VTminYceVfHAepJitPXkkM9T+6GI9XLU9JvpyQBQTC68t
H2KBevRD9q+BBXIefIG/TQnCu0fY75gBxvbUTnyv5KKmGTYikW8OsJpD2LzZAxoh
RhNnkM0yWVcFlGtmDAwZCW53gXtUF0S8MmTPFDlLbMRrbEav5Jp8yxDPphMrYl+t
G0Ax1YwVEjE6L4U3maSFM/xxwGaHO5zG8+iIw6sh6K7ORSyj8FfRXM8J1Bno/hxf
OYrcVPLWct1na3oFFFHyqauWzpv20TbvwAM24P534nt/mu1QiAI2I3ApXZAoHGV1
Y5g8llEvkNTIbLcxZgM2D68w6UsDcsSc5fwwsUNUH6HWfuFBIbc5qV5AhN2vLGq5
rJYk7aMdT1qQiy887j0khQs87gJIVTXn9EBVbkdVKxq3gOxspxWivZ3kfE2skKqZ
GAEkBAoDw7TyQm6nUN/CzWeDedRMc16PQSOWA3IQr3nR/kV6/s2XG/TXnanjNR+q
p+NP94laajbWXUQIsqD+ONXIhrXd9Wb1LMnB5E08gugC/TF24v91A0LdN1OcxNYF
Pyx7gJ5q3gXrytIfIBO4FRfzy08+G9zyjfA7vDH/jEIXWJbNh4hV/spVyUaI3zJm
81kr1qkLu9637kUGpLTZj1IhmIZZO2MCI1oyFfSHvyz0nTmO7wC7G015+a7i74vw
7byGfjofWY18gKrnsEkOjpbyVXdHSbmPzTGff2PakPsuJNrBosJQPnQjQVx19f18
e1MmoCWfdRF+6VMrGFLFUDFS4B4ySe+ogRTfysMv/3+h65ijdDA7Odd47MlEBarl
8rVaKjgj8paQilLx19n+D+oWNbhzmRgck+RvkhDkjDlWd5JzvTnriZPuZfzSz5+E
sd9kEOwPyR6OgbCmZonDaCzQNWc7AcLrnatDszBEzKOiNLOr3ZRmynCEHmgkDgif
X4SYzlHdewlX+yNejaL/vEbaS8ZZZMfoG9BOLSgIkx2pHD3eTdAMEPd6d+8ENpxm
cU196V5SjcrRkSN3OJDzss6G2VAcal4egokfZj6fjY4n49CojNbqIV7KvTNNnhfv
l47B8HMgUZ/Z6a/nU4sBn6+H6IJBH34+TKLTIRcvDnCIK0b6k1w1NbvR6vivaXvT
na5sdpRY4pt5PNYbRIlqPZuF9d11Ylw7zOmxRf4OTqd67XzVlFwB5C37wtuN0Scj
TzYK4t7mBfLhvD2DUunmUUcaXmYZ4IcVq6Iu9U6ldWMZmX6FM94g/P0wxlyYbTWh
eHafTAy7dMjt5jUf+J8QHSMJXL6Wkt9ENToYFWOX2Rec0uNIeEAdk52mzAizypnP
B5bYj3MTJE9sL7iWyAtvOQfXq2Y0lKI8gQeRk94wBz+fAbfh1JzD49TIbtA3s99+
tyOYVfFGH9tWcZH+5q8AlJCLJ9d85WlJRdjWGNletc5CzxR67m3zGUbOqLbmqm3r
Wl/4rF0wQ8iROS9deVkkP0iaf6L2nE1HQeRqiiR8fyvalRsZC/pke5Lg8sDvRaxD
bfTBxvZ3KGR6yhQC2gNStSLoQpjdqGYThnIJ+AalJf9BahmEhAeDF665MxgVjlut
qkrDjwqLquLXrb6ffDLDT9B3l2OT/NtyfUtZ8xzFoTbLSASkAp8pVRp1Ok5b8Z0d
diA1EsuQCAco9MD6eaR2itoX4NaOtCsFmW0Y5N32fuQTiWYP1+Ku0REWRLkDGKKF
d4nicI4gGkW2UJma1tuxmQ+X7WiuN+ef1Q+i5BFDTwYxSLmqIr2dYilyX47fMkS3
KivofjU75XnTAAhnX7+tjoGcavq2Bh1b93ua07eSM+yzQL1AJvBmaxnbDImHjTXt
FJ8K/aB7im2HA+8a+DTm0Jd87aZRkQrW4c7mcd6cojp9p1SjWtoLafQTZiu+alCN
HlmrDBdgsXD4g2Bny1xkFrNf3nd2JDmTBqRCYNjPDQJ5ltIXL2HbIv81G0jjYtQj
SrfW4ySLaEE46pnCbWCwS/2khmtA+ry+sshpSEZdsJrEuGHf1fPiGLz+y3yAtiSY
eTwCslP7ZjoHuxkJGlK3pSajeY2dilr9+k40Ve0dDIIsUFycYHyev6uxEHbrIm27
CQ28q4yDhpU5aIrsZQV9buIvEjfmPk8E69PTl98XCDIv8cHVdymBn0li9G6l2dDV
9KYO4QvvRwTpr306Wgq5+TpBoFh+XQLBDe1SCUrwJ8ZUJl8Ykl/2KWULBQNow9p5
EBVCR8bH44vHLLNiSqEfkndPGhVAAX3lxbbeQfnQfXFQccLSDDFnsXKQ9exP0b4v
r2OF5+OXDRKbrWDqe5O1CHT5D/HWHwG4w96CUAtx8tegOnoMLCY84wMkXSm3dwgV
hSZXpgnDjwNHCVzMTJaYuYpqnHOe7T5EsUP7zST27BGOBA0Kgs3GbF3RTehR+JJL
P/JbJGE7E58CArnT0qjt/kD6ydbwjaWb+fBc8sFXgmKwqLnkuNvP+1eA8N4gQfPh
UgQfvZ963FJA/ujGiz7EIPuqQeT4VQOd/Sx/bWHltxSVz7dTgWCRxYZqidkaSpC2
v3xkJd9dSU83ZE6K1XEQJZD1OaCuZN7ywA9mZHf0qnMcn5/fq2liKoQIhuZdHo3q
UhlrafxgoCLc5StwIdTTsS18LnCY6O0jyCXym4kok2LJU+Ur6zF9sXfaGBZhK0Y1
C6eXNxtwHw6uJAXzQK/mYGmW88gcgvRUCyKCcvy+7G+8EdaxXL0rYJhV/VG9s4iO
wziLD1oGCZj0AZ3jCZX+AN82p1aHZucEwIuJn4C5BUro0Djqp5CoFEZX0GgzHq2g
Mi36qNxkfr5xwCAInbJkzVdGvGbdJ3Zl3tAKhBb9JFYpIHkoNCvbp3BU0HA8Ie4i
nmHmtiV4xxOgFpK+Cm+ZM0qWXm58Ut2wgzjYkZ+SFSDYBgevAX9YFX4icOcXqxCM
+9bFvWiRB5EZ6Oyxnb+2kB/6Yfy/jReKOy1A1eR5/rfdxD9CBvo6ZR4L/Ry92X3G
cZRGRXaLRa+P4wgEqx8Nuo+om72ZAN8cBEtELynp2gaDMMqnFLaMla3MbjF8wevJ
wiaV88TDvibn4T601Xg9oYz3aEfyPHM3jvXXMwTrLbwJ7fcoz8lM8Uu5Ru/kHonF
oDtFo3OQqVbuVX7F2s+CAAvfBGhwPRmngTxkvbrU5KnvIuUmDV0kdbsKubKH190R
Gzy25NMOMDPySVzsXHyE56annhbOk7ynQ02B943bcGomAqD/wFcXGqoK7V2mk9fd
DtWvDAxG/1NgOiYTeMnsAVGhXrcp1BCrtV5q/IWHCgDPqSZHCzujBLEqdQFr46+r
B8a1BOOfsGxdzk29jGpJXYiPmv2TRLcd7rYdE3zP2Nq5gQPQielLJRnmTPfk0mmY
S5A2F/PePwDZh15hHr0K1NZvwESL/sL3voSRQYjS/r5IGPv7OrZJ4bh2lT5fJ/4B
3PFLHXgvExzUXhxuorcNsIp6EdW8UznEmCurNq8+c1NNQZkxjDBEO1Rcug2vm9HT
elBx9HxxReUAdQ8ffERpz74JN7o3JnFV1kliOByv+ICqr7Wt1PwY9TQrMxx93c67
2q/6bmVSayYjx1RfFY4JWNn9/KyMp6Nq4ZIoycWyzaEoyVA+CJ4ghPhCaEZJBqP6
mWLU0c5Pd1jb09p3VsArWbjF7L+2E6SEoadu4KXHxyWYAuD7Aa7to+ecjULiBq1W
vow+mUxJR7YRE+U3E1rm3hDT2J4UVwO0OmFSbubiCtmFNBylDy7dtqHvmE4zq24B
Eci2yhkFW8wg3+1UEf+5folsbxErtltHYndj45U3BA74nOGA4xVZVWw4P2JRSRb4
AUUGIsSiVEp/QJU6lMeRrXCjjEt9xMUafLVjbX4XEtj9pcN9sKlBHfd7jNEtJoCd
s5seqjNuLUKZrc1Amw0MpNkitTiyDcKfH/OW4nuVpiV8tWL5FFwCcsvTcR5CWwhx
jcnAxXQwvgqRBbw3c6pb03t56D2IsAvfUJPAMiCjJNvPfX/oFLdbY9L80npITknz
AjASJJjs+K/HoDww06RKAPApZEJzMPnHav0+0MnAhPKo83G5grTOrf61z+i5QDzl
NmaR58/t8h1WzqOAyxVJEftcvpMEPQ0wcuLUvCSVo7VO9mt5ZoC0nBL4dXbduFfR
vITINQ8rZnrFrKF46F68igiRJurqqCX5CKQiZAa4LxluvUVOKk1fwlfuQjzbdBY4
QcsRvsuSoy1vtnGrAotfbwfCU786Xq4c3bnW5aX0SOCdyMMEtPepTlnHQXUObiCO
YaaMlr/N/qer/N7tYotL8sI3+TW2uMqnjKL4PgAOIO+Jve7OoAVMizB9bLAdx3jL
nj4mYnFu6GDtDzwZ2Jyr1TS8+/LFq8u8B3io3BjQTGVJjS2BpoGlAql+j+10tR+f
5e4CkguBBS0ES30jS6v42s1vGql3tIV46qlMuPk4ZRKDM/hnl6xRAFEPcZ0v7wSl
ErpiLnyMB55dregnqLXEkzsWS2WUXRJWl+wUyZrVwFiwEkP8ldpmJLp16kxwnMQq
3Ezr5bxN8GhAUtuTfSkpJGq1AcHv5Myq2ODSeYAIpf8Pg3WUCxvO9DOTtBfXbWrH
5fJhrguJN9WbbSD3cc/rtnKVcZsrJuzovXyy0ztGJ6eD3/6HDm5CANj2GYaxHzXz
sygcdZV827EQt6NaWjMWiYRiypo0aQtm5qdXRcQEo1v487Zbytu2RzBXoWWJ8NWV
PglWdwQNecpfVfDJgNcsmvvAAVsqjU30sBnBnsIJsnwCOo5K5pbR4Yj4/64BkRfq
OMNuGkKRob8xBoG42ZRAv8gdvxt09NNiRzXqGksptl3Fb/zYFNJG/qMlCLqEJOVf
KmOFlLVeRyEj+gPuZk48bAqJ9y9mazRcHWqrB1Pv+j/cpMMlav+71WUEQ/b8Ip+0
wqNwKoUVFT5WXCR88ovKVJiLu7XiEVxKFSZVEXLjZIphl0a3w0+/Lxj8qwdREMoo
qzvPGrk2kQGjtPHEWvE7oN1w9ede5kYc/eTwBYnm/ugjCXdP7jQD6Zjj5ymSP2em
SXzThTh0H5QfXKRCOpxfz43Wp5bGvSR4pmRysoK6ANB3HsRUKBzzBzuvqQBRZ38f
fAVM71vAKlDGfZDial+6b046aAyetym4rZL4Vff2eeTAaXpRsp26niYQSAENqv8W
ojFK/RwT8+uljokMi8W2ZL9balCr/stN7beA+WS3nRpPWnurz78WqiOid0SaEouL
vxdipK+DofHn0WwURmzSxEgQr8/FISkBtAG3dVJe6adhCohJyozsnhjCgSEd2TGD
CZncDBakpmFxGw8d01UoM6xsTNuGCcwq47gFypd5gUnjgp81TTRwYAS2hdJ16pBK
mgjvCyKdLV9S0VodIK9cVFnM1H/tzdLDH1d1ArEhsOC9/9b4pK27HfbtWCfPkRaY
Bvj5IBrVHjLcq0uaiOaJ8AevNX/Mr6CB0bTlBYUq+uI/HCRV0gyBsUGQdDeR1ixU
CzxRX683Q3oy0rpqyJj2DqAMV5qIDZoukEqq0S3w8+Xdib1H6a7+SXEjKbwokTox
fIXJ1dgkGpNSMm+GZRK8+I/9O3pG95hVdYxPgI0gva6bnI+0PY/cTkSUb7Uzsk5q
p2YYnymiUJ3rRqDF9hSzBe1jS1X6jR942qalFFxANKmpK2WN/w+BmNzulvw0yesH
BlUIEtpZ1kGsOsSDgnYihZX2lA85x+c5bftx1he9mr+UnttM5Qc2RbRJEsT+otno
JowSsAYn/Si7PaEz0Cwvhp9nvY298NB3Rfvza1uWxYL4HC6BNFspp2VsehWWvxNK
V1OTrxZGdTm6BkBLG+FjHTnRAj8U3eH/htLtH7iw829FiDQ7PQGK7gVCjGl7oQML
Pp/77VrV24hmM1ZbvHLRrQCgThEaA55j9ycR0wmj0JA9thf4XVCqSOpDQYMvfXks
A2J4cepiYB/vcRYFm8iqgtOxHx7ZkKVCCkvYM6M0YWLeV1MIBeycaBKe1+osxV1Q
Sxwa6qYlPQIn40KAqHvfklQpePQ8HTswbWW1DPCRQb1fBR1l4gyJ5IbaHz/18v62
cT6Ogr69715DpPc+KUn88U42t78mT0NFZJX2Q5oc8eI+NsK3Tnra2E5vtZKGEOce
U6QbiKtsh4eylKd2595O20lkaiNIdox3BX9wPfKe37oZZO1g0/sn4uExMOtVzfdN
O+iktaQtWnlFMEqt94qtE8+AHrD8EGeEERcpaKT3pV3DmATcrbSISVb9ADB4scGC
mrn2RovoDzoxmjexsTKwDHWnsq8UvU8Rz+4OcN0TbPSnrG69as/RB0HqgsMtXxdo
2Lj1QJyVJbaI4ceHYORrfptlZ8k7XKx+G1XbhmPwzM8Kk4Q7y/OHV9TxMMG2MSn/
CCN8fQuAErK1JBAK5eHSQAgPqAsaikZ7kF7wvLr7LeEOqD5H7mzRShFGwOc4fpVN
YGHlYr7MJral2ScN4ASJa/JvXIm7uOqy0343XxUI3PGzsN2v4HY1nW1P9o43mMEP
H7KU/klToCliHhdrwbQimsnvrHuqG74ScQtsXJTSntXghv/nUQgSbkYCmTEsdasm
XxxxPpfL/3Q0yxbv90J1VTStnUQ6gf5iesqDZvjEsNEhiLrXibJOkopGT4iS6ow/
D0L0ULL4ZJMttfFSSDTno3sCV5kP8qFoLSu+hyVTArFe6kpnPPR+uIBkgFyti4GD
RqyizLO8WxcIl7k0ewXtzpJuyg27DkYGolFCEi6ujbHUa3f5v+z4410pe9NZfehe
MxBvaiZjaejVmBMjf+ipAvbmNOEztOnqAvHm62UlTjgF4YBBE8dqAd2HrJaAHk9Z
gpgFkkS60UKCnZHgJ72gMMfrsntMOwUuwyV8Sm7/1zYOkRdaHQ8MspobvjtWzIR8
r9BDg/e3OhBAkIPwI2tCR5VD1FOXdsrCS7eZsHOpQbekdYxTDjE8eztbir2yYJSf
QUGa//Oy64bA9mazRBbY6a76FJB4k1HNiQlr2if0CCa9Ld9rz3UjTxVkQB7maSIp
OBf2yxue9Zf/+h/fOvEM3k0pBXW6y5QGLYrpTZRRrnqnynKHQkmS6h6WaI6Q+q0Z
OPeBqlU+f0sRr0197SUZs3UJqRQMlUf6OJPCv6cA0MdbvbukOLgMqOUDT0LTmXEk
LhqYFzwD975NTXev5PhnTF4iN8adlv2gfJUR06YzhTbgbFjVZVSOzc1jmzn/TkkR
KPEC+vQH/YuXEnXfD7qpnhDpej3DDHE2LlcXvVVlLM8QideNhcKK/6zLSQTl0xvM
hNDGHO8ym6/7KCsPXx1Z4GHBBEXEOcnSg/q2IF0/eFC1v3X3aJtUDsaH9gGwR9P5
IkW7Wjl0Imy3vRTqqK7y4C6+chXyMGkV+rED45x+ouVToqo+xx15j1aBRbeWV5mM
JtedP2Tgo6GWfBLkmp96yutKThbt5tRxBHqzcl7xRmZaK6K77HJ8itBTh7FboTHd
lNBqi3QhZqhEbTDKdflwJIdT3Pm3MEioNOkc1ia5h9PM8T244NvHI8HADr0VP2h6
SKpdiSL/rbZmkRoNXYo0TK+/kblQNpnidUhvexRlyfYhoNIyVT35vCt3nusJzHnu
0eph0QdecWy2SmoyIYlGgRtIBYltp5rhnM/1QnxoMyvwMhLzZqo2IBIJVs4lc00g
YSBKXAdvzvRvHshkX2y13scA5Y+3K+D6lJqtISJ5GskXxsHa2R8v6Z3DKSVgwFjZ
4z4uyHrur0H/cky6MmyM8SyWQIekXu3poEg6OtogboOBKo2rlj9xnWZVSwl9BMQQ
/srgJd2sA/JO37Szq4nv9bUoQA8idjUnpjyFSrQxicojifIAdR8ZJZKfcf/vVsrn
3W0qaLx3YbE9U4aMVass+Bt5bZbsk+a6kNP/G05NBmht+MJjm9NnRUgqOeamN7Db
C7hwO052lNpxaF/0kpHx0dXD0Nl63ajTCEjKWCD7WkIcaSEtGP7ga+zokax+BNLA
hW/w5HOpqpYoG6RfTOrO46KoskktEMdpThruENjek+o9qdd1diqt/vSK5U78GLO5
mD21bSpx2ZljesMKpIo8/RDZqIgySCESYij3zOVtinJgVkc9KDAz/PEo6Ab71/Xw
4UKgq4cUpJJaWE8GHQEmqCWmd6xubi9JvjESxwxBO59wORIUXWvU/lX3R7th3fgD
EzNq4n32qEG+9wdrBnHxYl97uyadk4imKOWJPr9389l9juLAU1lNYtjNS0J0I8wF
gDU4Z5Mb551VuJyGGlx23s+TrDdfiTvf8+Xt0UhaLkQNXmrUyUP4pOpOjhBAptPv
F+1PNxCGMkA1XGDO27SpqJ/tcmcuaradj6cdFNUQk5OXseJBLNerlETIw3YqDqAq
zw7WRu1dQ0WqUr9dXCVuV4Y0jpJ2Pc0pgZG6Dtl5BXk3EcLoIiqSxFbZtjbDF/bo
JE4X+oEZCML3VZq07CtpTPL0gBywBj4mIodelHHiD3B2nEWuG33rChPPBshRnZoj
42JrcV6EN1mpSh0AJ9/XD4Y1ptTu9gBH7YN4QnLWRAXpr67IjkjhtL0I3UEf/TsT
G+GYlKBEDIREgn+SPeu7vvZWt9JpuRT0jw2Y6oLTFdB3IWMIu+mwmAszzCgSXWJt
68tC6eS2z40ZPF4lI4janNCgT7zVZu7mSMTVf0BO7sUfcu8mH+XZqCwhTfSgNuGk
JAWO/xF2LuiJdNEoOHx9X1Y4ueQFEr2EDDtFv+f3WRW3NxtvZkEyMX2Tp/8MEJl0
xD/p/geuPSaJTVX3l1zcKKOPXB+h7ET5ikFftIbfnY2+97asGqPSvTBChDttQVdA
n00WA/LfRvkeBOd8j7kqdsCYE1BEoGTXSOXxRgzIOB74G4Ixmu1hhGt1s2PyeZ7N
dq+Q59Y/ilSw8ysnq1l5Sr96V3rxxDMwhFucDnIBfsgDlibSCDevyiq+ezOJrIwO
3aTbfTdtIIVNZuhMdw392pk6/Br0o+PY8SDr3AvF+8i7/xQ8JwIMgHp7iDsgXhKO
vS6/udONeNgNuDBNKPqUiqxKZfGNFQ60Tf0/8ZTGu2k0vYYrOfwAseqV3MQfeIdE
dT+L6zIr0mPfaJbXtTP8vU0KbbIrdT1RPx4Kft9HPJHNUn1HREvSG80dSgFTn7L3
l8LME5oe7dQkwDbU5AMmqg/GDp4ApNla0l86WTB6XRP4Une/S9Wp0pL2vnc7u+Xx
PnTu2oMsIXnRy7wKKjOdb+ookkTMmgce0fyodzUW6L2j551sb32dZOAuXBT8lfZ5
TLQy+S0gtjOR4xL48ti5zAHA+D3ghpGyKjgcWeyqzTKFjvZl2j4RVuSJ3RbpsT0u
eNAZAR6dKMiu103eWK/dFozR2Nn6MRCasWHwU5mEyiXnPqtnaqbJRKo/kIy4FcrX
6wrAXSBjD57NY55uNMXgQwWG2IjwmkEb7dl5W84IEYucDFUjgOiHNXctrLtz+1Z+
53QJoUasxjrUabQHiJF2KccnMyrFICMjMu51HGNu9TJRErbkfncB6eQcPB6/FesF
45/gY/sv6OdV1JX1meM6PlHatxTWEmDY55juLPgEuTY0R4LmhBXQ3xhsHtPeSZvf
4qfhL5rtw6rF2zc02eNEtB7vU1etlIgw5B+2IT8q3iHaucG8KMgQqYPJvlXe2Qe/
xco97njqcG+a8qa9BN4KZ1atRJAoMmJlBaejz7Ez9G/8cyBumJoMlAt1Ur69w/Yg
JGfGyCmuMk2rj1eXwRVShfC3IlGTNNDyQL28xXxIO9L9nrqxqjzEqiCht5fptDKh
jYR2tKTVgXw3O1VSQsvE5YR3cARIziXnHw++lPz8YlgbX8WfqRX4Awm5XlgezGCy
oa6MJF6BRB8uH154Ac7b9Jr1SLVt+/IJ5+oa7RnCZaZBZK3bTC8lnv03hftFMOJK
X60bV0jbCa4OBwhARQUKbs55LXLSbUT1LwlMwU6spndH5t2kicOWU0cH2LCi2tmy
tkYyitsTr7sNu7BoDy1Jha1B0UtS8GgrDltakWcTN94yNmm66pKtaReMg5HmjPJF
aeajly6ne5XXS+5N0eDiZsfC6C03y+BrRG+nSE8GfkxypbNhJb1G3ps0HJPLqYyP
U1XBsQO7XiaLYckkvFgrzH4IijQY+muxD5p+16wJlPVYIeeF0LFOwhIZC2t7MWsW
u4P6HBdqoqWfaOgG3IQgEOvYUe/XzeA9c/vAu0Pymm4tCg7sFId6kbqjMtKD63TN
jXqxWP7jTUqrQMJWgXEJI3tlEsAiK6dXSN/o6xRddHt5NX9ih/ylSqZyBIjrSv0h
GZm07+H8i2XG6uevAIouQUmd6oduEDG6qa7hxXqJHvOMgBAbI0xFWdVHssODfnMF
2BYVmS48BjIWYpHq2Kpf7v6udx5Ms5TeYZRq/AMWcmEZDf9wvjeOJ6RgFJ0EswrG
bsIzjTGkdtBwgDsA+bbxFTEzJ+8QQ7/fyoUrOV2HGIpLGz2SyRBAFwfpc5hIhjjA
0fGPLL2b1SQj7r4e7Hm0lb0vRE1bn0YNCPtEKSEGtdzeUhMP8DuEAaC6UoPfvE+/
CjKRT/kDKO0cEjTNbmnrnTDNiESeKIoR7Yq9S3ffC2GK0j7ywL3v0u7ftY+I9JLq
xdT8MKvAVd9dvwrPNumPTD1DL8+KTyW9p8zHsqT7ApB3CBVTyx8aiUi888cbfdnA
kyW/aKQEaMj/OQFgYOgR6c4P9CmElBosiiglNMmlWZ+7lxMma6AA2iKXScK+YfNt
m5B/zYJwHq+zNZYunthKTHoJHvCxwTzC4QueDZANLzFbDVsZrVu/Cv1ZquJhs9/1
S3b7svg3l5jvIt/xMIZbgU5xQFQ6JiVwoGnlX72BOoKzuYYKmUmJwIIH7YtY4abK
OxU4jza+k6hjKPtwzbu7ar20ZSNvgE+Jo3UfivHGVdvm9n0Gz/E5wrvZy7it8lcO
ctAFcdxaKHgwbwoUrlrzAF/o4ZfVOilcbVrv31EQhAk9JgXr3BqIL9QhvHvihcvT
0qrDH9/rT/vPCBn0BAWeNv2xFkQpfWe1M9zteOEi16xycWLw+Ow5/WQquPvK3JG0
Ef9ntR54F/ajgodP2o7gfOZVVWFgIN4b+q7gU4ED/EVZ1WaDxQ4heIaDcA95WC1f
2w+Y0tsg9dlh4AQl124vlMfyO/kd+/c/0v9NBSrhsQWNnZgVCfUpeAZDUkgbQ5Rl
autq2XUR7qXybkxbN51vCB+i6CEpjDNegmuUnK0paGwODwvluEuTm0Y1OdMJMrji
4L2D+zKr31lAJCIJ1UCTa7Kso9hjktsSnA2zdskmwt0TBeyBJaZ9ErCG7VQ9nyHM
tCxiqeZ2wBozAL/3OJBc4vASkCM5T7CeAWVs7iVTZ1pC8paNY2D4plic5kzFhmCX
U6dWeXTtOAs3js1adAm9wXeiimAB+y/dlCIeLOG2rt6s5jANASuK7bs7ZT38kJKo
vXLfbYLYpn4GknX1/pi8oykQjNaSMxtCKo+oai+Rjl/K9J5NoQ+OavZyoSKh1Ram
7yLbBTzs9avm7WAsXXusRQ4AWvBfGWn0SsMKfbyA2unFju/ogpzeNw0f/IGWC4Nt
lNkwnT5T9zLKn6TsCEeWzqpGqqhd0sSjVcdKYHrxSLckaRBwqkl2Fw+IIaj0Bi61
tS+5eecYtuteSB1XMvi+vtE5ztVSvUI6+ZPyk/8F9uCSYNojKC84hx1gE0iZ8277
MgZn1SgI0vNp1Vlxs1xLm141t0N3EGFvz1cqyv/iXCmqD0cxVb95LTwY7kqWbocd
P+LbFAnBqtHiCe0TiByM3pvl03ACsH8u1kRObq9V/Rgn9R6jVyb88HF9QHTp0q0R
APHOtVERjznNRc2YyCn82djIyDvdPdCDZlBGsXACcCp+09ClBMrHX/ttn+DwzysT
eP2i/wQFmNu1O5n9Uwn0m4+Hxc1eJ/rCTdVlWbQuMAKizAc0izyFHnHk+6JTopv3
LC+H6QKwcl+yK1Vyo/VKFwu31K+EafusRnCxXawC66lEGXH+jwo8/fYpqTyGNVQd
Niytx/fVGd2x0wG2KQsv6CUEPtNO7WBDt4hNmuXUpC6UkQcOtjPx7X5hKQebeXS2
q6TBYKdqrwU2LGv6/lhykEBwC7Gpgz4vEVZYvAplO4OZwi6BmYGOt8yzyG+DZgCY
a0jrfBYdBPjjWQK73/d/M/tGLoIsQschiPI2c/XuD0LZ3g4pgVOm+gRNumvkDIrt
KTG+ySDZbZNgDg2UlfHuQI5uu/lTkgHjN8RYp1NIVc9rAJDToN7VGxuB6Pkx6Piu
84uUGgyHp0p9Y/169Esc7cxswdCnQnE5DiRAAB21Itm4CBT2xGskmSlMOx/9swG4
ABtCIdAmnd9Zk9DXRtOc/u2TUdwOGVdKfRHIh11WnEoDyUuTcahtMzcJcoNefP8m
oSSRjjPRYLHcuM+RO5TGwICti+qHQui31+zSmAcTceZ5k9tUB3j8gakGMqmSoMi4
j9oOFZPrvf2AzLisHiZKhFJWdzLTt/jG5ZXibDFrauZgK6viPRDWhUghCOt6KPqG
58eAsvJLSM+Lc9T4I9tm0fGhYLy/wE2qQBtkYUhTA6n+MTghJzTc7/02tlNZoSuY
vFRKOYGdnYbRO1XYBSBXCCpCzn9SYOUEATGkR0M65FKahQJkTT/9U23M7YGKhm+i
kPJZzVY6gBWynJuyf1pIufwl93LjfNiBNVJ86bkuBLXFX0d7DY4UFru97iA8BQnt
7Fuc3Ani9nrrtY259zCbfKU48BdfMoeeIhJYp0J4MvFXHzvB3IsbW9P1lKQrfZog
eR/TjriO9mrx8wv/fi+NWOuUDJqNydqGMRtxrOL6BAZbksOO+e/6F0HDtHezWKJJ
wtHdz1JNH42I9aJdzASZSF6PBBgSlg2sgc1x2xJv2I63ut2sATTbYTkstTc57gbc
RVyjcu38gZjQgm7n9H3BipqOcQJpoQqB+E+EAM/WK41EVIGcpfvQ+Kf+GaKSdC8Y
9rH1fqrl+EUtH+SVPcs3vBFXy0WdDmzhJRiZepQBMqFvYaqVG0iBvWZPHQTeuO80
ASOMt2rvCcF1MNWcX4tuz2LYIrfvuyRZBLFd5b0AGsIO7b4LV1IKl9m5b8JnZChj
pkTwHlhQ8JrwsOPckyaZfDuSSrbYiVHVb8YZR+WhebNvZjSS47M6dxwkzu282n+7
wBTlvwx0sGYdjfm7EnehP0wDrJHAcn1aE+5QIX1tm0O2kU+9xRHScXpctTmhcpVM
typBA5huGABfEo9De/rpmkCL1LC0gtG8ZlejBQjx+HCXzC/2m9yADtXBsjEcqMwd
YDMklXPfvkHJWY7Xou1XQIYndXCo/u5JUORelXHe9WiK0yYctXPP0LHgbIZzZqLK
pZ5ZjNjYnwFAne3AohFxAwC3csU0I32wgJfWYJqOPzf4VcHUpRDzrtGsJ7r3bBqw
D7UN32Yz+yST7zQZQ2aRmUWiYVpK9NhVzgHlt93ifz/aOPStRwDdyNL0JuGD+A88
ITnbNVXZ9z1/oi9Aou61g0ohPueLjIlRognwFyPRcOcJyPrVWxaGK222mRDVtFeq
svQVhu/rP0Ux5PhDjHFC3kua5q4+HxZ71eyyf3M90swEhwV71lRpoiiD4pqmWt6f
vOzl2NR0spfZby05lkE+2e6HyE4GIXQieWIPFNr9Kq3EPQPH6levrtXTCHtjQWZb
uIfraLjcpKgogY45r24hL7sONarMCF6CVvqhF+Dpir5REOikBSTmgLukTuWPULmr
UUsb+OX9CYiBSBlZTX36RALLY/oAjVd18KouSB5U0N40RuB/sDGd/9BPnSQWSvqP
baVvALLr9g7NswWE3GQGKahEeMIDrwmnKTTaUtThlBuolq3loVeQLHF3pP0rbK7B
fjeQF4yh9dpxwjDmT3D/uC/bb7QmnAXfU1cEf66a96GPzPFLjPP0JMka0I9oUv8f
hfteg3xREGzZmoSb1MIK7Dmee5n5YiQRvoJu18FbJ32/udvIxLuRuAH2mxAlx0NV
FPlQkN2Gg4JU2rZ60x0PYjZHqX3OMNCOnJ9b7k7NufMyC7qFLPSLc/vcp/eeE3Ax
wvIV4yhUnkeOTOexlCVoq8WQP28OOADVkqyqmO8FeYqYva2cD1YT47hWUtmS3YTC
hqCcOd7yMCBm1U1lrJjhDfBFImAi5piSHqnxkH/wyFtPa4JsD2O8Wqt4gge8jnsF
fsigB/pQijuTp+R026DuaWucsP7iiVuVP0QK6VPzL39eVd5qKmTjtKinLR1Ft6WI
IyniLZML0uTPb7jSmPDi4y35ns3aZ9pGMpUV0WVSeqa9YySMilekV9pqr2XU9CI0
c3p5hdYU3eq82+YfP2/gjdGaBtiD18oJe8WJJsx32yEwnRmwxJCOgZhSsJatE4hh
NaTVPRQ7gXzalZXaoNnWQTGuD/yk45xtCd+BK/OlGzNdWDEKgz8wXe4z061iXXTP
3D6+JEm3+fggWWN4NOmLJPHElVuYpx7jiPw+rTK1uu5OR7sCRMD3Iz/domOh2v5d
Nwq1FKevZ9qRlSjxNV3w0fuvL+MCAvYl6IKTS7nfEqrsP2yvX/T8ht2uE4nxJ9Tj
P4xfiE6vNVw+wFSEk8NEMM3nsJ5/PvTxrJ5qCgUdFkfAOfSu1g6Nqz5fVES7mGX6
i0D93B2plSalexQXmYGatNzL1lhoAj5JOYvAPCPW91BkWGNsrAgsxUtN0OnFt2mc
7hwKrci9RJA+3AwY270LzA3CKlLY8cLZvQGov7IAWcNqj7Vw5t7QpKSVhQC8TxQ1
Yjemn3evTyxvOJn4s2Fk3dNiFYPJ8fTwux9xQuG8t9yQJZTIUIzN1lXYnRaXoKhI
sWtZqePk3bABERl7Ih3RD53Cg/mAMuey7K9T1x2IRVnSbZk6cAkGC4//9Rysn4lT
qIzVR1I6VmYSe3O4RifEaWFSrx5+rmH9FH5OPW4WYBbIoaMMihc1OT04ii2hqfkd
eUw5a4tH0AGOzhfZkORORvQ+bpakBNrhjuRcjGHlldM1d5AngAPcSkLEsurj9tsu
tEK24gZVJySM5HulUHv5D/lUb/Xz23N+8D0N1VeYbzlXOw5VhL7szh1sBF3Uiibu
EmAApiupl9TpslnurHbXWeu/+VcuUIKKY6jVAupQDBwbf/sBzEmaDi7ByR/spWZB
cFUEnHP156AAHDC1M5J7oSWlevmLevu5IWlXCRhTjT7PVRcyN1ubDgw62HgeLu2i
HF7I2Y0fpho5DFQKdgYbtvZwByrCzS7xEhPhSTfi2+jf5RRCypcBifh3YjdsT1Ga
N5m1lOfLMiKx+o82Rbclmgr/kpaJC0e16m1WeWQu8cW4J9PrK7DQmkA5f/THd6BD
ailmF8sR7GTgUMmWFN5gERPOdX8iJk7JgffEaoIqlKa8KrImOzIFiLc7pwjwT1rM
85IPjrUsA38DsZSQbDMFTe/x672/6ikrWvcAjJj1Esw/DAhiAwE4SvvD8VaBkR08
CiOB2rHV/LD9lhkl0bOBCoEtQm6ZC+Cto7Wi9DOQz1/1MyYXteFTiwEN7gh45JAX
cCmvZ5KFUe93HLMB08/BHjAHz2zpZk4AW9DBfagmgHOYqaBMJGsuKB4zduYYsidr
DZQx5veEgXtN12u9KDVzPECx6e3qrSKxGRr7QCRfi5Ap9bTb9npaSBP/FCTS/dR8
F47hzJxO9DN9DXjovI+oHXpVIfcBZeW0p5D4Bnp4TApLiYv7lEi8wdtDrFUWYAR4
QMYsV77pVO3pTJSLP5/DbdmDTQruzwBIW5xczzeOSlKeVDwMPNtno7pHxYPxz1Lx
Wdr9zhPydqlupCMhFx+MzxhhslhMaNecPIx80Q6ICmlwBXhwhNU9rteg5+qrc5vR
FNSYw4Xnv0gTTWi4rjaBjdvWut5IyU/Nrq3OMnVrlCzK5GxJ6nPkkACcWN0UD30y
An+sZOaKcQaZlhk9K+WlL0QiScmLzcjmwzj6+g54d9/KPHP870BzYF0bsve89vNU
c1Ux0IOPuifMtVTrHcVH1qnM80Oc5nMBXbsgr0oWedX1A5BfN1GmknqUkFcruar2
qBQfv9dO5FuWAtaqbIVciVvdcdkw1FqwjwXlXKH+n6wc/Y3+DVNlpkNV/41Y3Gye
AchRrFUKk/FKE2pdbIlf7ndE+SK749MdxN/vRGwIrQbAQuZOEr41i/wBGRo6hDCt
/XWYM8FGwgwS1HMc30kUlwvQKCOjSN4QXVjGyLXlL6o6Qqp6uBvZetZW481QrOL9
iZomU0LM0LcnxZvWePQdc38knujVvdRBSbL7i4UiiKKvm5YRE0LZlYihgRd9Bits
4x/1n12uYRoqJfVcvBcqWctZdoNiBYoS2nPBUDIwMRGyu69GMD7a7VRY/feI2bdY
MgckHKLWTmsCqTZk8RqVRw3bybqry7p5QIvFvVh7P/a92TxWDhRDeDhrdu1WIvXN
mM/qL22EW1V/aDlySoZeB9ZolWZvnefVLoyFrq7HF8ARnwlnPyrNOqQ5zIkiutSa
3ayTq1ebAYQ4Vwal34eDmcxPze5Ils2Q67rNHABwuxNozPreJIbl7biP8GdtVaai
/N+EkxUAV7vGFOMtITTHQa0nwOB75PODG1hH6cUViNPDEUk30QBH83uFXmakCuCn
aK+wQm9IAnCCS5z9ezmljGGxxd0JoaJUl8B/wcQ8odP0TjnMPCxPZSod02ED1N2b
1VWoq1MrKe1/gvpvZqQ46SExxYLo0Ne4i8Fw63kkddavGq8TxhS/dWVDEfvMCUlT
sq38WgfuhbsmUwLiuHsl5aRCEz/NPIk9q+eOYmeDSPZs2zWLs2DfHZtvN++VlX6t
qElL4fvckBgPh0kqq4SJgOpGkgx8dhdrkGcQmxnsIzfp4anTHB9RqwFWQkXy02YB
zf5fLQoCaZli/INQ+L9bigod6hYvyDsOmk1FC+pLgN9IE0o9sCzD3X87e4gBuO/y
Nvx7C4wZxoB22YS+PW+Va0JjMbkZmWsvxixA80gPebb5PstCEFnzrVBd/1TbPDG0
E71cs54t3Xrgr35NsyPZsOKY8jg9isCiIc5oXW97ioz2yR7l0ubADBO1Vo+HyOTv
XYOZMDHkZSpOmOW9eSwbXrNFHQDuEGgw9ycTR9iCryekZiejYL7uG1HxhOiNWUR0
xmS3jwlXOEnTmObDRjV0n+jdrxkMpV82AGczjnvgJvTp+RuXbiMGfRRcbNMHx4pl
Yz2BaNMCT18fA40uJUSOIH4obljxQI6NIV3x0SpyUzl+C7Om1IzxBdkvWScaQ6TU
FPGPnx8SmAdj3m3F6+EFxUPaEXLIlk8ojnh6l+lQEdvBa6yOWoElMHl79FrbBF7I
jcuia1F97uSy0nCcgx4KhBoMeJbJDO6ys0ZoTPPlu7NZXG6NjggDdrnSyNeM6bkK
RhHDhpgXNtQA8HeLR7XBaBfhqpGR31dIn0Kgidh4Gat89r0Av+aiBgZAin1pVO11
Z8BFdiBECkGuzdqenDiVtr52FC4XpTG31U/+/xoOmrFBVAovrtEtVQqkW9N/UqRm
VzKt/zw54ok6HTM4NDZhD7pN4VA9Lyf51++Ky/QHQ56nCPTiHe4QeiXBZ8fGXxiK
BBSo2Gn84nRGDU66xcvKEs44zPgQSW3G86zEXxe2ecoYLj2leGeIIWvDJgnqNK41
4j2vp10NTB3afxYtb/fRYThV78d4mWt42Yn0e1N9K/vGD8yclsmhue43x4R3Jlhj
OpRktWdE03ZO+aFJhG2NJpyq/yhh4ynyzdgOZ7ZBE43qe7BlXtcf+QcwSZs8TnT5
gHseODM7SqbKLm5KH0+rDPIcR80uxE4oX0fx9aJBd5ZMpI0PQFIKgPRHDMPV4zyt
LT3j9gZGPBKfDVTwI7T7xeHM4m2oGuJ7vTAXeYQzrMIpibD4yc2kHfeSI8MDtl8R
sLp72lKj8ktHOX5YXKz1KbaMgDElBqXPsVP0qbLlprNKu/UIo6LS5j9XXE0w7miF
9oqYmrRsB5IABY6NHLlSGdNoYAzb90ps5QtkSWlTvylDJQ4QM+NWJpTEK1XDjuJK
mDBpfXFTgnx3ivwB6Yb0A0hjnTe4fviGABU4O287SyWKWutH2FYu4Qu4rgNJhZQu
OGkGrTKpf+fjDbW993o3vPD29nl8ETE57a5aT/goH/dYJm6o7lF0IZL/vUgy+GoD
P/47wbCMvxN1Hn0T4b0xiRY7Q4jCt3hvKRGz+cMFQW6ZaI98iU/cqNVMnSokkht8
lSIerPFiSm+nntxdn3PqDTgtPWGkkqxeZEgey+rh43gd+yvVns9NInjL5VqzfU97
Jz7zM/MDKODGJwy5L/62kek2opnpidSS7vx4wyT7v6uLaxW2cJxbYpkcSj81Mlva
9Gj4Bb5E3i7A6UsMUMlnp6MTF5sg8h5nnzBgFWekEB/YwQtO0aojImjZMJ8N5CeB
fCFxtlwqZ3LwgkWbTOTmnGv1vAjL9QOPIWhgRkmyCsMNXwL0CNdw9MsLijo2QwfJ
uKKmXJT9DX/tJkhcmokmmt4akavFyekhGpofUAxbMt9tple19jHkVP/Lw+QZ7gks
bGf+gX61DAi5SXpJMTAMu/weZhd+sQL5xKIN5NqZqhbD/JmG6a+9v30q9RlwCMe/
7MSVyR81WJy32uuBpXB5Taksp2fJjjDezxTFaL4Dl+rt9Ms5U1YRJ9DUZod+qR3C
AA4tWjnkCAgSx/MgWv3fDexWRl+rGEX9nP5CdO5SB8zNY1rz8NHrs2Uav9Wvynmr
NvKAtA36jsLHrX0yLoXLgYR+br+esloouF/Qq9GUR95THrbtniLlzdqSxcPmzRY9
RD+FF/4/ZRY0ptwG4AZTJKxKipNzZV1GyheaDL5Ci4qMDYqCh7fUQgfrCwSS71fq
B9QAvpRt6QrMmiSxvjHv8SZziF7EqUke1IpptND9wEVSBqn4sGlLJ61jBm9XqQqI
YfNdt8aufPchsBn2LX2KTyCZAPeruC7e5yZ88adOSlTGkIesDii+IxWpStRjzExS
aj1s3xJ6+zM7G8K5hvKfvTRbp6qXVq+Pq2gFAefIoQ875sOaFPCqkBCeVNdeSfes
2E5+enp4yzTpLWxmOrrSGHarNd7jfh29n7rrDTjGxfjhS7/2KzcWdVOFdSexNEWL
Kn+DCY8ExfezWl0JniEC23CcFcb2urHwgtGvVgB9i+IrHAVIROmSI4oAzZTIXfC8
w0IsuY978yd9a0Trk/JUfYV5VOzHRGhDdjDhVWs0g1blrcE1T4GkAlVur838lPD3
1HZjf4rtKApTwEWSiS85Kazy2jgjzBX7gfsjfSUmHEXxzYkwq/yeDxU/w4gWC7AP
QlEPz0o+Uz37Mhad9J3VvBDFKbr3dOjKPU7YuFDZcuALN2WJ/GtNqx9O997QBqsf
qICgM3pZGPFUy0rcpnaTQySv0lLbXEXtK8MkC32+xvl0MzbiIpe/s50l7ZSklj5D
vRxEUtc4ZHJt88J/3e9S3Hz7OsGQdGS7426HdroAf33ymUlBLIBvwzwvN3JM4fsZ
ejHqUkpGOqF+ypnxedDioVij7TT4C8S9dmv7b1vZgk/RGjoF/f9yEbcv5h5iL78k
iYS4IDDsGZm3SYpOcZ4WcqmPLpN0WJnBYCNZTA6VpXw2GboPL2U/tmyGn4013QhL
TjysgQhNnSYYixE63yhaRJENUvxEBC+8nifchcKiiTlbcX+am/VdoDvNf0WnVIyu
HUXpio0eQUH0mX9nuB66e8UPQOWyGW75nkAVkvp0WqtEnstTAqDv9kzwEPSX11JF
/hV2FuGOefGmO7/y0iPtXwq73KQGcY6I4CTXZ2J5wn77F0qcgxsZfIbUMIumWtgD
DSSQpCVrSxIzQ/g5afap8IjRKyfIaNvzFi+s8ehVaQh3lspmHBBTuj+PzGjVzYgF
UQCfNNU1aikD6zUgCpd8CifqNE5Su1jFXzD25269ZtssDb5TJVA6oGwoGTEmn0hL
At9ag4EImK6GUjCM+76Lg6ExYFWKfx5THjBtgZJ9g/whdV6KFBMORbD1TJYvSUa0
mPhgtQCofD5ubm+6H4p+RwMBH/gLT2UuKbFtCrlsVFSXH3x58e+rpiXgrmFnWjFk
f1nGu8r8sAAu8FfCnvq/RiuGQ7MRXD4kSm1hgTqStHKcH9sQBQMf+xw5Ea7CujtX
s5VL4qSI+nSmGpOMzjj9xUzJVCgNci073KSAN0yqA5U1lL2+7Xo1g8LuZuVJohZr
eHg9N0uxhsPRVMqGn0nEduW/cl1kbOrUndzdnQxH7CY8Jeb7hhIVaIvfZ8veBGX2
x+XDQQdaC42fmJSGsVsg2SvHDEFQECc6XPPKjV2jpwkFs+3m12ebv1VdZklvmEVz
95Y4ip63ChZZQj8jhBPD5uQTVjua8BVm6/83zkhSNbmrmzgpqIoNT0yjkmSmPyHf
hhxfgHWbe2oW9z5KZf2M23tpfMH5yBFABtSaZXPmKHSmL7avVU6hWZpwF6ZSTU6z
SgqfzhMwLWTIfqZUL8RfNFotizP9HK1ac3r+Ko9Cgfga3KKHSD0eZlWtUYam09Bf
dqu8xf/HhpVVEw1G1uPl0nC0v7xfnvtcMpnrFtsjXqoH4TXf5botWBpgMu1/NeyO
OrW1jY8wtv4E0fhAZUARLveMyp+6x27VGkXKd4qTco+9cFt4G4Z9zhHsHsZli9Pf
NNszYdxrmf0MkeCCzjGQLEk2mbwVADZEY1JTE63rfkxV7iJJY3wYDRoHr8yrcR6e
SVV9VwvovFlLNKjNIRl5aXAkTlWP9Xw9pAAJLi+e/H2GkRUcafWFbkE8Vw2tJ/Ik
JLEJsomtxZyKPd9zssmB5nC5BGztwS0xvDOkp9cfLU4qeOfop+rB+HoiQ1M/H9gD
Tzaw7r9NaVUs+IscmA5tC5lUkghHBNi2R7DtPAs+bVv2gcxWPUqpcAGs1FxsPWKN
5uS0MjwYkes9u+W2NH1K7L4+oUdbnhNgdqTaiE6V69hAJPkqUgJ2V06ko+/TLPt+
EF2UOJHfkC4lYMcvI70BRrcUpQ9Ud95BfGMbI28lrQ0Q35aqfM1RrN/q2LW3PxJj
honxH2SUrqWKFSxwI/PIaaTR/e+EYyXk6a+KcmS/Wqgspj3oVWgm7DI+Ql0oHSzf
39oz8YsVdZw8DM+6ztV8XG2WCquDfc2H4LmHDzjy+mt0KZ3RDp3C94hzRbrXDfeX
jUNkNFat4rhljtf/1V302FLkWbOgs3bs/bZrUVu6fsAUi08PEcuGrBndjxxEA9uG
f6NZc3f3EQLT5qCLXbtD1myowuz/7HFmUWShkzw+IaTd4UAr0myPOzAeo12r9W7D
2viZDKoL+ZYTpgE/KyyPciTBJ+qizfeKL9/9P7RYDEXJiDXLzpk/srHCsSCMvXcv
AFYA7QHOhkYZlBWI183n6uyrHBj9klSRkPuGLr5Le56DRPhbLLFD/NAsMIm4EnTb
MsIXxcZzqcd/QT33R4aoJrC+1vuKBgTKdJkJ3FjRaABM8rxaVoN7H4V/21Khrj8b
q9qJLrXuRi9K0I7aVwyuac0UlyG8QjY90r1yEpFnTZ0LFSvKhU5Hy31hTNBAhhjX
xJsCQMzlGAkmkXhyPMUxPtkeADQ777cfR1pI+XsCQ1LhPTsgQTX64mCN1JTDwOQC
KRKEFMDVjfVIoXL6pKJ7NIzAQEDfPH03zjWbYLPDtktGr6rnzwXNpx8KKD87cosO
8U3YX0gCSadnENS0MdIotj3YBzQsKFzKW9hhr9ge7oWHMlKsZGWj1L0VL1pDTdqz
jaQsui4sADCniUDyfygVyGC9ur7KwpYYbCwl3WZ+eK3//soVTXqD4n9hOSBnpSBl
6HTfLkju1JcMVca8NeoJtZ/rpNgOGbjCFmdqZIzxe4BVmYDEQfvNeLx5iIkkUcaX
sourU2v6chIrPRmiPFMSN+K9EKvWtjk12ZqOGKgW6co4WhIs9KEO6/6om7nicZXD
aA6yJtHkNChhn4Ryj8s9OBpIRmIG7bCwy4xldpz8EwgtLOk6uBytvSpniqYb2Ekt
wuAVSBYlkMTnx+MdY+4wI6aM4hfH+leEWQ60mR2p0TC0l7v3B8M5ZUQKk+P75fpq
ED4goGjSVUQosEl5ckIAd7DDt2cIWp5q4qXyF6g/1nT1P5ybd6zeYdp5Lj+fxFJC
YTMwh/y9hefiyawIG0sDzxSFjoo/zUubibaeDv5o1rLAaltpjLzFC1h0pxVVLHwC
zLhFqcffPzwAMdSphBHCwMLcXOICZ0catZvUPeEdceSMDHMV0IoxyEvHcQlysmTy
10PMuMEMG5wuSAmwWnh2t96NoMElm6nvopfyeF2Lmfny/81YNVfQhgjDucY6JuMC
O8azibNXyiB8YG++OYKVOe0F5rvtnHXgYCP21zd+Lzbvgokm7idrDV/s4zm87b2h
62i2nJsDZbtU6QTE/rkIMLkpvVdupFYymEzYJ7U+84lLvDfpBGJJA3siokn6Vcu5
Ar38af870y4sSk42mGEYM5ZlntBZnjCQ5UGkjg53reOBYUdaB7CgoyTtlX3w2O6U
iCOgk4cxcg7LUyJnH8G+NhytGjEPJp4G01km7YSYdU0vFmNrRHiVkmCH2XR8Fu5y
1Ybwn2sGUw2R2GQG7KJzENWDPPgE8E5msw14TZqg9bLn7wnTAn4KAVbIo+D8z2VV
BMIX5t4EErPPoYIA+mnIVUSJqjLcGl4YfipteCZlRTdhjRU4k7oK1hUH6/a7rCfD
q9bibbw5+lfcxfUSHT6nD7O9k6C7La0aDWNkvD4wXA2HvxMqtirR1DtorCtQO1IT
cFLOYNB6h2qSvCsFfwM09V/JiJ8b0vQr9+DNy/DlKV2ssbjjmDBkNrnzeLVCnE40
vIrBFckjdero4jhGSU3DeYy3Vgc0cixHahn0ov5jj0kJHjsqNhsluTFYRy2wJNiz
vmo2zulraR1TFogIyAAdYIV8RQz1zZrfgsPNHm28yOnsXw0LkFa455BFAsARBA0y
Ak4c6V5F4fqOdAuW/2t9weM3jEoh9vdGXARFCGV8rZQPWfJj1cKgghiaLsXj4SjH
m85cvR+pQ6UJ38NdYUjwz2lqlSz0i86420wIzBw1y8X4gpWEbbaUNc7uupqniewU
WbLcwmduNDYUjVWSpqLi6AiEq81MMTSz44PSxMwB0M86yVLoBKFwz4RvKW2qatsT
GONpCT5vJqye26W9t54Oi79AVGXnUOZfJLuPcHFS7NP8aj4c0d/CtJT/81EMlgOb
kQUTlySY0DIVPEY5jcy2VJ+BXyrdG9aWqvYN84yXeYjF4of+QfAYmtbOzdGHhnK7
BSQFFxdsMYD/qgv9U9RW/KgjaifVZ7j/u52EHJRBL8hyawystPGvsPUv1meoEhzE
LzLgXl6uhn80hmGYkVJRuqJvaqC4zKU1cd0AkqDLpI0mozTaGUT+GUc8eGsluAot
T2pfYxsqDh812JOwS6q2w8zYWhP6R7iVem0YwiLpXkcgKE9dKRHclrk4J0fcWWLc
t8qo0UpKjXm3xYA+FCRouDplQsRtKavWula91WxZ5crIwzLGIhHX2fr0DWrkZR+x
5UVsQV9CJ43oZVYgJ150xGkI9YzX166xR2110RO5E/1pV2l8JiMWR3+XKI+7O495
RUT1ubTUzk7+I+jySo5UeMoBxO8nBkngQD7eWWPKny0Gtza6JSUZQBZB9qGDOCPu
3tH97TezcXPpDIN9GRF3usRPy3sYFmGNdqZ7iVujKebzy0X9Zs4T3Qm/dmT0/MEu
nUfS8T1Ykmdw0b5czq1lucK0O9ghQwtwQn6HyxmyOtzT3pXNBWsYosuGhE+yCqEf
PFGSXBr1+8Dx/+mQ7lx5KoKaVJYZ0LqmJaZLCG2YqL1+zMmbjzTxuRATVJlN12X3
7lCQ24+htrm4Mz/14AJACErewmmAElXc1p18mLRdHupBNBYYF5HOJTjOywB3qzQc
MbG+ALGe6pxRH38XOVWRKbPawHB85NcbPkONdqxCdjWPGjGNU4WcNIVhPKfe7IXy
k7K1uflZ1ZvDD2KFIOiS8gSSyHKDtqqN3dGotxwFrQaYTRKTvIKeHPpLBYMpvXnx
62XZAtCTmLgTaFhuaJUwHarR6gi1FO+QDsGpCKTYzJe1FT92xOvEGoMK83Dv4bJB
7JCB2cS2s6+BTx+EnCZWBaUaUr+VcX1iUxn8xHKEFiGepHJKaUIsbgPdVyTxuM3G
c2v9rrIPQkynvMxfEKWogvnzeh0BFC6X82nu5nf+EoB6jfqOJ9Ukdw2/1xydogYB
EOG/0IuJmVKNh5NcoKFKhLnucFOMWvMjJII03s+hxCUFVFqKuLscQc17FVvy8Bg3
h9+wGbfY4d4GS9ppIdvCwWNH8YdCmFzPGATDBjqenwymCLZYBXoFF4uwsjjAVAgA
0jmjVezeaypuMX/J68Trg2sKCWvlTGVa4pNo2PQ5OFFroKsAwsqHYO5YOZY4urw8
e6GCym97euHdK6QGToBSuQ5v2zYzWmoz45ZRCufENONFBtFUDAclnsQ3BV9f2v5u
lKsNSzijkNmR3vw9uZ+r+uNEDTR4aiMiyOsB9zxhYsJEHVkpLI043Zib47IAHmZC
1yCCZ9nG0wUDXfAkSzC5jKs69nkDBxWvSEgVZdiDICPAbW/Rq/AkeecJSPpoAI2F
7if2zyf8umyd8DusCHfpLkYGtGpj+jQqV96fOU0/XFIGLuz2SpFgiRpRciMCEqCF
KsHCUOOq08krXh8WcR5KaK9UKp9WDpw/IlYDinvNX1qcVjOdnsmAli7sNjNmzsWo
1p3Y53YP6xaz/H/sbyjZnw1ANwsaaHFgei+nKkGgEOCOu+/54kdJ+nEkVRfUQdbC
TXfnwpGL4p6SDqU5I/AHQ9/jSxmKg1NkTr7lpXRV11uYZxDL0THWek+eV3p0BGpD
c3Tg3MYmfzXZ+mzrZweYZthtSDnuUz4JJWX8GJhl4QC8e/rHb3C1JlMVVPCcoJ9Z
GCFj0RWPJkXPdVp8fUSPoe4guDFk5iawjl911ooLmaup1iamxIS7Xv6VecWZE+/F
hWIsgmF1nMZzoVND7uLQGw6OtqXePFV1w7XrvR7tGVmlALI6m6SeselrPPex4UxJ
KKiZ/4CQqHTNl0r/6cMQQXVKhKbC8ngNjITfy/gR8I08zvgeii/tS6/ER/v4i2qe
x18o3PjyYKj+c2ZHKMxkjaIvBMwngKWTV7HOGZvOo/Re/OxOXm85BdMJFdGGdhxM
7jasaLCL4dlLqPCDlcd11TiS6PH6prSvMnV/Lvezv4uK3JEeVJKteGBwzcV3inGK
JI2vj/O3bBRz0/eVuhkCLV7QgktV0oSsqtBAN4+KZcqB0KroFrRb7YCzbdnAvfAm
rTsYrg+zoOI3dGikOGSrYxYgsaWK4KN3ETAys95wc8zsod9Ol5QyAdmJv1HUadGg
zTtFamfzKiS7ljtZ4cnrfzHNMagRh9XL9UezRriPnh7bHBdu1Nrpio5J1scHi3Q4
CubQZy5pkoO1oZuhYfEPG5UWk+C0M9v6nZwI7wYFwSyNHyBKM5eMkHm9b9DbwkA7
ybbnEb7uk0tNqjIed3I/NO0vavaudQj7eM5o6lXn3fmcmv7tAgq8TbiF6daTcFVZ
5CU37jzud+OxqdCwHItgLeNMXgNBILgigMC4V3+lO6YheSz3IZtYhqhsrX3d8oBb
R3lGPqLBa0MW9K4bGG+KaHfv50FwYwJv5rY+LJSNqkwXZ2zl9lsrFIn7IsVvIkVS
UmN3JMwW+3QUaqNjkOQsSRw61hEL5/EMvqMJba/daNQjT1XtNuzyyxBcl9Bza2aD
uXtHXXuiHC8/1zFKQwBmJWvmVfAQCTrwcbJEmAFCTaxp9DeQ1Q+gkyoet7XCbX2h
WwCfZ/9SzfK25GFTdEdgA21eq6TnSNkj9K6/CgNHnmprPJScdmIrri/nC+Jt1X/U
j6500BF1tqFkO0r/S6T1fYbuJokgcdcxmGtlVx5HgBBNOHxLuqoTBzEeeK2GYZPl
1v1VjCGBtmZ9oJ/VvXeb+0nMCO1Qbba8qr+uKWDqgJ8t2oxrfi1MB7rgXTvUMOtG
utlsCB7W6WZ7jILza9MUt04Hm3YXkce+4Wed5f4Ysd2r0zQ95lZQB5+KFZrVCFBN
jWTi8opHAB2nWgGeoVg9smC3Db2plEfQh7PGRSzfJ20YHN1J6TC5r3MBWJljzq99
u1kUBLrfTbVc7zrHdzzszyGE2i5jr8WxReIcANOmK5SsYgzdFymNUVc/Pnesud0Z
X8SF3KkJoRNxDpLVYPRn7/7zj1BW6vqv+LJrc4Wrcif1RB5o3BTTFUjVZyRyvHGq
F0o01fDkYTth7BFLxACqY4DN/wAhI2cr83H+XlEDt+xzRvguDZeMAy3GrhiwR+vu
Ctmr4nT6nWBfxnMzTqDCspsCAh6zmSpal1E8RfcAaNfrMpDcs+PwiQWfZwq/L1Wl
y3NSwtup+4Q1QYmJrTHgKej1W6YK/ixn5OuAvwjT8NPZ2uGFqFZ0h9x9/Om/yOtv
QL1agX3xGdfm2mkXZ4cSoEP25M9jTKFiR+WKzEZFmYx3MNNsOZObxdPSQRwzJ8d7
w3nw5XWZR3zGwrVW9zeNwXcspZ+J9SCRd9HojFuHR6/Hj25m3QaXFO1eLEjrUWDF
AULW1rfMgcoBrybYQS15IFCgKWbn9qp7DCXN3UfawIDF3430oh3HKeZxuEXasNMb
Pjz1ZCa1lxgIXoF7m2eab+uk2bigQtrFytPlCYx6kddTIZNVdj4ZlofZdnX0PUR9
lyw0QzlLf6pMs9VQUCF2hLULrLBSt0g7FKL2OYifUF2HaANKX5TPJ25KU/i2SRh+
x91jpte/oPA0fbJbVHHZnWG5dm8glo769DTdkswN8BeXOmQx0rUEY7pxRCLFnQZ9
Fmw03pMcmG/2XH8eUmOBxSECjtN6qgUESrAgQEuRQrJ1miehRjfQhByXe1y4uPDc
ia+KeDeANM/yyL8NWp8Tn2yrDB3zDw2LkNuzVrt9CA9p18iBXmI3r46KY0Yhc4tw
r/xwssmtSIjEVrwQygwfcC/9bhGTQV8CzkLoDE4j2zh+EAGcXKLppXq4EFAPGkaa
XwAiu4foYT8ZL5U6D4zJ4uKvEJr6Sn4JvdUh5MuyAlKoR0esNONifZwNAM1IHejK
ULG84O5mvWcGapr5erUU+qYVtvyA1KCC9DmzWlZaqdkkCLNaArDQSR25IC7vzgKi
1/6qFPWi0twsGFMLTg2vdfnYt9qBx4ucMiq1x7G/fSYUuM4g7iAiSjNiovRiDh6V
kYOrsuoq+7Vyw0fWhLBIOTLPuD5RTnBU/YxsJ/r5SX8H1mKxw7nVTCTnvcb9tE5U
KealbpwOB6nKknyTE54IL0+JDbwWPuzdsdbG8MwPKvPTyf9JR7hN3sb+9vMoQNoM
lCg+Hl1rIPAASqsUu2H5QnGX6iLEEsSWfd236hsxSzigbWSfmYHnPGIYCnpEFmsi
6DGnnsCb5qo5o3CRExhW541bXWEmlK9kWYgPUT9EZn0NnIYGZGBdOTiE+WNyH7Lj
CTQvvNE3EavT1fqlUkBhEZzYWcFxmCwq2D+nr9X9T9rA7qcMqilWWap+1G5cCIKH
1Pp36dCq+aSLmnq9X5jZPL7rgKNcumX6rZfr4bi6v9pzZ0YqmYFKg5ZIOBwbACRl
FlGAl5xVKNbh/lSI1nulhaBZwnJ7trxY6/xHlWcah0oEay6mKlo4dLN6LE7HVNhX
olTwa+RbYESWVRxNNUtAp6rvLZW9g1hPqRSo2v5Kluj0K4jaJ0iq4e7Lcu+4D3iT
TX7Q3f+PsaQ2BZTgepVa/EY1NfFHKOBJCK5ZvHboeuxOZUulgSE/GX0fL5zuBV4Q
4SuQvwQDluMCPFpR1K0X5TIaood9u0igbD2rc3nu/ggJ706gGim3gOX+iEXJposS
PrbZCB5WmXvoPEGdxCd/wW3GmvMwZyKsRvlY1yeLc/RgFsqcvKHgdOX5lvk3c3au
G3JTzfo2aTh7FZCU6EYX31o3maGZ9sx3Wd06rM4WEBMBbVHyw3P+5irG53TTXeAz
WCenUIukrQyM4iUooBjBOxSBxVGMgOA1my59kIiDyLS42RXGCeTwGvoTgdxhVA1b
hvPtLl331sgC1QOT/QPgiV4Bdi25Njko/uJRRDP4sL46BrpdSICrMsfQ3UEUMJmg
7oT57G3RPHU19pjbyNIUy2lmmf7PlnEArjuI7ecKJ/XTr6WAe6K5UzrS5GklVG8P
9vA4wZIsEdjiZFtG9s7BCHpQvpQdyOnv+zlJzINFgl55KPTxfQ/bpJrFp6dPZWUg
yWCzbn9sp/PVbsnmipcXmBP7PPGfAVlVWKrPE+rZeGE4qFKrtX0HrbsniECFWmZm
FLFkIo3aX+9CWkuPbqpVhR2/ueEblt335Mi+kbBXAAC9WlNjP5YwY7rv0FFla8Rd
d2xsGXWGZP+RkLjlqyOW8b6m9a13eebqSnxksxGEXjU5UMwXlfvQuSex3MS6jxxS
0pfECunETlwC/OvgzA1y3kcQaBuRw+XNqpqvFhKXxJNhsGDoicpRoa+1akR6qdva
wcD/w3yGByaeTsgKklbx5ned6/kizRk1hn8HByse2/83Spznk3adXEiITAAnCLjb
vCHD2VL0wwzhdn/KNYQJIZvU3YO8sbT/tdNB7e/xOL/2pZLu1Y5DNay/gMIF0SVy
nM5fN6T9uqlS+IIv09/sbzfzivggrW8KHrGBfU3CctElYK6Vcq3/6vUMSvw6FaiT
8Ej+SYp7F9cROT9lYCuaLA5ULWs3rM2WJY+A1djNce1VtlCo3l+Z9FI2Lvp6ezzz
OOOrWcYNttpC/2rXFqqT6c88xkSRvbU6Hz81ESsh1lgyTY5+efZb3BeY45w28c1x
+a4txxskWX1Rlvhpmyvi98tnYPKxE/Uh3EQyB2bGhnxN7uqVW5dGIUi4G/TuifXD
yjisrm8xM7w+Y81y5/Au8/YpBfKA+RymsGjZV2g4vyuv5qSsIptkDSHuLV6yka/0
bZXtkdAqDDjTj9CQSNLGy77x0VI7aw18icCIx2MM4cEXN75pibSNhlD+Z0YeSl15
6OYc9/SaoCF38x7foxhOgVwhygTR/+CVvgIyLiKo2k9Y79y+oZ/ZkDkc7jKH87Xr
IC+fWP3QpxlwrnU6N2uM4GIFat7mwUlCm/dexf4rV7e+GG0KGFsHbFixAr5eiDCv
wcVBb9vaa/nTHGOakF00R0Z0pOoU/3cx6cCc+Bq2tAdpK2cDnl8Xnvh+o5NG8mCy
qxBUZGmX2A9wkFSCws9buQ2f7lpwieC4tJWF4d4+gXQpuAeAEmiwMSy0cXWQUiBd
DVhbvyLCI70Jx9izAClVBUrptX978KW8jN2SkWJ+TVi1NcruNLOgSnuWQ5ZZ98tP
kzLkiNo7N3XT5RKZ5HpkTvqK4ZmQxI7Wdj91LTCjfgIItPLEKhkH3G4bb34zYBmw
cCDxsFRUg1DYoZu3NCilRJsTfw0oSOL5rjL3eD7OZfH07dApqZa43zpQmX7HPhzj
3dUJULhEDPS2A/vqc2Pse5WuEfb3/IAGRSbP9quUZ6s1M2CEC6jpOo4Z8R67QAf8
hXq3w+XCbzKKAh9I2LLxmToW0Qmp6OpjKreSQ7zsjGFDS8Ou9E2Ue1ANmKuZ66n8
Kvc8MqZHVC0h1PSieL/T3ZaaM7RN8e1hrkuxbbE+ODepC/Yhcun0ZBXl+XfnFMzM
IvcCWEKKrawjyy+94S5VWsf7r0jV6vFUfCa+T4Gam7gRKKeemd9o7sP3XCwdjCQm
US3fUAm7gV8abQZXl53yGoBH+yrjNo0rYk9HNCtK+7hcBFxiACd2D1risilC38xw
vfOrZIyZQb0Ff1mFDT7AznI0FYLxNv1ujAUaVcehJG8Wu3HtPeIHPDepJvRHANjG
GYZcNZzICaalRx3PrAilpeDdZmzE29+Nx9k24qGlxIceyaAOsVvDXhQybhywzu7W
9cXXApF4AQFlufRJOp5I/J2CHF9o1AAY6yz4AlNkyU1xApWl3rks3cdnDRGQclGd
KU0Sq27ShwidlmLgmasm4a6Qp7bXSNkQtTTylchA1Z8eKOyNYnRM/O+S9nwWHGBY
Hu98IsaqTs71dFGsUhuGOkFyPqa+mC1TlFaw+hzuAzZLqyaeB1nmh76VJUY/kGUT
7bEvmX7P1m1WGV95JbMu/f4qWY9643usVwXt4YHZAMyEocHlABGMdfK1nsjF4aOa
F9cRDKb6bxb/v4TX8B+cqX0c2ac55VR+hutZXdaH6UPHigTO+CMXkuT2Ik7klnCG
0QL6JG4u++XKWoIV+19m/DMwE+9GgCnQoXrFmhWQMWuaQmvw2m3aL9mqYbbvUyC2
IdZt/DpdIW72Rjml380naI8WYKehwpiVaeqcYv9FclfChviYsjJQNjoMsULMzV2/
snCiwtKJrhl5WWr2Kfutq5I+m7GST90Ji9LR8v8sIJhBNsmdIHUM0AHaZ91jtMrw
Agkeq+7dI55wxLNBMy8lVR+fF/EnDskDRDkr2AJiXfirYtCjDBoJNESclPa66vJC
dvcXRV+/WXWXQe4sz7ztnZD+VYYuaj1r/FN0e0obw+9kgH2zNSzfxNPQZ6GdK/F/
qL9/Nv0tAf+743buh3CFC7tOU00y5CoVaAKPHovD7Xn3nme7wWITYtseV6l/OKmt
tQqrOdrliQeOfJz0RnDuKsqTwEox7TpNRIfRstoa/Jo7rIkaKSvCcZ8yAvoIg9p3
wK/kwyLfN/X48VgFtEe4XAug5iGjJSrvMh478zA3RybjzbONttqt0zr6PK/ec23+
5KQoPRNrXCeBhverN4f1c7woeuVm0/rleRmTeZoIleZvPYNzKZSEqpCi2QLFjItD
3r8B6cGmA0A7UQJXtlUnSvFDMCKPcM8xJxoUrHlNS4UBIjrqpod12rEDG3KTaTF8
M7lVOx8Lqh2piovPwpbL7gOetaGXUXBFlOhgfizPVt8eLxJtYM+vR52jkiz+cl+g
rBj5aqXeQT3GAvNOCgpoY/9eHcnJgkAddowUX0fYROQ1XrQA5b0aNIG77rHe8Hjv
kD/Kl6D++XIZBGUb6F6nP8Sp2wX4RTXnqEBi1hWSo5Kk9SKRjSf8/yXfG56dB43S
06Tg294KCF6y8xNVfeEt53LTSREpOAs9bNMaZAKTyKz4EKGgFOmmkZOqtWHJ9ckw
ixHeRLn4nqunTjmUyAuR/lt27o2VOo5qTiuvZl6EGJkD8VFsNQMyqVzmcI6i4fPo
f+47ds8VOQZlVaVjrQ0W7cytMuf6+0BUu4GZrEoBbYKrtb5ZcpS8leW/S4Jnanjv
g0L6KLHOdNtIFbFqVAuNr/+m+PPy8Z8gc29kft9YXCC6/pP8fBfJjxmYiWK1DkXa
bTRbr5zZ6f3Z+2AkIajRoaO5e8ZlvwP5kaTiWqEi+Ycs0URe9W+3vF9vC5dmlskf
AaPqS0EBoDKqozPfZFPtizGcLFgnyuVe5BdF0K619/efqjW+LSra604nzEGkHQOA
4KGLSXKJlmWT1frTznM/KXTQDiW+52kKS1knGn/whK4pRFzKXJXYVi2ND8Lh8gUv
DMAQKD+QOOFAAL9dKLtXDS7F9blLZHiaoS0ltZ7Bwl1tYghY1Sxk5Gv5qK8/JAvN
6j5PInU3xrE+msOz8WUGVDcYOieHBzDrih5MTftE3uwdUVQABGvI4K1gs60j40SV
47LSwv0RxcCiObCMQmmugZWcDK8uJCmlUhdVGosv7uC6WXH7KNiQulqKoBKCpvx7
jEIvVDXiZjJIajKOPKJK6E0Ij2qYouM//EhL3Of5REUhVlSxxSu2+x477qGSERpk
kSvcJ8OS6rbz3zoulqFndnU94PKHo09Bu7PHtle7Un7+HS3W+MAqW8XIjParoKnp
jKLKHmMqay0TkyDSoG/vKJAp0ZaHfiq53TY3UJdy88u8GkJ28NSyLbFVpMsayn10
8tHozFsxum+IfC3z+LT4nQlh+F/MqPzkvZB+UNOZSU1kJ2mn3K0JXyKV7jgQVwWC
8dSc0muKVapQBkvLg+3KinbQpTw0w4TT1VSoYdy9nTE9HtoCqFxViGlsGDAH+mXT
K33Lb2vAbfA636PByKm4l9MFpKphe+iLwj6T/OQxkbEuLf4ZMMHRbar2HWF43nv7
I/uwPGjsZiKRvrjpcGTMGbwKwhKgMro6KbK4heFPOraO+1ZNsdFPUQsGAjpwk0F7
Y8vHVsJw54tfKqUB8Di/cRp9jGWOc4kqhKzIseBMigBOvOdSWi/FvXGHgaCaUZrj
uc9+uDIOLvYtp56qwgBBhuYb5CQwbnxTUpovE54/mAYZVvYpsjKXlmaD5IAmJSUr
/nR7/ifYHjnzeehhAl3wPXyuwElW2ukspVrp6+LinqNCt0UpFHGZT3wyM3X1L7NT
3fke7DHodaGnODoOnHq4q6L/uGb6MhGmd+eWitJmGvw5/k6fgtr2DMDglEy/7uFd
T5rbjId5hsQDT3pCwkkNdsTYs01tiYF9F4n/DWk5Wx4kf9YHzfe7CiXI7WjydD3z
n7BRdG6Nm+WNZmZ+8bSpl8DepFWIK/3FwxH7A8i0EdrQbUuJVendFCvlGRv0YBux
MNTGY3nWWrl+dWJFrucf0aUt5qQwlFz5n+TjO5cWi+woi0OIE1/AnrCFkqvhBD8Y
lz8LXnSTnE8gEsXNPHX5aBeA4dOY7ZTEsdKnrRNF832CDXYs/JOuBaLRznoswDM4
FW6xPZ6ScmUT9JiZTfvqsttPTSC0hkiYq77mAaOy+bZgu995cel7Ah7dWq/Cvn8o
VgAEhQziDiCg3oxEgkP1wMYyTxIYNw60SybzFCce5VWrCGKfBEXgcbj4Za927Zz5
1HUOae36BGnLvPHoWWzN805E6o3XmHQdjcGvAGUDh805NtwKeN7N1mgKwLFfiNAT
Ah0H4BZa3oolXkPbxUR8BPNt98puizRIdgYpLpCpPIE01MbB1V1+iNQ71hHF+w1h
TE15RWiz2EQf+GgLLqvWqGTHFC4vOuEZXtTtxeZoG8NwTWKFDIY0j4s/sjxnmC1r
Ho4FM5xGaTWyT625cCqZyAf50MnrS2RU9feJL6Co9KqQuCzZQkbSOTlW4oLAlJG4
ldPLvLthJiAI2LjCJ7MR6m8JF/iymLTc02GIrmyUl4gwZhm5wCeM/grDWCtrg8fA
fo7gJefD3lUCixzUy8mnudHCYgQbHkxOW4p+EL+gNpEMtRfSNcuff7tnMbdeQXfG
zAegtlFJ0lbkoDh3cFHoTdJi56wSOLipMkhvkcT2HXXzMOmghNbozE3YLNBrRQw7
I05FRjFHiVe5leq5h5Hp4ZQMLQFg9cW7FCaL0edR/VrdLvPemXDtPmzwguorpeCy
JL7CQRGpscRFqvfRuswKhKRYkbB/tAAFxE/FWFrUDxYXOH3vNXmkHTdNj+HnNvAl
7bU0WCFbvUsVhRCLGa8EM2X+V6jrctqvG0OdLetVTRnFCr5Gl1bDJI3l474ZKdW1
iVr0pQUJBiIhsYiEJf/aACI0u3J72K1YMBbFg5KPSP/171ovFhqCWYZYT2E1V9Rf
ipOwuaw7GAvU2NQJwiuqQ7RptdiUN9GepO234b+uxGCo6MB435r2I0HNQ5Xsu4Kp
W0p9qkLQPCEsBzyK4hXEKu/ovKZsv8eILvIIKdeND5Zm7S36JxH7FPiRjmZRt/SS
Cgr1CJxVOdK6PaLYnN9RCLnoYnUVLpMvbZl9CN1ybs+CARYuXu8Ylb+txjOpCt/Z
zJfbi5Y7XVx6y3vLgucQP5cfK7OIQOw3aDCMhfWhry6OvxfDXLH/bW2k2Mw6kKnb
hPoPZyuV0fCMLnfqzSfZJVv8GrMF3wQYKr68JV1yyEEa1IjXAuetpfDgnXoX6cVQ
kzJaGzsrJg9IRfAeX9ZAUEr4lgz/8YEj80L7+/HytITc93sYYfvxmphGv/oBrQPq
PbVXREbBHH7QBRBVcoqnYVzUYzoOYj3iWMmsswYxBecUMsLLucjtA9phyRgk+Sz/
vTszJcW2kHBlG14nqfv3A6w6NCcTnqUDs/j78VwWq8dfNfXPfn3RnveglL9kflS5
R8JNNWz1Oc3XDbIjIYW+LsCiXckdBpX7lDou1eS5wsa8LEkaT8WWceQSY5MAUhZH
zD0Ae4GRWlU2DIX8vjJlSWbqHeJ33nvZA2gfi/Znug8jrYMBSfZCZe9iMZBi86og
zgvVA4yBB4QPlWbzAV9JCU9a0ycpgxwnXUUyYG8W9XeaxEtKezui0ubNbCbBSSbg
XTdp8tlDTOUR6e86pDsqiiYZXn0LwsqW6FA/XeePPv6zbybnzq+AwrsaBZmnMX6v
76Yeg5UqkE1o76kOrdyUrf3b/cf7+el6uSf3RCPKlpJMisjTQyiKBSaWDvWwN9lU
m6723xnuqnN7pxvZ0HQSGysANneT2VV6IowAbVi+9OtHoCspv3JSJYHT2KjGDKq2
IRMmj26+aXzdcFafhP3VYUknI0SxUtgSrqljeRFEceKmwDw9X/e5xzqoqf3oZAYF
zMf/QQ3t5np6HRh08LVAz5dBNa8iaWERsTOFqdO70+fEClMl2G5F7KguOsoehYiT
2Fqd0md7+qif0tNDCT4ocJltyGFhvCBrIPjefBMf+5KqVbJTcQiAkvl2ABQpyEkP
Ge/J3LvFMZ4chxAvEtQK5kNwlQ/ftTfvpRIo9lw0CgEdzONmqxaNcbxPEiruSIWt
3/tu0IFQy9nJOa3u+xPlYPSjjkDsPeBuhB+OcT/gloKcqzIUA23EeInJyq98dONz
xrsLE0CDUJDWcWOjuENl8ASO54mDWl70LybOmUunztb+DYLezv6GH3jE6cFXOjGy
G8BxmlNA8LvxEcjJCWVr8Vo/n+oU6EMuglLB6aH93v7fw1y1VDPzdy64smX4bdzT
I656cR9eprvX+HSWITXbttXjWo3LYKRkqj6q2dIpJyvqcg6RwTmBNbp0SwevSB9A
eheneAj6EyaWwLoG2kCt7NWGJ0fDTPfy+g0rGNWJK0+JlV9tx8HhTirSGAEdTdno
5RRyly+eZlk9CH6J2kEcBZC430V77fbdEGLCkRT8NPbJNXrHVfZQvp5iK5T5dzus
MhCVlMdQte1mN+0OFaNtTezthiH7skt/fIbvBAL/WY78khnu4kNUT+ZcFDFot92d
7qMdCmb1ZLMszDa4BYDrXKSXa8QSmObr4asN+HOyzJtqoDknbKvkOMX0f//oEtH7
rq/eFZD1raz7YfB6WhlFwdeTmhGec+J7IEv+fjDY9dE0S/YfwO3E+gqA/p1oxUdf
BquQHhGr5uNj4iKYi1CSvR630D/QFgRLtX/JDYB9CtI564V6qN1YQiCtQ02JJzgY
nfYmvvzTESREEQab9r8B1M9g0bTc2es21ZQeEmbixwsIB/2OVoQi8rC6G9mHb4mN
v1zMSjaUBkCibjHD5HiRxMUSMveRd1ztrT56TOSxvf3yP8yyLAw/I+fKTvVc0cMZ
BL8wQcZMydkioNLDeVmZ3mfRCGYD3wUtkBoN6jYx5QXbtygp6TmxInkR17n8hrmF
ZIdDmz6I54QIulYtVYnWgZJVNe+wITQLOCR1Z7AsPJvU2G3uckHxfFnVw4y/zjSY
cl/NzrfYgUdCQIxK5/TTBo3AouUwVtWaUyYJu0Rk6a8XV7aSDAFB5g+0UmP+TuQh
nr8ix7hUy6ZAjyYo+SMLdAHjrKryrQNgwq/QO61zXS411vWG64Hmt+eDChKnBhnu
8QfKoNba78oN9QiVvvGZCoertcH5hp9U2EZS2XQ70gfDDQaII0ty4GbzReRNzhVc
ddaWjwNYiLy/7wghFnMu8NU6NVbLo9W5dO8aqCRohw+HQWOaKe+nlUh4COsBF+So
NSESKB3IUzqn5xh46CAt4vr/D+r17tMmt77Gkwh/SCRiCCW4N0CR4MjREeynry9R
i+DOgdqJ3xLA90hUkIAZXBYExkNFuWlnSjgiLoTg6pXIvFMuEPc63Gkc9DmCRGlu
MknV4tdeuaShsTl4No9jMYh9nTLxxEDeSTDcTxDJ2pcuHuBIikn7iw5QJCiLIF2c
L2pbzcSfDeb77Sw0J7McnaSV7czsMJ5p+4fdr/QM7s1QjhCYU6GIV8OY/MFrFlBh
fPVSPj7z+yelGYzFlpdCQdSZkVrysn7ZNDT23LYkOGiz2WkVyqi7MHxwYB2MY3yA
Ia3Nj5btYbw8mXI7EcpZR7eui1KNVQy+ESEKswgMzhw4L4lLLkKRJ+6RyxaMSOU2
lE87X5ahoei5Mvw7WSWhiZ3nWL9AQf79aJ01glyVDJGpTvGgWFqHnRKcw9TTM80t
brQTOCmdiD38OQ+NKevOpBXDoQEw4+u4Gs5+8B0AbuukVfMdccL2L2c+MxI0Llrk
SnvhhT7m9hF4xWmI9IfoF+UzqfGTj0XEWpuxONBYgkD52xYPHY4Ow6cicYIaJd6K
3VOCtsAsVevIEKkoLzORyieMxVC7WpWiaKwE3EiYJ203F8fuTAU6P4Ceh7ORrHbz
j1dkETNu1nV+BZKeML9IvxwIS+dWTVh4/rXJ3r8z483LouvIYpfybtEblHWlQKOA
swhTMFUOmb+yEhv+kaNEMjuuglkNVMMQzP4k1K5sSLx/iNsMcNtv7yV7nFMMMYAx
q/Ph1XfcihRddKJzb8l/tpJus7QWg9ADQPSX3ngrrjyFrjBuNH1TlRMf5TNXL3G5
9It3xsU8EQOjpi2LgPXsraPITOND7Xcnx2BUgF+A2Xcg207HXqI6XzirOoaRMg8X
yrwmh72bMySb9+xhre08U6FFs+kuqrx4W7pIhf9v0Ih+HSI66+6kN/5BhpwU4ZF7
Mpk8S+mvcoMJr5r/8jvrdJeDquvAHS2WFxXweejUEhPIPUVXEpqBmt9UL+upVvco
F/Tb/T5Ou5h4AVNiGAE2qnqewWZvmPuQishjNId2+B5Jms6F0G7+EKmzRFD5+IzM
qN75kNdYRdsx8uoCdHT3IHquBVkiCn32GXksAdeJHYvNXavSSYMDg0VcWV5hYpgK
inI+NgpqPvH70WFcCj1xg9I81rWH59fxjBzsTcodpFqz7si58EPSE5c0GPRFq9n/
+xGPfAm8FfjP8HrES/9/EHYArAaT0/NfOskkcrK+E73owCP4EsItjyflOxTsBTu3
JCAkqVjZ17GlyUbl83xZbAv3u0eGQIV8mEjNvJ3b+grjqCmOnBvX8GqqsYNBUmg3
yZnyA6MhCn3JezDUI2ZKKKLoIgd3G7nZlbmdTqJ8SQfsThh7ByzRUmguaVSCigTj
eK/ffEFy7Ofr8i/fdSH2U/T8yLA7TYlayk11NSGD01Bw+sboKImOOpxu4dqfaLEq
Pl/Iec7STomYxDZ1+Trpui5Bgu5vMZxIJMEPclOKspvlm0CUgaTpJkBZDsb0vxkK
UkaqaDrykMyViQpPaMIY3oBns1CSufalkzMCsBLVGjYKrumicCRUs+pyeDwF3hnZ
NzEZgl9esm1WNEXiB/sskhK98CvzygdF49kcwoBWz/kMV0A3LSh+A7coTHXfh28s
gUadyhnqbq4AAK5ElHxsJhY9TCykZ4/j3Sdm8huK/9C8SClYU++hEnQxOv47y5SX
SbOHt+ySSm8ex/hNrvUJyNxm4m+C4lmnJ1t9F3NCW1P6q4VTmVuvY1ui3wfduEcr
nDljmbAm/lRxoqZovU8nIux9Lds3sV/QP6BZLDNpZFgSZby1tmek0vXPeD8KXJ2X
pInTTKDfqdjYjaG6gsuTDJT0DRY91SwuEbOTzpltoMWCkXz18PVo/Xd5Hd+/uVwz
Xp4Cgli423AdXqaIL2R4MLkLGFuDx8AEGXOfN3RTc2Z5c4Qui863oUMHfslzGZfT
Rq9TlUG4HOUSRgLQ2f+HXL0uBzgRQ9R8AhNgAM2SphekaOda+W4XbGdP8ETox1wo
Ie4XsoA1DT+gM0O5k4EWvV/MPoV8wzR3OVyeX/HjcEEdOUvfURcgx01TaJq77PqG
KKYAEynCn+Yp4scDE1kPWgH1Cv2xU/FVJ9a5O7SSjvu3BXVOekfFyHxZmCHp9Zr7
zKCxBkvSWjMOAlYt3fXwTymTHlzLyt3AGoN1TKJhnA+hlCIUs+u9skHoR2YL+unH
Ly7YwvkyDm5m7s2FRxdv+oOcIIp+PKKbuUm9E1CS93fxFQsdPrJQUSlFu5ddmjE8
QkDu08De5J9lCjPgrk3pEbcUfUvn4VFWRr0mv01wt1NJfeTTrIzd8Kwah91XIr+Z
Y4cJkZ6j+79HmxUDfmsy4wrUw7ZOxMImyScm/lOFwj+r1SzNVr/zTqq2wIgLP9VO
Cvn1rtojXESY0mWOWhSB7cmL5GoAX/MZBLxqW5KMqMKn8mjlminuTRmOrvBrR9xz
HcyLf9folMhWzjnr8XTY2VWb/K5zfemv1FyVsxLpn74qjf+2T5e6kWaCUAl8zSvk
hwEvUV8V2GrBN9COHNJ65boe0rRxFne3duMFu6BrxYe1f8bmDAgURRsQZlFl4Ij7
HGQlI1PlM+ZQKrLHZClN1zy0adDpeXCI7Leq45ZwhyJctr7zMrOaVxr4L6uVSPy7
IJqje7UDnbCA5k9wyojhOeO/oLIANoNXPdI0gPvep9H5WWPoYmdLm08RolF075vM
tith/ihVuZuOOHjbGmzvgNtlXiIQMIGNQY/9EgdjENz/Bfo4vCDzqeKTUj56t8Ll
bxGZumLvd0jVcWT4TCDmMa56EWo0V1ZHDQpjc078d3fg9gw45rNHvBX07ztrAA2b
NENhPdr+HuqRB7VMIaz0Qe+pJ0nOr6ndPPGbnc7ekxGCTN3+HP6GUO55MtspkyYh
0JNrEhlFqRy/sBsMtcgnx3hmImkpHNMGb/O2Qit1GMgwAFuWTcq/9T3Lh27dVSCe
6qdD5iGxw1VOyIktGkBxLhYcmWkqDv1qL+PZR2KAvdfGFZ2WQpaLZeKgyucEgJY3
dCu8BWMF8Hp0HOZKFOiLj4o1pUaujZ+cWX2ixnXoGMG59PZpV3fBavsbTX0y+03T
zG5bIT72BRAps9wzdNjYPcrbvbDhEmoTpVK+MqH5aFvA9NhjOVCIN7lCcJgHQSGF
Pz3kOHZ16YpoprQ43oB0ncE2pojXxDrsOolskgxXPY/py5iO/W+m908dghdC+teJ
foRptRtP8nl5YpjtvE1uTmmP25y7vlQ7yLIjIFRN8iTOJdb0myguFrsvgUXlg9La
uGkGKcVfjeR0+15ycciJZhICwEL+lJkcsikVUjmvuTXa3A0Pe+sNLpqXK76BT8+T
dIli1Ykeo96BheghkOds9kD867yB8OsV98tvJEOLrGXeMhY27jY5u8uXRC9R6O3y
GBmXh/GMAp8ktuS1zPoEDGuqeVNLUOR8ljLFzjL/dnnDdoAJaVswEaMdGpZEiYA+
jMCBIRrMbYb8/Jt2qQwyVZtrX3IoaEJl3GItRbad0nN35OIPA388NlryuNbRtzFQ
fP5OfC0SYRXPgowYxsLAcwvfzwqivjSc11fsfRP0StoA56yMHg4yOen37L6chi16
nLd+7bzx1Ijuu1xG9DvV5i+UoSWOwMsYFnvNXlfLWpjIadbQct7YUcA3qbAPd5ey
Q368NTt7riJEqNTxKH175bp1rHPdmE8lOQPD/mm8PWZMXgMJOcS3uuIxAgs5Fm6/
WUGGrZz20Cnu2FxfR/ddOTQwMORK7QqsKmW9w2+KVf3U5xIn7Al0LSQyNBXt0HNa
sYG22Pp3F7bGGISiFwSa+JD9KGJOfLcb5r9H/1KbcEWeDoJY+/lUdI9W/SMnC4f4
hnNod0Y3tPeZ2BRdx221rJtFoKV6q54b48nXUKFbtowyrpYCkkCUQgby4N/wV8z9
bvzWmp3zviKa1CsDDVyy7NICe558oPdS6yJa+3XJ7x0FISDyZKjhNgNxuMOAT5bm
0BVJcgUBw00RPx3cUOUGxX9dxmG8hCPOGhpf3PM3gFJeXqT+jqXFoNQlU0VcEDv9
F64+oMETjm/0XEzBk2CPYNcH23LHLjxI46NBHz/Yldb5D9S9iRiT2DjIhds9oEe7
sm8cWzFEh7yHTyimPSblDCIKV3tnHuu2FdRmBHY89Sg+JOtWCQ9X0DJgRAByxr/9
LqbN4YcCNfUY3C8FVQGDP5yvL0lCGiwgqnLaIrR8PRDjDIecuqY+C6bjBPGBuKG4
+7w5SpEyKC0IO4qXaIPoSK9ehXGebRB12johFblLjk47eH2j6DAixrjrdUZT8SOv
1wBUNVg6ZcOtZ6fA9bfsd5k1En4WiWDqbyIxVTpIZyS6ZoXQvg0YGRop+EkEtw/1
kWIfdFYTM7Dyg0DLnWZLY/rjDCgTrpn+6B40+kOtnPo6C5HRQD0lWt+jIsO6o3lk
1wqeVxMEmydE8MdzYHzImRfegt1EfGg9S7igzf0cLHKSw7ikGtP7hvnADK/LUwt2
zETystwlzODXKknn9/H6y3I4trePbftKzuRBvroHNnJjpcATQZbtfqeo+FsYnVnf
9+huqKShzwO/Dn+qq5qKS40nuD2a0M7zGwROuvZXPn3Xel5k/S0/ldyZEVf70FN7
7X1ezKiO0VavcW4/XFgPCR4GKaGxsYkG4vdom1SRwl7m3aK8h/YNlF5VpnEGACQM
3+rarkg+uK6NIABm8gH26yr/d71Byjf7Ff22+VAfvlYwvG+KZRbcfzCmawCZEtnP
DdUrjoPyovTwPlSHQf0Wt4m6cZ40OxQOx6gSju1xdQV3DHo8KMUKemDm9CkeA0Wp
VRX28owU+3WjW39Mh6TI3zJ9y/gJLP8uygIUGm0wSkVNC7Vsz0SGyuk9u5gSuy/K
EXdJFWAxkN/tOwsclPO/KpoI1SOm0adriOb9E8HCekIuiDfXF43ncQ15FH0JoL7F
x5Q/SSYpQuUOU/qbKNgYsHiFzN+w0v6Xlb7IEqsIsHPQtGEA5WQ0jtYZTsswdEF7
ee34Bucvc04pQG5n09oIcVx3pAgEgMdkRc0D+Iy1SVVbbPzWRvasXwl5cC8p04RP
3CD3We0UILAqGe6aUuqqu1b1kkGZNrnYjrHcedTbkftDipRkthWySffLO1Vf7EP+
nzVAegZinLapECDTvpY7ASy350cmIx+8LJARP/1YYUqtB3B+UDutotRU0iy3/7Aq
s3Hh6rhzgDv6pYvGEnmfDDiHgD7DFYmoDmDtN8Buvz1IGTQDn+xlM9agI/e4FmBe
RTxcX7dvPPVoGAu9JKggPoNrTDuLmXSOWAaNLWF+Mpitl0ldl9bAZJ6p1Z3BiV1o
DMCM4d85pmYF+kgFX53v9NYKcpzogJklnSA6LiB2FpNURMojYoi//K2Q72Bn+fwk
fQhf1dl4ARAObfuSeq0oXtuVLVkXvEAHSv83YAt0myPq1bO9GZQEjzMizq2u5Nk1
1Hve2VrJxF7hu7w28f6ZUcy3LTok6UmcZguFD1n/ALUsf0EW+jhw8wgzkv0pJ2Uc
nVS4/kUXwlhBJFe6y9YGt/hN+PV27FRTAfog3latAcGIGrMCQKrZZr5+pFOvPyj6
8gi+ZDkRBU+UR6jpTzjYgVMklY+5Bh5uUrvUOgOlZZsDFHxP83ADho9kknYVZ/j1
/P8sSm5B2tmHnsMzmCKT7LJHwNaCWuodRu5wj98AVLqeYbY/3kkqp64sUWbSKNAM
FfUVRK0Eu+OB1Ud0vaiSIo/j/xOePxBswnYWVzG3p4BM410y3VC37Lk18yssB4CE
OYGAGe2T3IXrwwk2QvQDIrMXWiMpG0KRA0lPohrxvw/E7cSJvpWYuYwqrlkQ/Qk1
gmUmXYkU8diA38fD3MHhpo4pkh34cbnuuLUWCeiWowDtE6IGC24H41hz4b9tUNU/
TJsbwrzl9r/KnRpYZC+8wJIKzx213jXKlyD8ercPBGNVRO8OrjfdlpQpOHH8/V4/
uNZJmVIluEJ22CVzpPVPQCaklMvcNcwWz0BVcHac9QUNzrbKz6zUkQy+IdW3vrf/
uHXP32g+0ChyuhlwoHyAtN1VbB5pibOpGj+uny2uZUYNM4nZJkYwGXrmEd2bddYR
VmaaYyOmK1cyelBg3Ji/bHT+cISiDnXHtW1Xw33e+1qKAaI62w/BdFmFD7wzzO3Y
khWIRUEk4D47apGs7ojp+Edvgo7QKrQ2BMU6L5lOji8uiuPC6qG3JNMFGMa40z3w
9zW3zRxORmfi7B3UMYLo+ywHHwXD4wGbU2/nyNSVkPAVy8b5sv7x3Mcl7C/AFQQo
UHecKkMaYS9c72kPuTIvpkYXobMCTIqlHh3a1BZp9trSSZKPcTLdUfVAAPrc/fKR
zjXXEKHiBnrVwKnCSylFmAv4RrDHad77KBg/mpmPdSX8QOril8bRlqT0zO27YXjV
yf174PaCQWIue0J15JBnouRAR3spVhG653mnffR+Q9+60kb3ir0KUMauwaf6OROB
gHEIMfJPwLid8WLr3lUDySKjS6EFVPlP7j0N7j9Be9XjXswL4ej86is84/z4bvNm
zBoZbM8aq/exmQXwDgcjkiHoF9vt3LFIzYyiEvX/viXepvv5e8J+Czahe6fCdWOf
FzfOnQouJsNaWuvgBDEc9Os9Sm0vBU/GWxWt7+4afFbQMpfqLDBPHZvW6F6aNeI+
wDXgixz8aV0LJU8YfPw+qok1++35q09uv53G0ksV5pJZQ23PRMvhQM9ZbRlWj3jm
zS2eKgNkUlFppkQMqV2XqfKezg9MRtaJOZtiGB2M/2IkvcMz5YIPL5jAaADj3sjn
20zvfkOEDG2kqcl22DVYl7ePS/+aKoPCDnxylYxVxCcjZ3B3cbNwWawZZTnJRZ5S
1P2rajWuKxDu0wdG1h6kcIo4p8j8tDWGZ5lbSmgQ01OMBYvxcgawOG9XAkOqirk3
qlK7HA/ZRtDlND6ytbGlDJe7paVPobg3SfVJ03g1QsbspbHtj4leRVwmePdvrsqx
KCiEOMNUS7ktsen+Q+uw6JtVGIjxyNuEAs7C7kWpKsXRCdR69nqyOB5V3HdpLPKI
4hdXlpzwX3FlwyD85DTpdiuWTtY6rBeXeuP20Aau3VcNU9WFoK9iOux2GEWLubM0
kenNZJHCpUkYRQPzNjRqwDULLE069Lude9XMN1GtsmVo3OlTp5zVQGMQj/MpX9P9
wkSCZrR9knIxWD1a+2miOmnUavQowJ218MUNoLgOYYm+QC6vvLMDFaEOOdksnfK7
di//QIAq9elG9XqAwYyM92yihiWaVbue5NaHwb8XMM1Fn+eY4T3Fe69zi669uOkR
VcvhJg7bHeC3IbuhijUIMV64ebJbnmY4THgHmYHO1GW+ZZeW6WTaZFQAAInm5WL3
IInyxUHV7MsEjJDZTJaVaHh+JE/y3Z8m3UitB2PzFm8HuFk3Cjw6p5BNIQ+Ydib0
0CMjBbNS7qu7GH//SypppHAtxGxthq1UISBw/nEA3CaHDCnHeWS0CN9rap9gTeYq
7N8RLKghW1nF4H+8+1cjY/Rg83e8xim6uPuLX8PRxcLGkjqcs6uPJ2FWHor6esaF
DQF+WuVLkjMPvd2R+Jc386e2kly5hLtkCoCOPGZvpBzrGVGdcIoPXYlQ0xx4odl9
CFPryJePdmNyJv7UW5nCq2jqjn9/0PV+eBLZ5RRv7Bh9RaRnIFV/jpaWpyAU+6Oh
x2cOlDVJuvE+bZ11GiLOKFO5T1kKRuxnnpPzGDlr6Ko/iGdjbvxkztrmwvI8tMIx
0+H8QE/OfWTuxEmJCErd7dxJuHl2fpC5U+tq/VYkXFReFN9gSp0t9H7fXwfrVpqB
Wq2w70+tiP1WJue9/885oFodzuiNCKCua7A/uR59NuXkHMWy2xV1cdnvD+bWIQ3M
77ewqY6iyse2PnMBX90X4IJn3trZP65QyDSVpQc/xfKV/uUaeFvTMOWU80JQRemm
sXauFWj0D/lrqSsAzYbJ0ch86gGt/HZ6Cnf4Wr/sUigY+P/wE8ZbgPQdL8ZddYwQ
HQDFZRJM/Cq3X8vxPTFHgnEgl4efJW8VZZP/NPAj4yzAsVucP9YTiKAJKRRYYGch
RuMJyG9o6HUnJ1mR6dzVciBJmJ1xVmf88TlpEecC79jOnPk7oJOfL97528kGXEPH
NusxELe5fLZu35LaO4WPLI7Vl+Ed3hVX45Ii9QKfN7CriNFcsK/3oYe9q6rzcpRY
K9D3VLH5xbKLsqoiZ08MJNG7SwSV0x5T8w7i9qyvf1z0p34y77kmZDqwafaiABkQ
gPhW+uAp1V682R0mjGUQ8RyRdyyu82BSuBRdP0xDsYFZKQTmaUetzl0H93bz120U
txNgDzzeminrOdll6w7nDykHJrn1PxM1bJCI3L0OqveuZ2t5zfYrbxDCXWBZFMgI
QIt+bJDlSAmv2K/pvL6k75L+POZk+g64kCUlntZ8yHoIo0olffu7NiwA3+GZyUPH
GpONN36b9qaKfsp65jKe5+P4op2ynvXqmYOoWBKbLDw7O7txL0Dao9bjKhFGBwZ1
HEMXxFVRIm7AFt9USAhIspucGFHsRAvy10ou70F0pQJGr2vWhuHzGYnuWP03I5Ng
QoJJ5qaOUM6yJeGnxSlvxQ1HQhm1E558iApb7fxZuDDaOHotls087QyBQsYTtTq/
ZDMh5RC3mDdSHEscnx+Iy+Eq7j69tRwb6zGX3GGvRW9oxB4a4S5vAa5/VHk2kC58
DDe9rQG6YruTI48V4+Fc1sp2E7fLGhms50vkmxt9ur7TgG8TRWCBBi7bBFkpTIen
Mfc0QWhxXcNxbH6DDCtEUtsTJ0Upe8VLAith6m5+N6eQEJDh0v5WUeBCRmEllYPG
1WalvFMp/Fkl7tFHYhQeVutYsq1+sri8pmcmdeOEi7W/WZrkprSlnkKGdVvqQWxV
awYKWVqtpfgOACJ1l1aGNaOgk0Xvvbwlv2kpGk8xJcu+a2Kq53s6fwuuGetf6BbJ
hYNr+QNcB1ccgVPMThmrGEtkeiiB6HNxYj01cbLf5QJ3XYJ/jO524wuOj9Sfw0TI
s2pYqUzLE+ul9YmbsUhhg57OBLS9ZSc7jsxb0sRdOnLdvO8MZyIyEqA67l8wmYYj
vZOmQ2hknYGvjV57uBt01z5jOFHz4WRl1uDcSnMZoDrRbEk9rE/Y1oo5eGZA2+GK
+1DBAL8P8e/InrYSusBPNCLNaROIxWQAlokwzMmxAoU30YMXtmY5DiMaY0uQyxp9
wuw2O0UseOF/x6F6JuAE64juErH69vem+r/oXfLEQfQTPOubf4FOwscbVpj7NLDL
s1SO7+DsAhIiHTYDnC3eB6vWjc50fhqFRTnaSZEi9HLJPbOkwCIb+eloBaeGTgur
ZPlssc+noLhLFZG91m22u40RM/VKcTvTNFi1FGX6da9kBasROubC2rnOYrYGmGmz
rWPUXYlaARUOS8z/imRYUGGTMiG7c9HDfeCKzrAkMs1wHQRIT+EYeIbH/dAnLM0I
V0djc+aDYm8Z6DCUmevZLYDGiTQLLbOlFiljf6EaiIRdHRSEHMFMeheGPeX/nG3M
TwxxkuSoEPYB+RKdWGSenUSbHGd+HndbdkNjODs1BqyIDM9fVcBRZWtOefccZA+/
hO2J/PDAk8wEakC1XQ3VUqq8Zvbl9XauGh+a5/FN2FtITxHghMQRaJHsyOJ7qoi/
DzkUWdhkiRF15aAkJ64h2/Ke7QuS7GhMvyaQSLpmKMiT6Fp0iJxH8chcHypBS+Ys
BCdBlJCPAreXMc3ZXBzW4AWHxNL/SwdbqRtFD/uKhhhPHhfRwj6iNEarWAlwY0PR
q73LqFMT9KAXzTt0juoy3bU6layYfx3EkU9kCkoRIVdR50kJnFhMKTTAlvQyMy94
8UdYVG1wHc/yvQjcruWlkEux9NYqhsQItOpJe+yl0suf8hyyXCuvbPP4NBje9MH7
W/tFVoRNyUnTW9g2kNRgE/ze4F8h8RQeb0eWNm/GHpeIG2mTa3zFhkKjR4ywF9wv
afgIXzCK2nc3H41AYH+4p9KN4QHdRduBaWcBppDs4TtF7RJW64krtmB0SzIyZ+lw
hnVOnk4Xhgd4a+1eSqjJ5wjL2NzoAw4Ms7pxCh0wndeKaz3381xvG8oB7qExSVG4
q/4HaytuF/krFDWPBEdYhfS8hxBKnduZDflo0JyRGJPlo6NR2EO2uDeTG510peqv
LfbW+cBc2WoOJknax+gJ55K94trfLll0g+bTdnar1oU7iclvi1OXV5sINLDroBe/
QPLL66aPPlX5vWDw21yfwF9TEmYhHSnVm2jIlzh4Im549FMB1Wmafyo5ymhuNZ+s
T6iaxyFfLgJLBS+KKz3bwNx91JLJ45c4ykv3Yg61f8NLkYu3FJkBI5euahByNUTp
mppmOIyHC9GiXVPaR7Rtp5wzNDOPfOLaSSJjXXQryWqnWfKGVBVre4SwBDHdmhSM
nQqiEOgmO4gvcIgbt6n1rQWTsMsZnk7Dm696T/JvvNKoq7qe3zJ6jo/xdsQV1dbx
YOqFfROamlIXbS+hx0bjUrfo224AV/q18kzRAoA2xFFBA+Ajd6x7VHcdSh1fTFsy
vUFROkP550RLCUwTag+guC9kbONu5Gbk2AiEHoiXx/BvgLL0DzHOBHiOq5nqB8/3
SefB4CAN2IHTCdCKw9iIFmDRMQcrwqOzBGkX/yN+7QwREI64+zizfFZMm+fd+vV9
4DkBQYFd0n7DGR5wVPBujgX0YEYP2mnaoImtbnl7pb1wrUEcTMB+YsEW7n3H7T+j
advniw7+UrJ6MwYPOGipiYTtwOcdPETAc0jCucWpArsiEFmg+qsbbhK8fbFhKV19
rzARaKCkTfmtfmEqy/VHFiM+Svgbf+DkxqVoYOcE6I/hkjuKXmIy+hLRGQ7cdfd2
eZOzskdA14mEKQsgDrnULUqvX0fw5pXFArH647EhMb0wAs2pl7lWO5X6Zd6ManUH
DErvEL/xN7nCVu3oA+b11VudY4T3xH64/aGgLPlBmEN19UVTzMrj9ie/RyFhgfFK
2Dypz1h8QPU5sXBhaARMAyw+BZrdj1w4aBw2Vw6BVjKWBs6vgVLRu2O3pXxrfbwb
+8WL7/fSzIGlh/sESakgl4vzkZA4e8LM7SJKlD1rhDMge7mUP7Pg00c2+rAISLaO
uPgUvmy3Esc3MjGKqjjq7ON+DzElUM5L7KwGlb8ePmaytUJnuyGTzJ71DqiAvjIA
4U4yljUN7+4b6+z2HcPepu+p/5u87uP3cqlicykfGj4Zn4sVHoLyenZhVrVgt5dt
zIAyL+JJ0PyzUxDCwzg7kfVdPo8oYmnXHTqeFso2x2MIlDku+pwKTKKcw5hNFwDz
D+ox3YiaaLaEpACJ8eTNVhHT9kbbmKWqcW0aZZfkSWzDsvPRbQoRxUNgpG4Klo8F
C+tRr/EAXV0sLI/0oMdK4WL9QPzpGJdFo9Y/6soznJO8T5gc3JIvLGVXHpIFaqwy
o/Mf5rriuoTVW6aUfepM+aZcpd1jck2jJya9pi8Ia6D15s8dPCIVij4svq6jprRT
jq2lWdwgZ3FsF2TyGZQsBMnL+ZpZR4zJ4mSBBv7Od8TV9ZNwJFp4UQzNUS0btB5e
eZqCcE9dEiLaNHWQAAGmGu26oQRRucMQsPSjYLu1MiZW6mcOYmJLQxTAYf8egM4L
+DhKutHc0plX/BiXSNk1s+ZyLIfvDvWzYnylnUAhNpSMEDR0DkOOQh9O9qdPi3tN
4dfEWYwVcQ3jLn53UiwC08tY9+dC3wnmOh3Gyz1uUVBehZ3OLl3Z6LsDaCP8cFiO
zojamh2Q+brOKWjEXZsSZ+Zej0335HgFnIRW+zd84xfHrLzMj2V/Mt72NNl4h2as
c6RdOUfWZ7k0OGV71ciUEo+Lm0Twj1RyjyAxoF4e8+OT17i2LUwhoAhSP9Q+SaAN
/yvdhnboTTwNyGDbZd9S27DD+ot1Yuzoh2aJ0zORkXYNwyykIJps3lrOPT86Apx6
WhVZn3MVCInMDOyDmOIg2KzZtv/R+bWlPmeu5bSyxDF+Y+HVz0YkAn9lycw+NWsK
Vw/XuXdVGLGsb9E4UuLaWUTrZnYheOE6Gi7l/hDOH0YP0KlsCfJhI72ypBt95Nn5
coZ6N/+85I9uoXCuVDtBwfGLJzCoI6IB5AFJgsKCnSvnaa0z2avimRqxM17d2oyg
Yh4XsN8JfQdREujNhvhHoF2f6rf0wRWGFd0CzAtN943hGBFOPUKNmZW7KW6jDfnK
EQMOZRu0qJ4GJfPfN5PyahbqreZxo+N0V03L5AtuDUZgGVQKeSBMTZpOYfi7GvzB
Rn6nznx0oQ+JAkEmBLp6a43qP86HjRM1Tpe9LAZ3SdnThq14loukOLVqNYBKg0G3
ljFpczcz/bDc6RjV57mKX/oSMMYIqvCEK0qM9DLIC5Xqc3ZWzffQlFmtk1lcdlPa
jy2hmgqS6LCRxFiHmvMsTGwr5snqQ5T6Pqe+BR6Bcc6Gt3+rky5ewROQnhEqaiDe
efxGyntysvPAbhsHJY7qYvQ05wJx+YlShhHQKUW0kIuiFoqvET3QI7ppWJ0eu9y3
5oN9Rp1RLLhP69h60y+lYA8X6Ez+Lcqzpy/0hqi/r4c/Z1+H96rs5huIUIqpaY7v
HiPjxxbYL5+nMWRNWmrNn/C/E/2JwLSWyAifdQTcOqg9qoozDBhaltd6nJjG6NTC
y28cxdgSoBg9lY/YO7gZEjsghANxS3oGFcm3di5ImTeywqO691oPo3HgZFssbpkE
dmdZ80sMoaZCPL9NaNaxzwySRF5kJMxxS5VEV1pEVkXX22KvgPgk1QYBdiZnbqkp
eHhMVvfEphM/aEI73WDTWhyj1wVR2xKHP4e32CW5mxM5jjbq9bSGQUxrlMcE8aWc
U4F5pxtM8URWeHBiU7HB+GzP+38c6yUq1QCUaGy/7QmEzF5jzktzQY9FY49szyng
wJBF8J/C2uZIOooCBd4C9k6Fk3Ip+s9/lFJWj067LrTqHmdAyMyXgL2U9kofdRWa
bLj1vlSuEdt+WXsGG5eIQbq7snWf2FvSm5nLTfo+BYUilbPoHV9XxgYZJhJDjiiP
L2P47qhuTtyjLPNrfigm59EGUQm1cbZFWYX+SYd2aF12zMFBwDJ13O5mlv/5Ci7W
ieLEZVcHexVWEcSb50muG9YxVXvSz1IUbiruhRqvaf9/eSvk53Xo0KxdwpF9MGmw
AIhll/cp1tlJXCNrGit5l0DB01XuHMp/0VUYXKxnwki2XlpVlD0fRJpQUka3jM5G
LWw69+xL+FvABTXxnnOWeH7cmKUoLDlTzZkGv3FV6V+qleB5p1vjXyh6GPIpWEaX
eUDxfA0gTri5ZKInRNIjJYF8jkcEgysolrO3CS9K99twu0+zVfSHciGQAee+o3n8
qAE+wsYidIvg6Q5R4BRsfiLiXM/yyCFSx8a+vEtKAtM/jvuxyzVkhb/peM9VedyY
LCTq66nwep4UQUZDFEJWsrbm8DdViBrlP4lsq992F7yD1ruq1x+9Ew6LKTd3VyGY
J7vpOn1y0LtIQMAX/64yZGboRi8sy+1ldfjhD6py+gkKMqDiWMjXFx3qjyCsy3Sd
C3MGkwJWU4d5L14rlO7u+O+itGscISxaN4Wuhn6kRidAzR9ScrcgZY2uzqm72Hij
6SoO4KjIuLapE1F4MF8lDbdpH5SI9qDwq7UhzNdc7pdIVQ9Hujj36fYErd1DXW0v
O4qaJePsRPX57Be4bJXVxvsZsQRo5ffALOchZoYOswC6VkT/HgkO7akauntU0pj3
52eN+MuNzIF3uBGZxA1Ree36gYsvIDTjHQAws2tQDbnYUlwP/2oUn9FcbcvbEgRh
w146J+/iUuzocRdF1rDoUGfbZIFFxa9klFjr9wv6pLob47x7Cu/WIcjsa0B7OGPn
3MHkkCLQOimQZT5GkZgtaw1gD57MMfJck/hk3lCV8FVBqa/67Iy/rL6lZYhwV8WX
dUAQX1UT5ueuBucg8qeKR4hW+M2N1p643jxXrCI/i9/I+oecJilZmViGzWqu2w3b
C3hbV3l2W13l9wrstTmLhVzbFZBO26C64pFoZzMqxWWH7VQutvYCrFfxDTWbNUG8
u+F0/A1ZT5uNp5WEXZ/NsGrjGMaSsvpqBTPD5WMvJkFYl+HvMZH/9Ty4GLp1rJ/Z
lPnSy89UFbQiI8UBTZ00GWs3BRg5hMf/Wyk7Pnu8F8OMalMDRLjWvilf8ARY1FIg
I10aWGNMr3b+sjtQMVnM87OfKFrblLHCQBf8ZkAyFTQCfza3GLjM5COHwCZwRw92
T5BII4i9B0ZZ68QMMw7Smmn/RJqw2SGM78IJLVaVBL4mChfLi1mHPiXkQCw0oBdx
jebpMqzb4ddyIP0OdvJYHEQIP7Clc5DSI7BfZKEFNi6YPQAJkGu2kY288oIP2hwW
mG/so34YjyI+z7qgP7HI13/ujk4QWDG8rHLLclxH4iNAzixtZrGkY5XmsONnJwJu
mXe/ejWfzzqxF2OCMaphVnECWkIqbV40R8q3t4J/nMLaE75s0C73cxWhkEUSd9Hp
DxF4v9MsM50e0sCbThGvF8qejeJAD/P3ybk/7Bcty0dMNs/qOPN6Tan8Jtf6qL5a
0UyQX2yHx5kQhTt2A6CNuVm7n0a2/drrt6hiiQOQ9A0HA4Gl0TaTuoY73L9KVsWN
PCruWZAYdRSbpnOrXvNq2udKcUqRyie5lCYmGGJI3lE3fQmLOA5RwFsFFoQY94D5
RroAgcwWM00An0Gghw9pMSlz+IIkbG1/c3wArmk8y3XZwc23EpQqTaKcrMwJWpgE
1WeuQW6SCUe27qxe36eH4dkhmAac1UqtCRMeuYc2uPXEZQAdO1XCgzmZf43G5SHP
d2kYLR3IFrkqbvX96K/JoSILnEfAk+pOWyuNxixPl9uU7q/8NMKTEdOgxEEnjhn3
BWda8KNT4qN29+ckeOlOEUhH1rrYo/o3Z5DLstsXkdTeOvAAP5J7UQcJIXKtvi24
Z0L2bf/nrHmP5815ZOMb+hUUwCiaOD4dapArKRF47FhYIAGh3atCsEDZnmBnG4Iy
TAz55Qw6+bnwmOHWO/jyaRc9Z9zHqirUtEkrRT7GqDzTAiYBqu6qS0NsuiOo/fwJ
Yojdq+r2btAKPDrP7ynqg1DzLX0rb4D1qCYyMTlQHkTE1Ihbqc/G7ecBDBJUpF2h
PSYBqSSH6UaPiKzXO4kendetdzw6LYOPvXdRKNiVnMDQSBrbT13wTcEjiimGcorW
Fv35TLGuIe2eercnNLsqdjiKhNoVBH0We44VUTXsLFddq2wjuGxhOXY0t7x5H6AW
lAwrSsvd3YHKm896X5Zka2oLOD21LJqFvFAVh7AMTRyLgMk8UONLGiVvkxdiazjk
V1ZHLK68zpnry66ZYL+6bSY/4p4QYYbQ5gHCJr4Q/OsAApN6lDcOoTTw0hS8htJK
q5k2j6zYthEWxUd+OzZgfaUzqNITb7iVwXkk6TSIvsEOPFUFT1ZcOpqZIcHNBPCw
iG5DGqjWh0S8KMSx2AJcerHCn8Cz1lmxKG3Fn47Tkg91NjoYlrgKZQTSHNILmJGe
kHjOHa7QUhrZDLUsqQaTFW9cgwbeo1YgkyT5qzAeIhvLWWPtKdSJqBS9J1T2+wVC
5+OWF6nmIEhOdsqzsNZHzQ4+N0TIZjzs6Om93kiNO1kAUaEHuMevY2rbwHgVQsqU
oFL9g9FFI5r+c5gTlz0ZFTeDTL7+LxFiOl4xnPMcaj7aUrOnvCDcTIK8dUAUHJK3
dGk07tn7/iV+4AP990vfyVL5zaM9wszBm24DEEb8y/eVqMKJA+CYB57S4JcWeGOp
8/VxC08BaM+a3OVKDrcx+k1HbDne+2tIEDnwRj+bu519pJrbuue3ctBijLP57GQf
YGcTd8yLLVES5leBZsMPGvwqbsLB6QO2JjWxh+Ojkf0foncokchpqffBHU6h8L+k
x8eWkvoLnnowDWRR3OweaNpzFv8uLzHEKdqFEVbthFPhLagDjugYlq+4GDkEAQtf
UZp31mW6UGvix2XLI4OSmj6mhITvFSN5659OdpDW4A+mER4ahh32Q2kNJVW0TMeG
RZY3GeR3i14H6xGsRL0uAIamR462KoPDsXe6QHURMhB0FTtO+xiedA+ZkxNzAoDA
TTVxPXPZWzaPqDMsaJm1UpbflxpMtdol1GYW0+htLkIwaCxq3qnGJhXFjly22gGi
oc5WDzri8o99qNxjgHWe8LOJ+uYu9vMoZLdmkIueqeJftu4CKc0x8tdaZH3Q1sTr
qovE7Gsu3ApfmaiEL0NiFSpbA9erZf0N6/dglocSj0+lqDmmUhC55fHRAaLR0ZiP
ceR9g9MtA0/nbIydiYFyQnd7Yz8Wetks4/0ZvWEZt30qQZJSb2YulDX4k8d5Ut36
x6xGxOpQVqd0+uRy2KSf88e7u5ptxWbIbThzJRq4Pnb6gVi0noIXkls9v5Xoe4CK
mpcWVOqZ7b4H4dug/qK7x5ZwRkhpIM0W9O23xajyoqIaPjSJB37sPyOA9tGTRWTE
isRN3KtyKIAL7JIrQCM//AHCBm/mVRyTWUAw9MTWc6dzxsYNfi0dJ3TU/5a/ipq7
4IChRSVnwOrawuVMXuTGmofojYFqgZ38vBrPtq4O1CiwmwQU+LyB7gDnaZi7DcVH
eXxyrAVG+Lpv8dPA8irbl4L0/Ujb6RssGFfcNf0MirqAuyzb1fhkcbpTPaLDYgjq
xll+TRlftGwJMBM1XFnPvmSpwXbIT+0fp1HGDpyntbIdfpgdI/HTn7NndcnyJWLc
oqkCh9uX12oaEVLgZ+C5gO8ldNMAhKpvq/8gqXM5g85hUXL6C+JjfU1emNNWSWD+
HEicvXwPgzAtU+e8+BCUbTuOsiXfvaK/9R0vaYkhG8eq7tjsxD/83tVtdTQH01kB
oxE+O+8OCrNBjvCPtLlHtl+FBC4siiuMxm3XAhtpiDmSooXN6N9332oviZDLeJbZ
MpWjKLmrgQjDw/q0op65GZ5wOPtOeVsL8SQvqJBsLKXHYzA5AdSm/ultJWz1UGJy
/wOhJjFUuBPkOGI96aSaLIC8at+nB6au7+aFEXlnMmpNyrIRo9YCFgWvVbYIt6Ld
A8gzARuxeY/3L6trdF1b182xsCLkx91gTCuUoaprMJMdQarYDau6T++XpZPTtUF/
6zokDkxjpVYAkq5iWFNaNcVlzBzf9E+YqYjcFjWHB8q+pOFXbPGdPdKKjaLm7Mme
vFpVZOWZLvMuQBGkAdZRFeN/KiWIBYbCdheajXViCSD3jiMDTcxWpQzb1E58dccv
o/bh2qBANWLr1/jsUomp6jnZ6wt5a0ehy9HsPVL29q914jdOELiRDbm99zDg41Jq
RkNw78/yPxyPhso7BBlL28/Zj+anG8i+SOeAeKX9HMgDLyVsk/TaURbDv5hxz3HH
cYywD0A5QkAFc+9Q7r2jnmybazNoncSxsbQQeV2l+0hUFGLhtkUT7NhZ70wqEhJy
/jpZ0wjWePR4o0weKL5fS1MZ+0uRNvEpmMSpHn+tH3jVqUlRXRTRPQ0+gFFOliJu
uz+1WTGyFPowjFTzTAqtR2d+ulY7gXqEvZoFEPdbD4UPrSfbc8vnKxR4tTcOJpjs
fjrMg3O3T8zEvM/NWaJzpmzpZH07naA66NU5lPP4mg5AnFiHN3wBmGTWjxqPSM+1
YVF8sl/jpJUxW4MRGOygy7Yj8nwM1fkX67BLKaXwIO2g13Dcx9gV15kBl5B+AaGF
/ttuWRYTxmnzqLaJYU1rciqKahNAGeG717lCDlSerJEUru13j54M9U2+vPfiAnkX
i5eN5c8p+07X5aPfaNTo0mRmH8Tak+jYFbT9ZMqlkhL0sSLPZp5um2jdMEaETCy4
8uGf7Lp19eunGBTTuaQBohQtYmvUgYa53sFDw97RlKoGZQ16QBaGQ7g0J8It4jW+
s2hzukjq+SOmfY0UKp1/20qEpxlLNjQgNtNbzO0vAtHQHYckjA1EkpU9NIOQcEsT
O98j9OcdDtsXZNotyuCexK8fqie8Q6VtjRZBKfGMWWl6sSAoq0lbixPNL4AmMyTV
jh+gR/JxvpOXD0RwT2XBVtrZbQ5gQ0m4IAvie34SNapfvNHi/Y/6T+AXEVcqnNgH
9IgnkPRQrhiXK7SulsQrF3PITu1YXZsu+RmdTA/jbFw7TKfkOeN/0Jz8oGEQDVtJ
eJYHXcbXhZo7DOxSbm/oPmQvOCS5SRYXdomD7NVfcH5pFlDPyO08SsGmdONzf6SK
GdSaNcOPax/BG8XOLA7oXxzBQhmQKRqSoTV3TAr31xIsz5AWlV9lybjVgK+ttwVt
adCB9Ql6I91ngl2BvPs/XyYNwIbOwSUcVMGyvedYtKMfYS9GBKLDdnuNXz6KK3+x
eYEPnZPvQX9m2ASdHWKiUVhrmubDYZOMGIH9olc7UZM7Xyf6Hm3b9PuhOzxFfcgi
rBA27UUCRTflvP4CTDH8OtBR8So7hCa+tQcVSqWlFQD88vnuiN+okDE/kwXHJ8+M
qmoZwGNfmGjYN5ioQ4y8WhzZEw9ZOoo08JfPsgBP2dwESjmQDWFcpAtsB/l8xh+r
hJ3lfCv4KTA3XjCexs6mgKkLZ/loLfrjcCL8BaCYnrifuN+qyGa7z4GaQu6h1mr8
jvzzCu23aMFLOhd1UWNsWr1JZP53vjAsTm0WCFsaB/2DuwCg8gEneZbRr8q2PrqH
+grfQtujI/13ydTTnUS0Hk1PgntCfhVf/XCHn6xqMunrWW8p6g6Aj+hQYUOW1QaU
jViRTmCYBiFkHpY8DDEFo2w7i+bwRr8S0+LTwknFVGanF70Irg4Df6QA87TIJjw3
rqNVIWbqHTt0YWSMKwjrVQdjY69yZIvqtdyDjfQwpsp+K3C6EKIwEcEgwyT7arrT
SxcPQN6u0ANZFQcwpb8iPMk3uJtsldlamysR4ZO1ZWlGZvSRuBLEHPd8ULF93uCs
yUfwfr4/ba5PHtIQ8JW0+fjwE6vjnjb4YxwVPbGSk26L8Fvor3fp/vzjo5sB5UyK
g6krj19AQ+85JlwM2z1zIasMqIp7ksYvpXDPDODqZAJM9mNhFFic1X8wFREEjaJv
hP+8Jref7xrdJSj6iI9iUxtrI3uodGjNrFG+jO1zyv/QayxVQ7V0MjVYAMwuPoad
bI2nMlw6XSk7J4sulpzMNi1uIMVEC54KR0cOPXYY0Ffc5skmKKlZF371fkhLmq3M
fCKyOfgybagTZ2UUjvvV2t4Ji0ksSKfZm/dC+rtIo+pAPBhxMdBDZt0mGz7NZFmD
glwvccvRPKY4g93fGbeD14PNZZ5GW99knM+WrKb/AfTAX6fzPpT+UpzPSJTM2t/U
Fqljv1f2ypnsd6f4WbnPuin4eIQpzhGmnwrYZ4NI48op42tuM13F0izBzYYryOCL
pF2vKKQ1ifl6P7uLGSKONycEjl7z2fI2vywBwmgEruJOoQ/ukup4UI6EMNd7Aroj
Go1LXFFBIeKMUx+IDPLsN4aidLBO7BmqtfG7Ym8IuUFJ1GeX0FdGGkMR5IZrFRlv
WkU48yMlbxWwup3pFCGgngHcC3UuvG3TJWq0qQApinTUCOEfDPya279AMLdvc8NH
EYETpxhkypoLts6asZMvGZfuPMxjd8jm4J/g8YpzU+OyfoZwvSpNL6CYgddNFYVw
tMG7aqW7rUN1bokldvec+njTLFjWAEe3S8sgvb5ek9NNM3g/8MKaYXD0CeUQy5fp
KKJBlKnsPhcx8shSdwokezrEFjltgb+UDw1TyxbDD+wVe8QwAlO2TspP6wI01Cd4
l53V17abtetdXjcND9icZEFk9oEmwQvXz8O2pMFoMYroBx2MI6ooJe1RBeDKoK31
3ABjO61Z3cy2pSTacVWtSCGImIpA4LSDk4gNwnoxfB3MSnKsH5QWwJBNOp6DoRUr
7rzV5xVR2Y7Jgsp9WP0Vj2FEBuj3zKyanx9ElbnHjq2nfjkyvTdhoL5OWMTemei/
O/6f0haz+/CvUX35arWMDQnAmGnVnZhjbi2StbOY/Nq9mOczIy/o+Hn3iFd4y3dU
rj1PqjP0WRrdPjEBKpQ3KT/rw5JnBclpiHPbxHpsOALVUUDRMffY0GMtca0zSgl9
4NqMx+ZpwcfUzElyDNuVkSZq2WQ7yVvNBFImccV7fG5GbD/L1YyLEEHodHbURSV0
xPYcmZNk9ypWL7oaTGBF5+7ud1rualoTuMDDRG6eKz7NoNR+mUwtwyiNwGncGaMg
q3+Fm2TJC6BD+M+04sxADJwJTBxPVG64sfqtWbNkOrHIplHzkT6SSd14v/wZq9L8
k9q+4dTWbvsknKYRb0f3YbK0grT+rLECe42Rnz0n50WaC/G5d6VdnX7tNMkjg3lL
E5FF3aYgW+QFh46/60yT7I8TbLo6tNUv4tPARqBq8Knc3dnjhUobzhE1F1YhbIiX
QkdvW+MH/Ep22Zl/LuQ9o9N/i65cjabT05fkBWAtxKmHm27UF7qXGgGC8SWi3Lgi
iCqVhwbJoiz3noa7PjOShL1FWJVwnNNrlv9/zgMIgmDc8Q11ucuzJHUsqaR0ovam
R2NmtddfypipZ6m2nBN06OVXjMIYbooBypYn5Ac0wWBBx7MKEpBoyrUzcA8DrYHc
YF7q/BNqdBHmPQk3roUCzOIltPvcxHSINxD8XpWAYBKEY3jWBIi9NZtzt3TOpuA6
OBgPlsBcKzHQbO8K5+H11i+1B3OTh93zvDYUNMmw+5YrSHBiZzd8jE23soYW5WOZ
o6Nj2PwH+pzTCvumGLhL+XYG7IJ7Kw+c7bE6fUo5X3N3VLhKSHIRqiB4N96gG12Z
DfPQSJdqzM7NiwHiiiVKSPPj9hFjSyUebaf5o3EFkf0PML36krCnzjYvXOUlFzDx
GyxEPLUq4LufYv3CNsbcCg21wMAeY2x2yOMf38Q34dL36mIiIZ/8SWjVE+AjylL8
0gW5H2c0aJWSgPHY8CtVHR1A62DwOvCQUhZ1DPjs8bwJcMnO5cyaSeRgVnk6xgeS
AUJDMJYcLu2Fo0pLL6lx/UcKDO3AD7Qr0LzizpKWooM+jhQzRVbptdH5lTupboVN
MEDlIhD253gqGVpcOG3t1cpbgZ9gFnpSDzQvUpkPk5nRSMb/Y40haXkVRYEM4zAU
86WuKpPe9o4II26gBAsguxsQcLcvol3y8dlTXHjP+5LtQhqdU415WK8naWVUPySu
Q8L40zkTJUolat2D6MMYqed2MyEWjBGqMoisNEaCDchhgQevmJMyqfBMs3EN8EJH
P3yBn4GVjjaEX8zqctHNWVVjzb5TARe2838GTSVqpFCplKmLqjH5fOgzMksJXpdl
iPE1R20RvRDPe7GMyOqhuM7gPd8ukY9AKaHYkqp7u/oTGjvR+i8iOTure9tqnU2T
PRXjYN4v4f0vEJUCYV8RkgcfgcYa+2PggsMwFuC9q756WdSYwhE9x5FP6hkRQeeo
2S8SQOXJPpTmc6gQsfBmoRdIDmZ/GpDYCxZCbKPYnR0hJ1SrKH3chy8KgNXlZm/i
RIC89znj0t1+945jojQFI/JJvb92pkxWXv6yJxJy52QCdtHpVHhlS0dKGLiQzZc0
yPxO5j0VfurGB7Rj4Du4JGIbDzT3Un8whDCBBIHmT9GHPDb5sbpwj0rRXSiUDSL0
l40oofaUzo6MZOmZwqvcrLCV4HAGJiCMgU3ZkRlSZ8DNNrMTPLGFHeiVqXwOHujR
XtbrPYMczRNU3LDnvOyxXrf6roe6el73D7M40L9uS3piDlW5Cu9a9JMfdDCz2Jxy
79IlazSRkivZU+eVzkb7OOk5h1LhimC3Ve8hRdCI06/FS6ZjwjNtFsVAyaxQseGs
/xn+iOa0cVvX08go6IDrqE/l54J4XQkeXmfkmlUFknEYVlyUhCWBhhUL2aqdTwye
t97AA58Hx2shXkZ2wjqcepL0+ptKC/Q76065QGv3Q4ce24B3+mvDSnBqqbEIcqT4
1mBZgH2t8GuAxW8exXHl/JHnzg8W/buXn+eST8kzTJdy80C16HYhjVJ3FKVWOAnh
b+xNzMFWI7yWEPF+pL1nfgK8ORduY9fYS+yeHh3oB/yvd7zfGHT/6jUjI9SpHkn/
+NgDzdo/nd9pTwA3w2DJ4Y2g451f60m2Yinu7OiI/JKCQpLccRnTVLTn1nv2FLwG
1/xJchMaoRKnPf5pLfB3O/GzyeW6ozND2Q0CAZ2NKpE3V3pmEPsLHYyLKeIfE6gy
ddVBwvTHf3TknFXnZYiCTwD1ro/3whqy48uFTLTClUsOx0Xa2VmuYf2ZMmjnwtT7
QM0cZWqwwAp13mfbzCtxxhc4/7fGFso/IUCjR4oFoqDzYL9a0OawuMbVkLbWyVZc
cl6y75hkBI321t0h8jdz6pcVIpbAK55BWBz8ek+tMZ1+SKB5Acg+gHJxFa+TNTRL
ptq5Nslg0gG8VL2MkW9UfC7wRnl5JHANerGj/HJm2gvJokexezJyzZrDDGCo6uxH
cntDjpmp7gxbFPOJ4Pq9sI02MBCaaD/D/1I6ZKZJAYaILje9MAmtLNiE04Tp1bUx
wdONlQzeYhyToX8WmeQ037t4vRO0+xhNwOP4Vd6Kt+WeyrXuc3w5bcSg77c4wu7H
JNRqRlY88sv70w2lj2QsZ8QCpms+Mjb6JRwC5zO25/bDelDpL0UYii96hZWDzwiK
bEwQhN/9FxPFDelhe410TmYd+SemnlfHWblmDlx5VCECoybO2pubDjZmcP5e8Xo2
iyN0eylmttEzDcx4nP9gKV4axk0HEqGcWXmyo0n9VVusb5oQwb1A69ktu21DkuNn
bruVy2rpogez9yGdM2aXcuoEqc1TGvDckLaBNsSShbdLwXqL3L31W3ikTx/4aZYF
1w27OT8RtUYXOwXdaGFyICQZgN0KXxQjB0FxrGFHduhS5M1rDplE63TvP4Iukgxh
3snOqdwoSuAYtB/vfJBFx4vtwRXCcklII+Vu0WdHPR7MkRInRHCWPevSGo5QCYFo
YF4dJJocorSLSQuA//YkEdMPn1CKEdMyJlzl3oK1W8FlpAPSUAZ+3hvjpzgJVQOS
OYdTCuWSpF94A8J5nMhuNzjDWWmaAKNhIUg7Ox0VSjS/26LQvSzYD9qfwd+uDAdd
PDxIJb0bY2uINxeVMXtV+wgF/yBwvfwNcsf15ksAgCnKQON+JOfO4uEJ/1JenME5
tFoJShk3DNuCnALZYsANhHQOvN5Qu/DoiCOOrmlkLFyoCuQ7Cv2Inrye3yvuJbWB
PTpDaQqW3+n1DFAcd33Rii9VhqRatskcqiB+a6XnWif42v2exk/XwkIYfvYoEh1c
Dq/9yT1jV21n/gQ2wOl9t/5XpCmUb6qd9UoI7M4/dPDSp/WIdPUt6AkdJh+SI2Tq
DA+J+h/2TtVvjoTwt3HH5PCREnpGvRYkjj01pvY4I2xNmIno5n8jwtrbe1r7ip8Q
v0aAWfVWXzbg8/IIVSUVUngHWLHTImbbr7Xnx0BV6diTZFdMTOSyuviqBbN39Vir
ECtPz2ZpBuH7axeYG9QoqG9RzONjXHpmPztQUiQQJ6jDVPuoZNtBSR+HYwjx8n1j
1KDGJ4mMwg2dk7trS8bKfxp19nJuHPGWraQ6xmcA0kPXcAW2vUc+tFqnpglJ12z5
3u80FVQoLxvoxFhm5hoerU0u3qJF2iwWWBUDeC0V7le/lGE9gotOjrkswhedPJP+
rFALBXO5nhcW/AM0fp5ZGinue1s6Zkl3kv0wGj4mYUp+HM9H8N8HV6+Lke+mdeiN
1Vvw5lWdQSlslI6xp3/1/ochDdHraOaGsL9/brdhhT9YIAx8KqRc/qAnHCEjL+f7
f1+yRbICNRP95bCd8/GB95l4lgiypbEslbb5N4Elkrvvmgfo3KaPz//7NY4VSYWb
h0sbyNsB0I3kxSXyEaLmdbENE+jtlwbaSXmacEUVXFyb7F5Qph8B8U/iBhJQrtIv
rubA9ycRf8pLFhauN7xQXTO+04ncmCBq7+baveSvzb+f6eF/8AabLyF9gUSPeVa0
rl1j45i/sVzXriD0Pes9JtPk2ry7G3P+itzX2wUQ9czumL1fuHPJe5AMIzv4DKGv
lYFLf0HXKc2fCyAOcQEmSp8/kJF3iudWtjkCfbXt5UBxMoWbkFp5g27wJiax3whx
TMpFIWfFGwqslXgZDZeILh+lIgJqDsvDf7qq0jWzaHVcSh11C6zPhob6PoTs6pt3
baNUN7jBMLlSl/21cvoaCagxwz+jmhcGAZ+cWYwgv40qQhKRPRkfezlpQ5UaVuk4
bkFovxHnFmNvT2FacccFkn2dQJ50X7JTGfqWmDNxcFWI8yhVdlO/ddqm6yw5/pxT
s5FLTUDG3724g7ISJd8GhewCioe3GeiKyteS830cm4Us/pqLkXuTBJhq13rPAihi
7xfiI8m+YBbMkJilhfy+foVJwg08blS4YO2+Qc6i7BFjRBGUyQe8LztWabqcrcT+
Wp0puUGJCLEoOgW05DkuhyjEhfG12cLVMdWqcHqc1WCJ0NNkGcmkSuF6+QvWEJRA
5FLElv6L3iu+XWgT0tZEscizS8BkqOhc5+ENNTy0lRXeuYA6xLg0ruJGWQA1Z/7d
7FDBiDddDFZttokD4R3WtnS7w1ARSNzyixuY/CVV9J/Nt4mQgpzR1BqxgOzAYx2a
eq7p/BOinjWgEOzi5NmPyDdxZ9+sTRzMy5w0aTf+BEfpFAhoqCHHBJ7tThTHAlk3
HUddlszNT0Q5qIbQ+ts+37EwJb+kGPQQs0MZD1Lq1wjipZuOsEMDeFMqZfrR+gA8
krLiS8zG3yfgVYrZIHLrBFtco09Z9NN3gBtw4ddvBL6NOZdHXsYB9MWBOYERnAOI
9xaWuOdcSbVzBdaZ6jG7fzModCZ+mXHo4gt2hJOkwhUJyaVCkhxoUpBjuag/Czez
cYsdllwiNFYHEtk46GLCWP2Q/moLNL30QUt6GvX1WlI7felUvmZOuwjUX+EDwKxG
vWfFiyIJ/SoxINcGoSqp+QUoA91yJIqppx5tLVxzp/SQySAeXoo6EG4spqXjvpgv
te/sKraHojptV9Ae6wUYO691vRWE2FkyHsO+FIgS5zahfzvHnaBOl8PL0ycygenn
2mEtpvZex9g3n97G+CKMi9YVOculcg1MtbaYS0eVQQ4JGNjHau0tySQQLWdpsTi8
Odp/WMEf99GnNDOqCftI4wdZeXKSD6m0FvBR+VGwCWCO2PRJPYIxyArsFQ4hH+7B
UWECelE4e851sB90jeRrDkD4lr8M5nO2j+O0qv+PZy+nlT1lraNzk9mTRbjfyj/r
vhLMWapJMvlRsVVfkkr9aMyYm+1pyYY4Qd48xOf7R+bcVEF1aM46GIH6M+BGFUqX
uqbwSTs+Soj9kcDz5b0bbe+iVI7ZXm1iXrDfTr6qDkB5r9I/jlklsjj7SnFS1LZw
Bb/XXQOHfPo4pQEbxRvfCprTpAcqIYEvTTC04sd7veD5rkzziYS8hd6eF7RipJCt
qiDei/lP8JCLvZO3VCEGcECD1i+tbaqKNKX50xh5m56SpBUP+U6t2B9FcEEM4wJi
vJMWPuWqqs6S9gjBbHb211cSwskD2ScFJWKC+M1fl25fU31bK+hnP0XZULoNzttO
pvSA+h8FlmE50ndfN5kOrkFJvTzUCLjbJ2HHQbMJ6uGEnr2zHzMZlFFtMrsh/lEs
0AKvWnj8veuleWYMAfblEhfJAoE7Ni5WPKQcWQNHzYRK/6sXi8NmsG7fSzXDgQ9r
0cQjiVFB/IzcgMnbeC5iY7qH4onq74yQr4qsgcaKKebSVCY4XHqHHb3QMKsJNfeA
LUGhBLmtj64ABmzCry5Z6zuI2y9aN6uetc/asu2Noaa/ERB9ule9VG+fKArsIeVV
baqfHcWfJvAAZxBTN96qH9YBkJGbd8+D8hLJlU9DD+rt11YgH05g1fNQk/DgxJN7
y2RiKD7KlbD2A3jaARV2Ej9C+aJXbf+EdrfiTwYTzVNbN9MlrQkfEPhuD6n3ukuU
Q9THhxlK9FX17pYA9NykOHEC2bxJWpR4YSbLJOuteovOne4N6GSg9JUL4ojDxmsM
C1Ij/cV4Tnr2U7QgZfLP+uiD9mrWGh4mFS0cABcjjOUr5ie3ogxKvheDjIuSnl76
8OUfyEQmcWBjQx3567nO1QBSpXPXIkc26rRWymo6CvBi3SAnuBmIs9Fk5IcocoeG
z4xVQdHR0OIqkPP1S3COIbD4v0KEijIVBKrH0ISjD3KK6y18/sbpEuqF1Y9yJkwO
hQ21bRAtQ3KpeZWYp+VHCYaMtLMttkne49xNfFD/D1jjD/rjsecSC9A8qQFR0Yt8
sde9jrxoi3ZTHhNQm/LkAMOwJRiIYnFDtxOvsnki01thzBebwkdRr6lAoCmYQY/8
/rKaU5xSqlOm+WCBcL9UfDrRyERaoPEfvhEVafdjZffktF8xfZ17SSniikPB8nz8
VUB6zM8jNri35q23ZPUdPdWZvawpL7KxypvcMYjUCiOFYeHy7FNnwxVwercAj7rq
zrwl1mdazJezt/DCd7Ibp92WNDrdSHYjpl42/wvfzXdP90tbH/U9RUr7eabtFwEm
PatuMMhCx/2ofyEdwUVJ0MF90IGNdAKJbxnJfVe/onlprSV0yZMGbfRXVwcApFwf
na3MZZARLbeGcHIWQZLiJrsbSVfAphZZD2EsBoBRiGQLhetrwuemnTS+btLZMho6
5qx/2GeF+0qShIMFKaCGz8i3EtUDk3Mab6xaUL8zRzffX5hr5DI1My+gqAh/JnLm
FMKGamX7tZOvY9aG0O47Zy0InNBGjkf10WTECb/uHdyafC1tZhTRTvvf5OSZg7Y4
OsRl9HN8WKQ/JpNfs+Th2ubbWfqHIVVkvMQL0mjDkVjy5JUKvTNAUeydXoOkSI9i
jaD9lrqOb9xRx3v7V9PUbLfSQdzT0UVMDXquBx8T6sUxgHJknLfPnLz3OXKlhGaw
iYm+JLPu9bQoFKt2v0QZpbE3XsPeTYlTDOxxZ98AUgjOoo1USEm0SvqxHDWKy2lm
qeybgb/hS1F7FO5wp5RWP+O6+0kQhx0CtT9fyulUzlelKaqzZP3xFTkvKGR2lclm
gz01rKSVvAYQBL/0AtArys9q93u4ZZJnjXa2tu4qF/xGMFv/5Qx0kvFK6VNcHyH0
HHREYvjvWDAQ3cF1I4Ww7qYrfNKXUt+hIl5vqrjyzTn+GvLU7k4V7LL4JN6M0bYC
EWxKKVKoncJZx/v7J/2HBbco3wl+zSrCPZwJ1snwntzgdwSQl+PFKK5iM5W0nab4
xYLHFffaqlhV3gsyAIzfD30DcaYsdd58/DKjbq3DBKSH5NQCY09o049FAP4XOOTI
NC6qN6wcTxxaVj13HsGcx2DXyc5xB0O3UdMmagioTAMHQnKIRzBJjKKjK/5GUxP/
T8l828DMo9bI6+fZhQ74eXFPGRDHiMnUy/dPqcAw8nlAScnx4SSmZYi5HVsZCdPX
1bbGmA/SWREdJlJLjrA6YIbbh2MuJkG5ibjUZ4BhVblngjFtXNhfQziWkA2DNjRb
DT2nDHnCC+Dov4irGgmTN266Ct6ekXT5vdYdkOKRF8eRj0HaqvcG5M9eJpVLgZFD
V3lIHUBl6uu738+0kxpx7belquGkOGt0Cj6D2YTzH4jp3PuFxhF/KWtYXP7BV2Bw
dAFVgkpp8p5SQf2A1a6x7mci1AacT/z2kCD3QVo+3Uc+d4xOECkTPMs4ijWO0qg6
xRRBP2tqyB6o3xYKmpToCk52RKlWUZ1ZWH3RCtwhzcA8AGuQGplOt51EbxURbtxk
VSbp4e/h7KiNaxUIe1NJ92ISk6m+ojaZVeZ0pKNIF9bRbjXx8QmtuCNCc09cTXys
Q0iEqqDmezBc8bXF8b/64HfFbE3zFIdniblfeeKnbbCERQ8qrLSnvUpsnFnpRjay
OFDxMEu+C6EcjTglaEV7IpPvInX/W+vi3tmlmr8u5h0BtJVcuPprd8/1oE3CN5SO
8ifJHnKWoLEUsQ856Nw0dLCUN0FUoF9Nv5wk2ZdzZiuyZuzpKjVO8+a6YcF3MXYx
FDr808kop5jD68xBdBL/pRqlITEwEeDxEFX8Cgzpjn8YJo/8klo/JSLecUyr843g
XBcMnw5t4PtKPPjexV22TNJXxdJqt+kQ8YMc49fT4SEwpGpmvmObW9JpIpzqR1vg
v9j8Rz7L9KFvo6I+8ybkEg4vmbRSuiOofPXzuKmqpMuPhKWgDyh55Q/w5oCturDx
u+GhmDSbdAg6irXIgwdQKugnzTEb9Xi8ugZ3feClyUeFqLWfZqjw/IZPAM2FzTpP
8bGS5LJANQFCUAN8QxdN0ktMGreFO3JmpuASnlWjVpQSDK1L+D9aZbJrdSmfOi8Z
P5quGSyqE3AQMVGPhFAd5BmRkcOJRFnTHR39gG4znH8Df5fv6BFE7NCjpFmxzVmw
ED6tVmGSlRkN+HDNC8eopYDqYk/PhJ8ZXu1tYvtIQ6wssi+oE78+ZiKmXbTtq2X+
wZhruJ/XPbU1u4x2sdrrHZk++afVsTkcmpxUGG5m+JV5zZRiz1SqEt/8gmMSyFuM
7HV8ar5pPDzY72xgT7ypNhYbzssjtpxGhqV3WGl0tiVHkuwcW1cKwvZ1w3cpd69y
1Jx+3t/lTn7ED6LBw30pDOWgzUcWpouirsrVLXPm57RrAV9vDKSedANVlxZ6g51u
pp+W/+Yz88KMhbqyXOayn5UHY9hLTt3GJjyMGLuhVzSdrFtE7rKbYnVxMoMzHZXr
2lr+2guagDMI3eWtvtNdZ12byCA18NYrFix3n8JpgYs+vrTM1tp2Sm4BP01bW2mo
MBvlb8jtK85Q/cgswAMyKs1yyAv1ohZ3nxJkxIpGNIxofDRP5TNxFuNkirHXsNBa
m7/ki+PzLMZhepUy7GDqmJkjJ+uc+DzKSpELBgGFGc6tCpz7+16er61bVmumqlN0
z+YcWk/xSs+IQLWyMvg5rYfihPRTvFvNLc2hbUY3NfbfPg+LUWtZcWgqWs7zi2Ct
7MQd7PJUi8V88ITJxCoqTCQyS6uy+jZ6L+uJFC8N/s/VDs4AlP89YKPV+LrboQ59
W7uR3pzROW5Mo0mrkG1wXGQKAYyD9WAFmJNQLLw/zXH+3/wOBqhexOv2mzIJ2hLt
Ssh1L+CXU5G1uFK48M7/Jt3aBjp9ckSJk07W8bCelNMwB/ehHWxFpwTk/0+kRHMx
eN8Um33zfAJ8gpYCfLabEyJeQhYi6olJam+9IoaKHqQZULBclPiWAbs0Ej51Lbxg
+Xf1vTDr2D1r98in3dh1fQc1z3x8vJhKpUdLPbmfpipr7aVg6UoxLsN97sGOiDVs
Vqbx12c/gN6eNs6we9JPY/RzOnz0fk6ysHOZ4wOJ4thWTCgpA+XnOMSfhE1ljv8g
sTKL7/p7yANaeO1NozanitkmHhYgUI8uMFjI0+9nMMCilSnAvukRd3hsA+aM1a0I
Rc6bOzUBmZI1BURfK6SoWviTkWVfAHvEkxey3k5sN9oIqeVfS+EOXyCqvzlwGYPo
fsU8sKdNHDkeomx3Py2e/DtkUEVrMPN6EDOaVkz2SMUxFX694q3Xk11bj8ZpqBmw
+eBZNYrnMErAQStdl+/+S0lwj8bkTmKKVVD/W5/QiwoBYCX3lm9v2AtkwrKGUl1I
zLc2YptHgMHS3xPumtEd6JhpdtTpuidd+xEE/X9xpUKyyLBEKqE6svOzKLeb9Nl9
EVv6LHOS8rmZPBibiaPzqA2HFwMRmu3GM+WSh090xf/Dsfoj57VaXjF6jmXn3YSg
pPFqe/pfFBAeRefiAb00ZQzwvQLv3t3NFdT0hIJBSX7hjEeYSYHPBsejBwBGJwXN
S5erKSM+Gl/sbTwwTIi/zl2JsHX2oAipskE/0kKWuNZ0xuUmfNLouJ8ZXZ+8TdMR
1PS8HQfFTD+yJl3QraK8gq1aJbbMzwo3TeqkJ33QvyPkbBGd82k5bP4stCa+dyBk
9hyKJtIe7WiApSz/P+d54RDCX3cXQI/bcCCHOyqtxgb3TJnNjieBNZUMRwd2V5rM
ZFzwmcK+32K8YPoyWMBLSe2So/3+h1Sv2ykWczI1zwm+8slzVICqCtXJh2LP3Yku
VmxYfXYrBmSgRRW8Dd0gccqmgmau8bRYbMfaViQQwboZzaWU62oFYaLiMVkRcvrf
d5sv12OnZhLmrc/t9m0NqZPiFLa+N05QLb9JBAF64WP2aRmj/o4AW/3Sc72v0RM0
thWLQaU0Ve8B+dxHTk9vlg71XC2oJIKViZwtmufVJa+AuNUe4vW2Tp1bLei9njbm
g03mi2vnlO6okrUoP1zmuDduNQiN1XL7rg0LWppT3vEyZFBx7JllgV+mVD2lQe4S
Hbk0hyHGqrRRBQqr6dgFzzjxJNRtZEJ5ymu1ukqjYYiX7tT/sMCzp3GoDyRwoO8N
wAQRyJcQ6qwbRDiPdDx9GjAEq3a+M4ldC2z+dO9ZPhH4vXcU+t/DSQ+Npr55z+mp
AE8WpPUCMoVtt011HJ7eAopzYAb85n02Nk0jLmuPNgoQ8tTPRm/1JVJY7cJz6dmz
XTCyVYi+00OiQ9NNu1/icn4yKg55XrB9BzpJflQLxRbmHJQRMJic6FMOt3gaqGxb
ec6HgH7xxcG0KUC7DsF6ThK/aG8oC/YFB3uorvrPFn+n5NVGcZh+lgPO2+tA+3O2
3ECkAbGbV4Lh8fYwTACI2lC95tAT8kkmJjxcXulbxewHatLphUhc4jTHokqopR3C
GiSPgeLVyoGc9jwYLLkNbah1PdaZG43il0V7GnThWraMmejW8zSU9VWhaa32hT6a
xdPh2AG4MUz0IlF39VTb4Z/IfVUVxFIkuXG8iI0iwput04HJLLljlUzgyKTLnXx/
xQcHMmPtNnciNq3ICGOtAfkW7Cudiby7PyPngLc3/fzo4B8Lr6iVRlRsyBKlWGbT
GSp+QawkhmMBFSAEvcZNw65Ywf/mLVawn4Jgm66JUIaP7Zt7+bncrtW3bxHqpcLQ
VJ1pQ3jnNwLXWExAnTF9ZYqUT0QX5RJ8Eol8OcyhlmOHxsbnItnoJ7Z2UPgagv8G
X6LMDPKiPD0/JdDaSg8Cx2FSXuc5GaBY6rfeLQnkWAAh/ftjaw3GZeDUMdkilouc
B/rg/mneI99f7gfurfWU4bJzTlsqUClNsQwGc/IBfS8J4vJWbgv2LYTTc/pega0m
DNw/ajd7UP8Ue20uvPwO0tiVmXKuQAcoKe1SI93gzbWW/YasedRHovufUwPexl39
Ugjz4/nzc/7004+XdKZazK10SvI0UrKXCBz/JSEDYmvMVDioI0jl7ezDjVhsIc8j
Ia+8c2TDFh4zMdPgFaN4zW3tctZT8rHNup6FyMrSWbcBZN6ELBRdfB9As6PIsXt4
sIjAxs1sis2kEkju/Z6119f4wIcpu7mkvCJKHd2MSA5XAUeLRaxfIHJK2r2S6h5J
MbORw7jh3bTw4zw4df6wwnr2BMVaMBz2/UtKp1nUBJ/ok/aaE4zhYQmxQTE7Zd/s
rZo9zU9BjXxC9vbCqdcZ5Gkws3z8NrHsYlzKCyHTZvcGasgdCBzRE9ibisMH43u4
pvctLyT4kV+LNnzcuepIvbrSr87jXg/Ox9XySqMiyiT51p8wXfbRlHQqaI79lNNe
LD+TjrwZH5zFMpqrM3vza7+G2nji1M7WoKmcRWfEtk3BEWD4/yQ6q1OMn78biuhw
yKHVlmrLn9tqAHuZGejuBSc7xOCA83gIOyZ7o/kd2mY3byRXD1R+vrZ3KIp0PAXn
5DxAAwbBbM76X5z8tubT9nkkRlRb9kbFyNxdeVCqY7zrfTzcIekxWMveoFcaA5Uh
+7C0kTTjuqjZM4rGiEgNo9rkRH8UyBBPeQ5aHqi6NpZtsOFRFnaYWjipHwNbGcki
ZSe29z6/GhI5w3fP/otLYIbIRg7cEOj8sobnZLQzb2lcPGWf1ehbo+WIlRTtBSpE
Ocu2N65GSLKhcwniiYn/TtiK+d2SE8pq5miNom6QJFeArb7JKV0fZMpC3ADNuo+9
P3UkCO9uPu35C+qEMebvWtE4p3ZE/3aHMtojovGyfPJ28KF4oQqzSi1cg0jbyls3
p+vevwWa81wE9F0IKEDRzpcn4IwJo8XrcFuXYrcSk63Q+/qc00Q9DOputqBs0y+h
aF/dA2oIWasj3+QqUDqD+CAh7erbx8VO4uwf7K7fgwt12bW5+hYXSe2fKQYeYqE3
2exllKNAgS82OOWG3TOzA2ociyk/rRs40y2rhityvaqlzYhtxLdvUh8k4PC2emCW
vBj81O3O+Mri9KNQ1ojmi3+yFABI6WSox2cDX2bCLXJhUo1o1r3fVCzhjGxNor+A
lKe6jIWvYAVCX8YDTTogdO/lZjV6gFLSsVjSNCtvBSYqf5eL2QkkjuFztHIsZRJM
bYl2dUk9YBVzh0/+Fyx+SNWVizxIQU/J6x8p6o1wc9kf34XzlBd5REYiMnat7MPF
bY1M46WR3hLArYa/Sg+P1Xda8PrUE7xCdiV80NjwQvRuwu5i7G4r6Zh4dw/AQwQV
9o+dzHakXNYOEADBzKHkDRFhMTPazQYyXOmBXeHYXk+wAg9ml74darEWnO6nKjA+
1TXJMb1a4OFyXG/XhV9Lh4CJvF1f/TMR5kkdZY1jvVz2MYj6BU/1dkoGLzkVTY9w
miA69I7WWAdUY62biwxaPMzOMSGX0IXtCbtnodStMG0RCN9ORsCRIp6M0nJrTA7I
Y1b6vb0scELr0TotQWF3Sx4JISziLrJT2UCRwjBxV1yh1kib6Y7uN6qSQG0280Mm
9NfAtyobwuN6Xi6OLDz4ECtEMIWYUZZ081dIQPNSEAN7k8POFU/JvNFnEL4CcZJ4
0aYTdOGNvUjXoL9FC8kUcVfRg+tQfFkkM6VApRsIQFajtNTsa4/2j0pPGBBItUPi
Mep0I8a4JkyJhaNPgWqiVDeVd0Q0/vzFZ540Xq1nfRpnUVJoIKgl7Ii7Qkl9pgYC
wXi/nHU4NaT2ynJ6gex5pvB4aXCd8Mfv4qxvRrg03GV+GdgZVyrEfV9HJNmhOBSL
5naC6aGBymBbg7e3JzLLggJwnoElB04aYxzEp1etU6wbdsn6/ir1LR0unhb8ErmS
dGEmYwhp0wW7gBh0dAYtQGSM1TQjbw6Cw/uBZwfgwKnGQbXGL06rQWtiscjCF+KF
ZyxobVwC+c0+rO6DJbQBmbZ9juXRDXAO1Eav+KweGRufXgcZv3E4Y9hzFynr4tAo
6yQhFhPsAODmq5eS3yoiJtJRUqOAax1EQF4x+U6BtqoSsMKXMlhF6NpcaTTz8Dn+
w75qMb22f57/CdsXlIY3F/Mz9pMWlsD4kwkoWZZ8/n2+Jsgv4f+BFSiInTDFf1OU
IIWgNFkJ3o3QWxolx7m4j9KSHeSzhe86fMN4/vLDoy/pJP8G3xMPSpLwjM/Ky8LT
0xQ7oQydDy6nEYhcoGVlFbQyM4TOfNKq3W88ZF9s11nAhm2AiMyKgxyT/2gSw9OY
DN+RJZHOh5EOgPnUR1xe654N2XTS7BUXd8y1aFb5/2E8s9jiS+rQON34kxmuiAvs
tH2nuEFLv+6R6wmRY7RLYs9Ki48HaVJJFNvhpFnwQs/FIVezxKOjXVFH1hbHlH5l
ugyZQQV6KPhVZbf85L+QVKc+J5WKtcR2as1BRnO0qEfoWbhdHFgdUiMri2z1MEgE
g+Cmz1zFcZufyPvF2gTrtvA5ewjRIApBbyr1w8ubxaFfJ6I/Ti9f2g95MFuiQp4s
1adrQ2jK8+/I43f+LQ+Ivqxz3tuJjtSmK5G533qUiHClPj0oOjLt8+Jii+65u76N
9eXCHESVyUn3GlE5UgrpK0h/+3ytuebWqof7zC7U00Qai4M5dz/PmciKsXz4Csth
yJN46G4Fg5uM4kZ/UstiKORy4/ZlekRrh+fXEz9erJj+lMd24voxUovsKbbC+Iid
fPhyzLRz2h7b51t6vUeHyIu+GKRXqH9LPcdkHLIZEoR6qaEubo+2ws4GA/jZPwtZ
7QS/KIycidmDYWSm4RxS8MZ26ToDdNVCb368ccVltsj12IV0mHfsXoU7AWsNDtyX
dAUnoJzybw5MVyu3+9tYucpxLFHlOO5Mi2f/+o6TiXnf4ndtRKD/QqJ1tGdtvyvz
rCgvTKK8jvAe40WwofqJNxDlaFFzWp/9lEcmCWXF/f4AjjwZ1Iwx/nKLua1M3E1U
dqpGFTjjD44NYIA+sJOInR3lQ7phiKY1JOlWxmj+p8iuSI8OE/+yYlWrh75rAosw
sKXJMhg5ZHnplfuvksF28BZQ36a+k+PASoV/OK+P3w8/F6uQErq14NQiGsdOAe5S
pQc6LjhkH/Vn/1l9cwtNP3d7ulbO35cqprRrqzXP3Zekw/xoDi40vfaghzD+/tsr
DyjJDG+AM+IYVfS5oYGpCHwLgzBwCsuGGQDrZXFEvh+TTA1ri6sY8AtmJttCqk3Y
nRCivTG35Yb7yCxWWe+Xx5bgwB+OEgwIfKlL8exhqQsxeXJEjA8Vb9MVQif9BxF6
MfVYLp3RyBhSuWkJ+gltHbsNo8BUe/zI7rGuQgWDuXP/JFDezHUBHQRB8sznX4AP
AkeUtttos2o8zIp+EuY51tTyjCNnctkn0akdDf7miK5Hwfdg9UNIdZQpM9yAWf6F
/QWlgGLcT/cqnXWHprVQqey/S7rh2diWX3X543TVZqdqWdMqBzqhPJDgo5LoxMo9
xhtIZuUDBv1uSI/GljjMLlGNlS4dDxc8FO3Pxsl+iSigZYvwJY4ZWsz0AML+tM+d
nSQyqJu1pDN4G/VnV/B1PIA0/RmGndniJbuN+gZ0tc6wEdBBifBCsMy3UfiLTqFx
igGQDXteJSdmm8JftscI2FQcmja3sIYJoPr4mPZV5RAKMtXteHorumEkuaHKtV3U
wN+AkyUVhqk5OGs+sXJFOHPbEEnyCP2CTjYplovs5gmmRV40XoSXKzD9ViBEtDaK
uUn/UPK2w+sG9OkZVCovx/GL1WU07ETpGAgdc15+tglrI0qvoFU+W62gx4hk0f3Y
fwSiyCu2An9CfdqiTRhv1F2Jcaqyk5CjMgFT4yOYNwTo5KfzsivZ1cg1UAYvqQjp
ZqRKx8n4zucZxXM1jg00FMXly5W8uvZejiNJ9nYGIZ2gcrz3VH4DnKr+QhBAEYNt
s7eDQGD7R4ApZzUhHut9O0j2BEB/pq/NXK0yPVy2/4JcpAnDT6k7UqJ+Kwzax6eH
IsiVxETN0T6DeGeNH85jJv3TQsz+bLfHCIbJlzn4o7JLcRoK8SeKK7WZPHVXle4I
PmaSUR+MZX56E17Z2c9fjZLuZIS5TKTzdmCsnXmt9IFfCSU4cxirfHSJhAj84MT8
JGuFVWr/hthHZ4Rfqkug/+X2PzUQ989bR/ZiLhCX1ws2NDEfxn2PS9zMDSxl7FQT
OxW7wULa/zdKA3KrPpHWrMD4jK/MvNMqJgWQGGhHMavZVm+GN1JiJ2WVcXZNfkjj
sXWYG8IiL7tkiejqk3QNfQWek7FtkMT9twx+nAmF5FQuU5gNIyHmWdGro/U/A+1y
cEbS905sxW6wMcNweeMLaAigBrUY/Z8+YUOhGJDBayVevSwobtEh9skPeiFEMYid
b/dqhkkq1ksYr+KYbWLj6egRfhW60JDENwqNbmX3O9j1D3I0Vdp1b+UVV3Pp7bC7
Ew+7VDlJ66E1LKC4ODeEW0I2pFrAShqZTeFBtmNqm6C2a1ZB8xc9e131kK1fXaac
Znq0dKiWQ/9s0JYrwhkyPC3IxEOSl083NDPPBrYT5i3w/+rtARHoM3HFP907Blgq
RO6jc2MZk2zbst9bRG9bRhgO8z4BzFFnEY/0ADtNKzqaWBgJSvddmdPINQA5pQgp
dFu47dtN6ChZKrf2tjt0NA+totJ6W9+9n/lSS5xt9NtnbXBoNTYI7vu6j3x9GcAL
D5giyQCLAuIEK4fCrAJKVZ9DW0/c+zR2BUjIZnjinM9b/iThCQJU1j2w3gN8Bns+
LaK8VCN3FIWkhYNn7ziYXF1+0JZNiVZo+DqsjeuV3fHwxbhqSvsVZYd09V7QZ3zs
gUkB/exj5Rd1tOHc51rLO8JDtFdWIcKil6KHaiZFD6PhY+xw5gnsrxnhghEkVssD
6WUTx4UgDtn585DszWwSoPBZ5iS1QGlfoeUhTt3pzfPWDJ+23st+3Tzt1M6ZDNyy
lhjP8CHEiIHvXABiVMRuq/nEMzVNuVOcEvQd4LE+we7hhPRbHb6JGsR52nrLNfP1
Jx+jLjfLPjQbjkPsMqbP+/AF9grD5T/aW0cDSpiZ/H2W0bAtgKDyRXx/nXEA70xu
OL/f6NDOa0ab7MJZvARhQkA2M1ytWJBoRdF+b2isUx38qWUhe6EF97m7vtSkPhil
f+ST8yeqmatnkaYFDbSbOsknlFp/LpKBdfSHfPCCEK8AV+XoD75jARX+Fx+XVqq2
fxn6vfi49H6mt8WFhs0FCAMzY4jLhE9yRb+ShnE4qVX0VEECnALm9y62CepOEGzj
DuhFv/tWUYDpY932rok+hITV1mLiLTziECsrBmp9+k6iFxc5gCocyARR+r5uvM8V
WrQaSMzCXcmhlFOccU4ftthvnlOOf98vabyq28UiZiws60CDjTaSJq09ISlOs8W7
AZM+YlMO9f3aMJ7z/Lg3asHrvJ3eTNYA0vhAcqnMgAwu77mA7An5s6z6pp6ICC9A
ycUqOZWLw7hIU/vyVg0Ok9wPS1C/BWb4en/9fUPGrbe2Yu8T//HMnwHUQVLvQNGE
iS+Zj8TuXwmZ6iGags7itB9ohzCDU/oJONT6foLtMARcHvdNWjCpsBi/H7Izubgd
V5SBcJbXjYqE1vseQCMyAgYVPUsCBTjeezVy6126fFZ4s6BFe6YdlvPsMhnje4aU
2+eKoHn+pBP2le0gZ7ZoquzxkkPDhla+TnBfzs3cTjSW2UK+rDbNLKjFAj1Hu8qA
wR254uffmk5joYiYLgo+TCkhhe5UUfIZvYPNkWgJHxVHAjM1oCQU3sNU0CnLWg+I
Bn2Xq/sE5/eA6Qna7XNO/HDOXIFYrk5BBIuNzVAEjBtLn2u/n1KEPK3iFbksHleb
6C5M1PhvBI05509hhMheOKaVK94eRyerItFzRTrEA4dpwQAuDLcQVPpeUK29jmt2
YMRaOwq04SQ7ch396Quz3RXTT9qf0ysL3lyqtN6TKGr8rr0ZS25izB9wao3a+2kb
ny3xVkVlrVo2FI4jjMnSmfRnv2ZVPsmSjB34/AhDF9Stj+HWbL++SfsxcJzrwY0X
Lasoo93wZU0q1sMVI+lF4tCTmQCZsnBS7nyFYbYX37jlKzR3LDUsV3TdAKwKnkKj
Tgypid+wSSB7/h4nWRgdjz+4hlFZw62Mk93NeTi7fGqMskCx52n7umFO2nsuBCIA
CwZHLaL9+Qk+vvSk8e2wyU0Gz3q4mFdv0/jcqmPTyVoiUww4zv3+K4xB0H9BWzu0
AURp6duBAx1s6wV4guFtrOFnFlB+ZKfki4suspHzfLkCGMLgqqokE+0vNekvWjs0
qgjxFEmTfAAYOGk78+SNVVt/EIPXifz5O/BFF4ueBF7ufhBS2e+C/BRry/6rsJk4
fF7gCd/8hS/wtAOYceu8ruZvRoxET+IjElaZcrqJ6p3pUcqcJPBYgQoDd5B0QCbu
2pAUoGw/uc3qHDsC3Ps75xLZUqFjdmrifX/ja2k0sGP70U8NPbWkuDqVrPG1tckq
49Ctq+f20bbdV6FXVgNBqEskUoKgbNNrZ+m8RzUIIvT18lL9nnxdb0P/5dATzcKE
kCfBCVUSVXuB/RmAIgpktT34s6z+uQxG44XfFBBrP37eud2PlPGZQ6yYGFfPZ1bI
1za3AU0aWWTqJ4Y/XmYluVItACQfNVELsDjwc/DZm7UCb74fWqgOciXjTxRN2Rbw
4SudpANm9+qYCy4wTcxFeHHYzRV6xihYu0T49VyEsYmGpSVPYN6U7G1cSdHXf7G5
qrwCkHWP2EZ487RZGvnazZ76gp3zxhQ8V+//C9z8zL4vGUiMr3iCUhy8Uw9b0Hx0
l9nJBxL1B6BBhsEbpok3fAcFY0c8TLFGXFg6/erkQaWktNzAoqW4roJL+gQ3E2p9
fedIdwZJ7C17Itu4nT2MUzDEiIw/hCAiL298Noc+IAR+1qKTYdEPvcoCCgEM9dTi
FwKZEBU4HsbeDnY8Mk41wuKNa5ph1epE83m8DEJbPKMngbc1NdlU96q5UAU0SuWo
Fyf9XqZntmO+d0GowLvnb7gwjLBedw59pH/rw25ErrwS0O6eFLKW4hYoG9rsZg0g
4x90V2XGi2z+XZfwdwgXDR56yqLtfFLQ5X0/WDZmnsauD2KdzP6DZhIvTJx7dkXt
DZVO/UZkuLcq2Jnly90X+n1OJgro0mQ1lXCkGwaVy0evPQxZMdwwEHhggDnqGWZy
83Ihfy+6RgbleCG53T0+KJ+HQI1hTj5RvUEMnI+4q0cbTF7P3zwUW0lcWtu7JVhY
JUd/etj5s95v/TRY9uOHFgTQncf6FSV0BAOZtYIORf21TmRg1CyzBtEq5X4nt4Du
neSyIPccXtG0AaCt6vWbcVp8zKvHNnLOMf+jzVV808Zr72f5B2Kj6jf5ZsI4vvhg
MkWdIL6b8KO/4A8H2DUprxrCHXq3UQRHfXE8ihAhJOSDT1WlB0Gyn+47YFmnuwRL
w646ezdQHSRey8Q5RDhsANb8pM6H3bBCn4dE/lhRI+UqvsGppmS1ZtKbfruxlJqv
GKaKsGJG1rNzZa4f9/6hN3lqCvAc8Yp+ncX0rx2ufHP5ClMhz9kR5pFnE5Ze2DmH
47256SBa2MiJIu4uy/HivMjFs4ylKEBKToIw79IfFYnt7IqJ2EvJ1i8wwVKzVUSF
FGcIWqxPUFN5SdituDDrCtvW792eOcp9mOoeKhdFCO9HW6DRNCRjvEdNhaeh5PKa
c12EC+RQ7inPm3XGoD7X5R1mlWrYfOmUZKgJ72H5zFXSOX2yfKN4TadXnWn5swQX
JuP6OvTuksynWC8cICDf9/8WzSmVZ+zL7ZaiG5QY2cADfT+tIQR3nQgR9JBBjMKV
tzhwA4b046GqI1+f0bT+hNwTeNZZQzcayd+Cv925Cyv/VO9z8fcPFQAY92eBuXX2
K5IolXtiK2fp/KtP0Zp7THbUwc291KQO5nKtVZ4ylktsE+5s7+cmkw3NoaqJaC+4
X53LEb3zklkCoRFYE6y3i1QPdUOJHcnNuZWKME5DjJ4greRPrzhWfNzdQwv1TfK6
AbIO96B10ilKx6rUOHhQHTMnJoJ59vqwV3dr88A2HoXP9Qc67Ir2gM4uymmLUR+T
eltz13av//V2Oa5bUp4ZYpH6pmBdIOZ+n26DfPLCjTMiigAw0VOI4PuAbKB+mre6
mNwRl/JayQtqOT+JjkqeKj7qBG69crqt/dn2aVoV+1Y5WUuYGQKWdIGbL+sX2OU0
O7XaVCYjziEMBX7CWkW//TNTnMOppG1Es4PORIS+xWOQQzoKw1yFyZPgNbamwGxu
ib+Vo75TOpdlBWgDiqqJVmgj6DVmi0VMDeJLo7BL5wJ34F9u4Q6q6mNWOEP9g5DB
Cp6UxIspX01PI9b56zm8vv3qFP30ocZC2JoDNrxMMyK7Ckur35+2ss1PN68sMouj
NpAF2vHApdCemshmbZNl37uvNmGFPj8p78+PplfCgxo4yjgMMYcI/2x1SjIipvvY
yBt2eIB7sbkkgARWTz+f0h9Kw2DRrWxGHVPCMmamPkflgPlVOAf2CvpTFMnZP+34
uj7zVQYsnM8MCOtnHx7p5c+5I6NNJipaNl8enMqJg9nMuz5JdukmalkkQjaWFg7n
avH0IGw0nXCU3iF8W/qUl6gxdY80dRrTcgyWvU6IBdxTcnP+hZp8Epe8nQy50cvn
o1y469TFeb9mCriMoFHqgm9pBpeg/saRmNrexIwxSayleQ5YqmOeGz3brUePYNol
1f0sM4MhO0YUzBVIfOCIVcw89JROl3u2Au668zLQfrY6S03e8OHyZy8N864D5l3Y
WUAPaoBtX3rtcSCBBEDvyr+L7o7/lLwVQT+f8Ef7T+ne8COrBQfR4OIk82Ac+Sw+
oqd36AX/oMSf9luk0UqkBvcsqlRoGHEEyD1hItM+qmHC96+bMyBjLWsbCQ2jT4Ax
Z+qUcnk4MqcV91/Wwj6p4+kQ4/O9Em5uHckVW+RUigOzztXAD9rBGeB+I+QSf13r
Pt0GEaFgTOd+/hSg7QnwPhHknXrfs5HWxlLs/wx4RIeXL4ehrgFHYgWLXZme//A6
qB/lgxVHC9/A0tIOeo8TPc2gkd1WZQQeQKfGGqYrCD9KwWBKdFzZVo4qbsj+FxvG
yfnuShHLwL7KKrQb8S73xNK2I1Ng/40HAW3Wd9kcNJB6BP68EqcUtzhKAbTE5ooT
sToedj21ASdedmVu5knbaXBuQfwULZ8Jsc2ZLmtYHbt+VTGQsC32aTTJjfSi0Lcr
9O0dhNmfW1zHO3SBBwwAFoojOFId4JqBE/GoIHrckbu/Bh+/AVTr6LVEhcP3O5wK
LL6I5e2t7GOKqORDqTzxSLWansOpax5Cp0JvBa8Nn0xsH2m7OVUqSt5D6JBa2dG0
pi8wzkg7VbiVepN2VQTWRiuSAReDOG9uur3ykrAH9p2MUImVeO1RjprBaRHcoRjn
gwTErMNJQnzVpvgolJfFCEVmreqLL/XzuQSe8ZeysDQxPX7gwrGMWPmTx8l3ZuRV
b0zmpC9SHPsrDnwUko8NjZ34AJeZi8FhdD9TLCgH1ojGQYs4leKpWRdH29ZFZdbz
SYFTULJ50DXA6stT+aIENaJNlKXcHMHd7x8Q6NZkolVXfcH89oHCISAyE9/cDR1E
wRZtVSSEa1JAVagB5B0K+oyoH7l9aiKbIT2+DdYlTZ5am93stzIXiDvM559iHxc5
bmrKc/ENDxu6C+fAfCH14ofL490fCC/j14AtJjbui55DALcCpvKccOeCzr9c/DXY
ITjycEUNR9DFt+Yroyx+amxMK+9ybfZh4eTK0/CnlotUfc+IEKQM8dm7p91SvgKq
cpo5+MOxUZI8JDscfBqnu5OHidXFS+vQJBRv8gzszwbH1S2hn//fnEEcVLOrjFEQ
FeLuqZL+K6PHa3fghnqLTYmZvWZaxC/GewaldFef0lCRi1hTkhBiSVN4wWGCZdUL
XWOjW2ubPcmm+lbbwwW/RNC8o0smp+PNp71xqS4zgYtMsQU9xr7GhpQL+z7sCgAU
DVjrKnwfrxVtKAw844czVhDXmo95hWI6FjPAQyDVzqthsHJmMUqAeuJx9pdrTiI1
7xhjaZgOn5zjlo6K2hfBFZXMDJjcVyAlfpYVVJC1A9j3JZ2OrJtBChsK5j/e6X0k
tSbYLcMW+Gj6IopYjTN6MBaZd2Ty7+ykrZ6ntt2UaqKuj6RSHWDAzXQwGQ4V2ROF
Cvf5AEN8g0WZppuxdQOqIzYeiPDV7VM+DClQ2sw+N1MA0GJ/BG2aVzQyNOe1yzIs
AAr1N0H+GB7uSVNmXG9KaowgMfwBfBgw5R3U+eDeYc4Y33w1PG7CgFDlR/5CTX3G
eg7IYHn5NuFs16+i3tF3d3/qyJnegagg4f3XRS0m9m6WgJxePd02p50e1u835qHG
uIYU39WjAl6W1T7oWBURAzqIw4i4Qrmaud/YdfIhRBGAkwUz64IkNQhXxGA4AygH
bWbN6mRoeroGbpFpF4c+FJbqUBsApxlazi6fLTvKIcnl2m1MOXCE7wuff2c404Hn
3/jBhkGUrepuB4zCZmsCfpbO2AJowu/MTYYKuB0TVppEsvY1e2wIVheK2x1N2guT
tjYD/CjBZ4NDwO1kNGaNiTy2Qg5AE00KrbUtjxv3Jp3Nk7UAaoB+UuXv6nfmLavs
MMx30kCrIxG1FKuiyFRpqVpOq7bMfsnsmiT8PA5JH4m2DyN2QcYx5rK6bp13hAjO
Sdkp5LiYgyF3SxNQ9EdmJZJNFxy+tQWlqj32FF+qYmXJUR3Ev2N3vbYYscddCogF
OCbKS9arObrO8k9HngOPRMcO3MVDyDe6+ChOcE/+O2srdjrz+yQQwf6qR2et+004
eNph8xWae588LwX4KkTBUOXFSnrnE1vX/r/O/Cp2RkSuEvjEn3OABARhbjUoYhCg
qINKIujiqhQOT07LIholwHZeZAOYvzdRBKxEGKToErmbfn4EqTKEImqYpSz/Zy3q
/+T8v8RVEVEHZExemmzcodss7XXfqYjPbcQD4cauKvixk9eTS7wYHgSDTyJhr07a
ojpuxf97AhOML49Oc/EDXIrbMOC41T19lCjmz91Dldtyfy+cHX0xUKaflPKXG9Bg
cKUHDpipW55aQiurap5gx4b6VUO6ejjms8Zbqx9VLTTFS8XSlQQE2S3DEQunNoZm
DRVEqObCOah4a4SbwFOZD8UIk99auRho3AxitRwwgIIyDYonk5EB/MgF0TS468pC
7OP9BZ/ysd4CbY1bXecYpw7PF7Wb7DuKUl8yJvzN+1Z/j/Tdq11AjYlw9RlqdWZR
J2GjPulxXWq7/hyLu80nYC+6toq8CTIvW3Jh5lDVdMBdncyx/9fJ7SDsRHIgMwKk
WbTPKTvagnABu8aq3ff8Id8/SUVJ1N3OQGWBEW/X91QdJ2tk8Da2k1PTZcgWcqbB
2Yo5HNT7xLcWgeorBK5uJ+y/pzKSytLdCghTRfDzBlfCnAHq7vAtusK6d5xjDlDU
NT6ZzAUClCif1eI34tXtdFiT+FvKRqq3Rh8ifPm9m1ucIRlMm2jV8huar99F7xEc
0AnKtV48NoauL5NZ0gV2K8Xi71RXczAKmqIeaV8u/TXcOkfYKLrwpC8z/W3TmC/c
MPDitmkSBDcokfIQUAJRH3Mlb2Er2rjcRiJwuraK3QyCaDawRtcfRB3Ea1DonFv5
0aHNiToYjx1oCzm6/sOHt8y1Cxlk8bZ1ITf3Is+6RbfPMZxSXVEzfLFtcn3uwiYq
Tllx5taaZp+woa9TOKcTQO1MtnbpTcrUofhthSWWafplHrrPlvbX+peJv668EA/d
Dgz0wY19rvsr2EmCPELToyBp7GViW6FTxinrqFVyvt1hT7QNi/vPjBf5vo7tcUOQ
eMFlObfwVN9qim0rpLGhJuebZkEyNQ3JEZiOmiTI7MlkXzWGFSTF7XNApmMiP6tH
iTcitY2dPoLrkODe0thrW7QSb53P8A6S8ujLW6FwxAW2kVc5UMZnMM72U7b8WUBo
A+hdnjF5n4dOgCeUXEsNJqmJavRefgLINZalTK4TQYTnFZfRKnWjU4DLIssSc7Hr
/xHVpqivAqo4G4trWS5EyhYnvc44UHsEmi/+BqxCnxWPAvhvvTPT8X2rXmWpRu3o
RA+1Gl2ecN7PU4mCNqwL3ldm3D/S7x7vv/4VIUK0firqOMekhMrjJLypM1/Pip/s
Ba1r+a/cDQyg7ZFXxU5DfxD5bo0uaJJzeL/bLsrJmAhDZVX5H7KCQoRf94Dl0gI9
KP9DefrIUbVVuZSbEawKtjv6eH8LFNo5qIVSRkUATDLdB79JXK3bzYSXMmtITGNd
zPxAKgw/MZkFhDGBqFA/sZzvLnsK6RX0BlMQq4X/ymi0rPsJvCtAREHg2A5VHbnl
AU/Bm9wx7P2xhDlXQzLjT+orkiPKPFlkYtoEJop0XXSx6tnl02WTRNC/dHuNblyB
ozLwXdHRgFNwZ1AgMAWBTChAaPdJC4WPNfdgCia1bDUTcQfASVACcaWB987ts3oJ
lhgMhS6YRNg7f3mncE3uOviq3C2GRkMB7QU/Okprq6BYe3Zsjd5yEnT0lJDqia4g
jRdft0iBBaStGAHxsf1X+PngHzt5oeVDvDTadi12buarp5a2O4aX9fx1qzBIYZx9
tVt+1UdUUB+C6YuB2tszpqWnyga+aMg+IqbHu1LJTuD79w+Y7A+OxLJgFAN8YVow
XBty8qV51NVvdIQVDqOfDg0zQthZZ7C+ua84+nVQ4USQ7ckA/KzygNb+1Vh4Wult
NW9QdkVF1ULh0/9OEs1YbfrXhjgLgVDhRpF9crzsvN8ZmcZbjBIgGn/EqqJiJi0C
gSq5OJU1VD3kFA6P0LbY7AX9YWmbtagEZUcjFuh/tFbLthVuQAyKNeXSpnp7STbp
hxtmqpoX/vScpkjlb4jftcHcsyNy2mGdQrYRsyb2gj7AtYTmLx9+WwMYi3rrYdkg
gsqhqVe3J/f5nBAaua5AXOsMXqnEAe+455vnRU/zsFzseeyQYnFvQYlvGQawwOCL
Tr4p6q72DKhxM92jAMCZ3FnSZSDTugjey7HFB1KkgG8ZSMZ7qhL2UONCspcCcHXW
wvlJJv9GuFwbbPJwVaosB45ekAw2UVp8U7NoVxdpffVdvZNtVOWmXvpO0H7VwMR0
QLWE2q47qorUEGcrYghEVPJEF6Bad/q8pUMKu4dBBvlIJPdpS65p8rb70+Ri5O74
VH9Mb3mrTcLAKCyCVSSjZR5OVW0PO5BZjo+1d1jaG775WPPO50zdt8s9sWj4az1f
GvrY6hZLwUJoxCBxtudWuK4EnLmZoIDLobWDU8foOkabeI0sgormtTfTRvhny8ZA
R7WIP9qNutN87kxJWSnHPNuHxSDFfG568Dsbqs7WsXGcTd5t1tLOvgs2wyPfb2To
15oY/df1lFD0KsXks3k09r66P1o+am8gS9/0ZYF2Yg9ePJ4Am8QsjGrHjb2plwh9
018ee1SZRzRxB8FvKkFgL4gwTBCTgaMe+BDvZeRXb3BpJv6CUiOeQObI1ay+N1D8
DVN+RDMit4SQW9ZksR0WjRbai7mUzNRq8bWeIyNItr29mzaitB3ryI8ysmANSkju
drbOstYcpj+aoZhjLNr58ZQoe8RBoryuj+Qcp3Nwy6WHQjIyLjIgjusaVC9PGfS6
5oWsLddT9BiUJp2CM6NDPFEWxQ8QVvULZIyOZJ5URMsiAQOrs/ILCJNxuL1Eb0nl
9c9DZ4MzJKoa5WhZKzsa6eKc+e+uyx+H9PFRM61z3SlYKW2xPJzdMkI2YtLmwOH9
ee7ERzbj3rcnXu90b38fw1KUCOXyP1nQPglptGrR77zkpztLNlZYNhsSM2aRaemR
kGMp2ixXlhWzemjGRtwmZ6t+JWe7YCWcIPvunWFMIH6IwDmf26o60W4B8zyaL+03
SFpJDDVtchhu6D17K4pI0AOJtFUu9sUmS9pm4/N02yMDrxEwx5LigdfDPjaITSna
9LBIKeWbwPQ5+ZwpPtLAfe820ENONUyTMcH1KSYwAQwdfYuxqU7EnQ4ja+6/5T3d
0H/IBG9gUnrf3r1vXO2ltGrHGICdF2vc7hTehBp5OB+4+fJ35jiSPrdAg6NJ5PT1
58TngvuC6yjOvSZ8GkHLn0wC0FajtMZ2ORjYxFUJcBkfYANq7LI2NLy7lKjywax0
oiwOH1DH+HP79ZGtpnjLXbam1blr41TmrLV/n/2Qs+zWdicosAGv2J2+RiMZaIZQ
xYy+SuDmRVxelxFR2muFG5e3RZln9UqGhr5U3kxM9QZ3GHwmUs12oCcAmd+iCWvw
SJ1IX7JUDuyfCc+ziDgPQfxikRxj2kVKeqbbNx49swyqIslYlGP0mD4rpY/bW7FX
+ZQaJPxV5/enop8fpnWo2BzUKlvFkPSfvw0pVZwpdY3Ddodsa4/BIS0d/U8Nraso
hp4b/66nW3tPaQY57vpVSfmGOdxpqC5ewl7nVZzONU4K7Ps2ihMUkTvzIQekl5xx
jxNaRhmGk6WxTfC7OFso+BZ9WCcITitF7GjEFlS0ldi/yDu7MPE9ZMkWUmL+9RAD
QZPl8DhJHjZi2bRURxJksly8GH8JZKeA9VF2WiFKFF13WAhqwvIrQrWDQrVMKXns
rO5ZtgH2qI4qvRyECjGkNdBHsNKAmaSYHjjg3v1yCzU1tGqkFQPJoIghtl440U7F
TKyiZj43jY9aiSWy8dVOj5ZIbcsl208vkJu1dtw9Ur6hJoEWaWUIBMi/6XgvZX22
4YGzuF2rak4wU05OCLGVsBCcNZaTifSvaUsp3i30Kdq956K1KaKVBvAiT79Q8YoB
7vwuMyA36ecwVFiHD+m8+5Y1BsHkNYuE8dpCD24oJcfSVkRu89W8yeAEf1PwXP/A
pZae8ItSODraXpxGx7URDVpGISSVCOjDsXofi9QMS1qF2xtv7+zUEuHZ7ngkdQQC
bLmYVqiX7EeHy4zMLpwz13L2p7Y+3ZPN1gnga2u0ot6Wwhd/wM/7uaPLbqwmoFUL
xNpystHMdiTcmDnkkikH7thgyZerTUYSRQ/0I95VxD4qW10Lp8VVHGuMH9qRQqdX
yoUJadCvviI9r68Wu17TIbGeBVPobOwvKpFy3x6zNQvUvOh6pwAUCvJXzbbipTu6
Dic/X33uHrrBJo63RRDd60aCBAfYET5i47sAXXw7cWKF0e9Qsb6kn1e51b1/x+ss
F0awE7jJ6bBYB+ticKRxuTQ/7nA2QjacJ2zOEOHbXclU9Us62WGrzVcpIwPA3nyS
COECSZhnTUB39RHXamxXCqpKcNiG+NVakLHZVNY0KtKPdP4Ms63crzef6eUoSD40
Y52zYmongKnHe+dKGacjajWXYfhma3umPWKu3qgrNfhkgRAYhi5v2XdhZ764QgF3
q3rzExfrCSep65PlXGdJ7J0g98MlacfepzhngZBD4zkns3nBn+WKYLtaYPmxoE9G
M+v+cbE5ENVCjACMkUIlOqJPNhLy/pI3pcmGF1d31Mnb2umVY9anvkYCm5kE6eyt
6s9BR8GGuO+KXFBkPnhltRiZK66O8pJzGILBaeTCbXMcCs9ETxyuqjxzLw2rVMKo
28NomcCG4cLHYB2OzJO8f0faEIonBqEwlKz1EKQpoSY084UFWD9s3qPM1mgFvUYW
FgitUbWh7feYW7pnHDq5p+5n0Q6yfE3TFupUomcECxjUpHS13OnxAZaoMCO6c48D
6jz+xnsRocUmUl3r+JkVFT/aXagLPdL31l+ACIIuWBiz43SV3Zpr/oYbgJGgk2DY
aTfJjqdZQSfRttsm37YSfrTI4pUlfv8MvL594jEmihhWC7F2ZiCTCOyE/uO7NRBd
0a2SE/0LLBKTux1xp81947inx8eS/k/X6zX5MnErUwPH6EQdMsuUEiUEdeMsvXls
YSzAo3R7yPpMCNAPWGDlAF7upx1/n1O/W9MmNWTc1pqY4gBUgwelw/24MYPC1V9m
j45NtXgkz30KYv7gVu5/dBxp5obZLt0JDQ6aGXK8n+DCqqOM7xZWGqJy6TPUrUUd
lx130+OaoeZeAHZHdQVe3l0n7UVi9QIAbTFvjbfxsByfqUucOOMGnnWPWZaPZWaA
jyxUSwAQIiMGk9OmXUiRsYNrUA+Oj+BjiD8ynq5lEvu2MUuNxGNgWocpKZTaPknA
LWP93MG/TLHNF2zcqWBMi20job7My48Z4jBkgqWbQXAiMVOYefHKuPW2VTWp187M
n75qmq/OtUGNwTUS9IJ+l58vnVaJ+Tl+d+ebrZgrlOI1MNM3B9FgxuBkNzH/DqRf
gBEDZmqm6dXZzvenBI5ZNQRXE/zL7BHdkDgBGTnQLsc0NTdVLdTgQHc4gdbMmOAF
pEUBC5DPxjdPwqdNOWWhlfHGvH3LhQkaU8NmgKCA7D1kf9SXWomUgKC3sAfKFEkC
A94CgTNRc+SMC/ABgeyteoTh7oXYx/JNoAGsTYJwlAxFyNrX3hZuRDxkzmF12Obi
/Urkg2MmEcCx2aGPJpeUoCBm2qdTNVC4JWVYMLrDtctA+poa6r7SVu8fkvPhDObz
OjLVgONueUvNWdsPuRJv+wD/9/Ptd+CEyzo0vrM1FBwD1yqmshQejl8DXrv0m4Lb
OePmS3lumgI5Hf0aYT5+8Y6cXbEBmZTLQgQMsGl6hoHKP0Gr1Oqh0LxCOZryNZGc
qVid4ZYfWKZCJ6xvoWLCIlN3Bb97NCyx7Txl5CjurLYSWvBtJGW8NfLDK0RzriaW
/+6BVNK47h9uBXzFfHIf382gE9bHmNyQLU3DGrPBY5fxx9IjP1kzokyLXm2EqmGy
r3rbaLIUAQX2ju38U49c7kItlY4thzPA4aCCxryKbIBJKhRwQPG8B4+p+OVr9uKN
P648/cOtzCcgSHxF3kd9wVKAGeQsTbf2X6bNbGs1eZbs+0v2mozIN1SXFkMLXkoD
pKzFAo6VlUoyT/Xpp9TWxiQathtvPRnufTKVjgVgxwVSfkKnMHrYEz+K9DzJErbr
ctkIhT9lMU6uACjgbgnT5Q+67K2hzE/cqWOPu3f/VxjAQbOJRMXy0jurckaZmu08
X2eZ/LKSBv3l1Hu1L2TIs6En1tOIRJohbvoybDrZi89VyAt4AMBuyF2R+Jbg8U4P
ZUGnw0UYlcARSBoEwncBXsWVmKl3SURltu2LzaZpceH8uLXqEoZUKL2rkB8p5rCR
9nU7qExbqPioN2hafVZwe4rI2Eh4A/NmB1Ef6xiB23paLu/k9YlDQgxWUzA4Wwpn
Uz/IT90ZSCLUiCMSg/BbhzRJaME2OsQSPu2d9ElopYgrMKyrULlA0yywE3gG357u
72MxtqktLZyzfOsPDCjS2hTf986gdnKgP4x/TVoaNkRnJ2IAbbfpk/tpoU8g/I3P
wcmBkINy/Qwjx1I1+LJGocmXv1HcKgoSaLxvzdot6ac9O5B9XkqO+H6KUSddPby+
ejadrLhCE8WbgLXZobDbupfKXWEjE16bRfv7z4kIQY2WxRmDHL8AFIdQaBmm0dXX
vX/IERLwBGDfZ6/h1K1xd6d44CFz24PCEz9/7Z+8Ra4k0tCmQ8+MhmbWZ9i2Hotb
Aey3UEmTWX3iZsFk9+/2b8my0nq8VK9C6hCML81V/EFPGql3LcjCTKNeJyWWbTpm
aKJV9EGi6FPgC3UYGea2wC3puN7YwLoH+lYkNlLSrNHYfPstwOaz4qLBclGb78Sg
IsErtsWSrpqlcjNGef+cOwtkHWnnJqc4CoMWiZ9KsQgukdT+Z8awgYmIAnTEWTV2
uNAY8SxdLyKfXXq73gl5yBsIa7b3gi0vafCPGeA07bdH2LFJABdmEBuOjlRcIwlE
gnGgxugE3FJ8kwlntcX5jRZvBsaedQhh2EzAHDok5AuDhScXmWMcqh+U2cy1522w
3raDqTIQ+1g392ni7t1eXn9qhAbCNAxUJnoIwTGwyp2TLJPYpQbMKrBV5r6ImK52
bF+20wJSWtFatslgkjtxfabq1dhTAjeN/YQm9+6xwvo+qOgv9LZVM0HlSQhvK5iu
eKUbuue47ME9mHxkYEFlDgfOgSTVe010rElVSOBMgbtgxTBvLy11Aziv6X+E1qSY
918mOk/5nm9DKST9YPigXlGJIet5Cye3XRo+Zx0/JhIF/SN6DWTEpPa4pD5bWtoI
MHvYVoJpD80WOvxU8kpjQM6dT1d6Mw6iG8ZPbmfo+dlvkblr5Qu5rEK3GqbOVpkQ
pfJoVXkSZoMJ+38EkEwj5X/GvOVkGggyje3wJQD8zfo1Efm4nl6xs9d6jwfT/r5D
zfdLtoj/UEcmYqxhuaIbuAc4QpqisdWXwgM4Z21nmFKsbpDY63l5IDQESaQGbTvy
xtmccVcATL8bsOlRZww+6EHyxPreiKqkXqYz+MhEYbJq3TQmImZpptJ7bqTPdB9q
FL+sFpC1mM2vsctIiSf1swWDqm8iHcrxeajuWfPLVURdNjUnYkbz5n0UYSphpn0q
Tt2ASkIaehsQ+zRphP9BqlgnUdEqS/FCXPhoFgdoANdaUaBso5l/9lXmZBk//XeV
IP2loTq50v0ao1XBcVbYwTV70XNGoD6iecq+yngoEPkEvTet2ojDFsnd9U19d4Oy
rJ/WPBDQpuTx5H6JW/IkJC1SCCScXM13KF8QJDzL5elfCMCv1qX+iZv8K6x4hGrJ
vRNRg5uMAsryvFhJp5HUx6f6zj57DaMEsQNrOrnQvFBW1xVDRtloiMEQrcwU1raN
FcVXJk0mqa5R2Rbvn5AaD4RHsRBgqRYvAGBDk9w4inI1PCteGNd0KolWJoLLUHmF
EkbT/P9lzL9lW7aFYa7tHhlUxswd5G8L0xMucu2d4Btfch2ot1KH/wFjZou7Rj4V
Ja1QpbYWhOFZUQkKgIO+2qO9dqnwwxqmz1x+Nr3lU1+4M5gua3lD6zj6WpY+2c0r
2l4T9GUTphEOlBhn2AWr4q0/uaDPCujYOwqUp4cw0SiWKyr7Zyl6pDRJvzM+awOf
uA5ukE8P8Qvr5QBindOXkfA1sepUa26EFbIY0ZvTaQUxJKtQ+hnsPyGWENQlnnIq
GZt+RhKPGzAM7NvmqHkX8UjTZ4uR8Y5JNnjkcVA5cqxsKLLNThF/TBzBMpmsGXVM
iTHPAP7RKxBbs+94W6k5o3PBScHjt3ocVH5TQ1fqrs6035sI8UhNzSBMkp3g7mmt
CArtMh1/5urx5iXLYYk01v6fopkABZN8V5Z0TVFWwkwk7Yed+ghWGJPRZX4Irmdk
N2oiJ88bnKOewTG9lvqMez6vEE3zQyhw+YQRgDwDeUWLQzrpMiR7TlkV8c73kcSy
++D04goEUXvlIQyQonYRFDZbaI5Mgx7igbSO9qzDrBkZ7Kaqm0APVlRr4SlwPRW1
cArz7YtGA+zffEbaSY6kJRCWmBVkMgGK08wtHCaO6OosoHBnP0m/zvvg41l0BY4f
lDC1+a8R1JF+oWZD9cNRo04FjgX1TOossbTf3fXVeOTCl4SY+9xUOcQDWrZ55wgq
WW9xu+/ALuzndvMDylH4WWK1f66LUUzTSPN2WDmz95zDEfuB9H6NA2Q0Px61KH7o
+ioyJvjDAmsp1yiBLUoqLLCDh4bhNVMWBbh7DdJUPldOT032bNNEBy18MK4YUxcN
q/wVanZLQlCgkrd+W5asorqu11IykBb0FqGp8CDlWX5QeJWxfuq4QPB8RcmXgHT+
rgWkS73bR5DStE2BB/ahRrztZxnTKTBKgFtUpQUymWbPrJzNyGJAwTS6VP83I+CB
LusmNhDGzUfwSkpnujb0SeduIElbTvC46pbfAat1Oq8g/rWWnTL1eyKoBRqNNXKs
T9fmVKQGvvv02mE6D/MYBeX0PSuAQtK9pOAVhCFam/Bg6OpBW0fmeDtZJg9YQzNb
UUdUGb2f8EeULakFkZ8+9WAtZCHblDVZrXw/cC+YaLh1nrsfEcnRbq+jYzXEPIvx
/kVbWHYvCCsWWwC4/yDk4LzSDYwSJ14ly8MIg7GlsWLiEMmRso3ld/L6CQ+G0Fdh
rGcV2NxI+4wc+hzgfopnrDQcid5zY2roLBd/RvXCDappGQdmXsip/NrkKykmx1bj
0Tryn3eCt4rwMptAPvbzMfpPA70SUU0dQeMiLKHzH6MU8Q8VYrQFn7hMiCV4XZL1
QZO8ynRINSyxWh5KIECjE6COwE4gK1QhIdzTA4NF6rBcSt7QRg1fV0TzI6vvEloZ
OrpBeXPeGHJt29QQagD32rIqp8jRA2/h+3ltwxXzx9Ha69xp3cz/IDtL4n84xKZb
7karrI+bwQeLT+RNlpXAqVFnITorvM9M1Rkxo1RY0TRYhmTrlxfpzD1NotTS6YEI
PC0AbkTGgoN091ngkgYqkv74diO7+iL1+UvtbnmNA0r9fAV+Nw1HrqZsto3uDJh6
t7Dd8uh/kel7wodgRncpk9wThe4saZr0Vd9MWe50qI5zsphaA96ZG2oM6x2QczIx
/S6QjfdKQ65iZsrrKD1Xs8eHQwyg+w5efT5XDB/T6ND0FEX9Ja5e8S5mppIOock0
JTPz1mQJBG33s/yoZsabRW0iMmbdxjvF6+LG9toubvck/shp06edpGOm34u41K2p
R+qYZYbYT1kJKj1Gs0gw7MQhJY7rcrEpVyj/LEhmLXHcjxFQoWI6IxENiKfzcDbW
iivEidWtwW0MFNRbwEN500qS1tQWgpLDBl0IX4PMfjGjcMz2r87imZruwZEIOYTp
OmbktVYZ/hgAxnNjtCT8dgAxJhybVMkR3h0un+nmaDt2KQmGV7wzNBhaLP9GVJP1
YHEqKCv1+cptNvnyy0wDRCu9EEAql1cFw0BH+rMswVvI/q5TGa/yRnp9Rq9ILYVi
An8U95Aqkf3IxTiV2D2ngmI/WgeZ9OSwdRLpUq76HaCQ6h5jdEqpddlgaKBB385k
zToVFwIiqsIPZmLux+xUx4ccqvlsrNNZo/O14cDGC1mg/fxM5a2mzi8IWn7P09EC
UaWZRGqy02QfBLVBhNp9egcsjxeTFpE2Y7orK/0s/HuUZ/nBaFONyvlFFa35+cs/
5ji5EymNPrje2X9rjGUC8Z6CbMV76uazAwZ63ApADTB7QkYW1NIvpOh9N0x+YHbX
m1WdGNemgNu5NgBjV86XvQO1dQLAm8eBPr8YXa+KBfzg0CaYwZtX35TP7dQLb1wn
K9ooCftRVz+LReWxu8OhQ0N5pjVQMWsDMsClIuEZcgNAybLAMslc6a2WkCfgpXOD
HhcGsjX1fO8Nz1L//HAN/wzRNOWnjZYoyqT+R+HYLS9rZiJ8rSUGndBVDFP96BOU
SDzfZGJTitOZFilvzjv6MntTXAv8a84x7J5HWSuEJQmagriT/+VC/hPJEK2QHiX9
eGGDdcAwY+GQ5S0hjvJxPcYvfvk3If0ljxJUMIxz2XNIEZassEycJtcfON2m9cRz
3ERZzSdO7cZNimFmT/urkQLFZ2FTuXEibT8qztqdzaxSgvmOiZVSlvX+n/wT+PxY
BYpAeQwMQq9XfFwKNMMjbGZ6wJRWXCc8twgkSFA87U0z32EllAgXZ+Yl9FUWdTdl
61UP+4v9RwfO340MRfmgNKU3AV5ofJ8Wug1vcPMwsvNeIdW/6VNDTa8eahQ6cMnI
PSGORP3nNhSwYHqmwXS4OyxEkTclxnViYncIlEfM6Wc3V2GJi0UE47jpAGfDqDPA
0+/amTzunK+eEdcNwJv6+4bjQXZ4Loo59TP6xXeXd8qaN9YtL8B2DnMQDh1WrlG7
m29kyL+7K1FQAtMInuTzT6e9kW6u8IIAiP0yRZ1j7AuRL6XbdnTsy663Ttv5XT69
il4nar9YHl3Oz5yfzpxZmAOZcqL34LYBkkWzhTzS05so01Mghh8JeEUb0jQ5XAyP
UKkn70xhMZ5+NmQwq2xGrpMyFYkoaBcCfZMsBMY0bCGch40zY/5bjlRAUH7oLc3x
3POo+vLP8xjE7VTDG5R5DS1kQKPx13KOgzrmHJkLfsEQe1zz9+7i+rQ7FO5XGAPV
w4pYPMnThqZFWAzLvCqOzEnGag042IAMIZjv83ePKDaKxkB0P/4+n+Rf/y84PLuZ
thBhMn5aM0G9H36v1cnzg0tVCDiDCX6wv499YJzdRUg53RF7cJg72zFUu52S2z3P
XhPvCufizShuPuHXUBXMN4U3430OBJJygKOe95mudxjT6zwB5mrEDybPKVfydmxH
3CL8Qu9m66+CiPddRv4qkQ7/w3GTjnRCsRLQfE6jKZLnJ5gVsKJpMs8YHOugHSfx
1DxEyBlmh1MI7BAVVthCDy7R3oRLKOkUtkuTdAH+ih6KNeussEC8tY+Bq3aeSQGq
Cspj3H6QcDvKxMSTtkUYVISEGUK0hWNG9FFJUMubIDqzI3ED8D2S5AMIwHOShGdk
wPm6EMqmFv2dEHZ4gjnO5oUXPvLM8TkimXeQM4xJ1czRnjxs7Qyp+HPf65TIxxL5
lOMnPFjTR7EEkHC94g7a0T2Rc2+AyZegnKIUyP1nJNReuqMi11KytaRL3EDDofzK
OGhGmAuA7wTDLL904X9VhbYuQyEmm2gLfDsesPT1lMN2GS3HBoGJSd6LbtlmFtEe
Rf992emygvd3YARM/+SMbyYlMuYFj0MvXnHFuGsspf3nIYw+jMv7SoOgGdRzdEsQ
0m2Yi61e2x7RxuAiMLxICgjR3jQw8zBJrsEM1qBj56NxAmJ0q15V2R5qRiCsANQd
79llTyH1JX3FyazohRXx8zAhPqgVRydBugffJ78z+l8BLWLujaxDpTRWh03C2vJm
+EVnifnqHjyQSBKqDRXE6XtyK25e42j1lkbKltxUnUvncMoH2f97CKPnrcNsJIiy
TzjSd08x5OLPAgMZmjaCnR/vSA/Z5nKqEJFrCB7t1Ko9zkxt5+l0yqY6RMAl1P6F
F/m475Ql9kmpKJYa4hlbOfj3JD/zutSXx3fd7gSJ92S3r0qwybYquCzma/RzGw8V
p80HRPkiR8NS55zDvBhzOKQ70KroUDmKh2S/ch4m9GTZihIiOIsGq6x64OberH49
1hNiuxuZYNhm/S9s51chIn1ux1qJROiCSDE3ZYCbV2XmKyulTWRb8YD6gY5XnEtT
lDZJjlIGicEUGxzSNEhEN0FeSVIFQacaJ9WZolQvz/+xfgYmx5+Z/ApeCXNs2a0B
wyXFZQtpOb9BoTGDb/tdSmDV3FzxY2Wk4DLhwF+6/kUXjPMLZVq9niq9vTHEG+cq
5cflNftPasCNpfBtr0tRa/Tw2wDc/qDZiMrGd1y9QSs3+o2aOP2pLFaApBsg9+sw
ACdy+ys88fMvbkJtFcantD7HoX/k+h+qg4FqRIngwIkodvbuzRIDL7V21DPx8/qo
Lu/LfpPs/hG45BiVB3+RQYf0QrfLAU5F1N5QtzwM4/K3W/StXtT4BDKY5fb7LEl8
c5yzb14tijWmc/68FAlvONlaygytS82WQSGmRkIKjZVNJlpnxYJvSQb3/2Lat7SD
S8x8DQvLVFGOXD72TXU4SZmNah8bVsY9QeUtDWaTDwdnK+FQ6jvJOjcquKVtupFa
QY56buIg+We5e6U7wPZydE2OmM/qdyU8vbiLtSdJf0dvfYFdJ2YU8yiY3uAt75aw
0R2GAyzX5B+QzI2lP4/z9Er7u0ZDhxnv0WYfIsyVgk6c9K9w29+la3GYEWRoaczW
vRFm8Lrd85kQ5f0CG/Gvo4CVomHMy65I42yGdY7ZSwSF2YyD6KTmD94UJl8j3U6O
o/BqMpvgUJdBPRUKd46TeExVPIujQzGc91mRj0F0AsziLngvuU6sPmqotkGjWm1S
eQz0S69pBMaI42q/Fm8UASarUPH6sXbpyx8V1MOH+GrRJBjeFgsGxYDGkb338buV
F/1XVg7oVj+kZKGQthuZALSNwBNvpLU5ppc6v3quoxfPTEYqznH6DvF1iAJxjqrW
rOwI6hmT8DhIQcPFd4yNgBRZStyo0hcY/TuECFhZdW2beNigNQZsfXNLF22MZYMc
n0z0focjFfrQPgDW/6azRHQvtKPi05dHj/KwcpGPKzy67Wk3tOD3KsjwldEVP27s
fsd2BHYpOaJX+UjxcVNQg5+sIisN69vjBtnhJlHup8lgngVyYtJDTLl9mKUe4tsv
kKehGzdDkHm7hdPfeM8Au9NpGTW5tt3Wt7K+i/ERIGy8p6Ul56rTEsaQvywm72gt
onLYTjVtj4lyZ+h1KRgHF2IPDWih4iPu2S0N+Eb89qwv2nCpWtBZQbePyoZkfysg
y+Ne5H//8ZONcxtybu/sjb3kM6x4b+Rw6s4uVPah82lxDDFd9WboTfn2xBUXa4/B
lc9vsp1ET4eBN2MU2Kgl3PIQOxrWALtelYJbfcjWmIGHWCMdHNqeTgVW9vs08iFf
J08Gh0qjmZczhQYn92VJPiuOzMNaVHEIdRv5FbPWr/P0KkFRKJA25GH91nzTdEsL
lEBwWnEeJYwlUS60o9SwGWUmv2tKDeXkRsDojuno3PPRGSBZZPT6Nmg2tCOj1pPP
w9u668Tspnsr+4JYisJFAXKs35iat+l0kaRGd5i2K3hTEUJULVjneGkLYFm8dt3f
19lk9rm1ozUG30HVSGUBC5NFS6ogW6iwMKWfJ+Sv8R9WKXxB95Gm2A2t2eL5isjm
N826HKyLS/PhRl9i+7uIGr5SoMTrEy42D1qJ/MuC3JVEwTzQDgq4yCYlLoTDE5dl
dRBzHCA6SMPzc4stDdn+kG0uiDVkf0VLxJz5K5Jw6wbWi9PTPjt7jz0iSPTNqLwz
SKGcDzFwu260t42G/J/Gfz16HXsfe/ZZE1ha0WGvYVizMflDPusZcz7UOIVMZOaG
+F+Skj0Ec4NHxrkOGdpSZpRAlar1sdz/4Wz5vCSFin0AAM/O9jVuDcsKGe5KIMA8
k4DnyFyYSkhVRitjMdT6UomF9m7Pn53UGQx+h/jersaGLerBLqSZb4sXE5lYU62J
MIAfyy3uJSYSCYnr7eA4kNi1h0F4p38xTrI25uPpdwXiK3GaVpLy6g8Ik9ckzb07
vVU/soth6FjEItD0IQMS44Au2LXcqtRJPOUxheTSHaerRbInunUygMuDvpVDGWbo
+0SBSo81IE6eAhohwtXCXbWc0ai0rm2AP/JDGLcTEy41t+5vezSw1+WlV/rvJEtd
boJU3x79axa2SUMynby1pd1DegwOqLJitf1Iv3TwQ9f+tMJFC0uf0Tcd+N1fg5De
TXx/Rpg6ysFFUzuIvO7BfmZeRG8xBk9oXnYk/daoOLObT0vdHIiTaN/Yo9Jv2S7A
bveOEA2EVUIdJzOTfBc2cxt129sh+/7/tIbr3h5hKhGB5sluoFOq0hHxOH5CXl3j
YQvi0lPQ/bN1C88Lb64ciPeP/PuyPZpFEUcfTpXll0U0TZTtuH5X95lclXThNCgR
ugIBt4CkM6UH5f+TKkRf94qmjiJH67v+ExdpoMmcrX4pvndelIr+u1pfpv64i1y3
apjIVeHVkLgFDlzAetpoLY2uTMfPNfSo4a3hKR+VrNen9zHsri+rTfakWDpM/LqI
3om432MAFubVYyDN1D3AlHbjosQd2ywQsXfVs02wCiaYAXNg3Tocl9Vs8s6CEVlm
+9NyoVdUB1dsNUp3Ty5glOOzojyKAw54uaq00oafppS5aekwdbZpL0HhvokOcJ8z
1N4ydoVu+nxBup0yPDDnavxAAbaST8a4PeuPLK1Hl8wcnSOnZB7Y47PPBj7m4O2y
Ke45j+Fgp5zC01HEqrrlY+IwLZTPac4h5CeX9tgQoP9LhIhXxB8YXm2e3KpQ/ehq
wMnj56XOKpzA3Lisrr3kOpRSOz2CWzKAMJWKpN8nRdCW1mczyTKueEvTzHFBYyL3
t4c/vtJb2wxJ7uy4cnLyy1Jm6nAMbz6lfj9sZrDiaVYP6a9ACBjVCCQD9Cjiz5tS
8a7AlS0m3xDyFEpqX38XRroll3RN/KluQLn6+RLbXMcWo0G6m6aT0Pvfq31ld8jB
7SanbxNwwjpKpDVgh2i1lG3G6hZ6M2ZgrCwA5/5O2IVk3e86YApjR1Li40pF2u6N
a+27zQhH6/jBmdGGRKWNhJOfImd8GSoPI15rkXqkmmlWzEFhQMm0Qk2uzYkC6HtG
Wxd+9y3uolJZCyZuf+L/IXSAlUk1guwTz+QSgi5VqIC5lYQFXd6Yq0S6u/wKRtzw
tto36qJgEpaj/QqTRzckyhIgaXUPMDmbQoIUXI4510aL2EnaCg/qwHLPypZFeETb
QGz42cPlsOySRMX6UIhkiYprKuGVSrdNQGotXzXt8y4q2pQY60ut4NF+lnrU6Z41
eWIfJ3tUi0Yo3ibjNwwriJeZuCV1maecik9TSolBpwtP9iZK63Q1Bs8IIQvVasYa
Sm+DmtGzBFF9VMFrEew2tQhKrSWYDaBQ5IUKcbcOQCMGlcAYi1BDxVLliIapAoi8
+Q7yWUqkZuuFp5IKUwDSxtFccgPKNRSvxLYObqnH61gaMmqIJoV0w3gwL5Yy3lHC
4TWb3CUAwfCLGEXPLpVwyvgD/4hUi3Zmx9DcbvI/DPmv7CtyGUX5QQpl9OxalDLN
qYVybJh3+PIqMgmM3e2+0ZZZqsf9F9wYuXFmdPrTtsbx5zn/XPvqCm8hFTWhfS0T
AQygfEyRWP6ulrFGhWSwD6H7E/guOVPmDpfGi51XJ6XKlHfq3Br1fp/FAuN32w9Z
Msi3++NNgyYV1Rzd5dUtfmCqPuKpRcHW6E/Wwmh+La8VDN2Ru2FiXrMd+CXtjiPj
fC21oUyhRVrZx4x4NeeMHi3LtKBRuwLAgor/xT5AtrENb/VNtetD/B9859a9VaWD
2RmYl8Okt+dHFpRjK2JEGX9f9y45IB9WrhUsQ72Ks447rEzJG0W6U0fNkl3MC6pE
gi3ZifNi/pmR2yTF69jbdX+fRgx/P47LzjOxaAu0ai3/O2cBemBEnbWplbzLL75P
eL87mJ7MWQjIWpCXukh8qK/E+0L3bJ8s2KCuoA1Z9O9X+sJOTp218edyFTEKgJiE
SjbgLAdxAj8BkzCsqvHYuekNjJx8jQs2R/tYCiaHoKnmDgaHh8GrxQRFWkDLbpPR
B9kBeWRlt3No8Tk5cgsq8qaM2x6LJdpxPnbK9T+4kHvNi5yvMUHBfU6wqRPqEE+E
zhn2K+61KHBR86QYGwy0EUv9QD+aCWch3LNM2YtTfqZND9e4K2qohwNwFrwfPs+i
HAShwKYc1andmyCegqYHgbkzsPBs5bimFXzzGFjKGADZUNEnfLTxTcvK8gar+AOi
z0X8cc4a9f13Rsl2+hJoacoCE+n+iT5BnE52yhVSVvRZwxwTmfmry48lnbdUeWow
dDohRzkGLc+i2ER1T8Hfw8R9wkPfYiqRcYqG28PdRck00RXsYRN3vHTl81brGACF
4XTX57u8Pb55cDxvF8R7ObKc/ShtGDBAFwANCNww+vNKqCXIdfCvrarRhnnMkGVq
MyIdk7xFi8Eiwl1JtPLDDJr2NiH9keDki+h94qWyOe+d/us7yC+4+m1YEs+4cpMI
GVyVBifg11ERw/XQvHOweZulfwk0+StxFFSursPplxcsrcIa+3EODZ8MpkgGgnux
i4qVa1EKUV1md1x1Oh3BqhAr5uso6T2MzqZbbzrSJ9JcJM4CyRflgP3h6xJbt1xD
RJFyxv31+DYt6qGOVcJV7YAWKNsQ81GcPZSUZ+JIU8m29QDjwRg0ZDH1OZRBxToo
vBxvGs6WorIcOPJGM86lia8ZvM15SHAYgbCs+ekdzWBs3ERxB5+Of7UfOGp42yCp
+hnCXGfLKWmb5oDNB6KMbQJ7Hfan2MVhVGxwVXg8siwEmoSUre8a3bZglx/GEHy7
lwTlDYfYiMzt5gLW/wT/MH3N8erloBbFSuMOoSrrcfxSYQ+0bjWp0FgmdWDAzxeh
o0aBYIpVTpBRIKgcUKiJ7SuwwUKgwqJ4M9x1o0ypl+tCu0lgEVfFL7q8lx0yerN1
5lNMN20lEONI5kymbZZGH5uo9nbK4BZ29HDAxFTwmZBPv7bOtfiWE72JcwzZFqel
VmjMLTv+JNzLMJ+y7wedHdyJ71vqFOkKim5FnZuUILtrOfRKYY+okwbpalQXF5oc
3JF3F/OGoeCz6xoK1YYF0jLXRaffyxU7zMRrCVjd8k33gLZen9UyiYcKckmqKNSC
LCyxsSZlHtozz+2piakhmPYpvZneVFyqTCz59paogGgHQeOX6o/pyb6rQ0DjiaUJ
s5H5pjtNycgt1iMrC0HHS8BccHEICybRX0AeAX5vQZZ8imcopej/jJZweZK7MFPm
lxmRT3htSJnMucNymFYVfj+LeP65JTkbKMb1v0VHe2vXgwfzQOOby0qV0pUhk2av
nA6Ow7cz9rNd1L0OaLZwMlbMFser9/ZTq3Kjxr+rVVtWAhz/wyIJH1yHElR2PjO0
7cd1Hb+Rjjjgu2DSsJR1Wmhaka5U63WdBfXGJptPOb2g5Ywcccbc4K2vynDr2Gzw
vrq3OoN6hZs3h5ATWMg4WDrBJ3e15zNy2xNUM3NA1V0ut2nG5BpVOKsemsaSALqv
hyl8WPCfAS5PMIR8/gpQioDgJxUEiU/7bDa9l7678OMIj+pmYOgiV9/UBvcq77K1
f6ngd+RNJzJyDEfHQfoERwBHuBoIwx8sPO1bPKTTrHPLq4exOyRrDrKm+AY+Eacy
bk/39yvPBis927/Uk+BOM4cU5eayqJSRHxSxKD00n2jktjRvptAYy1xM2ZAt+Dff
2KBL+nUijrKrj/3K1jEgkw84FTC+K3lavM0wDp+NE/niYkrEdjDUGZEX3RHoYy+D
ulggBJFrAasaIBQNCX6Puo2wi/RwLtjKcHlNalj8WfNhC6p5y4QlMVkI21NRS9fn
SzduB24R6zkKqdtm89tn/owMTMb8uTFhmdGgShZLZl8x6FzH69Gqgja+NsBe7xav
67Qa8IkBhJcH9N8UjO9Lx36DFL86dHTu7OvuaqWdZevS3lzZ4ffpxnB8Yi+nV+EQ
E/iKwKVnCXzZDYcQJ+97rAML8npNg+/2mUsLAdfc14wjO7cnzPoHUI/A5f++jPKz
bWD4ZpXeVdvBu04hyUwuhoo5T4iqvgZNehdELQZYC6Ln2hOwE6Id7ULCKkJ/oVw+
P5lrrVgnO8OuIOFO9HnK4YYL31HHRg/s0kBOg8ud+OCFw8oO1jeVtizouav6m3Ot
P0RV1i1zB0uF4fJRv5wN/gjWM4zrdbwDcInK+Td5nbrhNfJGV2Wa0uC12MiIm19A
m8B+JwQBHIki8u7iffXg4MP6FvlthzNZL87m38QfB+VsPSmxlpPwCAWop/r+v+/W
K/GworVpyESA+lhVrBrwUvSpd2b/iE/A80zGQDc3GLeyKN+zov+MGzA40sN1iGK2
LIc1kDfgdlBWPkURkWr9GBdggGXx5bTnLTzbQSnaVPzHmWsFQfZX8JLaHyaN2MCE
inpuHF53FOrgwy0yjhoTR6Pw03ESCkArPKN3wTkh//uQSZAhxcYOpoOKybGzxyz+
vLqUkwNNcQMCDRzhVIqUv2wWyqT+U9kfWbaPC4/J2f2lTJu9vnzPZP5uPA7wxz3k
J/FQDwDeZA+qZ4Z1mz5IqiLA4+HfWwqY4NdDSOXE19nJdTTO2Vt3mOYNW1lrzclO
yavw6VRRnR8g6ccOhgYnFYIDrygPyLRyEApVqNiGTPGen4hwbdyAzwzvChdUVBMF
zzGr9M7ZCawGsniyNsn+tEwYzD0/0xreyMdEkQ8UbXUFgbb50oI+GutuQW0gnvuU
slIfAwDsEGEEVSk0TeF9LSVn8k/IvXN4WJ+AbqMXc3lwDKivyxW/zllreH/VYD2S
zSHK+IAbprR13IOOFTcIPRin0V16/gMErMJgO4JSiRANmiCxSrJXf1lbP92Jd/+a
PBe+DtBmjgVNfYpzl0dT372L1AFsGm3Mw39eaFJoqSwdWPFSzmeT1aj7z0peGkT/
cqh3EOKx/aHy6tImweqKLs2Vgvc3vG2Y/hoXQcSxKmzoKN0L1QNN/+tHK5oucCZP
2pOENLRJp6Q8rDg0CuLpxF+Dc3gXgY5enSfEE670e6VeLPLIEmPNqtV3WM8i/tnn
yXx07EJTnNQub2BXcAA4LRLwc+Q8cyjQG9QL/Y0keZNLvs6I+Kv5FsjYaUthdvYe
MMZBjJsG5cygpVU+Ezdr7BgZWaLpDRnQSFrJ6PeGVMcCHEQ46kf8uDkkboIDHsKN
vRI1rjdmiWxJKxIODnZmuFmtdl1G8BURY+mSkJrjb1rVg8xaAZAcN85USbyXKE5c
uGVw+BYTXFuVNQwxB8fomo54T64M0G7zPajtzeqH/ooskjkvvccu7IEivEmCqp1O
5MD6LLEcbuh7oxg4sWlXSim3lOSUnBqebjb+TI6HY42I82uYoE4Ngm9sNmrYLt81
ukVT4g6FWwu8ZZTnE2yr+Y7UWEFfwoYMx3EfbbYEXZ4usihTgJNfVDDP9g3nyHD8
Lq9UZNIpbZzvV78cDRT9c5IAgzP2LTk4LQOof4Yv9RS09U+4OBkMoVYcqGuYOkf0
PfB498xY/9gJvFXyb2ss33xdf+JLCNiijzVvbpceoNyqAkRazMQTyDxUt16pU8F4
pIoUmsZK+czoTzC33MU66aSK3lH3B665/6lyjrfbPe+N+0bot4zrxqQEFyjGRGxl
u5cICUk3N0Iure0ml1AwERXktRWMa6b4QAVpMwhGm/AW7UU9ZxRfB/rLnSS2wtBW
HUCAI9ClANRumPzyT9brmCNXPDIjXIMfhmp+u1ZJzEKx/lzNZXpRsuPnmta1FFV2
1z3ROSQqEtGwxyzi5gLKeZvb4UKU9kr060UiTzSqKY7seFnYokaMHkvl/+IIC9Oo
NUn1z9Rt9aXGaGgv+P0muVvfS/sB6rhXCVcDVNTAuSMqtAxaiehketNWJ148txhn
wWzzRAPdkN5K2U+1RXrIB5pfPMfz5016H/+/Tp9wWSZTt1gQjEQfIjs3rb0kuCfl
rlnwml+2vCMWZEhkXeHe9zVZyhTElfdoHM3ysoLKh+VQBem0YSW0NqbFXyvlBQMg
XkVpXAxPAv3XDx+0utKrNm0NXSvqnpFyZXmEYtU6FZuI2vL33SoJWP3axVUX5r7y
wHs8zFEkQCIzewZuoJWDc3TIw+eFiJyppPKWKNdUwz7s3nQVAJZHySClLfYQoSC9
OKHHIyd+T3jwo+r4e9oVYDO2wwBVNGKNf3H2mvsiwSO2B/VjnSy/z4KnKg5wcnjE
GyT0vJqzETq1YWZLBK3w0EFwxexKUTFtQZ3r5Ksz0tgE29MTeR/LPOmpe2GRlVhI
zSoOaHxwfnPFaKHWGldorjDL9hF1QNGJTB4BnRsBerqWsXPfpIU4koTFSshfMefJ
PSLhOWTr9dcGR+5yci3AdXioEmx9lFuBYKnEktTLN8qwWHuY8LP70Z/KSrUtw4sf
FOjHUnHBtaHlUVXd7oUI8zrkC/Ld2QLAFgIoh6y43TT0OxZzECtKyauc9JYzcDDH
52nuoo6uAGajJAiq/v6qqOmes7AJ1WGUw3sxxCcXWAWsF6UqZbxw0bdT9Q+tWx4d
JmCSlzCvlWrUq/GRNmFQMfZ9ke7CpxG/KbfDjYvAC9Mn8Fkzrhd1rIhZo/n0v5s9
YHERXNApTWkxiQojJoBIFl7bVTEIBQwM9HBt4YVZGY4mUARcygeW0Aa0yHHmhAR2
Aq4Dgrb/VEtU4nh//FLrF6QGlrO5bmWoxdGEnYDrUJFbP9xEDVC9jaMgPb8ISXR+
ntbNE7e0j4HH2VpJG5BEu4NUEEFbiJck4E18ssdhbB74xabDJNQrd7ciWhhIi5W4
AChl7Ihl/Y2VYmFEX3/JfI62/7wInC3FmE118T0MNWmK148nYaq0M4aprjEQegFU
+QjbsX17ZHNkaaTPEYDbhvVBHrdsAcFdBUHQa68Ce1GgDholrwqH1mYOUImodjSq
6ymGDu/TOeGZ3ic3GBAf88oGcQ8n1TjzAdGSszVfG75VEUYzu0xSiTCHJeuXoZ/q
FdxFSfucNVbEbzzc/SSdZCRwXghGLjCmEQ7sv82RNuebLW1xsLm/dEIKk/WRDfWU
HPbTWBHMamPcVbEhtLDW93XEQVF0r3dsme3O1Qm3/V1I4PRvzcHC2hh9aY729XUY
SM+1BmlXksqtPHAvjsc6SL/wk5tPwklCDKhy3zgqz+y41A9SKMVR6692kpsl1gLP
R77hmX/z/oWjELfYHQ5wa6+ArebnZUOEW6HuvUhp5FKkb2z8BspTmsIsrJ8u31vV
/YEX0hQ1Hwn/d1XRsXPKh/NgCk+4h0k+Y5T30D77+2Od7ANW2TQHAVUF16kbYcwJ
CuL/BnjX3CFAx0x2JESU3G9rFG3U5r/H9ZKF/a8k3yDH744HMXOlaozQ7cRP9o+V
F5uQDdyC5Ie44pfIc8cVhY/sER+PEVdKnxfiFWKJHpCzz4+r6s6mUtQ5jXLfuprf
TTbP2t2qvDlkn+fxJ4WPfhUpcHYCosA4zn05CUITFOSUQeqlOErFvUcO1E5D1KOi
qQ9oyAW8r6S4MPi1gvBScvPRNwMrxYyS/Y/lXxVBKhE99yPzZaRnN12Aoewz08PB
2SltIZf83HaKpgBnoSjVjmg5OZglKHjmbeW1FFYq+9Hyko1ncT1Leqt1HM8TNphC
v65GvcCPmz8bMjvhSJ5qR3mcQwpD/YxVEuuRv1CLhhiQL/ml2QPqFy34wC5UrKFu
xUjYG6X99rk6jg8jiDCc8jwwl2ZqFoVIvjnY/hM9zItNWvGrBeAde3r2qUDTFTFa
b04zmlBwoRInfIV8yuAI7NHBsUtUJIzaJrXYjy6mkoUpyF2VE8e4QFgtNc7RIWRm
BcwUp1oD4vbuJHTg8vgB8L5sb/nm9VPFZSiqxRFG0CQS1pOtohXMydkvA0lzNzYP
v/XtYs2I8ps2u0nChC5xSx23iwLmDlfo3l1PeXKUwEvAz+rqrX0GGNCcSMiNYozz
zFBO4TUO46rNfRD0DijIcoBQcifW8l3yBNA7bDVNbEnzkEu2IZjlOU8G98IWFpKB
wTvKGj8SsgVnrtmZXhU5JutHZYRKwWp+F4/QlODemIswy4jRMn87XEFsMStkkPa5
oDDTW21npJnkHDz+504t1zjc1SNYTVESbjU1URpvz9KyX1HzSqyK7A2zzvVRX+rs
QAGYKjUGOGp1llNXNPv4myOfpz5nfC/8epb0Zsf7BlPY1rSgnizIQZk5h2EMml4z
0nuLVQyWIJy5autVQB5vDY0TsVGQAkVBPtO72k/UVJybDszQrumC5ih9dBasf6E0
uDCMw6TFwZSOzyjO5h3HNCI1ZYE7RxOu1PrFsHEjc6rx300viGReTnbClWUZxq2/
zJZzParP69T4SJ6ACnXL35FMv8SDQH9rszRDxF9kHkC8McWxV2yQ5Mx9+WDcdT9j
EFiasYyP7oiNATWhVCmrcMhJHcg6+pkinbNZVHjsjnpyCL5wj9dAzqnPiHQMQ5ib
WyHO2uQBt5u3BIAwihxAvY4w7KxpMhXvZolFmAS19KgAqyyTUB5tr7jxsXwYGloh
8urq0qiLxgT37efJ/YPbfT886rM0In0hrbcApeeCIB+ffCV/Dd848Gqno5dIN1mE
5GBJocg6oDkPmuwD9o8Q/D+aoznHg3+H6BAZGsidCR4arPOF2uCRZmvsfStihYaI
2irGLrfyFC+T9PlaL/Il4VL3TIqfns6fY8lB41aU2i3HrQcfN0jlNMnoe6ehWIm+
NDY6LX1RiV2CqhQdxUMJO+DTQoYANh5xfyzjrueDmcnQ63MAjg7PLqOXxEIRErEl
UWIqsFlO7lid3oJtneCvL5boPKVQhoucalbGBmJbpN5vEzvO2zope+s9lQaaSPGn
SfLfcGywrQgY05/jq6FVqx/2nJSLQbHjG+anXbh6unZSWMEtjLr+Qn+TWh9O5mDB
JhpSE/MJq+XDFguh1uVmaX72jeX8fVFyF5GVBTjUjWSRhDx/0B9dYO3E4EaATUIO
5+yZwehX0YtY0BU3res1jfJyqEesuiGDuwUdS5BO2t5rZEOc5bQGMPtEOqyVmuGb
xHY6BhXBJBLMRORZmMfenibJGYi+vtCdjmFg2iIzd6QlIQdfxKNva1Np+bjapa2n
wVnhoiBYdyJLR58yE/PTZq5j3iuvymFpR9nwUkPsmAPxJJeCCIcm5NPun8ape56/
+26q7l9q8+8xAI6gVGLMa4fH7CJ49nVpPxq5L7o+J11OOAwUKIxxmoQ5cxc0Aq6v
PrCwDRlbYEGHxVBtfAkxW/IQK77Ig73jWtAB2IpeirokvEYvgAla26ftItNHkdXF
Tumb8/73uWjPjpi27ed/TLXTALdg5WmZ0S9jYujDPbD40osx4LLQliM2zLye5ks8
MK6QTT1wWkGbPT9HLpo05H9sUqaREz/FOCT/NscHlOWgod98wnHrtlehzmJaWb4v
gqV/ywo6jhPeQ5Mus+P0qeyFlT7ZUlqo6OCYVBAc7Mzhw6tjanlPyiR7gxZaNreh
OCK2Rgpw0m4+OKDzIVnvRbGing04+PbZaBE0rYwAGwuCVXu2AlqHSGg+E32ilVVp
zoVrdjcCZyEI7HJC81ICrK0NH9YGanoajdFzt8QrG4WV6F0T3+eJ5hP9O4Dolumd
765Y510v5So3RW8EMS50BYvO7KCpQUcsewN5sd93XDjiTkV59yhR5XSeoi5u/1Ze
1GlnVe+qqOURjxEiefW38hlxtbcnDMWE1qkJeH5De0aP76pMr7cDrkR7GTrcO7xt
N7QevpMkQ985Dp7tndN7m+aeH74vOEHhp8/UX8NpdDlPWGjBBG8/qmpvpa5weFHh
oWpLaHOJEMPpFAxeE6yK8g+2m+SVTYYJ+FK4MtW7E4UH+DVUuDrKdLvEDIFMDdb0
4a27f1MLMUTfWZ22j+/P+f8WkaEiJOk0qwjjU/eama7QFWsK5Q/z2o98IE26Qw3G
312tGYsthe+39A48njU5FFrk/Jh7+Si0MNTGrm6SpeOpv6aPVnr5p5sw/GEMtnsa
dK+dvx8ps13P1SAZVPvPHUDtDMUEDszEetPfQeLklqTkwio0ysDUAOQXaw7CFwm8
EVps4oGsqAMqAqaLvp6oHq1XxP4wtpgTZylDUsJbxLXTzq9x1U/D8k/Bkrk1JpWv
XtzAV/N+SQw2WA8OheR8C5DzB19hzopQN0DQdWZG2DF5IE7FMITy2+nb+DEnVMeE
a2IIkCcwDx4KYD9Ic4r0a7x9tzhefr0OFCR4gPASeUxCFOskoMrmetJ0E2LOTR0A
Uo+oj8/h9dG+MEx4vWDqYPk9dGSRozPsDuT7D5I5NlePcHxx7jAhvU1lCJ62CTAX
24uVZ5duHaA+hAyqLdz1z3aOEwUJ6l9m9b3/MjckoDdRRw+8FG/dpoc51msXNxJb
zXCltPNAHmP3avs9L1rh635Vwilbtc9C5qE7MsjNwpZEgGYODrEeZAiEBxTbRLYp
L7cL+7PaDsN1i4z2Sd1ZTF9pOlmWNfdbDSLRZ577RLjX5MPzL/Lx6f+Em2k8exgN
IgcyCx1Ce489pIn07reKVO+C/vs2Oo57h2OZPfauDiUOPA3uoRZWsKgOVyYVyD+t
60J4ESU3oI/XFaP675sE3nie0DpsK0x4ztbVUDb+1VzOnB29HkYTfbtk9B7WDjWb
SlkVW3bfaZCBj9mJByYofxSN6vbDjCZWHbk+6QKEaKvBb3pJmU8Eg64SEh6xcMro
u1FcgnzXhEDec98ZnsTF28VUnBc9w+mUjOJ6+X1VMzzNUa8flQAkjHQEs2POn45D
Y3Y/A5FXB3f7txW7XB1es9tDE6tfNsthTVofUAuhURyNMOtJRmWVwi/6l5sPWEVl
KM8ZCazGSlYbcOu9ki6HYyi4ks+6jCtbBBOTt7Uv2SDrzCSwrRhi28fJJTdPWhag
uvGbr998b36VzTdiC+FR6M4sBwSUil2C1pI0eZKJbqKAoBbz3gSa+4NoJEXnDrI4
V/pXaBlKsIVnnsevv07Vf0bndQo0hDBCIYCWcSoYJgtBYZ6TLTvo0ifWaqgTCZkv
KyUoKctrPrtTCPo8BcbK57IZUss3Ob+p4Gxdth3DwBmcEmcrWZblnuNqZVyyuSjp
DtYvQfYKbT78mMDScpWIrRQqGij9CqGGlH5skooAznDzXDv8B6mbs90F+h6SFx6s
U9eXEpB06B7EVItdn55ttzsUgHAsMuTtSaM65z9cQNzUZbqT5aiEmaDiOXFIIyuX
W5X7aeBB6Qno+is5Z4zZ0ybxCylUU7Ay8JYR3MLoS26IKyPdqyipNAJe4eGkkWvH
LEWYsfh+5iJOd3NGeULzDfMXZkGUyKwFslSU6mpWNyi3Ldki+AUqTCTt9m4b63kW
aw/h7aLq5EzTO4zkJ8TZG/EsRoiic8RlX9bU39TDU4Q6+AIHUdq3ykZgdYMmxKQx
GBm1JLwjOQXxvsO1eGMPT69qV2NJaGmXMtMqUUo3X7tXGeYTk9xGFZU+OZP4CLH0
I2omQiLAc9ejT48lR7k+MgU6Xxo9DLTawDioikt4o9gu4axCusW7Y2pVYu39GzI9
oOpUHvrB1SNfbDuEyZ+u+9KyGQsroZ17X7qS6yVjse/gA5R+xFNtcwHAP3j3aPpt
Ai5MeYcJLS7hsJK+kcGS3iFDhCKfkHUXgQ9KPtIrySDoRMwxIJJ05WTUmgydJ3tc
SHcXBXFxJgvdTp2RKLyytRbzlb83PqDJg2FIQPzJitOuplBZ/AzsSb70E80bLuXG
vSfDMSrXn/lZH1Q3XAckyPR6DiTMdBhrGpdldGTtjFGKq41uwzxQMJnF014d24V9
eiVE4UcR16cbUk3bpiPgyxSfJMoETL4DUxh89QVI/8QyPgjHN9r+uF7Uj96Se2oq
7G83GXoJAd2FZ5DShokLKVipDU/uhkCjBMA2Wc1yV1lEe7uREAOpRGa7hd1DgWTq
C2vtSI+/ez9Qw/hEC9N1R8nLPOwAcx65/KWoEku42elrlyworQDQLHoVkW4V1P+V
5aaoGupfGD4bdB48Fw7wEZz+I7fLXtKi2wvDBGbar3YTnxprjBMQSr0x+enwqtQR
ko9IAX7S7u70edFsuOAtIsogJA/FvPPlu8RLv8WkzH9LEypKBCovzj92PXlOBI29
a3ct6ibFzOCwTlkQqmYTtfB01dzPCxm10Ph2PeZd/OSvXxoV8vIZS54x0Dnmwz5v
VnHi5/m+dkNJVY23ecerXyDv5TM+roR/Xm4c6TdAJaQ7R3H3mP+fviQ22y00YPE5
7orpHWZRck6UneJ2bdRWgs9p4hfue+jo6zBP4oDusjfYhCE5aHXFu9+WOG7fq6BV
Gp06Af6otLMAeTThpk2nqBz9LFUHoFvc4cZVfLpMnJ20PkxiATMx1TJkL3wQo4hQ
BYyN41Iz8ddrcwySu8HDys4AC4afVWib9ytZiZmHgYw58J7s6PbAXwrJSsGGRSfF
TKcq+5qydgG4+mHs0yzxo5aMOqjaww6gkbnHrp97BjS00lwGQaiJvyiFmMee62hj
G+Ap7WlqvTrm4KURHyRfv/2nCr/yAWIxglRoA+coQ+sJMuCUeurXZRjZ7MphRHE3
Do6F6nZZ+V6fjOnHleSrKKqXXEKCybKV42EOEOiEBUQzEAjkS+OgCTsQ4nHLj56s
2sjuSZmqbkHS4kZXpf/S/r+vowpaurxOB4YJg1wJADW1ZOBMhbFK6VCQvaqFZF/a
ynHrjAImD/dJ5BDEgj80Rur6IpAfd8rpaLip4C1bb/7MtQJLtZQSIYQBPT5Akp/m
Q0iDXJDSybXt8+DYF4SO8aO8rfQgXc3h3J1ER8YDvslRRiGa9h2iHX2mzrHrWNbP
1rKkaG5KKbGxQr++Jkhsr/ElBw8Qksmy7biwvLUaBJn2lfo7bRg9o6kDBMVEQmfy
zRp9lbdCJC+4umrnLNmLY/iWKt72QHULNotBH3dFPBZJ3iBde8wwEG3SlZNoIb7/
kQ1y7TIVCZoNMfgqTX29xbiOBlBUR9Ffn+WbjghQxjWDuqCrH8MYB1DSybBX1vpD
x7G9fukIu/H6B5BNh3At1EA2HD/3nyDlUB3P+RdQ9Ko7zHmALE0h+V5SmsmF853f
O62wqCUaZDID36hoDial3IHOIth9AaGgPPvX238r7subrpscNBB1mis4HiYn06GL
xYA1RRWq02bMtJNWlZMN855KbYvxgBsrBnGbeFkXQPxsa5cmLnCyMp7/xwybiwpe
gXL9zK77my51z1pYnrjkAVCygxto3F1gGpKuJCO5GspLq1A8mUPrPRL7JYNVn92J
Zz0njpREL7cstvyZS/7KGiuSDVrxnJQhfHwJ9nexOtBnJOFYTBVyjRJRjrTAzDyk
cQ1fIVZJY593vNmAp21no/urJoKgpR6Ta9m2MDsoupAaJNWX3DSW/7ywZ70pbMkm
Piv38AyWXhrG6XcHdspBbr5o9L2Qj0TyrJaQEg5nci5BQKPQVMsvj0lxqveC8TLC
AJIcnIHq+Xo/AI0jQQVtj6LP3AvCSCWjImdeOGjXU1jujv0UzFtBZ4nu9l8LZxYj
lf6FqTGGHuRSBP8+TvbGbM1/zU1QBuWWFP3ydqJsCDCBeDxm0+CCWLMYhLLY2Hzh
4iUkKHnZu1wLdgDSgHH+DEPFQ3hs2CUTiTliEEi0MZs2wp2PJTv0E1G3XXn35d8K
l5A0YN46GekAp1JuWIvg91HgoOVsXAcceRFxCKcS+h5cPpuSzSOv1CZ4Pq03ZMTZ
AezFeelrGYb6aJEFBE41/X98yo2L+OBZQcKA3dWRdpk6+ZagxcvDAJcvGYbkX+HZ
/GJwuoiEv6bVequVKWjE/bAOfeNP9WBUesi6iaGqrHejX1+29UBVzxylsBLSBmki
xp/9steoLLyAGafiV/CAc0wTp1Roc3IvDDrug0CpUPQr0qO0gE91Tt9xxmMEPj7b
mvDyIAp87cbOzZBjkh7OgAhvoZ3E5pE5HHud74FK1EirbWOI4/XqYrkDu6koHN73
CyrtpsdtrILpCdaeNNfvGGMQRCj4/vWI2OIQP9wLuxQZMpCtoxOcg5hGIoRYW70Y
22maXbki1pIjSvFoSshAHpRvaEEZaC6ANALE+zQxcOzJdA6vjY61r0CnfHVAVU8X
hdQ1cD5KIXFg9xRcBAWo/fbfU/JiZXJ+Mqt7V7EQqwAyY1zwQ+aBmNlKFFpLf8IW
fY8mKzBV/3erIAX5DSEh61B/ozQQ+6560udv8JgO7b9lGlpfotO42lGdeVD7SA6A
pCLJGnDfm8wdmDu2MZcAPoneR30p/pAH8rmuHVJLf3nq2M9iVHQVv9ZnXnX8sFSr
ZvMlzYJapwCTYMs/JOtZ2aszj1VxGO64J5gW0xThkpiesHQEByMeOI2A7NhIW3iQ
fYpgx9lThL1SX70JsBggHiRiJF4WhmAKXv4ejxesV1ULgM9nbGB/PvVeW/2O3VlO
xdkeqRtzCxeMXzaG8VDckOy0JP3dM6tSFKUevCx1RqYW0vata1NkpOds9IIWxPZM
Yu9LcJY6zLGUg2d2vp29JTlVLkNyYiu2e2zQ+Fo9Snztlxpcoy4/Te/VEoiRz2Se
QJywPZpeb+qpWYelRvA+ZpYk/Y+rZsGUI976kdFrkLRmxK3yooqsgAs+iCM4rzi+
naok0k0olJ7t4Fkj75WRLhRnsDNSkgt2CNyGsnYBMQHZ+rmA2EdcNL8JaKTRReCh
IjQRGTnuEA9m1el4+65u2pHPQK7yGK7NhT4t3RqWoLxoWZRwzS69U4B4oOCTnCv3
jCEISB2iOlOh+aqxEPNcbBZRDWQ0DLKkbKxnj3IB4OTzIOgF66KsLFGsyj9RKS0g
O5sbt3i3mGrk8FZLqlw0LEhc8PwMfWYAdOZ4JPYh9kwOpFQoXsTxOotYAZbm+jyk
zQaArdbpz8BdmwrOopBLb2C+pI3ZsV83V9ZuPKGn0pqp1ozVr+Pets9IkUP+FSsu
Cf4dCgtcjYsGaJR6CL3RkWBYgVxAgDLND/ipRJJnabW9TfM1+M0i4p4FXdirCXIL
y0c7Q7fw0kBq0w0d1FjxFG00PJKfR4ih6p2oDybSb4o5q4bKr2+M2dqFWi4eVfpq
dK8K1TDVAcOMhsBiesejeMAE1EkWzVLc4O8P/n3FfMlypJ7X5oJmqGOE2/lUddTr
YdGPxD5y4NwmH6Q90x/r+oVukFa75MQQmZJ3YBrvMFuYMvokeUjLMobacCb6pxZS
uYHAqKDFajYORVGw43k28ceLfvyRZ8ajphUqXWxRAUJFbQ+bt/gO17U8gCE7sJoO
/gD2UBrx+7obbSUhTRrChjSwn19Pybc8jX9U3lPXHGWsfT3MrkIKkSuO6eMhTGJz
sWmgXt153dH4oHjQsgajieENO3DPEk43m6UYdqqY5j/p2vDTuG1e800nRv3Irzqx
rNFfnwLiuxgQcbxPtzGRyyqbz6RgWeh+NEJA/sai0ZmHWwhvcG3WiIETaZraGe1q
j48rguCDpSeQXixVxPxeeRgslU9KJF2qkyQ79V8kcGV/JxJAauTNXjK1EMBPCSPX
EkceHkdXoVtYf3h3HlBpSGj1QM8qo5QtUnsieK+W6n4BwHiEdItEDWRj4erF+Vq/
zy2sjBAilUrodIx17NSu3xDh6zOAv5m63JuTQsBWWTejzLkoFid8WzgLxgoWpp03
+Ku+XDmRvgfs7Q1Zk1urmI46UGo36wXsWoc/WyujNJwy9oRf7M9LBSI3M531m7EW
TEVLft60F37IwNLpucMDhhn3pRsCGDy7wcSzwGukarRW4X0nqT+xIuNalTwYzGdI
u+R7SjiekK0t1ZyS5aMFFaAc73isecITo2mWlbcExP0LnN3bb8czvVwsyBwieXpf
aZeywy3IHiew4F42/mV3M9HkorvgNCPCJAY6J4hhNzX8nnW4yMWxwJglCNH98/qN
IyTObe7yk6D+WY4qLsvEoUJT7MRcdblDBKHUs0MTw07ToqhT2tEmDEoNF1uxXmL9
SF6F+G4dle8/FznCG6gGH2HQjaZxyEdvepnbmsc3O3tCyyxcTiTIIhmDFbbFoGy4
cfcm4dEly+66nm/Yjdp90Feddv1bBDuSKyXlIipVm8GbMDm94SKzFRUZBjv3ckbJ
EOWMArqq1FNqeD8R7BQbdKnnyB2izjTp6wYWUKB5nt5UOv06v/lwDxHjZV10v3RX
zz46YqQQSeTFr+pOm0dl49faT8Y8FLIMKft+Yex0nPdDH3Wqe8hVbphD3l1TBDsz
CNr5SVQOtO2/1WGMLX5xnADd/6Phr2W0XanaQVVM7VASNowqmQ5l7gm1yNkGXXpf
/DmxOlixYPDFXBinYGjlhOMQIV+iOqJxE8Fn2QdTZ8sntScOLRAMH2bx5q7dqvXs
bcVikcif5M984tR9VNymLnbFJeMxcWLrhdlDrNJmxkb+nnPuDaV/uqsWtD0QvtwF
KfA1y6hsHO7MS++xYW/ApneZYBgUGNBqGanygVWTD9vhpbR0EMd+9OwPd5GQ5AKe
H5olsMkxfAjHLlFGspZwoYKx3sPFewPyJUEuwuIF6L5XM1V7w3yMzITQkl8ODE9n
PXb1IBNipcjD2s2VoIEejLo+rddCJN23kwG7qX7YTxZF6EnERo8nU2f6eTmHR29/
IBvY1cmkou9c12InrSjpBvw1STL7CP92dCR1grn8h52/AtvtU5xhaCGVyZKnddqE
J6VyJF2CGsT2vTUjct3sFZXH0sBI9lCD8cHPVIpre3j0Zt5jET5q4gq2XRwGbeQq
0XSiJfl0ixBDC75DVd44unQWpoY/r2ZEW/Pwr32RlDIcYlJFlXZ0xgpMItMD+wC0
OIiam/ItXO10wldX1kyidR/HpTYaGWEinaBeectrstjTzhmsZSLrmi1ZmKlv2547
WMgQpMpWCt2jcifk0Lras+GUrmU7gAn9XxShmuBDo7hLihyKgPekq4iyk4LpDpqM
dZRYpCMvKjNbj5DahHK0rCCBzgQN7vqw1hEtlzrinlO5faZLSoVR85UOEzbn2Em8
Gen8HmAiMJW2iPf4a8trkedvck1ixymDg6LjTGHW7PYXHRN+L9d4N8NaiMp2/vo3
QBaKHZfjFZrtO6jjC3w9XfUkv8ob1WIMwfIJABiHx7kFQNtOCzSW05lkS5jphb3I
6ehunQsRdPodHlXv7wNB8xmUHrKKp+vzbJSrOrKFmgyPwvJu7I08kJ/MfrMywTc2
NJVrY0FE7h9u8jJi3LyyU/XU+uzOx4K/vlVLNHVX88OZ+tuaclHJJiFmWSWF5xgR
MM/q+m5jH9+Np8F9G0SYoOZYQfREKs9cSOKCSQNXn3p8kNJGsCa8Z+PzITuUNA08
+SpxPeHuCPaNPXhPpFQ0Ukfr8w5KOcg5agJehytUm7pOcm5anyMEnnTTWhpjJwgl
vICb24/D2BEIeNj+6k1Q0CjrVK+Qdf3vDjg4wg9kHcU3KR1uUs2OmN9X4ZMc6eYe
RWayslgLngoOWjbzd5jgN6xHdBDgSPy9VIOO7z3j5KPuzdtN9NuAHCuv6aPv4y6Q
k4bBsWZ2st7Z3prE5nF1PiiTQ4OnfAvrYdgv+SdPN1utm+ZtMQB0qexotiXzyKN6
O4pNqtPEGa02HnqCquKUupiVJSE8qbKLPF5URKaoHc98yJKPdKf/TUBonTroIgN0
FkQTnnGzWuT3wh/aqlFH2khyPVPNqsMTc3j+euQ5T+8uf/2DOnN3+wE7FEo0e5Fl
z8qBiroP9QjAOGJZpEKDKfjWmMiCIP9vTcYwZqcf5Sk6xiX+TdESoaXAvPoGpwvx
XAHojgHRK0uJzK9cyV6yDvzZ9w4JyZXsxHyNcyJYGp8ruS5dnS+4LncwH7Asa1q7
g4B5DVdaIvLaPNtAyHyHeq4ZhicLLqyRaG/4Dn4kGOdhUfclTw5kWiDG2L1oJf/+
jSmX/DJdDLDQ5VeERuTNDg3MoWM8qhiLZPnw53ZYzZqeM01lVyW3o3L7K7FTwfYZ
NL/qTYJrhLdKuGnCt/yweNWXdoWxH3vVYfFhjSlwtx2iTl6veEHFOpmx0s7EaVub
Z99Xt5Hp149GWQ3jP3WTqKeHve5lwKay5LEY38AlBsy6o83eJPUDrelYZbmAQe4s
wcTrLH8xskcDK5zbgQxkSHYJoVSDPuMFCF2MqL+VzcCGuMa9gskRFgL8Mv/GKThi
gcD83Fk7cy3KU8xOyN278P3WEwdf8laXzQX70uicO+RxEO4mMQLlxB+Kvxbrphnw
w4la+yZB97ZVWn/3bN6NgS3XtDpih7eKQuwI/rCVHHxTcSiX96fwyq3VmYH9l1ur
c6nI2CGbydxlZRgoi3o9jdl2yf2fSj6SEPnHQP5AYJP1UzctJ0YXQgfATrfUFLM/
+yMoVveWzmYFdjMHBS4aNVn2aRgCWmZcR482MTPBbHednVMUSOm3LHkH058GS6Ac
R1JaTI8cB4GnYsPCFlsEafyUxzuD0uLmara1NNU9/0kkezJuYS8JY5DOQXA7c1J6
nOTPQaPp2BYRkRAjPoXBCenOUPS3rlf+zgBTzie4/oEtEO6eMUGD428laeZoDyL1
CjbI0O648Fpu2Le1fLAk1hkuuRhaO3bfzMvQ8Wt5wYbDRRRTPIbFpfJCJyRUsTM5
FcDq6Dxp4CLoobZU0tUCpnWoW/6PWT6xT4bfqjV56YP9jR3gRyKF02Nh083b9PMU
uKupOWZw7nrrkrWTRmd5PFFk0ynw7aU6kbwfqehDGuymtEmcnD3WKKIgKw/xztVt
84asTddD9tNShlj9PQKhRudNQSBvqoH1IbpqCRO/xwuzMDZCB1BgAzhx3nBw1Jf+
HAwkLPsbt2jIKAOuRkBcDQ3fLb8Ze9pbR0hghRfNbdld8wvsEh90Mk5MtHqRmlWF
meRYb7mChUHyy2r4g24O3/BkFUU129LzgqGXCXUusvlYOXoBOYPhh4Woc8YxH0Dq
KiFn5VnviPmc5KLBQ2OwcjD8wVgrF7V9E76tpMW+yLqa2OMsbQGQRa03uRA92LMM
wgUtlBWb2d715TxbVRBDwUidMFsmIdnWmwDINSpRDDFMgwSLg2gCWeT0hBbwbJm0
M1tBbIxOxqnfWJFr9ajsxMpmpX1+WKBnsKu8z/N8JVlbl9Qe9NRSyNb7zKpeveeO
TbEtRuK7fLS4/YGRlKWfa1qfnuQsxc/8mnWiulkfjc59wue2tEZJTg83UzWzuQI9
dKkZVBYKPh0MKkGsUPvIX9lJM3JJ+9oNk+Xnds5KsPAkYKWqs/39ByS27rCSGKo0
fclJfzxulUKavXIgjh91/II4D4EmhgNARM/qDpPfcY2oaTTP9SuIOhfmkeOpF0Oa
YTsRVwOCfuwEP+AXI1PunLrDkBGKkJ3W35rDuxpLx0Zy3YlSgueMAwGvSfwZ5E3p
IWC50BtwmDijVWNx4q8a1L2E+idcDS4atEJi7PGWzeV+/WBLPx3YFEIr5Hd0ewbH
yKAa0qGS47u017e+q/WMTtsKGVM4HhfeKflbAoYQ/8DuyFPKb/lzojHV2aw3qv9F
phgWa8WxegrT5KtCHZeZHPHEMkTQrR4zLcdyW/YQrhy5HmhBydMr5w5XkAC6A/ij
kCr83cQ7W3XUz0PYCnX51ahdv6hTbiSTy8/QKrCW+ns9YTCzgpLscyZjsMCnQ/F2
ryskxzMGEeYVduU/5PNSearA3DdK9DoNcxClH3n4vqs8bqCgMdbANksayzNQfovr
P5cPfFO/5fquEJFbkGsKjGJWv0fK/uuSe1uLMGTl9HzebE17JRgygEI25hJrayqw
WZS3l0VJcyEnw7BTcNp98juEY7sk4AM2X4difpR3JbQkwzxwz2Y/Eyew6JkYWWN8
K/1GfvAaAW4Bkt6wmc98OF6f5+E2oK1hUagh5uD1tQ/rjWfHx9sPNTHNiM9HlMHt
eSTvC5nwrjFwQgDaeC7NSb9ryyfTsUy+erd2YEoOqf3Zuy5nCPgrWhtk8R3Q84Iz
yDt1+qIAaA7sLrfwSL7YA5+UjpbkPlvLqFAEbWsn2zrzaamWL/DrRk741fOUmhIP
1yRVSBD7txvmFJZ0uZtXdR/PKt2ziksIasPs+bCrntdTMDaIxT/f41JLXm3af2Ca
qBvx74tDHWNJ5iBbDrSWSiZ+Bn3YZJEJqHqHWE3Lb7HpSrycO4WeLW94uyOGwd5z
VSm26PsMSuwS/Zx/4gf25mphU95nCDNFldFwOwe9Vq7rT0dNLPMLlO6qjV/uP/Fy
oK6TIOBkO5ZlZ59XAqn71bPM9ZJDmH+u/dGkm3zN8G0/n0ZOo6elaHZVut2XFE0r
qr1AHAv58s4ZqQTStUa2TzWx0BTpqqYy4/yE4nLgK56p4UMUJyE12Iuvflak6aOK
OLmIn/2pgzTgF2eM6/wpMsXLsLg4z5970vXyPlUBKnVv2DUQ3I7sFCiK+TkqO1mj
FxXwJHVAOF6n9dHfBkxaqsvIl4D9rDBxfgyCLNRD74GJ3X/aYX84j/cWw0JNib7w
x1DOWzDC3SSGDdC4AjmfQKCloaOWKEJX0QJY7b+k+678R/DlLHro3mR83RWhJMFq
sCF0VgH/I7aec+TE4FXMRkazrtBrf7dTDFV7aFBNkkVDmwIQD/7+Vq9LHp02gy+0
tb+xPZvVXAjoEA4j4JYR6rTkpKcYhBdmT3jxIW9XtDUQJ9OowyjVFZlD/GroNpPS
UDQ2Ninb1zDrNzdRu5iLhWnHvMgIYbkvyBjy3MmHy9DhBXxCCjqJN5N/vGksfxEa
xyIGKdcuLJihVKxtb3I64E9nCwOVmILdgOgmbU8xrYi0qxSMOu2zY4azbWrdWW7h
D5gLSLntzi1+H/19h1A6ffHy/GYGx5CBrD+z6c+lJ9FQUa8/qt9myAmwGii8aPYo
A8aDmzWIgAv/i5nY/+cGrrtTYEA5YX/VqBwWj3KWW5ptTGVHRTZyBQIN6zADVomi
RQ6TA7BtaIuzU1oJus7O47ZLMXSakRfvrRLj6zPC5xvnWbGjVV5jrUpPoaSV8ofc
eR22q+arkhSMgd3IhymAKcBWXx8dhUg/zxAPRn/CUja8ILl/Hptisotkvs/cBTMJ
/RRLAiJG8PtA16vhrJ3FdayZWSCelMMiAHaVpNoUtkbIq5MnuCT+QTBqvrKPmuaO
L8cDY6oJFJRLnIHSo7d5RCA6QaHPx6OQBTinzBriOhhtwJ+XtDcX7IqLwiSm406E
lkmfjCNePUx7C3TlSKgridgIrm1T4AM1PhgUblMNYdwwvSeS0nra2CXe3y1EWw1J
luWvlbaSTGIEs0DycOE5SypbFihlLvmvhPcIuU9UbAcvSfuAxBXmzcoN32ao1zN6
V36GJ8j7+1tg+l6WWAnaV8aReHy9KTKeOM+0eXVE+OvIdZWz47uMWAO0+4LrORH8
XMiZBf31MOZneJkSeGWUAmD75rkd4PiH/gIxSh1kFmH21j5Uc90e3miOZc4z2cRu
8yZFz361hHv6BeesqzAyxQVAeZ9Ki1Tkf/oi3QBF2cNUe62JX85R11xBYGwyrQ5Z
p4Kfg4j52/aE8XscvUodpPPLbCgwpZMnnXnEN8U46g33IMQEkDBnReUneCXkmxBK
vp7gtv3csBKq3dPeNYYQpLsHQmTmFoyJ2AkuKEeUftv/qDBy9XKnLdcZFHbHL59i
ZwW5HeXMu1i95bBQENBG+D6OM0cxi9UsolX31YFuU2QRiob2H2tahE2hKJqO+kBV
sAh/EDpNRPcgaaaasKFsl4z2hm8GjhvmFJckz65PGKhctal8eXIw6V/Xxm9np6mW
PHuXyw3Wa9Zhm7xwUBX7ppgYUFBYMNPAmMmhMwG+kYXgGIbH1GxVoVLEQYR2o8Pt
/ly0zd/QiAYrr0KDLYbc22c3qT5W9V1ygO4NOKfICcnL/+mWOzP5c2K6UuBNOo0J
eF9DsooqZMGxXtCyc22w9dLuBdn6FujMAXSihbbH88JabDP7QpHdL77Cm/qvP1k1
Sd5ZZGIDyiD2P41TKtOxM3NH3KW61ZIKlXLzoEXQUDeDprmnmclYLKS54e4iI9Ww
ur1iDNf88JL8LWgHJnCypnHmqgbP3xmMqrPlUl2HjwZoiPtjw4p4/GjjE0VVIMFw
BrNq1CyDkoR972Q4nuOrp/jBptM5OwFrkMsi7N/0aYji3lxLnrk1sQjjT2yNZ4Uu
69ho6awyu7jWqQS7LZMYH6hepjyYo5orR6qNIyYO5zjlqoa6LT3wUPU3t8hNh/hr
heUzXHmxc8uNLDXat6SA/7TdQ+SrRxOO3cr3bNWExRR4QmyvdY329EvDg2Vrsv+L
9pN+k/3G9dR0FY/nGmciqmAYyt/J6VA7z1rb5IkQLSKioiFLYs6MyCSzdSg+AFHN
M90GKgXceyEMObK35nekMbrl6zQENQjeKM7+5n0AleOOcmgBxsdLENkx6xaMaKyH
LJsdQVQN62jAgokWdJ+/Krmjbyli4dMNAy7dSs/SHwUd1JkSL7cPjP6eUKzLIIGh
s/4nKOBF3i41RrGZLATbZZHtZDzhKnO3dL3y/aw6JFG5Ak2Alx4pvLfMBFXO6Vd6
dlMFYismSqsy1cgiy1nb8AHndtFb06pZuoL7AudjtDf7Dv0vzpeD3ISf0Mwo1mdR
phR6ard7CtBc03JOpsFsvTIi9Uh8xqhp0NjajY3FKa3qFKn6cUGcYrpoQncuKXlF
8qKSouw5sKgRG+zyYUTw4zRaEhXXNIXwNbAFASaFjyCCNqRIouLm7Hm3uxtSO0Y1
oSkYphzej2RriO7gwxtV+Zu04+dTviLqK1Ur99Qi5qRNKRFPZ5SZbgLMeluo5Eri
ofaec05ayuRJDItZb6GBw5JConUnABDQefQbqKZ+zmnMXMvnX6lINW3ebD6QvBrd
d8j7ZsyKHTu1GQHfiKhKAfakUIMaShx01bipFuQPCzb/SOMgCGJAYxZvZiTY2Elz
NoyK28Ohco4obZtBHTJuF1ACMRyt36Faxt9NHnrHtEcEJSwD10Zgy9/sYOBoT1KA
wvoVnYAxjDA+2emxV3gsFXmI26JHq0leR8e/4ts8K/FuSIJ5MiZS2ccBk3cwJWeO
S++Wwr5vQdWjLRBxTrzQgeAeKtNyFmXpq1p5JnLNE9JLDrCZGQeKpSbUWO3tI/5j
mdRiL8ywzOx88/rPe4iZDkySRCqhIR4aZ6Mk1pi+dnslgOj7gMGvl0dkqPufSUFC
MdltD8NeJZTv9SF2GxCRvErfD4F85O6qt+yPi1fDuCbTwjOy3dYLuEXiXY4nnAC5
a4uDtxQdyzgi4/ZEvDx6910uzDvBANvjgSgvSPevsLZNTMq/nDurAttHJzOdcLZR
43sGm/Ls91sAWyzd4eDg18EX1Yn08eNwaVwwUsCCX3tmlsaRh41UL9cZLWp3yNzl
8YWTGu8+1DJp/9XIOByGNivvVEM6FfVzyhC9KD0PrkQsJ3n6nIx+fU+zfekeSbgc
R59a1MkKvMHMjlzdj7zCV0e+tK7V5YObYHL7ZDN7Ulegq1BadKUpMcJQnFiqev00
MTO3BYaY9Zs4nu5Wk30klwBfHGb9Y98wxXQymb/P9QzyeP7IXXqzKhEAF0KIbnO0
2hmWkZCvGD/B2bum6GYaMkUVWCmxHlxldtr1+9BnYEiBarNnv+sm9JIrf/SlJnRD
8oubyd2g6zfPcaCdRm+LkjUJG1mZzbpWQ4qlHjQRab4Q2DqkkwG+v7p4OIt8AkVJ
oeV4WLB4Uxj0EnNOo/pyeco3aY3fWRucAdm00bm5VaM/YyBdXp6FIhCz71HwMVNS
V3C8DHa0rObNdA40MIMgCvEB/vXSYVZbAXHEloyQmXm14VX+sitLcbieP0LlmAfV
HJtx1hnNyjayk9O/OIWDvP9/O66tz5tI4ZXGsmOWkUdkrALcybMJj7N7ajbh1qEz
XrhQCGGNCHAKXXXNhynrJnK0+LcLvZ93x9xlHbtOEUfYOh4+pFb9+AENgCYQZ5ux
+DDLLxUPqYOqGmwrbVaiWu9xKHZyEXyHxX4HqTqbOoPR9GqCoG2jmYiBzjymjE81
10X2m5toyTyG3hc5oxLJ+pV3g4aYQmxKliNVSV3PtqnATcy40LsxQxNbuRfWp0Vk
hmMLGlM//F8SeWlGZu79YQYLZGFoceh76PAF6j5Nwk0BipkoO59CjoA98cI88bkM
VkCJLlk7G4zA85pXMnbLhdTErRZGI4zsGpsobbFDNXJ0s2e9ytQK9KAKso5Soti7
Rg1BvRFRmc+P3EPvBwhR1a4mU35Z38FD28tCtNokfm4WMC863yKnZZajx37MPjIk
hqyDA332dlPieCTjLyai9AcGzdUDC9+GyHzqFAV+wTzRH2dygSMDQwOd8n4e8lO9
d1y5XlsGSHYQc031U7cqgLef64f/KHi87VA8Z52NoENmo9ttzU5XNPCyK/23yd0i
MJWVoyyfyi46pC+k5qyqJKuEo6+zwf+iYASZTlC2oeZDPMEoccptEL09skbb3G6e
gGZRpQK7KHK0n4SxpOFixg8UVI0QXXT+VMvvqbXxj2kjB2JpJbm6w3L9CPRb8xcB
fTA5AvPNPdfqRE/yx6/ltAOPx4YsQKHRtNAPPiBPuETurvMbJQtFgLbCm6Hd3mTn
Cwl8MxvKK3dm1IK5w8wsbLY4XR+okEm07WwSnSqSH2rLMivOmp4XwE0M1q06X8R2
4f/7qU4aJ6lnoP6VSP+NftgoRYdFfzvkexKLlgoM05R8nEzE/wh9kGBorMoyDrn9
7TE9tsMfQwBaL70MfHzyWBeCXoLqX+8MbQbZmYTyALwxCzX4T2sVPRgsrF3mfPSS
u6oKdIb3sBGSM6npG8/mZcwcN4rrm/g/4+MIHJnNY43uibEghoFrAo68NHV4qThH
ZQI2T5WklZfTL8/5Z5+q51S+fITz8vti/ToZ1ICsZMQzQrSKTxujR5+rJ70qyOZL
PTerrWiG5VEEIvQvrDnL20AU8zxbVWNGpb5MPIDlEwwUQwyyej+cuL3/kyLLnh0c
Z8XShdW3MrijBm+ZAvZQrY21//ZyssE4gQGJTa1aY85IryltxKOgY5qWw7xzXLpv
HcXUiVghIEOM4+vfEq/G/b7N/p+TJqHw1JWFVr779Au3bHpc8I9/lUq8XTCzH62R
wPzw2YgiFmvsd6pzoyZCubPh8YlalEUsB5lpNSgzJJWwCseOAqyLb7oJAO7VWiMB
L75ewY+p9Y85gfrLWBHVE07NwxoCxiznPcoHW1RSNdReBgEiPJbL1wV4FfvJYhYU
v1uUpthWSQIvYAhl48ugQA6XVirgtzbc5KospHztVHdHS36XCHOEz+7P5xBXGHmj
FX7VfHCfz22QQZjZdhfMWO7q75Pr1EoFLwevDrexRLHZEyP0wyO4GCB7sMTzS9rp
0gfdaF2C6YqZ8RyeEuasYHvs9vvyBDMxJs7VTiOCvWXejnSPIK5BkuS1lW8iWBm9
KT15XmaVFPAHbRtCXpVdYO0DCT1FI2BqKInQfgoypMLRyFPxgFGbzrsxrAt8uM7i
OIPG6UbR0KWri8vvCPMa9JbEqe1SqjmqchGIariCsUwvFZeII2xdHTDVLib5QuOi
H1qoYZJqEUFvfI3jLFY0bUE6RzA171t+WJ8rUc1K0cDCP84vU5Yv9h//tB2pTQRS
obTXudh7KEX3CwKiSNgJIXyDwTT856AjtFMpnLgnzbLNRR46e53ZXV5pKPZ4LoW2
vV9QQ+qLCf9keyziBL/+vQgkIc6fNInD7EaHm+s04juFKt2QebuhjKkoiCP6/ZoY
Ps0To4oN8PCc6jbCRpKwAma8cNnSAilBiADyEzCou4H1xKeX41n5+km+ai0yRf/4
DFTy/hgmyLz4KgSGSTWN3bwd28Sz2NgnU+3ateAMJfDGJb+ndzT7a/WvDlEA3rIW
nbHcO1vaGiK3LjnTDaeuH2I/3O3JXg6F5+mQFp0c9MuWyBicgFO9l9yQsdYPZCs2
nXB9+dDhM0mWHAl7dcrL5dSSFv47fhIQrLD/ef2OGKNJsarQB60Sk2pmf6crEQdN
8xy47SFPnykxp58iY5KYOvee8H1PvaZSSMviuP3Fu1jDSbdub1N83ehOPsyXBUmt
Fok0eMvWdYK57ttE2UEJkSlytUziI/noCdGq8xB/fwkzeVgZqGqkf5g7DDJhwxX4
g506vPl7hxHapfDsdi+v4FG4YcBOxVFtq8Au2McbyNHcmTYO2T6RKz+8wa8D+r9F
C5XlEl55Lj7+pO6Ueow/TQfRthuunEQ3SSQLam9iDnNFV2ygA0/l4WtImhvD6l91
ZNPCXXy+cXQgQIVIb//0taVfT78JmhVzM77NJWmiRIXemp1w5rUcYqMfK6W2T2qi
EP1N2IpxYn9s1Ux80aZ5IqC+RnLIANI58w3b6aDpqbJfqXsK4w7KSXjBMmlAhN4w
wYOQ7HyGa6UyymVYsq2Fx0pW1OdurPjww2cNrowlfBOz5q9bJRtYBRvA78rHJr3c
rsrzed2VdelsQmCb1e2IUojgbPCB9PrQZGplUHl/JGxwPHa1BucD8uvlvJukDZUR
0/NMfgbboODoycSRkPj5lAZuyStYjbQVqsThdJAS4HAQG7ouP/Za2DlDtlSbL7t1
h31A9EN+XbfTY3MCl13tV1AJJ2VaFBqTvTlS9sk+81pRHEQko+Qqnnt7B5Gh9rYO
tJZjFalmPUbYSBMw+ZrmIYrnSDwK8R5rT6vh52qfmzhyb+ybOJfs6OMwdfaqf9f8
MRNitzoUj7ntdi2A83GlOgdcNOCLlsr5brzRXVHEGbwRKiPMAuVLBswrdm7oT2cc
T/Xdgoz+IY6T9qnP0vjnqeWo1PD6pn60FoeVeh3PUTnlSXZMqkPVr4LW0BMphOs6
QWdEbH7YyBIWDcPJfjaw5O5pEGRg3nbr4HQTTdqo4iOB7GkDqsldzA1Bz+7FBnCZ
E01D/TMg4JjYnrsnK4EhA2eF3+C16rEu74uvFccYb+clASorc5n0i15EoTTYu7Q0
JUNqo2T6pWPJ7FP608GJz5HDgXZ5UpCv0NXoQ6SN9CeJ0yMhIYJzGq98jtrh2+us
l8uro+HGkeUX/Uh2koJjjjjHbI4RitqGD+ZqGHt+BTBd/zPRGN97W0JobDnWkNYE
7xdD5HlX/J/ijldViuxttjhrnI3OZUG6uNzEQR99egz8xtn87xn+wxGPWlt9krFy
ZqCfwW9Rc4G6jq6T9VX7JXODEi4h5jR2MkyPAk2kHxMOhSHvrMxH3CDK1iphmSw6
xwErfcGLmYulpSEGtb6LohAcENa8cYfA02FlvPJOyT0ObQdMVh3MK1Z5ic5QrsUx
eIVXi8vjNKzQDJR9rw8uT1Gb3c6ryYx8xDlDCgvdF+MF2YMENiDqD7/BEd5r70oe
ZiamVJTUW2EwWJAhNjOqAXYKyeQV8KSob0WKpxRxLD1hgr4DHoGqbN5qrd4KRccu
69FMEaUKojnkC8VbS+fluKfoXpgHtoNjKS3B3SUvyQrKP945cQBKMmbYcy6bV8Pm
T5dlj9S7Lgyek/sSdmQy2jM7cH8WKuRkGYi/m2uB2lsk+6JXnkRi6v/Ui5OSgPSl
f0VX8/cWj7ua7ypzoxUw0tPyJK7CVsGtnTtU/b7+3CKLOHX4n1h2ObJVsWPR2oHU
a2uTOSLIQO6w6EUMZbpHBC/89St3Opz+t40eKGLIaSoJZvsccwRO9RMCBoH0SPhN
u85XrAOH1LT4be0Cm6ZB6HDp5QgaoKVTi0oXmH7W6CrTP11/T53gQfJquJB7jICj
OWpjqCPlBStYi8rLyxm/MW76PhG5VYIS2NWK3PprgifODrQ2weqm13jQD1YXOsU6
QlWCuYkgxrA9GgjYxgRGB9dol26gVikbFfAaE4AnvypQEJfg/L0/+TZNDrZ1tKt6
0ckFfL5mfPPgxsdT4S68edWCthFhxIgiBxxCW07RphVkpj6QaZ95C+Xvv7oQ1+xY
yAuLl9FQWwFluqS9vKWIBo4RDa1uApJ963XIGAOuNns3PvGw7hZMhztXsEifFjY2
Py7x2nJncJTBJ3npiufGbOkvPreU4fpVUolDPjZhXo8+J848tlD0iPb9vY2NTJ2l
83ZrB5TClc7tCHGyNBgtu9hC3KbRrcl+OI1b2YD0aWPkbbA8Wbw8KSXz9/zGp9Su
//giDuRFG6cawxpMulP8+C4kg4Uipcsc4Hcdni9f/9vZnDMJLCwGl8t3JsxzbVei
bYXtY1gTUn+GsT9PJx7CFkcYKl1zymSd6OPb7bdOUvR83Pjf3QSYRX++rTPJvNid
4bPvmIgCH5eRjipQk0WGSxvqM48V2M0XGnq7UAGDw1JRIEFV4gmcTG2grQYMUXB7
VDPlaw+Ozdqck5mmZDvCtIDMBoWfI/tbo+LjPq3ZETbTzBPOOIwK3bp6pD87UaPU
iZ23/O3IFn7cQFpIvd3G2FSZwrpbPbcxEDIn1af+hk8vxQW6sPIMI80hrDPbz2jr
oKCIwviK8v51enN5BQneJNyKaU+SYg2dZi5oqL4N+up8lnxYQhiFvvtLkU7coEgM
nqHIidQetdQU9TAZbwosFBn1IBkxF8qeRQzvJjgMhsNjJtQPU691+DMS37tHrNQ4
ic0WQ+wekEwxCl0dilVyMccYoz30PgCndb2mKnQWpsWLgYtFvppVVkaOcCr/zy7u
CpwknIFSJTq34CM/RKSkEFUqP2vdLdSTZh8o2z8DiOcjsfxFArVuJ9C7+Ul+2CUu
QOefeMetsQjDdPd+Ay1G/EhdAZg3zjBrXQFJ6IFCs30pYOkRAHQyzrHoR7mwmySB
bBfGeBAJ1ACAgs2eMweEPBal9zFrqI7BgTw6mJ8Oj9PeZHJNxRu/zKWMtUqE2lnY
lR8V6/hZ38L+zIYe+IbQzUSfa6dUF+zCnHnvR8tYMe1zLAufaOycT53dZuU0PRzm
vpaJuKuZ/IjRs1g9O5+DFsPeaGVsoq6z8qcfpV6Q2awBWxUeMUJur4wTpCq14PQa
KC8431YdonNIideyRct86nCzBuC6RbJfdKhICYSAw5GTYBui3qTwJn3em4oFWFgY
kpyWX6nn65cD50Wtl/n3q1fe4a2Uf2w2uF4yLff/GYV3ydD5faSv9Xuluj3Cg1fu
zXMSMuAiP8LEN8/mK2S7KgTNwGyGodcR+l4XuWeYzRR56Dsn7ifwubNeiBzoAjUA
zKKhtCpsEqxoaJObF34o/IrHy4cnW0lI5EGng3TlMzM+Sjgu3bU5NLaq2Doc6u5C
0FDCCi80/dQLUQT1swul12YM0C2Bq5gqfs540DQkmxuFtdnjD8zmX5WrkvCgAwZF
1J5bif3X21EnjjNZml5UO0W1OP2EgaGZizEfyizYrnsBtz0KcwlWDnO9tTp36xKQ
rAp0L1hl0pFkQjPMwPwQY/otBS9KPtC0lxn/RuY7hNCrW+tgS/Bfdl4g8j9rGo1f
rndY7Zo2MEfK4Pb10Gm44PSGGrXSdPQFZGOgqVdzSymgZ7Zed0FfNMiIwXAsODKO
fVxdaEQ3wsYr3peSWrMVZsJTWpSUYG6E1sv4zDnkxHYWsmy1CdrM9whkuGs9U8yQ
wEdJ1MmcS+1D1SAjWY4G8zo/rxTSjGGshT/gcx97q2pIA68Nsby+QoVflRMYtscX
mkL9tBoy1Rhi3LzZMbxB6GgePVc5dD7lNgi2RYOdPwh0J7Anr1+MMaF18o1zkU2U
Pd+w6V6bJixLvFuRkbU1gUIK9PLLcvpysAhRTxbBVMFMHjZ6PDZzlSQL8GjqWTKi
pJ/JaZtYpWYv6/A8vyU0f8FmReyM3YBmU3B1tNLP4B/szIQXlgtkQxYfc2gueeX2
b9EGKVsuaMb5OW74Idjhmsb3w+kiLjmuuxvKZNOSQIDYPBIEOaexS1KRyLlaP5uW
kyqKD01ats/qeEduX+dbozC/Bc2c5trKk5NoFX2IZRR3s8045xDhuS9E5shDX+Ct
hUYc3LUaI9pgtzSUvDSDOTAROt+lU2h047JYnl4PD190ii12sfuzzDYqFm0erMEl
UZ7DIpNuO8lq4ma/Rsd77eOc02amfINt4IQuJdZ5w0FQx+KWeUf/8ccCu24VNDU6
2/nPRieXoNZ5Gi6v99d4UdscIdj0twOz28qzmXNVD7/FcWRC8uR7IuVdg33JVAJi
tJKokZFvQoF0mPs6Zakx6yDQBg8mKZ40W0MHRt62ypxX0b3tt1CdWeqik+zO0OJt
iGzdCZKlHMZAxVQrf4eT9TuSNftDCL69Tkj8ez2g6zzseoquJRDO6w6IJKPY6KWS
jXKClEnrQyZVUpNicvA6kpcaHgIUpiXzdHR0TljCySkFaPXlP52n6/W+sHzKjdLL
Mkq/xVXXf7Z9fCcdWfqm/qmkHnFxuBIyivIZ4/5rNxMJUMogd4hhYtHsrEgq8p9T
Zf3V8kFRiZjGB2kT/73MOiXjFw5pUiXY/HOasmvANR6e8fy+pFsjQikrsrw5zhgm
n6o5x/vP2jVcgRMSf5TMBRtUU5VsI4LAIzGx3DCd1TsMCbTAed2DJvGu0nVs48ML
wQI6n+/TWKiYigLKmQHKCBLjJI3IhM5vDDLl1LemvMcbBydMOrxWdKdbKOUK1shg
i9sa7UWvX8ryoto+bnRyuCYeBvnqFNZzJVJ9hyNW4wI5G7sTUeScJ33jxHxXWZ+n
VjM9nf+FOfNyCMbpqTYKH9VttOzAgI3JQB8V3SnLnCpQ2vzAzsy6zKPQQxlRJNVR
D/9udv7BAhLzi5powgchiekTOH8XP9r/Z5bfVEH3tONPgkBU+2U33kc/CM7WzlFr
EF8z1CelPnwbIXe/Yoy7/e54x1wl2fLEBbRm+23qyuKv+14TO06Bg9eUHwt+QFQm
wouFN9nc05wrG5CkRr8HOGB66Xebp/WOq2WXybJ4T7X+roFQfYNq7dU6uYTWRw3/
FckIOQFBc/tGLYUO1wbk2xlo14eZpmfysE4gP1jCvb4MGQE/KvozEkQa9rO/lrSV
LNGuBy4MW4w3Q973DFYeA/ObDVB671a7SJtgV36Dt0UqZCQtzGIyWLLdUuWDroau
41y4+0/xriV+WrRMgHgdiaedyyieq7YOgQdQ6amzzOXuw9HC0R7FfqmJja5Fd/kf
cr5XqX7VtapS4w/C246JPrPCSPknOI0nZsoQ+24OW80jTFc7uUhhc1UfKQ4eX0RW
ZHrndgWkDlwTi7K1ZNf6g0/FVDqKwTlE4lfWOq8zhdGLij3Em94Sz3jIkI66lT3p
Ie2jml/hzFC1G6MLyDHRuR7OSuDcUZJhmdECBG63lq2U9vmpHzjwX3k3VilvRaQ/
PgkhIAjhLDCi2Fp0h3rmrTNlOeEFiyZNJsYSxBONh+6Ufd8jQEZB0XmNzRqJvGMh
We1S8Sbh1+C+fp7hoLVR0sOIvHAnrULWeekA/mbPSQ9zVRqP1Px0+DtUC14j0IfS
66m2I1kznM/ENPpxw0G2YwLW06/T361HKidtNJQaqDrWDOSOoqedPi7CDizkVvYM
/buZUp03xRGMH/ovNp/nAvlK3bE5HPSTik4yyFsGhFgVBAVOCQLc8u6l7YEfvsgI
kwAIvwhMH42fdJHkDoP7eLOZu62LYh7B85wPY/x8lQ/7cT4TSk8IEOvriBBFKZPz
6j/3axYTR1EOPKAuj9reyT3b46TFoaizIc+rlioT0oUO22fCfbDnpL10mynbTMwJ
Eo96qHl4oZA1H7wBIH2w1OnEfH0/ji4dTZcinjbDvbOlOqhDwT7M7Sq5Auzh6u0f
Gq27NkfS/saWRObvSMMbjvvF0DCMZDtFk0/Jpp5SeEHE6wkzaEAfhAY/8LmWmqhW
0MkSPMquP4wjS1Zu+qEzlTwY110g8MdOXy0uIwEmlTUa4soWsL0w0qs8PZ6tP9AP
SkRYuzMRXpEBFruqedoZjuAAfnXaoxFnj+O/0+GcynXZPBe9h4do/lpzg0fXO8Cm
BWSM6IqfwksYcsj0JKDtnl8HIxlrIKrbmICDW/hDOHDDNZ9qV1H2K1QELK+obOkY
4m+P7I/+S9ijl4yEtBbXCQaqdJnOIDJmR0x2DZbZ7t9Nfl+Psz+qFVzNxOg3kHD1
54RWbaEb4uRx2QqwjzxoIud8FxzcPdHgv9pM3wOP089fCIgwjCkiSfTPDjX5Qz8o
T38TTkF2QEkO4nkUJy8VaepBSTtjaMkog9+uhnd6gI04uXHUO04d1jvqCz/86mm5
lCZRafx9+oqufrOVejW6W05UEZG+CxF7IWUDW6MmlMYFCTPhjNxVlQ+lXo6vW6La
VMQ4skVsv3aLqCGb+v3Lk60O0sURR+juEL5UkGIok4Je3F5BL4zjr6Kgpd+MYNci
H4yplrbQ6088DjCjk36PNpqxIPpoB/73TCwEtAtxIyByKWcjjHI8CucfVVwwdrsS
8lb2V3yF6moJ21pMOOLcKxyVw3FN/IiKz/m0hV1A5CWfFBTnLQ6q8BSyuktrWGCU
Im2LLSwxETlTG7kea4I+1wdQzpnduhzMgWctgvbg4CQpxYt5tZ5mZYx3HEL2QoI6
dSzYwNmVjHTZ6fjfW0gEZh82bVXeOCVJdYAWZNMv0FAmeKqL+hIfKvotM5gX8ro6
TsqUBaSfSGgb6VeN/Pas5hBaiHl8tjRAeYBaY3mkjgYLTo2j3ZnRPXr6B43qJD/O
QSIaWWQbgxRRReF5jZlzp4Xz15abmYs7CrCaZJCmOFknug6SZymFOA6SMlkW7pyP
PMkFvE6CbfmqAacZUf2O9SabxU/CzWUija4ooBmVd1Xht1cxbUe1MuN+5bGobMQU
kvrJntFmG6WuUS3d2ET6fNSdSFk2YueLDEu7oVwVkqG04LGQRLRBMb0BkA0S12+X
JA3VaFsmVech+JrqM0+MYnz/12P3PMvr5ldi77BJTWEBEda3SYBaRHatmYGpzvWp
l2GGNBdzpeoJzTR7P3ovoNOmkyt6PX/lDUtCZewv5n/k7mGrmdLv25M3yniXBTCO
0xLEH7aluW9e5kuHttbHFEK9AqeaUUXOHkYZjBHGLPXV5z6rtYQs9rhMnXoUQmSu
hE+MQz8BWKm7ONN3Zwpo76H8dORp5uYdmChdAvzintoTxrQHAtQCAVGkJwoDDpzD
wZimoW+u2EWMt55rLCFQ1GQfQehUHdisLhn9JDjgKypN0b0wp3sCPWOYRvdsyJOw
YzZu9xMxc2ZBGfSQUhi5Li8OEcdLSGiJt0K6/JOc7ERduzwH2Q5EL4ItOYLKNSig
F0MmpA5V0uWUHULcgxKwNaMHRJB78sGvs22KQ0L3xZTsNNc0TydNhzyFt+1CxA/j
QHw+NM4NtUc8vlHCz1Yw+9cVBWgzRNo0H2N4q4EWVOWBqcbcHf22SlStHANoqlzT
ntNMusr7nBBdKAD1JhnGT+CkyPyN+G4E+nXRnzG/q71lXM48vZdbu5hBDGE10H97
gggEfK7tNblAleL5wTph+PpLuNWx6GGJG62n6lKi8sM4bOham+V+E+rSDK7tvHBo
6jmHef+CV7lqnMqZg4crW9lerLYbPgEcE+SFpLwRKpDxVDh1pt0n6kmgwJE4ttPa
4FAMU8gS2rGVlSKjeNOzUaTM0D2cpIkTdJ1GZ9TbvW25sY3TbuqYhvYnSPLN6gRu
gQTLjT5CT1/aq/iqIKBY+nTvDuG0ZEdSDnpd0eH5xQr3TY3xEcAivbg7CL8TTKcz
k2hCD9AwTXUoWDZ6xaRRGvVH5UyCHTAuGPSfWw4DBizizKvBilm1WuCfkH3VK3CO
54PYZzBqzzdlCSiAl0g8nElDLHKNsaeRcFMa5iVGz0eypx4ePj4ie0jPArVJVIhD
UJamk/xacHp2iCHuAZXh9ELB3wjKb45xe3BOnwznULmv3CPHfVjncnRBr+c42ujt
i5Kh3zzUbvRwhKONGMFgPVzOc1JH33v8FH/mJrlKwFBGx9Q5qzK7dsYpIjNXrWJA
CXoCSDNEj0M8sxKpBzmMe09IojFtWezC8yqKC5IzZ0bgULIbXOOoK09+Dc7nPuJg
mmnpMxBgNOhSaJymKixoj1yxiASeebdw5G/co14LkZEEHIvhgiV4DgDJL8YW4Uwm
LS7Dg/zPGGtiDoIZOyLDOfJyL7QrxfKddhY8xpG6oXmHzQwi9nEp8lbxysYkak8O
DxnMzbN+BargEd0ujTXLA/ZcdCqPjYPrXflrc+d0X39v9Q/uNo6t7u6D5b4DS45n
c97VASXjQk6Ho7Ui4e16/1pRs7pezmkhrRR+96irjS1qii5hISTXNoCl02oakepn
NyvgcNtHtW3aU4HiYPtEs5nCAJNM2dKQxUFnj7nyySzeEqqDLUpaHgiz5QCApUZp
xjjACz2ZJ61a9cLOWPdRgAss/9Alq5eC4YcXU6sK4fvzDKKKa/oqG7HsqWpIVYcB
HLyQRopeutFPrJB5O80S7svJf5eOIhuypeANfP8Y8m/mmovy9i4SL6rz+NDZm2l7
dc1F/AWWQ8rzkSwi1aGOA0TepdnTZ4wXhfiYKlIF7xZzN3S5YUG22G+aMoH+jY7i
UwyuWsuFJdEyRHQhSaEiJJUdqxFU7SkDmAwcJhW6r8iaPG+Pjm5H/GvEq8NcfsmO
YrobEXcLItNTlVwF/27HHMUd/mcRn0w2m9r4chNtJ5r2xtiElqT1dP2m0Bw+lwvB
3W0sak6fhnxecDxe5vu4iFrQ4v8Ziudff+wjm8zsIfEZ2Ui3J4/oCmtgNEtaDbiV
kzaZNBpmc1MjW7l7BpYHrV8nqogb0pkeOJThvsF9WObIPOc9qINpFEQpHYI2rttL
89wsF4lccZFPixpOyaeE+DQPwac+88HWJZNKN77NoeYt+KXsJBFtc19IlXnZ8x95
NkwfxGfJS1fy9e9TvkxfE8ZopacuwhuSgr+T4GOkC34BNop43EIyhEH4D2ygz5q9
FlfnCg8YkvZpwGR0WN0RU0zrKH5pprSNkPZs4diJBKJ1nHE5MKGhk2Vw1pRB92ID
VIgUogUR74umD/8QTLucm3mZN2l+XVdrKCW+7TJnC9h3RiDKSdA7wbAthHHq4iG8
/CsI2sq3uIL9v3j+egI5oRq4KQ5yZv3CjWA2SFnhNfGaiF+l7luu7zf3nhkDrXWJ
z3hcjyT8sgOAO1f1SmY7LbefOm9+0leO+YgjUdK8Be/IbL0yRp4A9fIQR9WbLvM7
xqxmHex0tav9gXnuB7WXEk4oJZt4n7FAE/RIBrZYpMWoslDBQrc6u/2Vw38jT6UD
z3MoYK0Ggik8IhFdwfibCooVhnoS8ndDgEv2FCAOLnxwnyDG9zh7FdW6+ldZVqK/
5E324gnAyEjZbNlSLqFYc30W8jGdFaJJlZrVItUOi4cTQ+G6tk6Jodqtne2wdegR
pDnq7xru27DCMc7HxfzXNei3m+jBcMd4vvWZpL6I8Gu4dMdLC68mJZzUQzM97Ypi
E4vENcpyoIK/onVzEKMo4uau71IrIuip7+byKzgU2hQSuHX/+q32V3VON4+exODU
yD3N0p6eX5be8Ts38HELxi+kmMcqZ6BJk0mCaS0Y0zzOyY18r3wxZNzJq0Oy1zJv
oF52ahNHKH2s53nvOBVAy793jFMPRDlOwEEKq0sMdA3awwTBsejg4oKbvGGBpxu5
JychzBxDHHkgOgcjP81GbubTrsJTPsF6IAhxe1Bjid+kQU1PuWnMqV0LS5FV69Ja
NSV9HAo0kKZvdQXT7Cm2xfGSuqLjsnK9oB3/rdE61UDdy9RoIbw26hI+otacpPmp
WWjDbOr8AnWjSgDJaAm46Lh870p3lYDQoHdA58OuyvYDFfXbSVrKUSH1OSDheQGB
zEfxITcdjoEnEALbz4KzUZTUfcqAaTFtaTd44U3D1r10mbb8l4FBWIXmv6vkoOFU
jY5wCbkJB9OPbBEM+03w+8ILXNqQ5YzNyBaDv/Yavtpf7FxvU4+aRezVG9oCSauZ
VxQtkFCmPxPixGSwbQwY6bzh24XvHDJS9vBldBsERPv0LXWNKlik9SupX7uKjh6Q
hevLFObfqUeVKs4uqQoXV1YxdyWphyWAmGBqH4TIuUDloh7SzpQcDiYzrIyELxH4
tYLS0QBfXH/EKSPrR3DfPTpxRkI1wlhugHHx7IO/L68Jq4G8RGUR0nB2XDHIHmGf
Y0xXw4QQfAOLOsuAIoKaZiB8d4dCrSEpIeSpTBgYw32VTotUc2V6+xOBH0WFGfys
bQVj4OzNcW3MvDReSIRxt1S566JfcE1sYhr2khklcdz7LSjYSxoCoXAtOXzIiQUF
yj5XJWQCBlSILaN/2nh/HgESfIGhK8yH+HnM26t6D3EhCDbbdyAqeuFJsOHgAjjq
EyYUxM6eqlY4BqSaXxvliQPpkQd05EEUQHGWYG86zD8rDcqWJn0D0/zyCONKfOq4
fbV6FZJkKnxN7Ym6B/d2QSCUTQX3JJi3pESG+wE02yKcCNzbrN3S3RZyFYA9ZzrQ
JyQAj2i4YMPFATRyHCD/ClFx+4hJpteaiTYL0odbuUOsegUa+pa4+lsXRlLzrDvB
QHcldp3hq7GPS/2V45z9vaLWfxWj0KSHVX9aD5vCPe8tmB1XwukqvI3Itu2kYP02
9Zlv/vE8V2ijUGKFiWE7RMSp6D0vbH2+rr7wiMQZaC/1pFAlrngTBQuHhX6EwvVU
qxfTcfFSyP562tYTC7dMDzr8HaF+ozexTdumvXQlzAsZlQxrG6lB3M0COigiP0N9
Ej4lmd/atxHSyJFJf4q4whyEMRRm03vB/qSgOlL9FArsH8AYkdlxUM5U+HwxHZvb
3CDT/n7CIuYtzMm2efIPedQ9+lEQvqOMX8rVmxRZjPX8OkpldEgyvA6RgPMJN9w8
Yp/0jWALwfn9zCCXTvZnphkqmoNDL3V1zF3ZIK8nbUVur9b9W1I8sV9Ey+QcXZ1y
8FKUPnRblGN3GsN9gL7AAOw3R5psT6e4yniacrJ/6M1oKrUa5DjQUoOGVWJMmCJV
8xTnjZyGCo3rOZaNfnmCojW1flvmOZRkSjTF151qrFuYDqapKmO6o0XKEtNVf4EM
5h0vT6Cfb3/qDbui7Pb5VdW54VWcSsMG5j3BrrNHzEoK9gCQICyj9GP2ZvLhCyfD
qo3MBlHio7xI0H1MBPPm7hKZv7wChDnrIexnaSP7vKY4JIni724ysJJaWVjpaX4N
bjcY4bPahK0Hb4Encs3Urw8QcXbhKsgNzuI/i/k9kCT7WiNLPKKuPCHOxAunvSuy
2eyDgvJjGyKD+a7M2AsbBOuWhEhZSr4Q475UMUL+Ev7KiRfWr4CfHDAal7EWr+Lf
byenTtl9tiaPQEbvxoFIaRL584XGQSQMnTzKLT8+y4Vf8LU4l0GTxsPenxDNo0c+
tPiqcB9usxi/0MalFdpl9k83jcM3eVzBi7LzApdcKpkioBTpuE1LBv+yW8KhzdwH
AMLFD9wUeh9NE9JC10xy5NCTfddgkxohw4gd0u3nvjU64FB0DRAas0UYRmr66cwf
wD5Rv81vDkYoSCIm52DAb3xyWqVIyzrB2tScqzIQyWhOViTC8YU7y9PexzCPx+72
GO9JbDFIs3Pg+EltS1TDrlQ6q1xZBGs96RdJh5W7vof6Gavpb/A2AvdJSUVmoCIL
v1oaVtqXHjZ4dW0w6E593BiVjkg+0IakMPQoTYTbxgAQtXqx2BVj0MPu4X7UIbgq
3RCva8NIPbflxc/S3b7EPX3DbPcma4fHhTavQEpTotxP5p/55GpRl0E9F+efeyVR
NUQpk/RdUH3mzz0cjK6mF13e7PXh0Vc9bid6XQ3tXxKDnrVAE9wBChwY/i2nMqlW
KGFBB4id17jA08akFTQORON/YXyEBkb90vWN5eaKbsM6TzEtq1tvTR9Qb2dkDr2P
zVrg+HtENnZ8xHYFpnFlJEjgdOSTHMqYrHYcqZ3kVqRcuUYYESDqokZPIqyrHX4l
it/2PZHq23/kl98yA7eJzSU80sfvTvQHb3XnFm9mVZz+CyGD34cpHNSI6Fq8DViV
YDagmBy0lzrdrNu7XozlZLJQxKWK9D0k3EA1IMaP2iEg6Rfk6FWuj7OS/8tjMjr+
Gxa7AAYkaYKXFiv5mRf4Jy4z/H0C9VAFIWM3o205ih4LYGccJ7ILKHW8rE9XZoMQ
404USW7fnJ+/9NE1L/Nfkvx6ZTf8e9FoX45Kaae+GNyBG0/LBTAL+DCSf71D7aSY
E0SGtk3H5ZT9Hv90phPCnzwxjlgcrqWUETCmaETdTmb83xVUMHXlp43JLoJPSAK5
oxxiU85WvrHJ64FKrijM2ntl2re64KPhoESAhXUscJ7yUUqQw9rVc3WKKDpN1NRA
0wrMaDwBNg+Uew+WMeSQO/yDRP457jJZXkk3538ymTDIHmoYe/Pm12qKyh9boufY
45rzhuUt1wFPgCLg7cCSFRLuzXDeLPrCC4FpIELsb4P9uOdyzzOgjr93xM+19ZTu
r03AOs5HbFfGX1zM28JdWe1qiSwWPxpHciFX3OZtpNWlrMUYRifoM51C4m1KlFNg
vUCBqRJia+fo12fRqXs+/taKEA0aBbwl9iLw7F2e24Ulb39wc2bTC49KU/eyFtxz
NWTQMsP2fszESoueICkxFeliouuNJitMtVZhTvBz9c2v1OQCYmFD9HjVUIPikpmf
1AcHX55vb3UcViVHB30B29g6mhQXJZNLRzPv99h/mCY6XqFgbZ14uEg6MbGcXPQz
V2k44cUcSVAX65TnTV0IfL2MKMuruxBDSCWyD2vPU+4yC9x7FlQuHWKmDfXvtw5v
945Z6IAIbTKpjaugfmigm7r0KXV4vpMYwqnbFe6Y1uAiOUHKa8z/m4Vo6c5En8iB
fy9TWnyifyyeXgpX2CC6i8/ccgksiDQkUFwfseyGJT5yiRhZVUjVutlYFwS3Q8ex
XNlpQjZAOSTqscSWELGqSc17IhR/IqTAmU3FN7nWjtSN9K24LP20PY84+Uye36Wx
I2U46EN/44uSUHizDZAvsKl+4sRAdovzqpA/FrRQl6UMzpXznDpcPxluWjhubG4C
m4X9nxGMXMUGj/P25kSbagQGYifEaYb1oxhEBqax/7TEISkaMx8uy2fu4VK5gyyW
mtB05XqWgfsazkm9ttQK2cJZWWqVVS4sZeuQZO1p57D5dtuF2PFz/yKG5k32fXOe
M3zGfaU0iUjTJRnXk5JaE9CRvUtRh119aFqCfuLeKoV9Gn8tufzS9gPOfW2PM7FW
3II68DTGFZ3R37KVxAYoxPxIA9PwnJFt2Xs9kBAnV9m+UAidJI1yiyL1j+5ID77l
QCFT8xrVUhIKM6RQbMI2DQeA2HaGvx92kMZJG2HBdurdASCGZz9GKoyWkEOMiROx
SPYBxTW2TlH8AdkQE7UolKrTEl0JsxaE5/qpJZeHTAGdKBLQJsPCKd8g5gRywtHs
S+2RZ59zUoe0M7CSGediNp3htyJK1dsSIhM1ZB/lOi11V8N3zUmRm4O8//oE8DLp
B6EbihmZipk/AygsPE+Gs0Vsjxh6cb+JHme1TvJ1ecHT6E4IwP0Dxnei6tw6HV9n
dJTaHoUMYZPdLeasjZpczZ+lakNzNgBNr0Xuii2peJxFQUoR+KzoPfgcroMfbpKA
CPgFbvcpqak1GzJQPNkVq41vzd5OoUGfQz85CPX0VlI5Rt9HcizIax41Scq1yhBp
4hb2aGHTssEZXhQrFZA1t38hjaCHF49/bGgcINm16MKJ/7+SQeEi5Qb13onwgjCf
BnWxxajltxrCcLZWIwj47SWaH93PKRRcIrvxDDwhwExUvpeJO0bTuPWa/BIyYBGl
ngK57tOarwy4XG2PARRSyYTfiVO0bb9lbekdwNgNrmB1GgCdTAizDPNrTF40ztj5
I5ss9qYjnKzTfJVkYJYJzklicrKlBIdpV7KbSmlX8hC/ZDh3Z2WGU3Dw0gP+iuXL
6orNsXKVODU/O+sCJZmGKKXv2s/6YTydrtDQ8pI09MaxmiuayY4p6hpd2yaBC5XY
BENqQ64iUnauOGSAwm5j49XdUdWJcwgr9tufI12n4cQCFORoEYoLnId5QOnnXuB1
BS3n6wFCOvV4tKglBMibS/bdqXh2mqHxIMAlBhxWq7aBQvxrEtyO6/2Kb2SkniE1
+8okWaU/m8JjsOOc7rxj/SEKuma/jKv3f+XP4Lo9yovPnnvCkcYPDUKYy4VbV27b
WH8nbA+b9qzCThaqjF2TT5YFJIjat2dQG3PwgXEpceYO+fWuR6vZ7XC9U3KwfzvN
bvam+0Y4d6LLbsKmO0zi3ifFhslXDKGSo1Hp9Od9QU5vRf8Ujy97Evdvmdi5cONq
FJrI8YMFjia40tzI4JVj7fGZktqPdsnG6yP6gGDzV67jg69sUcpRRR2G60G5gCVD
iBHEyCPlEtRLREtEBaAKipnOCS2H7xqq5ZAjJPhK46lykj5H4YZ0G5t9BPKKXvoS
Y63EoKFlPx+GjIq0c3selHTrW0yZHbak6R9I2u/EhwrpZZ5HNIGoSTyYs5KIBw5l
zCis90v3eKuwhMzIb5B82FlqWgQp1kfeh1rZrir8S2O0EqM9kV45LOzgDAhxZAfC
mDazHrMNb1efP7hN3ZzrwoBsW0ayPBU80cHZH73GhfbMXeGN26C3DfFLBWzmY/sy
UqSknLN1ItnGlAscLpZwP/dXbCdYNMFhNsau4ELoStfrx9THEz+Ni/1BGQrJ8gN6
BPGgz8CeBgoNYryOMIZ0GeO4q40c9PH5nQ33umoGbg34sMJCQi3W6XO4uYe7tIdH
SDvev4MCyYjFupkUkQ3jzsvJAnT0O0B21bnXdA5xmOgzdBAqrKWn8zZnNHhgC77c
u55DAVS7FRIA/EidD7udroEPn7OunI2DdTilaDvIEgsCHQ/lClAWbcFRMcnWag5h
9Aby0FRsnOag0ALqLUOguWClVN+9jElFaSYChMn7Jh2DzROJntwLkB5ilhB5DXpA
0vHmqb+pDCazQiIeFU9HtGRG19Kinh9mYuziLFl2IQTdMr+FkgR2ELa1ZbsrzNxC
pTWOZBcke74pkrUYh/GbmPX5Xnp6SlGmBn1h5vMROG3yj+cXc75KYWJh6w6tk3q+
yPQNiqJ98fN7eqY2bk6ouZlsW+hh8mJuULnLjBvJupj+puudawAD2m0UR/Oy5iDU
493h7seQ4B+fXOoh9bc55yA9azHnBITElapNmCWFg+c8KvGDaD5TSAWHhuG/u5ns
Nf1s0JmvXyu/veIpu3zoKEYjrGQQvhfE/O79LLRK0sFg4V4B0mzyArdUJAb8d0Tt
WzWsTpSrHoes+NXFVfz1vOcfP/MVjdN/sZjbc+kk1oIB5/NmYxEyD0Kh9AFZaPu6
y6mXyvmKAxuHT8yauzFCr8ff3FGOo3wNVROU9n8TaQMhX2sDR3Zl9PEqYBa6SVt3
9mcCV94Hs4kyttxddOQXXUR/Ytzah/nEzQ/ALQAsnMtpot3BbOMIunilf7bwDb7t
bmTw1PkPlHF2+tEwlrUl+46d+07a79XGJHUTukCjAd4fY7dAlTY8PM3cOGpRt8vf
0P07EbmqVqMI2UpCllkOqZ4dQcCkdHHYezZIKtN8lbiwhvt/qBGRv3P9NZ9yY/pS
12Pzq+6dqGKAxY3/wyAKgMmlahfT4W4VK+ugIdFkrOyvCVxYpkLUIc1ucIGo0FwH
ygHWp7h9DPgI1+bLWT8iIIadIcr/Vvnq09JDL2n+oNBNFgz0otOou9EROk6UswWG
nfeYn4cmll60cLgchiw/cJ/jjmL/IIsVzUYwTX+tP5JboJaVXOIogQBm1PPFb/bv
m/SpP19xdV5C3X7bmwevq1iA7rqa5G5+YVF5qyrzJ/WOBI6vC5CrNthmTQqVlSXT
/hijglbRFIheRy/M8GCAUarzkIhfJI0SLa+cMR9XwyRL6qT4fL5lznJEf8IAfebX
bnOo/03+9w0Iug9/bVWudIEbSOKYH6xSo21KyU9NI1iDM+3iqBG8Zmje5n+GFkZR
f80q8qUPXBs0caMq9emkGJijKa3rUi12IEmoBcNC4IN99nlwDcCfLM32Q2pBHU5p
FnLBmvug8/fPDM9+Bw4fbtCvNiFJkOFLiiA/Tmrv/esqmxxOq04/G6o4OueL1CLf
zgKsuN6lJBNtaxZlgRCzAt1Gdbrluzhlhoh77bXbZGVmpQ1lnDriG+/CwCzbz3nv
hLaKjAtyriRHpkEOZpIucklcRNYixlp4gasCy7os3FL3pvb04ZTFX9cix+ybjKRL
gokIlhlJoEN4qPo49YMKSZDQXmoSCxoWDoz1i0TwfN7JDiyJapqMMPe4BHUiW4NO
qY+XWySoP+WoNiR31ThtMf7g+rGo0Xrw+NjrqG6R4TRKtFt1qRRsl60heuArG6MU
+I2X2XEShXKKCymUfsQtSOQYdzlV1j2J1AaSqvdE9sF5Khkw3U7vEQv1ovv6bBkc
JgIeopDM9OVmuq3Es8tnp1EimNr7Ie6VCF/irnyefVRkPVpgH8Wuy8XyKheICdqr
FgfaTRNd/cdUTzb/tP9AjjassKrcpabrXh+mLHYErOH9p3q8HIcQ/caWKai5kpVO
eiytYa3V0rlyDGcq3MRwhKp80OBIkw7xi0/Sx/Ok4qi1m1P9YUplp2CENm6x/XJG
cdp61cpUVIzV2v6L8xaq+nPLbhf1HSNnfrLQJJMKwtUrPvqhLz3gyc8+JEFRlSMk
lrrUstr71b3nkRz6hCup/NeNp8+fFSwan7Dx7iWAlbKLGsCKBBl9Scq12SKzVee6
PZTXtvhDN8teJp1Mv2g5PuId9XqEZk7hdN6Zbsfw3rh4LATENdTTAUgLoqmu+INE
qQcoTDwDdCAJWQFtEi3XxX4dju7b6iGbcEADnZOEiW3tA1skK/ulmdFVZU64WH1O
F+/lWKRx3BOgS2tS1LHylj7Kalcguus2fB93XSgct+SuqJwjY+sokXVrnYPWOCso
QGVq0GEziv9Ne9LuIqFUvc2rujfQp/cUp2hVeRIqWPK1JJ/9jFBd8WgXEt08KAOt
1Z5u1Hoxv9gqt/bGwjoIj9HsHHDVYlqZTuIAlDjGWQgOLsJLXtUmV9nHnqXA/nXW
oJGHVKRQb4clJb7YeCZmnL9099VvllmLfN0KoG+CTrT3037/boMD2bilT6L77NRL
GJ6hvvA2nVbFDqsbi0pMMrsWUqjK3c/DsHtKe6uK7OrywX5bTbX9dH5rkRP8oavU
tnwkdlfhADjUAQinJOSJRAxlMRCimRHM9+sYI5taSXkQhN30lJwj4M8mi3VDxYyn
cGaZWnVE3iFaax0hupMiGC1lCuQ5PZcXxfpwYE3Nagu6fv6Gb9iyzhuBprIAztxB
O7BpNkiEIWZktY13xA5CymEi2O44T275yhUYm/cpsOFT6ZEQAs8Y2Y6YKwcfJ9Qe
vtIT/ArKPTNEV/rrO/Glb36xFppi0pGQlUGcfb8jQ9KYQoFcxwCNHoeWB2Ek0KOl
Nmub8tIzPs4wPi/AU59w5iw/vvtQ5dNdFJPY1jV/pSS8nBy8GF+CDada6Y2JBamo
hXhkahlBz3fITu3c1gFMDz4nrfTXTcmZpdScNo9nizjQeLZzmAFlYbJoN8ZAphwr
rj0ecr55ZnFCdjrJrpWvYqbX8yiXN+L0O9b6cCEJGdHUhoBWFgLJ0FuVdEGgkpfT
24ub1VWPaCn6New8aGE+GR3QH2cDQmoqpehk5Igipeyr6r9CNL8HOjoG6QJuLO2+
kkGrGwHvP8gGB3PZDaZIUZ/Ts3VAc718Tuy1iXkXS4XLhvxEJIaNYQXNyByfqNbg
PLOaxwUbpjk1sQFM7+D5hPLoz37G1Wg6aFVPry2kMhjPB0V1bDr/oK5tcSIUN7La
3Z5ayJId0ky6wh+I2aRDC0QG7W5O8jsQHHJy5/QVB1UE3MUXB0Utv2SN59F6/AUC
iJYrZuktbJMloIbS0d6yRXXby4WWR2ssGhQ6A425QP5Mn3UvDw1oh7q8n6Zw/bUI
WVrvI2k+w9PuNXrUe0hmqX1+ER0I3W761yUkEAlWJl78eE1HVsP81ghXYYZ76Fun
/WTmJFs8THW0mdAFUhxcGi1Uwyb8hF0yjnzB9LpUvH0o/ChR5Ty9g+ezlRbDmP5q
1VrLgOpm8a9iEXC6+ed63bLPjpnudsa3Uxv8VDSYybJI1conceQx/5KrUxj3FSjm
kYIQ2uB8LW2fEelqggigZ9z5OPKGRML2JWSgWao0V2iUpQ5R8TSxjBABCbbH4A0f
DzD0q0JzMxZ0qQgU5V73rRXLsGCHbgLdSwb69rr9DOO9+PM/0rGczXfwPq68ihkJ
CLTEhOE+ItjFOf6FaO95ODvEc8zM/6qsk+fMQgdbX278zTtKdhzjy2uz8er8Sy1a
w2c32RZAozQXrDkwTrC6Dl1/XCmK1z+bgk98DYjdexRddjLPizFZlX9aL6ktCfd2
CdXh2YgRYc6+wXZ4LPqWsyC/F6hpxiVJgxaOKXWIttT4Av8DMQLV2ONx1wNy/oHV
+pR+Z8WGjlV+VCYrFbXWlMUCALLqeAWj1lTNxzmQLhJEso7VsYYHAIU86O2e7QmK
1I+09Dup8p2JaL5Dd7DGYZayKMbHmY3AVqZ/sPgLfgr5zI7mO9dDC1PmuBs1cz9n
k7xnEtVKEtZ6tj6c9tnMJjXRROmpJIHDSMWFwJxNu4HLWFLAUrhsEbqmH4gelNV9
8+tuKrMykqKX5PMpoyY0Yb7pR46ESqtLl6u9pWu3P+sPqB8rcLEh10nZne7EwF4w
YTcukNyAYI2P7wmORjE35/+X6mL30xuHUQbwb59jhewImVUpRCRGQIKQH6WX+t5v
YKNhdE7AAmqUqoU/5z9lp9Hwf0NhAcfjYCcgHZS1vW9b4L0paSgkk+SDVelD68eC
2q+XCKZ/FS/PIMzkCJdVlBy9+smUnnPTJb3fFKhjiLOH2T+mGOPv28bwcfTLaGBo
tjIxgUe5mh5tE3eUP/5mSHdkG0x9WQjDE+ZsycteBOOdc97EeneJpd+JaOfJ2Tdk
VylkuTcT+aBgU27wpKZsi3ZPxHtQ/qhYxf0QgmEB0iOL0jUGTdJhB8L1p59no6Mk
cufgHD8a5G1q0vqCNrgd2VbeAD4s5JYqUYy3E1S7PP4c0op5t6ksg2c9+KOEjN4P
idOFwNFbwicRvLfXfxB8ppovkSjUjbxtX5F1WVzufvg5m0VpNqSoEIF2nm2STcj3
VlvdExys4xr/nvc1kRdzm+u+cJncRJ9GxlF39r4xrHxLqEchdN3OqnonIOfXjJY0
/tF3mO6+YmXDUMiKWueprOMqrNn4tMh28uKeLd2P/eR/3adHQR6uupvSAh0oQhTq
OdCgtPiJbvc3B1vz/xbG2U6Kttjnez2O8r62Uo7J9KACbNy/Lw+PErTCoOciqYSr
apuP4QYtPc1AVfUiBqzkPVjTNnFPM0GQZSNOsBPXuZf8NXp1j7PL0AaQGmZmzqb+
6vcPsIPA3Z54/+XAUsDWAW6HEC+SnsdqwAyNqZy7aGYoanIExc/jz7QSBlixw8+l
u1i0Zpm2fke8RXaPLY823xDg3WnsthCosJS4QBxAoYrpB1bOOzBD96RAPvACTeVD
2OCeqyuhu2AgVWuMu31QBvzLm1UWe/iiIhb+ie/r/t5m2SIOSvjVHTPLz4UbJc6y
KSa9bDdAi9U26OjpQgozwek0GpYsWpBE8oJKu9x500/HAdvJuuMGpwCSPwXuSebA
TPDZZ9G/+MwtjQo3LDYv2byg1FeiQx7Z9LpjTsbg0tJrGOQeg1ccMzwSyshVRBRd
bf1wvhbiicYlXRa64/T+Wo/8c8A2ZtFwOHvcP2PuLaIY3ll02EbengyPIenOMdRt
uVRAR8Y815ig/StUq80+gI2Jg0LNn3+Z2brEwVTfwxMhKm1EuGHJSJRGFFLAwYHP
vf31BuSECZ4xxOMXDUPsbbObNIKe2iiMYNkNw8gIO96nGN4RyqahYs21vT02xHD6
Zp7U+LH6PAeuyGDLYim0Ez2VKJfdSn0PMn5O+3EPAXXUB4PbKIU7D2iTYjnMnhMG
ilyp9lDUJJ72LbBVOb4V14etro4/On8lRmqoa81oTcK5xkIhixSbHUgyzQH22XaF
Hf6+vsOav2KgSM9ocEgH1cYzfjFkUDHb0ogPrkt6CTNvSiyd0Kqde3T3wh/m8Nda
gcy1Yvx97YjPOC5vvKDMXVi4teSp032/O30AWSafV57YZykiImUs9qWS0c3+QgGk
g12efLx7jG288lbNWAJ02ZgPR/QUasWgGimuqK+z9iIzv331sYRYve0VbHOqHlEu
ufOmJmIw5ypDUdvT22eTbf45CYXITjuLBFOYHNbh7wiKuLMjD/+VL3Gk4zsHhuZr
FjUTlz5IUo59uHVcZrgy+pG5ZQXkF9KHx4azzuNqhbLN1gHoIwpyhPO9j5bJuIUC
Xsrpam9KoJtw/zgMfZhjj5SZNCvsSisYLjEYErfXr+cq+i/PKXhgWhCt1JM/BzVn
s0SVJPNzQsgIJ7ZG8rpjFWcpoP+PELAchXQ/lIbz2VGHURwR2PisgSihhwXJhbn6
cd72jCvj78fOHDWDwQLHs40keOwKcQNjjrYfcbE8Sg/0/xpBEdPMNZ4HLBT2FniT
NRg2Cfmp1JvLHKWCwk7Vm3VFLJqXLYY+B9hUCiP68TODRyraLSAa4dEX/m1dzAY5
1PixUQSuXnt+oA+/3a95aQLEV/rjmHxt4/Km0KEQSRaKFnVLu1AMbKA0RKcKA4F8
+dJ61vbC/n0HoUkR07zJM8eiDfp4djjI1LgWwcI9Ckp5G7qtD08QmJi1uwyOq9ka
4yv8w6pytz8+y4x0FB7RfASso+z9HlrVHwFb3DrPvv6Q7RGYxcsMZjYrYcGbjA5b
B93Sm12JT8W6YFWbdhEsfiadSr1gg9QHouHUkdTqoRdHZhF37Ml1+hcuRjpc4ttR
v6KYqAeMH6FPmJ1FKWVv3PK0Upuy5E6qggY6bHNNqlVsXJSmOgDlgybjQhLBdOPQ
zlSxUYa2hQ3dPm9yjvEMWNtGgIyRVPD0a+c5erfK7jJ7l3V7EcaTu5tyMqi6TmJl
7Ev/TT4a1lL/IX9tqhvjP7+1ymdr5m/PdHWR/kq58jlC1czJXymWO15bzH7X5d1d
8pCHSxD2P7YJyEqS6tYNYKlxxe0JVk+dX3kCQup3PGGQ9JBjdQU6SrAsOuFj8y61
P3iliX/wzaPRs04dPfRS6BIKwKRFVBVds1khEHjroLo1llZlvDTAIyEnJL4hnjIn
LLi/Jw0c7046kwY159ZDz9aAk5H/2zCi9vwAmmbRYHLvPg8j9MlokQ4lRQZ70eGF
Eqkb8uA3u9MAlCPG7W2iYSHj8nsirMZ1wUX9TdgEFsybTTPBUzleIY6Zc+t9yK29
GNjU+fjeBv5CSVfd5narhMixN1LMm3egq3egQgBZ0PGZLvzMrhPjP5Ev3l9K45b0
WEd6GErPqIAaLFxlWTT042GQucg2z3OzzQKo1zne3u0jTgV8ku9g8h8RutIhem58
nwHQCKJ/h7jgyn/P2hDrVaJ2TIuRhsbS2eZwToW8dPMxtWIzb2ilEiDdlY7BQ/PB
3p/JjfVCeO55NcOQoLV5HIAoJq8fseKpc3p7Hsdjtbc6vzaTw7+ijaMegijFFGG5
E3PFnlXjBnBFHrPP+uP+BO3Bxd+TvxD8b3AmWvDvbL0emLRpvCzP3La9sBk3re1X
ofg/eS7R4PVhlM3y+0vkY03VK/7FiroIdkPWOSpxGj5DNRQT3FGRbj+G5A2cIL/N
nwXRow3PItOlCz8TFJ+3lIC3v7x4/TbByZOiZPsU8QHP1trAHy+VnY2CLvoFOJMp
Uwpwo5Wk7UmWHBuyQIp5vZ4hoi/tNHcrF6UMplGurH4RZuYjRGDJlN2CBYk8UPU6
00eAq3jJaLnBCXy3xoH4sHUueCqnh/e0PoPlNrJ6fpu1B+i7xAh/XaxNmoGwPwqY
oi7TozW/iYbtvG0L2YYfXkqI8+UDsg7ULE8BB2H+V8I0jeUI3tmh4pTJgeNN0tMm
/Fd1han7hU6YDXNqtcw72wXSmX+HLkLxMTxs05Gu3u7M0LBQxFfzrd4UIJq75/vN
dayBqNcHbtfkxVHqx7A9F2nwKlcemUnN2ID/qsqorxKaOXNreLMw5CaN15FXBjK+
MNgxwCWvFFKyD2PQUQCJJYhoID4hUdmtGS/fjuWvB5qGeZIzPmPhaNbKxxvyMFyX
ZVHD83Cnhga3p3XVS/AuIrD05IXxHL/QjkDLUj6UiDOyiO+S46wSkXuRP54QQ7+W
VM+x262jhR3Q79yJI82VCXcvU0M517G4ekQMIsmHvEMoeajLUyBafjTHRCFoOMG8
oWoJE1IznHcPUSI1yhLVoAh3PDj2a9zK+3zj7JcNBqO8Cltb8f47GtaQ/iN61AD4
QxWpImYqaZIfEY/jlXaQFq2TUPC9gXkn4AoBb6MBbQyaGa6cjdkBy6UfP9kz3iqy
I6DsS6BmyIWnlxdnGEk6KQqZB8GMrE2PG3d4QBtGzHNDoJ85erkgsBRuq5oHvXlF
Zctgtw14abKTjEEp+8fA+HYbBTMAW+prJnWxBT8keNKTydQH8hxzoq7eekRTobPe
c89VOYSfZoqBksSkFOOIi5qLUEUczGBCI9EVIHW4/kfvrmmNtkid17yirI1jTwYA
PVCAuAZEgRWU5J25sgPSe//dhnWrCLCuW7wQ1j+QDUqG0ICVI1zHKERorxuNhLTK
xA4qSqu+cEmUOALkv4KrPCWEuksG0DSwkQSR5tjjjT2ECo2k1n8wf/YyUSwIbfZU
LQITeNzHofdQkCyghgzdGxf6pM2Q8xkHyZje8BCJqGZcsxjtSoxK9aQI0FTMX36I
M+wZ9Q14Vef9wqmCwgXfGG2/6P0rfHGIMqgvx8pNHxknmxPa720i4W/B7fs2//AK
J/+QOEkcQQ7ZtrvKH3L0KY7O0HX4k1/glQQxnqI7ougU4X3eOlFxqK6Fy5KU2u+U
DxYkyEVkGShKw+Sx2v50NCnwhF4q6LTBP/mS34kJUNfan/3D7mlc1YjKv6ki+Ty1
u5Och1u+nSeb9wYDz+yYT+hwZmCRwz29KvA84/M2zMZu8lCPF7XLWgNaj2ovSgHb
ubCUYVGMSEAzUqZQC5h5FsSwkg6bhIuoRWq/8wL1dwgn/rqCj8Plv0wE+l1GP15S
AKSU+amDhIgLxPWZJxzCcSt9eWAwmff6vTDhzTClVUZvh+abcgw2Lta6KS/pg3tl
qWTKhNiustPkn1wjrIozQlYRfAD5Lonq48W+oxI0aM4nsqHKQscNzfeDdXEkaAI6
QbOPyYJ9BKviug4QxL+Pz5IgXxn9qWFvVvBXtjXRoEBIX5OrzsFWCQiRdwdEU0bo
sKJ8gDJzdeOwqezIvZ9sGo5eMFJ8XXZLYcwcNVZAX7IIujUohSS+xxiUnfgDzRNN
807lu85MZVsIhgBZUC9rtMWNIks3MbMF3N+KGpknUOzrupnBPROztJjfIGLs5l5w
6AsW12XTrFh/yViPIEczsgGnyzjCtXvxuvHDLt1GabBSh72Mrz8PAUyEnXP/6c72
AyxAdsfqhRufzG4S8zhaSWGGyRHDA7oCNwl8BHoI6wyDlswh4QfnTyxBO+KPedP8
OLRFxFgnYEyrh3eUtGog/KrgRWip8UliUuG10HhTntu902h23ooOYrrVtgIfckDU
H49jWZfSCw9kxf+x+3o4cnG9yXs+fUDbF94OubskYqt/q2GQoyBCIH3JVyawS1Tm
cSWaXhJlWHtN3UOh5jXjCjHuHUnUz3hyDYneRZ/rubumk7QL/0nrMXCkB0XBFVHw
xh6iRtV9FCFNwZL37nhbJiX1bN01UjBkrlOGAoaFbWCehIGs1uMvBcIlFlii4P1e
TBLyklS8sS7mOv06TrMjJUzHgBwm1sUsJrFpZJ0o1OGPH/tmXXkPJ/BkbTmfSKRj
9b7Fakyr1jfG1OGpaOK6IeBSJykg8NrBmQT0iY0cDdudHkmhJhNajZ1LFBzTly13
EQag225OgmyFsznFQXu/HD9TnBOUhih9aKjytaemmL5D9AsEM/CA5G6BhdaMfmKz
taV5xCpcL9poItrPQLPoL76pMB+b9597U5vpct2Vp5wHhIVI1/iJY3mNBwkj9vGx
giZEapToqJFPtcWFxinWlUA+3A8HB5Iqr5ygKAzij++H/HgHc3OND3qZfSScnfBt
mylxRbWnJuPSK6nZ+tLBDpr6M7XJpnMOCKdaWwnR2uIyxjFgz1tZ2mmjWeiJ3Lrz
D10EXdqTA94hkfjDZ1z100VBa6Ssf7BUIsRiBSYwsAl/xHYBD5O40lWPWV/WCK4/
qumPzqJADFaa69uZynpCANUZzsGGc81AY9sJL/bGU9RvAS+Alhy4LiNrKtKCOcWm
2WkVUCbqyMgXIyNSwYAMUpg5fshgNOPbEplMOH2vcIPEy6EqP5bWsG2U4t4tsOXM
ADN6ynMD+s0O/MNRnjA09CxSYiAw5F2E8gpdGLPP+UKTZ+24YGKTlXkLjKe9MnAS
VRcCIXgK/QUai+bwehY76MxXzr5THZPRk27R0CUYnRjhRqjdqxBVa8Ej2SYgm9Nm
1tiLov/tb4sQ+hQtjElzZW4q2yVDgxqyS0LV2ut80MfpVnHDk2fva8c0ie1oRVv8
OybhXYAn4UStCLWBszNPU2cCZkQGLqmX1bxSdOeUNzpl2zLVXT+fsX1yBxteqwhW
xgJTosoW5sgqVga9OUPZKV+zb1F/VUzj2SsRwj5HiG759TZ0M46RFe5lbY/PFMbN
WdxvoFvwQjc0ruN8ypjdwmYF0WEzrdn460aNmYAJigm+GuMPTYcqi7SSTjJJ8YQB
mUYiSR84pEuJU9ZTEV+mDo5i2Plff9wHcTvA1YTOT8TzjL2p4Nadr0B8gGWVgqGb
YYIzq6ftiPgPPJPmG3g4cQp328SCl00ReNiNqQEDBhhhO8HjK7B8h+4nCtezY93K
xxMxwG0jew/xyLczqmbUbiXQ++S/7xYe558JrdupsrpMJVojA1qSt0MkPCZ+QuHy
kNHMKm7becRwZFendPa0wQMWYBY7tzQl63ak+9Sr826h47zWf3rroK1rfwnTq2AE
/PorNlnR/n16Wd8lrepZZWf0cE5BUoR9Mcm/1+3FRDc533YC2bJ3+V/3s3hKY8Jk
C+q8WTOh3cBlg/KFvMbK4H4o0+lBOkVOGrMVthha5dQzV+6gGYYzc2k2h6/BpZ/w
RWqe/6rfHPas+2OorF+/pqko6K/I18bcUQNRj2K8Meq/dMIfb6b+l5lCw+aTfU5Q
aOkFN4/UmM/I0kebTiBGhHTRENTdbBj1fxOcxRKmrgDceuOkv+vyfJrqMRhkpOhp
wSdMhGNOfXHPYPoA637rtOoK0s2dpG+L1B3hAbwIFvTnStLbj85hY5LpQstq8QDJ
0lgi60yOkUpNT2Y5xqeKwRzQ6peVMkS2pDRDKl5bIQigSPl0rMDgzF1Hb8DlBrzM
IH9QL2Ob7n4DLwl9A2FJwc+rEeI2JzDdUHpk6vJqWYxR6P3XjNvBIxfW49qF3cUv
Ly5NVGGNqUBZfMilkmDTBnJ2QxKQnGpcF61AVrA4FtBfM6TM2IJMC6Ajbi8KqMvW
HRRsEC/Fg//sh6Ejs6GyuW8ChCD9gvDWfsuA3lGkvVdJXI2gKYn9f7LDvIvQdH3F
H6Ll6lpxPVOohUTOKMe3njPjC0N9tPqPGRitJ4MjcoLENFMh7YLCPJm4Yn6lRUw2
Io9inE3HXcGibVj501Cgg/imaCTOfxbLSIRg+ZLvX/WDhVzGViVOQs0wbprVzmFH
jvFSFLCBGe155ijb7YkBAXyqIuRxTJiNZlNDyhvD6sGCTCotY2VHrp59RWo5PvhF
Bx+nwUxcTgAPrl514pKwCKgvmaCchpUcS7PSI0L0gxCcSOeFaGr9ecczTp0+oNGw
1pPzGR5McpB9j1bM506IM3s2P95sX1I4qA3mLIFVBtcmhCxSmUJZDZGBjSwSYi1W
33CSrHAcpuhnjs3+bRJxUgO5+TLtupjDge1iESnZk2XBmbacgZ5Cd9g7Pt59cg8y
UbVLNe+LXLelflnWO8+i33Pc619A1aRcA88b6pyAicpfmpt8K2WmqIPkusH3DfpH
DV/16rwswXkSFPR11OHYVcD+hpdlig4nHKT0RpiEVemAuxf7q5WmdZpS6MH7Ic8B
Np0KTwX3KsAKGmwQvOzz/lME6PuQHZLGAE9IOId0QN94IKyv3W0ZRnwRML4b9kTq
zUsZb+VUKThhMnhKRm9Xq38kdUSFUyRJ1MG5UXBRiEmHbUqYqRx11bxl1nrVJJ1Z
Wf3YUjguAU1FfEgePLj0AxzcA108y/R3lVAjYaOuGvpfLm/kke4KvTn7m/wsfrSS
dZlifx7LSTPdX8LpipADAKaCLcHzG7D/zUtpjPhmq5UMjXK7ItBeshV0UmvKy8dh
i0UBZhXeENHzaFyJ/HfrcDAJAZRgz6zPdVeXLvljg6DQ0GNdZzOMZmufnD4L6RdZ
0Hn45eGvEAENvmBBrOq+nPWKXUNQT8+pA3DgJ2Kjnet3qbPW1UaQrfSqdJ7zoH+Z
LGHFsMWCeDX/q9EH2Jed+wK9OsNWTLWarn+sOfRmza7Rwcm1njhlXDdcnmD5LgDn
wKVrrbZ++HwguRA7kcywyv+1OrmxuWTQjq37HHAmWQoGStWlOm/8hUiIzkQaoAA/
MGg7KeSzJXKm6PdfNm9AjAs8DImOQQZJT7bmmPzsBRUS9nooDNwzp4Mx/NWhE5kA
XjBiOPx28pcjvcNnn6qST4I6f21D3TTa/vdiKVH+ZQtcdh727esuqGdjUwXiziiM
JGGT8rOq/6GnowiGXP0SKSeJjJJVFvJqsTgTtV8r2NM2UK2rhs2J2jp64RDilpUw
/nGigfk/KZeZkPr6KNxxj5hhj169ZGcT/yxs0IgV/dHA2mzZCO5511lelsFfKSCG
gPXZPiHvsAPUJYqM1y9eonfL9OJ+4ovJDVmNOz24PffZl8SLgtELtjR9hi12jSz6
DtTQuzvdsoe/SC6xR7Xm054DoQjmAMgfw6/q0n1/nFsMTeQUVfZartXrsu60AxrB
QNts0hgHGEgOq4KR6ykpJbMbV4l0WKIg9S+t6mdFQyl6xCGVgs7OHxWDzmpdTZzz
KPKnq2flckEmHj7z91Ow/P98zOyv8f/vyhUfYDoJ+ltv4oE8eauDK/0onYWG+J0K
NMvWGPjFdZaPQWokMVsx82+aTU4T2XaAJMW5QnmLmMQWQAWrq/Okl1/6TmtyvBxs
uMXt4peu2xVtRKYyalSGdUtSoKEmZzO+JMI9I0n95Dx09U8amicaDvhk3Oe4VqZE
QN/+NMoAu6KoS6fasOitIcN0xOOpnqEkbTotTjwH58tPlcUpVrNiOpB2QEEX5glH
IeyXUoGdxwsP2HGCIR9iCd+VX9y03Eqplcjxg+jeMfeXSKHrm7FgocduzVDlcmZh
DTHN/AVXzu6Sum3NjdQDR3SQt1+6D7lFBAG5xRWRLTmj1cEtc14maZr5hK7md+h/
8DDDzXrXw2nNQCJc2RkaCJ+erPPQN/INH2mnxzkhTvY908Xlk2rFfldXqUG9kEuY
G1A8TmWVtlZ8+Yt/avexjqY8dO2tUsZSf6XsYqVKq59nnP8PajnYJMYKWtA1TkP3
OZ8UF71yHGPjXdNYBPYZsKk4NsZG+DUXE86GYYRClgo2C3jseLGzS0XFWeTCHQSD
8jadtwf4WIaERIU5pjdiVHqe24kqS/JBN5ngjNg/DZhrpuOwtqo+kuMVDvVfRmMT
NAnaDAlkYyjXMxeUfROKooiAOx3tQGeYVWCHrBixr2E2zqB0WdJWWMuTwK2UUggM
6GL/dtX7MvlFOokzJBHXZ3BfHhJjldoulu5KnZf98toXyUVnoI3WXNu8ksHQZ/JW
bu89K0zsG+vKFdpkFav4ifA+AwwgxqZLYpw9UGUksW5EPCFLATKQ76Q7Yjly1zau
ez1LVYUUhdwr1DQ4GEFTSxVvC5N/Wrsg6QdWj40ud/P+qqzF4z05/KzoEeN9fHkX
tOWMoL8Aijhs84zMOCcxzoms/wvqlcgVTQ1/enHcMMu5NNsCr+utPwV+W+t2n3z+
q1cIQdbw4S6YnSqdgGteoDNg3rv1fr6jqOxC0x4oSLHacvJwbj2VAEzDNEackKbR
tZi/OciAD+e69+Gj3itXDGUJmM4g67LOsgFtOOoJ5ItuaO6RZJjEqD0l31u7watX
5xWF+nGZdeZ37mMfNQb6dDGi0D5sG//gse1hieEibe2KRijbSTAIhvh7z7kPakLa
GeHxrYYNwtbTpwDW/Wpz1OAPzsGOiA6xwDGPgal+mp5JBmlj6VZccezGm/x37N0D
Al/xvuQH3IuGgUf6CSR7Gqd+IFv/Qo9OSYsOwe9WH0sRyR0sCeLqtQI/3qc11B54
l1DWQOU2fMlANoKofz/OqGBdx/sA1rCbhy9EyOtTTCa8osPV6c9R1P4qSmppnE7R
xYp9NslBQmOvdOnw1iaqa8DK0AvCaS9LfMOkrD9MTn+uSdfRvFBxr4i0GMfFuQCq
QReBPSHGCCqzAd+Y+07pC1fuub2fM9zC0Be/cQ9V/i0zNUHHS2Ibf98VBvINGbuZ
Jzoq5I7utZKfceRrKwZTX6ZoXbedcNaMCG1rl4E1j6JoF8Z6DZZbF7cfR3CkD72T
FgQ6PSmunY1HjcZr0iD0+uW3jS2xouxsGd8JpWsL3NFndYD2ltdNxd/OpjwtLzOK
ds63CaXKbcYDX0SiExkcg47yEvKNhYhNvdHYIu1HRZFbII2peVAY9stQJ41YW02c
SydmCKRGOztuh4NGSZ8CXg0nAEsAHA4PDQJX2KqpjzOd5JHb2poOxW3az4+TonMp
e+hzv37QFB3t1/QvZkDhRhO/fC91QPaK5VjBOM3mdrABm/1ZD3CdlkvQ3uXDXKH6
LNPv8V+4gDxv1LBFY8Nkb695nII6xnuHsOZkmWe49IcnU8UeX2EW+jNRxcAr7boT
biHCYMhu4+Y0WFQO6lLzqGxA9jno5GUPhxUjo0IdsHxScXeDVF0l7XFbYvgiBxYI
qGSxht1WlDkGkpMEIFMLFjrws7mMh1UgjH56nBSTQNvd72sU666dD+4seqjPGghz
+FjWtCl8u/D5ZW+CDMKHnnQq71f32L4u7Ju2azV3Rzj2p0LyopQ5e/ARZXvm9U2V
5R29XZ4dRn0Txnw+iRqaRLvg31LaRf/8D6Pts9+yN2uxiXvkCLZB3to5WRH9Dt3L
onT0C3n3eachh9ko+cZXcVtoNIYhZCWYKqwezvWf69gdB90gLiYJ+bxMgvgtrGOm
WlJFW8tIS8ptt6AMypFnntYffWzYa2NnSXa20VxikpRJI4HC+xlqUheJG/mrx1xA
k/xw3JYAks6B3mWKE325XFGNbkIN4bwA7cf/1E4/KGc/oOSwrgjq+KKl+dK36HRe
89t7zMMUCTGzCZz+ZN/URkLoSe8mrRvYfLnGfmjpaB/Np+5E1pPnxIET9sEJ4zhv
1s/8VgIneTmhvA2paYis3igfYoYnYwaJswXwO2PLpuBp+1fz/JB7U2sLIVJpaCDE
Ljle4kXw6isAZIuRqKOucCBy8AiKFjHbF5IpxkWgefv5ZMgg981Zw8v8BAHzD2v6
bUC/sSra+t2+1u48vd1GEijPagv5XOS9oVwuOw4rfBYr7b9nuemnKdouW1BHIUKV
6PN/mxDmdID0j8+Y82lauRVauk3H1EcLBzBP6Tv+KRSDhw4KXCKcWilt+IF/C4uX
8CtmG8hyEJ2D1Pq+UrX3K85Nvwqklaseo8h60lQYpSTqm5Xt+HYZfaAseDGiOxbc
FtMFk7GY2YEsLVNbEt49tiV2HmN7xSSyeSSrsrQN5jjjB8ncd4l1GBp3JduPjnzy
2jyTWD53y0eqOudgbz7aFLsHTGYyHFzgmK4qs3lbKvpH/in+f43xvCLCo0ZqJMB1
gyti3CqXnD8k/uKEZ5TqTIdXYPAqk1mpD9bUY+LFCw3VoCNW5uYdq68flCuaZ/jK
2QJmTYXzxL8pB0FSgWueEIQ3mua97idTAHuccEaAO9eoSWHBzSdi6GKcgD7A92Xg
TTBYFMYUKFEf/ltFAeXw22mu1Yj2BXT/VzU3+5yVMt3a1TufS3aL2HxVREslyJ98
6bbtrnujOWXymUuT9YD4buwKmBiywcmWWkO73mgIv1r+OveO+hEDe0wdPMX/d9qt
5Zo0srrQjBJJ6p6zTaKS66jTNTqURWeIGeG9F3Bwc1NaJC+sOR+D3pMED5fi6nCH
P51ce4wtncL31phRljpwpcO+FQAOXNxCuwLixN8iL3csDaW3VQ7DcGaqKyeMZ82z
Ln0YK6HvQMIUeu+PF0SpEXpP8JaW/G0i9c+U/R6VpND10+JSeGBUBq/i1B+Km+87
Da3y0MNSpyECWUN6t/dsUTAY4uiCPUV7avwrE57SJHjtRmw8v0S2cAPUaWH+oA9Y
8Wr1YCXwLTVtCcJU04yuwT6A5PwD4YCtKhTzig7Wvzx8PYkc1n25XE7ED7H4vA82
68WiUGuGytOGCb3N8Sdx+GE1ngViQiW3eaUy38xOUJS7JnCWIkAcTRF/t8eFhWKK
u11nwLr/A3ZFdE2sGYNQBDJOUki0+v3ndWpj9jnp1TUYCg23ERxnw82eAQqF/CGD
sKlQ/EilyJ2181ltEEUbs/LFvpTtzxDRv7XV8mdg0m5qN/DIalhAPU1GKHdfGzPJ
6I/XVGP/b/McA3j9wX8um8R09cS6lTPDjjI+aTRMsP03GgvVTM6emfq8/Txd5QSn
lLu3c/0KmDAc1LeTYz/nNAPjBbkMSELS4GR776P3NOxogjwN2mBM/JiVRxHU4Cat
o1Z6qNybxWNfPGcDeCjC5OKpfd8ZOcWLLXMF9qyvS6HrmK6+t7TThhsN/UZSLtU9
pNG7UZPva+By81R5ShcXtOXijnOlJjJlUDbOei+FF3F2kdLk+zAV72A4YuAgXiHU
31f8ph9jvS53KrLm9MhwSOl9930GOIEbL4XbwmchMkJHxjpWsLPH9q1E+uWLHxEl
h90MhnseSbvMPeveqiWnWJi0NP3k87fmF+pvapRonWgUPhqWk9XtQnABuUVE0aq+
B6EGB+zekHhkDHRScDAPTsC+pHciF2LhlzITn5bKvrgE1OibiX8fk20IuUUOuaNC
OdkeQdLubh8ZozjImsqOtZzlk5g1l1zB17qG14tM324HUdNKi2tEeVDmBcnuw18r
JlRrt0s6o4owILCQr8fJxh6cP7eyWmr9YJUR63yWgWCz10FTd+hI69lVLkVj6kuI
bbNPbIHhTLDnwBiTB4F+oguqSb7T/o+VhZsgumIPIvGyWkOAECescm4fZouH+zd1
AjAEt5u+dFEAtNdx1vjSuexZuk4NIBQjH5wXH/ljk92oRcsdMxlFDPh3OepEFI7i
Q+64M19Ejs5Rn0Rv9JNkyOF1eikGYoVyojvJKk3FEfvJQ9TKY9YC8ia67xeGALzv
zU+exF7GCQ6t5vUwwuF2GuVyJzUMczu/kMK08GfCbfZyfalRoKc7y7c46gkEH99t
wO7i4t08xjFNpDBLQQH2Z76nMybYH1V16QU3dUGXEY8nsnVJVV0q/FCreKdfbUul
YvFiHPa9motcgoapRSfC8K5vMX619uJ0rCASxasoInVPEmc02lkarHvStRg6sNWb
RlgENPj/BOPi0IX+wUzKuXqIZLXaopAcycfVmAkT2fOsF7CNemQ9PNRJ8HF5hVxO
py7YACMAgISjI2xHY8sEyl70Dg2B06Rk+R9CWgCwuMf4oB4f76ptCKULSkxHdDue
eX8zswH0t5UbxPEsIYVEaq3N+t4AIgXqv08Kj0K263aHonlbEu9Cy2Atbr2Juhgy
WfgvqX6UZzxAr1CICr4fhqbOXn1sASvyNOkqe1K36nf/kOh1h5DUjx91xKKK3zO0
5FNA7ctq/rLkMsc2xjYqR11m37B/GVgB8GLye8XVYIrBwH0uzjN4/qYSlwBI1IW/
E1p+pLrezwFjijhXoPc0MSf6MmCWv0QUzdIjY5+W5bAttE/Zb4cvOrAwFZMypmpA
8k8PsZgHMI4LFPPBRsK6zSuZdd0oxZt9rb8lh5bbkksjxyXH3MOFfR9sClL0ydyn
i7M8UeaxhTaLp608nnWtxEFOqIBynS8W8olH83oPKOTS4JYfwqvzokmW6LiF/jS4
MSmWHtVhSPOYr3jzWskPAeMNG4i/ircVsmagtzHMViy3+Kq6pRInKxkz2Mn2bi1A
btVfRzjYXbgiXMJb4jE9/sB0LgUSb3gqsfwnxi+8b6DUN4MifMBoALrrbThmm8+/
t3R1gw8sB5SsG5sWAryetsfXNy0452stY8Jonx7to22qoyMRizGCEtZmziNAvmBA
XO4sOBooa65duYzrhIHDtNEOossV2mBYGNv+KAFxJM63uAPrMa91O8tRISlmjD1E
Emff4WAFHhn7xu0RoUhu9ZwQwIz/8szjyM9nEOUjQYT4RdRgpGR5Z8SqJA2F/SV3
xw6Xmzly4OFN5rJrBjn/3o9rEfcvG9sFIFEF4of0cByr0aGI/GAE5pjBdSaKUtZ+
y2ZvwUZs3BDkq6Lqi3Hu9g9jZ7XtXpfh67/N2cNjtt+9Q/sxThhg7Ht0s2m190CP
bi9vq+L6atz7EsDybB7S7M2WpOyIeRWNszFhEfR1lnX942kivQBxCDivs941rTtk
9HrXleGUoIKAuUck/f6j+rYr4PjgWcdit5GhtlDSJe0q7Oc0r+spjX8y5N1o1HkN
fmrLeTYvQ5KpFsbgQRgvHJvjrxOOWCE0DqAt8zfSHVDEkEZxQhmEGrlxoahXL2gD
1JGhTJIyXahBlVjcUnmnpHW3d5/CY8zN2p62U1iPH4rJitQfQanQaLoIgCAFWboG
UTPQ5qOnzzxt1tJna7G89VATLApmEVYntkYLtm6Cr/SDjcqpCEFGbKyqamJpvYDU
qPfmjl+aOg+vDRCoGJlysTmrLqsvcEmhHW7ina9Uf0LzenSiYf9cqS5s9uoScHPC
aM7Ab92d8ZkKmhLK+rnHngzNxdKPHc1jgqsd19RF6aQ+8rUKogqhQ52hQ42alIqL
rm+85Jit7z42o2//gbqZohYGzC/73IVLN/Vhh7sjtkhOd6N/9OrEk3r6SpL76sUl
TbGiIh04JAx+llGU30P6BqB9B7RpLYmZNY/htdAKFRw8CJNHAlEZ2jcLDGtoEZmr
xy3bw7xCVFS/GafbvKGUUWbCeEEE1yIp/21TdME1os8UB+mi5tpTOacY+W3tdXgt
/bbvr+0AcjlKIZu7shVbKg3OAUS98XSYqWRPETdVA8gniqQ80S7YPu7E9scxxuPP
ua/bcNWPEeE/FqCE4jGq+ZQaMTI5/dcsoqo05J71Xy3MxPnjavp15kV4mJ7nc9B/
7xSFXgZsa/tl0c9COo609fLfHTaF/31wkJCPGsi1Y02Apw0FDDG1tABo5h2TOtnV
DV1wZ3P1j9MGlaxDSg1HDwU3GdNos/gGJZ2OOw9rrjAg1Iq0smdwJkXxCvnnpe3a
BgO9Ehs2MaG6SzTHiKEHKRt+M8b2TV2oiw04V23Gpt17E1mFsGwZA2QRs0pmp6F4
7SdQ8SscvAAti56ZOBLUAyX/7HFT0OYAaSvpRIYg7lfOU+ffBV0v38tBdxjjP9ea
dDjaX7NwkGhM1YpUqhk4dWKFIgLR+5FZBBzx9FV1CxMSW69vTUG/xomrvKttuPuc
zJUpKE1HDKspn/WN+rmGhRbgBIZcvk+Y+myKKGKZSgYPEe7Y/XD1EsEskxz7fC2Z
55g/6MrvQz9HSc1vjn1IhXCDGPZQZsRJwGI4SIjJVKkPLi7sV5a4b1dJsaIogDr/
0pxSbuhEEhLHD2DtAtzCQFfzrb00FCUlw7g5GVMzqzSAYE1eaTAYTcMXzs7fr0TM
RBY2maCk5AR0jdidSGtx+244gKz3wkQz1EKi2ASq//+8ZdTccRy8QVA9wnVmWnCp
Ja5jZlfrXEQf+Z+SEqjxxsFBnuCuNh934nc/6tRvJHYvt8eDjqIb+ynFA43YrUd1
zf8pbIajOPzotgqiB4r5RXe8pf2IlwM0OovpOOa3UPblS+Fc4qQtdMqAVNkI/lxH
3tVSpiwzu7r70fAxSyG2F/IUWqdpEgd4BjZrCUYb+Ix/8IN1CvcYjuT99zP5AD3Q
RAqAmXEzu6xP46ZwgjZAeO3Hca36qhBDqRIpMlNFOXW8o647UP9CD82pVeLSpC/S
et/vM+WtiPFY0JpQJ6dJXUCSdP6gqyO/cqErvFjfwUCp6wuVaXJfmZXAlmnoOMjv
3G8++uParb9VAMcBx/lFz0fcnxxu8HuFU46LQqIhoj8P5HoRewohzBb7U2X5WT4l
afKG9gX+GZJpXpqXQBSTnCag003ZUnC5Qv1VdywvTjVaU3yO5LSBG8DyNO9Scpn/
pZW/Itv7mrqdPYMB1UkcMjhyJHJA+5DFcmIVpULj8NBTHO0nZZgDh8sowXKmaxtQ
axV5cdwohJfW5tbRmE/OOPGLBdnYYQq+aVB0pUA2nFBNa8/Bg/xw2IBLkAw3zSnk
/jUld3XYSkbl0Gsvq6pTinIvW9oVWH6TnsxYip3Km0/05jag/pCDOXHqyXIzYFck
iiEOC1QcFtGeeN8erj5SIChkImyc1d+5fWBrS42bu/SyRGSh+7RpqGdFJ7h6Igr0
5Lmdoi5tjAc734R+utN71cGDcptr3SuCx+LirnNwEE1j1azYzNWVo5FG4dyJT/vf
HoGnvJrPaHkwpB3imGu3CrQvUm/Yg8d0xYxlTEzPugr3tnfJ/rVkVcBu7i+/pSYk
zq9qSUViEMSg9iylidweoZErNbKlr7tN4/BGKMJ8wBByqDYyndnoPIfkyKaO6WEo
AepVMtPPpVgWosa/LYb/LBXhf6aPQ4FGJ2m2Qb7265f6D4mjeuzLVF77aGQWHHMK
JDdfZLFDt8vUjmesDgXSWSk2cmg1jcPqJl/anHvQ0r8uczV5l+XOyP+9o1lG0d9j
s7PJIOuiWv8ZdLEyN3rQr6IAqN2v3s8UY5MOG5UEHtESTtgHtiv6hlHU7/JUMmFH
/hCdeQ/l9jh+NxV0brBehBf7Z9xqx25l1xvksPiTHEtfPlEOH+EJaglARm7Kissv
ehGtnogF12YlyvuKLYYZuCTaVCj1bS2mRX07jMjue+hUSEOsXg8Iqzx0sUNUktgs
Pd/xgJ5ivPqbq8lVPEcr/ytON/VmqaorOIM/KupHvEPYxl86M4TpX49hCUcviZb3
jALL9DZd+E1wjRDGd2aeFZbNeO0vsJ/wsso3I1H2BFj5ZIu9uOk2qW/ccUAytTKK
QEvGBbu/zel3dFKPlIq7CcWcJFvYTKVMEbafcEhOS0gSmiHmtJ4aG2+75tLLzQva
kVGQOw+mGvnsIXCYVKn7XqgXI+LcpxwRDvwhcD24YAqBk2FONinbk5sBpNJj3o9k
cL1qoevXsnOXHb7p+vWxRgiFpfajQ2dpB61Yf4b/vdiRj3Y6UJYBsVtLn5uEOa2d
AvSUSBaMXQgyTfH2vhmxkubAQuInSp7kveP4oRPzrx0b772Bt1hfQTIhnV3l0HoW
bB7T2GT+NMVw6JyHI+sKAhqjGJCar77xqFbWWyGpyUQNIQnt7bf9+USgnHgN07wO
pz/C0cXLr3jbOSqnyUMdzR0NGU8uy/ebRmdWH+EWTN0TJSSPX3GCwn3M/E+e9tJQ
otMaiSoVhZfIGzOkaTGZebC97Qlv3F2p+Ce+mrtmrXU6NiAL/DWM5vUCH7Yo+ZxO
L/Ebh/9ncZNJZaFBD6xJqnrWFW45j2tGhKJTfsctjslNNWgqzNlDcWPVBEftKk7V
Pc1kPQlFJweqhKK8TKKv+CJGPs2Uv8tN0qBeAEgN5zENSctfg2gX2fLMFSdQovS5
DXevn2mfy1Fg6mfz1HfjzslWGP4SSxldrzNOl3XvOMn3XhU8oHbW4o8l8qAWy5Mu
PP/JLoU3Hnv5aQmvdL57ClsL+naZdKDxRB/NopTDjXrBk4u9ploFa4n9H8BLDd1u
TpUl7Fq3bSa9qGgCxwLpFvB1lnGljg2xHLb664BFMwMo5dBiTHx8q26LH2Dr/Br9
HDY0NhY/1EcyBBz2nLra5iuHCEmDoY9NDi8fy0KQonln/lD9BU6iEKiLvNXS3nq3
1Lc/3I41bvBbw9+FhS39BF4dcuOYEV8kRk0bre7+g5482ruTsIoph7m0iXC4CglH
H6l3xJBrRC1XM7NT6vxdmOSatmGYjkR0uFjT3rz8DgCAfBfDCvMqCz33A7/xd/TG
7HH+JgTopKpmYBQ/6YJRm4kFPsG7vZ2/vZROOvAYnZW4gCV/ADqsoZqWE6pwZ5yL
3dGgvxi4X1eZiDfsM19VRP/ysoL1qgJWnN5ZT/WnSgclsH7R00T0iUNg9OwpBzLy
eyXmbSI47K9fYQqAWftu1wSSjmkJx5CrW8bRHfP+Oi7ykayh6SuII1mQHcvV7YwB
NElYB6QrnHhsjMLKbBlLFBF6IeMUZMgO9RgYJJfxfVp/KrDo1Ybnd9b8mQX5egwn
sN7D908dGN+rT0DpSbixfxJKPvQXKYfKHkYo3ObQM2Ir8p6gZGoLkG5FVv9xXepv
lBPbsEIiTyGLCoC3kOxvQrym8+XHtFcbAtESACm5vFUs3xZ6/YqRz7yc/U8tdlke
dePF48nu8WGyWY58hDHMl3X25+JtbGBoc3/+BuhM5/AXcESb7gw89DmvXEY+1DIz
NGDxMfASIWwHzzPkr3DFj4j94iRCIWd5ucptoZjsFR7mCZGA+YSrGTXCloM6UIFR
+JypKo3lf/SHixYr2DEDhv+EVb9UmItQNu1FiDQBzV++EoCk6Zr1OahCxaWZDz/Q
kw6PtYUqwR5dZVBVW4SGfKeAOPEYytU16SoQJkYLQQLRjTKgoNZnujRMoIe+YAEf
3U3cEHBom6q6oKN0iBAada0xtpE24l0oSQ7CIr2TQe6NNtmjokdsuyAk0F10wcAU
/hicsxBwMtgoE2yTpSDQvkK48Hl9hjIlL/u2ePKM6b+IIG+5vySNUTDZcLxK0XNL
7SXizp1rJiJ+uuRnsWGzI6fJ8rPHspgKuTvEVt5CrvKFfRkRlG/jK272SqfnTVYa
scvrRpd2sh+/rQjcK0awKRiMCfQVOuzwg3p+hCkPuGn+mCa5ZK5xKfBcNvtSisw+
ho5rehE4LkP+dq0kMiQfwWO932XyPV+pKKXYyFt6kwo7oTV5tHc5/AbnWf5rYG+m
M47VGareRYcx8D5KGvspEiWuA2ARiuSqzvbdH0KzSPgwmXPKP/Sp976PuWXUO8Us
HSr8+jcgEoXkGeMMjesHExh+eIxEIzEtsdYIwhnmQZ4T+wf1J7rUxZ/wudRX+9CC
c9NlaS2KhqCzpO1TeeGmB74FWhXO2p2JJuNo00qbDWCdxkUutrZ5tTkJ2QBVNm6p
Kch8CSSEkFvT/1IfLmiK3wm9uOBAwFYP4D9ETP98dNIm7X7dpWUa/GbvvKigTKRw
hRmojiQxmU3gV91aD9wzPfPQ/GVX+moB8LMtyZixVrIhosaN1k9pixT5FqAvBfaU
3Nb8XkxeW7+Sg6I50T7k+YJPHx7oaWg5Y4+rUtODv2wO91Mm4PRxOS22gHKXFfHQ
HfpAeilwMLnDSL1KNDFQh7fAvc8yslNgpSgB0XKC17RD6zF02R6ru2kt1bstXHS3
0KLqjip7uF7Y3w49B430Wm1H10i+o4d8TAFjhL/SJkCQXHVz8rnl4w33K/JdL1JS
1a39iqlsDUWCbK6uxadSfSLNyBAuvhaB5iwZVAXC/+4N0KmI0C7rMwsutjJreuE1
SlJzu7cHutlIuUzMsl8f5PEWX7xcvGKT0F2MTARTLpekSmN3EjdyTmEJThWa5Xrq
iCMayg/+ATNt3vxYyyDf5fVBK9w0/RdYNW3yMgLj0KB+tBplRgcy+hQBnrdjMZ3o
HmCMVbGCXOXBePZ/IK0sDhUS+Xo4FY/zvnEFU3d9WR3ORvNeiIBzKJSU06U0PPzR
IcPfM/Ec502EZMJRAtKmwgUl9G/6Ol82xSBPURTw0pyCS/WOj2hZDhfnd7FmjZ0S
8Y8zR2Nllflh77WbZGs6VVVzKSJ31kCGUuf21ZkoA9n4N4QFrCKS6azSttYQSA8b
YK7u4Sczfmwseyb1br2gPyioTOfT40l3iGLArPJjxA4jzoJtTcB6phb/qepEp3x9
CeJ3FKh4Z1djAbvKfznbzQmTFSoUX1rV37InFrJGSqlbqaXzIGU+fdJsL0WwQSQP
zPPI4u57MQFjIQdCokkH7+hgRmTSNHJyOImVTTu5oVHGMJiQvFqN2+EYKv0ci0Fi
kvWwd5Prd2EV20zIN6bECjyLYc0GnMON3jI046nlEf6pYfCGivgg3rkNKpfBHWz8
3/36wK1Jq61EFzhC96NZWEXP5uZ0mJijhN7/COkS4N3voQRIsbR0x1MQ5SAwEMia
K7kMb85xHQtz62mC0B2X0Phhtqjh0n7wMzWR7kG8BvYZAnOwvJynDXQYdyVO2Csx
+jU8osV+mGzEcgVmqJgttgrBoLSIMEmAl14e6iyIFuSzPGnU++Yj7HDvvjKkqk+P
gJ1urT+Wg6HQyNeOyfraiwQImgqha7mcUYEu1DRsfl8ZA/lwxgefDqMH9oSzJm9P
M9p/WqQr60xfBkTfcPj53syWz/K++ccPWQCLNf/OvdeRv1itNzfDiC3mA0pz4/3x
IMiD9t4N5hflN8rD03R6/9siEi7N8XFz4z7Ex8PHUFZpEWNWJIyURdBohkpRNGMp
P5qyetUMS7oYhZLeVyK6hgNoyTnlriWbdy9SyQ1cUI8zPknfP1dIVi/SxqpFZ+pL
FsgxCNkcXMak/3xTK/5xXH47bfFpMMUoKBxZm5xQwwWFE7kqVBUt3zruXMloAo1J
mgkTs6tjy0oADsFSN+5ngbEF3Uuada2j321QeQEJBEDk7CHw1d3VY8GkHqtCyv2m
dw1FeUSpUNSaou/tUUXrkz6pl1mMIyveZcwRQFlJ7Xmx/W3DbY+97FQQUKk9BeBU
4cwjaydgAMKM30due6ZXL3TuGtY5pbse1qT+43tNToN4RYI4b+sNG7vmhwBgyK6Y
CY+Su5XL3cXIitrn8vUu3hn1548h2KJwopn5/h73rBVWpSwtRI7qMkDu4+KOemHp
vfZww+B8tSvvWd7DRPOfsWf1EjVKSQCJJU9esvYBjkXzQ94EJVJmWszvBwUmIqwd
0W/zlbfqX5v4ysoMaA8OR8VzVn3UhXTkhtImZtXWcVcyQd7AdvMEgUkAOmU8Xk2W
TgMbvRknXPLfre8U+vAfgU/tBEURRAkaaMXDN7zFw+z4Csbt9gTGxYHTKkJr/abp
BYpsNqNecYDTGHTvmBHfvOtuD2Nlj91qNI2gdKwjRWg8iOGbLYFGLC+45foLZg1A
ZarJY7eCagMqgqv0UWm+9dswAuP+f4FmVMxXWk8GMIbNDuv2I9jZCYo8IMhp05K0
WN4KjegW+9p2OujMne3C4q+anv4d0Y8Aazjx5ARsnoxggI9uiWDeVEowcqURRm5P
QnfbKze1K5uIS0vdX/2WWdgCv6gBtMXD3bBfzAHWZuxMW2z3J+PZTmVRyo+vMAm6
+EHRvbcv2VM7dZo1vEFrwxV1cRwU9/jXaTKWgRjquoLSOLr9rs5RMluNWRKRhfPg
MkojUmbH2MOmANYZRjEARqPGGmpEDuJhtn4hgfAUUxZpgQZ+bs/UjnYmPppyp7NI
jTK1cXTqEKXPcc1VDle32YPtNOTMBgLyrnEZl4t1jJ+nW6G54lCHfFhVVAIgD+YS
W3WJWsTHC1qhC+wfJuqA0Mqqn8Vz7Stoxjx6HWxDHwU+0mIYSSR67WVNu8OK9AmD
CZQcnkh8humQbm/SFHX9qDry8d2kCr4VcscjQ4ZbHDVZ7FGM8PsWmDpiXMGI4kzh
kM7qY2QSJqKqTnztgO8+y5juo263Le/HxE0kJUrFDvEdIPtMWeqS1o6yCteThsT8
VEe/fWgAstakmQfgDgqY3GgjboO92NQG5WlGDO76bf1G/ozKDOT098lQzYWVE2gw
8byuN6Xgpi+L0gZ2TNwvE/TJNeYJ4MJ3/s0ZDsyhgBMWFt+WDtKh/rxUhjOzuRs3
Y9N8zpspwPmEgaQP998ffoN2HG2QJlrS3ZnVFXI99KQkjthJHiyMNi/Yk4t/ZaVc
QlxS/c2k1Aw61BwGEWu2TdV+R+v4iGGs0K2PaLciRizFxJfSogKcIZDlNcStItAG
GeBWMsmPinqaLB2L4he6n0S8kG5rR2tjQHlMkdYXT7/GU4YqlGRR73Owo4Onhfc+
Mw/jfvmulJZCbox9JYh1vJ3wMzB8n0uHO9DCVT+g4NXq/0yZGiJiklD9xn2No6hk
8UQQ1G47dcQIpEqp1FA/zbPbAPYI3KvMD39mBuUlTB2Qt9NZhuesfyapyX8PtsjK
xbMTHHZZFzprdZaxICa0d9h+Ct3T6S2ZmnTlOaNbWyeo78A3fLDsx6PmCPiLuj6J
zrguEdx/qZIIYy2mIY6rWjFVWfZYG+iJSrxwSi4qGXLNWGbPwCqceRHOPZKvh9uj
OMxRQcavTTLbDPW2KPNapzCVhCGFuBqSN+49PyoydMcvhVU2+0qw+eWjzQZdP5pk
g5C6DG48uszaQrD9TpO7uChr4TBd9kdT9hKWMA+5nfpi4huIpYtLBUliyZKg+Ogd
AztDtuAe53J+z98zAVbH/yRQFagsUrARaeF0kXyp3EMxgkJEkgwBd74Y3dYHLerH
OJu/iMMKD4jAYl3Bw0l9jdQe0Gslc4IieViMbrPTpBGnRKs5PMxEU5dLdA8aPEud
xuu1OWTxr+I9CPXZCbLpBgo9q4gteNQdcI1v4DLtv/EUtHtRbtLIDgGvVGhY5LYN
dBQL136rX+Dlc5Y466hVSFzvBDhrtZZa9zFk9rJVmYdvWe9e9XQYH2PKLD6uXqhJ
sN06VZA0Nb4FGNRca3uyxfw6C5YHt4i/Hao04Bk2+SMIYH02MlHijXSFbhJOuuqa
NHzICJavX4531cHLgN9yXqdOPp09BtPT91ypw31Z05g+CC8imfR0awTdt7iCW/To
zv2hxnU6c162ztnBX5XnpN60yu52dk473YaE+5KFgSIp1OlO8po9CGDDd1VehDAf
mMObjDsRYeCU11eYseu//YJ9sFGzm5f/5QN4gF8+6E17InJebbZiq09uXdbaapCB
j1Ux/aCCpeW3jiumJdcIYHKXS6/KR22dAK2oBpqxn/LPosjPzIIHpgHCfA30ZapX
Zik2nDukCRIkBxAEwMR6DoSRDp6Lwtwoaq3lo+AEKk2EThIqLGotFO9PANamm7bV
wMIOUHiyFEp8VhOl+h/COkI1GN/zdpciO21XtB7We6fYVxWmar4GcMTBqYcINXKZ
T1uUsk6Ism6+h1cqHwPlUfU1xNIFpqGWkCeKK1Jo+jIu0cSM5IglRTwetiCfH4Db
UAxh1C0MtJhtJpfJPbXtpzJSbNMigy7y5aHKu/UziNWySJR245csY/8U08b4Nb4B
V0wVTFbyHPnH9+3AzKgcbq+XNYEDg7c+6tqfdvWd+hICnW+voKkiumPRySMKzM17
X3A4Jz34VUrfNxstBxIeewcw2H79R0LtdpsThbO2moL4sRtqOol6X6cBhhuZs0Mr
jdA9+gvWaiNIxnl94gy0HrASi3TT7dbQsMuRV34uje+zs7mYmBN76uzOZ59GDUNR
REUodekg/2RJN9Ue4UJiD2zGzkN1rwld138xspn2vDUFHkzYYvpsTx8h697ZNghX
h9RtPkCK/eMxjmHAFh6HS2K2dEO4YJniSevt8ajlIszdh9EzQtkSlqT+FEEKomD4
DUsGHPNwjBIQhj3nx6sHOrGXv/H3oobak/bvOtP6kr+bvWfOh4+GMtyNGh9f9g2Y
3uvaCZsJ+6KodlvN9vdJSWnbUzhtx4T7DTETim+egtSb5J7Y5OqAqA/jYfqwqDgD
qyaknG4jJFlOnkZ3OZ2tCJ4sU2c4C4Q1ca43kAkwYFm1GZJFq7BVqi/Q5szfftWU
O89aN74KC4uF1CS3WMz+FQP/7HY+04px/by4Zpf8fbb7y8FuIFjTm2zV2CZh5KAd
RuCcWhrkV1/XoL6gQq46Ucwss1gPCDMBiItncNzeMtlLjC8Ij2m06N0ADLJunrIb
D1q34VQJ/w9U10TCEXZKnbN4jRI+PoW65iFuU5d+xMSymbQwfYb6uBDAKUT4QlSf
VsZQf6n4rHwUGnKMuZVjTeL4CkC8DVOacFVG6Vljs0WDqzm77zlk8KM/6P2VEbWF
cIZRXSQI95fCl8RPhqy1Knvi+27io/Gw9vy5+tyFIYp51o6XVr+TFHzJfkTV26YH
XgcEeEnRWfpJuOuKk/3tNLPLd/g3z2Pfk+nez/2uaIdaeaTGv+IEkwqrRKMxfwjL
onB6tPDhiqz3YnLid1tmH/GWUyea44oEbdNmYD8wSb0EKqE+kjx7ppzZ+mfRTskM
jFi5uvPub7CgOOBow5uF0//MapCUH2c6tMyBYrRBtwW+MA3iCfhGYRCgq8a9zIfJ
fukXnqfNFLc3xBwQVw+ScEsTO6gDUVX3o9DsOPyvY1Jga+xCRRyUvb3GYOk64h6M
/0v/Hk3YHQs7lw9wLs6Lsn4E1nqg8EvO0k5VDrsW21siiLVjmIbTf/DWxIQNHVcS
RS3Qs3iRDUievGCW6/rWFEFOV0UZ3pksW18LzAXpJABmm5wVFMmiQufIsX/Rdloz
P3GqiG5NKP3oPdDPuV8K6flHLNmFCCmSQZp8P5cqZApfGbFWnEsJzB8zRE1oI6Zd
qux5nsvgrWV/EH+7Sixn5SvBDLXPzh+Ys4wTwYm8R4Gwdabr230PGVRsopip9Ki5
zY29JfZdTT6ddx3TH343LmFIZFxdCcMUTqceaY8frZLWZmmgVs+fvAGzd16gcdh5
LH7vQsQOfzIM2lLH1ooyysmi8fceX8GIcSpXq9o6p82cfY5DDzRwcWo1rlBuWctP
eJ+MFyxW+3mhxK/87UzMVGExTR6UWPHp7emDh17rVkOEau7uwA0vcsWVtKhicLhw
vkHzlM3/8fHhnfvyIaks4nnXhU/DCSQ6hMqiUyyrSL5hR24Jm/uuw8yHU38RxcGF
bIR4QpoYmt0Spznkd67Kq5ZEB5MMzxbWBA1yxOl1uAULufU7ZuzeYwFgV6xf1Mz/
1FrX7Bd6YcH+J6pZyaleT/cMn8xuSbzlWIKWTm8Gisdy9BuI5PSCdLObtBmROXQq
DCc2e9WQWo/Vv7qHTR1I2jdServQCcf4qmiJI2UqIEjRafQQqfSvP0RJyL9kEHro
WBXqg9Mabm7dSGtHDdYwJgmswt2yxf+xCwuJrigv6qtZ6u3SvGIYyvyYpzG4b7dK
QrOnD+ocooZPme5i/6fg4MjIvNlnCrCscANkl2rITBr8xr5Vj79hMHJ/VVlK3Bwr
IXDTLyUxSgHf9aV7v6yB4cM7ccCutdyqPxw7a7F8RxhwvQVN9LjUEwmujQlU2nhi
A+7EfgsF/QOmECkTBDgb+20c0x/ZE0gb0qFGubMSMPsN7Krf52fvYJMJ5VKoQpt+
JVijHP4ADLEhx++w6vREvHdWi3M26aCGkL8ObvYhA6M5T0u/4h6/bPdlWwUkW6Px
Ml7qDK5zc6RHCxtO31Lno+TzWXvw89h8pfrV6tkDdTqJCZUhPxIkUeY5GiGVoJb2
zOKr+PddM5osOL1d2MmTkLoyL9P2GNpYBVNeuuk/VNd0zNNByqLC0phzgMfhI3Ou
rd5QtIUR9d0GdKNxzrwqdWL9sImtLQW1lO8RCMwdXRUqI6p1XskbEKwyvy+BPME6
BV+vWbSKx0p7Z87QmiZ15/vMsvlqGO7VeugFw8FccenXak5RTTf/0r/UVPrOFnHU
drhxwa9RPAmWNojilQjsg7eri3adqIx2jDEB1s8gopuDGlMWBb57X/8ciTAFyDO/
77hLNA6CgTEYKfo4XUkLsR13ZJA78L1PaofOxECkbf2qolWF59lwQjW7s8u5Rjnw
A4Xwpv2lcP6QeZ3Zs/vf5FSM5N2txWge1MhJyXD8yyIpvI8WtRB0f8ZVhIvcsoYz
0blmmu7q3g064wirfuw0fyKuFU5Ha7BQTaMGDZqirzcq9nJ7QHz2m498TH7G/9ec
KPOJnMeO8Lxv1Fp73l0DFVjcspYMR4nYhXMEm0GjAo3VrT6nOkCibQYJotq0MxJf
TNet51mT5RisgDN2L4fdYW68S0UNKk8Kc0r8LA0q7zteIuBtc5BvCz7MGPq2mfeY
zA42fci8Naic1X4nl70VHQQ39ivaNllpZhAEatqrOABsPu1tMuD0hblJ4Kr8qoIn
TB5c0EFckOZXfL9nBE1NJ7YPCXdl5bKehz8h/W5OJ6/Gjh5/pOJtMgvsAB3bJcBi
sAsVh7Ye8G6u2aUlVShkhqrRHGtpJKX+hNHdUy2gKqFq7vld3GPahGTQWepWXlVO
QR26liW8khLSXWytkP6Tbnd+ggyrlP2RuCYFmx7kVnrTQQtDPnIqGAgjqlel8oJE
AKkc1lFEY4xBrqcXGE6XHYjHW4RS7tw0P2skZANSkeDw83BcOthLVPV1+67ogXJb
b6qd8eaHA7i51VnQKMSMBQOX/WXyBdou0HsPfyCy5TANOOJLSJ3JEiDNfu4/ghNJ
o9eBBd+y+OMhPj7wQYnGeEp7B0P3pmWK7hSUn9iH2Q+kXFd82yBNDnLqLh8d7b3t
8udoGVRqFmorJNxLNrpcL1441ZykCV1B5qeEHcfqTFb+ytnC1OGF0hTq8+MAUMKy
2mt9ffK3kzLwq+QfMghM372dohdQ02M1tGyNL8sLS8nt0EksGRwQhC6z7v2GG0Ac
ZsXom1KBDT4QNl7tjNnSKNkeEO4OgJk41ZSd6HcgjKGEZri/h+FE0dsU5+5YFBWp
GSvMVDRuYajK35GI76aDiyEpfRtTSscuzEL6AYwqFLshSBYW4RB1WYQQ0EDu09CD
/oSGvKbqiy9f5ZBwVrsa+rnBra6To5V+LPduE5CubpjGyHjryhVWsR0vIO1QOmxM
JvAFcajMvvmXjiuCmVCf2Pg6xMRagNCJPlY6iJ3A4KmomsZsjiqCNflN+YnHWQh4
zm5YIudHOI3Sr/AuLby1BLMWbc/Bm6FdUOO2ABOrmlLDvTdjCbrIU6/0MrdO2q+U
ICmBls2T5WtFEHtXi3xeYPPE8qf27luo0dhSUBC6QY+H1JFkH072DT0WgM+K68bK
QulpP0hDY2DvLTcbu4HAQ58K4mrfofE3N8bd1AF6s/yK12wHsXNPufArsngOlJkL
PARRwZjbfeCyPoSqsaSHAan3aRNZsSOiU23UsFfypmAkOp3K6WppXw4Hl7EW2+xJ
6EwtcpDQOSYHgHttOaS5ItgpL+lhku/zF+A7iq6NFQuW2Sx47g3ay7CnQGjmWUnn
x7EIVarbqPGpS6kOjWujrxVI661OVgMBG0eG6OY4+vJuCspc7mEhPUM8QMxhPMsR
2h9BSgC9sn44SsmmF8xScS8FDAkKwR3XFt/iUfsjLBjtKJV7EP2lFYUpvVkDuQgm
n+13drGTFLLY7jq9gppmMerlTkWxuwtiGKf0GwpiyTZD6omx8DVcRUkjAOPBqxzF
2hT43ozqY+D0nXkvewmivrzR8xbRUlF6WTs6fvnzCLxeISRoB2o5J+4dS/EuzsJk
Av7P6QNiEoIb4YZEyxo50jXgHqIBddZ+UA5MExiUuhUr0Vzf/ZZXZWEfXs+1WvtJ
Tt7aNHxQ7oFQTJo1XlQlCHBcnaYExSiX7BKJetiSXnnZcrY/Z53/AkWzZw8iFrSs
f4WUGraOIPUcTbgL8wvXJk4BRlgK2U0hpvAvD+hxU8Lgr/hoySBqp6iE3LBfE8MC
doStKluxzGx/AAIPokskn2pk/OHi0WPGsBGw/9xyxc9ZYbBFFQO5Pb9o6AFEZp6m
LG36IxhwZPcsk7RY0K0V2+ohPVFoaqn0wQ+TvQZNkwE5tOg+YEgsHxS2iGjHBOZc
7fjm5KbmHY7k3DjSugH+4C8yHvlo2XSpIx+MNCnmYPXXb4YHSaDX0XPwz2R/6mCK
lZ3hhsHmkohAEP4w0VRcSwbQndw6o0FAJUjqmm1qvI9ZFh6GiAtgn67N6qFBR1YP
JNjqflyRjW1ZNIrkGaauPXvynefZ0n52w7GRtybx0MK9FlO0KeylzKQf4vrQC+kq
qusPy8jrTQE8iRsiT+d7Gb2UEtfoMPm8cKLL5X/eo+WN64m6jXTg7Eog/L3mLuh+
UpMpRXHKSfkzbs87ct3r5xYdwIIaN2oU0rdGSFji35s9HOJRssw01uzT7831ci7M
ZpTY8fHlebktmeSy7Qiw4A93oAAcPXlhlTBg1zfYdt6sKPhJDxqMONWlnKTT0Pgs
zv+BEfjAk9n0exxJ1zMeVEva/uwHlRMlzLXww4IypRIcK8wc8SjGlK1mCN7WkhyR
Lf0TzhnKW+m59iARSwgf/B3fnpkpTvwJVnm/zeQG6u8Mups41W30eVqHEN/iMPX6
fCgUvY5XkW4Ju+q7ERG3FcMNlAquc4A3k02Fzr+k+CXUCx5SxwftztogaEu0hk21
MG9gIrP/J2shmJoZHiFrvlsnPEg6FfQt9o8P8sNolSTW1IKR3SgntXrZjzmeqif6
n+hQIXiBTVcSt+PQEmi8iuCdz3L+/CUwSR9a9GhA7h7Fuo/g1qR0ugfV7/H/IGWN
LucZe3fhjiZ6DlMC7aDCE/DMQVNEJkDfwKytqgK+JbrO6y1eTfJDwqLsnVCNNhoR
KZjE/h/zTa21NZqF0Vta+bzXzneirfR1EPxn+DwQsNyIs2cTVe8vgWGLEg1nFiGC
ShtY65hhHbIlsv3qC2AgTjbeoU5DIDf6xModEf8eR7ZDq26BWurXlwh2J5+UOXB+
ms/Rd8dAzv08gvygwkI8l2zbPZDkBOJpGSKgV2xt0RExwUUtZT5ij5c50RU3XfVb
60Sc/G5cPRs+q8UNuD+Cqs01cq1VYCNvAGQ4fwAQxcD2pYLVPnPDGMZ+Id7KAP2N
htgzF+ayO5mbJWejDHpGsJTNhwSmXgx63NS/Ep3GC3bdvBqWM6TtcvlaEra99mnx
iFmzguDpt54OrCws2k9M9cq81NJkCmo0Q6Y5m6NyZfnlUoDpy4YbcIs6fKoX2YI3
RlRXNvsm/2Uxt4/zL0ceuyvbvr1NwTd09hKzMPmiwv4dQ8LHp5F67zmd93KU46Q8
WOvUV1efnODGmGK+nFd2r2CQYlmDnYVULTlRJK74j86Q2jjTaofvYzHOXOTj/Sf9
/hmEuo8RpWmh8EcI9ihLO9JtXGjecbEMfktgP0mwOVBh+RO1NBOIzi5OcVuVKFTS
jYT1vZdGZDY2vRKhRkGLzl4nkBtjmlUoMH7GN0NY2pKrLiki0H9UGnqjCaiKqgM/
9CnNrwbqaxcoE/BfjL6yrGHVQce5sc9HbeN6zsBdoXvTtevf98VL/Sj89PgmW6xT
2pRwqzaQ4aVH6w7vd/0QADZLYWN2peOhbibpaUpMFnAfIPfWUEJUs5/+OsYBYxgI
40mbEajE//xOD06yL196YIQofU2GI2LaVvWX0ChWKLYDq0MJBz7Z/M8LFeKXlP5L
pJCZZgScxadjsyneBQHoVslhbuolXQbssJWf54LdCFd2V5UtnsFaHIDU7IzC/Xtj
6BXBRoF1AJmsKvvTa/2xkPG5pIswig7nzJJpI0V+NV+e52nV9ojfw1Ewq1OylSOs
pIQdagWx7YbP3ilJdX1dG63Rt7sb/mcDEegIbDSgnU8f/2Qg92kZaJBS+8KHLm2w
Czu9+cZy+KwK3jE9rBF/8ftU4omUW+rumF0/hi3/zvHaCtpuC6rHVojf6X2qqym0
PgH+GBCE8G8IY2UNBQQoHMCx5okdqRCT47nfDhomJEuR6W0c2NDSHEydxE4egMRG
vZRgBLsFUyY69UR5MQCgpZMzUb1zS0xANV12ByqkMM0gxwhOdjaP0tOMm0Ivwuh7
Ks/H3sNrqVoWx0z9FiggBvCIdXOYiFXPciYWM9clRNMkujWNtPpmiNOPbVesEdes
tmnafYggy9y2TDnZZyYgMHufqlEpVjJRNjjkN4t5BAtui9cLtfDfHKX/HTZS2fCL
L+Ug+XGPGgeizrR1rpWzaT7SdNoJRC5Y5g+fIOstNGKEJxW7ITNsUDzeYqqQXGHT
YbJdKSrFRykkkHmI14JjWijSGyk8XPLnOtN8pYEzVXAkHwZYXIKh3+8U/E+DKBnH
amfVimurUL7B79SafAY+G1jivSRSXjntEHmWXdOSCx/GDFztKJVfHJ1OdOxK0BF3
NmDFSt9KfEDDw7cu/pzIzyUMxZlQ7c2CGLdXCcLuRbBylO65c6Cf5pVDiUNI7VNd
t/QVC0rMKpWZga7FJnAUVPQDQt1q5bfvFo7/ZBCdP5LW8C+yRbNb0QlmZqE4qXYw
K6KCSyYwtlwCVc9Va5j2Z22Y+j3rK8nx0kJ/WkcgmUwoVbEc2LrXoAnA0JVF7Gog
xMIvk2kn4nvCynplD0VDPZNsLFxN4gBt0qqDkMgW9Ca/FMLoTKpGviJJXK4JJF2z
iEOJZ38w6a2w9LHN/PsiCFhQiwjG9T2Uyz/fHwP+5jO9xjJ6dYs+vt2MCqkKvjqC
X/0P0lYx7ldtOqmuv+f9o4yJEi+EB0GmgER4pN4noJUnxxvyT8qO3G+hFD6wzs+V
HatWyogi0Pc7YiJYc+iuhtXyb4tFJrX6K/VwS5Zuk9gWgzqtd/fIszyg36AvNeVd
KajqZTnmaPWt2UfTOMzduJtWg/dPghon/PrjsjVhbubfNoxz4Y1V04KurumLwtFv
9Ny9BSo2N+IUa46ZY2tJDr1WQSxO4a5PMq5bIvhc+qTqStYOUbkAIkf/X2jXQVTs
BqIaUt1sTkGzmWIsjHhvcVqNlxQ3koxlwUeRVEWlCNlEpfxNojjuQfvscGhI7DON
XCxvT0MzeY2xtYFZADegiwUADhaFbWJdIdVRLYeoomnKcTqG/fESIb1ZAh5yXIPm
m1uwO77ePQb3qEYBv4SkQWrv4e84I9ow9fApnudVmXrqMFob0QWMz72oY8HEcCLT
guIVKeiP3DL+X5HrcxLbGqs0CHzQkFKbRbWTKQ8zLOMS2+h3lVFJ6cx8a9j5qlPV
YQbojXb4hOKOXuGb9oskbUa2mw9VUbSbG9KF31Vg4evVfJTlY+Bo9PFRubgF2AMU
XdKiCThvhz+IUDfuPYiiWSptUlDGyxLzlNn6Rhi7qNsJYArgpKPqq9uVOb3xbj9h
oGLIgwI0pMgyFz4m0f/HnUaQa6H0flupDNozpMv2iP+BFAmKCbHFaHg3b4CNdwjw
QSBnE1UbtOwO5XhUpunP4UHvekbY6gp3UGFLkEFB606bmNPOgFiv+i89Rod6nheJ
JyuumR620ysKAWbhn9W7znD0PRRISS4LFCPTt+cC3NB05gD8UCj0VyKfH2s3apG9
gy2V86bxfZx6NfbE2tx5VBcGeT5iXuUB6YitbLV75SnX2wOlZMIqqbYxiwoB9SLy
Hh8bRL5ldGpLJwHuRKFjWEhVc74l8w1z2qNbfldMpkavgzKIEzsmsms1YtajFX+0
LEzXnlHVtQTqkZWnUAiUSZF9eYXbO3T7Q3eQdUvRpBwN+Md6Teo3VYSM/iCGBai8
gpdbxo8O+JvEQZIMSoKY+tl/bSqgjN9AAmg4MlB8O6j0f9k9u7Z/+VhhQt8FDNTP
3/QKU+eYO4xAnHh5vFwy3KHPGIaAIF078cFqjoEjtxWdKzxWyzl0rt+WM5xqaFv2
b23lI8/tY8GB5FWCHpmiUmf9/T7xtuzv5mM+cGYqlvSTRm3osY4dnFrGOJKU9nZe
2WRhh01xTD+inIhsBVITP/6RPjDXWiK3LvwGIa8dOJuvq9u9VFpY/ZQex1GnOZYO
OmHIVjqtEYqw1oKSWf0rmoVog1jUfD/n+/qyO+DNdBiRuvBrZ1i1oDJgGiGaGo4R
jPwZHQwE15OghnvCZPXqaLx9vo/+eNt9N8f3jPBwSjU7hAfzmWNm2OLfVXinN6eP
ZZWY2zc+hrz2iwdS9TC1jm4N+6Ns2xQf4RWhXGlfzzQyAJlW/iZbMXFLqEdKmNoS
UTBpzpo/DpbXBugI6+VTnAt1QlbyA31e1W3B5q+w7edUtjPlIr0PL9vH+v+RxgS0
PFID4XPLPEEjFg7d/XpZkE8NBZA7pNtLm2JG1PHu3l+XjrlXZvXSm/GP4pcp6G6d
eH1P/gHv7QFrXkzrNWFVzcL/suCvka1l1A1GcyrYDQbtSMJ5ZeyUSE8eHFdlmcaK
bQrt4d74PLE5xW8kFTK6QqU9Vpv5oHLDVLm5j1Q3hor4IW/t58UUFCEyxJuknOBx
BIgeHrM+gXw6cH1JrQ4vh8vO28upvQ11IXZN2WSBgN04Tvps3YmRjgVDQuwtbBu6
DU60FebGDrvE1AsDV+1thuvnWHK3t8MHmsDJnoJM1E4L5gHFdyM6CZ7rznR70RAe
aTjjByO/sFvuHwxaZ+udIehIlNU03zqNhZvbZV8zJw8IAhtp/hF70Ft8lgrBketm
UMr9W8e5WnOIrmzZ9HEALP1wzc8vKEMbcap2b5I9tz0zf/whgx4PK6/UD/6zphjn
Wwk2St72T2kgn8DUTcXR8ZHfjNKPrkP6qid4ltV4As3ZSIJA7nW/N1NAk9YjHIFq
6TzsgC2Lu8/iqVr0/vfjgvUAUeXcg85zq8EaZ8plwpyASKo+10Pzg1DNLcx3TP8G
703ztQor1cEnGoROVHKQInryryBMweEe+XhFwJofxZl1nigNaYBQLFs6fVqmCG3g
H5eFBnC+r3lLUF07RoPDZ4edCN8EC8sZzeiOMgY4/4tgkPz2uw0g/+CWk5FxJtgS
gMfSXJx+GgwicG91A+11F25d1+kWRAbXZ3vICj3sGc9nIGjWjXdhge9X96+Pejzj
botLMqZfegA4N3bA1W6p53yU0FJc49MdQzwVQFulgSdGA+IEosu0Z5MFwZr0lXnX
q6zy/9BP13ChsCawudDg9yJtCWOSAkrFYeTk6KOhwwjyqVsd8lB747zuGr4XY6Of
dl2BXuhVRtyGxpKL5HVmXOu49gf8bQRGHWumzQ33hWHIQoMAGMmMsvp0qOTadYO4
8OvSwj+OJUovSBuslcwp6TDU90ckwdSCfH03e8XrX3bZF8rJrx2O866GWoar+7Gv
nrs2aK8l8wxrrIMaVYj+WFnIzPm5uiR1UILMqfOy2n4GB357FkcJbEwp3hDoaq8k
D6yw+DbAbLB9YundZmbSd5SrGgnmk5YzvY8QyeGAQeZm52+iLAP0ehITfzZ+lNiK
8EzCEp1VDhaK30KB3b3RAMoQkW3j74NIkv1zs/g45XmkKhxbdzxT4NO6DFAh+fJ2
NpKUDzEeDqsbFnCOrAhdsvcGrXo5OC7DI3WPRPpEk8rAzTZq2ca4VmRUYITPb6oP
iQZEzNjW6ipsj2adFNKl3zEeQV6XHODiV8ITRoG/gFLpHURQx7zI7yqwbFfpzdDA
ivNbZxkbHsB52CahM+C+kbl4rVp6vHOla2BdRzgfoxZBdMv7YGFNw5Ri6IStR7I5
O1jZfdFdAAWr/cWyERX5PBtnBwOCTf+mFzpMPuCOQOn8SGpdEI1R4IlunP/VRKWV
z83BzJRFQA2WHU0hg0I+6+CProNtduHDSjOPkdMv9pz6uA1CFtJ8ZvBWkxV9c2za
1jiI+rK40+ar3KbblKp5fnQM9yZxW+pm40TPi2bMzhs/h1quKfw2ph7vq0bvKeqH
KBcf5CY/FufmVQRttCVQ3iccC8EkE9tFbhxFCxRbkL4Y6SmNSTM209Ux10l+FbyH
kXKEx8y594UCvgPAzfk7hPcIJa0hrSKU+CJSJE3l9McivAMReFDo6zHBaRSSoe19
JFhkDMamYBmx6Sl7Ws9DmSE2qD8VNuaUmnYfFz2+A0OWJmmPIzvYxUn9FWO6ohh1
LzDYFPP83lWVoQ3Xxs5TcxFwim+mrB4lwGIAfL/Xmz30+dQjFvqrKpEtX/h5V77F
Bvf6Vw1lrXTymMJPxaEFPqYTiI22aq1NXlICbGlqSwdogmRPSJfEiQBWeDXJC9gW
vbenGrXbv6SExD/kX1D3EPoOZy+r4XWNtuEVS21Hjtg+YYE6CtZCp3Qi84i6RtIx
Z/K/87kDw3Y2dVvLPKoN5Azi8mNfNiDBFgMGWvjqZOR4gjoV40GdkbAqvZHf5SpU
KUonMbI0jTR4mBvJCOfAZwwzlMlvrALyyl3u/idHyx27curnbCs1JO0nSmugf9Ix
/WW71pw3bxfjhH4yMItoxLpyno4HDi3euNEHUCme3olpn+GnHT4P7oOZaem3xPtM
L++w3lBb4OxZUnmxGeBtFtt/SReJ4F4wsd+YTd82/5hM+iLBv3SnD8q1+6CchJX/
X0CDOzMrE+HgfcPBfcNcZw/JxJqUClNP/jH6cf/BcELMpYBaddRK/pTixOjcnOYY
Ii0AEM5aKRha6wxRsxUBpnBIuRCtspkw8VxJ0aO9bf8w/RIMtJOWOrxQo8HN9uUc
+5QDNqvrac+P+AoUGWpwMn0knunh74vK7G2seDKndngX0hTlJGN0AjWrZl9d8Sol
Rx8oaSiPfg7gEK3ORgTOicJvUVwAtE3Ig7QbJxSCdICwct3ilGn1VjPvHIGtVhxF
jfw0ps2timoaQcfNc3IKrymO6bj7nMyVmbrkpw6l803elB7E6ZEB+0j1m+qRb9MF
eTheQj4sqMn9oTF0I6+Iie8f91q/AaVM5YEJxBZ7CiG+Aga4poqEqFRU3NyGhwQO
rcH7EBBEHf1IviBModePAIWX+JNyqCYAc9hJNZCCcP0FautFyq0YaNn47YXvb0mb
PDTlGD05nc4jSnRYuF8EbVmA487ZW/xhE4kHVaEOkTKwkCyu75BzhMxh8uYc1ftp
88tRssnrMm7Lb7Vf2E2Y8Gsle0DgRlidna667d+/U3rZyg4WHFsM33z3DyX8faYO
lBkfpntX58yCxqOt8vk6K/krSOUf3e9YzAXa2iMnFpsPEmSQNfGkVjW0kJ+QgMeB
NBc4o27pWHH8vZcGYe7xGDJ7inMn97rglcTpa/MLfYzonfE5snrI5pPwtyrOoEjb
q974/0CluWmQKl/R4upQxHKEGowPljgEzw7mCbyy0punrMbGjZWp1n3oEDVHP1Sp
WslTtNDh6ih7GFkkZZBwHflHLllFI2qPmiUBcXlhQ2juP3e5Rn01aaOOwz3u71DW
ytdwujC/I5092KAv6Dgp7txjtackwmw+uXXtth2e+G/dPkv8mXIBajba+b+ZYDs9
Jb9V8fIfghvMf8zlHKHveAorm6DbzHx8XA8p+KL6XHzUUa3o6qmIOC+4Ty4b0DJz
fQMkaw6fXcC5C5GbWjHKQw0O+3tceqhzR2OHJvZ9a/9olQjntnpVPEMp0RD/Lycp
6QjEgWdX4hGTGOFO3ifX9McNxF83MSbgNAT5wFTt418zp1gQw3YlkIdAge9aPoGO
SH4+vRFG4fJd18HwerZ8wMy303HXj+xVREhpXppLkxZ5YgF/Nu8HRO633OO01mGu
KAtYeRymLFyBZbb/7u6P8O8Kt5BqW1QHEfKCz83I6i4J1XElxcJ2erjAlFzar5q4
MfdsU2qfZxCPn7xUk7pe9JryIZ5UV14q6VtBSQMKNawR5BDecZ+x+lYFKElPq/Rq
/R8b7/1yvdbilP/16Z+lKI2OEenfWLoYGu1fBq+P2uJQp1K/iuwlnbh0fxUCQ8wb
QE6pKITMfrlLTQ7ZFZVHNcQGoYMGOkqh1b+nXOGzCarA5ypaQJY2b9GWQnx+zs9S
86BWZ6nIES/HyAdAaRZw82cGFKTwnzbDe7jnc38cGb95vyzZBS4bl69jq6GpcAUb
4UESggij3xPiEIDynt86jh2PC7mrvHW3hycvHZGiKj++Jx1uVZQrK/5/Icb5fzxa
OX07U6ZeLicBTnzZmZDw00QhjZkMcUA1t3pu6Lonozcht4hgJU34LsYKpgQ7CxKx
5bzUcmLMvCFv8PRXMjZfd5fIceh4gpTOarS8O36G1LNlGmhLji/DYN2UHZXA/6cH
zQOL8H80QaLZIIkHDnGRg6ZdCJ4jHj9Q1BJJl1ArqiSCGUMYj57o/Ropqth/6vIU
lCOKxa8fRdUCb5nqm42tqA7EXbDRBYksYNaJeK05O86dYWPHZoYonnFAH7GXdAcN
oxIl7ZOfrssIpLHhvTOoAyDqs5zjqLoQV39sILI/8pcjNcjssZm4AhqZRx1Ca8Xg
eFwv11iGycFGSbIiuaQtMuoeBzvnoFq/628rtRZ5Ef01wC3ensLmWggsgzV0EE+I
ManSAg8pyG24e1MiZ53Q1SQ28ebeK9w8g+rOEf2UzSsHGUn+W4X2kdnt7PTQkdmP
KCvfGuLhQe1kIIPzOhffBBOQSNXBWCFHj0CAgjxKSILnQRMoYKUbZ0SHj0LENBjn
FevqtTLLF7YcaT3vIKkGxtTgWfRyg+xkzg1p2s+s4IygDcrAtKgpNOcX+QpsjwQ6
+IguFdoDsFEFxnXt8smgWtfXGQc7ynFWeNhWCYV5LMJCYwPwtkl1ZHGE37ADN0BJ
lpzkYGFPGQXeMRpUnyaVeFjdH0oiVVoIXwFVpgl+yaL07MiPLzmoVVsKy5pval1n
H/IIxO4UE6kdOtfc1QU/1o1K0zn7+7+wKdNDiZP3pg0/hmg/1AJxFMz9kQquuKPO
DEUawOau/OFJaqmUz+KUuZ5uFR+jMPZY70KdBljGrWcHtn5bwoE/eMhrLL6Ker/9
kb5/2oIdyjrhcKL77UBmuEbMcGTC89P31wI0N+5TbS0xcnNsSCGjLFJR2DNg+yEY
opwIe4FWLMbXLOYAN/8Mp8v+JOKy2i6C+xJ3ejWj8s0KKZ0Dp1UIfTyNrbPY8LSi
7HYQBdGSPzmh6TBGhHmTBBtivJwgkcgwyGthXDwfsI0N/l6tuZFyy5zyD4D+GAin
jQ1ymxbSd9pFHYJnm9a+GKqog0JLWxHaLDWb+szfX4KSpn/rjVTlKJ5xlyCuUaTk
v7wULMuxu8ygN92jIqlJYidD8A90fp254zczhatEXiupGTDCPCDlePiRypl1vFoc
sRGAdHt8G2KfVVyk6IRO4m6+OQM24PQi/v8Qa33tFwoDyQI50bTYW3CSKgkgSOxQ
hPYXJY1ZIaNK80Dn0I8cHmIvlhbJuEZkC/ori1G88+sCYhpeYi1UKUh0zD7stH2y
LiUQB9DwxyGzgEe43EfjcNdlSypqUdeIJ1Z7jdNBsiWRivE2+q6cIquxWqQOlVvN
D1wco4UL047JBZfGpBz7rRZj0QyM9kWz/f9yiNpV+14FKGnIjS6DgUcH0xTBudt+
vzwumVf1UAfgpQ1djRpPb7OBwxfoFLPwof+YFnjuNquaR17EYS83kLytimFPe/S4
afXug6S2kPPQrLXeVdgoEGYKXmjQBYC2TzsSwqvTxCxJP2uXma3PqmR0nog9UCjI
7KyqcSB8pYff7a46QB9ivRv+twTnOQmrxvSH7o6kQ1eXFV0MHSFlg92K7UCgT7GM
lgO7O6piF8I26Ih2nlwD9Co3gpGjIO4lj+XmATtrziYI38U/hkowBlCMN9NaxZAj
9Po3E5ttOQAEZcWlL2wtlQhcQcFSlUEPmestt391RUpMsm+eGwIGpWUBlfXBYJuQ
t/o86M0+/iJgBOPYQethSL/niSBEpLwQONsbX+Yrf2/YKp1lauDaQPDvpRhn7DFP
6jx25Y1ayZDbfcMlwu4ZREBJ+GJvJEaIVFEqLFfb4eLhHCN0JcTPaNdvSSQz1fEe
iry27pIqO6qA1ptlSgmKjYx7I9XpSyNLyDaazyDAotQy3ikar5/te6nMzrF8Qujo
46cxaalJithv8WmB4mRtcDBmAowaM2a+LbxRwhVAGn1KfhhA2m9OD7E1JZ281t4w
gCTe0O4QgK9NXPDakCgfPmTOsTIcyiSXSRlaDyIQokn6Wjc/HlMsMh/a3bi2PZIK
QBYYHax16s+835wljA0KE6Lq3wdOUoq9Dpqw/iO6PfuY07ei7E7HmvXbcq25CWPa
Wxof5GSOH9Fufv3CpqjNmwET6Bc17tNXwFek3j0erv05Kj7fXHGDpo/X7b6FUasW
jYWQwb5bAOM4omFrxyLJ3gcSaDxVCFHBbHqzHl+05wlcTyNWym0T+0oUPOhc0Qdh
8PbYkxZxA/G38TwJXYHyeZ5slXEzu8Fam7i5YvLfjkDajsJKTT+lnCWQz59xy2ww
NKXL3PlKbpv+VLakewoBi/Z6dIyDQ9wlGSRV/+39B858nDfo5N1NxDwUptaq6Yrj
JB6zhDxs4QUPYQzZPS7QA7Dxp2DIWbzjl/kCVGp6KHxDHjUJf4zSKY96GZlmNA8k
+oZJQfzEeJSWIbtddF8dKS06fYt2BPq5/edNNyNde44UP1R3bnbs1DCc4FR06ndL
4PG2hfCwxYe8+aNjM0JUFewB3O2L07ceZISYfZN5E2bCeV+aamCcgx/1rpg2/Dlo
0f0Ccl6Sx3pQM9DiE8SZgTms273/fJ1qUJs0n2pLtQTs7TLMzjxd6DSP2lU5NYML
26xFhR92lRXRRIpyH3PRzDcWnkZi0tzt3Mb+KkxFYa08GV9hGQxd7YiNz9U6BIcy
dFIGSH71LGvu5GbAdzgXjfI/Q/RXJpb8FKHgPfgGQ5gBCtqibHOxbJIQJ4gSh8VS
c8itibrtomSk+RiRPsAb0Iz+oG3//Z8tOSlfzspmSnDBqrvLqOCJrzVVAjuMInl9
gN2X3KL/R2s0o5HUvHwkVp4FPpuV4pZSEWE9Iu9y03GPoApVwRNVm80loV02vGn4
OTWHyZAsBYd9xUeHe7TN0rjMNMFObmUQ/LwDkHxeVk91BqrBEXXZAGVSDHhiD7Kt
PLeg6du28UZ1jnvJPzs75boWyZ9l26MFyTyJtfHXEtDJl+9if7UaUWVuI/4y0V2Q
qJSaz362NuEPRzq1tIZKVtNmmbLwgiF25zsGEKBSitRqcIDIFmtF0tQfYgm6drXA
bJSVYA8sz7/+vO1zIy4DgQ7RMGT8CF2RPQygKcgp47k/g8FRr5OBy3bFYLf+2BAc
LERIqDYoweKCxlUFBloCLZHYYzNShwk4p35ORyubui27YJku0DFEUIvhuByiyHw9
dGJY65ZbMMrw8bz/lqrgZnpwSxajjYd02ny2l4S2yVDelAeS2a7cmGU7D/g8x3xb
N3rIjCcLRypSyUMc4HVCmICbKnJ1zj+QGbx8Iy+EWIrJpmrpNLQob5OJ6P/AL91/
ABvIzA2SHz9B8rEilU2wuas9zSTbNrUzmc2Hb8YivAm+3VKbPOddt+KdSyWfDb5p
MEocLV0yuIPlkazkuHhnLAWhMYEGj14FwaGugrjWBW3xgkRmX3o3JEokVdiQeXLt
ISXmapEA7/W9sIOd8rv16FSAjDj4ZgOEE2TUoiKBb5n2arO2lMMUzjtnacZQVdys
vvX6eWaDjCmT7362MnRpfyJlY2CL8V/rPgdo04pb8nWdnsKWOFe5AFBE43L2xVo6
ODLST3QOyAZy4qdMDy1bB5CSt9IfZeTXdD7g1y2pT7j4jeQiduQ0rSTpTNUlnCF5
af5iYBAp71JS2/mfsbVup71v3JUaFRdMWJEF7EzSfYl17mXYd8VwM+i0I/79xziG
DdKUCi2X5divaDhpYGcJ3haPNGBeYdpwDXbq5GmzftRsl54x01sKRjpUlfrcf9A9
JelBoh37WUTwUZwIMuDR7j8KYvMvhshduH7hlXJGJRRsHCxKJbN3q9YYhHZZOlWd
7V4517lrn5NxV8hBOMwzwVWF1P08EQWA8NYoGNZy/XKfoiG8RfMLi+kpMtwb8eQk
Tp05r7eb2ECoxKw7X/7fmvHzAIPBqY8TiHU2vA4P2spUsI+wsz/kTZN+Ti6b9Atf
ipArtpALUQOk8H5Lbf3Hkj84ednO77GYGrevlztfhyJfEmK7pYhzGlV1bc8iZDDa
dkkT3sjLBxEiUblDJsdlfXeRFL2IJaI4+9qCHiYXTx4v0h1No5hlCW7so9KmvZ85
H0gm4Hefl0pPFnlpbESPyrG9/r1q28FbdoYPqIaKMSBZIKxFQlSiVmaq2MGEzavC
sMz689hDt5ptIiouacw3tk+ts6j/Z4zu+eNuI715QviXD/ue1tC8JkfRsZko/iBZ
rxXCRYoPhJWHEc5tRfTYirpWds9tpH5Wvq18ZK7tx0Fwe+gq6mbgh951RyFPRXvS
0/C4Jc6w6BIZcA3QVSvNvvEcmBcsWFN3jY8/fVeNV2x+9asmemLJ8L9pZzYOA2Nx
W728wDo2Zt68SqVsQhaE7XzYnn9ArmkrJftYz6QkIXjp1Z79JjnKkOAn9AmRLehU
UWmk9r7PhalN6/U8z9ICbwUIh4Lw5S+H+buzTP6b1mavXTGtDO7Fgj1pXkqyXymU
Hvn/D8T/TU3DjKA1BVz+19y7jvRWPi7sw8XIWW0Ymmj9K8JKuXcWItHpvpC+Je6m
F0zP0DZ5CXiZJl2Mew/s3CRTwfpyJiN1OKmnfZ/TYsvK7up6OUtapgRkTYOP9fK6
6qAAmURbFNNEsRzZm5V/eULMNNOqexiEGW99Bgdgfz6EQezNnFbzlXsciVFgu/mV
N3km4U4/lJqOWmNSrBAhOHtWhODSsCB3IDHIVRqKgY621BocUWSwnVqaU5Xe6A55
Hk0tektN+igmMZ1IwcivHaI1iP2aIUbnR6XD6FknR0/IrrOHD8sdoa7QHoU5oH/H
zji2PGsC40mb9uEtxe5iPgo9GGrkFPDG/aRpD3/anlUMQzddnKjnBBiZGtyAb0EZ
ju41oIbZCXiecmYCkQHmf5lMNRJfD50CNMlDkzqKpDQNGqQ2sYHcRcWkDyK67ih+
gr1wdP0YX13d7ZVrq/sGcnTAFRgOASWbhSKAVhaaqojnydV2kBqcnn8i15nxCyyy
WHJ5dWsGIKXqUVXrickk+GEcPq7Yelr7oyHdRHjeRyc0M7RmNYpIeSNHB5S6UdDS
N1/0JCnJKPGYWHU2qbZzbmGZEihoes0mz3vLD/Doo8gZeYCHd9bdNhK4T5RLMIy4
arrwfrorOU+OgzUnvlZ9tQaQLxjvbLEnFBTu4rI4o99HxV/ydD0fe8f3wW5SS+Ze
2rr+MPreeFQ80nevsM15xNwFLlVQQHhSHE9DivDtnreoTx9q2LUz+3DGq209cJn5
+ugBbAZypUMFfQGqmcQRqJtDHuEQyYEcd6eZ6KovV/FjFrWmdAwGsdpHqDm4LBok
Kfsb+24aqzhS3CPegBQLj8xH6c8trG/KZp7QpdlSrMtW8GSm9ux4gXZYOO/S43ch
6dxItCYO/StrbqLpGaRyLHr6gxpd5awJjmBckx1ZQE2omwKavofi2ps4+gC9HoSt
qvJsYp+yL66iH1WWzzkC49iPEJLcDRsbwQM8qIFG6uq9/VbAkqFPga3Bqe3fGKQq
NoWY7QizxzjTX4glImlhpoRmIJr2vXAVhN6f6q0eLCwU/ECwFFWFRxtJfxZ2AeN4
caohAJlMTYQQ7FPMPF5/nNVFzayTbvGXXUAOGWp1d/Tr/7CK4AXrrFqeh34HN76v
B+k5N+xdLh22JuPfNb5jSDlNwevJBp/v4Re21xxnbEL9SnY+u3LpMX3nZYZWRkuy
WnNIchq5KqdXaqJZsdKvzKrD5rIqt0CUwS4zvk5qbz0O0TslkGRp1BOt+bpGrUiB
1jlFyxrkgZAW+PFeZIKBnavAQadrxk2koFVPnoP6SiApSvU70RL7ajZzD6lRU8Dv
QOehm1DEnjEG3TMBGhthZAwJ4gYlnKeGhlt7MXHz/0NgbcX+A878n544Sjd+8hF+
djqTbgJLThfMVsG6ZEe42BOHZsC4/0zK8ONzYIdntVOVf/Zoz/2/Yb+GNEAlyNYz
7OCgdgT6KzeAJyB8GELlMq6tZtXugTvSj5VLfMuQf8yJcMuINlIptWLmEDYJHoVV
rNKHJ7yOyY0h3afOf+rHZ5rElOtbGYaZPECUNBKLjZHizE/2EGXza/sKu55lQxR6
/cWUUpi5UHPiCZ0x4T/thPvkPtSxDxPZ2a3+DilBk0Dc4fzH1nKDVinwy0TXU9n3
LfGzWEC7skwds1zABo0PaF233K7UZ9I9ziZNURxF1j1fiOVU/HvBgFTS0TETknUM
D6jTiVr2CDeFclqpeUO2HjYw4iVmwseVIDjMBPqbwv7Z/c+rjD1vHtumBiOAc7A7
k5KEqac3d36+5ejCoqW4Q58M0tES0cxXNStxLd8aOBrN/qI5d/OpDi7FZedFQhPX
nxWfAn7JYt2HjWEjZ0jGQ5qfIFhZrr90Xw2iGij0OlxPha+dBqL2E6Po0fdLB7no
C74JudLaqT8JezT3LarB3c/+TNTcYl+nVnWj3ZCSyWF6fA0TvprMHC1X6GtKyIML
phlLO4a5xX9ZxrEVqfFIdGs1c6dnOCH6qHmj+kzif/O74n2yBUMSoWLMWBk1L3cU
lkKmVKk0OR4tyYcFlvkqhAJOZl/qEZyhFt46mC1TZliXhOE3qOfaRYsb54KzaO6j
lHQHMpQOeIQDQWSFmaMvJPG9aUEkjreHPd+waPDyxSF61zKO0EhHZoktAoCi4oWI
rawQcSOt/6/6sFYBPBbD7CYJEjUwNjxdYEeE2oYWvJe7mx5RnVLgVvNjmTuk2d8c
NjFO/of0wpE23vhqJv80pkgHZuzYqCWyqOj8RQfJBUf2uWS3/5ASpNa0e1WaqL9e
OxGxHrh3K7MuP9arzMkvakoH+FW4vSwkX3Wh0LYLZ3hHZbhRDnTbSficPrW+lxVa
7oQuJhGZ/F9j087F58PFLxnCFte6/SFdRTPQfRxHwntxDjg5jrw4s3LUrgO5UQTn
zl/sjo85D8X9EzL+/lWoecMn6Livm//sjJhLc79Q7omvVymQ0XTBS76xMOv0nvNj
e4Ryh6rxB/2xozPSZsG+77NgMh6mIIHxss66ucQ6gw4CeXvAqAs3hd0kg/IjBuFJ
exgGDW/mF6AkR+Cd13HcFDcOI8oFD8fZj9L9oWuvedlFjx2JpgGVs8HY23wr5bSH
1EBpBiK6d0r8M/txgIkpAB2vmaC9mWK55xOD8hrI3FItpVMMwT3Wb8YWvvDhEH7V
esFZmRiiqOzhRwQK/UdSEifF35IXMxFWxJWYBGGFoStyDA369Uh4MCbP8mcBhSHR
myTldNC9ND9spIbrirPkSsXvFK6tj12gQZZHEYLJ/8Ckv8nVFODUzIbDSH0MOHLB
TKmzmiOc5qjXN/KAD5o87ld3M7WHxbWf/jF15istRJN3SHVGpgUw8I6S5iT1FhmX
ULUHaBzBhyW606z4VeWnOi3nCdBDwfJIoL8aEsItn9V0GB4UBOMG2kx96/qVwzJN
mACOzhgio2KrhaG4zQZuLs8nQTiu2YYvng9BIg8o7anZULYURkwQ2c8dfObA4XSi
p12RjunARB1pHrpzBAXgplc9Ma/Sfw+8g2wZkez3X0RE6W3Q5s3z/UuGO1MzNzBu
aEA6SWd2mEa1e9k5GWuJmvcox3wc7ftm8tEG+V2hPgb3DXN22q78OHmzY7qRRXMo
+sDcKOg7lMRqTIFWZpkalhL4UUEsRV1i4HHYaKfU6wVI6PXUdsg+LSkM4+IPj2fK
bHnk4pplu0c1oUJYkWWCUWA7rH5IZDQqPk1N3N8k/SLmhOsf4rkVuVDQAvTJbuEz
ndRtzIhIZrrmA+1KdtyZXSVfyG55Cfcqt7CYMDOxLD9pIEhJgrZAZj2gZOec4hHt
VYEhA7fwgvFNsApQuASUJPt4P98iUmg49xCPMm9ub/VqjQtzian3/TYz/nE8DhLb
zcNx+GaH+gTn74q2/g5zC+B9PgaKctBaDrq67LxVaf0OhMxyNz+nx8Pdr6I0Fzpm
/FNCRY3YaEex3D/DPLgXsFWx5cGh5eF8mkUfcTyriSl4XCOL1FVqJO+LUIRSERsz
/xaKFJN7CCLfzeaFgRPJ9CVHnpoaVv6hsJl82Jv90xBRmcA2agWZum+MGXRVsr3a
cSrtRSkYmTZETQnd8pA+y9wCgsZLCKJ9PV2jnLAmkYlxTlZSeWe2AJVX3QQTnnd8
LL1skeOKZDcf+uEdAU9T18ESlHDt69MDOiR+j0vcwwmpAE2cRvYKDsDqCPDo3JMR
RqZ8FfwY5FKFZTJZSO7Sw9L3qOZw59YdlQHpYGEsN4HnGIbABez+wNYpVjPjwe93
l5j2+UbKakHoKfwtKSsMFOsFaplkc/5p5uAHsU9FDMi+7NkQvTCSf5bcMQM58aHn
OTxsfkapk8krNirB9IJXlVLDvt+ToYz7nKu8dQFO8uReER8IXhuUkoiWDRtCh2Ig
TYD3jRCE9LupVmVBU+rJLE1cRKCGOvmfjNGDnjzpnpOnmNgtye1o2BBb9qUFxMoB
SnU0U4m8I5haBThv/gJ9bE6wG5gJiEaW8Vr9MqZuWwA5DI3vAGz9Kna4mzCBN/Zo
HdekpF/SIXvAmSqvrj3BHbHKujfPOD5CsZJk5HC76QeSaht539vdj7N/A/NGlv+C
+0SvS2U3qjn6A9zf1gnKalTJcnGhETZr8A6kuT332Z4rb78zJKVzkQ/ddi3bccTs
bW/fIMPncOiDnl32SDbAL3kJU4nxoIxLJ7SN56hfR+aFZfTEAv1RlbtYJhtbqSGl
UtCase0LXTHfSXT6+B2n7ku6wzLQsHzIMqlsycAJEA0QzE9XUl6xg4dTbc696Vpz
0LDPVXpK6TYc+21wdhJR0U89lYWh/4k3s39igJrJ8h8+xttMl+F9Q5qRYsQJu1rn
8Idk8MpztQEHbamhKIK8ZotPi6QChLTyBeHNVE1//erJi5Nuw8EQpcKP0iaL8uYs
YxzDZNEc7gk+JU3HwlGGL9tHmsW427TmR0MopqzbH7VMVtSRwN6QQHRy/MYj+576
GVPDfAI1ByPqHxsBJjFUup9iGSPzI7KdZhGoK8EDutPVSkTQf7l51KHx0WqUcHto
Qt756L9RZKkWrq1kJd1OuAAc+vZptAQKaC+6QH9324NJnftlmrnyj5T7PjLQ2JTP
zp3/s+zU8aqnMqK8YRBuaBl5B+xq4KpVcSfW6ShBAUQ2RIMZ2CJDyqIwvQDqvU7D
/ZDu4yYpNfrjcvyIyCihvAZWDGhd+XCjY94S9QZcDK7zuQ82pBPDU9zoxU6LgtXE
FcpHvfwzlG3vyWUsiPKCHfx3Ix+WAX2x3fgFEVyXUUY6IlW89nUklWslRBxpMWDk
Xzn8QslqBoUe+tHZSdQbCmNivA05oExIkONnv52CwGh8Go4LzYpglE9MgXa72Q12
ElT8B9Rz8WENDWHbaFOHr/7ovPdql96VW1gR83pp6JV6Imc1ClXMjK9PpFH4GCCB
9sj3oMn5xvdkUzWlqS506sC92HSlNdKUPqf8v6CXY+9BPLO1AqlY7sJM1kuP2rHU
D4OqY95JE+CPeOudf1R8el62XM98zyGReEDCNd6xkC77LUQybwJI3K0evcbcB1GU
pJNM3eUljKSIGwGKUR0yMnW1xJZGZ+RSc2fziG8rAt31NF980qWWD03ClCHHokCx
cXTRp7HaqPNKwbZ4HPvfTKoilEfpLDEtZTvkI9nXgKsYLMxy5a/oa7jkHa9MZNgn
GT3aodPoKiE7UaIFTj1XZ8ELPVfapfq2mkWqD1bRKKJM79g9d/n2Bb7lchI8Fqc8
1VI2kf50Lri+Dyq9yEUoP0dbqpRLa1fCcqDggtgRwdLpsWPh0rPN8Tprw5DtOs9C
Ogaa3UZMSdOJtIDlnfTIkRBto9y1xclXY93bewVwAjRI/AjLOwrXCvCI/ToSBRpz
4h8L3OekSTldZKF07Etmim0Wg9EdrsVwmkb+iJZma1aAi3KoYbceOPisTCtgoPtY
SdpHl6180DFmsjvMS291wmIT9+pF0pyTftEY85NW20+t9M7D1GIXhoBOHKhfI7kx
4ceyUFExkfJqDqHsAWtTd3+8f16iXKDX1oR1wgL5YeNwat2FlPcy0SwsctqSLu64
sIcEA5aVJq4H8Qq5S0dCKHSUyRB0C7VPDoM4Rf+yGwhpBxWuHstWQqWKmbc+EwEk
VYeqRxaWA3i1aXscePbSyfr+l2uuYk+nUazPvw/PUWkJyxZwutJByjfgBdDE4PIA
9dQ3M0nfZ7s/um1/i47N2i8WSFqx9QqqRyVUe99OyHK+71D77y6SzN1jmRB3Jbqo
eyX1oWfEmrODScD4yV0IL9p+VnIY79IhXnoXcbObl4sXJXuu0GAlz5upgSUcfY68
vUMURk2tFj7vK/Q0Jq8SGz1x8eCnXCLGkMniwAYIYNSXsFwPzDDBPPUI0kBJrIe+
hubRfkR0UcNMtB4Ym6MgwKz1FaCgXdWlnqUo/z4+8i0q7Ox5xLH4iUSuN6dKSO3x
J3GIiFryECNzLthxlOdyjECFeUKZ/qnzjOJA/1k/dgmSxDgITa/4LTf6asiFDsVL
ReX5Z29mJ473apQWD7mf7TgHRnjS6iUrIGKPIbDb7YgWQqeWsvuJ4VIa87YZomCy
1hlQi42fc4vxSs1lE/zq3ZJDkvG0wgYUOPvlnFe7ZaVi8K1mQjeaAuXAnaolyB+T
7/WlFYV5b+rKjMCkLd8t1itf8X4ZkN71BhKesXNabvhbnMGZv5ODDbfCfOkvPqQa
Lp4kPBj5lpXBsTdOL4w+fPlmnig5EtJ9drevuONcktGuByeJ/xNoC8SxIQ8uMMDb
yfVBwDAaIgzezHzIGGQJeHw3hAFBlciYLDzwZ//iQVlMd2sry7BqCXh1HcT3a2WD
EqsxD8sRogeSzVwRJQ95w1KBeN33FAeTJMJJ2p7X3twVXfqQSToxI03nQaI0mM98
ZUKBtk1diqtrdZKIMJscMbt0PFOPdEyFx5ccXafBJhtnBsc8KiTlwLXtcIHfcAJg
hTfqmuVWp2K/tLbgNKfRGs3KvywMHWWEuCJf0RvEodX6fKRmo5S5lG9EXVvxdlHx
O2n1XkCpd/CITUDmel9gH8PjHB+p8EVVNT+GIPt4hbAnN+cbv8fVlFl7O0O3Tt9R
V8SEdOEZol8G/LFO1yzFfO3FhiP0MExUBtNuBxIsILd7Pcqa6EfBxngwjoCxWHH7
CeHDpZ20fisVlNONXDg7g79Y0/YPQ55EgHyoLtOz7osDZWpZhYmANWx6LqcVrvkC
ohrKPXe6BEbZ8EYTZ6vXNa7IXAJsLRANuvN1Q/K1sLKZLuoteUHPq9DG+nLYpA8g
xCh/UHx9L50bevkFT8rvwhB4h9LI/jywYmwLh790L3OuUnl6Zcp+9rMbQCi/v4ck
i6frL4MZ/4eIwsBsw/kD8igptnIb6uuWsVsuFyE/TJFMJqSbj3PWzIL1lUoqSF+D
pzGFMvhyXzYU351n1dfcPiz8BLL1aWTBA0pbuU9lNyM9uTBQXXE2SGtmHyWzuWig
8yETraYhyzIgCPHQMUfXxotxr9zmqL9YTRvHzkS/NHfZmP9PxsdHeQbiaGV5Fwux
iaCWuj5ZITFhk62IrppZq/YA/kUfPLilOmw6PdSHq0binajSjGxsAT7Dm3kIicbB
sWiVegk7vw3Hv1o7+tTRljBcx9lVn2QP64o9wTcHbh469V5+7hk70e7ufa75G2WZ
XUtARaVRsNJF+up3R1YgnfW86TsMfqViU252YfFfltrRqteWr5m+wiuyW73T/toH
rdgkaLDL0oSd39UHrxqU7iK3C3yev4PE4PAHYTvcrTwFJCLra9nCghObhMyDeQGW
KGldKue0R7YLqBoIHm2o1E013GxLjDN/lJTJpiA9cW3VldWNFFEBH76+xXOgnzi4
e9t9W0k7VJySobsutpWp+C3iELuxOnbBeMllQd0oXRx9+QBGR7VqQLlTrOKHaaXZ
C+xIy/45//+BurtMzoYMLS7oVqj/HJseyzFd1H80RpEVlX4TwsxIwX8d4XGqqBEa
7j45H3JERNJsrvQsl6+MjczEOOPjDcYF1Nv4B63vm6Z/DnctCNW1eUQvL+pta1uh
mzxgKA5Q8eVMhqDHYoGKdFjj92s0QvkNrYNJYlCDA4Xt2JdSPRoyzyFdJ9dsha6C
gEtCrhijKpAI0Jw+dar+gE+Bz9Wl/OAfgWsu9TzEN7EwyBCz1HdQF9br+La4LXYG
Q7MitfTnfN+m/NVRkYvNJZkrnec3aHa54Z5XQOvvuMoXEy+aBrF2+L6bGumW92T+
VfpytcmtKx0fJYnXViZF7agM1v3zCXIZAoHzorGCO/+KUU9cEZUjXNs49XhyupbU
yUwkVEXQnpUSBoYI+cP+I8E5j5Mj/j22+Sv2sQLWcO+NX93hh/a6OZ0uu3vsNkTx
Q3Y1+PmJ5B/FmTPOZbBnKMp0KPTtiu37ykyLCHJf1Bu/oSFepYzG3chLzPdd4q5H
3ymd3GPDfpBvJJiPZhkTx5ziGUaVcEY83U4xL2yVjL3iJyrYi3EXbd/ZPFe4d8hV
UQ57CkEPIUwWEL1Zop8WXOgStcgqyNALdIUjwSu4nHwMbhLlXIidZFP53n0clzBH
MFXAWxnNWLo/uO84YLz/qaqj13RdKzaKAQjkM3Bw9B/2Bxuv/3YCq6tuO7KQqMqF
04NS2TxM2dkZfYolaGnZWOToTi31A5cI7Cbztd6fD9w+F03TA6cpYQjt6uRygzFt
I7qsWiRhRovDasInoaw5nlJLmDWdCAkAft/pYj7tP871rtQeDn9LE6LPnirR2L26
Q0G72cBggZPh95KixH7Y+OdGgTl9hSluDPRldfFeEwnZuSm6oOaA5g2qJ1XT41R/
M7NBKIWzhuJPwZYI75+V9RFHyXKbUKFU6P6hrxqI0wlxp1WUqHyZri1F56NZMvIv
e2XVc8cLpLrQ5vJYHCT6ODYDRCLMS+Fl2FkOz8ZyVY+39oPgdxWOtbfi0yUcXY+C
5nKmIU1gOs4piG8e63e6dZ8dIl8y9YzPpyQkKh2SI8qFdozLhHldgk8CZ1PtoJZL
ddxWEwg0qFxW7p442O5xEEVlqLlH9vEWDeulw5oNUFujHlMauUqeqKdMnLHGmhhp
03zXkkTin+rgbaTW59+N2/odX+8HEjsBpTwZ1sS/sjSy4gTqBBrJRn19k0p+078U
NlJoNvUjibps5uU+kv84kWJrjRencjoTWgQ/oObdX9ZxPZ8Uy6qsqHmVDX9mhpoG
5uNJubobz7M6gbkQkEPf4Ir7MFxk/O8CuW1pnrSQuRFhSoPLS6OpBS+DwKczWwvH
qbgvGJibv69tEjKEKbRqQtQli0elIprJoc4JBIwOYncZ2txKUgjm7UoXklpu2x8T
YEoZfV2Lljaz6I113AwggBRRnmsRtg8Rke+B/jh/3lp87I5y/zMPL4yaM8tUrGvk
+tERPERP+gupIGI3iJlGFTvTvLDpUq9b0SATFX2ax8xcWf2NMvpO/jAcb68yZSve
SpJp4J3orJr9iocPkz6OQo1Ye7QPFrJNOr1R8RwIMDYqjWKDG/h/aRvb/eFI/kR+
LhHpgkipCYuyBX/8ADxj414Ucu8lB0c8s0cxihyLa9Vw2mR3y4wiStnNp1FNi5Ia
c/PzGCDwoUm1scYkio+pgWcWFddwx08EnAtg76XyLj9vAVQ/xWlTSNGdwDpOeQ69
zgXxw3CHXmE1Jp1SRzdNGtE/wOxPMuJBURHUAqZpufQpdXH1izSvP0aFZ+n9KgLt
7ACnWM/K/XlH8InGYeZN6/Vs/BmSiGwj6p/EmHr37Z4QiVTOVwhuAy4EDD5HOo82
ta0+1VknF6xp9REy0RCD3Bh2FjfzCS8Ryk/5xkV3dkx1K2NdP5Mkgwv5vgl1OKRH
RAEWnXL5gqIZNRMwI5/Cm6iVDIO8ArevlL5Eu0DiObxpMFtaos5zXDLjiBLffM7i
aQLzp5lydTcoqh6PmF4M7Y13tXfgXTBFeK8OKa47VgOkImjWfXYj37LYtJ2SYnYe
Sd+2vj79QvQYj3bnF8u3DspiJi0zUcGCSnNbj0m5IWSUWEregYtTm2sDN5Ue4Qjb
VnqDIUMrXcp65ABFLdjMls14tat2CgI5btpSpxXHNqbsqCm32yXsUKetKCBX5GgT
HgJe8XhYZJLJw12z9+NdbRwijG49EueY6G9fAjVa5OGfnatiADe1P6/5TsfhjCyd
Or+uu/L02PwPzR5GhAukLBX0mVfdxEFFHLkTRTS6upHVuzMT92upZ987dEglmcQz
DnAaVC3i0n3kHhUfF+VlbzgPNt7+whzs4u8Yl9eweDG9SHSN1tpSxCWK/NhIwzq6
3ZdbsIOh5FLe3tJdLaHoDSoHLHUG6jmCDTqdYMKCa8aZCBL1xceqdflYEBjo3OVT
8QcaBT6YEUl8lyfeZsObz51GCIOP/+v2aVWDb32pac2KxSg5d2kDd6NhPg5xFrE0
yj1bd1MV6GJ/66BnUs89dLoDRuskhtAZ7EOSpuYXVgdPGIwaCBlnpoDAFn1/exT0
oAUyMmM2cdhSCQaZIffH/+iJC01Rb5tf5Dvv0lBATtxyWp8u23Vm7iA+dTPJGOnO
Yt0dejJpEHPqAwdubEYdE2bCzfUVp/IrHpAeoN6fKq34CSfSb4berNoo5ccGgJFd
ADHEqIudOewtWeIVeLC6tBmDaaZPzC7NQwl8YhskjfosCEviXvg00mePCjpUild+
lYXFFnCOcAKMx5XRrBcH6SpNevaOpI4wZl5Xt57X7b5Rr7pDWzwmyL29DycrquyO
AbppAW+Gux9TUqlABTwF3UI00A3xw3hGHXyqq9nIchat/HcbDvsvUTW5Vof2n+L3
uVQwGgt++VRwp/cnekJq6lxbFAWht21ETAifbMOXKcEx2lNY2rGEDs5AJOHG5FKO
9Jmr3reR5CLTUtcZuITOd5ONWtNBo8aQlEmTxapXdzV2rbz43WijBMeuU7Xs8WrH
+z0YLjBhwiZLRPexTp4qSxRO1Nyj1XgAKltVJQrHopKzkEESPnh8kChT0kbFXF8i
FR4cD7vcVtm3mXmZCLhjcJ+srCPyxuxtUj/AYIh/KDjwkrdJA23yZJ7K/KBDczSP
eOXM2G36ZbXqd6/r7Rvf9fC3dw9bI1GoNerekQF0j2ShhFRE4+kXgNHsUu7RjrrM
mGSKKrAOhx3X919jlqoQZEoh/6sL5Lw9RIZSpT9RNwcyWR1/0g5Ugv2URt2MSI9x
KwLeKBfMrc/IABzM2I2oWLB4Yxrx4VEaNM+WeDXR7n7nQdSvelo/w96NFfhgQvAI
ak6MB2GEUrWKhuVtWNv7/2KIOIrRNfMOwrj7TLkGqp5f0HWqBQur5GmlhIuWVXIO
AUF2z0z6nrPhyMy6lYQuixvg0mNedebAQx8cb6ndpFjRT76XtsfS5hudk+dVgZuM
Rq/sRJYArBFmB1i0xdq6aAbo8nTYi+kXy60RhXC/UBIw2qfsZhwIgcp/xi2HXZg4
5SRdvd81te8ngGAJ+0ynCkpFvvpm8NrQvTDnwPM6UXuMKkxwNATJceLNmWGFCqhV
gfdImkF+b+O5s7XfYZSnt+K81sTgXPV1agxALj1oRqVYnj9LIu8iWll2qJZTWTwO
mGPaccXtV11cEDiBdH042J5MdmEnV6o152ozY7tCeRC9hQYdEpcXZBwDdq68NudL
MKqBgCrQLHiKFHY6empgjQ3xlwoHYXD5v/OqaQHveJMQw9gvnY0p8Ywl6NCGnDfs
dk0HqXFzVgncdmDvEbqrAGC7omZaQVSWuYf9qoCQfFssxyLNlWyQcGh2BFK8wXoR
3aq/4M0seOoq2rjZKugIkyu0HP+wXj/uPaGThmUM7LtARX5ZbJHkU13FO8sqUbAM
gvgxzAyls+s0pPfWyaQdoMteF/o+2pX4l4h2PLLKWc0lf9NHMaKu2wfATWnBJdrh
k3PgDEnaTJ8OfSppFT9mrTQrRDWVb+x2TLmAjR4SanVZZm0wNhoqSe0uK4kocLUg
usQDEBAf73b8SSndV+fJ1uppBKZU5p9yux0Z6CS2FPiEI+q3GuUWHv8wDpyheTTP
e+4syyXyuhoXhfl4cBWGF24ghopDJ2bCkL1v3SHbgXrEB/oBbkZTC2nHDU5ejzSq
PL8jbB8ozRlf1TCEuwVta60quOxGNt3BbJ/ApT+WyV6vzB0XW2u8Fiivv5KYoIOH
iznxWWY3Q2Vjs2xx0umIPnh5xI3ndKdyiAlC8R3ZljXppP7CUBsfrMKTc+xPcBlZ
L5kNRpSOOOZKZkBs15GLFYqRY08eIn9lstiDy6ft0smBVXctjxZgfpk9bCFhJHNs
zrOYXObt7Jzd1p2JzCJuQzIGBLCS+RQsoaoYVJX7//FZfuTsPwJBtQMm2SiYD0PY
vab+oxXCcUGkNE7Us6BBZ9EebwKVZOo2ZD/sNtOLIWiQDQDyXRy+q0B2GEnj1NWG
PcbjFjZUw73J4ueg6hOC8nLOkKNXDtkcl231NeyO9eoeKRrROIhZU1Y6AU3hUwP8
2UPUr6oI6lQgYebxei9ZNPS4OQ7XqV5sMH4GAxeUb9FwHODmcNugsrVRpzSc4Ohw
0VkdINrrCCqgT/6ctKVvnfUpbY2600vN3Semd3xcQ1Zgd6BkQhIb8IjLjMHyr/L8
cq7P2Vgt7tg/Of2n49V5bDaRdFna331LsK//llNPwJolqGT1H2IO4sO/jv00hpmO
WNPV+Htl3NXFtFN72ODZyuF21asWAuPhOmtM6lgXCUwEhIiLejW6FXOALj5KtxnE
xGD/tbgWGBQxDG75/fgXU+o1fnX+IExcSVaSSuDwIUEr8Sx3M/AekIrSBd6yloYJ
BaYBPj3m7MVDUNwqGvFnzx2qg4eU4aqUtEQQaCQqn26/7g+0lEF4ia1XxsAsaOFL
sWZ5xlnbPXdNowOU28TbbrwP4GTUmCtkJ66h9v1eCmLvo1EdobT+6TBMaovhwFXt
PnIwtIaHdAaD0hyF6YiVouZ9klH6ACiSX0vqyifOxzwfrSn8GwlQqCLCNZnBVXVu
CCQYURG+oWfuNhrWHVRuLD4cJDbo0Drm+X7PIL6fuOys1rTentTxLHNdnytd/Bmz
g1n75NarLoGfy3dXdYdq/ymV2OVY3hgCt8R8kuLnyU9bvLGRMxuF+tXDCvaGXsIG
DrszPVNmnGfXp+rHRzecmKWWWciR6gdA/2LaZ33R0dOYcP3K656+6r0eX5bC0o5D
oodBjLxatrdrKJBOkmxDMyX+8M8ov9mQ87RFmmhnKMzhPD5ke7ziizjDjgBtuB/g
oBoyT2wPGj3sBL/V5iU/1JTlWSIRmCru7U6YuR7PyG+lj9E/Xa1yKc7mLo8v7FIW
LG4Pj5jsorDP+dI9ykmH34vo7ik/FA5mlU0cl1i5NE1qF9U6CBp/pisZ72L3gLaS
2P/pgkZz8qlhQaEReFZPu+hR92CflZNkPOMxWsTPfubIRCv2PFmlTiM7QZT2wil2
xXPDrqQbx5CkcuhP1KizRRGP8jog9JZb3i9GL6NgB/iInfgQ7+PNNjXEVE2I8E+N
w3YBCgaHf/U6JPe9eDV+Ij9llugyZmfebgcC7iWG2Lucfw5X1ZgKA0hSsWOzrtu6
k/cwpsr6G4Toj0U649I8xc8bsfH7ry9c3ANJ3C/wbn+00CZSmEez5mhL52IU7P8n
SPfq7zOitWecHBbJgqYWRFBC0ej3Ny4wYBkU7Nb6I4CEPXZLtjf7Zo2RZcD6Wxtt
yWK2raFNIP81+K9LmYiKe6rV/Q3Ad74XAFtN48vhJdxx77yUNxyIDqUptp/Zgoyu
T7NJKlmzbExwHBlJ1UnDMq2dhDOar4d1NCSEr4WknXbaaUaFyNJdK6MUpPUsvUqJ
/2S8z3SukgD+1BbpIfjdBYOlVe22bC7rYfLALecSMMfTPDsa0oQ4vfFhgzXicWi3
z3/pcqtRWp2DmIFCtjcqitx1vzVqcN1PEt9mw0jOS3JQq7G8OEl/wm6X+J0irdM6
gY2n60D8riNzpzfs898M2LkpCnUsn3pihWxIjTj8uziwMOCnYfk2OIzQ/6P87+x2
OoHjDk5bTXe2q322QiqDhPbV7rTmApyJdqRAmXPX745hG+kLFbPmlvZTCgVoFREZ
ds7kenwRseh+I5SmjFnn+Z1eOVrRJSxHlTy7rlvP3pZWmOqiRg7FgUe3mTdo1HcI
x7cM931Kt/sD26Kfj+MnIhcnwgtSiIZbh6lEio6o2QCcqmeYeZVrSoX/Pr+yNahk
pXh98fVxcGQqXQVIreW4VhItArf3IYpxEX9Tc6sM4/tQU5SCWsIc8vHbDTwkFiVl
thG+XO6zePnZzCwQpd1WfDi6/wtD7HqMDLyAv0RD7x/nQnJM45MrEaU2cJRPiYto
8NUJkza3QSteRtzF0fbPvQRnXli6EKZo7SoCEnVUDMuU9VkkxM8GCUCvrAnkMHz8
djwGDdQZymbAm306GLthrhn9P4Ksk28Er6VKsojY7neOY0aHpz3J2ZnchMEsN4Ff
1FuA0yNryj1FCr3SMEKhnNqwSW68fdd6OezsrQlyDP+ifT1N53jCyoWEJQT5/Z/V
FnH3v8JB1hJQImTqPA0hCnSwnXf44727lFnt3uxsRloYFDiRFoZ2XOUqO3iZs2IE
kvwcJTPvBAw1KS1oc0H/Kw+SAApvT4A+ECgsSGaX3rv6bgjTlvzikA9ull8edmWr
bmwUgJnZheZRrXZc3hP0NqO0pUx2qV0DUNFNaHTNzOySU9hfBuRo00Hl0UYStLbb
d+6ChRRvpNJMoyjda5NmAlIUyiIqRJo72NlPjdqE6w3Vmc3pH+lIJYcfajKEQYT8
De0tMYtiJHqpfNelMQEaQYmL7PrYvVi9symW3Ky2Vvxn34mBQ6JRvbqklBM9r5yY
ov1C6Yc5HJrQ7aHWSqo6KhTHtBpFYZDgSUdxqKBzK2wg4yRX88eQa4ZnNdOInQIp
7ztcLNYbwyr+GK9kA8P8RKP1tMJ+cvm5bmdUeBYXx3zy7SHwIGc1HMnE3mqiiedJ
s2NO8ZH8Nat8B0shXpJF4EGtsCCtEGaef/1oZPkwLylee/ANzn6nau9n2hKrxkWO
BUS3YFOZv45ou496cQDpRAtoLkZSlO3EoVMCpfBGvnmELLepb69QCJEYq4+gxBun
vU1Ca5/KWJotX0azhvHFn2/j5/2letkBstGbNn1/8qH3mcUzJcIl7ZP7agIPI3S7
dSvnPf8/ql+w/bWF38nii3lkcQuxhQfS8jogIBwxD/YcawApYPDVsXHphE5ibsdC
mJJzftN+MKz3T0iVcYiqfHTr2G/5cht1Rr1SjgWvtcT9hkqZwX385JkC+cKmODwR
YQpn5zwoigKVYgtcy8W6+paEEY4lfm9BPhvC6j/D8EWLYk5eMI1SJppJzEocsGbX
gWaMY8dkqCFQOuiFYP3ruQ9BV0LGRtSXEkLzOBBSYbSJCxIUx78YTR7p/WYEJtRd
i/UbH9K3oE29IdEH8bkXXglyYK+OnuQkkK8Axbstdkv0dPlmdZ39uqmMRT3Gga2l
WJX/9rzziJ1idQoAnWRdEV84P+Ey6pjDcDKKTXPAa9rs+E0Y3SNXiinzeZsFl3L7
uFlc+sDiFIK1EPV41IEnM5bCN4dowQr4wonRNmLBlWO6tbfLX6Jl1GnaSp9gTeNJ
IaiT0GMHst/bBPrwKZkZaBHxwhqpcgSiVagYuF4P9GhgzU+Dol1JOP3nqYTQbMvk
a2KhmP/kZfpuhsEy6A8lJAUG4pZjj/zF+5n2CsEbpPtIMS1KLgjROjTdg9YCLbou
kid+O+bJ703hFAJ0NMP037PzaiMLX4vw9bspMKVf1drWyFHO17xy/pjIe/sCEfd2
R4pX7mSeNEiAcASj/XDDwIWvGO49PuT9CbVpKWlXPGpD3grrwcLfJHbReuU30AhG
P0f3EHwD8P7c2K51f/MNLyjJu05HvDdm7dUTe9xHke3NwbLUuj/+fR0BsSMiBVCa
RHOHWeLu2iclRIpcBCOIeXfNKeQZvOpxjtJXvIVm47xAGbs5ItQVDGv8koPY2lea
Yoyo8RvPoCMBecr6chVgKJ7YXNJmPU0s1sjUx397wV2Goxw4oTkZR6up2jei/6Ur
r33JBNcfameGEju+GxGzO5tFlKlA7NNH0H1sRvBkNjaK5Ycphdd+Wmy5x36OG/46
uL4M+wMZ2frM2qA0OngGg+6JMfoRFIhc997Xq4pZ7CjGbBs5+GAzrHZB6Us7qiU7
mG+xnlcanQ3dLrzRzoXt5gCAZFOUJf4Y2MucinYZ36N57U8q6YWs1+bUxY/V4QJg
gCzT3RbWgYQ+KjMnX6H+wchpCAhF7lyYu7kh8lHHH2M2820RfCa8xuVbeZqnxPYv
AdbOGUQawdQ3qYIbazMNM2TNemsQo8D6dzJR2u4uCLjcWawJ2P9u6ozIZAVp45OL
/ta5pxUDqAzt1dnHY5MQspM6jLepur07oDeUJYMxotgDytyquf/RSw8vhUBxE+Na
PspYQ3QDc9YNV0T7tbZewaaoeRdTcrX7CqarKntWXDdR9mi9DOKULgACWtUm7bBe
dHHXs2UtIG2x96DELeCllME+4+mPaMSWImwWl05198HytMh4LGXIs1OU8kbVPy+4
RD00IE1M3dfQQPMBgFrGZhLtmIovxq0sMIgUnkrbwtxDHi6yYKixnUsl2NVO+1uc
iRvHXh6lJVc3Jj9AJacGL9Ft92ioFFSoaM8tvRnDLnSlFgAn14tB65uGU2RA1wuJ
30kAsK8A/hUXsMk0/YcTGx9QaT8XDK/1PNFuiQaaj9wiKYJ7SMip7Br20v7MnkSa
jFrrVK3nioQ26TgA/oGqs2JnCc8GHs4IAo7bayg7nXUPHIETgjn6J/+EgmWZLx6K
uGLQJi9Tp/jITL3FndxMSoEk7LEwz9foPdhqMkQqcOYSf8y2ohPoJHmKPL4dSESe
zJzPj+HDXh4p/PQN/Q9jRL/RTTtlsa42J/k6ld1YQI+M0r+ibHssV6VBin/xFfzD
bda5mYR4kSLDTqeWdQEikjjUeYDaGwSJWJ/PbmDhpygvmtIm2sod7JYBirYvDd3t
+rewa5K7l1qRQ8hdvatH7cCI974p/M0Ov/50IQlBdnDy8p7DkD88czXWocdyJUmh
IZd9q3yNPPypknVaK/+TqULnxaMhEwAVt2UcAT2br0WRttHgz94Zj8K5DJ2m0Q9R
/nplqblxPqFIVVHibwwAsDbTrehmuGZcRv81TF/qkdYmt053fBNoCatDDgX1U407
IUAgEqDsS5dmqWpxZLbvVes8SsDS6NK3E7yE1p7PXnW5LtwvYt6zCQsaTqwowgwu
aQmOI4+hRTjdtqYqEYQhZ413poXDXZBU9f+xNcpVn3WAb5B2u62Ccs/eqeW68Tiz
SqIfviufbda9UVSKmDmDa7C7VfTqdLTyI9zI/B/6vLUCq0GAeNh9wvTmkIPnefe/
NJZnlfIXzXllU0GGAjnhb2yT99gPdAaOW40T1fSKyxu5wFh2Vl0nsd8+zpraiopM
paNG3GeHLk4tuXSbH6Ea6M36oiyIbj/q3h/L40/qCH28qcsBnc3tG5edKlsHnx5u
8A5GFyF5EgRZwiUOZtZhMn2nc0qSV0O/uA9oEYPitcrdz9FCSAfvuvlLI+Dgxq4u
VoPssb5Uu8gRjhRGpSRK+3RkIka6fPLDN0gLpHGu9l99veLS5i1s6qYNd5fYJr1D
23lEJdr4eCESzPSKDjp051imsR56pnx5IoC7/BybJBlrAyf5Hq7ZYPeHMsM+o64t
sb8pN3k5Q2lOIxmohP4sSyH+tvFwqzuX+fZgQvg6zHALKWKs/TWfrUxaxiuR+p3Z
eFxlqL1Ju6eXGntKelufsNUyYdm9DNHKRbsns15DPjuUUFpPrRfJA1EVmUKGmSi3
fUc6UUVekGHIKmCLM55j0pDgdva01Z2GI7Jd/nXLblpmN3DVyDdE44YY4TiweLLA
iHNnubFggWM/YA8xSSWCyYzHoaNGSvuwWy0pVhNDJI03TaGDRxA/PrgNki6V3z8m
vQJZZqiGkOcm2XqCWpC19Ax0R6wlOZuyDNXw1OG9Ahx2Rvl7MGxr2Sjoo6dQmMXx
8TAlA1EOi+bfhhb0V6+oGWvN4O57Xl/NOzKDERhvf5k0YD+Dz6QEN9lCrCUIVmML
+3wTCqgg9WmGeDDir8WV2E1kKDvR59ciqyf76/gaPtXJLIvHb2+ureeiRHrdE+Gz
DPzab09qPc54DdZTTQsGNTH+/C2vrp/VP8nn51unNMDMMuy06wSYHU3luOWw1nn2
7MqIAw3jl4hr0fsRh4jj5u9pIKBnKMCxZbMc7qgArlDd4h4ewQ1hyMHh8RAIA8se
t85UPUvJqIgUgKJIzQjiav/9Zbt3hf7g3OEsNOQ74kf9dE0JC5fw2Kz5BQBqHeHO
U1Ym/aWbOPSto1ukewXprXez9JiQIGha4QA+2RDqPeMJr/hQOuiWbws33uuJlaSs
+MMhsUhzXCg6qkJTNN4K/9a8oO0OtarsjjR6s8RTv2HM08emYWBIjzDLHgBLeGRR
XiBoP6ZM74ymDMW6uk+LsLyQn4Ri5rORssw0rOuGx/rv7JIED1VZ2uZyBQSnPNQ7
sYmtpFbPGE/QubLax2fD3g2GLVD1IygwhROfX302uE2yoKyR9duP+ZWm3x8EpGZq
Vq03CTWEYHQa/7ZS5I2l69Go8MTxw0044Z4puPJkupzKX3JaIidYlqLxZ+/Xqgbo
yf93D+KNA6v1wn6wjqjR3bYKgbRWISF7nS5dvHTyAC4EbXadlkqmmFhtJkzwIgtq
PdI4EMVAyH3Z8nyVVRSyaK6Q70mDqktxj0VnYP/aYJMs0b35EyVW+wMNvZvrn6GY
f6/x+zTcwzo4Y7icIM22OGDQvxkq5LmyXCytKx62Uisw1IXJjLC9NuIkjEYXPk/T
piVOXnaAId1fUOS+xoPjyTBN1zQ8A+H4J3Nyk1nY1Z8s+YyRCxu/jTiCA7eGRv8D
ZvMeacozRraISKhHNA9CR9CKwyxQcSpwvINHy2zNWKJMtEUKGgI3l/lGYh4hyC7N
docR+0jTxQsbZhhB9Sce76f5jPgGJ5K1EdEHAYghvWQoz7E8sAx9bjO/XWNkZvDJ
S0mOdm+CyEgA5tivWUtTylTIMmGG6PR/jbA404BG4tRuaLC/adPxKVm930Oi8l73
b5sRA0ZbFxbC+N5ZNZ6ibpQQPQDmC68mc98HJbe+JmG2SKopjMNk9eb5Ol2f7bIk
dExjSd4r6/IL3zWrMLyxEqWmsHDOKXv3qsrXToaBD2dFifoDzhwtpQe/p6pTYvmR
lYypRB3B8K7zEO001A5DLU4ivt1NAlpYEflseyj/S3jcwMU8onqhMbhgGm5EClee
3/l6k/wl7RAQLNhzvgjWboKLnwRvu/qCYMflONEtZJvkYG/qnk7yAI9jz6FAyejK
h8h+1KfAQIzIXnog/KfS94bhwUo2TmSK6P79TdgX9neKps8aO/w40gGmQYL+RXtj
1rxOXIUt5RvZ7WqrKDDc1PM5Ny3zU4TiOKTQ/zPmSo9XxLee7kMWZs3OyQSKptjo
oPC3Jy7BsP2LwV8UVdz4aA4ETuB9Uc3DU1SEeTqAYDBOI+K6wYqE8K9T9GbFb2N3
VNuC9z5by3B4xbojyJssERBUp/PT15yNieqArDtGN9+4SMIyzK55qGaaLVQY7T6S
zJwkMhhjiPY0W0PnZGWeOXOOiugHRkqA59edaeYkIGB3Kw8r0WEOi/XR4XT5fIku
ykNmxuA66iyrSChSMfOUg+ChTBJ/wRrvdtJBz/awOL0nJ9RQWA668NazKutlT8tj
cG8/zyo8PNqqE7J1EruKHHuZgCF9MOHMvs+GQW/sSBWmbf86gGqgk+ntfG0c88rs
0UIaoPngX3CF43U7pbsnCmtfg28ahu5eQUH4vRvSdoPopHdw0JBUtpoMEPwMRLTf
uT0eiHoCFFazqedXnlv0FpMHWcDyuUkTEmxaBy0Eewr8VFk7n/dvztxArb2FRqCg
OjN+wood3/0/Z3xo7vOfIQSRGISIrb8sRz6PALAAIsIjCjlLjAooXFIzFxhVH7ra
A90Y4hajTIbd3+twpM3dWD8O/ovsIBk43M3T9l/futvH9uG0encd70GQABSTOufk
7pyHvQJNJUPudqU6EgRg2rx7xJDlndNfUtqJ3sq7t9kXVOLGwAK5prwxwncYwgwn
6WtSBp4xUZ9wswhDI1oHSfhoNYLmbPme/8DpswlSar4qeTaodwP+T1b/BPzBUI/G
MFdmssW1jjqxC8s8UBSsskDbj9lw8Wj1iABl1We1fdp0h0WzT+H6MeJEevfNsV+4
qOfXsxsnEYko3qvT1fCD4XgICvWKgBlUKBeu76KBHM4VjSUY7vAUSYLaPekwbJTg
anL2Zidk5FikD0kxJ9cvdtE1YHwYPq/b2SnFVpsqCJ162qN+dsfWXuSaK24oQZBQ
tNUjVaK7DYQXwU2UkqRphfQwxYdWUGpr/SY3KFs3sIK8wEibvnhicqNLvZCHSz4K
tpMhSt3US7byk9rdTJX/ezpJkOu2c50WxKt4hyAptxIYKbFJCvD/k84cdjVfzTxN
eV67cIVZC82CO95+NKq9ZUFcs/K/9XjRP4sbi3qM2+CQk+1dZ8/QTjlY+4wCa5/Y
5ZBnP6P52qNO4NtfgKn8Ltln05HDO2K7QYU8Bwxdt0jRAlwBtkSkK/6gxHGy5vMj
0ISZGIn1e+FwWJN8U9zN8SRtGyLrDxoWXPw56P0k3rlyOD7g9P3AZH2SN8dSILEQ
tUuEB5UsZA7RBXWhAavfkwG8KkOIN56h8FS1tavbjmYqEwd2doibuQqHXnKsfuSB
OBBDiT1nwvNqXqnomVmzE39uJcyFSJplEKtZpmGvNm2RnaB9vERUJ5Sd5vyy7fyN
A3l4J1oIPRLnmNyHoV0JQckvEQdNsYTKja4OFhYabl4kj3WTiXbA9rYL5j+Nk2Oj
Pqr8Dih2MK/3qFDLIj0tulL9xNwRz3QJuKl0qqJW6zGg/L5C04bgSnY2tY9vwk5A
kz+V+9xUUHtegk/jzuTtyXW/HfWaB2Lz1ETJWqrHKCvFbVJKNJq8+o42ZSq41uU/
hab+e70KuULtL9dBSSZ5iUwrHqy/paZb08KBouSg1SppD+6iZvufeJZEtNDgiW65
ZeTWo/QSdD/OuoUlCXBzC0sKYE2xzNI63tpIAUx1GxtKRSipybGhr5N2U5ywOO6Q
RAerrQ8pSNJo3kbBZNCTu5l7WNjjOEPMFCU9PzzTjTDtKh5Q13Vq/S52kfqSUufB
6bgzOAzM5K2/fZJwb48LMTF34OXGnYcIj9TPwVZmEGBdV3BufWeB4PDI27FQKSa0
sWPsEUPIZxcDhkB0vgFM+e9yq24pXv6CveMrfQ950D5L3WtPKbzaaIu67pG6UMKJ
GXtB88VUXEBihAhZIqPpvfJgNVoqIETyeu/kMwkK5LPOROcoYqDLHNiUXiXHkyH2
y6RfXpdcFjelpWkdQnMjgtKJn9Kq+PLNUEtMvSFBFiG/gBJcky/aKPkyrtMLvBPY
f4rbW7e675gIMylub7EfJNIx9GyjYe1Drs5uAMa1thOZ5BUZFiUOE43waz1wjVlq
sMVbKHcQc9X6aW+vek4vGP/myRpyPfllchqzBQR0dHB8EwKkDAoN+jPq4aT/g+Tv
+KqnTCNyLeszZpFx9Daif3jmJbmB3msB2rKm2/ewnbntLK1rzMAyd+vOuZoIjzVp
tcw51hjmDTkdeKNYXhzrawp6FknfvxxPn6bphB0obN5gdjlbkd6CYzhEC3PgltN9
UBaKv8WkIj7vdSgjHqDWH4qnqeLUYG4Paucb+rn8C4S3mOggZxKst3WxGSjEfbCV
Mz0kdsVWiY+cJJkSd9aFirNmP+kGb2KsGeU7QBL+stxG1p9dGEqS7Ffc2HrBJazg
IO0tobGOom0FybGWbOwscs7r+W6Iml8YT02kY9VP47x4KRRfVEle6DEU7MQiFfPd
frfa4zEjS+wJ5TqgKobaNK5wq3MxRM74wMiUOYv55GcvQw+O87rMPCgWfcRJSeXI
8vpS7wJjTnqP30DiYLqRlzuP/59/fMCZwNeS4XuBaVtP3hyCbX0r0PNlgv1N2kFq
254oDMV7BYWne+he71gg3PfSDcsxDzHOb4Q3PqouD1Jw3Sf3CRci4biNi6GQNodE
W/qBRyevHp3cZtq+QFWflNQ4MsRE1at9CWjobo6wwvLwSIgYKwU+ZmUwqj3qnKSs
lZd/Qf0m/wgi1vOKC8kRiiM0cOfRJS4VgGgwFm4vIYCMDY/qYEjM6bSglHaxqfLt
QuseVgvgi9tMeOfRduLsP/+8zvns2G8cfxSdQIu6+YPgd5Db/mW9200VcZDVR7fD
zAERl0Yb9RVtik0rFlX+qumAae9IxzgXFzTQt7bJ/zQjoQlKBYDCoet82dRDmz6U
sKUj+Kqd5IIkfSHgurZTFR9EtQHoB+BwUmN42D4QAU4fTKqaS1+/x5eaQp0yui0A
nWH2Hu+rwwx6+/bDsXkEQE3OWbFiEYc4gyeb904rJZcaO5u4TQo/PykgU2mSQDjw
oL9qnLuCHCGH7M3uaQE9JNgKfm/phnvBs9KiwH4WC1S0dzLdVCvMHP5Gp3rMYnIv
2Ni9BWui6uWipDJQLmkdNi8pw3XW9KetxS/EQFe9pfCaaW7w5ZQaDpKETzcJT9pS
HZ+rQmvrz5b1CVZpOp83l3SiuEhJ2+7bg33WdqnEFKeRxGCH2vWSTjr6YSLIEgYK
5gf8VQr1vkOzi6BljWelBgxYqijNjsjZYIP36efXnvw1j6SeNz5GTd2Jmk152/bG
tgAOHibJt9cwisjF3k2VjLgmYRFUUtTPXqryKHqKbSX+MqkFtA+Tj4JcNJId3LHP
nKtnng/Gz5/L4zbcp4glqKlXD7j9fT9hmeDNAcpf4qg90bo9hIKNkFmn+vJ79A0Y
eAwt9jdr3oGa8R4xuhco+OYAtWvQFiQ5nIN2XvNzDqzBZM4UwP93OdkHX0S+FtnV
zz6r3HyBp0uxKqD8KpoIlqNVXQ3bRrqTWvt5zFFtG3RVj5dznY/cB5JOdfKu3/Ex
7e2HJMy7ck3wieIzy/DgGKX/c0qSRx1QNu4J/dIX8uR7CJ615rMLadhcb5Pizyvl
+YU2jMPc2EQIbnkjsH97LSgkwSc55tOeHxwZ8pIF/rzpS04xrkmplUZrY3wPvnp8
Hm22+h1DTvvBqOrA0V2/s2fxllDnUArr1qwGcVZSz2QWjNhRgS51oDcoMpQwiFmK
DlO2gV2UE843JNkzNEW8RqVrsepaKYfeCDS+O77mE8gbcmhqOQPIahJ44fKDPX3T
O9Xoa++/3yww+2rukbMb+mmomMWwRy/SuF8GKy+9lsTv+GsIN4XTqs5C4l56oDvw
70zDdgF8KFr5lcxQr7fST3DDRFCxtatTossMYT9d24+HQrsKZfVJp/6YOME40w9L
S/LRXjgHwhmySn2dUNgcZJyAeXk9/KxXRWBDbCZJF27E+4XNpyxdZ8wlqW2782aH
qhoGXgVOYujU9nsjIHQqMPbOJbGbdjNdzj1Fi7FsCQXRj3hLmG+CnLgFNHc4PLy/
3rhvxIwYzmYJvJw+0v7+XIaWM/hEPQv7S0B3rWTgxv5bR9zUqgRGsRUT3O7u3j06
e4IqWFo9ANuM0zq5o4r0x1VHEol9D47+QE8JvjhCnRy+LU2J5bRPGINlZ9WN8pPj
YG3kgU5WNgw3PC2XXlcY13jhAl/5bpbKUzQeTs13iaOsV0uAdsYm71kzPqOH/MG4
8xmzqvOb7QoURZ0XTksRq0hXKsnfpvFr+ymOZrQ0NbuDz/iuScu8tfuc2t8dQPYH
4A4PAlCMnjk2QuR5WQXf7jOnKOAk9gmIamOfp0mYU42T1BIMNSx5Tsy2Si7jkqxw
H5vaDVH+gu0uKwQTUJ6FIY5C5oQqvLElpgO108p2WchidQvxDgopOiYe+3ouGY4A
TI1MguHViJIHN4J57hCL3MWBMvRkhbHoG9i8aW1fUX4gAz8QQ+MV6gYGhnQm3KZZ
TTAqhiUrTl7fw3UxhzxuuwFAd08Od/ZAl2sIAefHjcaX6ttbPeBfyIAqkg4Ux8xk
PW1x3qZRRtCMse1EOmjC/3QZqhT1dtrwW+bvOIZ5720eJksgRY6DSTbZI+/3lz3J
E7kGPBmvSFGdBia8qdnU3KpurnGIXesBFHc5t/dMlKkjU3Gx3s82YHHV7DqP6cvq
oeL5MxtKJu9UgNgtgM6rGsy4MV2pUqqKWn9FkQ+NhP8z56swszfV558gt4C0Vb8A
fSmZl4xobb1RYyMsYvCBnUgmBTqSPzXbTAqTMU+JcgAGkBz4bNisPZ8/7wSiNA9l
SQvdkZlO5yFyHpjw43wLtDMKDuy8iauOu/8bvRJ8vF5IIZ2C3SIvNE02RgHB9J43
jw2X2lfn0N72DgZwKC26jKZ+yn7UkHIDq6qSoYNE3s7FtOU9luIRzRAGWsTn18Ny
LIsbW/bj9VfIdIvPUZFGCpmOgNtuc+ZOYVeW4/P0qgHFXX35Wtwq19ttBsMuidgN
Mf7eTLe5FUU3rpcpWjmYTmaX5EBzagYYu9mA+2m1PHLO5SRbSlgS+CboUIYD8xm6
RWHpaEDFpPQQmsKTOWgzbzSUXhU45q3OP7p2Zw9L5lqxdSLlSvgWmp+3n+Ctsknq
JVLw3JQzb9IFFm+gO82ibpg7smm/6noZ3Ryj7SVlW9u5sxhi2G9SfchQjPK5HXcF
BpN/4xrpwqOl5sgP8O504hkTxSLhZ/Xu/bK5AdQrEhl0Di/WxVUjysHOcDoiiYQE
9aMEM6wnQeatmvGsEF8AdipSvQJLYb8pSzj8Vh5a0IczpEaPxvG/otrZayKWNIDp
YQ1y7iapz550DiRNgHsNFlIB5TZ7bdWjOjRr5D/NpV2tZx/hmvPPtw4CyjYwIl0E
NvKcLy3Er0aKc2YbPt0bBxDKpIBZiE0+PqgxJqVyyfF246vVLjbgCeURyO4d2aQC
W0R2PwW5SwDwfG7flDXolqHUP7WoRLTA2hSW/Sz/tQWx6uE6cDAgK7FVxm8Rj3C1
ByYRTV7f1YFaaZjZjYBvJwXfOitUW/9FJQe7edk1w0Vn25kJ+aKcx4tGbzTqzGTI
RoCo3PFEjbdstqQRgpiO75D0t1TRZuiaP7N9ELm2thydGKo1jo2a8qrH1KT7B9j0
N4pZOnU8iq0zcZ3BQg5HnVzCizySs8sEW0RZ+/R6YarwgmMmaKLWMhemyx5XU46i
hSTvQmgFhQjuP4OWKzgRxFI2AldoiU3N1EzOQo5nnCaDgsTqCDi0+fw6C7qzBKrf
IE8LsSQaXms86dYSFXZWnK3R8R64t2RkekJaIg0RQP42aovP41dOafDNbZN5LWUH
k0IdHkojPtmoLSjfL5tymSJw8w7vWxtjlJi8ctKa/SxB/8ruoVM00E6g9ISxGYkt
TtBMobsZPsY/jkHgoEuNVLjbXT1Wd1mL1+MkRVbAkTq9uwKoiw8u1zTaYYBMZHQl
+4cd0LDfPqac01jnudEAgLjzbmwSqNGvyeeIXEOGs0n1+Yq5/8AmvZvamobMhluz
hUev7SwbGboNzQbj4Zw3Oi5h9naZDj7r1X/jUGj9BGNLrgH35D8NZ3IgOXSXhmwa
pmqqQXqN6AksE4mBEe3UNxdLsaiDSr69f+XZMsoG4IHYG7HYOMVZDR9KuM9zb8rw
0Yj7BvIbHQfeF9VDt4/hoUl5TEJQIca2aqe/Z8zpQYnuyFylA86f215inwSQqYdu
rrYLlL6SIGztuuQ8lyj4ERv+UD2QEFj2UI3O6FC1WTtxd4B+7DavdKtqO4R14/vY
BLJ7pOZc9Gaoa8+VyoLbbHoGz+5BImA73rJW8lNgFGwyyVx2X2PNZ5XO0uQrFXkj
3kih7s/v4bNTBu3w3d78wFP2RmNKsBTJhgQFr2ZnUbEnBs6/tZt4VJ1zb35smNCN
a+MuM/xMJ7RG/KgQUHwVk629wdd020CrxjLdRcop8aZojASmk3TSmClx4NT+ur2y
44cpg42i34v3+aTyvzhgJ1TdSzhGD0Y+Kht4N2S8heTkC7fCTRJu/AQ3DTLA77/D
eim49YKpQiUihtdWVkdj5I4bDXT2SIqaj5xM9edqA6g3K6COgagtpBAPlnPdlN6y
TFrsM5NmbLWjqc8Y7dDqGBXAQn7L+83PzkUj95gzys+T4P7DsUjxMpw2Z3JhdqaB
fEVPlQ2+aZvJ6LV2tr3peCtIs4Hpoh2uq0GVyVSm14zlYp2Z8uTeY53u5rauNHVU
yQkyUwaup+Nuud3FiowwYwTe9+qsmf/aN/4ImLHeSvsdHktOx1oD3PxKFHO4dtnl
dkjtYoS9cRnwnWXVFxPsE9N/5I6q7fNDiEh0mgBu9WpcIVLHcO67Kd/oSobywzdi
auw1883RKQ/Tb5P2P2274WPhVvaBFmv+gwdNW8RfCOlsdhDJdj7G6GoTLpRqFE/i
V1sApKCounK9UQpENA/2o1L9FT4jxCxck09rKO7lb8x8aC9c8ynPWcA4BSUqG3RJ
TV7B1ureLQ/wZ9s4Q/LuQClrjx5Gmy1avmA5ZJWXl6IV+2JQNUZaUbVH3ctDeyti
HvQW2DPb+dwc38XZaacEg3d0NH/vURYMo5+yok90sLACx4ojBZ6xRtvrfgMYipgG
W7gJc0QNAvQ0PrC8Nl7H+hbJQBRZsqZqPUJ0Z9jLn6JJv5cvI+lZO1uiNz+qlhR/
c+tw77Mv0ilCDcA6iouzGCCduo0w9cd99mIBN99gu4SGj9zukfKrIsX7GlGvE4kV
DLhe+uF+BRxs/l/Sg6NpEQ8eWaRF0SzYbmMGEH/2d/bk4R00BxVwRB9MUC3FWelb
wMsjbcz9ph+POLIclGgmJ5+yDHpd0E/HEO359I06MMPHuLFpl4PJBVMdLaB1D6Be
ZFDd7abbxZ8FzoGAMR9qyzZshqLSf9ZE188kbnZZLGPy9KxG+LugK6Lep74NY/ag
DPa7y2GdOdoprvO3s2kA0h46cZ4Kr/xZ87w6liK8tPXY05tRC4E7R9b8PjDG2x3x
WNrlRxtj9jyp2kjmMnwrCq6JX23pMFea2t5jru6rBzjqRZN4lDWX69Pk+tONzbep
4Y0O1n7fH6XM34sxpUtufEgWXBeZjVzX7dY6ouIhcv9kCBtQp55sgHtWjtshj5ag
U6iP6XXyqbB5M9iyLkRN9nHqKtxRwuDAzazjrmREwjxPq5skMUcb5JHvaF05rDUS
jFZhzd1PrGhUUseXnQIoHjnRIIcI7pAtDjO/xb9Z2qb05yxXpRhXCnyCa2QYergT
Gm6Cffekf7xvcdE4Otz7JmiLPdIFn/PBPzb6Z4scXh5sNvViIxsWYKA338GJ0cGi
04RL1NrArztFt3WHQ5NUyhzwj82rDqNTTKWw3HYbpP1nXzhBN5+Gk+oIWDTW67A1
z1h1WsfSvPhnHaCTlxt3nncdJKDscUEAKICQuKNgHDoiucTvxXWHjyqaXOPP4yVC
/NexluChhYYPCTPyDkdYG5001368mXXwVxaJutFAkLNF87r3lax6fSy0ah+oFwIF
iuG7o0ScrFiasPjMzRQp1bDst4omH9e1mkuaGgSACaqBq/qkRHHVfsqovuMjGD/5
ir7m1QutBjSdU/4ZLTrsWfuQTaN0fVLNOUCVxKU66avjCetwuUTVy2WkivKQEMT6
+GtUAdVJYlj8/XCOvzy1vVdpeS+yjnJpoNLGy5yf4kA9V8+FMv8ApupoeS6+/mmf
yxYAIoQGgdqBWASj639Vhxqx9vlOejQZMAkbXwrxM4J0QxRWA3PdYNnsHPxlx4KX
5bO+ck3KDFmsdMPDV07kzRe+VgFiZbe4lBffi7C/aB1GR6lAo9huXHHJPqO9hcPh
RrWZCn+sl4SWUt4NRdt8Oq0Z0LhAG3LIE7RXD7welIZkKOVMKdIu0AI5SAkgv0VK
Tm5oXIvHoRfgMa6yRcv05ZdFWyrb/MPU9lLBOvfA4U1yyEZTocfFTXK1hGapgZum
5LrXSIsYxo4tUoUBa+1cdT0FzoiEw579YtLt35Coc+PjhivkHqL/YdnaJT1CW4Ki
XRk4mqDgIgUaSApfV+dPKrG5fakNCXeRUs/Hj+tLuCTMl8dx8cMbJuhzK2OyzeDX
OoololNMwQIgjKGJnR16QvfkXVPeykWkI9Kr30vS+n08kK9Wdti2LQcR5VGyDpVl
jGTJSR75fkC5QzUidOAQG+W6JwYeMWUU4o3vcJL17nWclLx1CbpydAdfzv7dImj0
m3eOECYRxDTR4QxwgrWGGL4P8QQDOyh/3qK7t+DV4lejMIAXT8VJDhM/1Jp87mL6
mZkbDERYMoLAJbZJkxxCzSZY8FVz73mBFJVtdkFoTrPBTuYsgc8WWa4b68SDXiHJ
ZCod87SvnkNFwRy8YHAxpqFZA8vKwesIR/n21JV2OoE+SQPeYaqqK85quPT/jpNP
NT8J0HTy514DPA1VSJpz3ExBn2RwFixxpgQomY0oUTT0FnFvAkK+1VrWzGQL8Sk4
qrF22+OOjzErBhaYUqO4H5ed/EtvopuZoWAbUEdQnlG1H3D32peZQxjkz56hO2n2
xjF+Uxw2wOq2jPnZFxxQZ6N3PCiyPa2mQewlad6UBK/CFDE4pedhuJBRgKXYwQlN
3rueUeF7/ckl5I8ily9yIV4qb8Jv4g2wsuh6NwIVXhGTp5usp7Nct3UqNUM++NSK
pf3B2XVv6Plr/U7RhdgTjt7LmQm437RWxPUmoPmlWS8jgbaX5DT6TF1oDY5bc5+g
P40WfwOSVAEVc+LDBTkhK61p43a8SJe4HYXy4h0SgDKBYKr+bz55GHpHWIcbfDgb
bFoIPjHUIzOis3jBWHU6zT4zkDqOVA7ZGOo13TxQcoTj7+PjDlqhkylzzz6JljW6
7X6gCfKHBV1DeEgh8yuUPyPcGW0ysjUMnTflU/Tjs0BGhINjOD6y70nxTKH9x+st
M8QjvRjk5bI10ZU8Gi81wrraJ39eiviYrteamOEZB9C48woff7q4dv0O5vCQAGjb
HOwU/CfrrXaRz/Op9ci73zI9fjQ0MkiNY7MmpYixDMir+CTWjWe8k9KVJyaZlXDl
ih3oriyeCLqJ93iAss/i+OsEvnK6GJfh2LkM0ihx2IGzX7QpgZZCNDuh4HiM2y94
yLWe4FxUpmgGJLXLgidRbyZoRjj8/He/XZIT48S/0zKmD7M63CJ5BISW+rJMTyxg
mIsIpQu+vucyCrAGtf+flhveOcYPIWC5DxZ8jQI0JIriwhor6TCo/7MPtMpLrESt
SdgaR5RYAZU1bK6HTMPEGL1G0im36QXx6HB0gPOTg16TCDhgiPdV2sp1SU8tRiH4
7R1mJNO1vHZW/uNcM1ZndjHffTe2+YIrQQQ8FliJbXQ2aa+kyJW6mIINrvCU0U7Q
EnBo9ckrUqtuSOHbnTQ/b41iFjSKa6OoGiCaUlCq9x3KcvnQRbmDuQzcKF8uGlfj
QSrymxwCk+3kCiqiY6wjYafp8fdJbG0VFG0dWVX21oHMy+xbhEmwCyXYKKl5e3tL
PbBI/TXumU5ndwDAKz+RHZYLYe9TCabEamj/5gHO3e1Sk3fi7aO+KfB7I+EmYHhs
pQRU8wJCRJvyspgMb1hrcfSIcelMxmPNm+IG14vGeJrBxUF52xAirave2/3o0SUg
0tLn+89KGDrju4j0LCQQALAaYqOlSwlSnY8fbw0kIgrflYOr69HNRvlr+AfJIyVh
TMHrUQKMVRsLjaRJeaRn9Mwn3Mq8VGJ1OR/D8VxHR+357sCxSMbtzemX8zwggXOT
9j91ogeckOfWwEPh39rJ5yoTQwsXkJc+vtN/iShgKoKJ6boF679AqyU3QczeFHD7
ZtUBP1CzvTLMW3Agk4aO5kTuAnDFtIcBVX2Bk3GL8Ao2yEvK8pLLui2lsrllXlaB
qE6YgvP6dqeAVzj2cf3wcRspQ3kMHzDZ7p3opI+63GWNYXBaYlV9guKgMR6L/Js3
aWn1PC2XVH1cYsEKQ/Z6/ZpiSBrWRNHU8WO8BjfOJod3pVO1VvkP4+bVxdhJ7E9P
L6FkigR9rTDOKVE/2RIn68/RCYSuNCqv7Ds24qkQZWSZua0KjiDvuGLd9w0ZPag2
y9Va8N/QkxVubS29d4qg0Fcv11qbZdgXJDbW3hjZap6YTqs+4JqAvMcqcJBj9sbc
zbZWNP0WSJzklpkBoPeUglMwEOS0qVcinC3LxW70tdX9b/fI0UG/IF+PjKLoYbtG
fVOF/HKX9R4qWhu0ebbUIicLqy2IvmmDSXh17XLRdBGuN4TwVENaevnYAjcqm/bm
vAcP1j4batjIc4GFHS2TAgA0XIJKLzaubdXwSae6dgfW5Yy3GH3hsJcsFL3gdS/C
EoZYFoIwZlcjZLFYMPE4/OGLmUHVIZsVEJICsjKTSAoGE1WzrqSgJMN3wyUUDyFH
tXI09NENGKCOVPLRi8bD5aWVlJCm8xODSENUUJUYQ7PiUHu/0TOMXi0G5NfO2x08
GWZ+P46+DkDsiO1zRuzAAzM7k87/S4fvKdHbTyeZSI5c+xpUs7do6XuPoSwDPq/T
G1Sge+LQz0b6u3Qq107XslCv5WTb5yLFZ9FUXD5SsDX2Ft9rk/Cz7ySCo7+ZMdEd
LAfDxpl8KDD980nJRk9kC7wEciJSQ25IW6jhucdloWqK40+6EvTHFoze+3vNSYHj
WEN386jz7lRCCKfrp3we8Y51n1mCpfKN4hloLcXD9tr9goGebF0bwyvgE1wS1bvK
CEEIdQlncBrM0FwKQPQHbIKq3Il+HeUfX6+P1DM+DfrUqyeZ9Jcq7IeptQz49Wvd
XdcO4omEP1CRm4YnOiKpN+RdX6dkxO+be5D7SrCtHcROjtsvjjlXH2g+kl/lchYr
oPghqwgi99RAcsdpDpH5zhD+RWVl+9ZRroa8gMljYpJ+hBshLQ7bx22qtYCgOeax
9+LHs0aLzoi9r/60+4u7rZQ9EqJ6tJ7hm9lO7JN9uTGK79a2D81E4JBqNpTAZ8/J
5Z56e7G74UokP1/KkDOpFd96lVR2ubQ4xm6mXWl04e3ptEEcoUJK6PlbccbgmBEt
+mKXL9kC3/rX+Cv1HgwrJBDz41hcJ8txK3qkHD3R+2sDdICxFHlbVr1KdeKYvck5
K5ySxGKELJnZXTRlwqJBxjgHfNVxWdfXmGJdtOXe0TYbx8OFTs6/nxRLsLCeLkYk
nQoXVw3bUt07fEZl3kay1RlC//7V6BrEEvxBjdrGJM0yDltgyK+a+KDCPi+4CRtx
z3Bb88IUpIyP4KleqLaGiRvkuXh+MFMLY2+SYZ1rk68NiBin+O1UIVRXrgOM3N9f
DZm24xsqqniwuH2Xyqsn7LQ8k7TOcVIKlBgdrw87L++FYMxTRrFQ8s1Fs7PNC+AV
XVPYogUvMocP2oeq3omdf1zLsi+emKaKOTNWnokypCVyoqp07jh7xOJUt8GX+yWa
ESB/JzvfWWMrbbHrISgtiH2srycCFpUWmcnvFCshxjREDrc3g4rt4u7MA7QUEyOO
qNuzJWhJmTqQLbJN+IpvNjGUXAxK8v6pL+Do4SXrNL4EIEpSK4Oj1uVjdhY0RJnW
IFmMhywMNqcw7N785maUqMV48Uk9o9QP0O37PFreVbuA7f3PFbW8Q1+632/WWnNN
Z2BZJ5jOqXGb8DsOnhlZAsvnoH50RG23wqflWpWpOd7MNkoIbnFD408r31F9vOIh
k/B1l8AeK/ks80L0sRbgsuYyhbQ6V2rk1H64tFY43e5W5yKpgmOTaEzfkArwU8qK
WySaXcWHuOXbc5qSHMzs2MSnMaXLGoAbfuRKOv4a4eia455xqSk1kYe7rM4dCL/s
G0swgGnGofc8Wf0edqOWvxfrJD8wtYsu9APP/3w6LwF/tZn9nvwSJ8c6sU09IZ9n
VSrrM0eBRZr2NtlLu5t0IDErSrMgOFHlkwwfchU4t8KXKzRGtmWF9natXQI6g5xn
lu4MxzfhcOntMaYxsS0f4mekIfsVIfAsmWbWWz+4GzRLQcVf4U5rF7RkRrcJJPwy
On5T+1WqZY3kwrqLE/H8vBt+vsFJMgf+8twwHNxJwE/glZQoslMXZCr3hn8pASAv
dDmqTCoWYUD/dXqkdZeLT7SXYB7EewOgSwteVGSgYv0RyV7JnYsmHfVJiY6tBwpV
8bYlLX5lwSPoYDEOEkuKBnb5EjRFtglzdv50l27DaM9CkvqQ8nmk54K+rO9Kpd4x
xDo/jsdsFzD8mZAQf52YRss1EMwxjtMWjwgypzYHMzBiXvMZ7M8NMXhQVFt4WQUj
yarSZtqkpnxMWLOymt9XZoeNe+pUEIJXoT+jZGWYvoCCi2o7u3imCOt/vp4eWNs6
v/gvUE0u0V0N1ogXSja3kMpI2qKsoKU+cM5Ivi1bd5qHHT4e80pQ0pqINxPFoRxf
HxLsQP809vmGcyCYRQLxPtQ3N08oBdXOmL+WAUAoawPvc03fsQY0IX2pAxhgt7t/
bKu8CHqMfjOFmCJPml/zCAHFsqm4iT869GBf3SZam2QLo1yN64ELRfMW2Fki9WWJ
PAXsMC/eSueELyWs14D69tVGGJqA1ttEsJqPc4hOYuBACy67Llvey5G0NQCuXVYg
9KA83bku9N3Fzp3aCU5HtcLTqB8eh91G+0rwlgKKw6HEs8EWjwomvojzfCuUwkU0
ZPt1LJWuGSrWP2LiApI+Raj4A+NGi+NcyyNwwwUtk8swv70RC1LtWhHEqORvTG3Q
bfgv9ucuvHbboByKVHbyZSz4C7036EUnKxUQTJVmHAoMvwhdvQL8srr8h3JQhxwt
o8LAk13rZFVuT6u5/BdPpw1g+q/76AD1IWSlZ6xag+tPk8X5VS6oA6c4c7vHpTkj
OHLSk0n8tpeEm3vitNrDaF8UI3oQdWnLWFnA/HpBd4CYJmjnxEsclfftHxQxMN/V
+/SbvHPiFb80NDAB++ScMFsqjm63+FprHPo1haU91VehDo+M95T2YqEZnqsXoldq
1285HCqg64xsfqBtiWQt0vFZ4HLjcndWBeNpdq3gYxcqx535/eoI0WqqSOr1p4lI
Efb/ODlEmaJ3GPb3j8rrntv5lG4RpdUsB3t3xNF9s9vSfTjeIfTm1F3UkJrV/Z+g
sV3GDn/zMyh0I5u+eLxUn/WdCzAX61c2HfP+oLSllzJLmge0g6u+VshK2hp0yJ2c
2hg9RQATqusObWSNube1hFfB2YWbOP4aCUBf8PsAngS/XJSBKDGDrSVshxDl6+Qx
7hyfpe7EI9/Q+KSEAMidL4OSk1tEHHDqVkrVLMCK/h03xFSLa3OUrtN502A3mWfT
qX+KXkptGfHV3p0PSkXNq1Jn0PayU5caTZ/t2Vct9umirABgrVUuRMy8M1k77sDg
mgmPDXzNcf2f6wNROJ2DaVpsfupnNeXKhRy9eD6Amm+i451FPoYdGZV2WIbIYIhM
9Y8Dkbj2MqM9oiomLBivnasthiiDoE4xWTVi/LQOB6XW3NkNQAJjKbOHgvz/n5RU
abAA/eh/Fll5YjafuTML71Oc6Bod6ELjXCUTG/SyIx9PrAlX1zkCcUq8LgduSfdU
G+VGKe8m9Zf0QrGnMAe8ZulSUBdYYqf/fpRjiASFa6vgxt7rjwm96zVgUWXQ5PBR
0fhUYKw6HQcfCqjYGj2eJ7fF3ebWZfCT5pR843XtRP+p2JOJ2XmuQVnyY2xZj8QJ
YwUZRIMwcWObu9INquEno98lDHJww+wK0/g6RiyHiVguAPSbL2suarKZUSgO7VmP
KaNbIxMhmLBnRTp0JO7EpkPZ1yWBz/cYP27g3vLWChOPovYbYcnBqSGA8TmMNWmJ
2J2eZsT1q2BB2Tis2tbkvq5BayJ9pnhf9uHYZZOAz0/k1FSPqoTz07gGssJy4YSc
Qze1vd1xleRPtf22UM/GpUc5x1lAXfPzOKkFrq8lh/VACCMtyr0+yA8X0/HxqRhZ
osgVk35Y27Irvp5UEQXrh51LwSZd5fBAVJCmfjZecHGxe3Ud/YwVcY60hTjK7YY/
AWYSh1PXFRZUTWvfHU2ipVR+Kd2Qw8UU14kNsfV4qSsfVSQ0dU64VS2QZFRI2y82
SplXE4xyiDmTuiCqAtPIdnAfdnHUcMqMtbEQoxRYOnfYCXtlZeF4NArmlaq0CQDr
1caBAw2IzfOwBQ6bPRsYXARlyCpTylbwVOIQ1NCwK7/cGuG4jVRfxDV1TF2soOAj
9aeQQX/y71GOWBa73oMR9RwFFsabfV0dShT4obIokJyOjGV7hnr8/MCutOhRv/eX
MXHXsJujQkX+6RixRCnpoXnjiTvWZOWUOnQolFHrXNBPeMlLzFJbjnOJLgRkVSDX
p2BQh9QjjWLiRmfyOIVMvu5NiYYUy1yxt7z6mL4iK25rNUBT4u5+/3DASI+bR/A3
QX/SwKihYso9VjpKryYiiKORN3FVq6HEtSnMcpXMJW+aHqB8EytBzyAQ92ao4piz
xv9kKnaGNTK1BWXECuf6BiSyB5rapmCJ+VYeODqt1W9YBqjp4pnh+cEQ1EGW65ZG
Iee2c+tt/z9+EeuMsvIqyX39Q5/JAEU+OuW5drDgh4ePN7Z0XOAJb8Quc/rNvOiy
03ZIQ6rWs0tpDrLLW0fNngqUKDFLAItLOjRmMgQvtHj2vkgyZAcuxzbgqMpkr4Y7
TIcbNT74TDO9yAPJJDwFvKjgL5aFosLgyaI904PMwH09T/M3MHFV/PtE1L6pHPEJ
8fWbWLIwRZZLLcUJ1di7KnA6nit6WBbp/EIkgIRIVjgt/FRm8YjO4dygQ2+61IJB
G0s/shdQf4WEc6jlaKAW5Ulhzm4MxJI6WYo41J28cfgxOUok16Jbyy9oUBAWHWOS
UE5wQz38N14p0KX1rXvROA+1RM+MnM4EymwzpCjYURtF5mNNzo7MYNV0gF+j3mz7
vSqiG0WGtY9E0/y2c+II2wpAcAY/3IR6WXeEs2MXnz2qYDbG2IfbMqgB1ACH9l8y
q0Eayt2ST/VOxbonK+a0Z0uyOuoqhO4r7ALWizN3mxUSmBhOvCCBuF1ZlZDMaNhX
n/icCOvHZhjTWFeaAvR0lyxPmXpGoNis2gnSDFaQZNL2agci6PwWWMLqwUXC0Jqr
L+6iCi98js9eoV6fr1Wv9T773mRtaiXDCBPwoHZJrUzDisSRhn+f+aeejPQYnOzp
LiQpIOPGcj+lz1vQIrKzK5snZNVKQNlnP8Mrnygm4ETsqEJC+MiNjfctnRz3D/ec
JltG4sjs3LJpNpiBkx+bxYKcKRdZDXdK916CffrMB3K6ro1uLsZWbco4A5xf19zc
u8Om4Hnm/wJGZrH9v39rxDpEdYW5orFeR1LVS1Z8RSeaxSrridtpeQEFkAHo7NwD
HPpk2SXEz1yGqg9+2XnPpIh9VSGHIMK9M3gNZlBXKwgv9SUvv4feRq+m+eyLBhQc
Y0Uu0REoF69CVPHznschOJWJ/V9ZDP8NFzPu3Nz39QN9x+Yytyay58cOpvpl5lZp
02Ibx6P3YPJnuxFc23qw8hsmen7yxBRVu7jUlM1wSbU5XpkM2oC/sn+EFdqvApYt
5D/JBcwoSHjRMrMGj0llDgyjicpqYw5kAlKmK0OAxb+xJEypkcfEX9kky+tmOYO2
on1ZKRLiEkWu13xfwPol28BOPZn2jxDY/BmAqKhZpW/CG3jlIRL0/jaYWEmpOGId
dKiJsHs28P7IBzOCqNX9phluF65fJJxaOd61hX7Q/Tm2czFVjiZ0ywuehjhqEfxj
5Li/gYeq+JvV0qnOH+KMmUH2g5EldJEqBFysU+S7DYn4tuEmtJSexooTyTmL3meS
Txm9BhnSQrDP0aNbKDIOFul4x0n4GFj2MdnDb4oJrxfVPn1INnl6mlqeBBoFBIo6
UWDHXP6YhHtwUekj5zVbC7ZoiMiXDUZNblF6f7yEpksS8lAKPD2Nde/aWXjQ5plg
pEutka4+zmPtWIAiml7Db7BExJU7ezdj/bCxUWGBJQY6pPUG9ZVgv8OExbVPoGNy
xgvr0MziSVCtV7ii2zSef+fHlTWVS7jx0UYoYXI8S/v0irrr+9b+tlE7XssOx2//
AQIgRfuji5ArurjZuXZjW6b8Ye/zBddskfGTvK6Qk3YhoQ0CO9fsO1ij06UaFpRS
MncAK7/TlMWedk4ovKOUTjw+ScPhnzhk//bbFnuDMLWAkRHsNxo7FChoODaTmXCA
5warP0UDFpBBORO++ckC+1LolOR2Y5pfwpGenOtnXTxqrHcSDYicPtLv2qxEWR8N
7X5qnxSaDSDCxFRiBCK7Uo4r8rPsmMrGsY72MNDgy6LdyPkLq/bbzw6pGNxlw3TE
+Hei+vUoSgtCkCG5K/2EcH2zK4fO6QmlIMr5M3uvAHowzNzhehplUScggtMT3Q6J
VOE64TeQ6nxe8uNuRy5WQVVHhtprg80MpNNGQOXUR3ZPLNehOGwk1yiC36gqfDR6
oYpyT4RG2zyqJozHGhypvtlM5B/SNjWvpVMJRXAMy5AoOB0Z6PVbbFwqWmFMxJUo
KBaoBDANN0/AsCtSXwrA9yOdpQIeb4WvraqAr4c7i9kqW0hqfITgGqE8PUfk4GaZ
EdzWB8m7MDC5cIIwzqzSVx5CboGqC03wmJQON5W8AMVOROsPu00Bkd05EfrXEOwR
OOuhdulE71qZNZAc3cTfKk1GjMybHDcYbbDPTySgoPwL1zvEQGkuZD6Cl1mkyQL8
s1t5321nMiZeuxzPQcmZ2RWeowL7alc5MzH+2skISkLw0SjrwvNhC3ZM3bSWeUWA
+85+gZdD392xKc1BTYIxpTsAN1i0AuujxS0UB8kkBKqYzD46fvUL0RzhyVb88cIQ
f2SO6LJ7bRaU6Pe5PK7IEgfnzJOodCqDm+G2RZCGC8j4P/wtUUfpvQ6aLbM8C629
KbnHwYxQklyO9zDRPOC1zZSix07h2TyFkjWSNCbH3Pc36CSwklLpearhYZdYJJ0J
/8diOEZ9gI/ccwsfApqO5mVY0e7YeVtMLKmxDlTx4g5gQ7oJtPZqV757CiOQj41Y
frB+Em9SfpokZnlB/8T2j818768EZh3FAEwUKzrCPFbXziX2ZqU8iXVu0gwDpSow
XbX/hb18G3zFfJHHtge4GjdWW5ijri3zbkHothE1ypGE17hnDZKOBymT2+DUI8IW
x9KLT2NjQc7fsthSSPLQKaqtpMJt/sGDLUs4s2mbn+P+VIVtuTWmPuRX/Ry6Jphe
BbQDxPz0FUP6Rf4Vne8Riwd9AEiugTnEviIOUhWuS0ltxJXCUk27/RdX3ynpistI
sMeSL9oaTMDT6YGWWxOVAY2Ekgtgv0edRor/vXcOvpXksVJFaPzfuwcKW0RBy2cW
9G37XjNiBkaJP7vUwhZ0IrmKPiomlKaobNiG1jgIxt4WBteNaXbF+i3cAsqLH3yH
8bAsY4LPrlKgQmT9HjLW5Ckb7seZeCsewkbIFbAOvjiyT7mutjW4yPSNH2QZ+BEp
TZfJ+6DIZTLzTntotPr4FsJcv0Uu+4l1UloUt/KHLqzYUkWUEx0QkDuf5MpAZ0i3
y53NgvMKTCxrrv/2Ah8hJLgfqZBrnmiqwATPPxY/VNmb0h31bP8uo+aOUE3Auud6
InFOxDe3S6vpbZPtKMUUFhCGUsMx0Wlyp+soPkq3YxOdF25qWpDXXfnjOmsF/vJi
seKyMxZCVNea1xi82f7VQeuXBZZE3W8c6r7ByUXhAl6JKMF6tvJK7l3Y6gCtqFxf
8QOvRS9hozPyNsae0wOrAUzXtK4tsHJWsCkW37XUZDDf/ffQ6/Q59tc8jqlPbrnF
T7YR3tLI6Z5RqM8/kcqeUcI2a9R5tnnEkK4HQbmXwzXyqVyX9PR3LU/t7tuY1DlE
gnq9makhkS2a2EIYCLn5LnsVlqDz3uvb+iGuww6+Y7Zj68FfC+ALGp2LwngS5HNb
GFPytFffttYD3lr0UuvFvjPmVQz8qOUw0H6ca98Cau6najBdZrW3J89GWDGxnKU9
AtN14ktAIlh3O4NKihrmdGur9pgVyCKfBUzj08qkG1MGDUcYmiDfyLihg4ImVrEg
f50w34qAtf02hCbHzClRAYLQWpIYN8bk3NylfHSyCJg3uwVk9J3c+YwXJ0y+pQpu
dAGAWH+VP/eZ14ssPwjfc7gjqx2OFefxu/DQokgcAlAtg//07vfh/5MsC3ViOHy8
OnOsOT9B+2N2eSr0b9Wz/KVBmJOTbSwVlpeKUuwKZwAdWH69tkU+xtzULwrFo3e2
X7v90bhOOuKUo18hSdO88IRBi2D7D7pzV6GaUSo4xP0HqhWk9k/WLLPCgMQkrMMg
5maJk1Dh69gGpKhvllI8dS/OJSoUjMaCRotMRQxWUumsNSdkTiBqReoa+TGEojCR
dqBw7ce56XXHgyBJCyo47Kqt4UPCiXNV5u9UqAchi57/cfcGnPlknK+W51D2DhgW
AJ28m7ii26sjbNabrof35MW3DkNH5JzUdyn3Ghb1zPsFxyDpS1+Yqib4HdX/ibFe
WbxFYToCK1MUJJuz+66B1G3jytDaRVLBLwrEqRTXWCG9DCmVeAsDqGUTHPIoTR1z
x4YQQUPT3XMsM4erQsFiTsnNqWSCsdkN5D2WEO6Dyw8Ep0zaXrGiLDObv/HJHHZ/
D6I4gZ5C83ojkb1qtBp/BdS6rnBELuKPYJQ7RInqBi+sAJoTxQsD3JoAjKvnBK1I
F5Pmy51cx6FmggpuEugDEV1AEEWha7/iqwh06eVOzjKnN2MmyfUIF7DoU78zLNrB
HwaqqhKNs3HdTez7cqHUrtxWfn62o4F+HT9wkT+ZODnU5jF0I+/Ea1B8AToXpjB6
kepl5hch3EABOv1LouqghFl+MIuHcQ6CEHGtiqCwCoHva8G17QZR3jb1h6gbD55g
RzJLcGElHtR7H/OKXNwKNwJTco/KIL2Ud6eR9Fz7gvLUFIHFKW8EsoBqQjDghC8P
ijhrnpaTyv8K6hOIDNeXJfNL+k5Rd/S39DagmyT2ci6LXHBmXD/43AOp3FcfYNnB
vztAZz7IJTGM5OfM0PJs1AgdQDwU2PQUyUjkO4pZnZ1rOgcfMJgJbJ8Od2Qn1M48
F335UMgcBeIEayNp08JlhN7I8nXmDRPIqemXVlbeJdV3v6MsYOx8wtp/qPPrBl1J
HxB1FIgwjTvm0wrtCKgGp9ENAZXSeUzlXiCtw0hjarP5jgj9/yN22ZrM2zMlP8Rm
bGPwoYVcszncFVzAVgK5QelpyozttdB7ekGtVQa+W9GicUebRD+Xm44J/ImVj4zE
JLcrAMS6TOeE5EIcrCZ0erxYrPF+sLiyfeU1+Oen8Rs5X2i6dm9TyLS6oYgu/0MF
7rKSNi0T3XBYfunWqummRlfliX3mjxWtXbrkZvjzI3W1kfwB+r3oDvmJOcaYiIwu
NoHF8nLwYk6uy9tb3oitizBLpB+VvB6WQleUc5KVRWIt1/+yVUUYY6YPtQ4UtjOh
o/8KXkdWflKRok2X4pCp4UulAvhiTcAHX/D8gdmOGTEBKOJV3l6yEcUYFJ/hklGm
fiFM2PNPvDt7yQEON28wbADx7WuyLstuV5pIeer4m31hWfWhJ4A+Szc4E/Bi7/BV
POnVi0PTwRezXsWvzd0qDlpAmb7ZZBtQxDTuy4jT35Ah58phcLWZRXUC9GmBkD2p
gqZ4HYiZPlVVVqRbGlFXxXibsVQ2kGMuux7FQ6A+X6tH0twk4MFYbTrm89ssKwJP
61inj7yz3/I2DCH7/yKmWSO7hj30npnnE3dIv10MFN1SLoTZ25wbIP4J99X9xk3G
MGF+Mkyd1PsdI7zPq3KteVIdA3U+eq+NQpoFVSER8JaDikHPLQ9t9IiZCRLkvczE
JxhSjlpKdD4pXU8MTZaTXXTuttCqb3Y08IlTY2KCRet1Gf6Hdx1tAdljbPFCPNjz
jIg1xl/O+Ll1+0HHJTlbLvDQo49EWGg8LT2INP2YjqVPyY2JIUnqvo12wwmLt5ES
pJW6UkLXkVH5gUdYPrHhSRSQMcNP5Xasa3k8gPocUnWsdfsACy6ybbB8k7ucczzl
bZXjo1gkKvfV/QJybmt3TTEu1+knyJ388GROwpItPB1GeMyn7mOSFYwcsCXbh53Z
vCZP1j9bV4m91YUG9gBZumzdSnFgVTYOeaLdgf5hckMbYGuknrA4LNlLaoP9kB7E
IXjjnMnHJCGqysENLVR+FD+JyFwnqwCKyWGX3K+XYa0z6neX40LY26aowLMNU82i
GuOkL8c3pGXMTz/JvEwJbifdS3yyogk/OqrgvLwBARKjFQ9DrmHKprC+fUQriBwY
nbReA5qwZ9FuH8NziqoBjqmBq/jCvoCfIo7Ff1Yz6DuSrJerajlPVNHIJ6RrsvyZ
NNg5kER+SvbbERzuNlhIqEqItbr307o7WhFBtzPLwOIWa5bzfib93a0I/WrAScUV
SXvTNbGSF0zQSyKOhUExARAfIKMggT0bwLDDqyjtXIaUgEcv7LICwv4EzJd4vFWX
IfwOjq+CIFgG/QmEFZot/NbRsgLR5r9hdSQWRN1tBTdSoUaS+7WGqOjrr+dwfsKE
pRXLVddn4DaEXBkMhbChIaiP+kknDnrW/rc/Ee/PUc8WPNT3J3EQrsPNZbeR0ZJf
sDVik1viqW12QWYLY8jRVm7mZNXddpoUYnRM1k57hpq8I24iOrnp/FvDZAn0H1ur
9+XcKaDzisLfbfLKJ0Tr1nDER7Ygf//rQXW3Sbm3zNCQfOAa+FgyCOQdfUVCzjfx
JqM+szDs6CXZARja4s7UBNOfq9uQOpPgmNugQb/RLkvuN60VQS9AFNUcxt2pLakU
NrvfjCGnoy1WmFJjJZ7pu3EsnvWajAmSacu8uVahyzW70fsOWh8Z5IWfmk5acgj2
L4GAk9X/xk7AMQh5tYuP69PBLPLSySJBQD1vY3QaHft9sk9H1EhDmVCDcze181nx
XUl+EqLDVrrUZpDB6xP2uMcxx1x7c963euK6Bofpyopy7dIwRG+i88al6vJ0oja6
OzDUEb7ZfM+O1ffd/OqvL7dw21jXNRxI8zCB3mtLYibTtnNukfFhh5TJThZ3JYpy
SN8iraoyUuibrYCH7PwcwyZ9X+arimhDbRY1MorYFX1mb5fbl7xQUgg6iZfVCp18
MvzNvaN4+Jyi4TZJQoyu206dyd43YmlfShAIPfOD1GdTGSEk+31WdVzMTnt2ab1P
4fVakkXsXOanLltJTIDW2yA7IccLGCuYNuP91y/itEqDvALSInOUX+JxH/oUNaWj
HHWjvxoYlCa9K2UFFx0rguH0Mj074wYbbwDZa/DwhDdU3F19+s864dcuwCx4n8Pm
EYOITdtXlrtCsK/4yb4GBBlceuxV6SDV3tJBeII181UhjI4I6LVok9iK6qZyGtwP
G6Ha6UKChv95fdqv8cNQGCoezmUbfqx4OoZDMvZ+0TVBDA6P0sr6ci75rLWKrnLB
kkWgr1yiM4Jns7dPb7hRYeGMhIhhkeYb1pN6hoJwP/vM235Pki/OcvBCeZnqIyBM
SXM7NO9oWgH5nqLHyfFQ0vb/ueU4kOlwriLDkIsZbrAWu/LFv3J2QDWWB0xzck5v
cRrMCAO4oklOyf5fRV2g/DiSkYDt/fiNetGGihbv7ef/e6ZOs0kTN6xETaYyaxSC
0hDeapCS3nwgqVa7Ig5NYC0aTRn0JatST3c212ElnQqwSl5OPVeQc2Vz4UKH21rw
nzcfb+9PpdApFA3Uiqx9i0sxfCKT32RC9rdzFWZRWEN+pa0VM+jAWBCINkjeoHig
gfLT6YojldN3YOlr8B7iRGA7iSeGhqwAWcrAX5AwuuQsUOo4z2r07Iucf2P9egjt
7XbXkyWLg4/waTBNI5uzoUYS+aGew2wkoBbFzLuAcl6UDIGMH6T1FN++zd+tlTMz
P2TgMRXf54hS2sgRxRde4w9TBXE9YYXNVm+uoX87FSmTx2PoYVErW78qXhNMJV2p
jzYNkgiW/f2ynfHT4FkehnGWOPQwhjXedcRP2I+S+vjqADnFYIsCevKSPVMxypE7
w7agJRj2F5EZLOQafoQfIcbB8LU26k2/JrwRQ4Jo/XEo/zJasoQLJjfP//hfRUeI
OkfUNmrdSY5q/cK/7M6gcQHOvc4XmIYWxhuGJeNJ1JVB8Y65f1BgZMTQvMBZkPA4
/ke32KqMtm8iMxxi61xtq6gy6E/yOhvxc7itWbj3GNwV7vnIZYodE2oNZ1at+PFr
aN7gnzWJFIl7SIUQso9rjsQ6RG5vTgrnj3RXFjDHqOfWJmHaPhtyxsBNxN0ojRGQ
r3IYIFs4Fgx0lNW/LUwOc6gZ85DRbRfdHHTlGUvJQkpfDoo+D9EBrMGTUentAqj+
ZZy5xZrAtT0h042Q2GHw+fxTWxvf8GeUKsyM/LEz7lmRbd6BBvEsP+x/updHXmuK
LN51+fx63oJxfMsKdVUCIjzfE3MvJYgIBM5o8B7m/yG5BAyaClb4Hyt16HrX64mO
7aV2jtmHP4/KaVERXCH2c27DCRRXLJhUWFNUXlhuzw3ueOHSUD9wYgT22UsAqgKa
XoLc8d2VfIHd9BNgW2WytspDoFhvlj8JNApvGvUe2pVWYim3wJsZaQK7RJB043NI
iv/ogSZLW3oRRKMDipCS+tu6KPioSOTIczmUHNEByR/L2hE+DLcdJ0+SOmrhFaqD
TvJOOiUSFivqQ7/HwStYFXTS9Q0Pr+B35zMSaJM38sR2lzEyiA3CTYcFPe+TITYj
ppFfEnO9GSDordHhAdiCjwgWJu5u7iuap0vjb3o3RhVpwj0DNv+7XzOLIwH0SIof
gmsmE3+KK8LwElzV1wAmtrAdC48v801R1p7O5cXyO1mbr4L6Y6v8tsaB1oEXpcTM
3hIFONpuJ6qOSNcmKEJoRnaqOE1PCw5+4oaatd9cGKlPdDsQk+/tV70GptQy0Wa7
QYmXc3MxxiDJCrWqKPa5fZhoHhCQQbagjAfW0XyOkYsohP/3jwR1ObaTi5rnKLP5
Zp/LseVT5xQ7hbBLoh+g6pAHZ0szKzOlifA8+FUpCKAm9ulr1WzD9HD6Pt+7i8rv
Em32AX+dYvkKQjciIQJyl/hMHs4DSe6gAf1s7ziQxgCXqVlx2lTwp9MIFxNpeGsm
bRPQaR3YuASqgATF5djT3DL+D3vEwlsXwRjzOHWI3paBaT+XszD2SsP4FtbbSkev
18yVCkvNB8m2l1ydAZ57Z8CQpOGSQGig6oGuguv0pRRFb9gIag9cePn59CP7lXhj
I9fGiEkkbGhod9TocV3yQfmND+5QGelDlXlQGIhXzEPjyGv9ZeMkHCzAP0gAaaTb
556VU2gSinCR8mkU6Nn7D+5G0JjWaNJGqH1Kxl7AYsCDnp3+uMKS20jfSbvt39TA
j5EStCTZGEWwYVmdiHT4vGbfGzB9kEHC7LogR37YW7kESzU4qFgtwk3cFwR81QV6
2iId6UfAhQFSjosJJRXcGENvv2y/p2grIqqb4n2zTARrk1eCM/2IOHcs0Pa+ZIqb
uts9R+J6OJzHeKX7r6u+Y58lk639jTV5OlUPRzYWoG4g0IwqKxegZ3wSNxGLDQEQ
4vN7157Num7nSXX/6xvQCizRqvoWrx694oLwJc4Rj1kBF39z3fmAQkpfEQ8LWcSh
G0zil3mlRB3NFp5Fbw5v+smWSW5sXx5rjXwnUgDkmR+M3+zluJ0AYaHP4otjMWhN
JrgIAuEWUSrcVnI9dMs3WET6VEBRvAvNK83d6DIqhMTe5kSyU/DUjaDyJ55+Lfus
L4AIMi59lAFGhPRl8jZIX5KuHk4ovqDOHfc5hp6dx6n2/sVDUTUgUT7fZ/8GFA80
KVv0iw82WxN90i44G6hDBwiNe5iYZqEcA26qjBx3q5zezapHg4HbjMQ2yIoN+fEf
kLhBPriKLGVnHrVUomrHTgyyx+qzLh/8a5A+TZp9SbeSIMvGAzlGlWLijGrwlmUD
TamA3DfDU2Ey/SwGg15QFkPEr3GuMNRjEa9sG6m+bFKlTP0GlSGD7m5DRKLtVs/9
/88oTB2CoVGw8l0ObPp2Ju8UF9vE4K92HSwnf5IXcKs4rkl0KNT3tMA4mGiCZFJh
RKGc6cfELAwdnOEdfxTDpzceNRDAhwS3R3cQOAW6XnQCpAecQ3Zk1iV2sbLjuTiX
kAQTyM8YDSa+9c4dsVofDXtfqFLn8Xx0Nr8f3CjD1/BR/dCsDvgsV8TRPfAK7Oje
b3b4+Ka8cgoWuaJrIJVDhf1zY8C6Ci3h0rd9rpll+e7p0qntYrLFb/8OwpcspJeQ
6JKzsrP6nzwoaKSjX1hxv+1mjS1hUQR0tT4tgb+/sTNZotwWScCVSsrEq9F5AywV
ipj8SaV0kInOfd7z35TYX2P8D1rudPc8ZuAYuWFqARyUL5fCC51geHFmOvmPgdyd
AWK4/QsAOdkmWScaUs1OtFjqBNGOxVnCNYlicDKZ9rLv208YfdsXBdM7+2wtpEfT
dy8dvmspWgCW8IiO7UMRf0XVimvb4CWew0US0CLIGkspGIwkScXPyssXv0iprhcN
zHphh6Y5KSZ8+7JJgUznlsC8QGX/JsXFV+wHCmUDzBnYEzVPBhJ8JRQ3e6c3OtDE
9MSNjIrdwnv5LNXcufhQ5KGvAUaVAF0qATApf3c0p5d83qkbsVT6oML0ApAYMxTK
70kkZpeDE7yC+jrZNznikkyvcna67U0cuGK5h/sFSHvQCLxZyo7VssUja+VyR0Z8
zrRt3NM9Sxp0aOb6BJzMkbGb7xdE2I0gXsQfoFSrfyCSLO9oJrn05zHpKdJZbbkF
Jmdf2V28H9C4vFEC6QZ9+KZ/jdj7wAbKIYrwzbOFCiIobOHucTSJJoyrXhyxwGVh
2So5hB8h44D30Nu/17awtQR2T/yrwIOLVHEJk6/6FmOh49YqZuK9eUQYMGoe1AHc
Qzv/563F7tU7qwrYn1dHUzrlyQnvfqT+AwNrha7nnrh1YDZvH9iXBx/oSEOGb5PF
woeuv67kvu/uj9bHr9Sl/JGsFD9bAxLKDc59jLH4TNGBSEROB3vKTzRJVhcdiEHM
afPbl4Ej4CPONPfy8gvuNlTQqyUsIQTM1FmVsHd2RvBJ/PJ4O2jR6JYCgCm25VQh
fgefvABO1DxfYoieTHQn3mFyyNCoN17xxhp2YJpM+nC4Gb7VsdnmXCAwqWNc3YN2
9U/vbtfWszQ6zgaeUzGjQsv0zjT8HByx16B7vvgoC7KE3PTs8i+JXZIiELpHApLg
uLu3YXsEPsQV+0hBgThmy1sRQkNmQs9gSgsQ0M/znJItPiQdeklL/9CxXaMLlTxp
DMxcuzkeVvsUJJGiB5PeyQoRbj3k67DdsUQbKJsuX1+a/Og05O4SM7EmHhHAWrub
FGvq0xmbDbR0P0mG86rfKHNb9WFfXMPy3bmjsJjl4Tt/V0PxZ9kLiasDLKzNcPEt
s+Pjihhl+/u06DS37O5Evbyj8euv+KyObZbMJwbmdZ/K1FKkkGDpiklzvEZEig5b
pwwpNZaks98xbCK6p7VNvmzd944sD0WJOM7AD60vBMgNg+8HlnhbvuJbR3zHSOmB
N20sZYMvYK5wNvJJ8UDuJmyhimyMcGmJpHOKKTD/lw1F0RWYsaOjot2jb0lbX/0P
IxogX90DYHNtHXX0KDTIItk/hS19vPqryiSmm/TP5ZQoWcHwgqE1S/O8p85avdcF
vMhcuIBL5SFx41aUOW//JFBawM3eqiW+rgSUx9/kxsC+KDXNbmKn4EOjz7DFax+Y
ie3sXY/sOUAqE/z9P2cZJ/r9BL1XJRx3tUK67eI5uH4mDTwxBagZypsdgPSSVz2q
e//Jv0YUIiMbVHkO7jLkNiJwGfUfeMvPndEygTlp0Aa500kLZz+qiKGEy/7Ltbxn
9OMO48XQHsXnkWEA3f6oqz68dxKSOn+HyNsmaJWkeH/0W3bme2hBNkZBK2wrcHSY
8y7yyeak3DpFYZSD1vakrTxyvInW20+JE4EinuZm0uvBVLS9KtLxq7YW0HVPTKdi
UAQ2PnPtw6l8pxa09VDDGUjb655fnlvlY/g0X5JxCbto0yJq0Ov8iA/AAm/EKbQq
+gforHutZJQiqaJIESKRxxRlCGPuj6DcjQmpkQqSOuL48piJixUPL+EXjNzxv/Sq
YW53l6cBK0ygYdPawcHsLukLA17JiYsu07nJtc8EBK9FHN8bPXvQk79QBhxhzPQw
Lsat92Gyq6wChS5+NqVa7GuE9YQMRHtOSScmWFWPQanvC0z240mN87Ob7/9gcFVl
QzZkJNdi4DAW6824T+oCsLfkc/2ULNdBkL17uJw9ttNvNtG7G/exx8uJzvqgKmbq
zrpcgxK0dQWRSyTrPgS5e7cbNe8vu/EsaoTmWI25rpfjzFy8y19xkorYPM7unTM4
Js1xAOnm/VycH30ogXZ9UhgiHX7bRVBMhQjdmpJCx9AJMNUoDlwAjn8MhtVLNvxA
DKqf3SzNKMhVMlj1j8xwwUWMctwupzg0uFaqQoiah9APHX0SV/vBaniavMzB7cIs
vM1YPQAkZj4bkTfZKdJ3bvsfa6IXc1hSX5zqWBnqvWku9AJrFDieFvvh9zW0RmSO
hvBylU0/qWOPjgUknqCcma1o53M60l+VFIie9uV85dAwwkcI2p77/YsSx09Jipa+
9xvhcP8FeoayhRB6kKbb4ZGz4rV8jd0CHfWqKdpvVlgtYD8/PZIBYthPGxvsvcp9
cyKjI91hpBg7pl7cZUe3jooOjqxeDWK9+v5YtuvInPKaMdYdle0R3TapuSKvYtJY
u3aXEaiurtXBgmTqCoGnKaM3+YqOoErqz55N9hR5RPXGlRlW3gN5t5k739A4CTmK
s2hZ/nNlr4XHyh7Vy3N9dqsnJLcZIwbnd6WrmTklb6A7GcykGllqEC0KtyVcGWw1
dBGASPdExmsr3OgMaDvvK9Y6DxPWWVIn6GLryDftVDa2FIdfiOR1yll6ubVlZLI4
w+wAkQRE7NUzC9vhuPqtKasNd+Oz0tyrnnNCHuOxL8xAF9GeCbmK4HJzuLRy2cva
OCFah55KyXO5F4mKbOuQkDlwtlOSMMEfhaAnKeLC15DJh8X3QIvBa4eQ4ocLR/n3
W83cHWkBTZ3TwFM4TqsMiR5qoLSg9E9U/1lsHTUqLOLVeGIuVAnpVj//Oxedap2C
xSbtI00zRBvPtmgPlU6UHNmh1rQi16lJE/3m6vaKg5Fynml5vpFegMQIV7LsVoPs
0GxLpo3P71fsYk4wg0+GcUNdB6kquRtu6Cwofm/q7QqJCo9UjQMEB6iNyKl6LbXA
onweXrteN7NnWDqNQ+OVtTWQm9zCssY+iQEEX/k91BZnHnv8kR0F2gBoUb8LAMM/
xVtiCdwlS4Rlz6CRtBBqPvYIvEVafVEp+kthrZQftzDw3CdDWkPbKlYlXI8bHRqk
7M7mOYVHB375IEC9nrca2doYeJIazUzylYhjqXyutv5DjRAYr5o9V4o6PrQDlZhz
yR8FT0OLIxs81qhAWLrSrqLpUZXmhhKNio3Q236R2M+EnNSUhqggPbSU3Cst4iNK
H9KUdX+LHjFdlQTeU5dNI8gHE2lcVV9ZzVhS/lYEf+9DP2CE/MGP0qAm9rFt7E8E
/yumqdUO7mITDFrq8GENCbSltgT+txVGi75g7gwjJMv/b4Nlx4AteVRvIJF6fFWu
3QDTlg5XfD80cJPmeQEngr4YVh8ARelT5m9TTObPjSkdQ5DiuAqmT9Y4IcT7LNZ6
UqR4nRpi+6UKIuSL0QMqvdxIoQ9GUmmWAz1v3bG3dETGhy8C/Zewc/uUVTR3MdGz
b/e5Wo9jIQGuWONQwnT06ccoTYq/xJ8/d7txnGxhUHKda5IJpGDKdFBw4LQgRe5I
4Q3sr+xHtYNvuMvUF3CYMcNEPvNmZuP/IG6kXis+4OSPBdrkkyX4cS9x9c8khGMe
/xF+mRl1Ms8qiNc5DqvwtYe0tKqMkS/yrsTGcQip9N72+3LIQEcMdFEMAgZGTTWL
S3yQmcMJAYDQ3gjQcoJnjGkbmGu1QzR+BUKjMR+eVyj4gLEVHwQ+8wiCcxqfTrbm
Gydh8UM8V0gyC/eVhGvbNV/JUtrX43v2EnvEaBb+P75biqdwyX65ViqePbvQ1ryK
Y1FkkQ9GK0lN6LnnTTqHt9vOubOhbuyunwMDfKLraM1qxktrB1x4gABIY6a9q8pz
+jMwCIUj3m4atybEQpAv2NpNEcpKBhdM3v8wqM0k78ulLMSRn+xK0UfbSq4fiZmc
P2ZutssnA9WYVCGOUkulc7fAhOCXM8R7Xh5UDPI6LYXk5jql0pCyxqNyT0Vk8okP
+FoYGTU5Ud6E1RRZNGD/RUgYtXq5k0NekBTSK4H1J7f95Yp9omrRJrAUsNlBeSTd
vBg1OhHBewEZHx5gBcA+8i0L/3S5hI9kxk5bsuMqcEl4S2+0D/9OihMTYLWjkQyP
KUgnqvAHu74180e2CCsNXkM+YWmFF414OciLUcUcaRtXNUdTm2XppaEj50rsgcll
ZUauUN17KN/L+clkefa2mhAWuBEVWuSoA+5/InH3C3mSh6ivOWiS7r1kT4hny1gH
aBUEgJbi87hVZ5o+zo81jh2GToe+1BVx9CMK1R5nQMFYuU2yiYxGORM7azCDpOzx
wYljai321cuOrL1ej3EliXhXPrL8mSZJ6vnH8X/ueBAQtGPTu6P7acMTLLbLQ3hf
k9lETe5BFom+1nH6d15Ko9AmGsyaptgSU356Xbl0OWwadK9YRgoSayaVig3xFHFy
kGnEgQ8zvh5nsKmeDTsiMW+t/y+IGazHPx6QmU6UpHd1pw32cEgiqm7Em0XiVTPU
bSfID5kyo+7Hkidy+H8a2hZP+XY7byZFjpQBNMIIPnwShTvU/16C5pBzmYHtBmo/
tQm7nxFIY/p7wZMuemT29IFsSm+kql4qLbOgZ86ndxsH5bCw+Xxr4orCe99uCdji
eOEk1bINQxs7pqPToB556ggyscmBwtT8Uv5Wbn8n3iO+dAgVX9TtZzo7HGExwiYp
ZmnpsBd14AEdI0CQHvld5DF0ncZSA2xmphTYhMQ6UczDTHEG6QKhQ/oNgueLFHlZ
8oclcVrLOLxY/4d80vJErYuCRK1vTO47w5D0am8M3rvaZHKp0WL4DFwmeu9RqXMY
x3WRDeNIucmpUfuIAbuqf3+Rd0FeJrk1QOklQi6U0dRsQ4uVQ3NNr72FPaihtg1A
SLLvDdBZM/J3Wc8hYlR1Wn2+8MDe0WuUPaFUqKZbNwfsrjAQeIMq9sD96Zx0On0G
ditggmHIA53QwA1wVzyRB7It373ovlK5nh1qV2Xs5EXoF9fojGATE5++T8BXnefW
peeZi0+fiQBxUg+ueHoWwehC2sbN7pg3wCzM6p24wkdjwSB6HP3P93MXJ5jtb74z
sqx8K+CGc6R77vcavt7aIEkChbWTzfA7C9W+Biifw2YQSh/7GuIhwx97qA3LJxTb
4I8fZrqAvcfpVEnVGqLCE679GXvkXG7aQVxWjwiP37ieITXTuN67Opir/yOAtIIY
j+gq3oy5Y8XICFMEv3n2qp68dFAwHWo8LFu4tHNgb8lV4pHUcLP4o50oibJkXdbP
RJymFc162WYgaCTHhyFOaHvtJvnGFZbtJl4UJ5hKmv1HtONQ3/plaUXk5Pxe5wLw
bN9tTkOlpujSJwtta6CgzsgkSrVRkkCGlRqCFYGB1PXtuM3MAoAHX/eRS5RLqHOj
XW6T+2Dnx3KdjJTAQ+VKotfxuJsYJAlfqEmDLS0b7YH8F3bBFY3ngragFc3Qz8SA
TwwpAeOK0NZOTZar1MqmasKzxnComM82oeU3WwJPeWozNG9F4eQS3U31pOEOSLYh
aMNCYBk8yIgjX2MaIrkE7GhE/UkCsCbzCiXQapmazschvdZvmhVcCn/CmfwKkkXo
5gOH4DEwdk6MZi3mngCooiCxGl32P94ifQXV/6djbEQCS0BKxeumM0kc8k7aN2lu
nMVXTN5LUucF/l8XRlWOwZQr5ylxlUvpvwLqz/iMbsKVlsnuHjWKMPZjqOn7CCDR
V8BrqXvVWTpQ1C4iV/U72Im47redV5JkRPEJrtGnUiZg6TghqdjcUf3aErgIiOOO
pydSgT9fUqIcQDVlQfp7ZTIW7GnEYzvmKHYXq6OW64mEkyCH5pq/tIxBr8rLO/Yg
lI8n4NKY8GNk6kZbQ5eAtC3XYV5uuh4WHpU0xqo1aKuBHgYFglcQ0V7Xij0XGIKf
E3yLqFStAtqQ8NZMn4+nBZqwgLZdiHHckBP2pcLi2weq7JrySadfRUm5cmH+fuLx
MfmLrs8hn1seWwtUZiU6k2OzTsBmej8skIuLjms6TkopLJPQkWbOLM9Q1eqw+oR4
N/qkfyQpNqHlp6npInONPNnUu5HirDuT6AcJhbo+7ETVESQjir36OsZpXfGPNvRa
8Q99njtUCB9EFzXxdnOFLMBouJmUCPfTQ/w8QHm/LliZhzEARXoxnPWDf22u4hgB
S4ai3Xam0CbEE1po12ZpacP+WZpkhtDTPo8tLhRzHBmC8SID9TPOmzyiJKYSMHXI
hFTP2wJRvlKt51HwP5mDClx20Nfqnt+vcD2+3sZQlPX3lLZgKcUY5n2atJeLAQpd
/6BMpfVnXVdBqtCiS4UtpcmIYFK3jT/51QnFmVbY/cAQXWjFKQ0wsFxbToQPXZMN
vEUwEYgJUaTMxg9Y4JVaC8MLDuj0i12OUhqYdCDrN7KPoGDcQO4QbrfEsrQ3EUud
spyntJtzW2iImEbmbU11goM4yWp6vNGsLo9CfkvS0vGqDeL8CnCVUYzNSL0riyYN
VyBM2EGQYSnAmIt9lF/r+LoGStsQhkFMMdtWoCBBasHEhikuBKdQyiA9HgsDACFH
IexRfgaH6e2QZDyvEptfOsnjWM9NSjU2uO0UqtgTiiLTBWqFXBL2tKg1h4aALrS6
DIYhc4UpwHhar87XB3AUb3N/vz7yNoZOLTVpUn82PeXkCFq2KojwxhugOdYRw3RT
zgVOw0JUrrpDQ4q2Y/lzrW+QRk3NL2/fERM3HlN1ndlHG4CXQ+pILtGcuDUqv1vA
6JZ3CmRGSWBJmtm9Cy31FPm1bi01y9WkJKTJL7K/xK4mQaaUgPgX23ht+LdN5cxU
qs4wl9H9X4oqVFRAvKry7TDkuLr2uRUaXD4cDkyj+tWLQtHhInoey6zxivm0k+YB
zNSpx6Vor7Cb6uV+/l3/FbJlI9L1K157Wh6mE23k0Q0D/3qz6IciqkHUTCwwq/Um
XwQ1ZJhwW9atNrcdrxP5nZ4AUXjgBg89J898xI1Uwewy1BkUF1dQYR6gv+dn/tqq
sTxQ5vYd5t3eP7GhS65ynLMBMom4897n+rzz6tcRCjYsBFrngAj1MNfsCRJ3VeuZ
Qrg4RBmUawkgQlegIZJmRAi/wTWGse/KWViYeiUW2bbqVAu01CBGcxODxRdeuCCf
H6TR7JM6/oqc15mPu6nfsXsyz2PsirskMGbU1uUEQoSdRTVcKcb/Q8GWfc8zP5Zj
XqNChXJLbNbr1Q1Wlg3RCe6/yETUBe0J1s/t1z2BNinXxEtKLjn+vW+JMXbm59+p
dueb5Ld7APU0mQasuYT8vbb9kr/D6m8v80owNqZksVlGRfRorOVew7o3b5qAEpRA
Gy59N27yOKILvSFa3HV7fDfqF5on/HfmMcmmoVe7ZngplOrCrJ27xrIDUPMZmeir
5vJ9tTfHV2831G+tlHU+FMBvBzcx4fSgCCvGqdh+J+DyzbhuN/ClLdQfIbsEBx4H
QQoL3u6ni9WjrfWHutINLde1xgrShFhysB4wO6w21ZRYRpftyonKjaXX7h+vJdQe
0qOtszF/8lBTb0kyu2Mmg5GzxxtjGGzy9QOB8cHKeJEi7VhjjBwZFzYRfovnhhKQ
MpwnKqb0Jh1Wb5cj74/QZFgK1vJtFEiwp0oK7xa8lT7bfY5re7HmcW1Jcn1DaHw7
oQqJpksUFqvLGmWG9SkNRR5/FIQWG0Z8hCpFPJDmNvvyCzGkbTWNDiCeLF75Wo37
oyB9mwQmeBk27BmDrU/uJs+Wf7HeaouWncvfJp+xrD5VSkauh4pMNkJg1F18Ihax
hnmaYiFtCMIjTCa45mxCsXGJoLWTWiI92RMpqL7psytkyOx6pF350TePIi8vqC/M
T0ZRdSQ/G9E+6qmd0xx2a/5U3+VJDisD56wx77NXmhq4i1PMsv3ZLux1bqGXPFGa
GSwZ/GpmBHnQtWuRR8lcSNI2wftqo/f82ZjLo6UrCL7p9Pu9hBo0dqZeToo6GxBH
wgWCUtrdHPQfGpZKmkmNzO+POSsHNokPW+17gAvpBMlyJZFeeorjY5RjwyWq5AnC
7POtXlh+OU0JTTfHMbmm1QKZGduZKWEsb+V+j4SsssS4RV/DzCW/VpmpsZoHfGI9
xW5kzkIAqYbJEYERmbAJs58oBRRr9wAPlRlBv/XKaVcOUGi93snJK7XgVonnG4OZ
gleUK54SrY3XsGjBVgMj/yE8eDQBp4J2+Bt1SI+R2uhVPKhNxgpzj4iKyW0oAwWh
hvQXccFahJNhPZpOebnUsHg5laYR+IoIUlv8Ev5Ls4u7tqV73kQ5HIxyHAG3orU+
fedTO4WWDW3pIyr6arGoAs/f3txNf9bImL/dbAKvRS/HyrukDZ06HD8riFRLrliJ
iPezCoLLmFZvunU3NBewPWrceB7oaD4PkMSfa+6M6AmNpZGagkgf/B0708vG0rmu
bfTunAm51KsrycO2KjInPc6yFNVvz6dOUszLYSGzi5JslltypRIaYKDH0jw8F9sV
zt0ATjg+0NbAAoN0Cy0ADN9utiu0g7oTkYjEXIk8cJrwOuID8z5oghRD+LECMmRP
savXJFM2U30paV49jOWRcurkmXe51sDOatkvnBpA1tQamwCA5AqpjmOrxq6igx1D
4Wo5O18eVqQ2IRwBkjK0dYMqTmkSSUh6MX6dbFvELhoywbNr+zyMoPZW9fzVpFIg
ohyFB/UQYFURmcc2WmxMfEL++oIhiPOjP4U9B0mk8VkUPBuf7gDpo3Quq7q8ahCk
6Uc5iBrV4iWonwtZNJ06q+MjX7YEMGyWWMzUYG3YoJcBIb3NjMV0U2GQJRZP9vN5
QQYQ7Ys35cusFFuMLKqaB7Kvu0L4Mwm66Y/H9QXTdStytx3/EkKVXgqbwH1JzLlJ
3aQEZ2VDsXlbVBgpkloJAlKCdtwoyYs9kNZogTfbqTPoGg3wRyXhjYfg/Iu18X/k
zp/OeYO0clcFBtBXM+y+TlEx0ck+tXsIE5WRNC5TXzZxfFixC9opwKsEZFSC7lhM
Lq9xWkFu3MEafKaBNribw+84BsxQ1adfdn3us7prWlPgW6GJxG5fsE5KUnS8wlss
HGOHySnLGpXiomP7Qt96j4/xQN56zeUL8ejQnoUVZdh/yRJsLYy3mSMkgN/+cLKK
J4OfJDNzguCoD4yrQZW/7ZceGgQWJ5u8Wi0Hgkb0ZSW7Pkt5SAy5Hy9q80zN8PfL
8HRyyRsocVvJEs1sDqE5XRzBOWHiYO2bqCXAIydEKyk34CT1CPjhFGl18x1Lbx1l
R605XKWpwsHQFBAFUSCTPmAXcwdqok2uJ9jWXbIJcc7bK+ZrGKA95/Sq5cmaX4rr
zst0PMDm8Rr0aqRGbXdQC1JLaxTEw5l2FGblFPDtL6I3CQ8GRO4rans1KK1tJwk/
8ZRD+Xk/0hdhtrE3Q0PuoUx1R0orhT1aEh/iVH48RmE+os0aIQa/zomsJkMJzL6b
4NL+EsoIa8/ugdqfig9K0deO5RtQ2d9tmRatMjbRRKnqxbdgUva4I1JGFMq9Zro9
h6mKUvpDDNUu9vhqXi0I2lGnuJ5BcJnLcfpOjoUAVb6LcEcy6pTuuYj6FmDiYRoY
/cFGej6e/ile978sdfR2G9N5aDs2MiDZa06qO5i0NH0a8JHqQPZ1BXaZEuFhQD25
Vqer82dcYjKdb6RM6GK1HuBCWBZL8frx2Wef21Dw6jgQ8uKT7/j1L8xmCwkAj6wt
jEEhQZQWaYbfH/9C1EKIT4oNox0r4M40PK0KI6C3z7hRUnODc+pItHxsmFm78dqz
amHSTNtikiKAkGpp8EMG+suqIX4ga1nZsj2tYbGZyOSX2HTqP7TKyKNhZYFLt0Co
Rzx9oG1NCFqY/tLUs75OoWEm242PKh+2My6azbqaHkqVc/bZqLN80705g1/Hapjf
fjEruztDD5hzSg/P2lt+v8agTaKd9VLjvZf/vTw+Q4NpC5a0rHs3beY3uOaDHUs5
IEAWF6wFpoRAuXACp2ge2TsOvm3hs1lH3dkD+OBXEVzW0T0+dbaiLrqO9XOvPBWs
/T+8OjOdn4SkYviRECLxJ3mzdCOBwmKsQ6++2PsExDh7CIIyUdq7fXNNIzxzhRqY
eyg1uYd68o+YVGoGSPuVr3M8b8n276CBBboFJT+K5hg2rJce2wGHI5buzCxRup/Y
oR0wBZg8JWDhwpznZb74WMDAG0YK+WPkWK2dBuEZisiQwbeNchfjV/IvERBdYLb1
gqhLX8w87vupmzouytSPlh19Y+VB7QlO2bgucoJ2ilAnx/tyTh6i2nV1SKLHJk9z
ZPAcBS1hYOupKyDvPKBY7RO1T6enc4HPpXkfbSP1V2/x4vpieo4kSMEyXO3Z6bIu
0RD+YMxn/guW7oANQzM6LV8G4QwzSLdty5iUcY2SL365YJec4shDPCx8jH0MLO8t
4SU4TIBTgmbxHUz0ckiREBUkNg5h8zJm4SVDVZHFuoEnC7eQJTIqOGnTAcV8Xg79
0Gx6WD21VzmAFw7HCQQJsdw5bRvTTWjwJdVzuS6fzOcC17zywW7FrVRKspz9mzeB
b5H09FlNGi5gKmGuu8kWYNn5cuVAAh2UgTfu15qXqqaKCmFG1pX0uezG2xjKjyoQ
Y59DD3KkMlSjlckx8OiLcA1/VKkL4Hq58KBAjOrWbbAeahneAih4cpSFbS5Xvf3k
k/l5z7kMHPQUPiH8Lf4Drd1WUZCtx7XPDX31RikuQ6SDjq6LiwJHZVbJOSEaHc+J
MpCz+7Pf2oDl6tuEt14B14BDtL/kO8Ja32lL8SjU7O8i7lCKtosGFig1Wr/AI/HN
kdBuewmz6OVPW8Qe52NfsBfReZGpQiTH50Z5nzSnykW4I2M/7zVksSWvoaxac/TG
iSvBaC3dM+HFiLLBhlpujnY5E5QkItHJSgw7Ln42DOB/zqsEaijoJmogKSbpSElC
WI96CQUwmTNzwurrt/5IpZmqPwXrUZbX0GNawkz1fYgiHCHBwe/i9rbPD88TpeUl
E4KMoxJ0aeuV+lhpKtIirfwWX+Rdbt4nlk+BxZUh68QJ+LaHSCuuuz1q10bcKKKw
efykKYyrT7K6cK0a0vex5MI/hEenYRuyKHmV1QInAlCKHy4+zv2bXjzPwg+SjHSy
EaJIPn/deGY9OVcEnc1QHr5vYnDvpKtrlQe5wcNgGF/w1kcO6krappHlJg+3cQkg
DZdgEIz+3r6OOIXzA693z9AI9trhNxxCxT1+bonXvhX+73T4RdDBgim8mw6eas0k
MSYJUzv5nbEJnlHKG/PEOd0wn4dS4NP/W3lJPerKAGqgXoZBfHVenIJXu96W8VX8
OdsZQcra4h4QYFKp/Fv7irqk06bEX/7o+g2vkP0xQZ5ho9G4rsoiTAbHdY1rYpyU
FdMWxr00BWUUtNhE9+AiiwmlkAaelk5STR3DJbGcMKXI1e6jKyqvuKllF7K6c0iy
Xc3yVObLSKHvoJhR6yti4ZSijPl5rwX60Cwxff+QHRpsDlX9kJxiBWXFntHkSbQ2
N+4izJX4GsiLbgf6S4s75XW1EQmSUz82h4eS/VHM0EYED/pCJ0v/CoNzriWhf4bC
ZcTqhgdZghzwfG1v61lK0wtE1U8P2eFrYlT4mSrAkKN741FT3G4mYScLU/RQCOpg
pq/9mu5H9hsOym3kBzoJmleUaRU9tdRNp6Z50m2PFPkI/13xyMTshLC2TufTBk0p
b5yADkqjZ8EEMAAR0GuX9WcdRgFrpHPgHGHLyXahk+8luedwuGcjptfzWQ8mU4xf
K5OlJ8e9OK/4c7z//Ohd1WFFhIIeHkGhnif682uTAcW7tycrDAPKkoE1jwk01GJr
WJPQCKhk4mNo1O3d05p5nNUTZoYmDPsQWSUO8J5ehd7yeAKjIPzMqU0t+dl/Phce
2HQMbLaKnQrf+a7hAcvGh5WdK2+KPTHDa9vz1sddrWV20XzK4vJzz62U/lcODZVT
Chie+c2ldgPjmA6gbep8vl23WH3xnsAU61n4f9Jwj8Vw6+QHEkBtyIjvDme/fxpG
LadcrIu9zBNIbfzI05JRFZqyMX0hn/5Fcd9x98Dd3Zj35sIS82yBpR5JfY160llZ
RVZmRChTP+l8UheD15Ao7iz1hBhcHAsWfiumsD8eRXwCg5nKeiIxXyizeVg3kWZY
FExC+VJOAhoi+EiT8vNLIiw7wShP3WtOiK4GysXkKEyeulE2MXLpqgQ+vUlYxTmr
HgUB0vkv7SwViPt6MWOaRseQkGqI/RngckxuxoCr8kIZTE6fdgn2z1FHCb8OEV8B
qNywsb47aNucjFXjo9TKRiLmZxwAe4qhsavxstziI0wAAa58Vo3BiBrkS4PuPhLo
4ikK3qhsfmaAhFBDDGLJsCI8Me4jEqHMGEf1wpXdudiyDCumJIDwnEtL8+6oa9s8
88bT7CMUdkRLUr5prb3h27/ny/OXslZzdPS1tlov3fIhL9PvV75ChO7DL9MDEGOE
J7aNwjqbzWgQPbenu2H/GIWCbvKhXGJgrcHnOhEUzdwrA74YKLqSR77cXMvDey7Y
RxbrPiNhooiUEJ8hgdOLk8w20lH2VmqnpejAJSj2lt/IWRbYUsmMVc9Lzls2p/eR
QkSY/cd5Wd6lJma8/PZPJlE7rMlkWuvnRbA/0SGeqTFJ/LavpG1FgnYmtT9zTKo8
gZA3y3yLDcx+iV9O4JZnNuXS47fqa1K+32OE8YiKkIyglx3NyEgQTVnRFNQUMzAM
rOck1tGE/Q64F1USab31D3e0NuihulhjxTYu7S0iDDQYAQurRUyUsqj6nLguzXQq
rAdS1rBKo52V87KBxre0VNXLSh8aKy+KwGDssDs5PGnUelwxgqtbL9B6JMT1hJZB
AA2rS9ZvjbOoWbSjbqxHoAhf98WltD6Py+80wjXNW+9GC1npkq6Ylis3uT+7Kgpr
hRjn5wQ5NBz972w+ZppSDU90hcv37Knl0DHbhY6iutxuOqp0QkJvf3GyG0cw9wQz
p2L2FcMSPG1HkHpX0xNtzeccp1ln+H2C4I0inzlxIPZijs1PiEqO0Qa/EXVXXENa
s3dGzIGabUL/SdP+EFg+Lze/B87Hja76wezfdiPjgfO2i0Fe+C1meZJfIcUTbyCi
OSuBZeGoxUFX4tNTdG+FM9Io3qBHHRBNRfOzYmbgoL2+62o5elYG5jLmjNGwlRr+
1YirNBJYGXG/q1ebvx/hxsLX7es9P8oIfSyY0uG6ZfoAa3jPt5jiDFKpwx5/J6jy
dTA8a5jlhj6JflBszDZ9Nxu43t9C7xkkdwvekxd3xa0Dgp3wYsnkKA2gr7NZ9mhP
N2/u53oH2a1XS/2qSnklhQtUqBhNREcdFE3ifVIpHh+SP+ayABsXrZdkRqDVxaeB
aTn+3+P4kMXZzOtZ8CAPuJxHePk3Ft9lcpUVZ3lx+stDfDxqrj6++4OZY2CvFxOh
3N0bfR2NDOdDYk267nJDoOjJ17epXVe7myYMaRZmGkC2ylq9j3JjVaWWP03Ms7Fm
gdSXR62xLC7x7IeI8mwc1DDjzwMWYmgodC62KMzAsozcuhGmWd3dikr/NuT6FY/G
2np4ZH5UlWjcMcWJHybN70xXvRFl4p12/Fl2PBwUW7dmXlFrQe44dPujniKJPCrl
36TpEDr43qxOWT4MmvwidM3qy1fO5trowGRbByKKPw/XdZSz9u5/z4jGQdwCzA+N
6mU6MZYFhv8PR36xp/OtxrT5VUzCUwoodgk8eAV3KvMyDfzrCwNyt7JVC3txDsoW
8/ENcYSVF7ncJXWGE4aKLMBmJM10mMjKzDbTREghmxNjZU/r0JEg6wpgfn2y0Cs4
kDXYq2zn0kuFmDZ082QGW+X8g6bwGIM+zgtO41yLyg7WUtrKyNY/7zUM/lRaRs8W
NWCd9JP5ThnFoXvApdyCvDK4c/pwXre+zqHW5ZfHo1Z3PNsVUfxDY2zCxW5OGrKi
8Glr/LHOc3tsZtwNQvwDO4YAo5zWR6TIcgWQpnmLi92XzKZLKJsE1+X50D9V5paL
qRZz54f1rHYbZUzNUBp77y8ZIfHHre1Ef26/VJaeXJLxt9dWZG80Cs2yagCpSYOv
SEhSAcJinRX3CPXOUKw1W7h8ho7IIpZk30Jdx4Bmsnu26au0em/+K1+T/P2MIEE7
FjJSeQWcTeemnL1GLHdLp6vAmmjl0z0By2ND8Ogw+lRyB87W+vDTxNr36B7/2JiS
/o2h9uGA7phX+GWx/VH5ipGstjd36ZUrJiqUcJERacKdMcRkWI3HuOj7Rk2fOUJ4
KiYPu+mIPN4kFbeDseG0q2W21T2KCxkyZd5gJb/3WsiwzX5qCzLDZMcixmgRXXof
P7nSJYzmUNltSRhhXwfNtCdaqVR9K7WHs6C9kACQFhiBRRjZ1hzVnnzOeFisqThA
kLLil3yIFlx3FSi3R0h0/JSYIRfXXVz8Feoa7Cqj3QW7hWwhsmEpWKU+EujfHUPS
QdpvteDObAxP1XfdWo2aluTmapKyfwfv0hwRs4sRT8HydDIaRllumF+SL+rmmsIj
sD6FXkUJYrnYCiNhE+rW8h18aKIheF85hGrHCa6F7T1LMurKg/nLnSGfNVQkp6pu
YJd8XxIbd+NPdHnxPQmYEQ2Z356ULW5n7R0iTCw/AF2pIENOkGlA6qt90OzvnMZE
SsGTib54xzzoFksh0G2oECPxQtoVs9xOY0eSTDbcPMGNcRd8R/eORUvSnGXQnzGQ
f+c/kWE6HOkUV7w1v7OGhMIS8dnkRi8l5c9vFQSFOtsfc9841vHedWXmlSC6WFYR
Gabx9tB1oMZFifFaZSfdtU3Fqj3jETW1+smb981SSz55HO+oXHD2keBf/hHltpuJ
JUqvAaOOsJ66P7xUiXehWVdWNUhOqnPVWI7ujCUYTt3FfmqK4ONHBvnSYrvB/a+v
5pHuh9C9WPYxxSxF7zn4BntXQ8/XfVqL7eUWpw6Eq8fn6HnzBcEmLm+Z93pazgDW
IAqLiQKsueGztQ3xebLUKEch1OLewLtQTLlI0RXW5lc+/uEEnnEVugpSpRIVhiCq
cbxV+H3a0hcUnH9nBnkrG1vmiFRc9ojO0VkdmWtvIzGaLrP+eESZXefQc0wprC15
niSBh6GpqEt1avhHo+fwLSx9d7R0eUhRYLqcZB+GDGUrJ6T8rRKcPtg7SQOuOFNf
TRLVJfQlOcRHSygufFNTShjKt6rZCZW/LAdyXaim1HZ5X+u2EePofhaL/9cS2yuO
JUuGgpChAM5t7sGFbFKd1TrB7fkie3JGFZiIduSUlzmWX1g8x7iNOK09JDgb9y5/
1VWjrHvkmFPaJecZum17+neZLT9BxewrNjeMpU3vgD8oEfO6AkEKpSabthhJMJER
nx4O/06yrbI3d8lUBo88zey8iHF+1BTEI0uA38YgC2eEmkvaBWLPhMqS2n8sMQh1
KCBBvmQk9H15wZzHINMqjVoLIosFktwXKGWlSXmIbXJWZ2hQrQs+BhhLrXbUZoBM
XbB8BV8qneZhXnbrRnTOjM409yxY/6qRk2g7vqrB/fdnZyis+5WIv4w8L+/fqrzT
Gg2+vxTeUVJwgfiqVXKh1dWRyPEwjgzWU4nIfFGCpBFDO298BfQ+M09/DkfVadwO
RFWM6rTghiSs+vlyGOiGwCPs7fNga5ir0c2HXmfNloL70X3JE/CeYMP4NsN6dNcn
Ix/di8LoIK/J5Hg7hXIbV4fw0snkOBKcEzZhrJV+m/JONYWZBYWU1/wgCZeV4dr3
lzG6cm4xggIx9BrsqThCC4jU1/AMqouj9zqCutdQfjRVZYxLlVVpy8wNCqN2DY0O
j1SVKQbmrceV3ffOTvj3YruaPnVzROZSbO/K79z16oUxBsAcX3BZyvnvceceLZ5e
toknhb3nrVsbwXU9VzOXqJRIZL1KOCFk1ZFrdgP9hFcw/If04d8aXSemFl6gRRdB
ex7zWJRzjYsU3TWIhXNZX1gvTEzJ2HV/4UVg/fUOonJl1K4hkCqY06qGthHu2hzX
GY9l13ncVWxCu54iIHLxbe7d01ktb7grqQTljHq/tME2vg/SXonad7Ud7PoyGqaX
X5XysLmJu6dwXqf9Tk5BIveU8pSrUz9SGMKh5ATnQIMeqOxWClvh/9DdWIsugWzO
7E2V25VqPJoGHQRKvS7TE5A3MJMDjOHy8Z19GQACXFvQufkpIJwhpHKygORKLG2Q
aimaFg2FSyBuMLM1pH4ULTYfnwtFhATShXh4VtiebpsZctXeqQEyP7xi6hT1F0VZ
DAWGCzlHRVt3XIsZST8nr5DX5G7T9XHBQTDSPD57JKJ6lf+eQ+bh+lLbE2XLNgnJ
jGrilBXB5X0UPGq37VkI184exbXo7shMO5IZ7Qfk3HQUwF8aCtPaDYU/M+Ll4C5f
JDQCdZGdHXuIrAw2VKuvAoCqJbaz5tOFKM/iq9IReWfEQ7D9hh1vxElktOfH8SBT
UbJs8PtvtmqaDdOYs/lVV9YIdZWKF18FLNV5/vIWD/otmOWqWsQwZXUKTqFF/s/O
hpqJgE9YBqxVm4a+LhgioHtFocMP0GTYBhwHN4JbO6WblEOw6CE7pPT1LmdR7/Pt
uapAAQCFSEHK70hjRCEHtrU9WgXaYLTaHII+jPCtBfyAMyjj1z6gCQF0ssI/316X
ndTjIzw768aAmmSKcNto5W3bPVAd1/i90kPCB2drI7pELjdHD3nITFqqmIpQB7zi
1Q9LRN0qz7vqdslSDFR00nUrGEfU0toOvlwvGx3c1/cTjxWL++NTYejfiLkzhViR
ZJEZpxdc3zGR6qpKzjx9ojTq7q26DEsx5681MPAABZXmgsq1ZCrjeVAOZ9elD1h1
I4FSSKL/4BUW9iiHWz1GCenV9sQRig99r8J/rYmtg8Lu70YRIwyLOUFxkBf2prgB
Bk5t04pWQOJa9nCW1S1LzyhCgn5XMFnsZCZAGN2fxkdksKq47R6TTxkV9dqG/MZe
Preab/SSQNjJtwGdPwX8bRnWDzxVhIjr7vQvLnU3ezskqKTIsqnRkfAzIFSmQvWn
30PgDpDt8+9JSWmyS7H4ZTqkN3xO2cDC6MwNazJHzEaAvYh7FeUYk1dB8GDi7lSZ
RgUzCRtq/WVV5EDYkW8H7nFANvuLkgzTZD5i6Mb3Y6cLKZcKo8VUJp5FfhgKxxae
PdRDm4J7Mq7wfRFta2xZses8oQtKYcvLRaAlMsFIjKmUvDIVL3THwD9f3m3Rg/jZ
eIiWVcz9/bdXwVKoBdkli2oFOyqss9rNMo2Xiqvi9YyoYdVkcWI+amAvlkXnQF1s
VOXrf2GrEc8XluMirGyCl2G6yrEXlYXAVwJn8yBeNXc+qxXoTtvNT7zUME5jULfw
L+3CffNPKBroTIFTuPWOH/mfev1kUO8vXNh2lfVeN9oLMHihzCfWDQ8nA7jHQdUr
UzOQMPyZKGVfe1E5htpAlCSktkw8OoTdPbZ5Xa8k8/aPr2T5qzUThC2/fLRwI943
r4NVl89Lmbqc9GwTWTg26ogzTEc4dKBzuaknrzUykDYPFr+ZrtqiolwFHW3xWpvs
UZ+mUFG6Vrm896TDG7xsscK9xR813ojG516Bw5z3JPQJ8if8XNdiK5Xs3Cwo0KXE
Rm59IkodIw4CMjMj/Kud6Z6HN0wNocLYK82QefItPR63oxshdMARj6Oy5UrFcMeC
dd+UW4AO4M+TxUPD0G9KTvnrJDax3eUf6tALgNDj2WCwWWtl5X07yrFarYUprvYW
ScoJhB1jcitZiHlOLrQ3YrJl2tlu02a2wj3k3ffgNoZzLyLNQrEiFyooiXMisA6r
M83Waol7BEFl6IwzgBo7ibNZQxZ1fNIwCIQ0GtI2Csv38YLb+/0a91uiWIXruZCh
Prwca8EbNbqH4dqHjPFEQATnt/gDzm0LmhRufYS0MScD9zoVQAcoX0l7vhhFrw1S
8tIbXre/4Sp3gKhWM4Ew3G5G4zg/OUPw+T4orSVDZeuW9nVrHGJWYLajpHh4NI2U
gLCritiQQ5no0Z9KI5kXC6Zpq26GSgmFlIVnmoZq+sXOtRnuEjeZ8IRM+kU4d03A
FGva2FNcQaTYsmCzwOHfBc+2dSiW/m6k7St8/u5CCnadonHv8K7A5OWcj70sOyzT
oNGzL1+U8KPOyoxh8+6Rv//kmKEZ9BhhoPJWPlmTz2xmXKOhu5dEcam3w/BZh6uW
LswiTKJoD6sciLt2Z1C05dkq3wys5Na+8SDCTsl+WWI5E3Gsa7xc03DxHvoS/IUw
O6kX60zCBYjWgK5ws5sTAR0tdoecBVbt5WitUcBwLZc4evgJ3Tzrnm5GG3cki4xt
9Gaec7qgc8aWV/IJbhYlgXQFOr/et0oGc9WNUB09R47i9rvT+QkhPTeKT6SK3bZu
kCyrCml6YAxeP+yZJ8z6+wCN6iNIB8JDjqKtYYwHASWA6fCXn+z8cWZa3CVubGrP
Uft/FFYa9oIkptafkcOCcfq44hMRsjh1atmZgWrY1ESaGHbmna7nI1vpqBwKjdEP
upBKbRCQlfxk4FkQ94x+YiaN6xhB43jBrBI2bq7h172IKKsVP/kR4OXTX0KemBd7
vdNiM7KAqHd/TV410k8GoOtF/SaJ2y6AK+MjnbYiSagdiX8eRFmjgp6o0L5bgPBg
r8p+UQ5uZShDR+LMsIznVfw0b5sIgGRq/2QTkfi+WaUK8M49x8am/SQ9NNWFptX/
5/+NRgbPfW0AbYV4+rro1vODNNcINhQ3Qvp4QCNIKenMq8btRes6wwpKz3cG9z9R
mfHcMf86elHbykgifsixjQdf+YTlnzhUFU6Nz103LXJHQGy0W9EeIYBvTR52227X
cpCiq+2gz3s8WmCScZuJt83aCxFu0CNlytCm5flF5LQb0AC6uWH+24+j6cYgAgwj
8Uw14LRy5xy83AqdWNHn7ixoFa/pyt0Zsjf9N7BuMJiwgbxUggOl7CliVR7utMPs
Y00uB2cMUy9TVTKJc3ZrH1IAOZAyl8Y5WA8FE3Mzv3eNdNbkbjJhzfNAWk3NrC38
9DUo49yRY24RIuFvNW92cuisMvqYO7SPIEfgKuXXqj64TbICSL71RcA7PY2+j9IK
m2rbp9oQ0SpGsuzyPRLhbTrjwWrVpXzhrffLrPqYOMaFlAbThtYXt3Ot0iwxsuxo
WOyESKZW7WPGEyUkJTiQiaMe7WT4Xkf0rrQIOH8i6fj8oHZMkEPO4J3IGeuYkuOV
dSmuUoCQYhh3K5/Bt9o3c1/tcGkcJLbPDik1hI3b9K6B8jjmt7JkNLimVBumEb7O
+t9zYTos8TgfG7hk/Fne7cJrVcZye+bCatGhTUvyl5/LXMNtUnhCtXU4bGW1k4XD
nYAkK3yhgYh98ap0rMIRn7yroZGvU8mGq/mq3P8/EJJr8KtBuixMlHPk7SA95k34
rIfjFgEgLa27s+VZtlUHSm6L6WMgtMIBC4cibJn4qT3JsY+1po7LA1PREIcPvYZE
WEBmov5l5jYM41hQhIP4Z2YU0sg1YwVfTRUX3SADYMYTAigy61oEWXmbfMabFDij
rmvfyYeQ3RCcYMcqK12nqFCunnly/5OhwkwLKLW+clK70lIw7jXNAsJQMSDLmJ1d
laFrYRFM70f+oo4USAHTJgY1ZjXmiN0xfyfOuLZKBnXY4PfmbobgKYImx5IDsplq
fU5eIsNrVAGbBn477Ql6T+jwwMK6a26fr2qzkl5WIY/FCaXCtXAqPC2j2RxAFg6g
k/uLLw+j+upYM7uCWeJLFc7lsNnU9yIkQhZK0WlwhyhcJXuAnEv9B89JZfL472Gg
DTbw78KLHSKN+p/fquwUqDzG6J2f5gAH6ALLoqL5LBtxSog70aoagyOu/KN0vfx0
oU07TzVgwWgfzP1D63SWiLOYvmlfzv4gjfm1bGv7Y8exAEkeN4Qd9M3L56Aalycw
Er+p7mTNQxZp37883BsuY58W0A74bpV9Ol8CxqQx6e6sZRBFjYRfo0cZ3worfybs
HM6rdlNUXnUdkGKLdkq9oZ6L8IGXZyhPRcYDprZx4E8nYoayph1X5IAXuwAFlppU
xuNf13sUHP9uJQphtckc/v/VqSeFnmpscuhUaoeaCfzNAbLSYVUPPABl7Yt0vkEJ
4wosfr40zjj1ooV1T5EOHrfUqgy8HIje5kSRnCX8jc5m1K97MgIpa8uXPwrB1aBz
sDUHFb6iEUDEbC3TCBIM+oo2fA9OXEGXzsUfn4s6x8raZkh3BO5+0btVHxpgMf6g
pTO14m2i5potGg9PVNh2yELBuwhjBmemf5bjHyKO5gWmtvIVxE8jDxN999Shb49Y
Z2E8aFvVi7z70qKvqSts0p5Clla5lEjNKz8uYfq8Oipv8g8pN0YlEY26XXhOClU4
lOyXjWZ5el76hx4ImJluWplmEIqmUAViaYLxaDrg3/hmxPbX04KLWpchWCA4lKwk
9QbGo9WAaDp/KvQWFyNQkSFYevmMTOkwaGtrgSGTbmidybcnrCD5103CtskYrkxd
yOstnf5Xll+8w3RXqSlgYGttuzN71s/fl6G8/YR8DHe9aEQ+qPrbgZ4bymdqpyT5
QQ0lSooREvt1YeVvJPmzBGkkT/CmxoKogq5cAf87/DN40a0lfE9jDVhCZH7dKVyy
UGFrv/pjKBmistZpFkaq2fBxny3X1H6QMC9gf7VpGmdxC/UB5Il/hdgIDM8hGVKB
OssvGoT3o+85JUMasK2VoCcKtOxy1V3rTt2NW6isK5QUHY7dhIDNqp3qRXCArMHm
D4A4/1F/aHAUJRRekvfhXqPNyVpoedOqIVSzVDrC5zt0GXcugqgEQySJgUQH6g4t
B8cSRf9THjncwe7Aqv+lfYBMkS+Wnaw4Wz2BJqS0gainDXVFHdpUoaQrt6s54QCP
mg/gcxF0cskqa8X/0Qqeg/qvkkG9Vjfoxz1BDeq+Om22mXFAZrxUSAJ6u8fbCDpf
PVgp64U2B266Xnm3WmSe/LMLLEY/957mNdhnHmm0MVjyXdgW3qaXDuTZt4dO6KLD
V6SZXr1H9m3m/ooElyDTgl2U81OSnylPfTAhpf62ok2Bdkry6qVJ6V0DG1Ft+oUZ
cjNfOJXjyiPFWNU5PJ8id+3E0lhP0llr1f4V8bCacC52ycGOKewASkk/x9P1PXQG
AIoObkjpF4AArF+MMacyQCc7wjm2KSZJTG+DBCxKRRp0qdV8pGQ3HBd5SkOefyQJ
SdNQic+EkUOkCL+y79F8duG96nMCxg3wzIs8X04j7JX47ScLNcTuPLE8KJrgjuyx
4HlI8UJmktvm2wAhGS73hz1AtGMfJnakK+5MeK4i7e33fqZiA+7vL3Kb5Ixhr4W+
zVD30/YBB2wppzlI1LypLQqAa0eK35kd4I27Tb1SIkhOXWtscfqPIL7nXH/vbqlh
d7pVrT0VZ8oskoKSd46+LCm9342GfgsnmPqfHoC3Sfe/959iHkd93FwlvPLbkPKv
0oAA7kikfKQZtuXFlX8EfLrPeNTnL79bpOLYMGNKF/1F1pXXPswu02xsROgNB/eH
L01rTwD1UlM6TH0G4OmaeavxKacKlbcrG+O7OM3tuL1/82WClxt7geIBCrtQAkDK
8xNddv6jx/9gSbF7hcP0MWjAhjKaE+yTv1/pzUgeVoZm++8GwKd0imjL+Hj35L1q
Bal/3SsV0nmCyVQ5khitJpuoLvzseuyCDltJcppe5NcRNo8qSh/HiAdnmd/8OyzZ
9Zp84ky09WHIw06jUvg8zLs407TUvvDk5rRrA956Y/w+KGO7gDN0oWzk1SmucVeV
OOSFKF/5LU9DcVS5C7ki1zt5ZppQRdetXcYmcKYdOIuwnmjT9wF/SBFYUJM384aX
5KObiUYJnIDpYS0iUDKwmsxBbgMttf4yTEPD+pFvdBgJJY7s2nWuiDM4YRYjOdyG
g0NixG1Uf5YNMt6F3oNqF+bW8H53e/Ia1JyDghC/GCqSLWCpZEGyADs5Zr3p3t8r
+DQWQoszUfq1ZTXto6J1+1o8yRHa4y07dExoefkEvLR/vQQLh6ZUpJ6pKqqPEkrB
eBMcJBUPlS+h5sfIN5UE6ze6JxjrmzZG3O2n5jSIdQ61V9PujsA7VXlW+WmmSTA0
FqLROQwu4RTvGOGFhDvdRhuc7upTlQDIvhfyBH7zPSHmy75K1yIGKapqre7jkSst
qodJH33O0SX85E05u3gBU9Mr1Paslq1iKvowX6c47c5++ZZ9qGmMlZ4X0X9qAMmU
1ot2HOBJRee3Qc5YkfvyIjdfidFq/PGYos3MDud2azzo5KZgzxJxUJLjV5RwwmlI
N/bwAn6pHiwRiSasp6ceN8MS2TWkMNTiSJLtjbgau37QtrVVKsOPBudTvC7fCg61
rk0c9hFWcSn1GzgtFGn+YdyfZ0WDE+K8ZZNIrFyKaQTsV5Ft0zuqZNvPd1W5O2Nc
DQB0adcBSWwEBqIgU4HJ/K1aImIs1+TjMh8xz7PXJJXFbRdehQPus4YM30ycjzrB
JX3GXbX4nN2AmrerWD4Xof/IkYJmAKqA/siSBPvY8wJgmcpIKeGJ8hbZ/jd3gvTL
BQS2cQdtUKIcUskpx9e7QdBqB9g6HA0HJul0jPhX8rP4TnJjMw6AIwFj78ENP+iE
rYxc012r+SgzmuqiIqNsjTpRpjHDt0UcDrEy2piFBiZAIziqQbDidhYQfp5vbQ/D
T0Q+3EBUqm1thQ/QGmsX63W+oZzROGarNug47CKiEtA8PwAavVcg48vQjOZPeQzv
vmhi8XLf7fmb2DtqN+ig6qKQlSYQJyOvtZkRgzoRtMzSZ8YcUKHZTWfLZCBNfYka
zQaJSllAebi24H8NnMKA0Ce3yfMYQHDcCkUhYCCEqb0dt+l90Ce5ffMilWdW8jmx
H8Y3uHJAuyTrf6JvLg35AQVoyZgAi4BzcXo1e+Fss8BGpHE/YKkSHnjGt1g4Lj1/
bJvD3p6guP1ndjgwuZCdSEixl0xV8ryoBAsDmGilUwyUBlyoFsjEFnNW9to6xZLk
z5wKhf847zPKA60FO3z6Mrn1UDCOezbGOgDW6zP8D/RyAjwy0D36JFK4p97iTo6T
5FqKBzbUmi5bKfAnZGUuLIXLLLQA3P0ghavhUC3gqOPfAipq4FX1njTJ/geTcEun
/wetVyUNbm/85lOufYMOu52rlfzoKb9XegpPebU9+Hv+BvI+BVr15y3MRz+9VV+k
jFFiN88f2+3gt34fqx245dUMccgz/K1OD2qm29NueVmEUgXm7DwGwGXGwLV0e9D4
dmy0Kimy3XYlBMsBgksW0LcUSSH7FsDu84tIqK2sunS18+IVyudUa2kva7vNQbmy
2Pg1ZWb0BYR+U8qdru4s0PIiQSqdzhselVcM/29i+xXmzihBXJl0a0lwqWzmh0n6
34cQu63aRZPe2CSSkNZsiosqMVGqdtDQW6FLDOw4pIxKkq9leVh42uQkO/4/Qq7i
ZSXVD5SecAuLNgSUqN/wCVDGLx94ezpOXbb3uYOjB/s9Qmf16weNeknOuIW9T6oB
J09gobG/rx3e6YT5+EcL4vzD/VqycKfF4eRHuc9l28uYV1EotYJ6vJB7YPVaTCSx
LFP2cL5Aafnep3cgE+lL3fzv+tR+QYn+16ymhIiiW6CvZ303iv8JtTnXMFETmUEb
QQ+B+QaemsqcKuLoF67BGo0lNFWgWW4hdgDvt3Q+yM46/eoKA2bYGkVCDJ9f7cXC
qqCFJdxI87TQUcBfi/2eZHQC0sQPEV4V4HF/1ztqgwSSP/M3tVgC2OWGqbVICZB0
lnMWVLEARLYxy10uuD+DaOK3SoLyRgRhNVT19AS0y5DHZV8X8nGJLdiuiQ65hySU
I3MgFrwxGtOiO5nOxcK463hJxkytHjuET+Qs4T5bAYVV+wsqisAPyB0AA9qefLDU
7G2gmIme/cyEwfsMF+ZuUxxFRhR8DmHvR2HzK3ITewRkSZOPSFS38306ZQmW1s0r
N2tB5z0t7mfAyC4pfsBGy6nDvT/hy6uAAUZ/4V3TwdSqIV+799w8y+nBB3FhAxBm
9APAjUks9sqOnphvEXcTVvztn/vxtDBMjJxXcFmzaMeFS/4RStsdQEe/N5TKAHnG
eTmqEANxXzVx9BwPUzQYRZjK9AfVk02uhV/LkmbrJh9Tgx7Ye2QwbegXj5rjP/7V
cB3QgHL0Qmt40Bb8aclGcbcwn4KxZfJXDqMGayWvY0JVUzWpRTT8272342GOn+PH
X/PY2QXhwzk+oDWvxDBtyFw7Y+dxYrrzbiPq71v5T1qqB+E93Z/s99uqAAqtb8Mg
eUIhLqc+f3ORavh0IAM2/KunFum6H2XDYjse20ACO+leWS5kPiUr8p3diVI8BwhQ
NGyn8cjeNfhouPBWCsID7q5jOAzfNH/WxD7SK+o49KhyaZPogaibFDBjjC8jEhcB
AIlwszCKqBHxI7HlvVih089Ff0R9KLZ0ZItBE9Y51qy9NWBrIr0KGn6nBumCHKjF
MiuQb1FX9Brt7YG5hoAGQtjEYiNt9cz/yNnygFB66GwEGeYl1+MFe/ShgoNYfQQR
3mEBsbN2PBYT96q7nAtnj34Jh7w07lF2PQedDrmuP3CZnbUTgJwY72zZRvYcPCBX
yQ8kLA9bsl2kjnIzVvzbzkMh91EdA8fAIvvrRRD9/LXa5s5m8PXDSh1EvlFbvFDJ
kkP67BXeZrjfRrVZ+DouFUdOrGp7HZ4yWbZZ9vscyNA6Duk+8j3h1OAXPPL0HndI
gCQlU+dQLTmZ7tLzKi5Ji+Ov911DWqwtjYQKijk9HLHV4Dvjlut9XdaAkdYVGmxY
VRGMyOaZt8VIMCuxmc2shViLZ96JF35ZMBMb23u3BCWwdGRwVLc1Dj8awzZqTSUS
O5Xa+sShwgynDsDNp3dsjMpbAWyw/We8iNBYaqNCYlqXzD3jrJFMtkJyqthhRF7a
nmoNkk1BlTGCcxdov2lv24llEfqnvoUGSMeUSdjgk5tJigk5JWiozcoXRy6MKLOQ
tknDGcblnsECMsRsNTfoy3mCXwLVb555rCAd+buZ2XFpLaA7ZFd0EoL9y17jw5kc
Ef15UZxxjsspwT5KOhNM2obg23XZdpYlKy730Bn3B6FA/GFL8ecUsZRtFimFrrxl
CqGSz1xPD4cPi9M1m9Yt/+ySUq+wqdpwnLrL2UvS4bSGo5sWYK811Pco+Rl52Smp
qAp+NKKLjtO9ughx/Sjb3KuObBcxPXo9sXmxZCiRWbazb8yE6wxeDDD+myjvEpM+
4fTQ8ptMkxSsiYTn7ArW+b1+NTq/qkw1SFR7pOinljg38Rmr3KWjpvCgfBC/WKdf
ntKg6tPnYzMggpcf93G1zHmW9ldPc1r3M276lFk3uQ7Ax4v7BQsE4YWk5Kk2xGSS
5mN/d1wIF6HyoiiZxH0x4BfUaJPMcmAYPrk4cyZwyL6Nbn+KHjkFHwbYaqpPh9RL
Ibi1FkbT7qE4BFCCm8AXX2gf/ItDYKm5Dl2QfRvoUCgjoI3K1rgeiSRqCfRp9gh+
hZIpbGa8jTmKfctFhpMNxUWziM5y8bzO2qMDLNOxtnQe3ef3sGs4xJpwPxbf03I4
+LR9m0l0w5RSYSfyGskCMvLaEBA+ZpB2dcOxejEtFKHzV6Fy450WBvFC14UczGYV
JoeknGZhYGR0nPdwFtb2NvFW4RQf5J0M3OFuOce1BtN0fwlGsNCokUJsGXJYy+Ml
h8haFTd6lb8hnj8DrR3QdJnWWQHaM0CTdrSGqjvTQ+/pTpRUr3VvdSfQ+eArhbFN
HfLer9gw60nVmsJ9slnRiYCqB/n+0fg/gUMcFdqdAIkEPGwaAHaHLieuZzDgAOej
MXDM8GKkkbWc0AaRqmgS3E9WgHPrO1Ra31fbTuLhAYivxYa6HzaHhjPIvb7ZRPJB
XO1LfdJaLcMB4eAD+wy6whMZnN5Ho6iHNE+9zNaaBYqCPjZNV/ZXtSrdmZiRe7oY
oSKzksm2NLE6GKFQnhlivOEGr3TdPIMecNwcnMeNGWkfHjjQkdrqeDHMqhk6W5HO
zP4U2pFneTVrWW5XEFfD6kVvd27Y4BgF82gIG3mGPd4HV9r5hgNd/k0DRBZpgkyr
o+P8GvVqi/z/CRYI6FfCwNHS6TaRVNyZ1uKgpGUR4cH+igm1c/HmO//jbbqklo7h
pbJ46GhnpVzNU4JykxgfpC0usK/40GgIXSsMQK+drA9wMVZHvXBsNFaX7RpZ0HEF
z9DcazNxUiY8jn+pi20ZjEvsoORVOd6+o53vsZmUOseICp2M2EsJq+/uYgj/UJP4
y/XTse7FmIESnQ512/qKrRAUFD8t3bU4QYgtk9SStTZh3nxB9qWZV8OaH8VbqRdy
AmUQ9r3p5hAGL+ZJorOyTaNt73a0NeM6yPmlPwf8zLkGgu1Q68qmLRbku2PhAWcv
m2+17QR9Wk8FvAR69tfVLY7ufvFDiePfuq848m9zQ4OJo9QhtKPRgwb7kVPF7aYz
/kRHxCGFmTcFQZYBGLufq24Tw34JmpLDyFHWG/LOo0W9yoHKniN2AaxXtuVQczzg
F43Ir1Nc5rHho/w9r3HqHGhjrj8fAakYWhhPINvUUxYgh8dHsar676dyLcYZf6xK
GNMJ+GiBhJAIo0e6UyKLD0tIjoUJjnm4CWQZWLAb/LRIFy5ly73xVNS/ahR6yK08
VpgoX94rUjiPQA9nYby63dXu4NOggiEaz0rHXVYvIizkbgVpKW8Ebdcuz2bK7Ie1
6AAbjNFPbt1ROzkTi/AEmAy47Y9AJD120dCC/KkKA0PnZfUXXhu0+TVbQd5sDxrB
5/a6/HdbEpNaVnokXPpi018Y76qTn7Okase5IU3UM8uDc+vUFSYiYoqXRuuJf6FQ
ZwqSLeUZpBIHAGCKNB2mCLFtcc2otURtg27pHSlC6BDg1QtBdeNDA0URbZcxwTRO
x7o9HeNYe+3StuPymrwj3jTv3QX7S+555ehzzkfJCl53+SzjxfaCCLhrbAfhbdw7
ZyjB96E+UUkmmV3l8aNXyxcRvPVCWxr8t7yxU6NByrFPYS+4TJTmqzDG7i1HHWNG
Hc7oTHj/Mgxx32IqoWN828USCnwPxFdzZKtMwvLwjigQgg94Dvio003/0Ok7zLuG
4raN7ntTsxluv71mTWChkgf4OWdAx12ljJqjABGgbWrEIKECK41uMJyd3OwOwX/H
bgrk4j8Cf0aTPzIfFz1NwqwfKRAUcV5KaTMClDc9v16c4hv5PIAnajb24L4JX5Eq
ij/Tub2I18MIlDH9RmHBH3rOTXUvdz9S44F1okegL6EobsapUkkTfnKGN3j71mQ+
M5L/T8CFoKqPg3RltfXd8UyPF0f61XM9WlIEvYWPFB9cSXmC3fLQYfh6Rb6af3Ae
i/tHzfyhz19DnQqqQ9WadxbQybsHiQ6UQ5jom0FhXwSd7LXP5CE3bhE51NdhFSXl
U6irQCbr41GPziYuw7uVgYGarzHT3bzR3eoQdMQzccZJbV8z5pWooFBD5VT0OYLi
hAs+CPxvTGWWjgYn3LfSjdF9iuX++FbH8KXcwDW6oiexfxazyfow3HUAEaOON+pc
TWWfnushDXltR8Os09bvBGzaOfUnylEjskyUZjH+axe3BiaXGx6WTzRAzXNSueJu
utVNdtMfVo9uZsLkb6ImvZqfBHKzz+gLG94TVlsRAVT1FGeb+lxq2D139Sg8wzM6
HOvtup2d7NKxmqPEbypgzyMQmCCbbhWjrePc7/nJR7iSoNBs0X2xaULX7WyjnqLJ
VReNxWOkL6TkY7+m7O8Wtp1yMsJdEBP953XolyRBND9QbCieeFfBK3b/IQfNgdwQ
xPXyO5il3s+0eaRx5u6XaFwAJ/I4OLWjcWeSrm4JhHedW8v7RKui0wxo1ooT8fLT
apSFTtW4ixAO5dUfdEMQi5Eaq1Dee2Md0Bd5jIZKHZ9cssaIfKHVgjgub+Yk8FbT
j3HwLORGbE4RyRNWeFoonbNRP4dYzq4IcKU2Ls9wexhlOVvUbKyuSbetVCVxpnQu
n+EsOxO0ukeEP7OczrYyojy/qM0sCqf5KWhxnl1BnS85P9Rnj1RDmXHC6QdAM/MG
4Gv3aMl+fwLNaNa9wiKGOQLPAZfYFTcyhvqYye5M9Y6sTBwRfzrT1XN+2N0PIAQI
3DcYEl95kQS95/D1e/AiH1PTsIgRA2myCUTrzVrWYGq+/UOPzcKY+dKj7JRcbQP9
FdbJ9uEpEVf2TjlG2g5VrM+zt2VV6ypr4g+Q2062d+tQC5FpMs8/pe+nO9bbgHJV
SjhkQQa2SSA0KG+BXZKRtOI7kfAKGELiOLmVDHORmsUCXo+SPtlARqhmpr36s2zl
2qBI1etvfZHcXScPa7VEN2IhAi3YPfeAWRTwZ36YDKcPdEm5CLFU2jTdaRjBdfIM
5VpjwPdM96Se+92eNwCRbk0B3wzAANeD7Umukt/wWUXcq2OQ+DPI1tMr3Xm26H0R
06rnD6hLoTlXCQAj2QSGGfoFhy+4SiIR12CVwsdX1WXXInyOOVHwDU7h4tLllAp5
ffw9WMOf+kbu1sDzmJAeKG45VoTY1naEvc7jLvlkHpYieOa/Tns2FrpWpP0kvCjW
sTfB6s3iyBYEs3MDPuWbNIe1zsxxk6wm5iBXaAlNGvkbGQTKHRwgvU0H8VImzWC4
zPkN74r8YbFrbmYXuS9F1uU7XiZcIl3gHCckIhCR3dFUL7YDD1AW96tFL7nCl17w
8+12TJT/ivPx1m/YTL+jANr7pRBX2U32UqPwsUFYKcqCMQl03G+rMifdqm0avFMe
DR7O3PJUXNZM5yoqZOFunInT7c9pWsWxsHDiBOQx+ZBrpwY5TrXup044MSyvFMV9
x8kLv4zE3nTeRvaWujxEURDqRRsut6TepwPP4YG0cj1ED1/1AsDTPjrpLNF5SLAn
MehUxE1p38wpjn1rl4E0JEqPLJ76WvNmh1k4A6N1U8JPBaxIMpO4uyIB2AxU3NRJ
tFmhxdnX3pZVOBgU9oGxvjERR0w70uLamEvWBePFqUkBIIWYJxK1WXAhMnepqMSF
AS/cCfDvvwOtT57oEVsYiYXEW7O7rFhuMOVNpjMGbywOe2eS5er8X9DOQXqddvZ8
iP9Yd7+0XInvKJru+jvaQTlV18GuJffPNkPDKcWf5BIz6UX5CHEp/NU4m402J1GM
0cUlSiDV1A2c6GkKdGTOYZRw42697eDw12Y+zzBqdHlDso7ar5J6d/7Y1LTW8UZN
hG/gA+Fkp4XZLcqe/y3MOAKPwoy+qQQV9b1apBdnmmnC2Vvxr3cHSqKyZRVZVnYa
r2phUBMCRgDLWsfNiRG5DXTdXGQw3SCwf2dd5UtAFBxZCF0eF3eyBV00E6/OgXkB
bIXWvMRhcWGRXSTdQo0b3cjLxwpccbayGywsexpC/1tzgHhlVJYuWBQKJDdHWF2L
iZh8yqlbFr+u6vGZTdLQI71/ZAIT1W2Vu0m+R6TQ0gOOvlWouSqM6hZSAvq94h7i
0WZwzSGjZuxn364RwiLQVsNin178Vz7NcG8gbYTJxZeuXKvkeGgj6zOIlSUDR/8T
GWrZE1xl72Wwc3fW0X5s7maqevJfc1LBWWQqgixjUpdCAEJ0H2LSUk+3Iu7a7do8
H0Zl7u3ZvKLz2yA2GpVhVi2ZI+JghzOe2yQkoO7/sF2vGlsH12tPKWIs6k4yIGVL
Nu5DhtZUfS1Zv184bhKfKeZWjs6PcyrB8GC64dAygUpGPRFBaQdVgZ3/pZ9p0lIA
ZBGAEW8FmPa8nU5L6WQp9/M5ZFGKWyolBTEsVgkzAXroV9gPTEfsfueM8A3EUrvp
bqSn//h0VCSHAohDDGrB6D2G+X/XxCo9pQ/5j3tsseSRBOvy3aDvwepjx6eJpdhp
lB1x+Hv66mXOPG9rFIH320G5OIicipFx778BlLLrtLIBzfYWBPt4kjsd6/sbe3zX
D3NCE552Gd+L59XPOnf8wLtoNNznBBJp3tzKXhexU+5IDtQPGVw40kBZtKCMo6b9
kcma00HsbrieWUbQztpKyR4+RHmnc2aaB5qyxtalGhf+HEO4OF6hIfPbsKhE+Aq4
I3kBiGFoItGj4vGNj6aaRIZTUQAHuTQ+iVpoBIfC9yqJDue50gaoVetveytR/hx+
Amipb/NnMmpTzTBEtWFsCgXtYypvS102Cce8l/bnv5AT/fMrlEJa6a+Nb6X8QvEe
qMSfPCM1dbJAk56dEsX147NHgL+wYvy/12yMCZZ+e/tiP6dmIAKaWek6xnymp4XB
qxuCSGM9YjQCL8bFoIZI/qBkXQsUyiyqOxIgu3DbkMVJajLLGkrLYte+RzEMWRpY
p4ON9ekOJOrbEPLHav5f4FNW81zV6fp1fr+gtlp4MRGkl3rCFB41US2kWCPHLsKN
Nmx1wQZSk518YGBIij5x921EeS3BTOg0Qq7awBg/ghrRPyDA//wNZlhHE5HQvvrc
q+WFabRRG+BoCIr/neurPCpYz9qrkEDibDwQEKtYM4Zc1o4vXAstFrBpLx8Ss5UD
9deimLIMLHRNc8ErO4CepqwP7Id0HTaCFhi+knKUslsjBYF+P3IplJ7dSvhnwZOM
x7n9zcvWYE/xy1EOgzTrorihCjs/7bbom+emDNhca3IJCMmONFsTY2aejxXNIEB/
Py7rB3VkLhKiq6r6/8iCifk0Z7ZVPhbMZPXV6ZWMpqpUWCmWyzpW1EGnqVPdxPjY
lBgGGvKx6HQBDGmRlLQcXpfDdV6KBr5Fkg8VWHEYhfEhEfk8Sy6tP5p489wEpx41
LbqvPONQ1z64Ndkn4iUZL/GvRUvVYpVekl9BHUYdeWduxcC6gN5zeEONmHW+qfGK
eZ7mWJNMEUEb6yntla09srJJQ5OULnmDvCi7QhDeu8qQLeNIKTydX4+VZa2yj1ya
Knk+MCNvHIdHEPFINvL6FdI5jxclZtykf7vahx+8mXpLSITmYrMIW/bVOnTQ1dCH
5lER1HcXJMy0iz4sXXfWDmIqWpPiUtHkIBIJqIs6Juu6aG128Lwi89307zW/sBP4
THATHSeGcPEuJODx9XLI6oCsMoigI45o89FdUMgul4vvf7muvSEsc+G/ugC2IBR8
xvVFp4nIju/KJ96Eeu0bjyGV/0ZI+72iLgnTmw8VPA13w/NRJZ1Jifd0ZWtHmioF
lsR/EiYbcxMFalZv0DqCjaYfVUoOjVg+1C9QAyL27uYqZzjVC8fHG15I+pdYFpE7
KJMyIIw55+ZP1WY1mIZO7TmZJ6m0zF/bxNjwvJC7xxnBv4qQSf/tH1kDKiArhj+v
90NC9YAXyOjnNtAN500Q1VTb6+OGbFrco9/PFczSEXT276ElfqkiEryqdsvyT75t
H3Jsss6JxMBL10FCZl7hETbmO3WdvNKeOpaJfi4itWPRfM+DycPHUc2tEzKnAoDY
EbLTYHhJ6TJDxhI8UXAlYH3kGk55EhOhkzP0tCunnCbMWoKq1gz8QQWBWtjxNDZY
o2aYQj8daPq5sME/uOWXl8jf5lqWDgl9DJMs4qS7328HGf24tA2tRIAGGkO7TWci
6bbnrulpswjDxBT0ERhNh35F6+DKt29YLYAufmZ6qNXakLetwIh+zLJTA/nfUmvC
GDW0IkpaOfltkzC4K4PSwAzPAw3ggYUmv8hNS8uYQj0RNWOBj3O7eF5duWuwOUnI
ts3eFpWZRnhqxINjiBmD+AWnJDPPsUCI51MsIdgmKYPC1LXZsa0NDDmGSY5Nni9T
SwbQnLu8A3LwLIXtpt8YVKh8LLihipIQVgbRlDDhs79b247BBHRuipf6OHgaBvws
+pkzFNVg/FLjW8RTnC2BeB/Alp0XWFOctgkr2wXFRntoEHoZZ/Xlx0bdhobCA365
OiP7MiuSshwteYP7MxBVUxJK2C2/TP7UosQoYRsTTfwG90uEiGsxz2kxp8YtwWkf
W05XL04db+7fLGjp6B94K6EBzGc/rKqyvgt4Y1TOVdQKXRBO1MpkNJvnzT8nqR73
m4P91Yzbp06I9Hfrd4FpqVJqfhvD89fozmDTs2dyawv+j9Z0Li4pZIswCUDAJtTE
gqkU58ahiPPZ8MBDOeyHsPP68hRLt91U3PtIfnYQu2K3Bz6jD8KvLAAkCYR3svBl
7BAvoUUCOtcxhvlmz8KB4mONFGeJ63my5N+yMpDvPYtPM4/4u9DbFdpufkK0PJ7X
LErMl1LRxRRJJicBdsw2oW7KdxrCWRnC2hgpIbYqjCKj5xbjJklFeR6i9XK13CQJ
oMgLpD9Vg/7WCi6a9aLFxuwKDFlChuw8KaNWq0+HopLEBJ+kz1ETR11XLMue6IqS
yX1tcY+VVRJcgZpIcF2XoA1U5/ZWqJy+ED/ZkmmT7KrXPPgXyrqVbogtnwopTqFr
pHHre/To/GQxjAGeOl0jcp8iFsyOqhBaLKJZyi8mi+25b57DgEXcqdjTEtyaziOZ
xetWA/6IvhQQCR1JDWWlbK7crJU1k4jbouGQwdeKbpTwaUBVlUVLESJdT1Wr5fKj
zx2Ykvr9Nl8ws7p0eeR8Gi2MeNXd3IN0RE227p26wA9MshMwPqzqHg9Q8kcYWnLI
9sn99LiTBHjmGVFJVmoNyOZZVllWGQvaORjLsqmNNvfAoBcjZYKxJ1kCeNtK0RgT
V7dtG0qDAt40gvv3yGl2b4D/boDL3ACksHiLeDdTvtFOks1cQBoa/xZfS3Fpwqv7
gbi6k6AKCndUyKg5QQNPv6jojWd/M/Q9kEV2Sb/25cqXtqqIUEKBvvYJjcZbDoyJ
mM6+fWFKK2jqWVrS2tZBCF7xocp6h03whSVsPhJ8lR+7iMxP1DDOd/3zoKd1MiFk
lg+DV7nkhgKSyxXPV1MFgLLyjZ2YNr68LbRXdIvuM2wF9WCsItu6suAibqSxwx0G
Uys8z3kLWuZZ8G9GFCJGkkYYoi/3YPGrB6QQaxm1ZQRH1YA5Vq2Y4uVTavafGFfI
2SJZSS1ZBwCPOsQEPsUtmckHX3nJTC4HYv7kusZP0sZQfQKK5+yMTYfzm7xY4rcA
HoGQmPsoDjieWRvDQYPfrD01cwjGyu0h/uuJrbZx5M6IxZfYl7LyZZbcWKTLw7Jy
RxJKmTfY+JOj8NZ44gtqqaRZWvNf49w7hFDSWbEHE55FGXXed4vGelQEoa2AgmjG
xIWPczZ10w4aAOeTg+sAwBPPcBftiwE2ru287vn5BNKZRgQomCqjoOinw5dGdmZY
ruCay+2vSdQ+SudnE6chXAPzdMACwRNL8SHkN4lDJp6MgD51ZpZU6bufF36jYhVg
NA99Pw10flssTlfDwiYWoiI28AZC0i9Trq2HX4zSduAaH6VTxB9XfTNHdRvfXEUs
XfmKHyAl6GQvcyH9uKi04gRhSpmrmBWLwWxKF6etd/lSYJDwKTZ090+rHscF6MwD
rg1RZJSb9hwJqHWjCuf3ZJSNE/w/oq7bjUIkYAu27cTOuiar+0EXnH0H9w+233x4
9fXjrgHCCowMvnd1QAKXxz/N+S+eK/gYhzmzo4CkE63EXlkHox3f8QPgy1pX5IsM
IRqrbHzUURjmpjpNmlbzU18CBGmdkdXG77RsTfDmH0jNS4ooBVQSf/53e3dlC4aY
udXNJtVcPv23W+ytHqINwye3LCjmjrH516+0i2sJncd58zTwQygiGb93mtq0zUjw
sm8Wo8PYErBjVbMFvTaXOSRNnKISy+qFD3napBZTvhmwXlq7415qMFmOq26+8obE
4SwcacDriiKDoIjuyjSur6BJaAybLyzmlFea0QqqcB3Nxcur+PUNu9UGj4I24laf
0KXO8ZxZc9NTXuNHPhG6vV3470U/UKzuULDW2Sv8CaavtVy8U6kKqDd64txoOYi/
ME4WBAQXVp1mTrgb43WTWE4msPpzzELokK2+I1xM2HWLhFfF+q7MQ8J1fqcl0ipa
8pK7upG9c7CpczwiNsMsCpMShHyzXS4R+VFecbqzahZvEf8o71vt5NxunySZB4uf
asYUaGpga4FBfq+Fm6VL15FJ5g5MPCX9ALajGF/CAcYu/iCuBMiyW/Oo7fjrVjSm
oKVOQuGSMl9EPQV73Wa8do8V8vOCBvY3ho4TB+/JgVUXX8p5UFOoyDEUiIirVinO
IaEX+QV0WKeD4PjpUkJ9WkLEqzEo7vnK3C5Zh2UUgvQDqnTnB2VozrTmlv8GVr64
yuJIuU+eCZ/mQPkVYd6FkbXvwKK6Wq1Q5XqNGCm68pc25cSCJN90LvM2LeB9ALxM
uL3w7wifhsxF53nZGAa+ZN3S5+uFJny2WYCsM/VHVb4qA6R8uGOvcEqK++iYC+Ex
CMAgsdcglIneGLK0n7dNHIazYWfGS84usXj03etU+7lxA0LoE4Vkf462qoYgxYGO
K/7fMrNto/GblXlecrTJvlq9nKKIK3InXvSEEFfn7bAjEhHY5oPFPjcXa1rR3Xlv
6U+xboKAGlwwHwPQGgiSJKi6DZgq3Ib31dbOMOGFzn40temDG/0MZ3/XdGANO4cr
pwm+Ee399RlyrE69DxGSsKeHcouHeX5B+VDNEJnaGbdTBCIM11gPlhpcFNldwPFW
AiU/aHxs1cNTrheKaswEfE7nU2hBmfE6E+dHIGDpuUgHUl9MaMkShGdSmcpba5Qk
0GyVMFVcfsoszH79+l8xw6UOk9Nz87bgMLYQVUk6d162K7s2vl+SHDv2xPxP438/
Q6V6Rs1PqhADzEv//PtQxC0LNv4MT46x0LhXBiZcFZSP0asCEEWmERMLBkGR82Tk
s+cDXn2k//sk91vvkGvPYUmzZG4q5FLrAc8Zwj2sPvUnhnXR/TGzGGbILsAYTU6Q
R2Yw8IuvOeDd4VyIt4tkg5XuiMCUeHXuLWU+akMKCeGRZ4FFPfk7edD4AO/cT8CI
jHlXG2m0XPNXVG3V1SB5FzAE93gVL5iSNGBy6FNkHpPyY+d0EmhMpTykQj9To01H
xcFxC7SuTgnjTooKDvT10zP8tZVr2bwzkZCq12dIdAXpEdzqKy/PBcFMWTcHXuxx
ri/HsNlKlTdmDC/wR0lXpiMaLki+u61IVRrHWT4W7hDtpdZtc81/YcqtjBtgA/gi
Ydw/6vtJjbQETZwDE8bz0ezdj/taPXtPnmRIU0aZ4ZBki2Ljdxlg+538/RutTgW+
1MwMkIIsQwU6P2FidPjSH2ZnrzUYv6OV4ynW3d4qvYkofLMfb3RtXn+J72LDq2Gh
KlkuvDKsiA6kNk3643xlFBawvXLFgUKFr703EjkA4Yyi05cXVwfKCtEpLPcuhhP8
KQlVrSDbZxTZV0f7N81dKU9kKBvNisByzQ4tUgkAfzb9zNr7d7n76vCq8o27eVfl
5JN+UBnsIlBJhCwo3yGuBVMulCH5g3WW+Y1XYFO0VFb42u81BLcTPHxq3eMmci0b
pz266uuyJlColzflH0yF1ugf1Ys/jeYyxXe8mzLJ3hBAyoXMdGgOyqCsSAyULNRr
148ylGB9+Xr2wwrEQiMphTcaGpr+JXyjg4RfJoM2au5ONNtqy7pGv90UBCbCPzgR
znoV+qkCatGuLfwHEUqeyYYIr3BHwjlrJXnl6knkB80T6u+biVLwXhusjbVU16sC
ukATaEK9okyP18AE8UY0PLPba6czJdPopLXUxjAFHanSpxOX8JDOmhdC4iIqT/Pz
6z7nALm3E5jfurT6Jn60qKppy8BSGC0bjY+sXVGFSO5ihYA7ElncWWV2nllS/Pqa
usfKPc9A7ctaNchLNDf67SQu9D0IK9iycr5KUtQsvK9iheV3pMFfESCKhdzpqmci
jlN4/eie9vHE+W0s8Cojq8CxwA16HLVEXpGSn05KDFabhfCyj8Q8TI47BDkn2J7z
cLCHeO0H08cAm4Dvib/lchF3uxXrXh9n3ezFpU+WnBtrXRWt0TsPh0su0Gjws7Ep
MDiQDf/Y6FR9rJvrY18Ov6C/34cBHKiQUQGzasvN4ASaimYjOprPDRbxNA6+lC0N
O3XBmeObWnddpQrr/P8USQA1Xqo1m6Q7i/YqlAz3qlHLADyNGsKKXk2t+77JbDda
Qmz812nTDAmyDoeNsWzxe9TCznGyfdvoAa8Oqi+pYQnHjKqeSYYuRdfXlG5ykCL/
01bjHN9z+ERsHyQZv4s9Ho5WKLi3Oux8xUf7hqr9q6DtMTEiQ7RBoGDxBS6t/lsw
h7UX9Dw9Fdz0tSKcmJ+k/fyHdGuPjZ35Cds2aSOJwaSLxAW59dvGrDHvaeZJeWMc
rh3iDoeBvUMXsw/mWxAiQ6qvXbK0scbWz1YBVJ2cpT3IwLs/Y1P93UfdtsXEg12m
ZA7Sr3SKdiViommSyIVzNhajWqPkVAFmodh5N/Mviu2FGHx68IJiHXvCjR60bG4L
sM9h9P1j8MomddxhpmXcIVZui1OkMFdKsAkH1vDuYEhw12gLjaLt9dTrwioRNutT
kEwdNweF8ZuGI6kJewybs/d3syh/74ZKSdmQSOyE6w8tddoblJkBjCo4YuIqtraK
41VRLl6rdra2SpMiVET5+FJMTA+iwJETW41yEBDdV3R7akTsUIT+irXDfn+UTTbk
48K9Olf/KcC+ZcPq1XqQy5rVNRS6velz2WEw7mqTUXBvB/LA5Q+/mfqt+KFOmQ+M
JyUeDXsWVpoD7Q4Uoch9Flejd2iYnKb1LCz799BzH28Ay66aK5waC6OD37zompFk
k6H2zK28XUsEzOVaDR3iOz3/RHE4zbM+g33u2Vkz0R7/ZJ9i8f+ABjc3jbmIp3xV
dhGaH+PMWNB0O3mHAxnKddqGyZgCFy7a5idHAwCXEE0msKbfExyhOAvA5Zogo+Zc
Xgd2JnCxgnskN7Zz4AiVPoJguz4wLStuR6LMYhdB1bPDgAal8wph5Ai85ZvpbBdh
KG81+H4sJNpB9NybQGUlLpRcrCqhB0o2ZT9HMvHzW3iKmnkShFZjnRuSSkdQFHwj
W7LRY6RMziuvqQ4UttCnwndr0P+tu11ecoQm28ytLN8E0m48ChX+HKV7mhAbVs1j
QcI50uVSEe/oRV6KOsAK5OruYEAXtxfbAyLjatxkuRxKFi3oCXmgn9o+hAylp1B2
eliZa52DRJ2F3xZvMsRTx+xcmkEVaieIccrs71eAcQ8Kv4KBy1paHx4f/SJeu+L1
RgemCujUjDUeMqENTGQbNC5m4sCN0hxxrTZo1mjRN74KLTgbmnhVHAl60QG2CDN4
PnavF4hy8EB5unLhgFQaxLY7IFZtF+zh9ztWEDIrPDLjimC8w3INZ+0daFd/5DKf
bpWPzV0Yx29BFrxDkW4HFLG0Kox/dGdxcMXo1pg6O8KIV1o/yX9Rs+A4/yJ81+lc
y4i6PrBXOrE9feIGdjdw7Z15xWvQp5bJ3o4JJOgkvUl6xCD9FJERxrA5DRvZW0Z1
oIa9doteFuze57N3BzgU0TPXf2GY02MRwnQhnR+ZkpWbOfyDgIKoexXGXTZBlrEO
SABwY2PWDDNJn1QBzJqVoK80bibIeQXKsOD9nE9BjTPHoVBWO5tZemEVBLCI/qg9
ObVd72dZmXOwwdgRK6hzzrUxcg+BT4g17kGNvEQ1HI3mvXuLGY2q3xZXBECarHq7
AzX4hY2fezbEeoZMF2HO9t8Q/b5l07IK/I/YkT81GAshAJRvCKa5wMZNMDxoK1GK
x4vuHtI4UeSN5uNuya+IaFahLsVPpk1S7OLYFLfxLsE3nOpczf8jZFvysGa2+zpt
YspsS0NCnpiEdwxIjfPXYsDpUiycZBxa/8x5OjjPT0PcyUfnZDh6vbLi4VoxdRDV
aD2yDTZIzjG62ancKtoYx2dBLjsu4cRx0JLiIBp4uq/w0LmCg3PZk6X98vzqlmSk
feuK39JD+Te8Xo6wuMxksemgFEYug0WzFalPCSvRsM+jkaIoSrSoMGWFvLVDNFpl
XVYixoHE4Xd7/JM6sTnJXh+OXQOWvGLJ7+x7X+cNzeS/JJ141KK3nVNL0Oi3nCLx
Kf5+QScPUwDoet2dqaGuqj0ViLoVDuNb+TGOBfcWUK1vCkJepk5z25BfW/FpoIyx
GpP6CsyzWGQaakYT7kYKmpHCf5XW5hS9yhvNGDOFcLvFUOZ394BO2Qhb/CAsxiRq
jQ+cF074AEdob9t1mX8Svf0327f/GxWtm1x5524IoAjazCzRYkS+ziW8andsr3yq
NpZ/D1y1HibmwPuU6wXs+BkQeUgdkEMRa4PIxPycrISPSQB4+k2M6tcBHJ3l3I1L
kCGTQDkjLDcjFs2beyS331GRv2LtQjVtW97eZSXn+veRWwDgSZ9pIq6PxB1rgzcJ
VyEU+Ch3GJexUZ9xJpqWNgZ5lTwJo9UI1EsbfE062JmecaooKTpuItIw2smmaEOX
ENpqqVDsoGYxg2bzBVljk/58x1s/oLkWho5eQK4cfOfHp/iDGVCWhaq/1ns3rYTv
TaquNV+03Z81DTkVSmAO/FmmidgZZyeW9q0DFw8/6fPg+p9yKS4mZoExXilGVsKr
G3S/Vs7TgAm4psz94ltaL3qYm2xQJVwncod2uAy63dGTXaWAGYOGs6VmbMcY82RP
YSXeOmi1cX7c68Vfp/XPhI7ZVGivX7pxBWhJl4I0wRjgAe9+s+sEIR9yIFQoPCVa
Zw01Bu8ZUFZvgMtH6MbB15SeKkmCia4TB5DV/AayFn25QS8B/IzNrSWbqfw0YCVI
CHYEjWTS1L41QQtkzr/ZEH7ynoibsfIvTuOiQKonzV6215BqekjiOXs9zn0YYaiL
1ErCbB+evVRuHk2SGqQCDRjKRFuPSyVoXE5OLe/Uu4SWwLcAo6JjiL+MDfgwbaLj
WhYVPdzVKiWerSV7PnMoM2CsSFliVia8vSUrREnyFvI2DbHPsx9WTn3n4sGv0yg1
YmyTnjrfSs4nSdmNQKzUro5G/zzl6RdtwegJ0QbWpDXkWARZ5hzGQxf7nUwm/Hp6
9+JZ7HZzvW8dGm8+xdlnp46bFTDAwuGT/CLDZ8/kV4CHhLPhGYFOVBUzMo/U9xib
raXyJnZPvKpqgzkH0Fgkx+ufK3oz3k0gqBthSdoRX7W8kh/E0eocRE5ZXiSgQMLM
AO8QQ6eFU+3trd/Q+sVZ7tqt9/GaDimy1ZXEkcNIZ9HzmUs1n2S3tJwQ0roXpery
+go6z8c4o1oNxqySAD98qbqdv58fZqTKBoVu8WJDpGGgMWceH9DptL/1wY9AEzHW
2d+HJ6cF8hcjnJxmgeuPSaczCdiDrIXrELnYoOznKNetTIhFJuuAPsWMuCdsbk0M
Vh/0Gq3FyKa5YFnZh9bLeF8tPKwDtUQR6USLXJtkFvJwbcurAIsqflh81dewaWYO
qiF/pAxobU7Gi9wKLvzs3Mpivn/7ZvFVWkeYXUlIkU0cZDhe3+ZTXaqHHMPQ+OXb
N+otvulN4i+vXShMkYsMYw7orsyrqVL4mZWI/SHxF5tPXydunrnV333smJoLlZ6D
Urbl4jMkxiLzbYecSWqpzGcWCm1sZzhc6ZC0bEwyMmEKacY3l6Bml905yu5GeJ6Y
LO4UMYcR7rMl/iKYRevzABe40KPuq1mQZTVPQvfFVvEGKJNWlIl6LadSfxH4POqV
w6EQ9JrEY60keTAgSNkD077tz84D02vyCd5JZZn3c7nl7fYPNvAOrN2U+vP7mrIe
hegkh9WjoPbbJE7SAc7wRAHv7adJZlRPkZK0LYClgDleyuPjaIIg/yLNq0vYPuQp
x9vE+6f+YawrDsoH4+dadZ/CCOVkDsypa9xYFPo6dQDXU1ohDGcA9tFV8Ee1bRiw
u6rY8cb48PrRHhEXQoSm3VnwVhU32BFpYBX4+mjDedhar+t+UbLDW1rbuVoxQ8bi
RpG8GhNNQfCNEOMNRFah/Fy9Z0cOm4gLCQoSvnIK+oTidQK/7Ic7q0oUorgzVJjZ
0mWO0cGjuHBWhNnfC8dTab8puy+o7BPfdcUmK4EAOpiHPwVdi8AXf2f2HVD+LQUc
BsqHnn0o05+qr1ztLfcHCUlyDNbrV3pMDTs9eFX7sVceq1T1fWQzWhdCCZOva9G7
UqL7BAkp9TzkvwndO0/6rTWCHlD+gr9GgL9xF9uaIf9hzsyn+NDWziVN+VddqI5z
d93T3VKfeAid2f/kFfDh1i1Tlf+K2SHGxcfFjx8+WiqHAaUvBcj4fPAE4bJ4Dl8E
X/VKhkbu0A6vbLUZJ5VpDLCN/tNjQe26OVciz58nM5j74dSWYa4eaC0MF6ZbCJ52
7KhzpocFafRC6HI3TS2tCUT3fRipCXOgU/UFhvMRVupA+uyxgz0ODI3h690wGc4v
4R0ByZ3L6YfSttpeALH27/7EVNwE1uxnLXfgPSdipkomGAr1NgH0mZ7X7e14pxg1
kmmPUa3l9uYwHF4B1ApO7OXHnQAHUMcR8zDWVKUYK1/F7ta/eAL9zVfqEHMbFLsX
MKNjae/oeSHq9ne6PQuefkaZh+I+p4uBYXqpd+ew7TapSQGF8rpARjoRJ/Lg3hXW
/KCO7rp6EIEWg95rH1kSyB+MC7449osQ327+L4pcp3iii9kApvB8BY1or7Ljh8rz
EIPZWyHBAy+cb88K7XYFXSZtENGjQwx85hHETPA6PW0aPqU0B7dfUEK1ayy74By+
Efe7EMvY7r6uN+M0vcJON1/V8YH9/LVsvNZL/Hb9whhiCYvSRn0bPpcfTJYf+Rvq
rN9Gl9xe6EOZpzc8GBbgkP/isJRd23a2T3MbOKbIPo+K5QnTyzhGuPtTjQmGdw/0
etUQhHesVUHNtlQXEGrfoEyb0FcBXZ1TRrVyCEzvBgFjAC3lzucQmvXjtbbqNUS+
YjDu3W9ic+yLZGAtKEuweRD6nMWfOsGlNTOTUStsmj6eqeonb5VjnnABBtafHFBI
h8PaAEWdVMcZzS78aG7aVerCDf61lCpgHOPuY4/lKUsvoyYO90ZtahtVSXV/UVz1
UUJeP2vKpGcwV6w9f8fNbhVwAGFSw8LH9RCFRzJmquocKCqDsYJoYfnXK91qzUaP
0UgcY420ePzQMzNndQw5POCGE7GupuZ79tFjVI8NOgp8+abB/2f1BUOskBzk+G9E
oDw2WA5lLepUfJAq2JD8rT8uNXLWV+qxq44tw/g85zvglunypKRGNA6af00lO9aH
RHSg95wZ2DIiZpZ0M8C26zj9HXpaNFzzC9ZDeXmIs7LnnLImyptlAlwSiMYARVby
nhwPUjj5CCkj2cDNVN3J9O+EGz/Rq3xh5GJQAMTlDZKIfhUOgLZM2VnzjfMUv6DE
EYlf8ivzdQ08cgucBLfrvqehnEaerjOSh/J6g5GsBENuqNDaKFCsDBwGIj/g0LSM
VZ9o7JEBOFP09gml4y7hHd3N9QaHeWh11FJI9DvZ326xLBMZJJsZSY6IGDlyFMT2
/8F4I6jSXRw3y1VGEkEV+81/XvlgRhlXc/fkh+3TF3kztQU06PKxJHpsH0K0X1fz
lt7fQkeRKZgSA9AcQJKivgUYQ1/JgoMWR/0YOsQC/3anm2udfDHM/ZY4ItneDR3o
20b1BeNuxltogYOOlonLFFT3O5EBUfD+N1TljD4O57+Rj3jTiG+r9rIODcDFEdCL
AvW75GHI1Um3SIsDoUbvbNSF/dI4tHRfRbbHxaEj7q0oANz82qCLLBcTv3UNN2mN
WDD10M4ws0lRKcrUTYztHrQTHUIJswbA4aL1mpelMZtLMDz1MOyVFBFuHqNj7V89
C5s8LZSLzpJv003nU0HJE2hBmznYloH3HE/ylTDQNK3gtmPSI9aLf13NsJFIANKQ
yidINMS7+VjAk9z5J3ipaOZwj9OmwzFCO85yl3H7qDSfsTky+2L/5B5YwoQvXjn+
5eP4JNtqWhmCYb3nIKWBAPGf9YOD+9jpQldoumyasSWnR2+gU/TFcXm/kPbpIvdm
vS5GeuJxrt7R3RymLj6lztJLKQXsVyw82hFYlqoNBrwNcfABlcWBeBtvkhbcqrqq
Ba/yocXFOnpr3KGsoFZsY7MnooOe/P3v86wwzCQNr4aDaKmTCBM/D6PTJl2/qcLs
6UexsDqqCuYtccaS3D9CpBzlnZ+NCtljeBnbwFKjaTlNJkexxnjkA052njKLHSaO
gX2sjDI17KS6EYJcbsERSFLFyqijopxfzgMkmDJqh9s+26e92IJFjV/9mhYHVxPi
l8OmsO5y9BkKdsp6feOHNXjac3kqUPGyCWOritCyqhrrS6UXecekFP+kcT/65IKi
3pJoxLNkM4JElXS5NszoHhahDOIYlMHhgTj6gWAbqkHAYMluAmWFg1G4W165LwTi
hslqHS0cndFgpiACE83W6JKte6C0pBJYncwiDgUEC5aJPVsqWnN6eYehjMFuyZlC
8lytGASMmWdh5IkVy3nqpAoWD639vQx4wjJj5fWtCItZ5Nfzktjbf800jofvtA4D
vbQoDVygruc48R1cRaTyoZ4EbRup6cUnoNLhPYkbkQTfCBLIcKft5U2Ia/cCm45x
QyCkAjGchcNbnqRu04mSPgFWVTlvyk6HQRfhn67VJ1+0Zf563iNtoCRsWiD5jo0l
JAjVs3DfGBDO91IUdot4ukxVGgDaUd1v6Q8+9NCdA5kuLgiwYMZ4PhvvAHL+BM/h
3M0TnAjPqzNCHuJtXNnN8TNtQtbSm8Zf3/jo95Vy0iSzSzHCBcgFw0+AgInm0heI
dsMeqn815Bwt6Tv0w8PVSjHjMHIWijitlO7gs3DkdpiAWBFursvaOCqN+JLfG+cg
dwrOiKJ99+gmxDxnXNxB5/0wrHCFUqAd1St3bT0+fagq4LP0u9/mTXIDhrcsqpaG
FMpJMQ687Ps/AG7QL1r3Wu1ChtS4F4p4kfCCBDGd9b/J3WH9yiMIz4GDHVmpaNJm
L+6B1Zr1qPq4G7ywbFMEyixI8hUx/V0Zv0PkNoFuh093Wcx3btncv7wwN8jDVMV5
CvEVdp8CyUkRGmJzz6gHE8JbeQ7AqXqqY7gBYlYeygK8Cdl0GQD1j4LxzRWo49K+
AO0wEzGeTPEFnYQGeZYSrFFUmY2A8iQ7cthjhvCvVwVH4Xs+MCpgc/aNnEyONw9u
eQfO9/JixXyimX1IRDOlWtQnYHgmKDtp063wg1yKLnGhVXGy7d4KzB3fVtem3zmu
Glce1PsrWaEUWDwqa2bfSi2HpU70Yz687NBxV/srVoE5bByeB6KxHiqcWHi4fjbo
e0+TfD6GHx7aqj6v334/0uWbWx7oeAuvIsjR3uOJRp3TGZWJu4CMtyxOqOfk9grE
sCLs8bJ1Rr1RHBnOTwtg5229/kAE4cGa77PalBr9/v0AfGWnDzLZMzOLREhN64Vi
ZkM7tGe4NTaty08qXW8dV7o9ns6SJUDeimFNlcMFwe7AbTLU+lLAJt9Mn0Yt00LC
dJYBLdvQ8/CSy5f7F+xzbQLjnHAxLkUAtt0u4Zlq3+5NUfbmkBmxz0scGoAkqAwO
cEzm/cOFvxWSYBizmeTsIo9vGQhtBaZQpFi+6xLlVszwWAnD0MwOFXAQSD8E9vN/
yUMjC+IKKo4lzfkfpK4/qG964H9/P7EzaDPw9AAU2q2X+xhnNOM9OfXX1nbPfJu5
whkb75DpKoeR7qe7KKrJ6rb8YKcUbk+MdtvCAGPNNDW/HqfH0pDiCnwxiavjfZMI
mOB+Xl92YZNsqh1nhGV16JEnt+4q/2mX/4pAau/p+5iqPLmoIzz1NBeEQhd8YrBm
k2qPtuGT6UrhJG0zME7W6uJa5S/hBfzav2NF+zyZqS6NYWZ69FpvECFcFFBso+vs
MZ6fuur7Wl+uAxRnuj77Bbyrm0ZaFvpwhD/HsYX3KwZBLcjD/LbWi1Mvts3GgNXc
HvghDkBx7YKvn2kwlmSHSiCKZeCilbCqmZiMozqaDipAMGf1e8fawNOfVEIkCxzf
+SwFraYUuvLFnKCFFUnKNDeaA5Qu/TDwylaU6CXaEF/TyCy3qJrC27BfGEIIDFnX
doHDvBWPIfSe9q2nf/L8CvhrkUdKba3kqFjQfcT/nmg2lLNHkfhQsASGlCmEBB8C
dp8N8R8Ywk/afiviDe0t1vhG2mCxkBstPwENCs0+5hXChyDsXZDhxLo5FPR2VtA6
vP8JZjefZ1N56p/CWbCnb85UvntbhDld/ZeivVpDZhmG8/pGRTeR/ba3RSspLXLy
SS1/NpzK9WmeB1zEqQCa6CZlNguL7BG2wcHRMETrkwFFaq2h/hLOS9tJT4OF2Eme
zRBLplYU9FlsF2wljL/SabX4iGJtJPOLCTzSj6gNc0Atdrh2KHAawZ/2XlZYr+wa
ges9PEokAeVGpcQtpre70Ql6pKCZuJoDC3qTK+A+FWSIIW8rOGWp3xHVFXqtuNOk
QBCnIQCx2P5gdKgiEV9Q44sYc0XZfhdNuwY0MoCC9GIMykEr1baRBjVXrjBhYIYr
yXX+5HV08BFgM3uTrCy4DyPU6Qtx76MsboHbv5pKZB/YgBRe7PU7wGfgCJwvLuC1
jaiifeD1M+WucWCDGmJFJssSBbctE0RINVOyuSbU2Kq/QUiCwP97lXTYnYPQC/Yz
m9h2UdUjf7DB/hwM6uzURj1f2qspkgjK4pUm4esW2P2SNVLweX8hLghxUbLVV04h
ymwvfmBgyWr/K8TI/tdua1TxaEyPpIz2JQa8yGlgFmQnu7je11ILNtOTGvsGAZni
/g7GsnegHAfk2xXCoe4UyTjBTF1nkn+j+/Mc1k/Y8J9ZlTyeOaLC3emZRZuq/rIx
gAGX55pLCKFQdFPaKxg4s1LvNWhkJME8ZlUrEwHJi9PsICqGj5WTMPsXHd+LDGfg
OX0lZwHnWQ4xNE0l+TOHj3x0bpl/OyAQnE/UhT9+umGkER6CUpEJ084GyRc8BB1a
zK0K9EaMy5b2QJ+hFlT/I+boNWHt61iX20ICEuWanR1YVjZaswFMLsjqtLEsuX1d
JwA4dlMC40F1JmGI3T7kN6u8rE5Da2dp3u/JApzQZOC+6bTUv29uGPdTTdMLW2WC
+nH/NtxYWTZM82WydP/k50punVGTLBGZtJ2NgYTlmm8sTK6GRLmQEO1bH6xvzbeI
NTJwE4Oy/mrhcyunDdh6hM/ZPkI9uPfZS3t570uVqdBGwPBzj6Hz1CHePHRRj4gS
y4LcI8vOeF/Tujyg4c8+CNAamnqlr9Mjb5KS16QgbTa7xXGH7s8kVg2XnuC240co
aybdbdboe223kyT42VrGcALH1XnYVYgjMURbhGPnpJ8rtl1eUAiygZJZ0JxwUDR6
gqewcvK5TyiF35TuiyeSNa+jD7WkARO4Ega7Xg6VboDL++RPfeLTE93pcX0mkRoj
16gTd40RIMAsJkNgNJwRKA7ICej3KsixVkzhRCmid8A4OacrwB2UT4uZKfEXEh/e
rQMYJJCwHjgK50KSBFBk33qrJXzd5OnIbOhAwohRpY2WN53xUOhA9NurSivpqTvZ
qWBSzD7sxFUAuKSL+DP8usGfiEb52962mg8Nkibf8fCU/BLEho6SYhfr8BJDgNQv
+qUciQL3FTd1/wVLaekB8+q7CGGjtfFWYgkDsrxMddczroOAaZvJL1aeboHNEAmG
1i4hD0kBKHQL8v9Me3EXLPAVtLjwN1aDGfVUfoNrhWG0NouAEtX2Ohzs3annzmne
x0Nrvc8Yuid19AW0Wu6OJtFoUGeW+o75HNvlQgD8j7lnmDjRTWgMfdqbfnjasEek
aS0BgtMUxdtfVnXJg2VH7VSMSww3QTQ6O4IFnqqQ7qKmgWjOZes9eyRkXMKTPBwe
x0cuYfnoCtU9b+9v2fpaII/71izn6WGb/UKRW4keRsYx3xgPKm9nRsuV+lKxHIYF
OmN6MSdJ53iovzMrFBvaOHXYQvOe35l6yfEqUeioAeXcwTf5hMK/w40ioq3LJ9Yk
R5vMnDhE5IV702uIhZFpsik+52KZo4IoRdHktUxhxHZEMFdcauK8dIWNVF5idinW
YBVZZpDAo5tM0ywBTvqOXDorWgtzNLG3YMXR6y0THWRJgTMqdLtJRw0jhL4RZ37e
dJs/GjIPM26Hr15B3F6bcIy9KTGxV/demY94rsKUrPs/VUnHIATnkinF92D83aPH
dI2VMpa3zktRkje6XCadUh/Dg/PSqA5EtiyORu5chfueaE9q3LAxp1CZrPeliP1d
Yf5cVN343wegnwm2BanhhPBwOeUu859Eo7CGywUs2o3vXn79MZNxoxGqJJpc+OMT
LcKg1rN4i8n/wnZ7g0Y9bzeGIxMcylkpTNFl9ripu8KtVSNC4dKFCxJ7o/QNfkfR
Ye9NmwNon8qXuNTKqkBOa7lCBhcHRKMPz1t0oy8X9w7cdXzo1239NhZpLdPsb7wY
da/wiNMXKM7rBxU4BwLGunCFI7VAxh4OKKCg+D4TAX1Xq/nmbTxkYr6EGLbOA5sc
fg2Hg9WLJXAKNHpuTQNXpRLEFbsSa8APpBHxFAhC5k3JY+lbnukwUMN27ugPP++u
E2EFqrSC6dRyKWZOQ8h76ZbpG92A+eSVi8ybUU/kwbKZSptfg6x12UCMYfmmxu7g
q2o+9dyJPxU1J0WVHqJHYoJvXElMbh1cmljPxq4KwJYvi50LLJ8OLH33wVa9Pb66
mlY7Fj/mRljqgReyR7wzUgnooXDlXCnmuyIc4St38QxiUjMef+PXcrZ+TjEMllgJ
MSlP6B/bqGSWZAqpb9HjCOj4O7Znt84ZJK5lZ5tN3jv/02deNQLF6kLILTrV72Ut
R3JC+MEtAhqcp2DWQutjbsd5tPI3ZyP1iHOEwbxUFPuXuj0+a1GZ60E/G/mOXa7p
S0IVOpJNlF25FN1BN2stc4C2IpZ6rRojqlebE4/rytZtNLUxe8V+qBKdxGl9WM2z
jWmKSD5jx/FMvp1XnvSS0BFaOVqBCz+9dmUnQk6eNkb2V2pYgt8ohD2yqEhe0kCa
G5mLGAQl6xtXfcBq8eWlptE3qGASJaiBbsnG1If+oMzHEnD+i5O5kPSYSH9hEWX7
W0XHqFchFM6/HZTvL3a3GwzeptNIDT38LecSK3fWew3Wsc6yIrvbsTP0APu7I1Wk
YESa/+Ig2q/rbWr1RjxgMKFVs+R6dT3lx3h1eI0gyGX7v5ewVdkF4HvJPAq6z/fn
rca8pvduY3+wOuHAD/DIaUWwkrXs4mGinSrgb0dTaczoeguiYyyLto0H/0ExPwxG
1mAHwMSXK7EpLqtcAcszr8YAkNnRINS34SqSusdZpjwTQMePT7EqEnCZFL8DKRyI
56GuYxC4hnC9ADg2DhNo1Y+Knv8A+NN2APf1SVIBUWTAjzwvZR4537kGpFhhTrfN
hFHAlnHL0D6yFRHk7JsIe1DySV6eiJ81/VhXTrd7JBgJtwH8cZpt3Kjk42DNkQNQ
Ww+ni5/U1VaGPHfYacQTOH1WlOCQJvW0irYJKzx0wBtxL09NoZeJqrCMcWCJrR6U
mC+2AIZJ2D4xfNx5yzkUYfDpeeLFuNEMwu1IPrgQPl2VdF7GI4UVQ+plo2vdZXew
qHmUtkRtyI4WSxCGQY0/C/numyPp6YBd50bs5fHy7gmixRno9TWeew4ipXXuQ8wh
p7m/2jXIJ+T2OzJKjw2pLd0lCyt2KPHLj7wfZfJeohMnyoFsUlug3xyVEVvFqEIo
RJjmyz/Ho9QBh4KYEJoxDM3vhJJZzDLq4Lb8hEO7cHxQeX0pGj0WL2iScdXoEQVc
pMcjPapQti3HBkpIx1jUHe6KahsWLP7p6QY6BPHPwbgy0UW4ESa5vWjCLV9fmqDc
uLraw1MRjw4ZKKG9n9L5x6K3YrD+RZU+D0VbS01U84PZIE0wH4t1rV5FGs6pnW50
HBFgxn7WIkLfVEVtOTdcfK5QSCz0823vV02lBjcdW9o8NW8KcnMVzGQC7zJvOi+7
ynqxysXkvQt4/IQ3KX5KPscXEOK/XWaFYmahF03gnCZyBi4w9f2qAwhppIt9TjIt
1+t0HYHwFaQwyHWTLu0hSFkEIZkc/kHGbAqHthEFqTnGJAmr+OvgfPFQ3sHUYucq
XFK1HHyEVqG2NRkTApVx8Z8DEcIUQl6oyssZVWyadHMQOMpHF5wYpsKFkO42YNEA
3WssQtsLGSVcuwv8HTCCV89NKGnUtVx4w6F+tIjc3qyqqOzzYJCMSOhGlUrRWuyX
GlpZoqlryhwNhweDybbq41Puw/aFhlD4ErA94QtaxXdbVNKjOmF8+2ogb9I9MX6Q
hih+ZNIsDyAkXG38mUwrXrlLSSRQncuoMTtF36qqzxm6Azczz7S6A07eyChFXzMS
TaFZSAkbln7eU0YX7x3HySERFxNny5lK7lPyMx7xp4NyOQrEetJ4IGU1Ufc3wFnM
uAQ0ETpotVP3ub8w6ss2mmedzq7vdLB/KCboGgSGj/zsiQV9phxA9uMyY3Ia0HxO
uqh+8Ulb+4+kHncmWaVx3BZYn3+1PPaY4NVDD1ng9bwWhitzmgnlpEJCnqgq3SAu
LGR4z0iPMHr1nZYyupIP/K71Lfq2/g7Umpzs6qM2O41xm9F/YOzP5wGktOr9pYYX
OuLVWVmMwf31aUp6QM+pEdQe8Igx7cGVTJ0NQ13VwvsorEqIQAmAPX5gjCu1D2WJ
e3dxacA3AakX+6TFFnvnydcKNszs6+ehKtCiikM7W8cVrCKPgwXXxe82a0sMwzdD
xdm4IOZfbJR9b9H8OmAG62gWXRZnN1iTt5LLYpqMkSL1T37LbhOat0cEMPHtnAuS
UjW3HMbBCMYIp9RNZcELwB7PN/FPAiN9BkGHXa7s27zWNZOc5K1Ihuvly2UdaWQh
Gfn63/PNQXxVtX/yUcc93bkKOLGp7oQrrYAo+ZztvfeXyAvvTf5TPF/FlGK+qXH6
dGYPlJGUDGZbfD3O9NA0TbALrABHk4qpLxaKm5B8AW9aAIIxm5aUROtP3ITj1VZo
sbV91BYvN77n8t3gDG42d8hVU/WPyrRUXTEdKCcWoydudRSnJy0yX70gIhTW1iZd
8B/PkKefNBzh377oPQlkae1xXeNyRPYDhoaxYr66fLDt4M95nhfR2PFOyj6SUYiT
2Cnz3zfOYqkFeUhvahHQ/PHXUeeBq1nawAnklTF0O1dH9LIfOdLYaSOSaAzLBn8s
Zmvg4bHnhtMMtMjN/OFF2x2ZlxCSFA1UykEhzNR6UU9SzqFX3AIhrEaO2IWtoAXS
uCdfFRsl84g8Nvnoa3E8AlSOq43o1kQbeFgTmpCBNH0o6e6fRkShq/kXI1m7mb34
cwf5hkaL/+TZox/bdqjM2Hb00HBZ5eXgrSWVMc3m7NCYzWsSqieQv9KSBnhsspqo
gpZ2mV4aF9q8YVhnx/Kk/11wRFTdOErfUDT8mzUZcOR94p3isszc71KUKtIFp3ih
yVx02HsDJ1YpQYf7u/QYZm5HRYakS43UXN8Zy50WrqiNcqJBinaPD2fTwuxaPO4v
FEyoNEOeOtPB0REOasx6uWifNJcaJXTzeujazvOjeli46x+sNmuUS5wTu+Rl7me0
NC8zacqVZhJQWwC6WE7WOcvQG9AQBlCU/PhDx51HzkWVNZgIz/+qixzPcwi18Zen
JP7WyJY0FuSkxA4Kw4YuZ5pT5egBM5sUqt6E/6TpSV9m3m1xkthLyhj6qHXuPRl4
qfLEkrh24sKJs4U4kWPzO9K+Fh3PxfcWFn76rr6QuFuYKBP6MSJPndwQIlk17+0C
X/GiqliP1w/gIhYoBvv8Ozt6dMc3+umu28Zw7Dmzefo7M3r87PTIJWwslKrhpHn7
b8A949z5IBixdGDaZZWhQiyNKtZ5Yp7/HhbPzEt1ja+VQTcZjJ2nuawvwXRcFVXG
dI68qBiwfAhwOQqNBw3Rf43V0erbqvL3Nbs9dAXSBVbA6doCqWxEVp1U2Hi7YbFf
X4dA9eeGxjZmkElQ6kDteEk9dH2r9NGqEsiuNO3PY4otDWCjGp2tuAkJOt7xq3Ko
N45WCV/T4fFXwUNQkP+6Wtk5ZOt4bYWa6thPtJNNDuKkS3tCMd+SiE7yUPGo+3G3
wyAlYVHFomD7iYbONSwmSzuW1LGWTJTqPkjtd9aN5Camruzc/XYM5mNjjz0ccthM
6226mlY0cpb+q6qQV0fLgOm5q/4ae5ZH/FpuATlybP5H5IZnY/Ay8LZ6Eru33wbt
LIDyBu8caNc10qrsWzpIM2pZ0dt2PZxSwi0TTK66DAA8hcAZfO8WckpyJm58Ug/A
OCQBvRnbRdLIdpyIzPFa9pna7jWrzEfqiANk95GYcm0PZUrgAzT1TKaHrZqqlzYG
9IOB9mxmOacnLdV1+Bxsi4frWSHlIF7OSXyogNaQFloxR81OWNPWhqwe0CQLs+Gd
TAjC1iKff5ak4Pm3jgwhxIhMv3Wye1EKCwUspD+NgCG7LJ4WWSmmRLAFlP618I8K
ANeANf9EJWJNO4u/0hciKNhZxvVgjkzvnARqULGQKVCJOhxMQqKhyRQCuRwry+/b
JIcoBCcmiIokxsqDdrcxmp9DX0KJIvZXhq8FdcVauoZfsXaLqNGufSlmyiQjDT/o
2HGqW912/FNO96EWNms9GaYm+H7aziXBj5o4dysxaEwBXZrJexF5Zz0wDonDgzWt
InuxWx1gkpx8HOc0nHC5s0Cpv+AJdpwn+FJGaBLdzkFBUemSV1cAPHSib0P2tD9j
lwqyBcl9y4jB5LSM+SfrGN78e77KIOc3vgFiuhY3ZM0eqkArUwSywDhJRAhxYX4v
jAyj2CwQfwmQvvm+NrniWmF+7Olg6WP3NsSUCzarFOEyjW1pudyfN0sbBVeijwX0
wcluNM4NmtEi7b+bk5JR1nCUPCDdhvr3qyQVvSqQs5uQVBdMkkA0BOnYHThZWpC5
gG/ssqJpB7EcVXgpz2fmITTPDRo16MdskHm7bJ8aoxpez96pduykgE62EoMOcXcW
vtJzKENfnes4zN+8EEOfLUikP1bnksNwWJjAvxTeRYGek2CYeOABjRz8RyTl2VJ5
jgNYIkEHuKaZtVJiZtZEiw+brWE8/qIigbQRM+lXL2mY6Y0VhrASCA0wVEuS1agM
3Iy0i4YhU4i4f2UL6yxnHElS1LiKkEBTuMnVvpw+V6omxYpzmzyOjg2mu1qmW22+
d6vWRZd5EayFVGEwc5Q4jjKDO1RQva7eh3PXsFhBTJ7X8lsmU2xnDT4rldWlYq9g
o42+6fIg31mi2gq7S5AllaGwb1BHFsIBJeuVCtyFp73m26ZCg4FkDRiCdYTT14yJ
30aVvYk/deZfppJ/34aapUeMRw8xvyYYCehBvTpyvqWGaWo1sVhV5eAhtu5fwnNX
6+UvrqMAs3IA5RPp4NFojPvvkXK0/2jaRSINC3LB4NEAQZ3VQX/ZXyQ44p9Iq5zQ
5DlqAPcmeX9U4rbe643EJN4nLmFBb12MH3aQuyZwj7GPR6Moj950l8m0Ohon+AZ/
2JfZaCKHbPtz+OSEKmuPIdU0KsylNTnSTJhH5z9KoEKc6gXa+TT6DXlnRVt+ZCIi
1ohnFJsbjuUn37t7a0tQiLEuQvsFTJhqgLRBAzJJPvZXUGffpxNc78L+t30W5dJR
lJFiRPXm8wysL+465n56W3C9QOE1Jl9JNJPNtT+Vfc0ODwkqWv8mLxIiybnG1NCc
l9R7gtXp705QZ1l0LD2EdqG9E+lDENitWAKitrc2ynoNaSBhqDRlXMJFEiWOTAVa
KZmINE4oEtXQZtiIUEQdnBGxzQPe136QJP/QzPrK99oGDiQ8Az2RuFFKziMpEwlR
PBdqTaCX/jfwGDUZqdwIpYkuBUDbbfaDxro2OYQToVaEKoGxjfPEAnKMRuYUg42M
qGOCAPcVWLJveEHBQ1Eacu/Ga4Xu6JQUE7L8HpFfJaxnuHLuxGTdND/BLHTsy4YD
jRW83SZQds+R6W8DXgTrEApdc73OoM7T6V18P0N7tgGdk/XBRLQAa13sAPCnHiCA
t4Q+5Xf1aL+cmc/XsyXLuypUMCv1/Vz/PC64irAtB9eFS7S9QbOZppZHgIrb6fRf
LEIGQwGK8zjO+kp+bnThK6scmm0sIkDEZULveTp+pxDDVMJfAx0lt0lxWkWKB8GS
XiDsvJEmXaRBi1nu0iE4v967kyWYNQVVwvJUHNw19tqULKbUb1rd2n1COny6nhVh
ct0oLgoLEd7aPYgJYRSWozIzensfGkpe2EMKD5uX9j/QYB7MP0AVkUMXmvxbRChG
nDv4LrzqtbZ2fzSUgvD855bEQsKAef4G0FlEgaBnBdEemhK08hE+K9osw39OtAqc
vLnqeO8yxVMGmEZ7SVGc2k351Y9YV4HkHfvEsY4UF/R/Pyg/XJXIFxprGATwsrIJ
L7khwuVWM0mnPo4FDuDNkHbpkLX9Vm+kTf7HssqUXqLMROIrAWiQbnhWiNwIZVDa
8IUs0+TpYSriAS7FCN7fqhVaFXighYLPAXr8eMdT9i62bvCbySpPUka9W15ZQS0g
Tm2sBwlUGq4LsF0t1OJSISIr8YEsF5q9ZRqyBch1MUQf1GBFlCj7oRkKePv6msaD
BPJqp9Sr4L4MOz86U1xE2pUJ1EXCwCOX1Cp1GGkt1G8tEfnzKxu68Q2WQpTrnPDt
Xhp0mtNyCLaIbvF5BAL/qk/GzaUcCpdFcdgY1vhXeowLsVRC1RihCmao+3vC/BJD
cgmijAHCWM+2/eKKozdVyq1GExqDtlDcrKI6WDCS5M3pFe0i0FZSyWQMSLDgu5MY
yBRdDAho1Cp2jupB13ohoB1yVqYEQYLiwNjppgthkzpgfQkhg1z/GQa0CQ6Ww9Sg
3MvF4hUXUu5uNldJmeS7M61qu6ByoqFVG6fQms2BiY9GL4wvHYL+4p5oSQI6hZL+
gIwpOxPHmSivoFmEs7GO5eDdu4fKyR6n5b5AngOn0m3MZ+yHYxNhQGbnNYwFb+Sb
ZYOswd1uhQjeYF9ADMkHqToUwBXJcbax+a9n6DnWek/KXgxH3aDKR05OGDMFlwpR
IZxZi8TrjtD0epcrCXHd0h4GPf3J3u5cxpmJKSVgrLk7H0+Ji/vrCEm9Tz9jjAc6
R07FPX/vAztB3l0IVdfpDzaXGjXxk2RYkPQbpcKdYT/9eOXNPqX+Q+pZSpIrh15C
IMk9pawEeb97jQmx1tQdwHpN+JuDMis2oFmeYfNbXnnWlYBnuvOCBHDaRvfTuzOm
I9XP4HjNKn97xXf4NQOLRnfLQmjQtyiidfl+NMqypS+ukGbzVPXCYafcSe7XIitu
Cn1+nEcVzQkq6jTG259zafqRAPvJMMD6iDWzyMbyutMhNrnPTXb7VjckM3hW1+4A
bynDEL6G9SJy4k5Uff3ZNl7+PeCr8SibBIh48T97dCfYIwuDvj1tHDF167pU0q+y
lNxPE5Ei7+xptWWQTNE7m+w1daUSSP/v0DHHuw/jIhv92YVDuqAjXqNLfYFLBaqA
DElFm26/XZbEt5ugNlm2i132F6iCiutSgEwEbkdjNDuJKzPRJAm47nFqrwig6VfZ
Vj28rVP/MNwMrsl9fzPIezg8YrmrdgC7UONdBj/xnJt1QGmj2i8pCN1Zq1E/qqtF
xT30t98UJ3ubJIC06U6fQWMACk/p1GMH7dwDkaQczakXYrl6bDOZwiFeBTde0q+2
Q5MRkW60fa7ZfFJcebwv5wVG7BGlvzzLNXoi5+t72R53v0qrgtfrGP0mmpCqLYkh
0PhSZIMQtI1J0QJqVxAF9vaSQsz4qBCs1SZ+Hp+t003LD+RfU/juRgzzVUuc6U6K
/ZOJ7kISxZYE7R0pZTkolLIGyVRl3xPBZXanH79VOFSW79P+9oxMRcqcH7GLWkH4
tiT17KIFjkYq+lDjMLKDGxKnewMUClg31HXE/pKhTV9y1wxEeGYdFS8hr+3iezRa
3w3iP54XYffD3ov+t+E5ZqWxCDQAUAGe+8BvouRmAjybbbMnuG9jfaMqH30mvxcO
zwChd5WbmXwgyTq8FCGGAeSghTgi5dQdV4ax2rfdKbZHlhTvoEnRamckua8j+iGQ
ryL8duDb9JSPaAYgGlwFysGweAbiQX6h0Xc7M/O1om5xSi8D8dpy9zHDng9EYHPm
wnKqReDOWgBDqpv30SJtoJGH7zbZgjFIcGFFuHK3LiRQRhnCsLcsqp45BXvwRZzA
KZBvfIuREzLAmPKdzm15LIsALa4+50JYbZ0PfWVHIr2jPOkRsKcrGmD0NE+xVyfl
F5HeuvfjfiDFZ1X45UiFWp1Mn4kN5qqm8yAueb4cUOe4uxmRjpiRO5M2ARI7ZLfI
O5TuLH3p4WgiDciNuCb2FLXD1vsOcjPl0sh5K6doQ358iuqoGzFRSg2CMCrPXfrW
ZYgerriSx0Q/yS+bVfeaj+6Lg334cO9j1xBJ2trcSW8KnYuZ/pCe39+Dga2TQCEC
9tm8aVg+/mEEvRdVA9oM0hvhMSi4QM3hLf5NWDJP/qUisDcd74YXU4oHz2rreSr0
XGesZ0fcPi9dAwFbjwUennFAE6l4FT+Xtn7bhdWBVF0zfUwlzj3kLT+QX6lIoq4Q
x2ZahrSmeXehfqR+3eunWGim7BGoRxTs5asro3wdDg6y6DY89wCcc7klHO+lI9E4
K7m2APr3ps/sR+aPbwBISuePa/AMtRg8yED/G2g3zn64vWsBpTdvEFnRNfKx7o6r
tm0INKyZOrCANFTNw3xnnBIDKGB1AEn351geleHlLv3RFRMI9e8ieRthRxRNm6dm
jO+oqgBbJExqDfV999vurq/qyz45i1sj+1sRXRVaWE+nGYKnehvO5bET4aebcp3m
BP010jmnYFfhRUf+P7NTPDtHc4VXHSE4Yxk7RfJhjwGFQ1NUBZn7t4oQICpXsnVX
BVG0fwGBymGR44tl+XNYowrGQkSSFkaamSW44ahz9BJ+DCiox8GzJFBnPnPJh13C
9uj1/LGVjU5kP5OxSDfNZXRfab7fFRVR56gflyglb0VS39V4IaKFyKAujQJl6PUk
PKNMPJYoxj6jveUCkNfTYj1HufZ3XeHe1QcfXTMQRPJ8dYTgCAIBYqjGEkMaxxuZ
GvwoZp3718nD879G1fZekPBLQWtGQBAseKGOBQ6FzcmNGxe8NU2u3quENv4p7tw+
UOdrWLKZdhXusyt6rg03x0jRu/nX8/3gSp5c8mWipOSewBt3WbOYlvCTehD9ww9Q
10ZcWNxv18y9613XYFAdKPn3O/tbsE6NjGrZjpUPncxKfUCI4a7MtPRAX7R5lQ+k
UqmXLZMl4oM3GfeI1uIhsNEfHIZSWQ6PBGGvHG8AO+5ej+K43OGIOurA76dwvpQU
ysC2kbiwAHgYqZ4sMZjshgVxg4dqTs7mlHwSbHWyOKAOTx5atnjjWkihq0wdIEEG
Znthv1kCW9djHp+MWv7CIabD6R/qRGLW2+RuxIQahIS1pWeKLpLWTQhiGkSyecND
3wAOHDxABmgMyNAYq4lnFbC0Kmcx+CZQJOEpp+RMOAIwMM0ahJ4uUmJ7ustDhlkb
ksgQGHKcx4q94PmIkaYFqKmQS9Njt2FGCWadhfR07QTGQUoUEJmhiyJEx8+cJif7
zbao/NB3Xd9o8Uh4PhDQTh5nyzvw7JbizMUeooeG09FWLe7JRxfSdlhIbm4Quboq
B7dC3EBgcIP96gFN6PR4dY47e2Oc2a9eqY9yz31nwKIXyN72mrg+JN2g0mUsHxou
72sVI5Vn6+Lr4CfIRsQGgCHe2HmA9GXRZVwwgXP5HEA+bjk9ggsqj6Q3QZdScNin
758AhV7k65jgmpALa1lCxDU4UaMERx+CDcEZ5HMMDf2uylqVmsdW/hRdYwqT1Rr8
FngkIkL1XIHKZQqwJJlEgG9wmqVAsOt7KZiN6stIQodna8HYBmdBb2m6S1QgmLEQ
loyaRLYvkEIpiqVrNfAfYu5tie+jQ24AeFbe8f3YfjgCFKnw17XxdGeddzfQ2vwa
n665NGXKVINf+XWYNVu6EgYVfNrsyCrQqgkT7f6DKKbKsR2Wvb7GppjBv1LjtlYb
5J5MFCOQmcjF9mgS1cTa1PYxifPRK5YjwcExAgrv3MlgQcflOmWeyOD+FFaNu9XL
gMERdPepIlGwvBZXMWV3n8sDsNeZ1QCIgvxpgs+G/yVZ9IsLsgTvYDg0GcGzzqzf
1Jp+gho1aJCXjxuIyIMNq5qQFpv2Lqrvp01x3g5vqMgHaPIn3KuAc7qKbSpPoqGR
UcSWdUKxrd9wMBqxoy+byoHTIT6mzuuo+c9Qoym/Hno63lrGohYNNcLbjx152Vb7
LPrsiMGrGx2Zt41nIVH6lswwiK0dGHsK3UjAglMWwBnJdh/9EiB5pB+8uWwh2aWD
NGv1OwcCEWxDx0uUFyFHJjEG7tc0CcE4tcxuUpTSFvLvAGB8HNZA9qJk4S1i+a03
y2fCOU+zPiDTKZ+bu1sgVL7Pkg+E2qsEZiu6wrUXagFHKe8VALGQSWJZBSUDQiGm
wRn8yi9+V0X7Y7l0EvNM8t+YM+qnALaubq8D2exfGM1RvkhabJLNL9C/wBJlnpV2
vDLC087H1t6mHTWINzzlwgITGFskvBxq3PCnq/s5SERMJREAVyIPvnYwmfffUKiT
ONZlKObeEs0oE/ymDbPvFif+GhgQL6Nt3F8nZJ4XY/KBTU/TFMaLyhVNT1r/LXUn
XcUJTKbgnLxT9A1R78EibR8LtKUxykoDaT5NeKDBi1rNs8hR14hGsp+xczaTDbK7
WHWUtkk7PqTofV9rIq9RUqb3kyzQWLZhq0H1+i7dMRYh9Y1B9T8yRDWNN0qg1j/S
ASVVb5hv9V19SdaM0moVGuOcMtksbriLc5fy5cmULzOl+D2kHjOK4gTynP4qr3Nz
Kyvv6tIVKMHCdkO4oGVkoV9NH/DKlE551QkMHXibx3ECtHRcZSnaJTtJJ3uo9YRP
tbv1/5S4WigM9oqD8UoPjMILprTirYl/kCGmNHR7UVXkAqwmkkbseJ+UKPF8wRrw
CKJV7WB7BYChv8nzxhN4iXpgQiYx5z8RZiQsIfpoJkNZYCitn0wdFwWaz5AnoV7d
BSnOoshISKYJm/Whoj8SHTj+FGu3YiXdfeqEMucMgdy11JZvB70+EIc8XyCFTJ7y
hFEMkQH5kw7FvePIRgpq1uSKaKjIPv6Ii+ET64jXHLOfPV3CDW0QkBQAmxoZ/A3n
vPJrFAUlhQ7a0thGgutB0JXEAoZFG7hfsdgtPzTh7OZ+KOmqRk7MWPULf47nz/BS
xeqbOexlPYKgwduXHeUHbmIXnIN7uYhcdaDiF2S36Mme39pvzYuRbXyL77iwn5ZU
d/T/SF5BVkLybORdQ6p2ojhjckg+loGES6UvyOwo68JTRrxt12XRFbjSbzxM3VBJ
7cpceQWRriE6N/SyvtSU31a7rkLXk1p5g3ifMQmSRU/TgkfN06c4zmKJNg6SvEFi
u7N1W/UfJLw30+hztIzSyH3iYwBWfjHHm5q1wLbv43TtsnUXXUTqsfWYSXn2VIDt
Ei8Yp/nou44kztNzF5ll3e621Gof25ORarV0/JZObMesVuosqv3AXZ8s+fh4AmAN
wfItyHz9+NnkEGk2eEow/hR0EguhrnhEAkBXe7dcTsObLuUgkLeRnEJSojhZBvK0
n9DVudMALs+T2VzlMeEO6j1NMN/K5quQz1C1K+mHrGGftWqqZ+5OyZCqe3kIlfbF
jf7uziF/C1odZqgAVhOkql2+BHZoA88TbMgG1Kx/MEUhNxpDzCFG0ANExHdakQ2X
XpXXeZaxw5GBjw4KvLi84wVrH3bgDGNJq2SynQPLNLKUZTYVRyceQmDDGl9m1O55
hnBjC3Yd1xuXXrKJoIS1AfsWZnBoJ9x+4rMAXC+bfHQSFX3RVMXgHZnIb4Qc1TSz
kCsl3RaATtXBVmbVTLO/OdzHywXl0gBViaAxrG6OCe/iWxRn6CRb61L3l4efnaEu
j7HPS+ZmhBTBowFcf+tHIZ7YYgc3XwFnISru/xk7C/80hWMMuIyeYhfa+VPoxzYt
040LqlK4p0DW56l48Q9VDxJmhyv1sRyQSLTpaP8bbrjsdXM3OzAKSRPw1PzFqWbA
r/6JjECEnlWK3WH3wCpRWV/U4ZezB+UsOPNGmMdDUFg1cwqTkwwAZW7DdC7UW9A4
6SM5fJyCYSIGvw5Bg7d1e3k0z7r7Hrr4SpAZTuvL7dyr0rz+Kv1kFH9wZNH2aPm4
oGnw7cpCCnesmmt6CvLEgI0HENFRQTi4qm8mUc6aKz5R6wyFWV+Y8+c9vo9V6zOX
xCNLxgxBuEQ47S8H7iC7MGZ6nImomdoTLp0iwPkZzo+PNkUtwV/1NiMQQMS4cjQJ
jeu4PKePUsCRLHXE3cTAG+H4k+LAlcRIVkEAqueF8TY+0zQFwjRamSBBdUNG/qmC
8Finr37x1RJI2aCXLsWt9ZG7kr+6sBfNQttVl5ErslAJvqmgCGIiQuzFCLhFhBD9
kDaIZv9ADFVCaIevrA/PGLjXstm5Srq+40/zmG+1YQoqd849DE7dbw9dw2DGN71A
bIxkoxk4V1D7K9oIjoEJcvDz1o1bjy8+zaRrGLMWu8qzi/MCwlAVBhDTlUWqJXQ1
3sWb6reUwUKox4e1RrhIBFAXgLcrjvIbmWrKhLNVSTVo3zpaVcLq9wh8GJQN9FLU
FMNa7SbQpd3Xfw+3KxHbyvxNJ8mmMPhmTTmNFQVK8UCTmUwBIw70rb2KcXW1wPal
pX44piUyMgC3aXpHwRMDLp2g/SCHp8cPWG20/P/GmYfA3fUIcTv6qhFEj213q+Ef
6BkcnC7fpkpLNCrQqURLqo14BCvuFSG9+hxk2A1r2NLBk9m1cZQfCJwvvkPMXtxB
8sKtv0dFqY55A0JWVpufd8YKmMoi9gLeaRIVQHSRX8gf4asbB4+08llBCl5I38m8
iRBtNl54Rj5O1wr6Ck4L+qNZ+1rmo2GYY5yTy/9wOaayIJjTkh5EuWNK7fIk5a/J
9c+MbImDkihViXZT7aC11j6ObPvYNuOb/ZRM7+pMC8NvuDyHB4vn1XaFuq8tItKu
RDQrEQdDpwFtDA44/NDyLN2yOpfSqqvbh8tzazBU9O8IIG0ocP8XRJuk/08iCe0R
1M4omyfA5cyllR5lKZPsRMs0JGMu3A3UdRoYH1VKTSRmkEz7evg9HG6UmPKRBmG9
aOOXFJtOJRjxnTKIfH3bfI758fOUB6644dNM8F99i31czlryYE4U+Gl3ybTF8BW6
ACHLMqyQ6WMZzIUp98G+D2sKhn9R7z1OiN73oaOxfQTqW6fsrRKwe/E1mslx2c0A
wrnrA/Zx+MPMGABBrBjrOHsRbMKlHqXxym0MKpvgnSMZAba8qTJVwzWAPaK5LhON
w49BuimfKuUq3Wd4gVF69zMCflmx9GwgiHDvar6lSxRZo8b+vV+zDhf8EP+uu8dM
TWKG7UeEnCzWCsKk6l1A0vtpfnLNR4PRFXn4P5bsHnurenuwGlI4sZ2wE/rHWLBE
VxxZle5cM4EfwbfZEztnrreKQKTQM8Wo8fFWBwcQifnooKvDYqalLF4fvmsaLvLR
bdZ/DTvwhyzA4jBxZeb0+xivlEMAGl/jUk3gp/IniJ78DN4MNu51vH+LzXShBGWh
quf5dad7B3F2edRiRMzfnBKlwFewr81+UTLHcDNPaIibGu2eflO5BIzaiwjytc6u
IN/Uym6A1PtbnAE+SyRFINMVReagsK+th/Uzjpo9UpPrs4Nrohh7KvkX7aCzV3Rb
xXkOuQys4p/ZgKoLcY2eE9E8mDIdxFJo2dxwqOZsqVNVRIHw9X9z2vyh7iajXWkh
4bhlwHQZNhYsTe2YbWsc1EgExHDbD0HzuNmr3xxwJpt/VyjKOgKKzIYBB+bqg9gM
wg403agiPxFmG1IJblcmw1l9CRk86KHDFZ/iknJ8ZOrQLBrhy/vTBC384b3mAVc7
t73sRKEghPofCtiSRwSfM8L6kRskkYpiODc687SW507nwgt+Vy7TLUBs/vslauC5
mPVylVIQv8COEvCqF1CIFurcDJA1Apjg6o7VVh8rZj0pnQCea7NfKLgWHaY6N69v
3FE/6gcVABsibl7veH4S++V7EcJ5CdPcGInXNjQ1HGNaLC03DdHUAI7f0fB2KhYf
9EdaiSZnNCzCEOIgmwli9R6bbICWSwQmD9d8xmxeQCD6RLypt18yTdF72Rc5YCgX
uB7hYMvlar+G+06zxqvnm9cYnsZw6lo/13mD+pcN6/lLF9LZQTPXez6pZNJuqD3y
TJsADnZ7ezXj2yoL29eUsi6lL/7hwHQdXBg2HGWjXAXs/srT/Yy5akUu186mlvvW
WVSuATBlM4dvi7wSTQtlFTdty9OXe/R35sjVhxvful5hVnZrZ3Q9zOhhFqyu3Ltv
6Tzt5SmVib/GirQnDz3Z8kib0odlknlUUNyVggpfVB6sWFBwT8NM6yibd7V5iWdY
YhqjDrTZyfqaZboOo5qlsJMIYKGPm4fi4XhK3LTdWHY2ePIYC4r9Ati2a8GZTyoo
zVSKpZX2R9mjf1hLkmzDEjjqWXL9PrlKYswxb1SRAEQNWjyawFUHXrACyb0+40vZ
SqV0ZuxcBzDcWwjcV70Ye6qRzd5Bstf9aHWu12IqKutQ2Ld3Fu+YPRC8UZC+7ypU
3ogNEYDH5ncAO+TA3iJls7T1JB5S0LilSnJ6WZCu0POIYHFOKYiAm48He0e47nBu
Ok/jmVv6UskfhHZmKBCnKD7+DPqxeOsHZX7CW5bAdh4/XfKSG4lEG40l7ugcgHi6
zZvzqTtlFkJqLZOktSzyJCG1ypkVDQLMhmb4iwxQWYxU4AqOliTtkp1EY2jKWBW1
IaUVa5AEaXi9/SHQcHgF+A7ZIMJ0GJ3ugud/kmBgwiTm1jXPPohXog32URIyttHl
pDm2hbOznE+FiYGg5JYtdgPcdJikhBmx72Qwy0j5ahfM+YIWp1T6chEV+3qhwyrj
Adj6zZ1+s+mGXBQwm25b76VIG3+aoyS/iOzbUs2+XryxNP6DYVmEGcoRcwkWhrnd
KazGrhy5ChR+tGb0qHB28h2cLoJJhZIPPE7XhrvU9bDT/y+zahj8Pkq9u9JmiJbb
M+zRUV2roUZa8d43RAD+wVauuImBdSZg5DDEdNYA3Tg10H9VDKchpXNNJuxQM7gv
5BBGMqb6At6G5cd91xW+ukhxUHH9oxCnr+GTm9p8duOKY1HnlWrtwdIPQllQsEhx
deW3rueJW2918BuZh6Z6QGOUIPAB911jtJeHhSB1OifoxHAI7ovNucjqGwW0KDCt
NN+5MDqxk8m3GDINeSTbwLQssvPRr1rf0eEeQtEH8Pxhrq5+RMf/XmYcBdAN4AtU
a8Ecj3Lb0Ohc1nXgvmhymYezJUWO/w0TTbFFHFnPbgijNTvldWLYTJBNpAb/ZYu7
KcMyTvXVgKAxVShVp1wCPlPrPRyU+69PWZXyu0O757LvfYUVCXDRgyRLjqoqGCUM
ZDzuFHjrLSooYLHIjzZvUc5/OOFI4nRsTEnCjn+qafwy4BSVbOYikkyIU0+WFWfV
/coFjyBgMh/gfcyY8HjtMN2c3N9hUspOLRPv37YNfSryn0fJa8IVbq/sInUaMZq6
1A0RqBcGBqj7ahPh7U3YycPTUV6Mx4aPjbxiUBiWds8vOVKTtO8gCFZ1phwXSkv9
CDosCWhlV32bvUZLxY+AkvbTvZ6pTkfy+TPOft2TTNTjxR6QQ+/F6zhfRThB03MQ
JV9pz7Bu5YU5gb68r63PYbFEwpLS9/whRDrYwn69BOsztM3G2aQkb9IzsHJD8I6G
VH3a7OyxyHd/dlotCDVDNDe/6p4oDuPnk6KOpaIOJou6opGsrwvcrHF6hAPPQcbU
0sNiegL7snZ2l0kxwqe/QskSCupkkQ9OC5sIh4mBrhozYYDM0FsoE+lGsA9/NPf4
Aqe6SYIk4fhhYIL9zaAuyUBURggSohZWZOi75Q+rSt34PTEoEenkCGkNE+vPUGG5
udWMzgYBL3hghOoVyvPfCwV9hrOmA9r++IaUhtBHhaCW6WDBN+2Hn1bjgv/nBPr1
wKuPqUm5Ddt1QzceDcuZ+OCwZsCaQsjW3eeWObMLDo5zdg250BPitI5wpMxaXHZ4
4nzgXNuCuUBU0ptkxcnOt7KSCYx8gYlW2sgNwva3bwXK5XFXXaOCJOeaMDTaeOlm
j/1nHr5PgEhIN4lSZfJJKUDM8UipEu+06xSxmMA6NxRdPAQT0Kn57e3i3Dtw7WYZ
CG9eI8sYTxM7xsjHbdgOa2xNkh/WnMv2/6QGrBDE8ABmYl/o1qBED/e2lb3FYmEV
up5jps97WkLH0bFq4PVKJJretUAUSahIAV1rikrWcHvpDWGr8zPEMEZ09OhLgl/6
Db5u9vQ3fkaX2sCMakVmEWPbSPP01rFCAt990fR6kC6bpFv7saKzhv3WTl3+AkNL
izDUxCSjPlDo7jdxGRNDy7BcpnGYZ/Uq7IhXvcuURbn/LzwZIXi7UOj5BHNy1qZX
XaUy7Pryb+Z+KSCHbXeg7AHr91O+ONDS3SA1cOxxj8G2fQu29nG7ELlYGKf79f/m
kHcsFA7UGCIN3UyNBh/RCnfbVrCeMTtrhfRBZaqGrv0PZqoibCXwWQ9sANrSieC4
BRfAUV0308an2zhV9zNnTPAij5tSxAHNRw1N5XyK5vByrYGoJQuthmNewNDYXHMl
T2r/1E5i26eGxO9i5CoAG+2GIKdJj+jbnDlshzfLZlX6gg2ioKD5OV3UJwl4VEke
6IaarTIWKvV2ui96rvT2dPBZRfyoGfBajFDOPk1Duu3hWhUXDSkCvB4pgD3/qOp/
hQ4z7nvh16hg+K4wCENumIsbEpgi3Q2tTFd35OqLKglAzwh0CfB3yuA/u2SmqXcD
Nwi62oGOifPZv7BJ7jmmiNEDh16sXcoLW9ZFrj7jHODbRJHS71z2msfvUyw0yz+B
QDETQvOFr+aHmGL8m9apy/SgDitxy1taJKQV07LHImIrplJejYi0umjFRhmYkpK2
yxFJ7uYVxlIBls4Z+mxwYVHfHe03Ta6aA+Kg/KigDADoYgixyCTXXKligyf/fHgW
41Rx5dlnbAdaH2/Y9qzcSNtGvZCxyshxb3XL1+7g+cW7pMwVIkO8CclA5Z95KlnW
1rHvEAkFRSN6GYiwOTHSci2Hmo8K/28GEOjURFzXwKNzQjmLQ9Q56hZFB2mkrd7X
mG9X0jOqjvtEFXSr/KygXo4tV0Q8ZcWZ1BsEjbLEOZpX6knOllJmtGMBPYsoBb3m
cAteuDWdxGkYYYEgyEw4MpkYdhE1otEuoA87vqF7mGU+ozGsbMWcnR7C/P6T6mNQ
Gly7WgNc0ZICHm5J4SiMAjPxuzFkDfK5DhWNqV0WQE2kmJqsu68t47gGQi6XHxEY
0Imqe85dsBNoiBYcQ/GYTCzhzaP+9dxjfnUw/9k4rgr+StS4X9Ezhanm9cW0WoTZ
HDA12yWk0v8sN8vN+4NUdtiqZR+rgo6zy3Vp2TydiktNzRjk4BaEDs2JVVdPXIiF
t9432U4CgD/AatMx+RxN30TVBhPsL83EKQhq+sHuiAr4J5WKgt816+Z4FycRLXx8
Y92mMyE9BCQBTdtaRzs406krhCsOZbfQEbS5D197DXcfUv8EIRkp1mrvkp2ompqU
DkZba911sLNvC1Ol1I8QszCrO3jzKUCPsHVVrKhy1dF1yxfSu5OToe/qV0qzh5oO
GZ3uh9XZqKd5BifUeLOMnabT1anXPQrwqu1FT+se2m++wiQslTqtVyRN3aQkvNpj
WoyroR1dwIUhTnac4ytYc6nlHtO5qFWKeG4hD89T+To2oN6RtZYktqYmOqSRNlmJ
T2sP0aeui873sXaKgdx0d4sEVbU/oyWviI3jfL3zygtV0S57t/qoEpwSYf/wH2R/
Y0NhHigmI5DGXyVmzBiXE/XFxgOQqi4fcjK8MN/7Hj5diAc8+ILqnAYFV6ByQeF6
LaMIxrKB3AbfuJdxImdd//X/yx4wcREHgXnNg9QKVDvR0R6iDlpceNQcrqMVHeu4
TfAQsd6LGYs5ZjfVjSbPPAHEUk1E8RPRDmaRy1rW7HiRl2aO953ecftuFaMVwv6e
7FbMWl7gQEmzo13vnWxmhj2LIF3TzPvMcwjqeuhkCPN1HD6dlRDrlm8qko4Tog5Z
Ia3vYmGmlt+mJqTqcI7a8kx4jee/i4ku8w87BQSWMmOJnnaHi8DRgZgzN2FLBpQi
hAJoD2i9FH1YoPMigrzDihz1E7n54yhBnRjB+5grXR8IJlvgGrXm+SmEw5H91gy5
OXOgUrumucfiBFv+S0m9kXEICXamU/AfrfFYmMgXhs8yd5P0t6EUBkoc91Iun3rF
Y5G/rpoWPU8aK8z2FDM/QG+mQbHk9cHt+b5CepLH3b1iAIIM6GrtFTh3efdmOfU6
mAtMGQDUEtDFyYnJ+C1qy6vjGvk9k7t453Prvj3lOdFndk3uu7KGHtAeX3RfOKtE
WsJLyMI4lxWgmP4eYlRG2MiWtHH/tO2+vn/54lVZa23Jm8m86XswJWy0vFqOR03L
9Hl5OfQIZFABrJTJiN081Php6nZDivHuNGABZieF05lsqbpH5rQHtHTRWs/79CqQ
cz2XFir2A9x12CFbHQ4oLIxcMc0MGCVp0I45BsoDqK6Tzv6WezcXrGDuBIgSKOSB
oqoWf6SUpWd3SwBXj+2swvGiBDj1nbpJwpwolkBKJtaSjhKJHdbv9eEgAbhXlx+3
/nWUMXGCMit5JFfPrNMTi9234tAR3s4XjBJzgj3EstwJXmZlgCdyh2nIl6+/Q8+h
NDPvyoA8tH5UKYx4nFPTCtk5tg7Dvl9dPlJDnpHWtFXk1It4fs9NaaaongLWvfAc
+i4w3/Od7vIQiXDS3+2V0Cu0HuUXYqswukQ6D+vKpF1yo98LRXLmdqvoaZy71A9K
ABbAST6Mg+pWT/xMH4jznwSot3FR2641v2IhQayB4QGM3zMLNAEUJwJ6LT5sfZye
7dbre7UMsWKZ2itcgs4XmP9vExSwgr8Otxmr2NbayjAI3ckkvHW7m47BG2/0Gokk
5uAdUckaknAiLrNJPtA64MsOqRtffwUHoNvg/vvY4gM87dpkEYoUYW7DiGN8X0O+
jEehNt7pe2FBasrVIHY8jtHoZwtAwFU4swUGiRY/vatv7KRaMvFnQg905xn2w3kF
YzVvRJ1lJFkMfknd0SFpn0jPsI34mEpuQzbv9bhrqjy3QU+8nhWdgJouGznUvhKp
wXmS2mWTVKjrDjWZvtwQLOyo33l/pHQM2vtbtezJieaeb+xyMZFWXpgf1UVzBWWA
mMRLhIwGqaVI9WE4DzP5MemG+Dm7dEcXA/vsALaKvOYrGR3S0/XvC+rLwYws6qHN
OLuZJej2rommqOVSG0bAyAW36WOTKQzVQZR9o/Tlsy45jOwhXZy539YStOmFtZKS
0OmP7WBfNxd0YlF61rWzslDLBF9tw+PvNy1AEUZd37H02FfXOMTBo3hqhOPBYL1h
1whKyOe/ZT2tbcftVvCpKfsP9nmpPEx6gxyQT2By+Yl4J72YqPceIAxdOt7HlLuu
hu2CuCOHWeGxnmcFHis28/suGoGmuEnTltxaKWo9hg8V4QFJHAjYHLk1bWfK/T+t
KQdCRz2fv4TCubndr/jS/rrFUfBN2/nlAt29T0aDq6r6IvFnOdf6d/MF3VLFCeJl
mR77Tq3hhoPiOBUvhHKPFI76/AWinoEF7Jc55qbA3gUf0Z596vFFAu3EpPSuAn+T
sE9VlbXJnhGMlwQh3VIvyiHp6lkGNiPbJauDfOY+3+BTJizhRIvYUijJ5lw9e1mm
H/v4ML3oQBXYA6YJAZ90JNJ3mOrCtnmH1lgYu/ylES07IUwxVwIyitNYV2BI0Ylt
kCu7J3vtnEypfMrb+iA4j1qQ1S0yhIna7TObdTSua2o1JXljbNIlzeqNsaB5MHev
U3Zj1O662AzmS8pFAUzW8jwRZEaQp8tRtqyRkYSSG64tD97kLgIQIeo+UrnaO7Xh
+Hxk7vFFc8vCAY0OBXJb6nn56vZ+JwzxtBxOa1hNHbP8oBYyIQ36g5cOrhLLaiCY
bRJ2/eaeYLWLoCI5Y8F1FJQvYG69vV7ruXPEjW1XwoLPX1r5MPD1WR/he7rWbYDP
4Kdqc9MDocjYAVEtPIUbL+rmw8LVA0nMgrPKmhAt1q/5Mc5Qtm0MNbTTXnOlQPRc
NRvKjIiSGlhoJUqf1UON1yQIYuFPt8qoeuhVllRLVW8uXZawWYTBhBF1iUfTwcMW
N0bRbamMjMudLU68ZgSHr6lK0LMidDkzB91eaHZkHJndh0Izj5s33QlZXfq7VMCe
g93o1NQ3B6C/sF0F3wKJAukBeb3VExA89Yh/M8RTkWlEAh8wZ07PZMXQRZphEoSb
9dXGDnwBIzGh4WaHyZEBfCOElnsAPoBDxzQdwVV0fjsoj7RDEoRNtduoq/6a8S97
m1yyuBLhHmbpKTYStKCjyCX5VWYhpBzzELc7u2oSbo2rjqjvnpq4TWL+pEs/iza7
RtW2LOnVZe1tLGFqp/aSViZYrCT8nc8RMUYLqqfr+1jzNC/LBoQz+TrB/TjemLpW
XwVJzjYOMkDO6TTM/VHA3hhq0+roUS6iwilTzRYc/PEHhnJe6oddV6gSZXU+AQ4p
P4JgkWtebhz4zo69nrJCSEo2F41uLpccY1nBvCF+ZwEMfxELRvFnIPyfvzYpiy94
2HA/sjts1WKT1tdXOdMkpKzfBUK/EvGSCBtoz1QiAAQB9ctbJNsOTEBWJS3B9DLl
8oS3UyeIzZjffnAQhC5zpRVak44+Ehl1ZHUQqxyYroCJNIzafrYCm7RJnI84rMMO
NK+nJDsLbxs9kIK6mYloZQCUIUOEdF1mBmke6p/rNjuUOj04OVCJPw6XtRblIScQ
Sj+foBAOzEoPYchLB9bnTS7wRKZ1OrLNbMV9r1Jm8rJelovbAqWdqPZB+eufBB5y
a8RvWk2SlQB2W3xa/yTXWGM58G6cDoIpij4w7WFPkdlu7MqN/2f113v+vk4ffHXI
WTFfqvrAHlS9Ph3aLjvw/dxFcDaqf3c6Lf3i8KPJV1deCPAYpT8skBd+GXnEhUEl
UwK1CFVWgCF4BIl2MQ1WsYhSAaSQ14G7gW+NvwPf4luAmKRzF+eyqkcr1BKXOdKJ
es/+BfQ82041AyfHx+Ln0l2NDs4plHBCSpR+HQRRT8BUOng072W7OSQ+83OweapI
5+Kuweq7u6kqo+QJAVxb8GN7hI2YWC4m6Z2V4sC8z7QGH/S3dl+kIKe9aOB9vxPe
OUfAas5fLtDFKen+ueHLd3JL5ACcQh1wmh5/gsFP7QmZkEi9kN5x+x5D3NJAuwc9
gLjtPqP82UrBaHpXVMwVLN8KghOuV6uj0acVYURiSdtHIhl5fN8qCligmK2Ti9rj
dyF8CSTXGFPMDwE15l3UJONPhB9KP/YgHF4Qf1qvRbx81YFJk+2/z1BP8aidM6Bt
ChfZ3PsPaIDEzkWWqgZqxhk55dkVrQlvL0LetcupxX70cT1n8FbWgecxm5sllyR1
B/tGUiFMmDIGsHr8Yn79Nysd4cDZ8kuG3YeTkiXpl5/PuHfku/OWeqlVG1zVBZy7
tAPosxhMCfkItGF4lI+0XzR0+IfmnH50ygWm0m2oenFcRQZYrPlIHqXwQcoYib3h
cByZ+4hiYfZa2u4ezVvkkI/1ov0R0hi3Tq1G6o1+H/d8T/ijyB1/BJiMEYfavDpJ
3Enuah11+1r7rdc8frkFZ8BFHmpJg7smxw9l2Q1PLZR89FYt1wUS3tDH8pvrW1WM
j/+LcfZSxKARnLW8piHQBmAc4kMO4JWpI+AxXrSDSimIS3d6zPVhlkAcqNfagsQq
fSx52a21OKejhe8tLs5uB6nldbp+5YXXIJKIh1MNuEOmSAWaZvRBB+E9F1+PiTfn
Nd0yoIuRPdpdVtUzR4TwHAsiumxeyhmUrxCinWj64aaZpoQs5q8WAiZRsdRhNz4n
zsU30daxY3jROo9X6C5NcVywmggaqoLsq+VmvrL9XUu/WmlyYCrEvFUVnsRJz25E
VLyauxJxrt+NfGLI/ogPMIa0RvCOTnHLN1eRFVrtbazN7Xe16OappeOEVUGjPeHS
fBz7vXqTKotQE5NWS3vtG87zMozerclvue2N8ouithildViB/45qXc12eaKMS91H
+c9LNY9x14gIsKFhcjIx3Tc+KCGDGv/K4ZFqXlRQT6NQA17rUtzTn/F7uV5U8FS5
C8R1G+FFidZREANstTpsbO4cOrBo2QEgfH04DvnwstORWkYIWXB+cTlD+uNyvPIP
eHzDQPruNG1BOBjzyQqwqL1jcPzxWB6NPuzoM+NBDfkagsSayh/wGISYPsUl21qa
Ag6bqN4nPk2ivwnYKZWGJX5DQcBbvLrimyJLsQy2lMQWtEPnSbY3x3Fr0NgsPN2s
c7CfDw9DH9T2zXpPFO+MVcPZYwXbq2h2gpm0FtmopZIMONE/Xkq7ZVYROsRZD6G6
cZsD/3zlMsqp4a0WBeYWIXDY4LWXu1yYXOQXrWtJBOlbhMJjnqRKa0EfqVn0u+eH
AD6NP7PJOT85+jaoGf0OJLwQWfDqm/jilvLgq7eINqlWBMsnlbTXrYDFuhN8Nazt
8FpRqeMAgzjJnQjQysJPZ+npxZRodwOUkM5DXo5Zjt60pCJQ8c3y7nF3CN68RoSA
xG7lJ00jwHKl0UQy1uwGGz/prWeTAE/ODEyC1FoFJY//AHjdEc8+eJrT+JVnSboP
FzFfjuZTMcRjyBLf/5HvSwly9jSPjaP1Rpk4CFRjTxgutP71FkZt9W5FOhHlV7U4
4XKFQ+2ZYV3E/faFUd6QnBN0l2iAuUWRxS+NQ346m7Z7EZtdgx2K6GWd2imBz5w1
HmuDqyH3gucOq01dJb80e86doYBN9SpxMKpzqJOt5OjJTlcKJJ6dWlDm5CYJRpIr
iGyZPqTBiziDt8YKDkNNaSRkfNmJ6rW8lFNHaZs4sVTim/t4+An83cBsJw5ouWS+
SERoD2E5rXUFFmVGjGmgp99MCmktt6d5T/3TZnWsAuNU9hynyJPe5bJ8bfB+KTOi
qN++gNE3UwZq7KeI3nBIe4QG03OhK8vV5rrHzJ9YajfFtFzuNaONhIPKloUIyY2/
KJzr1fXohRGYkxq2iDNq8RCBtKHt/l//yWGsaYblZc2WpqSPMDFGOn62QHmmh8PR
D2fSz1rloqlByq2Wsh9dQXvm4opHRD0wvz8RqcHDTtWzWZk5hzNMFlqMQZuwahOd
XGflBpp0g0pFN0tOLuEycbOYVmRgnBBftdxIqqlRL0ba/XRg43ajZtxsiUo4olb7
iF9nn9Izw6qlnB4zeWmZupXAJcF8M/w24yc5h0g94LM5KhCcbgmkImkqAyAbC3EQ
US2qy8Lo76tEabz0fol6yhbHAysTHjEdUfd9NCNAB9o87LW444Rrp5EQBBM91YGP
uugen1fFOAwFfIJtTMP+rRDxd+Jcu8c4khi1UjghZsr7oHtkZ81cCLyyeP+cAfAa
SdOMOdxO1H0gBNC+71eLjn2Yy/2x25KZyyO8wF6Jum0CYe3fShMW3RfnT3k/tuJm
fYVJB4X+UudQP3bNiVF8AIa0x7435BTWrIrpEZ+llHA0eQt7xKrlaEBlALBLUr22
EDiU404mN5tMzix8GwhyXs5UsGkvboyTMPXHhOzOUWdLKgn2JYy2vthpjNm4+2up
DY/VLKwlBFJxGrFbj+yEAIgZ7yU6+E/higsY/asKQoZfC4/Kgf7hvriUWnbdl+T8
gxFBzYu9cnujJ4k94VpwA8Rwni6/wj8jd6FqlBuPXg0oHGCNew/Y7rWx3sJ9KWIh
UTTm1ZbArLxpehEIPEiCYXWN4rZr+1s/AzmTqR4hD7nr3hD2Uu2FUvIEysXSiJ58
k7D/n1s/9LFimv7BUip59AVQ6gmdV4q5iaOcOYSUnxmfNw1tXws5bae2qHQk+fSu
ICQj1LmIdIUT2R8oUtn6Tl2Iqg7/dg3DNqcz3b7OwnngVkE0m1+DMeDttWgksOku
2pwZwEx/2HzYLKrfYRkSJA01KESZ/QnIW6mKTgwhHrxarNA/vryU92uECmoKiTh0
61eVzQw8P+EkjFUXEOCPqQI2B3CFp1khVhqxE3HDisCPTMidQYNLI2WBO1oWU/6G
B+OAbdz2k8Jflf0chja26KlSud9FevVGid3mQVtLOaRL4D/jhUziUPJCcOuva8F4
ORyoywdD4oXQBe2oyGR6bjXeVseTp1kwErafM8uIGclpKAwIXbCkXycmt6vXBnxe
18YkEpFfV7pXAtbovnKeEy6PSL+R2RMBGUGLn/bdyc7DBftpVsW8eswn+1Q4RY1R
G+nz78fNCL1lXsdeiQi6f8+nhsZYZ51kpjf2aX0gHtygJ3oI7m68n0mnvKQGsc45
P4hpiWzIGH8Rv1CK8wP6AJ0WgXwyFRo2VNwpOKG8TDK+4ZPgWLil/8HzuLcH9uxB
6BOCIQCfxbyV5gj/4JVb8V3xjn8KQtiOOFxWQnKspjDXxE/dS4SLn6ZHUpx0s+ZD
igM8FinJXluUhe3X5nVfu1eznz9E2vl3EFP9/d3rQJjiyxITOirO/WiNmNd8Ekbn
2KcdTmAVcMdwvcu57ySDA11oYhwfp4KTpdgCLcy2Xaeeu0Ci7SmnGNwCA1x2/vml
UvVviebnUpXXLTyON0kB1G+YSCn4qQx3rvCCZjfMeXB2n8wGAfvZdNch9Zw934QS
MUsq39iHsiMuGQBUwhex/st6Q/0tw+PPw5ZYdE9cDcdImF5lO4e3BN47qKAjthHn
zC/hb+ijwld5uW3qq/MmU8AgCN826qyeRfw9xCpwnwFcJ1vOf1VFFMpzqZP6t1xt
RsurQ8n3CZezjQ5Z/jE5W51xp3CJjDbvBWQ+guJbee0E+dWTwlNjEj4pfZgWueK5
+FC41f/m3P8mgv2/OPFslzEOPWC8Hl3LYcE9nYurqNCBtl6LRbMd20XDCK0YFasW
/xoagtDPo4iNghRU47ARPzEOmtDueuXJi2RE6egzoixTBK1EzYf8IC58QUDJzGrc
6NpiSaLM9uh+6qVTmlJaK3y28HZZkR6XNWGwh6DwMqNe3C+TjTBomDHcHsgZCCrr
fB2QamdieFeE5i06M81fVrC2Eg6utK+xwoi8GsYGp33myCeB+4Do0ISbBkwZ9Uf6
YMP3Is5Pbkss5e5BQ8RxpRz3JzwrclMjEQyuYEVJU8kbRlAOrix3zyRXkAssFfjt
SwYeilFOekXi7TasoqGE0q09g5AVcgtk2RBb0oQgso0AFLtJFv79p915eIEjPUTW
9VOXjKZfvPUFF7BzTbfMhpyTZz0reZYKOgvxQ0ms4e+k3XO+13FJv3qJFx0nwEqV
JhbiYvlVdlx7ibi6nMHyCwMY0DvEGWx/o9lQZAKiN2qFa645Q6VUCHW/L/+gF2nH
hFlapNOH5fwHogzc5qRv4wNJYt2oT1ai0xNM79zsIvNs5fT02Kb5hauQ8aXn087k
aCNHtWbZECWUdYmfudaVe7McaOrRDgZgLsNGO7DxUf2IwJPyR9UY4GUQjhEzvQvu
qcC67X+bY7XlF4w1SA+VX1cZ7iwqYCR4IgyM8e8cmR+SAapxbZL7Exc5E/4QuhYS
eGB8cuINX/URDMaOPatpT/baDM2RoCIzFde85uHuPB0ADRir2mk6MwcQBTjOrA/b
sgB59yrb7H8ERh20yKfHMILPm5kEe7X2ZnpD4sFjxaHuKDdlwJ0FQ1iXhYNx3hqU
JPXyOdWKPS2CXUtIWyQ14KqC5L0VwzeyIudeVj87MJ1OlI/6bxTDHnp07qhNPsNB
lP93rW1GLizwMoBgvVBcj0G+Uu/Hl0/XZkirrJQKYXsmiqbGZ7H+dwl51J9eYuMB
aJNllkKrX8n/K7W/bo9SFwrjQemlg6R+C48T1xpZqzz0+KvlptYvAYLvM8Rbx44r
fr4uhTgJlBnWxFDM1v6al9BUm93yE0mxGNWsVyFkTEZr8D6NeyJPvxd1J8VlAqjj
xR6hCUzq77RrVNJ+UL+bVMvx9V4e1Dq4SSbYO66TfsQ7DbBsIJiY8nR+sMXZqO6U
EwRXAdmsNr98Qazf9yaiICe/fM/+btL2xy8NBbHXMeF8oVsK1eQ273clBtHGlEgl
rYACRkA35JOVCOlJawmtNBPQVuMFyCDh2mV2lq6HjrLxxqTSGwbB4AIIQ77dflbk
yr2y4mWXt6qFuEssKTlOBqWt93dmQmUrQptOJ7rEAmnXjEPnJGWVlrrYtcRt4N9c
h0NCPaaZAjMBnjbPcnJAW3+IdhGiyecxN1e8xYpqdY2pXjkpfYw4o5/WKxXb+2sC
EkFfU64qZn/8TWTXCSahscDfyr6EbksqymTCBWLbO4tiI4Cwh8EZ7uq4gEekPI8Z
lSAwTlukeAkbWiIg+yYt4nt6QWE/tnSRQQNVNL4nJPZBrsQNqsBff1cSGBkhR/iq
8x4EpwKgZnnCNUd3q6YglnnIwThJDHRAMg5QTJsX8tyaO38IexOU6yHVw4Vfnn9n
UkwCGYeViqrAAXVGQM3XizQJsHxYh0/n2d3dTdhovL46OBsHwh4yRYIGtJtL3iGP
wX6Smorop1L+lCk07Zbn9N6VAvzAYi+9oBMqbdgp3l2g+X2ZgceKJC2rkL1zSqR8
H5ErEWwTCccv7E1tMSbyKr4VgrfkoG4n5xJ3Q0RQ1tTkgNcMFMHCfy1p39h9fPlX
zmLqFUgw7ryaFXnTd0U3CNPmnANreeGAwqY3+7KR2PygHBEyN7AID1/6ejUDh6Oe
uP7fjCOvoSCvi0JEfjAzW8g9WwJ3TM5HO3favVDnIFbj5YbQDs4MVH/oqIEVl8N7
NpC1TUtXXT7AdHueS1P6LsuF9RZi+7lqlndOVcg5JfKu/KXLbIvK4fqUHakFyitf
3rbf/SutOC8LaXUTyoY3TAfw+Vd4Ao2mi0Jv7MZLx4ne9C25RiFr3YehV95kua0H
H50B5VcKemUd8suQ7bAWXjRcfzsDgeMQf/sJWG8hM9++pBQvRpEgR8m4yK+sfIWY
/zQ2iyZ/mrZRaMOM57QWuKFF6KGNHEg7DntvIP33Y1TUKe1QJzSXS1e+lx/eczss
Z6VhkdI0Zz0Cqkp5t9/liBFPc48QVFcMnMcjhHFtQyQ3QhlvKs2+i26Rs1exLIMm
fAFjMneQoXVUF/XMr8ZkBzQBZW+j9a7EOn4VQqrVIS9hCQxXPZVpdNR6yihKoCGp
axXBSHXUnu9J0Ik5Gioa/9is7YKE/vG439NF/nULatIdMFzJNnVceLak+439P7eM
HAE1BzFtv4v8fyLKrN2Qk3gT1E0vyEyDe2CZDggIMPSkA7BgZ+/DsqniTEak6ZF9
UggP/nQMx6vhqOK98mftFlXnAv9iaKXqCu7mMbSdp3u+5E5P+vv7ZzYtNw63iHMG
1KsnNYzcxb4Gp4xZKs5oEJdJfL6Y+XuuN7LGqFmDorkbJT0ztv1Z9R+azXu4yoqA
Mn1s+H6irddLCJfTIetHC1jtLRctUWX5y3FHvYaAufFRhmBCevTWzQT8+YDTicoH
n3UhP9on4F2pUq/hV2a3kL29j+F/QIqavXeoNhExvVRL2loA03P0l2eCxOFuqSHu
MuvUJ5ac9rIozlhNwlh0i4ZxGxpFXizYjOEqSHiWsqnDvSXsSnyhHb4yVIq1GliD
GifoScciHwamF1j+xqw+7B6A8jhZ8DcfLVjE3VlJ2RFxN9bZ4p+CE37okxbLn1yG
P5KtuTJu0eZ2JtXT7RyB53GUJ0NLYLt1PIbg7w3UZbndBkXqAAAwql5jDS5bAzWd
W8RWLCRpMClmH1qzKayYE+4aryCpYu+qDzACDDOj7J0Cs5e8Olwo1PaCq+KH1eGd
35fanJud7681nTf9jHYxBscdhFKVEfS/Lw4tmQxnXKaUDrCc1G9cx6v1lO6gW7FH
Ie3ZsxLz/RVzo5OmmPt3gSzVFqeS0DODGOvrijdBYFcsM3pu+2/a+Qc/eD+rwE24
EBG6+2DgMAPK4gulYVqH/5MVR9fFeyC5RyPnDxopYYdfRUj+aOhEyEDfcQJVVCJR
CWB34P1zxiy8Pk58M0IOOYay9VK0Msy+HqoDY9XggwNKbn6JQ3KOiKnEUCUzLjbq
KlVszHhXd2bgOvjPqsLum2KdbQ9wgke+dcVHfHdGaackDXNjoGzGV3Y9uKjSL3J2
vOjIBGkp0YPtsn0Oh8TTwpMaNDXevLczcHXOn98uWr8Vokebbh6OU7ZhbQpAAOv1
wclHHegjr41Ogq2MledAnhoLJd2VJIcZHPjesWkyVJybtIrJJiipk/ZDdwt/83re
Vjd6zyjYUIYwqhOHXq8+5wBXDORi5caBBCdXNCfelxdDHzXtMb/mbG9XT/4Lswyx
m/fWy99wIjBmcz+nd2HORSdrmQYdnAEM/HN2ZETRkJI1snPsV1bF8f6groljOlnC
1C0zfsYyQVPiUMR4REWYUcXJSEmbeIKT43UJcHBX6PQPA8wcnjPMkabAWM4rugQK
1jHD3j3rhRNGOPRpMD1ho+D/zOBL/+NF6NPI8giy6qlmfddf0OPVNiRMhLc+s6o2
+Utd+GPfgjyDqI/dXrpcIAZAA/WbN68VfHvaxdLxmJhAKebBrIVm+bk8N592/OLe
9l1uqp78FXZo+aCzu3BSMRm/xcNOuUYhvtPxOOSkw8Yil2PBLG9/Z0GmZNekOMkh
ONGGQ9wwwGGbw+XjmWYLPgQ90gg1ZwYKuUehcIdHEp2EFbs7TpIss5u2+Rt3fZMQ
02/Ydi1dQJMtEG/KdRb9GxeYZRqPxmsAbnk9rsbrzCdBmHTyFOkEbILNPV15o4yh
Kl6sjopIC5WHSeXzJjmS8zWoXNJS+u8anmvKbUmxFWN3+wlf4c/mKO3lA5wDS9eb
/abcEbjDoBFrTnfl87JZrOSaxQ++XcGwvY+K6S9S41mS8zGK/qC9nuJVLItICMcu
EQTyu9YSMBxz3Sg6iq7m0tCGzU3P6BWnI/XT5rOM1wGR0pyVSz6DhnDFHlDwDeWk
9N5Rly++S2wLFxC83RaVbGqDWR1u+82PmvNYS7tBzZdBGjVUqiyINpVXo5IDeP3z
LAKmDcd6sRONzol3YXYnuXyt5uE2l7POGjmNBVhnk5ZLw1qx7N0lsRbx1yWzN09F
2t4Xl9aY+M29CS56ExaYENCI7sefCydk0SPY85Q54mPfzMbzYT5xFa6Ho+2YTTLq
OzYYBYZeWdJPimL9ugC5SVUbKgtB5F0eQfD3wnwshySpAmjvAANoRxtFIIRcP84K
ZZACsAeA+DNnlTefm4KrPxj7imeZUkVW39mqbm4kYSqdQyIZ6jR5p4dvi2oel8A3
TD1fKNUOyjka0AzCakvtIz4bMprlvuLoEGiS+HL8OuqMR6iiHDONu4ame+aqKxLU
YJJ8+i45yFYCSSXo61a1TxlZoXMbYcQHpf9JN+yzwlui0x+2jriUM/DYr9iE5owQ
i6826h0FuFA19pZE1ddgyatOFqmg9p9MA7Baxbqx1+t3df8ZCJR4eXGoTBELubWR
xP06Aqry0SV4ZSTMEMc/QvyWwZI5n4mlsgcOm1oLK1eEOOj2Htjs81NiodZEBEfl
0rq/gyW+i86yNW2ecWrOMwvy3UUN4iJSVGtATXgJMGKQXJMkbfxJ9U1K8Ic9OGft
9PERPrfOlzB4drAsV568xvJK/yJd3DE6vuujnutiP6D6T7NZCUWZGM44Bo1ISnW4
EAlC35HMV6VX9fdXgxqWQuo3Z5y+Uab236q2LA3BdLFC2h+V7RZVvfp0r9rD7tQH
0l283U/E5fHcBKjtXip3jN613OPLPhTo8YcclG9t5cO0kuB9uRswOAxnJu9Hk6ZZ
EIS2ALfzcPPmZEOxjC32/Igd/YqW/PLmxOt4PP3tJR6Y2AmJ3vhxHPBAOXGavUob
yBnfxzqMTVpNYnuIQcMA8sFPy03cSfkj/2BhicJnne2BJJTh2zloUOJTk95wyJzm
EDOySpKySEnsEr0q61h+Q2RUTB/SWXI/UUeWIhZUfNUFNcu9nwetepIrr8HDO3tR
hHaqDeg+IySiseKViaUcWBrABnux6kU7/irQMCXeTzFik5vV8QB58HvCUkX6y4G9
20AtXjf0HkNCv3XWU8n114PsO7KavumFlxpuRJQnqnfYxG8RL1PeLs4isWfTURnz
beetMhJDK6mF7tqMINCICfKVWqzWvw2ndIy/fNUhb28AcRL69jCZazZhbsuImkgE
H5ZgFzHr4KazU+GGpwqq63y0uOZd1WSK2fyXu2rnAfyHDso5V7xFgtRtwiMiGLIl
Bn49S65QLz3/9jmahm18D3/4600+QjAosdm04nUJd1Tdcq+97v/+CVb3RbEGbnTk
dbP5auuSiFSH4uEWnddw9THu2lWqkxyg8S2MragqZwN7e5FadeZ5eFQEmshJssEA
SrsOQ8AVmL1mWNSYYwwCunRvfRFrjIk/qi+mvQcimOPcmB5226Y0oZdsX0Yuyq7a
Yc6KvQC0X9c8inH0GiyjccgyN27C8bJyaIepugNMYAHqlB3ntw66kLACg+dZCiGP
c3IY5cIihiQ+3hWjEfp7hwZwFXIQqNYSITyDCwmUApargs9AcAvLyCMfvq+4//LY
vuSO2o5EVLYyyc8lkqTKMw3/KdTGhOgQzgsM3lBLv7HDlDHqbGSlJxXEgMN7+CME
qyW0yiFnUGsdR6yt6dhzrtXx9xJxmcWCKn7qqefYnYSyyzhRzKUotyxkZI9rnGIk
tN5dQUKFi3Y/jhxIQnTa2xijAXirjehiST2aN8OSWPp1agWvhKJbuuelCYoZtWYp
1O7Dy8Ob2G4966qa1AgcVLBjxxyLzRTbuljHUV78w63cM5ZHnnMbTwGl0UkviChk
d5kKB7AkBoBjAKbXhJ6HEeMG3faSskE8erk6+vuwriTUAPbACue3IHdeSeXUJttK
fkNbn6X6q1RlSZ8m7ZWU6kfXTw5vGSX5VWWVy9ciAE9pf4ovvLhq39DOCX3zIEUt
0H0Wz+P1XUCjn1eJjMrobsbAQE4ahR8/5KIqKtoqBBIqXXGL5xRwqhVEItanyvEk
0fbf+Mtm+M93GOSaGyQReNOVIpSIvEJa08eHiT4BNRXi2dBRdLJUdL0BEdYQRBJ7
CK+GgR8CIS9Ed7QW95UzbEQAy3x6cbVp9UAJ4Grhr7xoCOC8yQ0tZPcSwauvTR9c
TMt/WRxTzOkkgaeh/ielnuSJ31rx++17dBn38JrkiRSo6hs6BvVOq/wBE2JoMDZ+
+1BlqiPZLLpyOg/sPm0OnUPow3RBFTk6RHZP5wC7NYf08t0BPTXEa1N173Xv5RH+
QEBheC+8EvSVHxZQmB1X1Fw+61danR9W3bFDAAP1sTCsybDs2nvZG/bEhyo7oiJc
GEWK544jzdZxRSDrGtaOaLX/Y9Gk7LPWUCOock71N3skpLvLq3M3109PAyc+03hF
cRahiBeFigI30UAOIn4q6j35FN6sdyldUvz3hFs4jRiiVqOIAkDVcRT1U/3joCBO
0hCqk9u2KgGEVFh6wID7iVBz41mlKDZ0TWlx0tWikczP2GOggclGt5tl0Vl1rqju
0ONVJ3vyjCBCV6qBUoePXjXssFYy3S04jKKDkSYOxVSkTZq30xGixWmq7XUj2mpE
adgHsxNAKh2RAi7bPIpfNL7xQzUU6aoBotcVBESkhfuYKKwmaF3X0QLOKZBZVvJ6
XF0l7IMX6YcUqZiRKSxvu5baWu9yMc91VFfwJ/zF9X8ATr9A8sRR2i3e6JMCrpPA
EEHSCdVXEL8vRZghVr3IKTf6dC4I2P++cSIKt5z4fzeSnTpcP6x1vx6thL2hpuhP
GuEl49PjWhkaM6LTaz83hYL+qbS9I9VUaTkcxHG7yG7FSCIaaYLcmyuLsd8dF39c
1kayncSUnS0YAALmSYRwie7/9N7E4DLmu2OYCv6H74z8MGF1nADcC5t1DNqT+PK0
AVXYjl3FROUw2xjPQusmvp5J7qBOFwJh29f0oF/GH3rjUgeeUpCoji+5U0b2ExGL
lT0wqJzxtGljAUbU9FGr38r+5E0ND825ci0vpS7TlE/ra+tGqfhcRKi4haMr7gKW
c+O5pGi2zinHuAHvh0jcoww9PBBJ/MmmXnh9+pvr6y4aNgj5QFZY13MrNS4Xkd16
zEZsJ9W+thubEaH0PFpmjK/lpNrfNcN29KFzFIP6zf2W20TAHfHpLNs5rJJ502MQ
K12aq7pHoIdUkCCA66wrEzPGW4P2boY/fTzbK55kZt3yAdp0RHboaF/e5B4IMSEC
HpfytB10vR8qEBRp08Z/vf/ylcBXVksiRcQQIievLv67qTL1UhfVU/p8WHN6qc+J
zfTuhE5eRTExpg6yEK8xLlcChrEcC1tDT3RYDSS4LgTy0F+49rU72Whl8yyDY5jN
ZU4uY7mKe6rkroVLIAfD4V6TQQri8ULiXtc8x/NUOF3lUJda+i5UMsNvfbfS4blX
KGFed2rD7Ao4YpY+GYLzazGkbZjwOQp6nH0GLxNJ8wAbfLa/t1XPvZv6JXUVu1JR
huetPExpCNldqttbzXIKMFkLJc2JrMpgrVED3OPMpHlKntV/1N0mkjxcDsoTHFfL
5NWdP8VwRuNIL52VOOHOL/IaJMv4ggLbfYZyUjbtBb7KcJuP/Btb4ckyTSOtzWM0
wbBeWxWCSQkaLSK7GGSIkIbuPrdacxn1U7n7bxWJ9+jFaS8DUKL/YZ1twddm9dEj
9K4aBsPrtDojoWQUn3vJ7F6hDGPGaIksUBgx6BU7h51wtru2tvIiqRmxvzZbgJs8
dp+mhaAENlxGf28D7u2Nc9x0K6RaA6jEXqrW3EVA0c1be8e4VzVbqmJ6wGmo+hRo
cmWmbm/tKAe5XK3gv4lQjL6rsnlIko8Iwi2DfupLXAdB3F60MMz9ufCss47eihQn
VZQD1coCyjSb5dkkh+474BLmb/6ejumsL2mnu84MyEn1jaQEllN5Yp2iZNVF0H3x
oZGDTlrSx+Y86INi/A4fLY0ceE9lfL2+dPMgiDXBOiSxiZagP3be4ewPCS/+3lyl
g3iBkLBLWhClumB0M1YUcAYHb5xtvT+cFu+fE3DEYg2KWMfcgJSiEqt4wVO/j/eP
NrtWAzak9v8dAMZusQoJie7NAN5S4B2jucXE1bWH6JyFqg9cHzt+4di0OQpRJWNw
rp5znGjUyVKaaMMwyuqlOb6z2WDgT1tdtoIx8cfGyViEAvdqssEaJYwBvF6mOU8u
wqTx67dUFNf2gWOKeWVawCR0KdbB178JKgTg5OTFItUlbGiCaVdU77oh1n4INxHF
cQEJvgBW/4FSv6vn2OMz2Wmzw1oaD/T4G9YAt7X1Y61tOkhLCGVeNhAwKktLmsZB
foSbLpe8dRdLPNJPY1xAxSBnxRmCq8O94ievGrswmedeTPCJ7QE4DNlwuSFHicbT
cTJlUo6/WJdTfsoULXBiE3Q9UaS389rytePz/sdNj65EgN0EDskSbYY21mKe4Jno
aklqqQEkCuj+igXwSkBCRlxKCmuSJfgctXLVbaDUzv+LQ8jzAWKc62vVaCewBG0p
nS0rf9S8blgVh3LzsOz2nl5EldCGBJ2Ac7Kb+sniTrVbZ3vbAPoCIGVwowmoP8uL
2mmpmvqkTcDY2oXKQ18BNi5gQPA6L6qJ9DCQimNfJV+TCgMkfFMWd2g0qRT4q/UZ
T+O9lRX1xBjqyhiilROevoFcXmZL1DBB86e5RubAzQjdTtKmtluBH6n8UBLf3h0D
X7oCnIDKL9wvd01S8MvpA5L6eVl2trOaSxW2wcMOBynEt6hwzR5T89kODhX057SM
lO6WXaNRPS5U5USkyIh9zBNdgnVcEOFCjRLaLFAUqzZ11to7aYXuRn6fQXdlCCMX
xsLcew5wzczilPxzY/mVOA5e2WYdr8RfAH9swooywEXoOXsm/K6H551XInCpC//4
CHX/LIqU5JlWDnPfuX4T9LtQ92sJ774DpW/3mFRDlHXokrm5GHlmm+t/JMkgfq6P
DVVZiDRBKTHi8Jn7zhb6h5hBJ4XbfcbbD9Hy0sDF5FN86IenIXt3kIdpIk3VbwEv
743VO0N6++RoRH23YdHViT/k2tvzzlKZ/HR56XBZlVX4jMWc53k/SchjYeY389ac
showYb0N00jt1Uob2hOhymd5lmSXkUD7P/hQz/KIDxzQoVpfdEyy71N8cpU5Lv65
dOy/04TysWEGpXhjL3I9JYmbpjjtTJzAJqCG2bdjDjby0l8UdRvGMK08+GYMy5ve
8a0kfvZDliIg/Z9vsZFfHcTZLE0uq0CC43sc/PTiWhwm0iQUw9DZKKSUqTu4Wv1e
qmqgwVpUnAi4//kOh36vvNbtBa9M3Zm4mG3mleAEx219NTvyFuzPe+YqkbcYYBXW
gvkRVT2INhtfXGGZ8fpKi9lELAo2ruAly4xKqqJibaOn+QeAA/4ZfMOOOB6ITdgS
aVWi2xr2oq9MAuFLA/oyQryPXVh0AgiSW1c3tk/Uma22SS2GpTm6r2dOopnyJ7DZ
YtmRCYKXRbCAALZWMftwv4wqZ5/Tl3GCmrJPU++FTQC2G/EiPheWZ+o7uV1sjrER
UVzTp1+mLzyApp9mNJ2XcwBXMZGwU5F7rd+yqXLvV7A/mMsGhsqS+VGuF4dmu8no
cW+hBWGqAG1y3mBVXiHEFjoazwr80GV6HN6ticoY49GupUFxWKGK8i/RTqgG+zJY
ZkDiMqmLuSIvP6WRkuVdvJuX+XGoCLYNpJbxVBU8bgkPQFNxpoXpNC6M0oevyD0R
NdpkhZ85w4zF/0iQ4Ao03Xv3UsmDKE3pWvMt3H6mb8ESehLa5bba/rq6Fay0/ggb
UkouwckUm0pthXEWZKWf/wsNA/ph3XVOD1rTtBHuAs+67yIJo7LMWX/Dqt6P9CtA
KMPxcAfx7ULnFu88qY8ttTA3xEtxWwWe9n/F4Hr6EjMwFC1xobOZiv/r9b7q5KyU
p9G//phXiTzC6YPBxI6sHjMUf5yoy9VpOrcHLL4J7T2NxHhzNztsGyVphVkEWjHp
IBok2ov3IFlCeR4x1Z2+/LJshV+BYTuEBQQ2GFnnh+gsv150HJara4UrGt/ThnqK
2ywy4A/2n4Le2zS/0UvwARgNWG2z1P6IixOHK5nMm1Z6MgD0OnyeV8/uPyWtwCSy
r3etQi6rqNF2dnZTFiWxdETVm7XkYsauhTUC0XOYKa1mMoUrZrS4l6FBJnrT04RR
jEBZON2evYcQDg7V5XQuqxj3pxhTYs/cjXpFdCI8ViwBItPO/sSEc3Yk5LrBZnSs
bZJQ+Lj36GLfAASfou9gxk/TF3zFH34jfJ+j5rCXygJ2Tdo4eV3bsHd3srCQeVwp
NLQLCpBVq1lrt5oX31BZwt/BUR9+XFhduIF8ggq2vO5ZEatQpbcb1hLqqPOv9DYf
K0CTZ6reSNyLBi3Bn2lRq5cTwz1ENlgHKtLaPfn0pqK+oFOQ2UxhurFrcrfZ7XDh
Jhk6A8MP/bh3z93+mKcrw/D0aUrnsNQIc0EKbvvK8IhIpdgnDxzfauQ1HTNo3+H6
OzaQRrmoNwJK+no1iK9wcl9jMSoXEdf2G7aLAdXAKpPd07VlVsLtVkaSwuimzLIw
cKsqe64+vcYppri1nUY+WyORwgymD8Je1rGPPme7qd9Dm43iCWv74HzkL2rlhzbd
1LLtW256jqZsYbRvC8ONDxJB3465uVzLDwnnrU9D+ZJzCasasomh9eYlDeIQitT4
MQW93WeT8VYehKjeZ7zSb1KJJOuy84Q0t0NsZbhFakRkaW2FEhlIatg7SBX41aq3
RAJNc+YIn6j61Y7vFqP/yQyK49qV9ctVYa1fe8GY0U7mdYNi94ysHHGcGYyZxphW
n7bxQx0Nk+wB6QqyAfeCH5tdH0hlcn6XR9K5rRoYcWFuunlsUrKhR+ym0TBVEEbE
0ACzKUpO8l7/i8jQkg6l1tK7GdikTDPetzYpstdJX/jnFOvpskIbUPBpSBdyIcck
hBrj2ClFNem2Vozwbi8XZebzCto6q0kq4trnmueHPPSvoBNLAhxB5fj7LF4dEzXB
9g98C1ja5FwIE+zi0ifA7BIRdJKtCUkHOeulMGwkGoNo7Cl8Xa49Wd/TiiOo8Ccp
SMgoyVzv8JGs3+DZ99tgDcXFWjySqaQJjFm6gvdtbXOsJh9O0OHvRRErlJ4D9IUU
kqFsV7vDpS9NVEcMJHo+VCt/4QVnmJgM3uwaguW9Cyz74bjPk1gRt4BVn4fOR4Rp
WsGxtrg+nFCdzxS9Ovb11O8m55xx6DSI4qtdp/nqueBVuG+/qBLdS50KNjHLDBef
F2P3iPnyjaAqEekdgU5vpAtOKZ3XvWFPWvsprPxUMSnKQcidpCrJ/3Wdi7L4PX/b
Kx8POs9zj4G2+ZpnoEsAWqTRh0FBMTbDrD8Hrz2fHjsyUCZOIAo2OjEgHcqV6uDn
XZbetnDD+aDBzloi6xnCu7gMmJqwWY1NMW9ZLnS4nCFrPlO/O1jESYg5PCTbxhQ3
n6yvlmypdhvMdZS4R8I0/IJtCDDw9ctuiVO6qqNH01HlpsNqGIbkwybzebFUnZCd
nBQ3hCIzwgPisIC8dAr5Lmd4dYAtvaHKod9gpl0kfEA9kcaG9AyA9RPJzpovkXO3
uDwxiOytqjI+bGsPeWH6YSfZ6fPOdG4lq+O+Z/iGvRonG4+0HqftMLTCmMekbEdO
JYVJaS9aCdGfmp9Ix32LKnqwO7LjsgyzC58FOrXZdDz2n6vBEjvRIdyZJo0vo3oq
JshkA2ym6Vs/ya/JYQUoqA2zH7QIGaDgacv9qmaAbQzHgeqLPEUKDWM3Rvx5Xcb9
6VwZocgGqFbWqHzMa+3Kvs6ezwCBX1e3WHvCh2+ZimmZbNpsNarmwFi7TOrz7QYR
RMoeTXr3itA1icSwwRXou/sp8VqvveJOqpGJLKwGJK7ShLB5CQatedXMcKech3WO
j9mko6VvYHr7n/2uGbRG/UTOZoQMZkIfbTAlvXizaP+e8vCQb7Ly/qR/dY0Q2p91
tHlpfhdZus5tQLPpZE65y1ya9nVGW5Lq4xjeXg/4Y7PNyW4qhqLMKR8KyUBYKja9
qtdr6gxC87XoMVE/Y4FpFds6fkcItp0cV5eLYHX7C08VX3kRYGbAZQCadu7lak6d
jGhPsvBxXKxXKwwDxkP89ejUooYMxkmfT1QgMjDkcLmU0cIeL6VxA8g2eC2u66NV
A7SBxHhSNWTIVVG+p1/75WraYuspHR+OlJAWXPVY5a0cnDiMrfXSndkPnRSM+yK+
lSbjyeFs1TnjIBfVFsnuWPp/1WF8vitiqg70ChkuBABgeeXLmETJ+9Ysx+BONqJd
MXKWlgz2nyaJFlspBH7MkwjL6Kzl//13yGwHpn3DFBzvZcZQD6ushmlmzbjbS6Gd
/uAHNaJBJQLnl/g59WS+FGWVGmsLK0r073uNVDgdJeHD1S2vwG/nHevWEwVw6noX
0bK9zu4K3tVt0aUAhK0v23IHl7mCz90CxrEo225hQYq5CF0/QI9LArqASLN+KxKU
uCHekJPGQeDstDWStWaTW8SLNxNLDzyQRN8qNQS8PW3O9nWpXV9m8nsPp8n9soBT
e2887JgpT9oLvanhA14lSjrm+t0+c+XptuTuzSGaY1Y1bDqugEwPVVGq+jzAGHW4
64U3dnyvT02QuJXVzX/zgQVD9FiAp9T87qF/basq6W3d2aHhnIY1/s6YeLmF8bYZ
2bIkzOmgb/qJlQvIk+0XVkZWcl7cVsJ2qU5vn67uCpIYejaw3kuE+H0S6at/uqHY
uQlPyHSUeRBUQjDZwVgAl0hVqdEwBPgTBIL/9jcPB/MDYLN6ARAdot5AwhYXoLXN
PVZRZ+qhXz2fvh1xlMm8cJWn71wIWFYqfzf1SacEFSuPqEks2cfPJpJMVmgxm0kx
fFPQUCtihNo85GASqSTc8h0ruXwZzTcVvVFddm9EoQ7odr3lODn7zjGg1v6Itvu+
p6sq6MDgLqGqPKn55/WGHdpL7GDGMOl1blwBPK1Kv9o/5TFkE2nFUUW6t3H67gCL
mVjE49Cbvygd28JnWCPyFn708ghxiQHpuRpW5bo+8pU03/yMYMCaEPrMnEpZiMi6
5SYZlU+GAwk0EVPbSN4+6i75JHfPfzw0evlzHmfm4Nt3Y6VpfjSivhF3V0uieItH
DJEQp7CfmTQ2EujinYYNyKR1iP6qriXHmaIR5sXPZ/DjOMQHXZqdk3T+q670kI5T
9ERYRnTzFDEQ9SNt8JZ9MDCKhiIT8OEr/BS5w7KyzAw3X1nN8J6Miu2cpQymSR7P
0hUN6g64m5J3/P7PMB2HHc5SsXRuWrAs4Em0IK+00++APswUuEKa4uB9ESMt1CnE
81U3aTi/7/6EE4j5eAhRCRJrtltWKfLwNt0KgbSEBVB2+vL8gsQ8ctoNMCBzaFRD
LJB3TJMG0i8jrOtWsUlvwr5y4Jh/GcY3JnsBZ4NgFogZule0ZxS/f5KXtHCjyEI9
1Vut+hMviHZpVSJ+VIHfTILfk6OPuTFiH3kljyf0UAttlQDBLqmwrMWtiB2gAkFl
BR3vWHL4gJNPqSYRdOcnix4Jcz6LaRnlAwSz7ealYsc693DKFq0y5cAcowKvsX3J
EOSQ07ayMiuHiQZolAhVpqdHy8Yt4562OQ1/RFRIsRci3WLkIhe8dMeQjxWBJ30h
1de+2ahTzC/+nbUs58iwmujuy19Wmj4A8sgChiK7ruFQGiiVDEEqX8i82QnrrWsd
aEh8jXtb53C3D2UZqA3wbTs2a+v3dDZbxmYu7lK62pgBrpAk9cFyT+ol3/rJAcAQ
SsGw0bc2XL3Hoo/zyMccUawosQKlS/3fzJCWcc6f7dr0TZrOc8zOxtv48lx4n/Qe
xrhHoMtHVTSlA2WbDsxlu1bgFsPuFcpns348U/hPNNZ+aYb6o5dbxlNEY1CO2o1E
IVLeRUVogv8YxLaDZLYFd6pYe8cEFe0kPmpWQIg0+N4NMuNRvTXI3CK47qQjwyts
nojQOIKe2W/Rx3wkkUETbGQcZbSiTxq67gpZ/fI+dDppN05J//xk8SKxdAw3z0Sm
5vHYhLhwnW98UaNOSrDGwaCZZpBpvUeJnHW5Hb7FRFVLg69KMvv4ZALWvV+6P5Br
8ZMDHt/359MG8bcm0EQTD0urSBbq3joJIOYUWxiVn2e/cNWMqMZMt/sdmiAthSuO
qUqw4vIE9Y+oFtiyjQKjZZRpvPBaSam8ndT0nfzIDrWLCXozKsyUU+nfyObdiqEr
x+LeXXzH24mShlcfsMemHJNYSoogFN4rnGxj25AbKfcK0bXPLFhSvXFN6A9EXIqy
88luZXtZxeqB4JqsFYpoRB29Wqp5st3EY8huOl1hbnQc8nwCtUFYTo52CPvXmVml
SI9AvaJDQ0fh50MUeWsIVA3Jl/qJ9rr7s0NBzdlPG8Gp9+yqAYyg+XslxaCoa2nN
hF57nE2GCdR3xWZMNDnMWcWyg+hdvY+6u19thAsZUdETDGRUcI2H0tLgwefOjwWq
npqoZ6XQrfeVCyxP46It6e7R0QQ71Blrhf5YyaZMKGf/MrwrKgLBckT+L0SFZDW/
0EfZszuofRxLA3a9HUZbUi0IRVpcBfprkys774qwL0ST4L8M8mETmfmHIMRCsJIL
Ft50NR64cXSCLI+DGYdEL31wFCuEZE9JtBgLuLke2xg0PRKHtVt4Eb4ELkCQi4Mz
ZeMrpWBND5UcOnTWZKpAxOP6PUNHABqo4k35woz9/i7YnyjGH6OBmD8hTLPjx0HX
rIFS59w7u7PvEwrqhJbA/cfyzP6a7Xk4BFBYt3JpcDM9vh1QslebqGONyjh032w3
500OGF0Jo38khFp/Pzx2KQRp42uEFzLzpaIJhkRdz6uFsZBfjc2LdPFoNYunTQnw
OFVIyEbpIqkMHQDDZyierk414MOgkjINqJbJWU6anzYNLhRhC0Fxl2pOkxaooGLL
9txrVlVjMq6jvj6JgqaA5gLvPbHl0b1k8+Cx6BpuPmiuX7Clei8BKWaJiSjDGi11
fy0gvqJH3BXcdr83x9rsfm/iDdCEfAWCJTTJFDtIsCWJiFpkGTyC12w5i5s4BlxJ
wMAQwQrXsoBQeVm8ejfDkUhtAH8z8Jl0TuBeuVmeveZmMhjELoABd44Sa5P6Cxz6
aKt97ZcZT651w67rCwrHFdv8f6qLWdYlPUJySIIxUXAUkqS6nuJP4M8jVJQr+IKl
zQ56UYNzB8Q4tUg1iChRbKomptR8hNCkyQEjNwZpaL7Ym/+hasBv7jYl7Fqcq7A/
3jZSU9LZYZzw2sgmZJA5bRDAcOM1lBTFCsxzADzU9mzK+gtw8H3+6uWJphJ1bOmZ
aGbsMh2tCo1RjCtTB/UyGBQUYBy/OXw9eNZFpbesGBjSYUT0jJKdVju5biBRgVO2
kGGu5ln2gDsR/qheh7SWM7JSAvTPI6w7zl6izj7TENN1rA/x0csj2bNfkdiiF0se
OTBSOtYtsJN0r/Phz+PoCogGMNR5d+9tg4U0/7RhG6USrljzIPtFICTjpmvj1J7T
fdHpJqiCoosK0HASQ1fJzZ1zJAOL/kjIX79Dt0bSePKDJnV24aM0x49ZlqueKEYR
a8sPTVoDYpbqS7/lQjccFb9mn3/sQz/WNMYGSQpMfzAzZtJ8VAE3CG68vI3np9x2
9gn2PWMOT4uQgJolbdmzpcoQT4m+SgQ6gwyNYTHPbWKrzX8Gs59NIViXrH718+jz
HKmoo3aH5V0shR3pY3pAR1I6TvMsQG9FqQdrJVEU8zVNNTV1wJpy+gMtZbnfa8PZ
c2PPaPvXPbnCbaKwnK2V1yPMyAHLbt6cDu0sSZHsfIqUfVyCfRz9XjI4bJ5LPzh1
0VCzQZUOKpd4qLLTUVXJdYNM6rJO3w+V/7Dkb7mWwWg3tJleh5u1EwFNdxRtmenO
C5BTV1Q/lKReJYempdoBVQM+eGU/a2K/25+vd64x+uOp9a2zAc+zm+mGHXy7ITfs
TRLFk4DKBQs50Hb91R440CNkmw5OjvmqSSbRD3X1mokkcDa4CqDqK+PAE37OPCSf
5mrO65H2SLtzut01RqS84T0yQ4iLfLNy50aMqph3McyOm2h2tDvY4eQYjnpum72Q
ToWbmzNuLzkiSeUDNtTr+aIVLrTptA+/B5WPGPuHwHIKSo1PhqyRIQIJGSQuL6dS
D2Oj67HmpIJJ4xP4N91jgtpA5PbnpTo3xxC58jBA6Jb2vGqs9mDNCEnhFNb+PFXB
5gF+cacB2wnxVVQkRBQ5miPRPRD6oXECtPhcFosZ7E4WibxBkeRvqxLvlPK+NroH
UQWXy72cosg8VkJC9Dn3ekFrN78zGHFbuK2XHbSkuAHSV97J9XLxbo2Vm9vmdmrZ
jlR41Cmost73MpHn/mdJKTxUVQL4u6RxxzVwjl3lIbJIuAdAqMvI3B5ItRoPQlMk
3h8o55u4Zcx0AvcbDrSNPwjCqHdju9Ier/y0rhcatBh/RF/6/MsBRxBD60QcW/l1
KiRSWu84DwJ/lnC03J8+c+cVeJkD//eBFUznhfpBqfIdwyLh9jI/+T7TiMusGgah
w7CgJViJSOqxKlEXjanPBOmQqrt60p69P3ku9T9bCZMKk1tLzNnRp24iHGDlVq3e
h66jsf/n4ry+y1qKkaekrpXdFFeyFsJrWUZajOZFpN0dKTKQcyzJPLOSIkEDV7LJ
dDuqByn0uVJrrsjpAqFdI7c28bmh7jccvaPA5CTKiD+ph2koIMRhRJqjemhEwCNA
cIchTCKqB/JK/0wns6vn4XAeHRrrpyUl+GTVg4nlgm1Z3Xgnoac9GlyfTqYfR7LX
xj7PcjFLAHxHkmwUMHYom8LUmmvpyat6YvQ7P6lCDO4dgogfB5kpV4dY/UYarMHm
ZScomywY3caiY4/pY5+hI5kDCdSp3E4cvp4Rb/+Tc4Q9Qsctb6z9ZbNFYxOX4X/v
1hzFZPOy9gLXUVnbBbo3WPclLqyM8bgjOFtYwxNPYRdA4qtE39eAQwFtuhd0Mr+l
kDIyL1SFDE+dh60ouF7UMbRu/FUOzPsYX58XE1LMFPvQ/kbNp6OxerzCfJG3rgw1
d59wmz8alUWDH9YsL48gz02lyB55hZg91/CpUfYkCmXBZqFCHVWvBOlPdJ4Dl7op
p3kdJ/0pGECUFaikUmBQeNrNkSuQGkIst/EleJLSvKpxOH0/Dh2XZDJOE3/sK5L6
k3LDMH9eW1sv+qAPqyeYbmd1w0JKC9kOLc5z60NeuHFq4zs8YoHVaby8gl/jSRcQ
OZaUO3dzleMPuG5c+Hg3gf82NFomG0i/yYqVphKfcc2TydigEoEalANdZt8RlWLW
lCU6bdgjuHn0bFF6pEVnQASy6j1DhitFe87dx6ddH+Lr6I5D6Bjt1qudJg8wH9g5
a/jenVp44ENZ2I+1g7EW16lzfh4ll6HrJsc2L9LBquljDjzjrFrfVnwwryUvRxku
XzZVlIvoYz44UCCJKc6wdZIc10ouB1IPnpmDbDDej5sPYqT0Qaq7q3w2AKWq/Xpx
MSB90iUXkDlrpWgnPTtmM4K9camqkaQwZifuXlh6bhP8nqO/J3Bh3reWPdUFJksZ
TjW44F2fMtj6Xd1GRNQUz3yQf50YfSF/NbHplONJKhu+2iRnfMK07CGDq8N2xRwT
Cg0PShwWNG3eOu2FfNTjLpvbwte61lJaABvFl5tWyOnyojbNNGmpXz5PSunGlpnd
a0PSbKUVEXNkFqLyGNBQwk9JHPbXiaj4Zx08No06Z1d0d4JUc4Z2FeUC9viU1T0z
NPbBE/SJiquwvYho0rqDxjCNx179s3r/tYsinP0mbG7oIyX0lFOqoRSUeKbhAtLk
8ePnYBftaufj4yd8ZwReM+3XHLl8vYbOdpIxDb/DorQar9bZo9Re8k2QZhKD2UXP
+PBNT09guWCWh7/CNOJ/QjANICw5BmxlVkj4jqqjBAa8yqcW/ychqJdVEncQ6Qc6
YfM7iGurOW399GSnOLsSksCiHFNZGC3VlCnZsAyVmzwLE5yhjFuaaeSmZHWXn7wG
jqzbgicIj+qw+MguxigAkDudyd3xe5T5Fg1PLC/uHRunHQzJbXZ3C5WDoId5lETf
HfOjdI0GgUh6VJ6w53/uBecqwEy6TxhDF6jBBVagqgrPMdwnAbbw3Ysogj/Zowm8
BAE3/oaY+/RbpTg7R+YhDgJ5dURugKRm8G2+vIWAvHFlFa4Hq9vnqjgNJXLtc7lm
8nwmOnsNGePbNVCbYVklmH9ULsjdR0qLNCkITDCzfYLDAc7qqoZx8NmVjddZASyn
Mm80Ew7xkR3aFVtG4s8GAnsTTV8NgrbmKnIkU2GhCZEnIh4n0ckcD3OjsYBjOMAB
CAd2EwhCT80nlKCeuCFPb/YX9A2UyExSAQMM6N3eHs2q4VG3LFQmqCrQUFsdY4Li
3LHyahKqzOqDBziDag2GCVU6a+R1YijtcfbCEg4PflAGfkXwiN86I8dGHto5+Xbn
Xiw3k955sfSA011zFYXGAT2ahMe+dS0+JSTJRlwB6XEp7W9SxEZNq9jsr14Jz+Pq
s9rpQNTQswo97kKvrmEQ+79zvh3tAnlMfJczG+WCYJ2wDEIWLZhShAUIEYLIdSI5
qvfCTVcc8oNAy2dLj8n7QoMGsxlF6IcbdlX1D41nXqv8GBpo471ihySNtJyP7WHm
e6H2Qh6hqwUaXmJEdRME35AAx7Bk76qqgWtkCB+5Q25KZIFi4B5efQbeMdVIK1jB
s5DoArPNpx5z0yg+3F6Lf3oQHhCxUapKxegqVTuLvqc+hUmTiSQVpHlMMzAKZNw+
I2mKpuBX/3k47QJ09QpLf/nvbBuF7oB6ZLvWFvaMj3Mmtb+UiogxLH48F0WZkd2e
cpzmGo+zBTNZOZD9R4b2vlfR0Z0WSwvT6RuwkZM49w2Vmd40pcXleG6ENi0UCt2G
WotH2GDqDFSuu7HFh92zXNBRmX2uz+ZTmjJdkqZnGYVWA7WFzevUiVQkqhvznSDL
VslkjV5yD7KHZGu33LnPXhEYTzksrkZnYJGCS3nvZwhg93CHjNXNQKMgz4KRcBf3
/jBA309TE4WiMjMYxvokpQoujP3HfKQ0HdiSoK4toIg8eSNP5V9z2GxQy6TDAwlT
uMLcuBNNQrkYMkay+dGim+ByTl5J8GSbzO5pRBMA9g1XVIDMsCZrcheMcy5mabco
ggOwVznRVxNLjkRT9QBFUKhXovgiwWq5xJedgaKQYmcBGCPYK65iogk7Otub6nB/
rweukjKPn+ckDuNUiNXzrJ/Dwtksv/NtwJuh+my5JDqngQXPx2cbjMOdjlxyCNbk
ZddJ+wg8vIN6ppyV7SsHUSWTqLx8LCwDkHrsHcr8Xgyn+O8nNL2WQodEsy9mrTqW
ufkg8APqfcClExxE06U5ncMbz5Xm0gLyKZBtFtbWwyZHesl36tsDwyfxAvC/L2cU
TcIzYjf1N21ptEAS7nUjXgW1XloVD1qPxSJKyVt/6bkLkglsyyfuHl6LaZ9l2/Iy
FKG+ZW4QOf3Z8gJbO5kFR3/A17ZRwUQN5JntoF0Voo5tFFQtttnK12tIQ5QOasW4
cjC5FvEok60G+2iZiwi8Rc+bhyckRh71j/iItqOhX/+LEiXgRV2BNqpi0HikVSjo
N8xdhkdsPJCaYT7x6wH9jPtv7zmCUJ/XQ2/i4MzdNUODkGf5gunJdttEy7w9FSDQ
oCi79v0GfiLb0x4SwS/V2Wr1cjD/nCb04eqgr0NBhvmzL1NAxmkMrwntsRAi/PYr
bUCgZ8GQGw3IvSARhvUwrXtIRgKrpPWyVymfNyBLqwrbxoynhJwAzDhQydA/CgKb
BaSMLnFwBF115j/HJ7h3mhIlNHAMv9nHG8fJlxmO1S4u4sXxOhS/FOjFVk3dG1fn
GTnUakygYbIRwdm8D+aqzKXOyc1W+G1qKUqrAblY043x/1QUVaps4UUu8K0QA2ni
oLn5RZzOFcXCAGyUrWzhLyNVmN0vvtBYTz5NkCDidW8xIzrzp//kBWRsWw/5ouKd
y2ZF+e7TF/RNqb4RouT6XaXQaB16d+18ziC8jWLPrJEq0gUr978pmEK/KWtg6o0X
gc4TWkZCOfQtdjdWsDNmUkWtM34AvmYNvRbXwcpuU+VxbnWUc2LtO1hfKb//xA7L
3Cs6gb1mBcg/QvBB7g9zJSnskIO1hRszevU1F3JczaIFUKKqRs5yXslq8xk3a9XF
pN0Z/8O6vCx8iz4rJkRbMBoywmoE3rsy9oZIGRdUEtYzt4Nn26H7IDK2SbfPH/Fk
mYDQHhzPGC0+w1F/arp3+34E+N5wdo1UH582Dpu0W0YvyD4K6LDmSipuov7/tRyi
i3jRzYfuxKNkyZbZRIW3rv8exqFb8eNG1UvO3PxVMyVGsXKVh7lLhYjtc4hMeyUz
rVAfKxWUh7b372PTJ61wTBgKzezJbtpnP0gQHoFFo/e0+CJZo3EjuX1cuT3V3aXW
LZF3GHtJcPJZZRKuKwmCJKb4J+WaBzxgPlm7dlWmWKbvz3Z+pQSMnmEwfVUIx/h0
vT87pMzn4StgThI/NhYLl+FufkRzKwtp9NmvrHPvfrc7ZhAuDUNRK6KhaF3BudcB
QX9wdf0ZM8vX5d5yY/vzoaWIkrpbX90CXlDbD/9qckpVEgt6FmyxsWfl3zmd1jhy
9z6QDKgtVJr8hLoKEqTkmdj/4gxQYXGmiCPQpsQh9ElvFKcnUXJG0byaGG934Kgd
YccRh3gZQ5rmV4aOxiyV/JvPkQDNN1TUDtnBYziIO0BmhRxzN6ZGSqOxbYuSna01
IQBtbckiuSX14HVt5FenfYazHHFZZ+5AwZGN+jxfqyqDAwwiZpF/R/K7iZNreyGh
jW2D+BPuSIBhxQcPzVk49aenBrNvHatUkAgiLhiajquvgVma+CD9Vgv8d4N/c7dL
WkJgHs2Ju2kCBGBqjouVnC+qqUqbxyWdKu4oXVFRgZhsWW/HmRi8p+reXFNb1Rva
2EWiJhPIHW/AEpnoEDu8zUf8ynpz85SwR1RgmbG3lIBJgg64qnEW27XgwTdW0c99
nBtwa9FjivrI7eF5W3RblfGG8k3Ar3sAOCEv8s8QN09mn1T+ywfxZ8AjJZNkI4jk
d6W6gz+uJ9OY5/9YFnh5f48TvvvF3u29UFJQsBYkmaEISNZmdxt4mQ8ChXLHXUUH
vWq4VaOZmZWjpSPRHX9s8Nx8bQ/oGsoDQlCFTi2l1xYPnVrR28KVnFf6a3/izXb0
4Pfd1Cj9A9iR5LvuvevaITVJAn3UIJDPkFVh/qm5y1FWk/l61EapyFJEcMqA2QmP
zgvDS3BNzSo4zGiVBZGXiI8MphwwdIYbfpyyuD5ssbOxAXZpVxUt2QPQSOlQPkQK
k9FC0/FOzp6ZTpBwBtPXsat3Iue2FMZcdNtrnizffS8P/j654qeObsv2Sukt9K7G
dacgfBRw/oRaI6aw/dQWszRwl+xmVYsANaaHC+tCukz0kNzLA6ym4h9MiegiN44M
yqcChRkBO7JDvh0auRdP9Oa03+XcLqqdqFDitnAy0ZJkZWkXk8aHxt+d19eg3YdV
dliDuUXt7wG/rsRrrrSlwRG7J6a5ezc4Qt1kL91LL70ezNv03LEtaq1z2r+nhNBw
40A4XGLVKn8taFKYeZPfXPVx40IxYpej4fyktpcplc1pUdXx3D6KxTMEIq+6gJVy
0Kvw0rMYPAWUcBemxRK087dZKSzm0WLD6XIhyWWWNzWkP71kz5DaEMcPPO+b3IKF
3A9QaB6mAgWoD55F6iiQjLf4KZMGZhn8zio/wl8RTtQj9aexPKcPEmsHgBjyjiUA
NHljlqzQWlVYI3wpJizrCbJGGEwkClcuBCRmesa8ovsv0VLUY9EtJsS+v0eaPom4
J2Dg1rHaaPTvo+p1vWnx08Ob8JZuXrl5pOfGCPc6J45kpnit4tvAZ8PpO+9pLdtR
wXVBK75QVyTLwVGCf02BKv4sS6qTnw4ooQZv0+I4C0UcMlDjh+h/8X0A45CWtuct
IxtY0sAoQ8vt4s98I4DPePYjFqmpl/lD588smXsoMK+WGYxxSY53sBtOQHWB9RSG
wXVmOnOvCdyYsAaHMJo+Vf9ZCyaUh4BqqTA0wcZxQ/OR7HR8vRTIIyUBpbZk775w
IQ4uehWeGypyqNv0/lYbrLUyt0E/albDbDD1p0FV0hVU6S3L8N8lj2G5WOlAkdOn
9s7TtLSPuB+lMpCOBF6AnukvKqtRWds4e1xyjSc4xfCSOSrHe8VbzWPpNnGzFZDh
HAZ77d9IVhdb91M+UL9jpnuPcdUvz0SytJfv5kc9C9WfSv70yuxlKBQr1DM5KD/a
dJe6LK8rk7Fv4BA0qwr5Y0rfM/RdPChj4du4lQ1jVhud9Dv0iY0JsXBN800slqB+
gO4HDYJb6bOkOY3NpFG7lyRd+o92WMui4CMGoFvjpSg891dZJOyxQyusdpphWCUb
XsbI9cRk4/HgH5dUk88SUJGtFDAmVnmblRQeVmSlNby14mB4/H41uFqK9sfstRpX
+TzyaGIlCcJqIXirVwFAtgI15HO4+1k8LsgyWxeI9L4irn9SDzt/ugL9ellisNa1
yuG/mjN120r3puAprJ7k8HpJj20gZDD4wGcR8zE/xGoyujABGWU3Kc8WjCs+npOP
eH2wtZHYFxlrifRYcxoDYgH9qTw8qecOtvkexCYcYBPkp2sKUA7QsFvD2SFedcjb
ekT5md2v7fl5fEOEeFPBwzdj+sTnYp19CCWnmKN0XPbOD/el5B3d30opf1jgg72C
lggLvZF++wB18o32isFMDmVWpYxTdYPbDRQGhJX8LnJdAmYqaR0YdV8q9OIiPZ3W
hnNDkqjPT5wXpJX7Yz7o2wfMOXgyrG4naQeRBZVAvWKD7dgPihIc5qz9Drun/p2o
tmRsiwzFd/QmaQt1xC6ZZ9JKz0HwBbR50c/YYro3epcuTd6IrqYm6umio/eKAkU/
MsC3pxzxTsx2jhq3wueBCCufI+dprfudnRGGHgQrdMClUQdkrMGpY+0Nb7CY22wL
/PyBpqHeNl3gmlJbaXOJY6IwpwYDAsBskti5G+wHT/hdu1XUD7oeD7Ueji9u1C8Z
cwgq9nKcUBFlQy443kXOcOFryVKJ4B19mgSsH38WITFMGeNOXDCFtVOxp0A91cRe
jYpjfMt9kuTCNiCGjdoT50BzvBpm7/FkOW5Wuj7OV3LKyJcaDIBJ6fXAK+SR/53Y
VPb1XAdVQ218OFcEdU6Kf15xg1rJlY0JitAlvzTVg6KleeLy5enu9bVoO1mGG00C
f1bi6mps93MgLoa6W7CsIv5o8s0KkfZlgCKLMP02PuPRNOmv7Husv51MOKWTsFSo
42vN9CWgc33Blr4Vgw6rvIFBA/e5o3SGu/BjX6ysms8Kxto3+PPu2qvC6BliwvFP
vnML0A1Fi01LsB13Rn0QP7NCkAlf+71Jt78IOr7kdHYKzltJbjpiIApWLxOBpF4h
iHu4I631sr8sZfr2XGmTTnB0AkyN8JKC++BKmjYZTsTOtTrn/i81+AeiSsYcQn4p
gV7Zwe/A0WfwnHOWiy5hZ7f69TAc085Zg9Cnp4y4HpBGAtF1sN/Hf2pMejidyR1m
8cOydZomv6cGYVAj6lwd2HrvpAQ0zwz2J6TqHRfJU1hfsPYP7JiNp2jgYpkqEHVN
oVmPqdKGHuC8+2QBkPN9J9fXbfruuh39k1c6Ofgw4Im06yuO7ATgU2nM7S7KyUiv
pyNZ1ue49CKNunGgjgtpyi4b9pWIBzQYQdLEgiA2e4PxC+zzAHmZi4dALV6a5EMr
/b73gQzj2lFTKovosdmMdTXCzyQnUn5CAaHEO7nbRG7esxCLr+JZR91PAMbMEjjj
D2/L3KLWsiMiMx97mBcwUHc1RsTHDnuzvL5Q+0zWzTS7uqCbTK3MTMY/JDLSoXUo
vY+GaWYjCZUKIphdKHbwFC/bNt6tIEpAdSG1cRjG+hsVQBH+vc/bNJdyuB1z6xb5
cbIMCT3rbtZteQUmTikITRv4des+I5fJggeEmo/GjBg3R7Bw8LuoxOMA5BtkYHBX
2PIxhLcBMkWnW9iBz5mPGQ22ij90No2mlq8b7tQjK2NNwXdrCOy7TIVxRRnWGF0b
biCecIYv2Swx+2aVGp1L+8raFWI67zdAA2gwCaHBMsw9J94Qv8xOZixLlZ3/XRSU
VTqK2qCxKv+I8+8tjlmZcRXndTwoTPu4Q4iOzUqiV8YOKcp8cHJOQpINuvp6dQPI
6y0kknSrw6VgZ0q2ZJbnjTQnkV2/g57VlKpFQPitEUjgHs0E5v8WLrmlQsFeQGuh
EHlKwP4NwpdXvJr6VKv4rPFaZ528tAZgcuzPVPsnLnqSqf5zuUFVraFddkIdjeDb
g2C0A8uv08cy37zXhYZiEHlL6w5tNR/Uq++xBoe6Cm0tufcKCNcTEc440O3sb+cJ
hFnGIcuCwdwKaZJb5Wn0uSM/WWJkQJpgPD8NGQOsvtbzgrV4JptTYkXxkLHz5C9u
YFyseRgTDsLCimXuvIuUE9idMkWZD5J+QU8g1ELDKzrCCMTK83OVnX8qeM+7CnYz
nKFSiP7xn7fEHRBc7kfeSfzoNvvhcrwaJXfIYikv5Rm41TqNa5D0JwSEBjw6M/3J
pRZ+1xEqryRASVj04+/9WWArlWLPixRG13kkIE1T94hX0cdwbL+/JPikWslqpEVi
hnJNrU9n0uunj+PPQPdcs87EiIX/aV/sA6kBzhLMeesJt8VFWp1eDZq16WI0ZZPM
YhARr0AWmAwYv3UZWi+RTOcEHmQGmu7xi3OTsiM+XJ6NjbRUue9ncpqPfM+M1mPF
PJEGA09rHRrUZT1dLNvBd8Yn/9PSUABYRZqh2WNLQhKghL+jcyyIMFdgrJgszxZu
Ozc/UjtD1pWgq2aNNOvG7qiUIRgLZgysPHTDFjZ89Z3eyN+F8wn4yuy31AKKqy9E
m5j1Z72ADvBOcl9lsc3SsASCGomhTecAiEhaX1zeEpJDb98zWbl7M9+Av/rQFUy0
iVRPRSHr9GSphy9VTd0a0nXIyo55h//kZlSyPHWSG0yXRtOHQa06gwA1fqcJf+8G
JrN4SkrPucZHJwqfE12/s5VO3VhRS+gWwNHTh42Zz0fsKaSUhhfNA5x31TdPTJdd
jhW6LM4JSwjTfllF8HuCgdEUfjTLdOOY3XW5ffUbXeBxNzxNhSOVSKDHtMIRC4+u
VGJBkf8U8wr1D9JGw1QCCcKfKLXk8WUklwuxb/Zqear9ABhWEt6m3SAKivLnTJuv
cW1osFEuMCW0mVAcThgPjSs6So5wnEz3qmj6LGgxM3+47/wojbwZz3rLuoDozlre
91sjre9O2UUH7mxwkzGvV2ZxcRyYhRFJ4YoSOeyEhHseOxV+AkZE1t1+rNMaLf/v
mqIDE8srVeAByGEPeG609ZfuF8RFTIIx9j/qslOSyIPxYPQP6VT/ZYJ4Z9aSGi8O
FpeofJxbqW7v64wuxZZh34PenZUB6XebDh82G9Rgs056bu5+2i66Zj01m1RHfSNe
1jWUvAonhq7aCMlYSEuR/HotQ1qO66yMx7pvng5IDn17Cut24UpG1n/EhzsaK5uL
XUvhoCYqmiTzDgMsvDzcXn9+djjr1QgPxkAW+HTIjWRfkcwAPIG4puhxqug4z11e
DLjrM202H7LxL7WRvLk/9qJXQBPITrZaW32zoiZkifKAVGJ5e8n/UKI5OqGfTctZ
dBs7O7mFdYOKKYsc3oDpD3zOLy4BW8pmgrDVB8wAzlar24cTspQav6+C5orzrLij
z2M46HpyuoJsiKEm0heSZygrBE+HRjGXZEvdiTrf4qDhwA8aHghlo1kffjDvJjEL
JETGGKr3ZzTzMB+7A4q39IPD4k1iS9kNs55aPROyrciQJ13m2pQiCeULhmUerSjc
q5P+NSotzcqCiEiPgkrI/5MXSb7szZ3xKub5jFAmvEztTDdxsfcLnjW763ClTewY
2qawnTUaCEHljn7tVmEEclgcScGbfeBkOQew5XEqKiY6orlyfXkiLvHYlCVU7+p+
X4GrK7zJXcv7RTARJ4LOMUmeCMf0IdxBiKbiAFNo45uO5HujhkwSSGnyKb0lXxnc
ceQ7QQ1YFj6ixlCfgpcQap7GSlCzBB7ElRpgSUS/suD6oPqGfNpAjvHZcn2ElX3C
M9ENsLPXVheF6kGUQIzAYLE4zwl/gn1dljHZ88utykjj+sPQQTHcvCyfC3HGWZ9z
KiuAIGEouMU7aJlz6QAZsGTVO9QVC2KH3r+SvRwwtdgnFpS6PvqZaEyExhm6sv4H
Dmy35jJrpF9G9Pjlt3agVCeKHe508jiP5ks0Z4Uj0K1nXMrbzXB8ZRTKzenecKs5
EGJ7+1zLeJFE0Hl0ynDU1YwTIlC4PaAompEgZPyP0xVFklcmO3VHGz7zcGlcKrqr
Tt0F/L+AF8H7n9W3t9802LCcTkPRdnXNlgQkfz5PrYbBmUMumdBrwyBFtZ/qUwol
5gl/pyrSo0/YsSbbZXBfkzr5E4rp0ItrB9HT2IqZYfITajIk10CL7ENSmahrKnAx
46ligfz35abtz0h1PfXzqnH6cjPjp1eYNHkz7jnxLbtEbc3Ce/7F41/c0NmfDN1z
8vmknB5zEWDSWQUP3tTkDYdjJkVhWclywH0/66ZZFbfbJ3XkMNEfLVevwiT7innF
WGC0nC0tzN3zInMVSLdGuxqOVziSvMZtVAiOotXFj9ElyvItCV12FyU4IWo+K/Az
yBwihmZDXEtHgEaDWsUk/x3YBgkve5x02De97f1ruHBYcoxh/C06CU/y4+U+kNiI
73Hg6ntX/4BZav9GbB2Fmj1ioIjfJ5nihij6ibZ9CnL3j3mSYZI6iJE57U5mfqSg
Up830JwcMONDo1VGn5y+ZWjfQAYPrgU+S0EoDUufQBqudb1WXuwIT91FSeDUboyB
nIBAVJNTgfnZR8wJNyVKU1xQKMbJksZa0Lp8gCEfEN0Ili0kH21OlI2kwJ/EwOYi
t4ggTSV7OTlssoFWZlelNFgct6+5enmFnKCFTEpRx2Ky53Osma9F5/sZO/DdJu+E
qYAmJcuQHCpuZc9g1ZcO0Eko15SKfQPw7H0IjeBMYinGV08k5UCZDfoHzYuCXVNT
6OqRh9RaEd75iWyjDFEeY1iH96oPBLNvudy0X8oIMSGMGUS8hzKRSizQvpknx7iI
bWL+NO12/U/XHAI9CUG/dlJWWCpXRvLfOWIOHbU5pE7tHKuYS557CRHZH8GLRPLK
HWAdTVzvmkNCAXqJcjY+nEcMk7yQUAyHC9Q9ATFfugE+RH0a8mOJO/efrldI4ATh
R5ZMPWGjiaR70xOw6EF8S36jw/jiqPlKi6w0olG3EuVlIlylQkCqiv7Ypj9Cqi2R
ig0hk0m6uLr9FMHlwrDpktwW5uOZ3XITeQTVe8XpC72zPkbGapRPPnk4kH3uU6xE
2a25TxFBY2ewAJirt74HV6dfdDMTO59BefyNk7kjne9iCHPQXBAjllNPw7Z2T8zq
zAsX4RzFCPOxcAKSeSOBturoAer9/LMNdDX2pbcSaRBu/B3iKUyKDbEUjCJcaamO
olI5R4JF6GP5Lv7GRwSW5urrQ/47dKW/vKIMylKGbNBvTsE8qYBZa/cXzDv93t2Z
+7YaoDI0uW5KouhQl0PFxm5tOYxAO1zyp4DOFT7jnJMC+Owh/ymo0FFCEI5qx3Vd
xOdHkdAfB86jHgcXwm/Ib1o3aAjQA9s0Jlx5VaOHlVikWi7io7v33uyWm24IGB7/
hTmiwOjeUGztvaAWvwV+8Xr2xRHRbr7WGiojw3O5V3C3G10k0lvaazzREd4SpRYJ
CnNCOCVuIF8S4tA96RnoneTy/LKdfRJlxEHaBIbj5it+l9bUDlzrW5Df8hSVum7+
HQid2XCkYjU7wIndouEOEcrJ6xQ7L59+nlQdTXT9vTVKb/wXs8zpogAoUj3gN5nY
IAvDoG46gX9iED0PJx35WDb3HwjmNIWMW7APT8VSPNa3qpddfheyU3r6ezO7sxWK
3UqKISwVvct3yMx43cFnXmCERAljI1sNPoI3swXbzzt//3nYAMdbySvbP+Xrnb3l
hm5giehTCIie/2926YF84isb/by8DOC1NF6LxZT3SYao/rpS7Lv/9Fa3YfIK7rTm
1jqejyUlpK2IG+1hQY9CoJR+ksSM5psp1rwIMHjkft69/HIS8IibH6CBYwA5+iZq
qcFOH2MAduBp/jSk5FAFv1cNEPhkCWbNhUrcmv/bvIqNn+2Sqo7Uutv9wQ7vA2xw
LZ1dhHvWLU2FK+bqj3ZUCgkMNwGdKEejGq98YtVfmThJYgp2AhLl7qnK39sUX067
qT6FM9Suw3xSc8WFn/jMQzYGvLbvOwFLM6wX7Yc5DvBOrb6QP0LBBEw6bATzs2aL
LlLeKmQUTGyBRuvjLdXAbO73Y5mh79a/Y3StB96k5IHXHO/+N+fa+bR5YV2d+G1j
x/TZ9hu7ZdJnwQWBjGW88/XwQ9dhuow5NauhU1B/qvDxJpSYPCx5vOqa97P2WPcj
KSgkjTghV+ElX4rHFllvv4gmlBwZoakRT4IJw+tRm6kkCflgNbdAK7SEdaDBlvh7
HVDdSgD2BJKyHgIoeiE48+RWpc0tbnMoWLeaJpSDfQ46vOOoEGg14ygVMWSzmTS8
6Ry/FanWTON/tOM/Tei4GZNgy3MmTnJGIS0sGAZrEn1EG+FHIwjjXqKKaoo9BUi1
uyHo8/cW2Ic+gKds0r2RegN5C1zf9E65V9dLJgyBcH7nouE+dsGpao7o7jpIugAO
YbcZMDB+2FaCq/Bg651LUYLi3nMnTBzkt+f+h7cU5kABhHuMcGT0TSVb6eCzYppB
QfXB9MM7JdmjrsoT2dPmsO2o6uVjQlzdkfLPLVbU29VIElpbQNi7yKGJ3A8IM0UE
GAYGxQpmFDbcLARUo+8Is8VPchK49Gfpv3XGxy2MqsNInhVlanpGZXY8zl4iN6Gz
bW4tPdJWy4WA5mxryE7vExdQXv4rp5D5gSKfBRbslPnrvO4cSvS3FnUVfDwsYX8x
2dfLWxWs+jJ9HKJc7xXOkfO6Hlco9r7DKDvGGZZRcjAN9jDClVMpGJidfSRj/Kt1
oQ35QI+OoRUwlHTMEd2qLB0ACIAfmEnMJjzr80xeGdPcSlp7od359woOzhX3W+OX
999YoBbWC8NOQGjJsvP9mnCWvEeOlzuopjzoPfjizigSUl35wbQNXUKll5xjrMhT
OBQ3RGe9Hyj+lEd5zo6A+o9AXnbh3oJYAXvoGoZfa1NSwcoUJeKq9iJ2lzOKDdI+
Zodwp5rFAzQZNb0eHuV3oMhZJ+PAColw36G33tNvEYhqWGGjQFiIb2IG6zGzVLuw
8JmfDekK8YO9l42XwdPfceH4Q6l6xFvxnzXObXN61nsefK/pQ3fFatD7eJ6fKpN7
QUk0hU5te108snSNQXwu+Mq2oXcDGXSQrv/fHVA0D+AgwYrmq7kKhaYOLLLhsl/w
IdkgV7TnE0Cr4Yg9K7hkOb0jBp7QPfTIFB/S4NPJi8mJoy4SRUXBzUvf5l+pHPPK
rHwFvQJAXYYLa6F9PxHFgk1tHU9lka//P5/jaYbxn2PDZHKH1vRZWz7CoeLiMCub
PW+wVGdHlvVDsd3QVN9dQOrGzqn4msgc9dmQqheEjc6+dmo5K2KX2HMxWWCGXG+A
w0jWIik2fj+nJxRxtzkFd5MWoDrV85bmA2S4j85SrjB5CgitD6G3T4NUydBWWtt1
SiCG7rKbhF7n9gZtr3KNesdkFzDoRM1fC8JYOWrtfbQjcWWoAlkI8ApDhh/XupQb
ZXt1E3txzz0Cn1HiulLElGEi2iOEbxpdLaGYPaJAtUI3b0o3Gy4h8W4uHw91BjVJ
UC5H6RAsd5irdCTyHGQKR+cgQRgC70lnvde/5NP1oEGgFuKLK43DxOnUfGbymwMU
BTucbHnZCi9fiTDDQlyd4VGTOs+TTNfRb8jNnWVYr8u2wVgwTLIwOocpTWTAcQG4
da1J0Wk3MMK9uaAZAiNR1AJvfa11qmqLYjwOzaslw8915SgZgOGaitDBc1hWH60p
f8d7HCDY/vU/kVZlh7oIB1pDJrwWbruLymVv/iI9nbZeUPUtBr5qmxQywUesh4si
/rSJJ+wYtheIDt57vCNYcV/MrO/T2mN/WoYN+H5uEKZ8FQyA1SbMAsWvHmPwFuaM
h5m5eTf2/k2XUyNMvZGn2pTh3yfPe8mAVQ+Lb2B7b3zrAGAvw4wjbdEiI74MpJg2
puA3Trf37M5DVupbMqtv7SctzfWD2QPj9bQ8jYbZZuesAoXZXpjwLWSNlITzQ2M7
OEEqmpNLI9QdoJxKkdublUb5ZFR/046FTIz7ph4+8ljLYh8P6QA9jx9lWFTYS/4Z
Wr1iCbLpXio3y5/pW+0XEjTKiAQVHGuH5/cAiX6QsPCMK3/bKtY/xculGMbcWyS0
gHRVgTwHCYBxHiIhabfu78WmlUuHtV58iI72/alYBXnizq+tBUUu3sqKLKgBCdLH
UNEbDe4JtDWnIBFveafOq8s8x3iRWjfZl74WDCjKxWkxFMLBy/4BgnPpO9aAj2Va
8mhdWfu8GVJ8//ar8E1qAmnugNbJoi4Jl8FjhNFZvsLAnZp7L5mfu5U+8dg2Rpq/
4MUePrdDBvndqmlieKEV1qCZgGJ0zmS2PX4HRkrDjTMJNE6mDODwmyK7STPlpYIQ
rzR9MQJ44T/2i/k4KGi5dC+J+BvfDaic4on2fgdf5yYFnrB9Hw7EmzO9dmNUJ2he
g/D6zZQxIDD4uongsiazrrejdcbng78kS6bO+v/5nRiUmOhizRRfJcMOLx1MuqV8
ZH+FztPn+jBxpF+Own6LK8WybX+oP1ezw2KmiWRfvbCoIjl7RRb6E+p8H7lAhYFS
j97X6XU+SODUJbEpzS9MbdSjCup+Hvyt6G54IDT69XDVKdoQROcXHyFi1h/WXH+R
Zg+08M/Gs9gZzHhP8IuVyoKkVqedN9EniT9VA5E1irEUrFxUXKaKjz4YOWKiqlQs
eBJHiGG/hwo6n9SeIudQHr53uRA6jgzHYIGSexJlmQT9TCpcNAtARXuOmOQl4aLY
+SzjQGgixpTJtGlmFWvv7JM86v/kzhwi/pV9uaG2mqEdBezGhsFOv9ksRdh8GiAs
cdEVbQyaXILunPWf5GRnZMTDwOaA0PaEXQQfR2MG3FLchED/2SrK9cBOFaVzLhwv
fL3ehffclwxDDrpV7YmoV1s1pJybUGBCtEm3LLgIwxFZnC/38GL7455RmIdmDVRF
Zp6353La0T4jd0sv4VW1LKYm4NMUF86t2b/WYiGCt9Qw0wHGwQWyuh1+4nlDfMi5
XjxOrMsUyjLrwPTFrFaOWk2nPLDgtBrj3h4ZjCoi+6mFOpg287q9rAWgfS12Eus4
2zpzuyHGT2iVfh2XmMz/5Q72xawxoY74DhLveakm7k0jRbz5k652u1rWYwQ/2hTb
4wwVRa2XcNtTusbcwJsaoUy4kGAwZGF1+dcJKZDP1OZhjbd4K/Nh9t3mKmgvlhYT
y6MLctIWuadHs8PL/AKMy0ROv353GeNPDBZjpfEXHSeTJHwIV+53BbqNzPquveRt
Ec//A0jy+ijYrA9KAlsvRUxHBx+kBySY/KBFKKahX8fRjnsBB+0SDlIPixFaS6Gh
DwbEQWpTPDLQczRAq3LjFs2EUyaEAtqHM8ISxYoTy/2adqwDhAGYJGXgQGgfODLJ
bw8Y7YP7p3pwDxHg6bk4fXbv335cMj3x1S4EQ8NOMsNfaBSlpfB0iNRi/lmLzWhN
KTsOXbn9qCFDIGzgJ99NSW85Vbsr5YOj3z5QG1ukm5HLQOG628xcdSrKkiw/spBz
GDokgKFIOeErsYg9WZDPssuMaTbST9dwsbUzd7cBByTslWkCxG7nbj51Irltra2G
J8Outkx7XXPo2bfBhUq9Et9GUJomrU+gKEfbE24mMQ7xezFzlTfsxp3P4cprd6EE
h15B4UBK59jHviZfad+vFkCgpwTXLKWNrtpoKtdUK19kik5bBjYL1zis0a1CWQzN
Co6la2gb38PGTxOHW5ip+600ZeWy8LXYUhSIfSCitmKY0pw+cMJY4gkCgA4ol6Hp
mhb7BH426YBXP1kPJb57ZOxEaGvu3u6UAMGu321kwZ950mmH3xPFZsKPiMR/QFxT
Y0tvkfstf1ZLgEXmicjvwTQ74aX3Rd+spVuuIDMs4kT8FaEIfLSSeBGFilJjLnDS
l5bGnu9rJWDGG7RuHv93OEX42Qbw3LipKxVot5v+lJbV6ymMw41YrfxKoIiN5qZe
0JnVnNco5y7u/cVdRfXLrFWCfeEgNRGKGdBUKCuF7oakASreWPz5Hl/frpm+J2rx
uP8gUTkduiUxBvuqf5DNet+3kIau9LXz8TXVnDxNaKghi5N/W/Onxcg/Db8d2bac
2FR7SMqnOr/FOOjjEo34rYpr7sRyF16xcrd+EyXpUgFYJXdIPbciHD9xAc+5fMGM
P6kKmKFoeAd9CPWJFDTqOylACYJM0X+hRvSw6IyH9pzKD3MAPvzClhMEcobdZnRg
N6F6RbP/B4VtPmSH0Wb6Lpio7CRZnGJ69J65Dgu+yD4IRQxRo8Om26oLqCP/hpTc
AzDqXzcbpakQ8WvJRAySiAhkmGDz2d2oqZHxOEJ6YHZtksqBQkAjh1dSFmkIZ1q6
DQtesZrjbvEQMJytlcD30HvP1hJYO2WDXADvS9harWWzickIheFr71EL1lKgbUFb
xwFDVyKAhooVM4TKJQcbFfsqnqkJFvtlwjwZgvvhJ6VL+Eap9GGEkotMD3aEX5af
1k+Q7ewcaB857BJfBSgO/dVHPnA4wgD97DNZGR3qPzjx3Lld13mzGvubJ7iFgJin
vTxuRMJ/nwXzyAaBKNK30Fm57hm45SGjZGs8JyJMKVxdlQzbyy4XS1/UUWUPUIkB
PE9yLXiHPt65If55LztA22eGY10auVSO04FcjB1DAVNU8JmWpKILpLv/GJd2BmCd
+Ry2eskOvEhrf1XEp9fshVXkO0gH3N6+9cUv6DhM82ceoHwuXeIA7UsyyfC8L0G6
NfH7yC1S8q65cbtLcVWyXZOvK9pTlPg1GYQEyHERNqE4PSx1yT146VTXS2Z5q3tS
J1u3wor4yDdIOAFBLHrcoCHQCWJB+4IN5MFa19lv7S2QHDMaQh0djPAvcXEXahyR
JSIEbo3+C42HereAS2KsLHis1LVzbxOTq7CjgFP857qZz3Wi2SLgUGp0a7yK5daL
qCyRO2sxDv5lgcjsMV3LANJgusSTe9UYUDHftOn9xBlYl2Fnxt+LebLt6XwcT31Q
3lt+FUCrAscJOHptw2pBEaFcB9Q6f6vXOO/EUT93BIdYecCoGMDg5xtJXibPjdp1
wfQfvsn/ICz98dQVUKs5t0Z2HADLRkQjnv2U/o0T1TrahD//w3U6RVUqfXKXwbfg
iaE889vBPnOoQoPO0/Q2v/6tLk2z+uFJfSGJjBbb5oFwpdHmIuperhP5xam/pHu7
ATFo3HRZQyz7vxJXpznfAC7UcxZyTThFzkSUyqUUb0Yy/zCFE7/CYAltptyHgkT/
rf27oba0P3SsDJQIqVfidHUADDeUG4wSCuQ1qbYBx3M/8CEhGzkfwNuaaJHEXgyD
E04NPBjTLY+982WmzPY0l2j93s5EbHXQhoC12Ieeiv9qzIJNDUJzgB3YiY6Ju8xG
vSrBqJWox9kQJcrp34FnB7v+USHXdBMKYcazi+Vj26b0f+gt+oqwxNj2ZglaaV68
rTS+s0IOWZrss2znZ8yAReqZFdb6/syr6oLf2+gaYmLNQgOFlh2NMV1TflaLW4uu
vWYYZgK0iDKqIofhiv4Cv32qM/PfxJGDgwEz7kf/Ay2ZOvE496BZHe5/vfXvM4Fi
aPJm0yQIhyfH3+QfWkPtbmI8wfb/Ui/MXvFz2P4FrlW1WYr5JZO+Bg3fzgJ0vXR1
hwwoiWs2vq1SDYUgow2phhAVnDK5nOqCNFpqZGHGzZX7onpaXmjDCO3yr3bvZ6fF
g/FmrhUP/25Jt/lV9M6wR0hxaFTzGkBJ2W8eX4x8xWem/d8Chg27BcRQoLaRI5gb
hXDR6n1X7Sk1mcoGpopm8VhDXtDkoQu2G6QU8F5xbgCH5rDj6Mzdzof1pG90UlFr
AWPnmTE4EGWqEmayjyEEz3RmYsfXFXRmimyIxndZPecKisXwbk/Hpdj8fQVxsLus
DHUSUo8gHLCqv4HpOezjRebQAnsCrhUwfGm1ia6wUJlSnrpG1Pw6DcI7PoJEu9iN
DIRYxL+bi7BltA0UkARBK/8PaPVBkrkfgYcOArTdHOcZ7+dOFFVjx/Wgk4D/R2i5
+UNfnzi1MNqCcwULFhu0QUZB3fbzpjXCwxjSysro8oD1OjXzPDbMlASdniTbvHmk
dEU7wNm5/5RZpzsEwDmn7WJPuG8ASsnBv/TtW8FVVl5pBIsamUWBK6Z9ON27uW1h
pTw7hgZ7z6fbRP5n41hvKr919LNtferEd9149l0J42kyBd/u7hc3k0R2/aJhTbx0
vK4JQmbB59dOMq/JHZyZs8JCZpXgW7+C6EnRcFGPd67GTUyqbtGuJjqlfWX2uxfj
OGHqmabEkSl7irKWSiF7emcZxxbDoaYYI/J+0xlADz9jIg9E20lKVmaA/qRxz+4J
ZWwLn2R3VvZypqhDI92YB/ADLKPR4v4lSwGboCmaRAqLsQh/4vpzmbaqcEJKVAZx
eNekQ+6+/YhFU9ooyercGK3kEaUMb2uBqbko9ojcAKtIstCrJPbWCDoYnrRqZ8SV
xbEOnC3KWTV98VRZughP7dxNPeqHHp8RuOQq6I+xuvaIEL8lvZ4su7qMNAHIQAFp
1yJhYLSzUMo/bphQw8JHSm/ZuoIJ/4PKxoVmf+ZI2mx95IbhKNLG6J2NQKQhJRSe
v9neR8M+A3owmQxKfcWtcc0xo36o+8+hR7SnupoCjh+NHY6akcxfchDPRtG7AZrQ
mUiKb2vDKzwP58YWswKYJ/Vqe79+X7n60QUsFG/uOQzvHpEEZ6wgBQc4b6DZvwCJ
tIENGQN9tJsz/AGlzhQVLvW6gbK02bXCvUW7Wh6bcutFoSVdHiOC9MqbaceOTK+6
aZBge1GYHEbZwFLWNj/9hek8VFjQqu0+h5L5+gFIdoCpv3JyBE0Pv3Hg+sMQeJLr
q+rLeJQhyWBiclhWHhwC8iowa1cRxRZYZ97LWpGIUTe43DgBIksVHBzx+c+SC4Dh
ecf/NAhozVzSir8YBcgsEc+uPHJwDQQA0kRxE35XpeskQEg+TN3T0JfaxkL+W82D
YTOvCor28tMV+22Uie1lsRGgkI3jrotPJatheXmK2VlvSJ0yFrodFDcktmQjSD8E
29wwoPB3yAC+1t/PzmJjBlpPRHHioTVVIS+rSGnvD8gjNGGWizqWowlGkoZXeujx
BAUswFjMeXK/cOsZB15btk3LpEi/tQcpQTM8dUancHiDNVJGwmBEUzRr9jd+AMZ5
rZWNOMkubQA3ltRyGXxNADx+XIZ1DyO4SoXA8siCWDjZ1Ngvee5j0HQveFdC9ov6
iX58Xx0+yG1kxvLivtYa+mS/5AYsgI0QcbpQMMwYlNLKj+jWG3AwNUAnPtt/VqT9
sq80RFmOLDgeZrDdz7o9MWDV7SfSCW2Q6z7gIjJFTeqM9gp8sIIx+VZrMRPR7oQm
m4524vLO/pIoF8GaKAlSGEv2rdu9p9ib2ECnzLD+aZAyd3v7pwjyJ7FoJtPKdt1x
AZWHhOYq5tsKDfGAArp849Yjgsff8bE3bfNJrpzjzZAw8SRcnpwtNQiI2k+8MUrN
NlLNfLxzfRz5hGKIsAj3nyeS5XZDXE7sXX2H9Pi6TuyNZa6OW3zV39Efxq8SRius
NdOxTZMxUID3UnHJsCKsON1CcenNk6oeysi5r3KGhLmYg2mZu5AcfagyLefhTC8P
SruimbTbMGFBTBXpnzGqTXg9HI/oxNgDFvnfg1GSU66Bh9/dvvqv7CoOSvKCYaXe
xmas3Erp7K0dVlQJzXcaqcJF1Xuc9rzPEq9lSVRdUU87sbsZww4fJoTxDB/q4X6N
CzR0lplLQOSHdl6J1piryl5TCaQX0F8iWxt4PgDGQwtc9YLFWMfewJ1RxUI8f7KD
HsprHyjPtm0XTJMC0NGrVBI7aqmiNLaRjNnKFy/4dVOl36mmmqBl8Db+pUrPg24r
co8+KfKT/L4SYJIuYL5oSW9uN0wIg8fMjXzEARzJ012FxIUvZVMHBFPasLaJKzKd
ehI9CPfEeh07HqSRJ2yUCzTOzd1QgOLupUMoUyNPsmc8K5z7EB2daHHxil4kKSBh
JxjMfFo3jh7ydvJGIkmz745IAjoFwhAuyFSSGrJfH3DlP8kXbYn5RdmUatYweNIU
VLtxOJooATT5dU4ERHS8rQPosJo2soPp7yV+yjd6UsejRXTvp9Iq+F2fMPLP8QUm
Kbx0JkYx2+oPEnXCbZzMYYZQzZPlij+Ok71vE1UfUR9TB5lP4jBooMpdyD+EetGi
2JxF7gXega71bu26sxIy3z6r9fD1JLSHa5mTJ2UF8uSqdh2ubD/QmHQG3SpPYWbV
DAaLz+g3FHbIIkOTXxmpK0736noepj4p50mChz8dR9nyry1RfFEJyVPvdGHVMFzz
wDn1FuI4mTE1wYHdwQo2lQpFINIA2sxzFdghEnFicAarI9B1MR5AzFxZqQWW17b9
oCdNp4AvOufgx8ljIIDpd2L4A+dkxcLv2p0jm1ZqNOpa2DSDE1GR40UB5s1dFK8q
4EemAemn7uUs9DGVLxGC8InPVJQpaDwqijpe35axS78d3iLzOpSbodHsprHVHXJ9
/yzkzYHqSH9SmJIpWvJvfjIxvplNBZJ/HHBxyKmeOybaq0U6EyyGShL3KlN7RCCA
ag53A7jS1URDKDTmzsUdDMAFM2dsYHYHnK+GIKJzVUp0Odx4ofEfmwfab0U08E0u
VakkZ5ihalbCxggPLHpSA1dk6SggByaOAGrVrj/fGd8cZU9b7yPGQRkDiIy0CaOF
lKY3qhjLS4L42aDr4hg1JhHrgejSBOf2Woo2mAWYfEDK63x+ZGMi9SKT8huBVoC8
pM3eab+xWYjRaUMnZplPiGjj1sIJxEkHVEOtdafJuy7RknkSEN7IW8vd8iCcAJtf
Yy/4DggfNZuCSvaAKdhxLtHcVFCl1NPao3II6opDWpoYZ87GdubEdViX6dqpuQQW
MLTG+JOZSD4Q2XIJOIAiIYPao3SppVsp9HmfK8XclxvV+sszOkmRErGf06IhK5Hh
+Mb706YyvHm0sDp5gqlCIuINLBw6wZId+NvYSq5VTLj9DSwg182TyI0z4udsJasQ
AJ0DqNnlxDJTFHC38P3UWVvsIEYnp1y+8vEasosa1JI+o5uSzVXVwsfj9jIrKJ6Y
HriBdQIcLWrJtDlbFf/qozB4G+H4MCqGS7lBCqjfZWpGcZuqxd5yR4pVuPumSSpE
iNBopuzFJiJp4stJJITkDCjlKliB+Sh7nyid/mrJKh1kJhOF6f6TyD2WXaoikLds
QqrhWrC8a9FjLdFEtvJ2sd1G2qPiHgEW0KCJv+1mXTMEl37ZwPkfnc1PdhvYoBP3
cd9XWUvZe6d2a+TdptRPjUwcLXMo6VWKbZtD1rD/bNInB8mHt/TkZ9bJm4LbCqjt
TAWcF1rxf5hRPXnnR0lLEq6er9p+7+cQ9Nus7NdPzBIAM1xszRodiRq6EOqjBaLA
jA/mDiHeOhqFfcvLQyDCAMY1dnQCfN3NvP0C+keY3HCJa7b/o0T9ZunyuCIk+jYc
cLyGEmi8h0eXbldjsvaQdzfrRtWIqNMIDCxemMBgCKewfcIgZ/CtfTHxa4qdOcOW
aSE4Q6VcGwmWMVeLlaRZKtVwCYmfwc/WKMy/dNwtCMc1wkW4kAIPq3EPoWZkFXJY
vTxL7/4W/8JDaG5M+D5RhVqVuyk4RM25qCqoVgfOfrmDpncSvkvzXNj7pxgvWebg
Z9ogqUsIo6pQrqatQGDgSvdicJaOd6YdQ9R2j7NV0go6ZY3l049BzMdQ3tYmZD0y
+G5NpxFCX8GWpQpMX4aEgxii1VLCKOiKlXa15TQ9+T3nW7crjG5ZQ9eET8jyhDLM
Q7E7x3LvAIsQX2eCQch7TFIoKLG3Y6z+AOsyIL/Nz4pT8D4hVLAI5ANBek2NiFOX
LJ0SAXHS1qqdKtiNdBtnAXtR3SbE9ACSK/lT1q/iaZeJ7zNgXtvhUx4JtdQjva9/
HVfAb1domh/jn3y/GbEPo27yla2Y+uSbfmdQMRjtTQUD42y2IvQCRHIy5+hzErgA
/MjyHy/9QzKQYckmYH2RtzrKWdD4Ug6gJzxnkoI/OuXLgRcGZP5H+x7nAvv/oBu2
moAS73Pj6YdK4CbfPTq/OuNndAJGPembn0F7X/yyZU4UJBZNMLteHAfzavq242iY
nepnN6GDJRYll1IKkeUQTNGc5EowyD3V9NQBP3Jp/e7FWyAJtYAVabn50jChEnBP
4AEVhxI0kNkWgbMofwwjlK/QQvaqoIeb4rD5DyEyF/NVNYMi2ncch23RijJ0grrN
eBK3SUSYisy42uPWIInGLM4oZdz07UesUmETiqMmTw+hzCxQ9gujCNIM3XyyQGNj
xS9eVopIMRT8wdd9A6qvJvk7y70fqJsBS2YRBKVg3aIdsbSu/Odmh2MmNbNmPoT5
2wCp2iaC3+L+frSaUf5S5Mhbvqc1ombx34pxH3Pn4Hb6X5FuhIaBXZm1C3/tFSDQ
2+QdpNON6TzmJ+75xb2K7YknTwbhvWZn+1e9nnhXjHS+Fikx1fVXtP3IAWWZ9mee
wA8eJh/G7hXUAnoY/7USm7YeIiXbXOpaxNxLDNI1vU0O4UlxWNYOLYK9IvGmOJt6
r2tgDuKJ4MVK8VYJrnwSu/n2Nz2JA/vB/KeTWREBKAwDkpNZfM8WkK2+VKRmmHU5
kdmJR4EIGksAH+jQxJjMLxU4fYt2R2qdtwM620WD66CKbdqX804xir8Eqzi4uFJ5
pL9a7UKQYeC4vyniGKIltBitKEglpRyHAUubkqeZiNmwUlwbZduzC1nRza6OqXn1
rq4zKVsFQ8OxsX/vrclSqEHLWWkUseRm5Zm+BC6VuNtZaPML9xCSB11A45fINBiN
d8zVAwwe9tnPMfpAP+C4u/4WJ3p7NtSpU1D/+NgDpBhedtgjXiKouuQTIy6nGGl4
rOAnEP0DLISyAuKL8gz0Qr3mkNYt8llEGtAeJyrWOLfr4Q1fKHxN6/ShVMwuIKeZ
TMP3B8rXzkaeISvEOXQEvqTPOetswyrCY1lX3nLpTBzWUr/VlD7m79J9OvG5XPry
BUDZVdNfHIWNeDN+f7vsTVATlWUVHas10I2Wt8T50uFVc9a9b/HUNr1zaoc9n8yr
z7DCo0M8Ma4YDdOclTMu8B65V4jlMxaMhlj0zTswO4rGUZGYGpoM2H8FrOoS59Xp
7tvq/G8StyhHg9YhP+TZ+Dl/ZLdPZaFHq4x26urdb42t/TGgcQStQmEQL4SOVw5s
xrgqJQJNjOaNJqR65vHcj+IPktm5Bd6nZMVWHogMNFo1X9TrVNrh7JyxeVKGaNBB
+1OaMWFJumIFN3rtyno9ptQjnamJOu1LPQl9bNM4ngkYXnZRJmvh3uEV48/9uEv8
/lzhblMZbdY1SdLT+R5LcoqTZr7HRAH82eqAFJdyPFxPNPgfGaB6+ycDCIdXf+94
MH0C/4CYxhPUeGpyvjEgSFMB/UpHsDHLiNTPFOt9Ht6wp3KOeGTU6oLM4xLjWCEH
vFtafehm/TfY52mpNCwJoBpdmWGCfcNE/RfcQY77UIa/nsBZRalYpt98mFR+6mE7
/rdxZO6jBQHNf3PKRVRKHUVZFe7WfAveeI/Jm5Gvel+usN7tUJaJP4+TECjoJVA6
Zhi0inHsl0hRL5wVf+tEFuGHBRlxhxLqKXxOhilNjyRB95u5ow2eZVkeRboSjo6C
7Q7TzVNc1DbxzU5Z/jX8lHtLPijClEJYu9H4Fs19edjXa3xrvQkR4YRwu21n8e6e
VrgJudC04rH5Uq8uwisgXwZf1uUELg/lfxPCQibETRyA7VmQm3tjW2oz5z9cbL2D
YiQ+iO8MfSzhw+NWJxcPH7x3WJzUXfiLgFYSlki0xfdhexCfTOW5bDIMed7jhFvW
xz5sgTUfsJSUE1CIpPKuS3DmK9CwaaarhD3H5b+vzUmQvvhk4g6ZLPbXufwVyYDH
4bRSVrW9uMDpfGhEy5khyHLG0+HjBu7a8AaommT0HvnHnw4IwSqZfwUeX4aqNbrN
umZ2XtRVIjfIj80LVSnCjII2S7JrLKxgYp9qkZYT5FFxxUD2ZJFwP6dVpgrQ56hL
BZzJLFVAep1C7nnvYu0F6ovlUP13VClvBxHGk94yt/HrSZkFA8iGmu778JcTmJ/Q
NNa9UAKtWnMfa45/oFSi9kox2HFH2AenSw5AtJy0tiWByhxNizy9Vx4E/0wXnSRw
8lVk2we2xTXirT/p/YKAlel3d2/ucNvqRvE0CEqoNTo8Pu447tFeVc+QoX8lYhHv
7w5zlqO6j1nk54AKu5g22kQgbnaZWamk+0jJdRWcdfZuT6Im/fP98KHHIZLnBdRE
REyzLKX7IVgP9BbybjDzYIqH1ampOJuwtiubJtEDtO8BrHQe1uCPKHBVCXAl3rsB
v/rbWg0WOChx8q18LxIvhRb7HMoWN7EF4D38e9QU+/sbqrQC52yXjJYJTjTSFN6n
w/BQBC4F9T5b96r0E0OAV5/9HpEk5qFntMxq+IVoYypij71Gnb56fHXYmalI7ro8
Va8P5TnEbvgOd/eO8cif9jRyv56pe6pIZ0Yk84rh6iXTVPsidhCfpcZd3iLf1BcU
9IMaXARCRBpJCEsYyMAcozJr7dnRek3UDH1/x2RyLZTjmkvLoIEmRcv0MU8F1ZpJ
DMML0gbXcgO6WIdES2zedSEyE5iHBED2ehXnd74WoNl4nn/1VOmgFWTyCdxNBHwR
r9XofzygzNYj5o36JXJx8z/oNxAOFhQSAi6j7pqPnmWFH03mASd5Ytlrfg0Pjf5A
EFvxovV60mRYuqsPVQaR+TmsRpD3BzQLu6K1M5YTF4ePxKemFnDkEm2vPNYzUD9t
RyfA2aQH7hWh8nBMq25/BVCS0kFUdNhvYW1DBEK4VEaszsn+ybxkMQKNgTS+194Z
FTHSCKD5uR0MJ3MnL7gZeV7MEGq5J7LP3IPu+A7jp8MgoFb4Q9107/Xv5eCHdsSQ
NHqzv1rmhKK+3X3+i0lyf1UPvZvcRMl5gjXdlsY91SXPd6DEHiZ1lLiXtXgtTibi
rRr1r6/iv2gjgfTWSAGmzOcXQ9NOpPlLRGBZP6NEOBifWLB/H9Z7kuP6cdtboULc
HoSDkGl7n5/v9DIBME7xACdSWmFcpGhQWmxjBxpDbUu9m+7ijxvjJnKfmciupDSR
QPoMjdUUR1oNUVU7+id9Ia1LW/QVcOHwerEiUcq7QXcQ2DQbyfn2WCLsMCNVdZy1
gEwJHEGKgg+T/CVLE4QKilCpHbNTDWH9aQFLM7liMf6+S6kbkm6LO1Y9WRMN6z9A
cFG82TGZ5aWEjHZ1nI71ivCF3UXdIrlKgpOeTwnxQUyBCzZnxW6SOpnAaodbofTg
aqzBpVs3qSA9niiw8KlByztp81BqmFZ4jSpFZoA2ap+HLjWpN2/HGal4VT91R87t
QaXmgUlXr/Hqm0OVd//1IZFeXsFjKduYGetprxH2Mhk/OKbwRVNu/bGY/56LCLZF
sTuSb+Jm7+k23p9iYvu1CPpvpl8MBYxiezEx4SCHjZgC2UYN7xODfu3f2yJXhP4T
7PJx8yAHG1qktKp7xUreXNO0Dqp9IN9D17OKli+C0xH/YfHukCiULmrFdzbmfUfY
v1+lIX/OzDaipJNz17vVoLbckw3ym3pVX4m1Ttb+wFCpcHOMw0+7IsaEjsjWr7z5
5qoOi8vaadxkrsNC7qWEnJb6mL3xxYfK0e00N3XD7dS3cgKfzg5t4+mz9tRhMawq
dyzCegQsZDWaB4KVIdg5OOOY9iGHwz+U3SyrG/++CVE+PZXCwi/pe3KROQ+pWOtb
CMgojCCgiN7aZBEUaKwdyURf3Ies9iwRAs3GbBuKsWi7SgHqScLjw9v304I1F3Yv
qmrV9BcF/c9mm2NCVVL73C9gz1pCCWtlwB1R8a/zHiUueOuQM0V0/24RrOamBE/A
g9IviSfbgUJ+Gau7R6Fg6TRmcheG/j+lMhXYEYEZ9gwK+vv38EmgNXCxbxglLWXd
ew5KnrW5VxEmxCJVr8oM3Tz/DFe0xsu+ewkQxnxmPhAa0o6noZtOjMaD4op084im
HNjDAPhjwO/U0HHjEltG9ylD9Achz7bmsMibNkdGSDqLnaMjqK9JyFGpA3suz46Y
AbIozKQ2rDsm/Q2ABgqQX5OkW1TrV3WMQZj+xUmTVa2ddvjHVU/qBEkRxbuqREOV
6Z0xo5su91yLXNxUeUIrh1Dc3L8j8Kb75qtdcIBpVzPrOqjWd5CTuC9EXM0fo5p/
zOlsTH3Q2UDbZfPmdQzJ7zhSvPHBXWEMNwj94EmUCUTYdiZX5vlM/cF1mGa4++DI
M/D+H4LxUQ7A6dheDATW6z46Im7Ay2hv6VxETuhVk1Qx+z0ANXr09IzsvT8qajhx
wxhJWtvPQTrZx5gDHelpVOr8g9AaSks8cvbuuREDDWVUdh4c8kOssxEDucM76U9T
tfMJVT9dxJ+zR8+WGgN2r9gcpuYDNVm1LTM57lhwoMXAov4oQN3l5Flrfnnayn8p
ntPzjMXnCR3B1DSKL9aIPz81oLGtxENMPkmDIBwzX9Ab02EiNDDQNVt7CFJ4JRVp
YMMOPlak/bpVkCXvivDo3cjqo3eUByN4aOw/3NF/lSsODKOUJAU1ECA9NLtwnkH9
Uu+pzGabqa0lyYAevn0Pgejkgwt1mYvO09LIOp/697PTEKiEsaSHTA8j/t9b2Mq+
ToslMeMNRvJoJDtJhndBp2q09W4i31OXu1zvsYqzaFG4VBWXE9XxgWwl6V5OAYyO
r5qYuY7eWwBL/e5v0zdk4+5uUZUU5iBENmGgQaNEhc3VqPuKyxUNgCN7+P4nyc6F
kdC4/Q6RD7IUj3jkQPUfU2wLhid/7sQMm0qc6Mo4kVocBhXzAS9wZ7uiGnRV0ubo
DFWLR+LGzkeCh6aJyiw+xt4bRW7SqPFYZEPZSN4nOWVkkMdub3ebVba9xwgxuctN
/Fl+VePGqq308GC+TFWUbuV5tDFNKTeG5Fn7FXdsGLJ/LMURlg4LJ484kVA66a5S
rLBKkr+p3JANlBWQyPRBMu6EQbDu/M4cmC09i6d+3RRGFW7AP1fkP1ghO0arcm6w
ZW/55mA0YNKscdTOaFpNHxq+Z6Wqh6JagXViLKJKBFwXjqKj4neYkaLePhxIREBS
cWXdxlo77r2mTqWo5B5fBgh7PC78Fy3GX9CN16A9xtYhVF73N5EVr6G5HBUDkQHE
Ex9pZAlCT4982I5Tfmh237zV4qIXW0xeM2lc9xvA1H4NnBlNYiLsXlwV5Ba1hMCu
kI0ZYBB3xIOWbpkAWKLIQ7LIr5c0hxf0onLWpp3HY3dMOdNn51J83bFfYJr0jHL2
l4a9m9cDXRRgfhYPQRDwLiXwxVHqVHKcNgtjXdAxCJrjmxDR0nqsMBRTdCrmU2I8
q98itiTtujOVZ+unFVAuYuB/JsL3zVh3stxoCk1DGqbb8lWn1rDUfA9ufUOmKhrc
d/mdXqqLjcIjvMWKJ155e+s/YpwO1LE9eyaWdZnuxnFPuS7RPenJQ4nUvnerHjxI
mg208a1UTD2XWt7WptzrC6Byz5sEw6N7H978mxFUcXCpxXEBI84UWnEDudRgOO/g
5TbEL8XohM7SCsWUcx25ccq3L9rpO0pH9K/VqGRZ8mEVyZR/P8EU98xsD77BIaaQ
BqVUjk47IashpSI1nnp3RBowwAMoB5iXphZBlXGBk2LlDN+0wy924o19i4z4Jm6E
eIhkpMnCyvaD5u3BvFIPNfi3Ntxha3tnPJ4EQQxH7Km7/OdZEehNZXJ6fPnsomzN
vbDXCKFicFYc11Cgo4uWaVzK0u+ji8x1Cw9YiWwW2ujPx/gxr8YvnCHJ8exnWxe3
8Vsms7cpy2bzMUkonlVvpd6jnivKogn0TQMpWOzlQl5cjTQn49FHrI6xiEKtMwme
kb0yFQvI7lW88SB+yP//dagdVMgG6QrXrOAvTrDZknQI9T89Vn3yhfaEVxZa74oW
d3Yah/7j1Pf05kdV2rP80ClA+Z4nXW5bAA9zo/w7fo+twxJhzkdriOMn4GMhEReF
UceJ+J88UXtqWOKFUV5oVVJUz6Y4ivgVaTZT6d7RTcl011A2CJokvujh3wcRUtUQ
bYt16S+w1GULyYDeAklwknwZUjZEXfEwRiRkdME0IeOfsJofigb75iB4hGB5NaSp
ibmHus6qKPIcB1LfA27K0sSFVGov5TiIwbCqzmuei01ebsa8G2VAuNgVrmlrasjY
s/YWUCAiTs/d1WT29KJRaeUtvqGc/+ZSXTfwkBT2pbtT/NnODOE3Jonc3DvraAjL
FQLrKAOiAANP+fv57R4OcVqy5FfQwwL+1JNjg0O/IHCkrluVGRGShfygiaIPxVEZ
7Wa87nsfyZZITFqZhDF16wNGop0SSYl2h8DDGuPTaTGWG9u5PseNvkkdd7j5woim
riiZOB8a04G5u30z0FnrkbWKJRu5c6J+zQIXwqTBUgA6QQ3SMrpQlgeBx0SLxLNN
jec2dzKMvJ0XfaxsFEzgfPffc2ghFNDdaCp4ymbyfS37I+P6i+jHd76Xswh7Hif1
h0qHifyQPBSexYA5JebM2BCQ5PBx2fuEQ8FGxWkaWDLkXWZUAgUpiOEi/mrsDxgz
AusXfA8crqqu8fRrtdLKu2Hk2OVKhRvPAQq3lptwSfIH9sJz8SecYV+GwiOy1VGz
a/veSjnuB9OC6Sr7TohQPxsmgC3XSamGSZ6Cu87osZF21Q3DV0t+b9rP9Jk7jyEF
NVxq3hYDn+oqNJHfDrLDleJHZeH+wS0tHUWNg0CZ4Bo1MBZh3TBV0qCm3V36T0Cs
dWoJRickwHmuMs5aZDZFuGEs/M30hflsUpN27o8aHFOBTcSXl9vcY0Ty6DzXwGym
kA+NNQNyrJxhnnyV7uyLWnuHdw0VdT8Vzq0Hj0sdRJ7hYMRLMcMVLWccM56YEtzC
CJ6nJyzTucS0r589/f2RpkWKtB3cB4v9b8wc+MaWDbLTpvp8uJNF/6C/St/i2KG6
1sRakYRvODTpTLl3LFd2ggffXMUPBK87AFJVyGZT13yhV4rqyFwM2YJUVKrca8F5
R3QlJvXh2mZs9vO8aA6EXINY3jKk062IF1wwowi3xDnsvLvwAO41jm7d164ICIpQ
hrJxoo8ueS9AYHz9Fjd/39h65QnMqyY/9UkHWXOwhu+fl4hKj0B6mPBm+Q5SjZ2L
kL7JGzc7YfoRwihYPlmUP7wwdzXe2mCIVrJnMH0kNPmwoTy4wKkMWm42nZ49Y/pp
//IEy4yzw5XUEcY0zLSCSQjcgQkwrNN77W7s7rKnlZ4TrfmwzjFkY82vU0A9cPWN
TrCeMJgZSHaYnBJ0qx0xSjP4fT5DYnf43e52vPeWaTyS891aOiClmzbmveTmGgtH
9BM3lqA9L9QJR+XKLSEsrj5/Lno14q5W5l4bXfIz1VI8pNuwDzPHM75pUSkf70wF
98Ap9phpOZXb0UKe8IgYobaUHxL54nitPnQy1kwX6ML8v2uHIxGYbgQUIDP+hgOr
WoKsBKI7093Xq6aTID55JMbqCi2cHFd/BthN09/9Nv0NDHICe185p0MdheqJzS0f
8jdPMukjaEgKwn6D4/etTNIfClJqG59hZl6RELPZnKEDWUBLMRNZ9pRP6J620Sm2
aP+7yHGPc45BvFsQAnJ+Jr0diQMTSJXaTbidiCVVVhRB3S1poNtSGM9qmZnO6xry
f7sI9cNzi5wXKW4xvs/bpvzt+5ojMjzlZyC9rmvz8wpNkUjjD7iYI30xC5kwTYUi
xRSIR/dhQLmMJY+R9ui0wkkPIC2qCum4w85oCgsxzCb8sAVPho/aFQ6tuOGAkyW/
UwUR+pTZ8HqhUuTAFTSB/k26oO5xqTR7Ujl4neQYYqJSgn7Vk9F91vHagyQo6APE
h0SkeTUGnxYYw9/tnUeMsfrKltW6+nBFj2JlbOT+DUN+cjNKWxtXVLmbadz+qUQD
7ITVwp+RFWyIgLyQDj8odIAf191P9G/mGnu4o0yC0LYf2+H6rUjcs5EYHzsjoogA
J0bfAt3Brz15S6vuealXzKjwQ4kJ3hgXjTOE+wuwdyXxdN00rU11esTSCaxAoapS
UaM7f7dKbN0oVHFSxVEPoZ59RYwrWcmrGW3NvIGiVeUuoyZEcp0KOb/P7pAdn/sE
frucDLL1cBDfJv0Wt5fCkVVBS0OVvkE+vsSLji0DfxOyIvsRx12K/ljHpWcNgwFM
lCEeJeNigWc6+se5fTk78nnbWMLsveNggNe+rQh5uTnSFHRrXWmVfrvaFHpMEMAc
9pLimqlt3bd9VCycK5UyOqm77UlSOms/dH0EjFJYxhbWcN2fIHy5uZ/fROkBO7x+
32dq4Fk4ajkEthrRPmLao8Ws7o3IAHVCpNt+bktIDDPpFjWWslFcroraOw+hF7NJ
oeh73cDI2ZkK/dadAmfdjgRdLJh1Sin3/Y2BJcaFNNt4ZUik6vsOO5egt8/EJEp4
VcSgOTwe+ACjHd+/R+oCiaHl/dAiWTUq5tw4e0hm1yRu7ludfzblDCpqlHP3lTR5
ClbsfkzbrTPDCFFx+0jeRANiGXPJpSn0Sbt6gfJAdSO/NWqmVtM+HFRrAcmMoUEX
FowmwyCdDap25plPAXybwAj09padpUt934A34tQ4ePip2H35+CT7vnd1Ch06uQrL
TnPLR9MJhOX8LwcgN9i/6S1e6yeTsiMBHeLeeUAm+N4eN5GQhNxY9OIh9Ia4w7qs
yH7py2/qT417nrSCKYMvnwjF3pkDX4DAx7L7RuCaSaiPpQoMpYZQbcdGJz+QKrYN
70m3OOs6OkFDnljjYgbyn6Hh+R5W8vbX9//dLtRinHE/p6rRf3tP8y2UvvjxNxiv
hwGn9eTHMb5JD7jmktHMezWhbwH83mNUJCvIMru5uYVpD5fT2c6ZeuVD70+0n1w5
pzcwCq491S3X7Mr4G1DWcc8RXwkm4vFYTgelY1ufCVGGvOhsnFFUlmV+VVGP1I1v
qLV96UFIQaLgR+PmnaP2O5IzQSNuGNeZUm/pJzzLWGVC/RDAI0n6+pgpow3x2pIc
nm0crz7U4/eNjIL/wNp+J5fK329IcVRZrjVDkUgwaKFTlc8zM+Juxa4k7ws0fpdI
TdQcDQQxnP2qcqJ5KwROqVTqSyjt6bpsjvPAXBkemLwIVYjJnxWDJwWbLyAhc2cl
LMAgDu1NHyoZlOS+naFu59BAUyDd3WratEz0CWcDpU5ASyaD+r5yOUUFDTWtSPzb
dOO89jyE8qoCrf053vPBRy6jMlYAzgWu4dgLOYMyRC0TAQrduOPvWYqQREuYSI9g
B9AoCUF1zLvP6PITkBngc44PlJLm93VyHRD8yLblVlSG/EsmGWK4RtA0qLF3ow5T
xLqqfbuJ0TyCG7Vgh1o0VA0t/8r5371QvrBjDj22bdvhj3rBzXTA0laQgk8/Su+K
XzF4+wD01tewX/iLKUaCMCreaV2sKdjAfdVFf1dnsI7XdwGLLdPZgKXxLkrjFE1q
ylahGWV1O1jHF6L0CExs862N4eS3zAaGg7ZDLVYVwuYbOgpJWk6BWkvDz1YQ9323
+p3rDEjObI8JlA5HjVDcv8bOyh+yrMSXEIaMDfEf0fFAVX4an1vd0aE6NE8EtP47
qFoQwVRWbSdxdDsSRsrsx44CIBd7NuCKHjAWxz3rCQ3Or0FjOM8o2wcKU7vlHtW3
yyw2nvsSdZgxpRtvJne+7vr91vRWbK5WjeRQhfgSvYIZ3Dq8VgVZF3Vi6F+Mk1jV
gE57qG/z3sIdmlA4Yz78GQnUQTiVbd+ZzB1TDE4NU9qRDAp0bKMJtaC9zElSH7n1
mIU/CzuHT5TqgwAFcDmQlIdC2oZoqefZ9XPKu0oYEpv8qfntlxXnUWIJ7Kcyrsq/
R6UlpUoCEYXbkOWOY/PACcban/rzPkQ9bGY6FYIMmDkRGuhcwXEixOR/jjZRRQtU
Vz4buR2h5B6iFC1FyvRlWtBPvqdCbNoaKD+FbyX+G+h7zkkYab6LEqtxb++CoGkA
HjUOJoX4fSsLvE4iYZEPUb6v0ddc37U/lQ2SJuUP3OcJb2UhAP/tmApyW0PC/qgP
/LpLGUtEoT+Hh3Lb9VWgbo0gaT1p9Q5byZUFFF3KjcIZ7CUk0b9+0sXfz777iE3y
cVkrHgLpU0LyncSwWsvnd7kj/YsmttuwikLOFdo5UuxRmu/1WjBmrKI2GBqJD4oe
Q27rhdrNG8bjbb++WycapgH7kzl1WZCwI/jlvNXHNFdcxpBSAI7M9jcvSEFzrt+t
jFieGxpzbk7jsUKNoMeXhnMh38dqyzTAwZ6fCySklw5YodpHP35k/NpoqdVLFR7n
5evjh7k10Olf1NnDIbB71lbjU7LRRJCtNl5WCPthn6Eph6dVSQTv0ySBh3y39FZY
V24m4t4wwEkEtFTcybTjlZW46YIz8I+Xw6TIk9Ce5dFP04XD/HqtbcBdZyDzsOi9
S0puDLC3nQWWHkL8gjk8Txwro3X5F8ZQ61zOSgLvxPUXnFG7yxNdW7n9nkWXEOk6
NTlFyS0l+8oDX7L4qrAcXj7cIRe2JH0jvftdHN8lQTnif8VYKbQk2o8xU3koV98V
B8aCyxo2dYtocGW3sRAD+x5z64MSF/9FWcVHAkfLmOcORznnAbElECbPg5ttVmu9
KGmO1XuX1WStJdoRfa+7AqbG9qzR9MW01eU7jSnk5hoJawtW6oVrecGdrGL6uRDZ
DevvETartwgIN5Cuf/Ns3x4lggrqfJ/B+vvDqF/fS9xvVxsnK4a23WY+BL/aNFvR
fHn2VdfgV8rtEfLIfq8pzX8ewuFxfBGPlduc+lKjrjFFGOydHXgOV3B2IMW1/zpb
HC7RBMRGyyHVTewJenp8+3Z3Ge6AVbTraUGudawTnBcPnvgSeq5aoPiOyq/xbNtH
rxxR8rUhkI0b+AeaqZOBHYS8X2xqjisAeic7DYVUDgTBhLZiKp+0Vko/OpFsonjA
G/y7e7UysY0q4/afMwjgJ+TMFU0GeeRQl0Fu1W8847Rf3ysbOKTvuCSKbPmEJt63
T0bFVuUC2tTZZnXaYuZCaGZRHcWHKyT7oot0Tpufd696hYlbFIIkigbNxiltTnXq
QeU/PmtG10lw2LsmAPMMcUVcGkP2VhO6waULrswZotTZ7XmbLhA1gEziJeTK8pCI
Syk1/smWMQUej+DFXs795fPXVNA8YbozAIoC5EyiPT98Od5grzNdptYTx8HoGOeC
f39LptVa0GtQbzYEzNfPf0AAVUoccb2htyyr2nGW3gntprjiIHRTMhZ5U08wbJ+V
4+GML8+Z2IvcYgevASRrAlk9C8hwasdOmUi7DPU6kdsyGyi7X7qm8N4RYVi4IRaE
cGHnu5Wf9G8OPgWTiz7jn3IBe3hsgrjwMm6IAAQ7azADo5cl+7uUK2rUVRz+6lr+
sH761WIFwQSuGRY7WGtSibayN+nX3/VyDW+bhL5Ccw6MAXc+uWvHEGX/4sHnY1lQ
NbXa73amNhjqyoNnnI3hI7rYXSDeXLugb6PHqKv9B6OkIRfn/nUs8bJJ1sClsOht
iWmFzRtgdJl/A/fWXDOZz4MIFV47Nn3i7R+ZYHRCMJcVP9lf/KxaSRPeLOO1nGVZ
8nlr6IydgQ5TgH1ygxKu1C03xCYzAsVa2m9BmNQt8uqQmOlrqw8IMrWs2hH/4QsU
b0dknezTDcrVIw7OedI+kTq4V49dgb7ks34CDRdgKF6ZWhhTxC6JySLXwaOqGLrK
r9rRDxKsLjvV8kf8K2WQaP6LdoRndmmjNvB02AOBvTYOYSht7EVPnSMU1EGgl952
8xrq7GZqDJ/n458mN8sYUcqOxZpRGcg8f8e/81L0Bb0rGIfeCIk+83iPQjQti5oG
wQ+XGX01n/I/dQsP6J/UqHylvNzMiSW3Xy5DOcoVi1qcK7BBKjA0DaKKK8fUzyai
DxySVMMX9xZRUFF8a+HOwZ6nxCfH9Rw0No6/QiLG+EYUvECkuAnEAh0YyrJc+UWH
JDGHAmo1VFARUu8prR5isZv+t3K/LDxGCKowLd08gDhMxowsUUcRYIfCHgrvDLxL
3f4Bl/k+0djcMbrWg3aEp35MtSJP45CpHTONAGf+KooPNGjTx+N2gRD1uAUk4VLu
cXoQrBifIm3O6t3z0jKnsvUQuymRzU0Hl+b0dPj0Ze1gFyyLU7yitk72ptzmwt6i
GBILYKPsvPNtYoG7wIRgRorUOETryRXsxUAjIZavIs2qmPEsMmPUM/YzDxN8t742
MzrXokZQeYCtvkWtG2PGD5dfYkgQcYsOgJOtkR+bBRzJqFdRwCo0R0E9p/XU8jFR
COhl7knRFzQT87TDRx1AD8xqCsn69evS9sEtWC0wUJ3rjkcc9Jz5MfMSIJF5t13v
cTSbwmOG5xu31ExJBtrzTxSEhkZVFwYNygqbtHpOiYmWWac4/XA0Ab0mH1rFk9N7
Owbl3BxQuBdTXtRU2RpnAn6xSVJwkNHzwiD20o9PejBi1VVHlJHJqqKfrT0whxqX
FtSlnaBRZkDk/8Roazm5nYvIqTUJ0Bw37Sh/IKJKj/FP+0IGsJbOvDk62hkdqzcw
4n/dJKESpeAKMcnkQ2NUAlTvPMQfT7+Ignx2Iyp82d+M/cIwOKLfYeFqsXUjTa5B
7rhJbor2uSkHhTGgFrtiYsl5kHjaXRGSjHlTE1TPl2XQeUQYlc/L6sIZEHFc+B++
I/tWmqfEOH5qZO1X0LrscpO1bllCpJXGv/r2bM293S5pajz8DKHFGUjTbGaPp0cU
UbJ9Sa25JswAdMPBTLJs0XuVBPUjlPjL46yv91OfInL7CNGGy31g956JKvGQliQT
2xj1Rq/OFX+hNpJJYex1TMpMZ4AZR4POUzJuRlyHJMho6V/74JyIff7UENpjrB1M
yw4yZdEUq7lo/dVw2+zbayo6qzLGKtemJpoai+MBmFjzRvZu+AfMPMqeVBATHwLU
+YJXF8idbw3RVcs2jAvOj1zKeiAz3VH2hvoLxkwExOgMM8Gr6LkNQCK6YOxHpvNs
ExXcTwevu8waPlDJeMudLmt3Sbbx7Ih3HF0GuI871KsTnx0Gm98Kcu8Z6HZmxrcj
WGb9oi+m0wNXVe0QmYTuXJaJ8pcOHEpTGl+bZSwCr5qhnHW8G1Bo/VlV4YRXrrca
L5z3Z1/Tkk9/zgPDsYANS7WtdHRc+ksHmJX++5nNh8d0unFemhiF5XcKZds4xg7+
JcH0DNLN5XDYsCCQYHxDl+Aow66rk8v3uMHhF/SEb+HeZ14Po13fz6m/aoit1XH3
mtKbWxhNlDxsXzMmerMAqQMHC3Zx71NieH/fbidYPsXjSZ2Sx/WqeKv4GvQdZKdY
WrN3x3HHjE+cgqL5a+IR1qAwhvum1l/hh7hEqL12nM+4G46O6qTePmp+CDJBvX20
PTQPdJl5YPvikpDxd4uCJijTa7/GenjOGkbLZoyTk9TQ/rtK34wjP7C9D0KA6Kb5
4YRYtL1sDghMu7NWyhmIp5ROzVjevvNyc/w7UoP3q4L5xvLHbw7N7ySVh7CfyA0L
BpxPRHse3Gpz5FnmdQppR6Yo094+hkQWudMV9FpXgHtFh0S854/d2viLU+kL8YTG
GaxAxIfxYU8Ni3qRxPiJdxjuWTa1kUeLmBFSeGNeIKJNBAE/Nw380fMV4l+/zYV8
afJ4DY0iR+jAfFPhL9HEjzEFB2vo4F7LaxX5HqebHMnxzH4/N5EMNaSsB7jDWcDS
Ac8itgnLgF3CuKHgVaddlIz+iP7Y9RkiXCA7Go4JCAyC9rXqUZJWEpX4owc+Kn2j
Oge0ZxjDIh1Wf/jiGiTG7xyXrdN1huq2POPKlyIkSpFxq5MOySZGjOGQa2OsjlLa
5L/96jc3M8ZID83ebuZraVvTpT/gF6yoKbu2YZZ9uOfA2n3nxRRD1K/KrxsZ6kuN
gYweedZK7GI+xzMha5r2k6H2UaaaI0p+24iJwln9edaGUVYOVViwyEOJDxCX/0XT
h5R5vu0ckA8dXzrWExpSouebeKr464lk4u/Vk7kJbwim7IM4E7MV6JyzSoTarpjT
rsKzxwOvXxh8j3Qkz9ZWsW0gYKIg3llU+AqYIv3m6LGEJb0txwUC9dvDVyx4tzKP
hBtPqIrFuKP1IAwWfRNZPsjUI5vU1Qeg18pSwm9ZFkKnJjvVOy0EWg7N8aoDtRHp
sdUTn81WkborICLcWO1DSDdZqvwR5GwHDnTBPwugKt7hbstz5d3Ms2t2uJLwZ28T
GbVxdZl3TicBLyglkz2iRKnYfs0Lpfp9RQbkSMfKGpaIFDGPASSzGTf+lrE9ACrd
zCcxZ/M47wEKoqKgNcH86UBx/b364m88oCkb6TzD+Bz6X8ZyGmvbhl7YvN+TkRol
MX8ywPklfxako8xPkNGa1Pt/XjgAvYqe2M3SRb9jcdQ4xJYybWKP+v7XPt8oIEae
YerH5dxKb6Zq7E1LgL9dH6SjerCRg/NOZtP8c9hjoUqiet1bP6iBb5/Da66MpZTs
WU/lWs0KoEZHiVtEmpebxrP9l+/qQjCLDIEcjhCC7svn8sTr1ZErUQag1zlht4oX
X1IodFrVWJV+WVYYLpQ3FSNea51n1YEBUSdl+HuHFP9Z3zB8GzZXuEDO1blMoaqP
ZmRp3Ot/aAJcSGhhDGEbBpfREV625xIYIwvCe1bhqXCtDTEPkm33EABf/uRk1hgG
6FVaxemrws/smgPVrjVeR31xZxz9UA47HQ222wKp53jf4Yvh/ZQlaytx/OaWMFwf
nfLIgcv4oq1iIjoFCCPVRM2gFxhrCQ5ULJvHfxEqb4XcObKUT/jJRWN6mgMGRJFS
zYNlarLGA+mHVplr5E9u/XqCDSl4OhbFr0Carj+ypUrFK1uKm0i4UsCw4yIa1Po6
yAnfxa8RxcIJ4NIGx9FDjLRRY6ygv+6KQ37JUXeiW5mpmBMzdT5VxzoKtMiSrvtU
MtmSf0H4RLRh9pf3wLZaiSLW2emSrEAgiKiQnzvR0sz4cGfcmzrpnZHHittc1U1s
QCKbrDveQNXAhT3v5LDikry5wCDKfMSTRAJaZe17aDKbb3RpU8uJrFNQMHRlcD3E
6llf/OqHOX1rF19Oq06tGgPkTvotMvDBVqETBMcOhK42lZkqClHM/4yAJFDfalyF
qYaj1Do19K/2TYlAbuEca1EB4ziJ9lGlhV+poR4xc7pZC43+GXxSv80MSi7Pxo9S
qO1P3wheZcmeHtoYAFv4FLdXcekdagF/LTgv4QKiYnKl3SOO66nZ4NNrvUGuzjmM
3A2Nwi7D4j8StmNTs7bLAoIDYOcqrA/0zN2kKRA1rF3KVDMLN8spIB+fOcMjDjlZ
h94MqkqeZtghxFlBPWIC1E87DcMd8NRgf09Rt5FrirnF19cmw/5uGAkeNczze+38
ONZPZdHlpHeNrK96a+agavvk6mIivYW1pbQ9xP7ZztSbvoHL1w5Fc3ps1DXuTeFf
MR9c/fJnGlF1pIcwIVuyqVin2gSXlAr/xxAKKXYJ4mtsadOkbivLv30GooyOd9Q5
bIRTMsqj74ywvwe1jBk05eYhLKs5rOVmNvpyFuGISRosUJsZHbBGOtcY2jusiut1
pl35OVz9GWT1dJR8zqoYrt4dENhHoIAaKecICWJgvvmcPoOyxFXHpxalZH8JFhUX
dqBtWTxy0DLw5Fdj8wB2Ipc4A066jKNJJPkYRu8poDqFKYbSZvpq3pBmjGPolPCd
E9wKK9vR5KMNrJlxeoVmvpi9z3kQGQEhOVf4L7fk/UQQ0m65npo0k72fQMZy68zx
OB3pscgyhEMOeMEVEXC3zG3oxz4ynVVtyQQ284sd/hK8c5QoGcHnRjXhNkbw14Fv
wXAlYJcGvey5JBVk1WeX61JVeze2bAs2WxqXOtaA480Vk5osTW6xAuQU9/0HCsaU
Rc/1sC2bvnDzQ8V6JF5X1nHGeXrgtG2uCiq7OXl227c/3EtGstwRz8oATRSINRLJ
0S4ldehcCinz8zJZRPWoYHpVUJXmzS3/+UuqNagMC2h8NIkv+Ecs1dJGC6YHlU8O
y7pa0dVoDipW7I8vtJ3wlagZfeit1WCF5qMHfVz3pqlQXfSV6OFGjWechf0HgVni
bNWYnD3RwgLoggEmqFZuW0443892eQxHkX9nAXy3D9akV3UlIuAtRF6f9jlVenFu
PW9BpWuaWVyHUzIgAYaniIoJM/7+XEDtTKI6yPxlMEaVuJ2NA5elGC1PTaW66PMU
YdpQUi3LbB9SzDp+914qYt2DormU+b2VENFJCG+IqN43GBogb8K4TjCpMNdQXqNp
7LTlOZJW1ZFIcTW2zapKpmu8ne52jIo1RuLhjCHM1MTkOIrGUd4QOgkmIrRG3AH6
Vswcaxl0QATTjVz9v5zLzgdWsg1yR5xjlRZnNbosqU0TUMQOljHXJEIrTqqIo+Nd
wa1Ia4AAiKOdjVN+TJCm+KjVz6Tt7Tmue9Zn7H07PYxNd7f4jBmlhtCeNlfXTB5E
XWlPt3HnfqcP0Goan3H7+eSUi8Kh5u2nFJ2tIdQ+N1HO9Yc5ZgkAjpwJ749VnAQl
Yp0+S3/cIzUq5B9ngmc9jVLBIiDoS7ZYm35Ae9mAeLG2nXz+4Da6z/a87vb9KHTX
PpHeUCy/3A6EDBoh1wt8iwwSkrH5ikzLCs03xPgRLkYUa5+w5iLQAAi8tdQAnoVc
2UOBZeiWDuh/+t3bp+abqXDYzvH5NxolpWQYr1b7151Kij/LD812LWm2dAAcgFOJ
q3UpfpJ4Dr4zf0Y6N21Yc3bJcGG0QmTF3jQWzc/zy3ykfo+Cp+oxv3HvXGttYyUI
nHpilMeCz/0PQQFj4HOI6blhrJ5yqe/AavPb3X6UtbuQ2P7bDpdRG4tasXk7e7T1
z7q/lCNrNL9Ovnnl1DUmTTEJgronR4UUz24WPZ4c9k5ibvHUB2ZUU6nworB9TEQ7
KrRthKep/D/HoWV0Iq3Ge2WVYGOzNXmgSQztRJap2j0Yr5mM/jiA5+5Gakxw9wtK
adTKkvKBJCsUU9GdjGGmFUADox7NRNc0pHcXXNPLu0F3PniZgGwgS3jg3NdUIH80
I1eCxlENrrua7omglkhKMAjnS0ijLd8uGpKgZeTUcH5WM5Ddy87KjQDU05apJNPb
Di5/8SCGpG+2YTEpw+MPjY7CF8qZtNa3GQpvSKN3JvzdtydZ19bH/z9HVH+Pmmux
yOJ5OjDGc37E54JlwWr+Y6QF1hVlfuOHgCwIpgx6smKeOgs5eRHyU3E3kgg1J6Ab
JBSoS7i9lUsTkh+i1+vroVGxjb+Ifn9f2Cbyy3NW4naDuGANSnrd8TfFdY/accFu
I3X8T2z5Fzxo3paR9vinUyM1bXroXiBqZ7QYUTgzDxhsRhgVhZOIKJZDEf/nmiZ0
Rb60LmiTiupUFDYlRRIHLd1iA46cPhArqPrVF0uRZxai2GnIxe4uAkLY2Ck6STzT
F58bvAEvXK+KsSWWqRMdm8btjVAzKisNpnUgO0MndT273cq9xputT0KXWGytI0tS
ZDAYLKxtQnvbHpMMb7ezDkNv2autT5jPfyLylhafWCd/NFzVDz/WWAaIH9CPifi/
amHMbkSA/YCH4jEPLEKGQSQ7vjtIimgszx1FI9axXMM1G8I5D0hYxQkJk19dLtEH
lY4f/gPYOhhQsGGBDSMcm7PIbVcIACOl5F01ovkj3fq/OR93LDhWYaP4HnGvfx7D
OkBLNre+rwgZtZAPhPuN38+ecb5QJJ8eKC5975tmMyLPDnKd7C7ZBAhSIH9zL2tP
GSUXs3JZAVuisqy42Su2ekz9PiOK4EKSGaSxRALlC3AokzVUsRK/OCdj6a7jrnZf
8uhXJ/VQOQljQiIxulQPlY42BotwI0v1O2ALRB8R1mVr1/8WQiRi32qgmCzNh/9s
LJAk5Kp+61TmsgztZDk0PrEz3WCuYMmy/eBgFs55IYYGoW43cyCLl8eFTtCnGLtc
Kivu0NITJdjEUS61jpTYk5aEjB0GYjR08T+bhe5EZl0MeA0blmEpw8rldcqW2UsK
xeZOV762co0gL3Sl3vSaDxYJspyKq1c8V7sC2+t0GZchxtDqnHToNhPt4o4KYSDZ
umQvLpGpHDpd379jpzs1/odnVRWD5o66PIHHMVfh+dbsPtAHI7wPOlpXLO6ST4Of
DFrNoDvGWmJhvB58ZSbvOW4pwbUW7YuQcTi/z8w0/JlmNHtSEcRRhO3yMPLdH9Yo
YvaySxrd+Aev1MY0TUPLY8mzW66vRO6+2Ni8heG75x68Fan/1Y6Lv3yJGvs80tXs
D6V9jvxsXA9MMsxNiwEWkr5gMbuP/LEX4h9mLHdAtwC5EsvA8e4zU7Ip6681MIxw
OkvaadmdyXn8s17FpLPz+JyA0+W097Et2z3/4//boabQrAqGa5h8aOjsT6WDV8Iv
gi4sMPrjA8bBOBaHJ+nKO2vVVu/AeDgpZGp2cDADArBMOAlxVOVGBU3zczKohsJv
5eU0f9waw2rSALmni/yC7RDoSWLxeI+RlweEP0YYMOAHe8eL8uPOe5MboE4OM2rW
R/vyj1Tp0/vGchlIDmEuwmJlddKm5cYI1fey4NcH/u6GRzaU9OILOJ3KbmUp7qlW
LWTTBtk/DMxUoZqM1GzbJsKeiqKskDn3jeqVXFnmdMbO5GqYH8l4NgIXksuUueEk
yx1fVkAGjmckaaLklL50zT8Ri+jX+qf8VRr47Hk7EXTWQCXe6I+WbPQ9/mcAYyRI
oIQ4bBGoJDydp6VR8KlVfN5+pE5w4kuOKPmROaec/xxK39gMaqk+713pQRpRrqIU
BkBnn8zZi3MEHEYuvK0i8UTUqZpwZ05j8fR5JPlbA7+i3L+gIH8aqT3W/KLWa+fe
c91wUerbEa7elfQ33cS2QU6PZSPjwdbmCi4s03c8ThWlqGRSQr7UmCdT6N2evt4F
CaYXnhTm2izH+/urv4tcfK6eS1DF5mmaIasWLhJmtAdcmZeWuwFqdLcoS8h5QW5o
zwvvNQVidFxahzi9OL2AuAg0/7qKRDDLwxWrbxHB9k4kxdklDziHEwc1nPU2wjmc
YNphV0JfdHjOAOTzayG4xmdN70SA6a/B2i64s0krsx3QYl+c5NRzRU03KoAjLM3w
LuadDkLAlbKInyABRL4FPJ26/tN4ZGxQw5s2nq6R+fOfGFIyYijFX9XKe0lRKV3Y
a3FHezufuMmVfCRoz0augTD0PpPrHSF8trej/kWONGOwrNpnCdT2XuNnpziw+vOx
6Bk4kX81f03aeHc1IUyoksn0Ele7pJei2f2zoyLQdIx1zQGT6U1EuDUMay/aK1JP
XCsGdgAMl+OUkXLaKzIrnjCdCXqaD2ptu+CifgUp18wNjPgffTldTUQnLEuoIonW
eOs8gGa8PTz0n492SlNVBJhXSeD+Fx4C34Yub9fLUmb0/OHCpzfWcVqsfTXnDTT2
pSXi4FUGB5COa8uGmQ2HYj3UZC67lWxQJyBnbUzLiqQGoFc4+P132PWwg0fljcAS
nZe5+QjOmyv7tGyrjAp2MWyKbCtH1KizKbheNIOuRM11Lkp+84sOk/JyhBVyWaLm
4lf1jqCbwuTZVQouivaH50pqJmycWBhnfd7el539YvDC9/ALyaD/NfBxoHSyGuB2
d67Rq0kfQi1xBNNSGpEND6HPhsXBl99wEtLjwRwfjVEXkjIKIpAzTIvem3kVk2U+
ZlUk23dAlCh595ijO1MGk0Z+sB27cZJw86B2ma98NqsEkl0nJmWOINMes/f0d//u
jNLaLx80eTYHIuGJUJmOwr7h1b0ZeEERRLEIh6Xfu2X+uWFcO1d4eFZ4KN5BCakT
kCjLfMLqHsun9MEgtQzwUK0nHovB59qfD/soOzmzMw1moZTHAtbbpZHonzqdYr4/
FBjT940OLqhDhRwRxaOIgy8xud7/Lh5dMTQWprTlOQNYSe3Z1L8YAoj6KEslBDKj
mnWhVbj/3vc0WJOOA08XKn1kl/lqk7RNZOmp0NS+HvIw08H+VC79WcnKRxNpT4Yh
JDgRBrDmaPU8uOK8GTb3Jd+HwleSSK6m1C6H+yqK8B24BL7ER4WN6TGhJIm0aYym
DnKPdTzLFQKIVNktK9Qf7w+6uFUaXEpHhs4U1WwxQz8IYGw1+Bpk6V0bIXop7F18
aPJDKqigVvW8rFLv+w+ThbY5eAiF0iDn3rgrmEC84qgkCeZE9Y4TsONyVpikSlvG
Ss7h5n+Q0h02wlgXfWZ41B6PC9rooG4+ovvgh+nmSOXxIXu4694FanLt/xXMi5gL
Y3VWys0btf1FquYqcbz4x0xzNGt/OnAoCaZHm3zdJaP+ft7qYTq7r5yoFFBzzb8W
cMmvbXPZBlATdiL0hLHPRpJWNh8q8zMTiC8q8Ah100rQ8Wu4QQgohB64Z+zH7cZv
nHXRLGTqfEjY1ZHCjuCku5/O7LKgk2jZr4c+IRiTB1PnIBkvihl9MHakRMmvL319
Ur4q7eFQ3XjbZZLsskuqyOcQKetsok3l6efenDPtuZZWkDpW+0tQZu0WkhRJUCnY
TAuJaizzRg7jy2Twc8C6omjCMKCoDK71NRcMILI7OzJTWztqjwSp3bp/uMgxaUZq
AYjzoZeMfisF6LF1pYul8pnPwlqencsw+rVvP7qIn91AG9/MOT2hkfPBmGE9YXR6
Ksr42qsfuZAzBLquILSZvQUp2DMQChC/xR6QRH0u6FizXHoqcp3obZGTygA4fCLb
qO9hdvqv2Mvau5JV/W1vmJv3lXocMo3grX6C5aVg3iv/EChChUJvRmmrugKBhXPX
RFUu+P1WNBBH8TVd+Jr4ap+dkOZKCyyj5t3zrodlpOKNwgbysatVbmEQ1tMHyT03
KL0kHNImUVLluRtk8QLxM8pR7pNgAlNdeB4+5e90YvGitkr9XplYqqGduNuU5VnV
/4EfvCNIuia6xhFJOGdHCJ74iomAqE73q4pXe+rwxxAsPZw2wE/BlT/BcpCVk+oV
X2Sfwuf1qlx8KSqS95QMJdFtqbHpc6tjqwfEgD5kg5m+myb6QsEuFaM95jR7a6Rp
1rYlp0P+vMSnHE1zZNAKJwYci+1oJwFn3g/xH0JG8M/jGXWpDo/+m6s5ZBCHpZng
tI2+XWEIVQdKLp5Zcxj6bdCYCyVYS6c9LNhvFLqeR7XFTolqJWHXybQQZO2GjRzF
GGaSMJ+vpYDl2zfsqYgMpkJc7YKV74mfVpCLdYNxyWPs2I72GEyzXXMKKF1s+lyP
8dh4FZN34U0YJYK7v1AbCtvswz7MFES6vJL11+CK/QObBwGCoGCh7vw957nwDB1E
HxEEB6F7K9UJSq/TyPWGQwFr0LGVerGKPc8RQeZNDuXAxqdB5nAitWsYh0VqWZ0m
qHOvtsb/aXAdb3J9PPF+q2tZ+GeMDIGOHCJK+SUCHR2oRUjyylwPYUsKbniqHvQj
0G4sZEGn8AqzuS1FZRZWFtUFsrEsYF/lTtMmiPE8VVmYSL+3oakP24jbo8RQ2xD9
xCLTYx/p9Xt390IbGsOIKnfvCKqPEO36Cn8ue1QxUPTt3MQvSrc++0OIPmvMwP86
NAKoI7atUd5kHJcn1VmVVLGmW/RSfz0Nhg3OZwAnmk0SBVwURpcirYE0WLjfPeBS
6c7LZYxDGVQET5AU38krkRRrmRxMew+DF1JmO4H7gHgwojjursP4gaChep4tJE48
vBri0STuEiVSEtkkSH7J2qcGNdmbFs9KTg6a7Vb50aDBXRbKzZ2XF+XOR5++R4ic
iiR7a/zqoRYyz9OnHUIOAHDnl0Bz2r2WH2vdVG2n6dFPfpyd7c52XJtO9fC+R9Gq
ga3a+jxkJcTxOF0fbE5ygjogrFalhISBBDRUQxXqIsYtFVtWY5Pe1Qzt8qy94otN
WoN7dbM2fH7EbtY2n+CfhgZ/oEFEv/8kvYFN/7law3LXa6n/taqlZ/0KFItT5r9k
SUaVJP6GriFKatzqZUqS981PGWnRrkahfka0OqXWbx+KDJs6pzMi0QqacGu+mnCv
DkyuWuRhZjGOfjrIo9qazCPvL0N6ZZEVFlXF0i/vaNZY/ZJJQlqdSiM4iifGqR69
TxyYwLQ134ISrWYP+vZPKojN6LeXZxSP7ci8d/aF30Fa37GkGW/BG6eN5kxIXQTd
RTZmWGKQc9a+PrLKqixzezSahfDH3lc8SnvpvYZcAI9ypVjyJIsztkG5GgErk2h/
Xry1BJ6l0JYdVkbquS++pbKdRWYCEo0j4IkORwiMHxb7LuCPv0/m60tI6zn4WcAi
vHyjUntSsNDHZrLzj57D8R3D3LQjRWp+e2FW4mIGc2vlpUNfksAe4vZuPrZMqx0i
s1is917e2rgptfBr1HAJn8UGepB0vR6GpArRKbaiyIcnDeyH9nummYKUtBn9Nc04
bh1cj8Fzc6DojmCSy03ZT0nX58EiQc8Im5pf4PS3hBJ068pgUABGy6bDc6djVxjA
6nSmDvfGP0yDCE+s1+MG9mazpyYO3STXA9lgr61A4wMk0Wwg+tuqlcEfHhTIgWKG
hLulR4Z8sO5ftVou/HESdG1G9/FDUhCtkzgZaZXGYkJni6RMSVjwEkyVziiRUbPa
4k0DlPOWGIbELBX+XkP7D4nxX1FI2GWS/GyaKFtqeKrJt2zVz7vel56jsJof93aL
KCE+uBB/4ve3FJpcRg1JseVvoX573hgVDo51rwWX0lEE9zMylVe+hLKya5+V44C5
CtbT7p/ZidV+OFNp5bdFTz6JVXRyUJ3ped9QN6s8tgJ0oiz9ka31IHdBMzpRkCAr
M9f5Jkf8CGkvWoaXASJhnJ9dbMvzJBP+7CdWAuGNKrlgENwkv0oaFXkfZtSifA4Z
bY/Tv094WZLzLcBKEUxze2xcSW9PZc7LEKBC8PpWDTBmRaAl6kYJc7+wpS/slzLd
imXZJcn+La2ejrL/k7buigoQkWRZ3dj1Trc5mgu/3Uw0Wz7RtI9odQOZxn+Rftap
iNK1yMZ2srrC0CCiaf0wkQvgD8OhTM6lV2YRSOWXNIan5lIo4DJqrcBsqwJWLYeb
TNbwBO+4iDQfmHWUfICBry6evlR3PeFxnEEAZb479bO8n7o8P7LmCZAfEUODhF7y
0ANkpkm3W/XLG9K1usjp08t4usaDcjWzxIRrPUPE6VmD23pDyEpYt5bALMa/zceJ
GxWpcI4zb3zCvbxOSsXwnmPIueIfPGkZnLVIQgnNGcEY2CCyA8pAYpWB0O2b63zf
S5foW8fOE/Tm2oYY5be0Mg6nvdaP9SA+lPZ7YDs4sgOkVf2vzusF7cAhC9UV/NZA
riA2+AZCld5RIfXU7cDtKeDGyHHU2uT+Hn+2lq08mTB4YRqclHYfOS78UXtClWDs
E8uAJ6rh+3C5uho1Ayr95hPUIEH2WNnrsttYHeWfEZ86GGo3C+TIkPgjA46BIPvD
5vBHQoMV31FhV33qx2qckR/M4eRxO2/AaDHu8uvQz7efghctC2I2Pd/rjJh4bJks
M8RriIRpGbnaKpKwpT/Yc/YEN1ejQY7wCrGgIFY15hNNUzpqFxLbGlytjUORxhG8
dMWqgXiKOrnaEUsEx+b7eMYPI0CFJ7QH2XfKWACwWEwFUPl7pOM5oyeNKlDniuCi
f5WTt8tTrk9jWXd7kkefkam2rpRau1R6P2G/PLHQAyxl4ZdIGjU2+/UL0BHVdgcY
tt6WTAesi1qlLTQ9qqRIFUCEaK/2eUETeif0eDh8V0/SJnJG/2mPFn6ysxZW3XQU
HVJg12j2cp3vuEQkUVXuIhORlTle8pXkDPBSe0y26oM7sd/Js/ioKWO/W/aaEG97
ytj+qXcmxD/NMUB7OvQuBvklzOmimFHsNXEZmati+vrPI1wcl57k0EPt1QB6XhFO
0N0hlXao098ap75+jZVApzV/r+NYNHR5e6JytV2RntCX6zargmAUyLDcvQdNPFY1
JDAz6wxPN1kzkf3Se9OzmqY9Ys7n1B9pcO//uWRuovTZPPzitf/VgPM1Jpgv/Z4Q
Sw2o9oE+M7P5Z4mgR/wTzUX/RBCNT0lu1cqt8/j/ou0gf6oI3+P3vdAKsApGR69o
mVUfND4iY7ZHYu36/hK91RgocBTVb6yuCQSSnXp8S//d76Fx+rlfskPaef7RUMpz
NBO02RfYhaeayTac+aVqX0oSeTdm6FwdzkwD0H0x+88AKSi0Bs6OP7nSiPaoJmNT
MQpsF/seXiE30uLXPsrELCkY/p9f8Os7l90tg1wh4HuAT9hSxGdoVUq85Lp6WioI
vO8hD8xz1JjlSiCcHMV4CTXGnCKMEHorYDZ7I8Wuir02x4YvnKYBbuKuRBUjkjXr
nk0HZjlWlSoisFZv8Y5FAvXfEhnGI6n81bRmuJ+PXVqgeXVmcH7FzmC5kLRHctYw
PwFUoEXUAOnxDS7JwpYQTQM5+uiC6r4zUSR4C2DxPAiqRoCFLkttqk9nIC2dsyl9
rAK+stDY83xAUu08iDdCL0Y8LyT2YKb20R15MB4RdgQC/LBWO0R/SSvxRxBQObIc
A0AthRdjjNs3yb0usSF2cO/DiDxOwi7tLxtzv6UEpdOTmVOkdwBOB/fhVc5SN3eO
3L61rHg87ZSEAUQRlTfBOw7YlI1LeSkWGviYOMPkxmhPjSseHcSxWe5bhBPtlm+V
4OgpwwOH7brFY6g53veqxFlVRpLK0BSk9+YTKbuJ0/pKspYy1fyOQdgQd/0x0/Dz
7AtFg2SNLKY20WMhqvMW+EGu1TCSjN1DWAI2nfLmhuMgDEhTTnLoNi2AmSrXeClU
FtfZQqPVoVcbHgF/kKfFsV0Z52raCzpzK0MY91z08pV0ItfHMVpgnTPEF9+G4ozi
MAZaWZFU/EoIN1N/LU2OQPFVt2rbb42Nc8aNY6m7AMFcLIfrBy57k4WK1MzVNJ9p
KRn3Ntc8OqjFci0M+gBplEbhecI5qSaVyOB29IZFvQpzx6SxHVTMbxaauP5i515N
2y9nOZUawfY8A8iusojSxS0/+Sl3zsSbHvHZ1ZO+ykH8zs1R8dBBWntl7zQOY3FO
CEZHzNcEhWIRL1YyjrDRncjxh00ZKa56x5hF7ZVGYQhRoSGjWwFT1T2B/2+9im/b
qoPUm/AZNb+GE7lbzlrg+F2qbDMiXudSdPeMYvypUHx/qflbGNMviFaDZseQ2AjG
yx5ZVOO1DEKM+y8CkSJK5fFwWooEvy1Wtk1qbJPDxDq/oiDovs80TGVgKTsU35VI
LKppWsCgRxdu5Ckt/kecO/Dv5o+tqIiOUVjQsGpjUoomtXpWCMkQ0jHHRCzBSCkQ
EnF3KYMIJ2+kHOTYixwP40Ody4hbNAR1S4irWKjJN6HnaydiYzZLMQfZnaHGFT2Y
e+dPhWOBkIJe4/cq7FDyAltVpNUNKaBs1hz/+qH5Ri6fPUZ8gSm0PhDsZ2LJQAS/
ASlHlByxHWaicLmsk8Cpk8lDth0XWeh2pV/yp+HIl2saRoaEyltiW1wltE6Doc/y
4RPVroFN/WPMJSV0QOWiokCbrBd932Rf6It9a5Jy96AQ8AfQEYlej6iyGOSbvx3O
Ei8VwVm0U3rYcKfrisG4RK0W8uwFdexYsGAtDRL58l1wozBSLrTVtyefVzj4Zr9x
g1ukU4R00JVFToKDbNJrMLgQRDosOJta2JVHaljKD/SiGoqZgf0w8KrgurwvN6qs
a5pC3QGIcYAUPnl3PHZ4/yvsMjFdI7EyKg9UeZxqVCAz/t+2YAJ63R30I0j6rK5h
vCxkgxHiPo+kHcOa8VWLD6j23rF+UegDf3638pXSZm++FtEQyOhPZ2ErU7fcLtXz
tnlp43x3NDJiycHJ0jWpFZY6CIrKF5QPIMv03pzsQYH0fhOYvxFbLXQ8ZAkHtNui
VPZ8c9sDuedUwPwgrjuG2OemVjAXLVevDCSp8Hz1qNzMs3rcqAWPtul/DkBhzl7s
9ZQjW/P9A60bmrEO3TJ6JP+ch35aApaaYLoW8lL3xaablNxQ1KjYoQE1Q3rgszwX
j7Nl00sEd1gZy95xngTwswctPZKXG7QSOmToMdpoRLZcHZK0WDRjEms974cj280q
iwDy77w6Od3N7mbp2eIFNCXf0jPq4CoAT/b+Tqy5831eP4zN1S1IhQkOVTO/1fAA
Xngz77YmWGgXx17dpWSSFNOgY9qtzMG8MykelVwGrEMs+9ShaJF5Uo1auizwYkFc
/Tifq7cfxunvJpBshomA9VtBqZvODieH5cKlIZRCOTBFWuqqU1YXr+rI/qjbgjUm
/0M/mlW0NWxR4jMxlFUvWbUXWBjh+br50TR8+bwFnIITZTqbq4qO16Qa53P2HWjg
X4s/j4oXHicO4iN0pH5/En6PAfupoTl1SomNyCQ6M9dlS6yerUj6YFnS3wyFahaj
rcRLLYmTuI0XcmyU0ERI3PS/wSMeMUSPDqDVdmhcrUpsYhFtg08Hxz4XdiLm47Qm
dQ50AkzJUNkrbE/WrlG88p+S0CQXbxWzMOE80R9nAf/tmClWwwZl6382JHlfY5iZ
jLMFl7SiJf2sgLH1iL3uTrgvppxw7K8dFVFctXUlNG/JJ9YdHAvNyUfv1i2uYAhf
Db/22ouc2cLUk+VGX5OFUEUohk3t6A6jIBspLBXD4HrJwWe0TpL/Pq2rJxXgs8wQ
/8us+aeMTQ+YKAou8VRAQShJxp3PGeSJWs+vZ+muEZ1Z4NWz3undw0WhOKLb+Bqr
RFPuFWZ5sPfgPIjtrk/bdcqDn5J3SFHqbjchgmS2wDJoj4G4pKlDJsZJzq/Isxsp
Jc/y4DIJI80vNf+NrCv2G4vrI4HSrW1mvs0VzQnSQIWCKUQPMBzU9kTJBJVYgMNA
5QARKaa5VdlWouEzqK0vn0ySlZ4Z620MB7/rQkwf5bcbcWdjIyYrDi1zQUH5AeoI
sNlpEAhx3QsdxmL/mziaocoyQgLPTgzC83HShkX+q60nKwOkScp8AlQu2g7PLxx1
fPF83MKqHgL3EeYcUJOIm2ZJwsA15mws/NMSFuZyJ/yg9P2uWpKf4jdwDwgBVp07
NXaCSYqWAiPl5nFeJqOyX9L1bZc6seTWrFlx3sCknyVGPO6ax9maJSvBknBNO7Um
Up68rqNGK88q3DTnJKg7Jmv7k8jXuzcukkudQlkCY44K7Q5it+9jV3ZiVBlsGAFa
/dqdLSj+m7FQI19cWdIZHS/+tNPN7DhLaS1CWax/QLk4JdAWG0ytOGPsNPgcOJ8P
aTQPMSb5sqvndEDMlcUuZl72gT17nWO3VfhMX/uI015Ha3qtJ7j5uzBO/RvNTqZ4
aGT/qglwqvGDYwYvmU7UDOe543fWHPUeWEblkxwJTusZ2EOu4uOj21uF03Fu4PFk
Ln9D3gAf39ORlTG3HVldbSIrauVUn/9qOznniaa9Qa6P5sq+yioKBxPG+kqprF3C
eg6q4N1eCRR9S2uR2dBptQt4CRpsFGbnJT7QPPKcyz7WcW0ukiao+dRXx++pcI4G
qVKEjNywXfn+gX8NqU5z18UGxyHPXbn5Fk1urgBBnykR5UnqUE3mDFuZFEXeNcIC
iOeFjavvKwnBQJk/UPeqn2Gqi/z6BX+apUrBqo0iTUuBdvPzvrHyPldR9AFSWwgt
+NLl/aA+3l76APehxSDuN5z0IcIM6tNlmmU+nOfZNj6bSz3mVz8vKHSn3FSjDh12
J5Pz2hsaj4CZfKCq4xEXHWvg3vbk3QZiNlXvr1xuV3k6JOiFgmLF/FpzOt87yrX3
PHGeuFfVwY2ADvYa0d6POa/K2hDwJyjv7bRl8BC9krJ3jsjiUjRHmht/CBKfI7fe
DladhPV9Q8wcTsF4qtov8JzJEmYYOUfpygRrb+a/6SAIZKgVRGPJgMmRD0qEYfU9
OWSPymx9e8TcnPzDSkFFIle2nmWPJW/56MMoDEPlynyQOa1CiHrfWnEwfZvyD+PD
B3vlyuQrGhhg+ZW350Ob2xxCA89k4wecWV9fUstVRyAUJ5AoMzhE5iPrT5ZdUied
JvnXykwJZHxLRecF6Lb3Pu+iOXJR/xWrZhPwxzvNvPAVwpiJFo3B6K/paDhDlYgr
dY51RGGdKIEu46e5v1ngNL0OvJrw/wCAYcNIgv8RRQdVJDJtEtKojBLAtFQFCOW8
pyct9MBRBiyOROsmrRui30cNz7e+uTec+VS94lPCAWpx9sIIjFYQlKN3TO80LSFq
i6L7iCJ5D0OE8m+3nbZAb1Enedv9ogAQyd0830rfZfez1NCUFm9K9AmBNIWv4WYW
ZKNQsjcMCFbhOtnFEZeq6iyXYhX61iIoS5srtoP0jyS2Nq+Ed+3vthvmbEUw89w3
UUW06Gk2jZwEqcd4D6hczc0MfCsV/Zja4AKGi3fd4eKtLJqAKUEZjufLDP1xMpx0
+8lgfyO+lqZ+E38zUAEAryKsr8DKYnfSu8RFxJ0y323TF4xR09Rz77SHA3pvyoMJ
ifrblOc67pxVfKSiRdDazppCNX8cbtS5MWGPxE49HnPEA0KeHhH3K/XptyIVUckW
RnG0MYfVTzfmEmJQrFHpbZ1kZxY854Jh5psOp1D83qxP0gCCzm/Go8MSLs1UlrVL
IL/2dQx1weJZ/uqvp+DgzVZGTFVkf34yt/E5MGcU/4ezJspFDtJziXXG24uIDAQq
HrL4EtpSgw5nPwni3LShSUDpDkbTtFtP8GzSbSSmAODMFee+1+A1rymLxAXQmeDt
GtsGgXcFPmZMpSXGSVh7AkZ3Xp4EwmF5849MPcyNH1H4u0cxoegQZcjWsp5P7Zg2
4jsawVvDQDHLkC9GElaMteaq2L8x7QlilJhaFHCoqiyIvbU0i2posjM6FY4dNTia
QrIn9ZMcpZ1awBqLjJZct3yKiLmI+zctiKRI7mjYe1tzomEYiZC8GmoOmEiQ3iDI
oLm/EC6iVjRj6Kpzc7Skn0VrpbLmPDLTq9tJe371rN/sOvOt5FOgnpAjkeGHPjoA
ljpk4P5xlGOEBGkE6h4nVJ9Oggz8peJbEcZaeBttZ8EWehJ2+4MVvlAW6M+KJ0rJ
RJTns4hav4d+M75AwTGSk36wivOD5NuvRGDkHeGbyAPZto5w0M1kVp0/D68NC8ap
DTd6rH3hCG7Q2fq6f7V000uV1H41WVym6/ivRdWWVWtTmpA833oLNOJ92R4P/g5C
Iq6QpTS7iHdWRPPhMV3te23GUpUt0iBYKFF5Cr3f8POwovQ1EKbkimonUcg7B2Ez
Aqg2Br/ItPHJRueQNWw/zLwg2BtYMdmMgr0FV4p0VFQrBUzTmhe9hsH4TgP+Qzok
QfpwrG/EdAnxz2bZRSemzbyAJNw/ddFk0mIbyQhxnWsrNhKcHAdB4PMkW4deqAc/
az01fis7SexDawoX+/TxLf4Y5j6lKuYKfG+UlIEU80JajKaJGgRe8dKQQ5ozKwn7
QeLh2gSpfu+MnRiP7G+0xUSXtJiNO2c5aE7lhbgahRB7/HQF3c1kIVHwbqRC11CF
d8GYLy5PIvJjKUYyqeD9cxdnPt08KzLsg26eMDS/Z4kENFf8rSb+rWhRWqM54ka5
KUtVqik/Vg+eRmEx7WeHlBqaBpJ+zdvnsBICBIX/47O3NXZVaFqr706LNNoqJfTz
Yjl21IyfILhIlilSHop58f5rHDHDDlYnzCEbGCoHJoNC8N3taCqEimDi3HSVXE46
0Q1GsFVEUZLagLem3ruS8Per1hF3+cfYlxQJo2V4CIo9sMV2HDUSA2qEqUNEEMVu
TkzgPr8FmhFOdqakTlw6LZk0C/RJrajxQjSbHTrEs5398XplVbgjllXYTWVkBLMP
JcgIK/4OtkeBvguHKBSWBEA2Ij4kMdhd/6Ouv5gULRSqvIOMe1SGvgb6+lNn6XtD
1B43JIEhOmQk+/qIcmMzXEiz1Q8isZVCMYrpalFACWZTdm/rc6C29yTSelXG1dz+
b82B72nDoxqPfD5S/T2yOYLONX/nzlvOjS4t0Wdj6a56EB8dm52jCocAlnDKHMMg
Y5yhZbgEcyiwt02moNX5Kew0KuqqwWG6DRxpdWpuryLN9iEAC7ExYdqEz4ggC3oy
X+fm/43+n6zqqAvBnXTl/Hyr85RfFta7j2l1mh9blAawLOe/U8S7/67njcANkG/P
cxdL7ZI9BMz2wO1t2ldUazdNqjKfc/zWd9lzvQcaCO4i42EOcj9JA6RbEAuaDINb
6leJK4W19GYAl7xNc9b+OKMTf93+7RwRh9bE03zkBdvGYvHC2mf6e8YlhTXbP9qw
O7+5ORMuCuhjTxzxR3ta8XkHKNNRYL/B3cBEXqxfg70bAfGTRDHpgvPVmtVsB2TF
wezO2ZueCqXX7+tCGlURALfTflqJWfiAPRWGNoCO7cxhqsO/uVQD9IEu6VeeUHCB
SY0rUg2jQiq0hjVPqaRiUsN+cYjBoI1urwncE5RYEzzJ9rSFNiDI16ya2hXa1gdb
lT1gJJSbqNmQ40MN7kTKrfmlpGm2vNTrOFDJjOiyCKBl6RiyxSAP8WgsknjmmVSK
rnHzHqZt2MguAQDLLm2BW0Ywm1F5exvtatoliSzGcyEn5qdVFUx90jw8iOsUmQRJ
J63bbTaAxraY//+8bSQZ/tGwaKQCLOsypEe+J/6zSmnjCWVZ+Ccki9KmHd30p8Jm
AF8I1Kc4BS46oCSNNua5K34Hws1KQqVDK0TG/VG7ml93y+PDdeld1NWPBXFANRlK
uiATURa9nnNmze0LWYVAwNREQStIN1Pi8ZyhkhfC7Px3FlO7RzzNjlhKQBL7sLYb
k0CSUrjPzbdx5eNstt+BjZXMtfwotnq/PNcobEx32w2XdEjKmy3pbdmiyKV2gj7V
nwagFAc8idXNQL10p1EIs2tqkYnbpL2G6sZ21VmdkUpvH9W2svX9ifxzQe7TrW/7
iKOcINPovP5BGugSOQS9I4lbdD5urvIyj3G3cIdglTBQ4UqZWLvBVWTUn5auEWlK
GBDjPjL3ZqGy5jaL4+oPHv7Y1WCLewIoL0vICkc5JyiIH4EjW67p5rYC+ApvqNj9
GZq+RFOICVRWiO3eajs6mbSsnWg80xpJBxaLqExaXhxROkP8h3w9EhEXtRK93/Hg
DAStHiS+LUWEeZnTlwObuIO33xzO63Pz9m747cxzxVAFDqqmc6dbouaVWdmL9FDf
J4ZdILjxYqLAGnXXL8zvY9EWy1qEJdkUPnajUYyH2rrbvwnCjswsCaUDrQ7VL8kS
TsokcoYB+MbPw2vkP3TvBds38eBlt716Wz9Xu20mOCglG67FOC0w1cH+MdcKkKcI
bAApLJjSNp6vCFLpe0ue/0xgJfUE40j70ltgU2GwCVTSR/itny9+fR3siY4HwZZn
vkXDTxTP5YsFpdX8VlEeHKH3bgUPbrKI9sp9zRXbpzvRPR0bKxp/H4U51jKS9p30
uzKOhoh6FcQTq6GEw5VKphCiFjCGqESMxLUOTde8wCBF0tyvzl1W92/9fWfW2U92
wdz7OhWtsd0G6fEdCPHMmxHQ4GtkxI3LXk7JgxHB53v1QwRxyX7P05ojrYiysi/Y
uUDdw86RDC0yd5C6u8SPDKv1uLNKLu4gZlaRk8rQOVJ1JznBxxOWhrIwT1HIVadS
Svd1SRYfNcREjXGAl88kxGCxYALRC7+a2zd2eQm8p8UcVFXiNAs2k6PwQtho60wm
S5AVs0JnN6JuXR7GrYZX392cLCXgPnwWBMTDfdtS6v+hUkRx0VnWtRX11rNlnnto
tL7UR2dE0JjcMCOuaqWedPnUpXaLB/2syASuX+2JEjPP+nyzFqpuIoxbGzmHGpAZ
ywZfXU7cTdmlNJ4uChxQ0OpK/ZjY7k/Olq4rX8GZ8LKTfagayiaGxtGoogCuqriQ
ZbUwQ7H14OroNwZWNvAz1U4u+XyvyP6SkkCI7ghkGl/GIN+hvY8blFqy2qMBT39P
3iWLco/g1ihiV2sPrVfiH946T+5t1EUiu9NPw8NSlb06T+QcuDQmE72Nx+RGiFQZ
2UMrB4N186o4zzs2c2+u64Ulfoe5sWPWWL/a2fyrUVJFg1G3KmkaQEpDC5UiaMTW
Pawh4ZFHfJHixV6riUhmjTf+nVDwx3/BAlqCH918j5/BNV6lgD8Pl1AsmzMmoDJF
4sZngJSq2YRVgSo1LCo8fT+uf4qtdOo3ST2uP9rkbOPC8aqWMJppKaeN7+pFSNqq
9V0QUlqYKFKa6m6Y91bI3+bwejDjL7fx5ye2+DYSaSvT3+nsLZTtcNrsckv30loV
sY0vZvsCh7OxFxDaY0qvJ4CwxZrufu7IDW24bws6NIvK6+DhMJvLGD4Mdx1DlTCe
hEawXCNlH24AMxxTWD5W61LUINfKDP6moV8bxtgOUxE2LzqVUrVQ1pXACc/qyfOX
0WpTW3bSUgPQFlKSiKlnDWd4yDxW2N+M2A9lJLmW5Hqj7sZHvYAF45Xdv8ol3EwI
HV1NStaKWd51tX7oLq3Ga92gk/nd0yn2RM/Q6W1HGycGo35HsD9AnNms2m1eZw03
ED15yaYARGKu2M3E4e7OMchbfhoMbGoLWM9QWamezNQR2XaFI5Gv4nSlI7vNl46C
rdB0KSmJJGvof0kGBrjjfZi8Axs2xiMvVHdb5BjvE0cK9ilEpP6ncfrISVlTq4MW
yuQ/CAOW7SpzPFTIegBR6iPRaH5OwUb4iaifBAmsCnslBP558HwrmMbMqFCqQdG3
pkQH9WKM3sntrR+Dk+lpo+3WW2IC8BEePgh8koCHP1TY+bADPuRmyWSRCbFevehr
pQOL6oGnnrhRJtaZzss9hGUg0++odUI+9R0HbWILD/UVbDyt6AxhlAwSll/u864x
ANU7sAKuDKc5A1S3esMFW6WlW0vT8yDwJlhV3lk8zDk3xZp3Fu51dWCdk4ZewSMx
tJfW01wxTzYAZnqRR9b0wcwo0HiVHAW5s/bfMSdq8UUIZbGe8KojqcLcMr3UYQr5
twPHBB4Upt2jaDbhGdyLmw8KJu51VXi1TSqd8oAwDgacj9RcHCpq069yb43sDRil
s+Z+eY0Qw/NDU/M/mkLXuoB3tET702lpwfBn5FlPNUjBxryq9cTE2o/mZz/GQNLi
X2VQ4rCeHYbI2Y7ho8kvrtix41Rkx+dodTSTNXBE+1UudPioQz2Zr9Y2IiYDIXAE
Hy+3u4hG7AZ6xaC4p0HVQFjP4xsCS4ih9su396J+Jo+UPff+nLG3kA6ZkDWFYULP
eP/GNs9WV4RmQsd95SAqHVN5EXMQbAq9PJ1u6puPiBAkoKU4yx0geA1u8XklAwQv
iq+egEsD/iOs2g6mHlLz1Vx8f1HFkAilpW1bQO2JB1NEQ4oHyU82cdLrNx5hNLTw
MuorcugmsnLPqGpvGN3a2VWj7eryFCSzflOjwCLhp01lGW6bUGhYmUKqW5HXNPld
3QRIfHLREPGq0bcEB6yF4APk8liNRGUAyZSiFEZWCHvehOa2mqLlKN5TZHRBhzGW
rC+nT6BUr98zh2j33SOau0PtJFuizOAwJYGL/osroa2xeNhWy5JgFH78p3ECCicL
vla2C0pYu3dw3cucWU+TrXjvblAzRPGXQb6bRrnSHlPzJHfinlCC1jtEwnMyFFMq
HsZ+InBIWS/Xcj+Hjoh3koYKxWMxHvFEOd9o1Ol/GXdn+eYXmN350GLTqL0zeZrl
6Z2+ZZoQN4rejPQP3immPH7qmIYSN2h8EIiwlYSNwhfLXVTinfKlyyrJfV8Y2yb6
dlt773RgsYnKlL4ZF+93Ht8NjN4OKUv+RVlTGgprfp7CaN52SLgPNwVY57uEEfiJ
3Gvo1wVPjeN04H2udo4jmbmrceEax34bAmfJOS73ggbx4GOo/15MAFgohnaGOYvd
fdX/yFWyJs3fNI7Cd/SjaI+1+E3w9sA1t+dIy9KhLaPOTNi8VPFpLhZA8BuhZGrD
LkZo8RAlGXvtlVxOi496WeRiYYUBodpGagY6QEjeQHL7PlfhexdhuvQoQLWFTNJ8
0IaWdC4LczVMrbWgbcx9BxQQDNDlRpM9R3+lthw4w3LNxkq/UsL0nbCU9hQHGAN5
GnYQqVaIfyZ1594rrEMI+KQYS3bNcO2+nAiYclVb9+Eczt3imJ2mblNqx7GHcatR
zRJtldwsDt9EB+gkMHKipupA4ZZrxapg0Vh6KzrWd638Mj7v7mAJ1TZBmtgKXpSL
Qx2FxtFbSMAVwAlMfz5I5/mjfuC8m/wKWn8aUqbVfybu300qVWuvCOMdNPmyfBnP
o/TEAC9ncZJeLK7OmUTCZ64711cnY1L0IIyAE1L9IJQ/E4Fs49xCw49ZagZEtD3z
1gvkK8IDfJlUatCsdCEsUjE1hsS9vg68A7bklAdfvne+P/vpzirkZ7+23LI80aLf
uUp7UpcTJf96j0BbdvsKWPnqKDSsgN3IJKLazX9q9oQQtRWoZc0sRt3nLMghwzqF
LP8ImYSglHu0lQzG8z/inuU/OSIKvWcEJBDCzRS1yRHHuYSFo3+jn2+6lRCePlJI
McLrM6YAkPJODMMAyzvRjePhJkWbBoUbaUTaDsQFN+QkE62riYUFcZhBevJo/sCP
XSQQJcsQ+SS/OOYawUAhlg9Cb2AQVpdrBJsozgmpQynRRJiZciWVWYsnti+GtkQl
BAArLa/yV6wYsyAieTp85ExHNB5MZA/zU8sVUVegSnGH5xGzOhi/JQmBPk7+XyZ8
XrS3D8iWjrgIBtl6VfrfFC1Nd8bSClGyzlDUOD/inGTkUOu1A8cdjc6cuJ8obYIH
D/QhlweqjlW/BVCfQUP6KRoHVHjcAfv7ppWhTPuDtLRL9VC99V5dFvBx76ePnMVK
o0MYh9/jin2EzIw0Q0bq5oAFNFom4sGqlZqNJHwEdxMGh6c8/Gq64fkh2Do2XB6v
e/M4wQLV095peKTsr4N0nbcdajwG+CktGGgjYx7CYJtftShEuw3lsZujNFszBrBK
SWFYzyjkFZYjae7MfbeRfYy4AkCAu/FF952yiGL68SK4UUTES0HW9MVUPEZILGzJ
x7dnw7nvCeJ9clFoQGZ6FrArfJK7lquYiAYlCYE7DrEiwqXOs6KOq0LRQ6laNdso
pVTC4fRcFbhNcNJTNkPmYpMCjRdrmcOHyn6DwwKWEGO7ScZWB9sFYduM8dz87IPO
TxwiCnINcc2VOWA5dtHr0QAo77IXbPeRgW81QM3Eh+pe3lI7bvA187oVKQuKbYjV
IkaXqGWbkQ5w4u1jw8oIlum4lcb1eh+gKS5v1bYh2jI+Uf6YPFhaCb416eJmQeB6
vDFxhoTI4Pc8dyJzhTYUYwGV0gRrKW2mqYpUIMkMLeqBDnlV+oHWLQMxaO3aZ4ku
J+6/S2VtNpYvu0YPPuQLqC0Zdha4twoORe8Ds4ySG4cbU+N/mTeBxhmjU6+UuHhH
sHrrBsavDpFRXZQjgeEPtASF3Fb+CfNAlj6W7t+gwOK52BUX6PSX/b8rD1L7PmsU
zGbz2RUFmwlxpgtkn8U1o05bt0Hd1N2834BNVzDHbl35yxP63H4lOrY5L2DPTi/z
ci8FrXr5jWfSa7uw41ob5LGWly9jOh+9BScTNR/wHc2IuZIVBGYtkUCWcDWz9DDL
LSFKuOxINBAdjq7sTVemsVFy3kTKifzWOFfmdGJjUIPf+XZVzU6+bHl2qFozmGcK
F3w+FiC7HqTkarujN0JtfZ/0d5XYB5ltIMOHSSykSFgfezfFmnUylWfCxgCHv8dT
M8TI52hhDT9a5zoZDUIOTn35JpjCrf3tnu0wh3clPg998s20a1GbcCoqJ3ulZWdc
H+Jxo+MAHP7Fkpomvwy+wjg7C+FEdCQXAl9lDXdUKIUBU7xhCtpRRxGvLVbBzXbF
Ss1Bndfojf16CB0yUMNvcsgMZITNcd7CgQTVL8MFuG8HtxvokMjUGBe9K28p2Uxz
OXCygvu7bmnqJ6Q/ndB+Uex83YngCzzoKsbHGgJEy0bb87kLVr8tOVmYxXt6ykR8
Y9qhC8FVHW6P/j0gCIOOkkxjYfZUoSJcrpAQgHapCCxIecj+yChKO5+yCoYlmgkb
H1bF9lnWYkPnsUZyfFLSd48D9YyZ/xAwHXG56VdzE3tWKiczS/wtC3BL+QWNYuV8
LSISlfYoy4GNUtICVbajkgSC94Iw7jjcIqHudXfiTo3GFLBRWctQmXdbah8crN7I
ZAbYEVDP063jhYzQDeVTKTF69kbaQZ4vWLrTsw37GSswWiwoSNOun1bFW/li2cVI
5gZd6Qeci+TCWAOFaVKEFC6k4ycQjODxt4jTgqywoJ7C6jX0ff2c1sAAvvwmZEV5
i952Yhrq56SDenYXMHeDM3MCoTLU1jV7wXWE8tCIKqbzPqjwnJ8K6GMSIwvYbGaW
OEYnuQf5Zc1+WENyePOeaCm4e6cIQdXPeBc0KOUy88ROU13/zGUP3ekX8JmKwrsC
P7gSgMJf4MasBMF7JWtsph+IIR3+RspDN5kPRNNYAjBgDZw2fa9V4ZB7flZXJEhS
NXACnK3q6WSilSQ2kDhV/XeKXSmfkjSjfBU/GvAKMH5/lpxc80G01x8JvxhOPIFw
0xntkJ7gg207mk+F+/9kgXEUHlTVDs1za+63tqzSVPerG0P8qe1euG/8ktTCRRdA
I8uS98iIcoqeRVifTU/ztIaD67Y3lQhnmSs519BzyvkgAj693Mt/ag7+uixH0CT6
0ayfJSZAa7lKyoyHJQkyuURLxVZp116r2Z3b6fVwaJzGEqnmIjiBZxjBTynkhmjc
7fxzH/ta31XB8QBYOLO95VTdDDiuWta5RoMWEHjT/751FGQpAjlCLxt5ZMxpgYhj
17glDE7uivmA03s7O/xCxpcjaOEro6dFFRy7qxPRu/dyCUekHHpd5y2m9tA0f4/Z
R65Jfjr1G5c1gmx6LDxOoIUerb5L4MrdpuVwp3iRtA/kOrtehpqM1XuPW4XCf4sb
c5aNPvU4Rb8I+ixqwbWyddVVQG+ChTX3CKRAmqcaYBxdPYnZlbhOP+47OJ/wApId
ZUsj+RGrsiLLB+Ab+ke8CWueEX9DC1c4f5lr//4pmsyj/e1bp9nmYqyScELQ1bdt
sknXiFLGwdyoKp1Dunlrf5hjR10kFZM8v9KoGMWOmHPfCTB37UJDXazNjmMOOoVf
DVWvMjb6QOgnSW9MLb/4rPlD7r/xKx78F/0tUut/SZ3o4hByDXRv2K+rs70Sps5J
BzCQnm/lySfp1GKHd02peNyAluoCv1kST0gJOmmffzVmSvVF4fi6g96LA140ghaH
E8k8OHYGakaWBBN0I6XOE7/VS7NPpN43j+g51ctdehWSvyZM9S25i0mHThKyYAhW
UpWnigokAQYoubK+Rug6IpZqlYB5DfbCP7b4dPzuDYh/rgLADB87XEocZ0Qr6y03
PlwkzZttOTDgdMZT4yoOFfrodKwqgVgDheAV1c9S26RdkrO0VsxelpEUmqJRioG1
nVapCSnB2j7CiHz+4OivPeSzahBt5Y2mzhx+guzQGRVPXvLE5BbGXotACMmonR5d
V8tQViID49YWMgL9mhNez0KZM87POQE3nypIUrIGnfZckCDOP/JZ9rNITsTAdWrr
dzXoFWhU2frwQQTBQVTiy66w0COQku6ChcWzpV66jciNwOUfzLrmvAg0qEIzfGpm
ucXqaG+Cce97c1fVwxp7G+INZ+vmL2rW0aAJgcAFQc8SxzLb9aqS6lcEzQlGNYR6
T5/sNELzNxyiXcF9LNvxj8QAIL4wLruMiFsdAzWStTWEhc8lbSWpI8x8IbOW/4Rd
nvNJvRVWhpGf9TVfOnyFKoyUlBPXke/DWlzlok5Ztqzi6w7n3d3dRnmTCtWaxyux
H49fdDqmFOI0yoOKNwu7wq1Hrfpzauy3n/pr4oQMyRW5siTLzNNmhWaU/e89khzz
ER0IIahOLogdLjjSw3MFPiduXx8XTwHqYJZ8KJwDHJu+o7LDswREHzLE3Xi3W4m8
6sQHZUts0JpxJNA9slaMnYSAZoqOicblTFr4jNF2EIGEnNYz1eSMrc4bHwMDaHrY
G3HnIdpxQSDzrff8uzY0OTJw6RPSYAHwz5YKH6cksx7sf2l418Yh+n5xaJttVvbL
9vrnNVKmyKmE4WPfZN496Hoj02cEVzdhfOzZsSMWGq48CeYTbQ8kggPmaR4ODkNi
HqmlbbTT4GiHuuke1gRmtKd02+mCUvaPfOX7gme9NQwAnevya8oqj0r2GFSLZY8q
cCyVUMa80P9z2kS63/iFdvYjk2tT/dKWgzdcX0QWsp+c94k5TDiKU2CxODZOSbO7
ChYJzR6VGHDKut6DdfHlNOa/meUa8RnkeEpsbfQ7vXWSRtgVPDqWDJTvqFtckk5y
5GCxXCmN9XI0LVEFduzk8DNjw+nGxs1fVva26AaIMSlVnd0bUXJT4dEI2FnAuIbt
vnHhQ9HKQBcQYiWByG8Fa5oj+xQL9LJcIrLW17pkE1V8N85FU18ByAM7reuCGPuQ
Mmu96Kh/w2ThyMYCIUUu7slMSAtHGyok1BN2IrUwX5g5kO9kfR5ikOspSw+JC5C+
q7TD96xtHETUWadQ7X6165oQVbs74VeHcxOZaez4tlW8mI3we1dl4R0V9pP2e9s7
xVxmjuV9phuPXpHTbl2zheCuo9wFFFVtWbf9ziy9SFA7eJBj1Tx5q34MsoCPcakr
4Nqp5Z5EIT5Axsl89dvuXqrMKgkRssFsA6IAb6EJIRG28tjcd674MSL1XOhBD+Nh
IE2ovl2u8HMNdxyWBNUSpCsK5j9cL1loqBICIZRxzx9pKGePXndOV8W3AcySvcY1
PzY10oCBVOy6G5u54L/vkjd/nX3lA8Ypin+P8+Mvn8CV16kZPmKi+D6DmukvvLAm
WoaJsHx25SsSj9fkr2NHijEeullQu0G8nYNeYIDHxMHwEPk5o11AkMYUaJijKplK
MX8Ggrpaqs41TSD7/L79MydS9bX05vFVsTDuwkdfZ1M1crCkREjmWL+bo+gHLHiQ
WKzUmithrX0zdXcyKDf+0bo3JXEpGrv1XQhQ7AUxYMAAdc3AjgQqtdBxcObMdFUi
gR1rzJOBjzml0iRciYZk8YEjtMo9AnJiwQ+vq+KzE3oyhSjBKbb+cQxezueZlc/j
uCxrjXyMFnxeGlmQl1dZ+l83J4sylld0BhD92H3ASYOWvg2xol2k4FyEBatx9utD
fvYRb/aTy7m9sTSGKbPDbmmWuN3Mi1RKd79mSQKIsKj7UcqV8SXpvA41IfAoIXGU
+c3IHgYEqNHn+Bw13GhavI8mTxR5FW9ot/MkXYxkWwaZSmDQTCztsIqkpylvJBLk
eZK2/Syvoi5oIn6XGIfwdyADCb7CjqbCH4K6eU8jWnIDu4mRPp3x8h3uweDoJ1ZQ
maD8RZN7kriAMxIdzcmH+ZtvdZnLsbKmH/Ti+VrvLKDEsrusGl5w92ZtceOWhqdG
/SGQUMA/53m+Wa7hnwDzXs7sPFdOEzEeuDjtEhDxv2TLLLu/N8xvy74z43UDlXfn
35hA5Mnty3ISNv670jsDVJQdsFq9u2zR6YySitOuUapdbFDpjSCztBJdF21v+7+M
N2X0/pME3Gb/ND+TWXLGFku+Y2BOAWMQ2znNOmhZljDerd8SiwZi6zPA6Q5HU5rD
qXQIeMnQKhaj5Rm5ta0wOg2tZYaqUIBvMw9nszQX616fP5vNdLguNpgUZxy2jkhm
06k3OBpWEdXUpMhQqjzUCDZx9QA+lgG1H2wIf1SgQ1PRYDe45PfgMq4Zpdixbcng
jSn7VAYDW4lrvdyL1Zh9VtMyAyJRJtS/YXmDpxBHrKx+Uc45H8pixFyOPnsSIdAe
Pq085Z1iXpCV3VpwIpVeGqmADQz2r6/h2BbQcnozUTdAo56WHAaqbsnWUdRb+8nw
GgmscPbI2lqQ5Dxp/cv5PxuHuuKU0qK/Af7NAbF2EwHUr5snk3ol7GoX4n/xVGFF
eXtroKCsg6rCAWX5Ooet4qB8Z748L1zozwDFfZ4DFhKawrAcqnNbhl45Ka+W8V1p
HVsxUPGRyJdiMnUS68VJIAvdTo/FpqhCIl7hGsX7PeGt0Rb5z49K0lKpBPH5r1rY
Nju7yBiLmBOCtjjfyw+0QS2bt0d4PnZllF7TwOcBwbzMAPzFcZu/b1mCPzWU5YEZ
BAILWWatIRzE4E8JUhBf+imbF1rPo6m2i4EbdQ0R6MCVE7EKU1Fu6ptIrcnclNAu
xgaJeQe7ZQS55HfnCp27bkNJ8HxpWSJxmAbrO6M/OCBEkDgjwc6cTtvA0Cv0M6xg
lwXSvg3q1USeoo4Mvd/CAw2tUW9DeFAJM1A6il6Cf1vquY71H4vakGnEEbdxd2Ld
NiSEgrxIyYh48H+T3gsU6/yUQtzZ+rDxY7XUZEKiicXsbJ4YZrWUO7PwIIQ+qyLI
wzg0xx9/sUTMa0inZOUUW5rDkzF9TcLpa6Zlt/yVTwOOv+YwTzU0z8RcYypTpzYW
6mxcFsFi50ePsvDCEc/3NIZ5wxRJ2hWdo97/AXZqo3tI+ZZ9YBan9/ag3h87SyMd
apC59FXgfZO+JCDtPg9ygRLksSiADJ0Ij6rl2B51gZtgr3w7/KjuZA8mbHe+uUe6
N1NB32+1eB1JxB01/+L8GyJXNFsb/lWEAFgVIuJzDnkzV+dft4fjo1EN0hy00D/r
S+H3AD6ut8oFy/m42tF+LgFWjt1SL+/4gDwR+N7n55FgJrtxxdSNgNjtfCVl4qa0
Pt2JxlsA445xv3DAWavqixmtdwPxyvp6j/Ml6K9xDWIQ730/M8Ey1314u8mZMmDW
NA5P6ek+XbPYMSNPYucUATnpGj2QJOX19Gs9K2E6cktx0A5TckY/VhW/r5NcPJsn
T5nEm6wgPcNt6cQbHndM1pVIlXzTmIzoYU5QrOKz5XnNGKnNzsf2ctqvKzqaetP2
0cH0svkVInJrLeuShQfEUikpFV5Ik5SH6LmWIduDTzYeaewdq/xRBhE8smBVzziT
/E803RFC2RM4dxXHeC9klSIccYoZ+tStz48m7VsxdqIO2yZ3D2NwfHL28+NKuNP8
jOhVEBxJTTPorXBun8BVknr70VX2hhkLhRDvW/yUWYexN8Gvagd7qhgjfMk9drku
flwwFx+FqVQ8JnimPpBiRSti3EY+HOkgse3zW6+W6dH/mb5t9hz0SHKmOFHvOAt1
CMXiP3rk8lonuF7KPApPEW8u6cVQsddh8MobBBYKcCybsxT/FNCnSZySYeT+G8J5
tAihpFiIUTKJAZ/nH7iCKoMGzMJK5qPv6LqfXTbJUDW0R53W79Zej7eWalHAXMNT
Yso9JwcucYv+3tKg+BDq3QvyniBUm81+eJurjMghCL4IshO2INQQpYNWy4Dxgnqs
/9R8s0GRygGE2ekuCz0Ga6co2cSy8NdJA7YNVJdlpey3AWipJ8mpskqv1OK6tQ9g
7p1CLw8fzVOEcXaUgk/kA8zJO1+n6dkoRFvdi4n+SNzHKDrodhbTg2W/NJGAe/mj
C187m3pel+McljjWWMIL740vSxI5NblYNZNIaJtKt9AQjOj9Kn6zStvybGHbPOMS
YiYmkdyNrndqmSYOg0je2oMLvvMR6rNa5xwZYVjvvknHGv8OEDsvPehWGvB7O3XZ
lUlcFTdkm0/SQDyJnANKqfTgObgjMCKn+VGCmXETGjtZ+L6CgBFGXwQL5FNpBMYF
HS6YoptoD8PxrF7+p1dWMMT0vFy+rP/oHii0YJMecD+7qGt5GGtYqV0FOxWA2+/l
RYbpg7EA11YDex4oP+vz9BxpSFC+89AVXREcQH6qDCASj+F8jfzgvAQUdo2B8Dss
ckX/yDjz260zzfwtY1a6R3F1GYhy/1nfdsDBQULBKMTN//ui/ko6/UqgCdAdSBM4
C08gm0NR9JIY8/Cpo/sy75VPPeADR8g1gGJHOYjmVkAh0jDnsv18tvJxyMPN1YDb
410PD7IYb4hfbhtl8i2DegCmZxBsJlkONq9SgsVRRn8up0bwCwrt9Q602WtkqHa0
COIEjEkehN0qzlYGeJ6ze+DgjznCZbGgcsEf7lHnNczbE9twnFGYT4wIdYM5w2HZ
b1ZgrYjnIU6ELy1DBgneDl60S6MxKi+KxpEJI3KTDZ4qeRJK3HiEf6CQXRTOdRet
6NDihVmgSOu9nguDSRbN7uml7KYiPJUPsv7f4MLGW1hWVp/Z+8dC9nMRHZ1ql9WZ
nFaVY26FCvy8bK8xcBhO4BuEMoqGvVW4LjRtdopFEUzY1agd/HEhXtXL02KpkzsW
84kStJ62g3LAmUQrJb2aEhanxIJh2wWS1Mu9d9niEAjQl0nTtfUvYWuLPuXWYp0J
2J2gs28ZNZPY5dsGzsoegqvF/yza8Y223VUY+omJ4jxhVFaWa80xHT6V9oKX0kmu
/5+ZN3MfRXXPWLPCfcjXJAnprUB0K9aNP2JXXTlL8pdieTgVgnXDuG2CMW76AO9S
uYPs4faPv3J6Gpb5rpbJkQFUk5IzETzld0wFssOhvcMl+U3yxdaAfzFaCpKdvJio
kHVj8Qux+wnBFNcqn4OYMzR6DVuXQtm/1cmFIg9NDicveJSs9pPmcMjhRzlruTxU
KtIYBC+09Jfip3Ec7Znvo/EEfsNnn/Nxv+7+6ATHQL7UalK6IiGkNHNbplWhROLi
wS+FAcBtT89ZDvInnkeiiNJDRuySyeOy+EBQiFT406JcwnLeiZHgfRtAxEuHIgaM
M4dgo48X0X4ikGJ+d0qriCmV5/7qUtTLLJ8XjBhTaXzPC3hcMGPmNCl3hsjg0vFM
Sz/0Ye9dKtPr9gFLEHkHqdyzJ9D3ut36o221HB5j7oJ9jxbz16sZk9aaNj4AWmE2
7uK95dG5X1bQO5c/F/87y2BvVZDYrgOB3kpArodw8u03jTv2DJu83MMY8Y6XCNew
UnW2a+ncKCafHk4O4NYjA09j77af2dxYIkNoQH/Y7vFXxQiweb4qzNtfgfRpMFq+
tVrsaz4wXsYbYpTjIEB5KFc4AOLvbvODrU/uUeJiY/KC6nVE6ai0cEAjiJ7Bd5Hq
HL4VIh8lf/9m9mw1VDUHKK237kyFSWt9fhokDsuJfzQYTLUJq5Iq71k5F7WYcfdS
2TCj8b5FiUwLz86WQ6Arkf4mxqMGWw6+1115fo9RTkZsMyKEVLLZzMOJSTWZBn2j
/5T5ABqUSOlyGjIGWY282gqxDf+FyxAQdXjfkunMcY69sPv+xVKZojY1sQDJi4Xr
4pkgGLQ2uZMHOiW4dp4qKPXmaQoyC2mM7ZiZpKO2ko3zOX3qXxQo14GtVW6f108W
DWJFO5dSLL4Fgqb64S8AHAZxGni9ePjPyzvh4ALZ+HjqFjPLLPhN+xGhQulb2iJZ
OzF94OHCbhNAQagltNdJMHtZ7+zHFeI16+8owQQ90ntiwtDOYqkPlP/9zLb/UyCO
ZA+mDymbevRhzr0BCEFBHyGxoreeoD7vBrvAoxGgoC9PITTudpXNQqcXFAlBCrrk
YZ/UfPuM3ZepZA1cJmFGBAP6Poq9TwkRHANnkaxeWWvflIEAEunZAOaWFKPnbooS
JNXw3cDb/lWK50vMLw9Yrwn24v8jYkYjY7GQxuq9dmn4vWhxzvson2ba1gZWUAR4
yiftAVI1H/SEp4+3w0wk+bTE3+LdhQO1/c986iznKnKAzzXRS+HAcHxmTgDSJVl/
3O9nQT4z9SL5EUbbu2NT4oVGGO+c5XKOtOR6D8ChKv6e0t43KTDTcbPoWhWicEg9
zUC8XSnNOlaulOkkMIZJC/fv2oVCY4Jj/QnDLiwxLeeIEk5ZIwimP5ItY6QX+QXo
IubBox0CiKg27poiIjIXHgC0xMV+wNM1ezY2i3d8NG8FNDxX8ywTl5sf/VEcepa1
GQxyQPTqGobEMhFqq3zeD1URACP4xJPXJzs7LzgP7qDAuSnHj05xyS1xBhxLyHX+
N7yu25Fgbv3nCsVLHt+peHtDthIfxJ8K8zlqj1L8RJk0wrxGXmXDhZs1/mFf7EiB
+EKYIOSbb61PwKnJRMc4Qr8xWIb5Z8oap657BLTXfYBycAjdFsCZfNHBbu9zoJVp
izg6Ui86aIow2cIazwY/T+4yyJv5v6kfBVLnF20Hfb2TinkTLXuYjeJ04TVFRfxS
b9W6w1g4RJ/vg29aVysDOEM+sW0c5JN/iiKWqQ9+w/x+dIhAcw5XWImloPXvhG5e
q+X8p8ztxqKSGDP0xuLOAtawyZyw72MXO6JmUw5q9m+wK3JG48lVSSGbSUZjkJsk
GtRjW0zVvGlMZ7u8nNOLI+oxe3HX19QXhmFSbklsRuqKyl/4+ZFHH7uUNluUWKm1
aH5oL7COSU9nLR3LbJZ6gr6F3LVRsxoCGfhlMjrrLr25etfqFdPPP7sv2RXdu3b4
19WwGMqCQ2P8pYCo2r8rWWsB/yHs68ZuzmKP4T97GKV+xYJhEU7KbjQiStLbaqma
f+0ocEIGT5MINmxMb/ZMN9Sbi9r/CetC6MEYPIOoQ9m0tArZbgPGmj0ML2DJHbsn
SGn09wTeZKx3xrbfqAu3BsdTr1nwX4GQH55CS1mxIXtHL6t4IzZGE2Q9qoHnEfgS
sas62djI0ERI96T/0JNVbzj8sT1JgcK8zfZ+OdNRaiq7ISMtQhsSHqBvG/3nKvKM
koY0D7DQTWSGUaBfcMpISZpkhvaxhnbAbHtX5PKEFElyYEaGfBElanhEjCFWshCZ
Xzu9PJEAB1RezTDdQX2rInIFuyeOzhyRYEbtPd5Qmd46ZMxao8GeL8eujW5okkRr
pGuSMGpjdnVynd2MAQ553bni1BMeR6FZWs00FLm8EG/GUEW/xTvvW/VQ6ehVQ5+z
lll/UA5+khZfqCUk06bNM6P9uqKW8Y9qQBGVY64OFgjBf+v41loWrk51/lQf/MgC
6lHXL4P5TY487b9ZS7C+mt83fQIASqCF48ilBojZ90pcrpVxlBmBk8wcHgKCTQ0L
sMbtYKIQOkfgwqS+RYn455FHuED+EBXnCqBPkArlagiS7Xva1oZTwhRDK8KJIz90
2o1WnAX9z05OOyXPWyRy4fhgVI95acg7U0FH/hM8dG0ND3ZRWTuSJljU6vwopB++
6GIEHCm/B97WuAgGpGlmR1BaG9sMC8TbLsMReJwBNYgRAFjyyTne4jD7jX7n1RI8
fBsi53WXORVVpQfDaCegwl68+MlXk4w6z3y4GmPL3LYIavydahFq1of/ccuJ3jXb
saHqu31ff3CNoqMviCloM8ZnExxtUlm38GX+RKVWFIBEGFVwN/b/oaT3i34bADG4
XyatzU9gtZLS/wA5moxSU66tBuzazYRdc5fY/W/fxFvcIPGuKysiZr0hPs8zVxVN
1vqdHjRNo7YLpGphjKWOc5v1XemRzJFCsnWsk6TLn3ohlA4l6LDp1d2fpXkrxpBG
z1o6zPvrgjBs3h8ikM9Dr1Kl2+RnGnxKj/G43pecJIOlKHK5gKqW3+XWQSypwSCG
lNYnI/EIufbfBPDxfnlQtC0u7W8YCtQaYyguYo+oPFdl+gvp13yY7plNusHE7ssZ
dmhc8J6PUB48BBv0hI5bAAHqh99hYcgyOhCYJxDrW/b7GvTRV8nBCOsy1GyQff03
qfZx1Wuvp8HJGV5mycDN3/CQnZCr1xT0aym7WdTdAvqddZlQn7Rs5Id0oVfJxvHA
IINaPFUklz5jVKkUkOXmxBvRePIXe4xYmJC7RO34TwBtca9GK2l8cxWTZmPJT+94
Q2Y4z5l5+22feHrREXotOEqmh/3XRh1JypuYi/ZHPW+JpjL7MMfw6HRfz9gkk2Dl
vwaSHKc6Ay8RU2FyOB81V4BYYJRr7qAjO+3dOb6s/9CQrGr3bc2DFnYV7NJMI3D9
+Ob364Cn06vLGUM0J8frVzuLrivbgeFfW4e6z9iUt0EtvKdULqaKUnhhUb1dpYS/
1fRQMIzEqsIF6Rmkd4BUEH3jM16xiVVGriRSfA+VxkJ4iWd37Gj+zh/xVSQJKXzh
uC0tXE+eYYvPtlnm9QGMCIEI9po0Ddf90V2ZARCO1/7dZlafgllYDslej0a1+Wle
5u69ZnHKZBfFcu1AYQ3iHJEqciDoalAZRo9hmIW0OsVH+Bm1ZUWwAyRVy5YhBVmf
pVYUN/kXVMzHpMtrrcYYoQU6mNudNHb4vBNDdgInDafXuPtlKbWZ0iMYIMwEMN5u
fDaAZ7on6sd9Cfrdta/8hrGux90hW4cdXRUbygYdsUqdCvssPEbHh+xZcgWW3vLe
lm5LTqeR+nU0Qesp49mv/IHakscEtulLcqCl1Bvd3JE33Cp+8UJRP6wxIqE0d0Yx
DLRcSvCw3BMtIoLYB6ELhq4dVu4l0Jm/O8L6pwbC72QeBmcTBPPbtZlS4uswrH81
MO42u9pMpktbsRHrCjqJz2FnxVLUmE09nWKZ36wm6MUUsmngy7vIjn5iYcJ+d3Pn
NeG7Mn7SFvpCUJTzcaY3Ef9QEq7vGPrO9t+Cx0bBBxhOcyG0NLm//3/StVHsFFI/
c3xTGjzadVd3QPxP8uLDc0E8BumF1OyMFRna+x4Ee75Fq2cmX+j8XFdv4zjrBY01
n5ebj8as4bKuZu4Rah5fAodlBgeooiUMxUrVcpTl/yRLaxK8slxmNnO7q6YyIzwN
EQgFk8A1RgMkD+H7auq3CKm+IThXNcpT4zZCPSR5J5KBRAvy/aBVWOL5PqP7YRDf
7/W5t1z8ihk8f0qrlkkMqkXRdh2aloIs+m9LhSyk5W0IrJv9E3c8fgM76p6HYVdC
5GOJ+CqUlI+dr2SvCp/8ggZ97hCy82qGWsGrs/27S+Htf6/nLMfydmqQEzVMZIPq
E/EC0+v8J96Wbhc/LO6bjSxvqlRxpkvFUZ3gPwwHs0o1GEzXPTkwrlpSplkw/zXL
ry7NywfBUUlDnvTIRVnFKI2n5s0qd1LokL/M7Baxti3U2oJwDU5zkmZlCXr66qEl
Y/hAYpb0uaTQF3jNclodtNW4SpceOP4Gh8weZVfT4mfCwfQL99K0mQxhOpWFBli7
cfULCUZHZpa0mD4QW+kEC3D9hKSAP48gNL3fdU3uauunJmBq5kExPH5MGxkhhQ/k
OzZTPli1Xx68tUhCdujiTx01F5Fx62kA7qROEPrMmTtQhQF7+9Q7gdJhgzGWMSdc
XFBGysbOughtUES7gsPv0ARnPe+4AVwRj8nqB0ortVzCO7toK3gMQ/tZYbRcQbqX
r9Ob4tU7QkQ7MLOsDH/R3z0NFasnrlyLDFb9AE9L+XjdgfKAUlMhQ6lZVWsfxevB
TwAaUgBerGyiKSbzKudoIwcMYOjM4CxGwmbjTQ6tgTJH60vnBjrcgJBAEM/tifyi
MGBw8udZYyfTvAxddC1iVJaRS0NlRJuzCzFN3NcPlAFkicx0fqlkGJu35yaAr5I9
XpmQb1Yo5Pj1GwrAvaZrS1c4Wo9gI+Ybh7h4kTVKa3rc/cxtKCn+7FlHVO3MB88H
cxpMk4sC1r0T/znYqxQHjHWMsFQ3vt4GSb3eDbZdkV8lVPS23tMCcfOpR6StGaeN
s1+2oFF2ToyALe/sQ6ez/jMnv0URkpOg/MdyuHgSXm/mMuAa9IaTGqp7cRGTC53X
QzrYyT11fsoyQ1p5++J3RHikTqYB0W1+Zea4TuUGADYeOFx/Kf+LwXySZCHBmP7I
UPU/O5OkKcNzlkVwv55rQF1R+sQgEYX3h1WqXqx7bJpPkyevfTXQJ08hmVbtavwg
eynzSpCN8NTHSJTH9KiHXrvtd6309y+gnwsItF6EpcDYJpGhN3YqUKBnNkbssYUf
7TvgEnU196bPQqZZRTni8ppDKcqjKsmqK+UDulzUR3zxFr5bTSbt/tT2B4cogAv2
UgANymm2WRHiBq4TheJBeDOB9w/JDbRnnyXbjkP0c8V6985WQsPegNDUQNlR+l3N
L5g0mTS6cFLpg4DiwArzESUKfTldp32NTYge9w2LOwKJPbc7+TodT1C6worXzclW
kH34ZAdO3hQOiBQ1vFoqZNZACUIg0DvGdgK0AgjYD8qqyPd/99K3SIxMTrqyPriq
H5UQ6B10vIDnLUUesnpOxHD+D3hUjD8A6WRxFVoxs+vqL6b4UU7JNgMNLOHVj+31
xJJKSBMbn5sIjA9TkexFXQ5tIQ/6pOsA4rpf7/0IzDVLBxqrzyyoRHOrdYp/BlsD
CgqGSxBmfSLiaiJJNap2v91tnTo7WTQn3JdofflrMihG1aUmLT11YmqkfTNSUdRZ
c00UIktC5gBU9Cm7HgiYVsUbFKGZ/xRIXS+CBzPU+TxymSeSVA2VPInwIUcM6IUb
nS80DzwlPjoJ6DQTzBZ1Ee+jmmAQxyWI9NNg7r0Ue8hv07L+thsIxY07cN8Fgwfw
Z6TqdgczczS7D/l1HBeJ0Fl6aiZkYUH61Kh0P/l5KH2Ksb+IjtTPJ5NVfbAHpoDF
4S1GPa/cgL6vYnLVi8Mol8sETIdpr9cDgbjtmdFlMoQwRLee3bQQKlU9Ig3lRvlt
4qcJlLJ9xehMxrsneT1JOGA59xcXFJwFk0wmAfXeclFvNOUqPOZBERZGVEoBP+vm
g8si5dHZ/qaAMfNf9zhsiE/0+nM7XYJi8aTLuTjITVuB/RudtDl7LFvTU+LzGIHK
q2PvLsTkOv4P6O2K6vSgbGNygbWersf2v94IuDxm6ySvQM68goVY2Q1I1WSWV79y
u8HtPydz5yBN78fqWbZ62eMUiFBrrzfn6KwA6ioP0ALDD1JzVOshqyHEnivMBGkG
rE+yrDvdQe9cGEgxsi16/jNcXYy628CpthrOtyCRtSoYfpakItR5nE3xYpIal3lD
LN/Pw0WZig2p+YXxUQeSa4xbkB3ce4RO6LPWd009rFgMp95uHOdVdr22zHV21OwX
DaZMRnDWUGhvQGyWypvH06GieoTZm/d4lQ0gjj9NxS5rgrQ/V9w4fTJGdmS4MWcr
/90498gtcwqxsGxpS07VWBm5oARv3PR17WovS4zpZbas1KMjvpHteEuz/eHx1/FP
iG1/GRigWd4Pn2sMfv3snTlT9SilGh5xsYKxo1T8sSeh7v5kQG9GqIQph3WRlnLv
jvotDkSFhrLyT4SQRDAAsi2cDHjGRfn/yMy7TT6xfPHXWAvTlRCGL6y4pCoLCnpA
HwpmUwMgQLNl3In7MtixQz2wwejub88ORVZRItAsrCRA3FAGngrQnQlq5tC642pq
+sS7n5hvfyrM75VefSxkWjfPQZpWsWn04i3gb+UOkW97Tyyru5FArtd04LwE5b6z
Re+MfK58HlHhmC/N2XLrbodMYcjV7xgevi3E35NXrP23gIvWw67FcQEdu6Q5maXc
QlWrVlFYVDVv1N5xpIJx2+p1TLp6S/QNL90uOp+pbIK0dpNZvf+UMWzRu7ts4K/O
puNNHW+hXzsTw1xXHxdA71rm5PWfzObjf61aI2Y+YmKxn9hgQiqbZ8fp9ZfxKDEt
Q1CULwubiE/fBi097wBf3u/K4TVabVBiu4SpPdrr0lo9Dbi+BpayWBV2K5Pzz7p3
88gtLCOGoAsHZwUSLgTBcr6jNyQXGcUUc7kNdYvVGXZfV0a47spV/W2rhv+qsajT
+1Hvoir7ltUwvqz3sr46cwqzgLH7hLC6IGJVDn2eO1r6w1A3FF26rM7G2g0c1ZOr
xBSwKlseUbbIdq6EiF339TGnhqsfBfRR0HHgrzifzW4AZZfxEkdZsCHePAaZiY1/
EwXqnlTh4VsRpZpgmLiG+/UY9UiLSRWqU95NJOJYc2mChG5Ybo3dFSzR5B5ZdOZC
YwT9ggouGDNGVMQDFIQ9kLAaRHGeOz8Ar4fGtZxQnskwzeFd3A3Y4F/3ZlPB2sva
GLX30Z5CY7pJy9y9IqQOIJy/Wh0j4wtvlHfuFO0214wUpEHVBU0tPFpBOBn9m8fI
iFAIdp5eZsgqEl11co5IsnkgJF8Ozejs0PMbtV1WQJYjB3k7/TxYybTIjhofW4BW
COGK1fh5D1mTRPFJ4kZvcY8oxo5qwzp1/4KYbrbVHjAkLqlLopM326/s8hIRqaYC
zuuzrC2E0weVVRpo8RmNfNhAtPlmJzMtF72uVmPKLfa35l1NnNPi5zdHqT1VpqBM
EfQeeyZPSyAzUyUOUna98aJBM1yPVcNkzbPG6EfxNeThz8jzm9pvcJjdHy6zbl6v
Zex2PSiiO/6qcw20nwVNhWBU+ryMGgerNPcuV1RkbXxRFmrdI6m/bNi4mskM7ZWG
EooX8ESDlGbdiYl97bdM5O3QxF9FMBJOE3Mej4FPcA/qpgWhmJ4tGsMTbW44AHRR
QVcWTbMcR+wbppsjCag8VkebWEeJCoUJlr5Cv4ErjcBPdFFjTPdW1gtgjgko+JGU
wq5FAfxo7LHDhOpqRb/dv8nBwEplWBxjm5zR131jYRfA9TF8HFMgkEsb4d/00Mdb
arIIJZmoZUxepISSG/x9PfpwCwexbAQ3qqKQSJeTIa1gnsSKAZKXkDawNunvs/5c
mCGxDzF3WI2BzKKIhmqdo7g8PIbzkad/P0Vy9UpYAeZIiTIjOXvRUaz+sHDn+fXF
yAa7R/ETpyDlyJyJeCgX0KTYY1/s3NW5rvLzw1k+j4fP7sWIKSclKgG7iDZwsaI2
duQH0MMXxDKOPxujGrKxBbwvzAAGFgkqnIegDgWn1QWkaa1VWJxXirNxhijoeoZ1
gIG8NJ0AoPmYHuLbdVJM6B50LWKG3MjNzfBfeRbyymewIBHC/ZgHt0FFO8e9KGWM
6nw1ceh7jwDVPcPyZbH/H4j6DfVipLPHdsW7d0QQKYgvNRwh0cFlpZFLNcDlf0Em
MPCBSXtHwaT3BI6RbsXEYnnEz4WfKdQLyl1dd78Xeoo3lfJE39sURx87t7wLudQ5
u4O1T8bgvp9fcDQaWBkhACEYDx4vS9sXdDX99EpkDXTiFzoeOi1/RHIe+mgQasJe
ukaqB9YL3ptJR+ZcnSS2jeFvd7AzYcvUdcC0C1120psegWbr6aGOeX0XEGsZl/6s
RSS7HORjlUh/gJrD8UiwEw8JWjwbVLu4lLYNAjLe7CFCutnb5G86mNNXbWhAJ5Pd
fWdOTFbl69UZND0GLb8AArx0iD28I5tD36S5Z5ui3kIQiCfK1LS56v7W9xB2o3lx
ZYCxxsZMIyA28rfqrOftV6cuE7E6w/tU/b/qmuRspzR7Id6mCGYnJaJrSjIvNmdA
SGXZCuCkgEm0bzNBk8mHLsWxXG7/Moc8GM7mTim3btYxnGFz1vtRPlZc5snoyElZ
Ay/GMW3Gfqd7+CLZ1+qlN1vsk9DMe1LPnKprMKLNBaSo2wmFVIWeZIrbwHwnHq25
Af9g34bitfGJJ9a+Vyoy+p1VVFS6lzRaVKeYLBKN13UBWHhvjfqQAanBX3Ggei4o
BxbQaUs6ohHv/beDGMZvhgNAyDwMaCdueaNsEw1WuuQk4q8yRefkbDhCAwNsz1PS
iVdiiq3j5aCW+/hOKpSBOZ5oETY9HeuWMPQUbSEx3ljXt4A86p3ycy7sfN+5bGi0
DZJNaDcofDKEzafAByD1nDuKnCnlzr0lLp+gi6zpivvb8RmOza3omJ8bKsF2x3x0
KBLAyxBNxEi5reKxCMsB4XOsAeVI6JrAGHfR1LJEOXa/ma3IbX8l543Jo/FPib1R
f9n5Lke6gGGtq2V8gawTeELYC8RbdWLonjyOX/SO9+4Z0AnP+9hd4/ufzyBaWVq1
BrwUdn472VVECkJaPpEXinW9Uut/OvjymBFRLOFjbI2So2MqRU2qvSyeNRSsm2lr
7S7hNK0pTm/NFNNPKWfQK94p969D3+7kfGQ2V1mTYMEZRuvlBFi6hKHqthhj3cSE
B6XWcajj2AIx3Cn+DtUwdBMR7xe2xVp+G18U2gxu7ENrEmMrpOtige/ctrTgxUZR
PlxMTMui8+KxZ/pTSxmI4SZwlcXcx/a1z+oG0HKAv59Us1XMPaEzwm7et3Gpb8lB
ZrvuoYhY7wwrDOenus6SlGq69AxY+G9HhWNGV0a+oOWMzk3YmN9613hVqYkY8mFr
1uy74BmtMNnpoIMBy8mzUYpS1w6jNepVCqGn47/20GyLSbmG0nob0SoCzADvywu5
scW+iGzqIWMNX9DlcIJF++DoYteyZcsCuzjv6DfWfA3RDX0HKpyk4WNfrjzwtLM0
Fm1smehiUdTDICZKKTUA9uHnLYM3c6Q7V+aQhPHtt2dMmGdXb5GX19w2cHOP6PdC
UIUDQ79pqQhbEr3Cbs9u9wqLOtdb4NS59IkEBIqVrKw5atTWvmV/tVvXbVuPRVY6
9AnLkD2GAnMeneo7vNaHxSEB1rK+NXHNss3FoyM8xd7dNqEpE4EEThCgLaoB+sEM
jUkhbk4I/4QzDUYqqYmyP/LjrDm1M6QnwTS7TcON/CULDEX2eWWP+W6HsGaYzaxY
bGcDrGEtmO+6VwacCK8Ypvd1HQ+wNUlRwq/7Ao2caKogmH9FXrnn1iDVS1fdxkrk
zkYJAdoq+Ju5RFWv15Y9OWzhLzj0ljTdqCPd78iFfP5DwnQMsP5P67d0m0zAvXU9
b+pyThphv9LoZod5ndSmNOsKA8iQRXa6Lf0M/YXj/YX0QlGoGC9wAofyKjiDJNSN
tDlu0V6N71m7Al9SuUv6noOr05UlD7dDegOSBDgyStwn+hT3zNmtXEaZDWjsLSr2
qfearOuVctorc+wQjIbE/RVP8+Ya6v865H0MDBIuxhhklyg87mnXv47Inhjq7BGs
SFEtxrgW5hICWdNFEsQiZbGLR/RcXIFdCP62ZjtBzW47RVA1DcHuIP+coXlaIAL0
szRTkEm/KUrXyWe/2UlVqraQfz3zuoem2rXqXMN42zie9KY1Ev53bofhMFkqrgE7
X7GCNOtFo1AVOfBGNPX3vdIbx00MMZ9idb4xCr8Pz+kCGhsJGYEMTlqA2tcuvcyY
QMvA7f4uwcCMI15LlRVqnNFR9dp+enHthFsaZL2jzXHbC6Sv0OuQ1PhiJK6lLIlR
DbdbCke0j+Lgos7bOYUpC4Lh4IYoWixtcewA39vNTHdR+ddKAEESWYGrTxP/E5Ja
IudG7tU4lYgYMbiyUKFcls/wtNkr4naLL69/kk0MZ7QVgvvYqiagFrV7+tLYNkrH
92U/SFi0EPer+4wSTG6MyRIwfnPR1uwgOE6G7XkUFq2zt6vlNEWawQokFtsrIx9F
hFL6dA/T8i9vk4PNogT3nwuM3cGmaN966QP5Uu6DuivzoXE9wz3FvspXzk8Oi07c
KF/x90DDEdlAq3b2nnu40Ch2hIF7eOejEq5LLnBL1cbeBegZKUpXbPwmsZCrVCzY
zbonjvVA44eKCXOJe8pYyaQcGSUu13nM1475T/HsJmvH/dXAXrJnoo/ilTNLdgyA
y7zI0ZQRMAWDvXmpwvIUCQFxC1Y4NSO9wWQFnrN5wmAUBd4KftPyJJzqLSXJ/+Bl
j9ntUSaP/HjHvwIIx3opmJeUcx3QPuAclP2P4kyYM36YLm5ijBOZbmiyx1LtcyYg
fZDrpCBcEn2Zzqu8AcIZUPSxBTURkHInl/W5wB32aAO1G+m/F28YwR+KvRc0yDmN
aW9ciLwEYZylzoA5oRPw5ePkqutbsuB6lb1PPl+O2/nsVVi58MzOXjFb+TI5BUV1
+IWgJA6qSoRogPhO63S4zNNidJfqewIeyx/4okTeb6GE0O0UpXdjxdMEL97GXLRS
VXSzRL/Smir5tt650samCl/xZYzsJ1FkdxNB6cFKYKzW6ja2uhUo/tvOikjQV/84
9UvozxHYNH61EOehBxaAgHql8HGCxLdjg3f4M5B1RD4wPt4OVrN9jr/5Vhf72YMv
ASEKZhIhk0NahI+T5QD0uyDlxcH4NkRzWifh2fv8BxfD03YDTWzX4cNjgE4Kzi+H
4n77D0vymnrsoklMlmBssRcd2N++gGs/uRyfrDfOU75Qxmxw92gjtdvpY9pTUQG1
W413orJFQELZWoaPK+s+Qp3jkUVNk477uyq7lWcomIpUaby5t+RP8/STZfbs8h1s
3hZK247Z6bAirVENJ4Zw9JYD4xYvnX0ideTW1bUDnXB8FneRDusSSzV0YAS59++s
AoO9gKr2Fz/VhP3419oKogRr0xxVK1IvD2ANH5P1bCZopzGn5HT+eoWxmgHwUzX4
JTC9slS4FOrczfYTTWEnVMqeFJwvLqyCEZrz8hcjb0HIspE3wUz4Cms2zeiCwHvU
smU9I2qXYNnSp7CHryx7TCrfAKwii7AvSdZWPrrTRiU3PcCJYISMNCpO6DbH+q0u
32mBlz/e8IDwjRuKd0gJac+8SZ1xQm8xGDV8V+kJWwup0OEvp2x62SLtGbSEmF9B
F02aYJcbowaYSZm6U6KN+UQL8bBWDhJLcqxNhfEKVEA18RzpqUvysGJ27yzoI6Qm
xtpVCv5mLkWtROJo4qgsY0vSG2kuhxfpWZ6nHR5p1esYCuYu56ZOWm5SAKoA5Mie
yiEgHw0jJtSmi6oN0gidWESVmxVyAWcJS/3NMtxKxYyUFFuuKOfSrobD3uIVIHhX
0rRpV0f35m2ybjRoc+H21/DG+y4pSFhBnsOpoTzyNUp8//98Sl8TJzEth8pXenG/
V3aspsSBlWLsr9ZnKaZyb5WL1sVpaxtu8X0truafWmmETuyVmI7iow1D31tSa+De
ON5NEEWbPpz02LrL24x/URkg7n59rMGKEjZfHgJzjMyCrj5SKIJFHxAN+WekFtpo
M/nSm8b8QulKA/XG0p9e9/x4jLS08SjX7f4Dbp7zjbZZzFBHC63TTJkBdwfUXEPl
DF6hq7yOX+nuttZNGNYLHQjtDYGWMW0VxKs/Dj/FA+O0HixZQwatVE+ODQdyEgcF
eqW+MDM5HsdIdgCt9sG25Q9tK3Mfbm0Kp1FU/7/9wPPz936j04F6CQjrWHvcnO10
mA0QLNRyIgSu66oelp+jMLSDxYeCurs4dArDFKza7WG3Vm8hm4jmVUCKngaZXNWM
HKIRlZw0PAH5fCOoHfmbML6Qg9ZQEu9u5mRyX1A0OSnzsijPILLKZhmoO6efMUI2
d//jdVwgLefpFKp2P2u3r9QzL3h2T4j+jWHCfWPXvQR3BbiJpM0fvWGeGHk8Z4Q4
lzjbTaRk+aPHLy87WELdpXrG5I8zuoH32hzeZnhe5IuRRVsFWz1ArgkexPem3Ce5
LuRzgV0GNBarraTiQSNao2pZOyEA6uKcCYWqEPVkArvA6gavwn1txd3AdZejt/xm
4j27GIAXoz9i0NZslDvzLV/hqe/8DuSjrq+4/p8Lqp31IU7LYXlhC7YPupiwTpQN
9+oQdW5lRmDTy7gaXlPGm1N7lZ47iZaZHyruEIrXz2Af9eSW+IfjStDa8iVZtrhE
RiERalFuJykyX0aQfn1LmBJK4yTJ+ymayi58eKQQFomLZbCRLUFa/kRZqKdUYjE6
7YDqvrBu62XeEeum6MEVlZZCr8SOeg2DLIE+2VS1s20EPYm/qP+23wr9Xi4DWdnl
oPKsKBTu1IXvuntpfCzQOx8H4djmhHARzxjSCkX7gqsUAp/1fOTGbDJaZ0qXh40x
jQMb7jNmn4ykSqcUIHwxd8D4FV8hgTy1tguK+hK+xyb4PpP8aVvWV8QZdzNd28VS
T5pkurTdsgNMBJviKy++P9sHRvSfBlZ8BiI9VvJzEWG5C7NjqiW1mGy+MpQZEEzu
nGc3srOGFxul6tOFEvx3V25xGNpvmkyzdd+41WTRF1DKN6jn4a4DJ/ibGlgZSeeD
P9cQct8Ng2F7sbOcq5e5rZpVQ/soSNwBAvIVaSWEaAha6jzZr7hq/Rt9mql1P3xT
XyyA317A4sMQaPa2aTc9kP3HSVWln8z2jdxLL0c0pxbrUu4RhmgrLIznf+ZLRSW3
EDNvTDN7jkEXhWoZJvHTTHsQIEzmI/BKSIBycFwWiJfw2utvdKDUeb4ds1KZGWFb
Zd6K1kDAiveIBbw4e/PApM1H/FdSDatGhgMqyTX7yJ4WDZoQbnHS6bahjV8ah6Xl
TeNJPfx8qKWOgSzQwUUzhhz3oEFKzFJorYb2qWRrXLZZhsPC7qtycv5jWMV4IK5K
8+ISJWlA7ofuA7NraUKL/27r6/Id+54AAaIXu2glsTKfCo4Z1jVGXcrafx6ln6n5
L+MLn+wHRJeSOty/M9wj8m7OgFDn6Mr7pfC/cTfkn/Wl7G6nB5KwhqAnO6RiD8X5
DcbrmP6Mz3640S8nOaZxVhNYn9tX+YhW/X67KMa73pMDK045eBuGLtlYxD2PbhhP
gG+RyQn1+lPEZVOiuNj0/mD5LNa6GZ39BNaSuZQKoh00e9O394bZTkW7clvPo12S
byLNApYkw94BgoJe0p+4Fs7YI2NP1I1XXB9YVv2Sj40TuWMMm8n+ZZCYT4ckDcaX
llsQI8I4EXSFRXI7rDviMfwkCmVNUihx5UxPZTbDGnbfkafU22iZ0gCW54pM5v1+
LyFVTZSZfARLogfIf0VG+tNZOElULIuh46LRCxSg1Bzx0GO/K8UZOIJdXkbllJal
g6MTnVrX/5S8D0SzGYhBjDtl4AvJYzg/f+hxaXIcF5hwA2qBwbfCBQghpNH8L4fR
K9ePQxzYtMAoKdDJq0uRLfE8t/8KE2TX82y8w0m4zTxA1brsRAVaMjSp9gOkNEaT
gpDX32pDwMRPZixD6twMYzeoPPmWlo9rHe9oEZGu0e9yZDDmZObw77jW22c2N0rH
45B56coIRvl9h5nc6H3p/w8OzD3p77fqjtKf/RF8ZEeAom+Iwmfxsq/cdgvvRVvW
FrY8KEcu6gMOicdV/1/YsYAkj0YXWxnr7dfvp/Xm/YhKER2gvzCJT69bmOcbJdti
5Lst85sIxQ/kytfLLE5sWD7fGs2dGyfprhHbN5GkQaSH+Hz97Z2KzZVBDcq4/NaC
TXhCtkWloZyJwyQ2SoPhJzSU4GTnsreNSNPnv3SToLT+UfX/rhzxTwWqu5m3/xDE
Id7kiMQUnz1dpBh6YzhjClB/rM8oYoVrt8IMJXy2M0Or2g8tWvVUmWU4aESxpykp
qoyZF9/1T7TWRp+Llcirbvy6krNvokhjh3H8D96oXXFX53fZ5mEp+fnwtM4Bpk+H
kypir1penrfWIuQ75htFPSvVErJ2nhvwz7kGDquljoJzZL9Z+g1InG0tKv3HCHcS
5ALGUoKAX2B67nSY/ABrzRlncbgddo6QWryWpA+uFzsQWPVVLpDwQo/IfWZnC+uc
6nYUfJBlzzPaPsAq22BzOnn6JcmsP8XeJ0PPvCrK4oduehjtVgYuZ4YeHcRwbIjx
7oAISllNLfnH9rd50hC8YvhU+7+ys45QRmiV4zxyA2ZNpZbaSi3vWJtsSIiYkhx3
I3fzA7EYbVgCQ+84JMGzLhonCM/tF6HKg1HC1U1Pp/KBPAdvubsE83ozQ3+b3SHZ
DLLsfkflGhfOJc1TClwVImzLbCVltQ2e0UZFB9p4dfS3sDoKpr8Xxt2Ck6YYf3j1
r/n126FcNC0kgiLm81kXK9s5ZtCErf1UlsRFGVSeQ2MNPPPD5x2kp+BYqwAKiMrt
FMSEFzleanx4gA7pltqnZT+887J+1X2+RtJOWeQ3SURPZDKA1aONe1jr7zSR66G8
ClQZC5ekS9hI5/ZsI5TYQtF7yM0TZYXPmA3B2umGMXnp40eMKJFYxMDubwteW2GU
zZPUgTEXVBZcGOKzPstmzGHbCJf1HK2LFPMl2SeG08eM/oDw9Xqbn/cZtNnLdenR
PdEJr+HLFYPOuF+lT0HEv0JCAGyzBhH2cLjObpvArwYAk9Xp2AuylKJ4rze/DiEN
ZzkWzc0XbP6J0/A32oRfzDCNDf+vf6a5FIkAbcELkI7uf2pdAN7zXz7wTw7vAXE9
uP/zBJOz/NBmg6EMJEjgxf0YLnRQ6uMCJTfgSeYnu7S8YhjEskj7erTaTtLWxFg/
BE6WQesw79u6S3a+T3ev/4t2s+MW7VPeqOXzKiVmYm3zpshAXHj9uNnztatWC3Tb
09NzMdtKUX+I3cP38qFS+xZ2QAcBU2WXebnQBlkQDGtWqqDnZLSw2BdXjRvCsOHw
0ZWQ0uJxx9pKnV0tqove2fPRgu0NNX7fl4D1GoPcUy3yzVpV2YT5c+kqhg1Qz1p0
DhKbL4UqPEylGz8LLY2T4KPp9wneo7EOWkK3VznrbHboDlqQ6pNj6TFuAWZerRaF
GP2MBu9s92f5U7J7LYDZDpaqodDrzdwTBbhe49t/xNUzOEuYm2+1qGAhrWqCwOmS
cWhrI18wgfad5PPDZwbgYhMIITW7Og9FKUfiGhqnWwpDX1sa2ixh9d0rf7l/FPAY
iVgC1MQYy3h66L7AlPipjpfKMyQA+8ZLTLyrrI1CZuflCnQ2LihGJDlXVwEDOmin
+DyNNxYcf6o6Mjk8BIB8w61qN/rKIu/RmrrVvkl8CS2L2wgx7KqIr4jthZM6AZMN
H9yzT0objsI4AYsBGZpPK/UOePqZtO0aWQsxKYZ2CeI4phtg3AfiqFS7I8UCD2Lo
TrggoqYYK9H7zHC4cfkycBRveUItkI535kNBZWG4+DMM3hhEU+/oM1M2prGI9/4H
UFG42NQZrqoqXU+OgYDA7baIgTOgx8iDuHRFWYwsC8LiHV3C0ff71/9cJT8LX6qe
jBrl202EPGZqEVpb9zHs6l5zpzZc9fmEuaRIqNz9SupYKyR1WJ6ze++3o/6xV5UW
pg5gRlFJj6ayuIE0ZpCJMVZ82JF0zGwqxvJ3EBY/JykWI+U5UbvJGyeDvO5RVcGr
LiMv5LfvI3qIU9YpJS9OvxNzhqIAfWBN7EPjbbnilqH/KMZi/ba0mfIVWUsudJ8t
980kq3amRM3cTZbZ+OP05OSkt9qZAlRfEBNqyyIEirBEC5c+/UytH5mWScFeexd9
cO6g2mV3MFvHwtoj9JU+hDHdXhBvF2yN1XymQzjeq9Rf/5znRAKG0o3rXCwlfWei
G+WByetQiGNjaOpVm8MKutHz9r7dW8hB0CxgVX17rauXiykz65idfZtWX3QvHybH
7n0a78jKuHGiPzLjBPctn9cTWnSHc0wnkNF9ncZ8ipHOe8WhlGzDBdlXd2wHK2hU
8lvoKOI0CxvIoeRQ507g2rGqIXIrhcnznmIV0ytNZM1YOAa06TIFz6omxsG+WT+o
2FyQj/cXCSZcyZqFCaP5SMtw5zW/zN4gzRpsxyWicglJn4cp9YVVZ/HXr11IqGi5
yJ03CM8TkOVR+WV9Leaox3oGuhTn/WR0Y610rH+IePo3efvm95S3LPBYYQQ1Pdsu
MOtiDnqwov8gY09ooYCx0je/Jouzt+WLZIByEAcEKP3+tzcvsqUDnlF6AjKhiazn
ugfmJ4B6jFRYqGrjTnzH1bk8DcXhLrWg9OrOOLTgYRQc5Wvdjc6bD0odDZO6KbW7
2S/7R7oeuFbZfTCbd/nOExh+gB4vxfr9rSrFnE0XCzszVyc7AcwYKT6z6LsiybFy
c6HfB8UN9LbVIYmjLKYIfD3L2ZjgROvFP2sBlHMscTONWFJ7VMagfldBrl7hMown
1C+Skmqhjyy75ivO5QTlQM/vDlxjMfSi8j3g/YQHMxP2xgb8c3N9fdSxGFWoBlCd
dbkl/hvspJ06dSdeozZAR8C23U+XRjNQGhDSlroC3qOnCxhlIjyk7h/Bmp9jcIpi
zuxKXImWOjU+i0jFt8q/9ueIVjxwRNsDsYlrkXlybLYwH0zHW3mGFXMd7cOe5frb
R6nsQp4Jwy/fnLbgug5GeSq2swMbJ8vredB7aD1IbNdk1q/MfY/yOA7dlkUjhdy6
18I311ksp91uHPkWco/wIh31iWiGPhKZe/okebfAtMFmMHdNzD/C6Wa5iFOkfSwE
Tvx8Uy4U4gtzv6XeHB8P/9f8vD4bY4gjFFd1e9xKDevkks2jj/Y/Z2EpJTsd20FC
hbOTmsp1+lQ3B5I2h/GdjJk5INBhCm+Rjm5iqwUp4iMj0R4pPuLX/uPCVC3EsECc
RyLAOPmoXgzZflB+Cq4Sef/3tTyumDpf9U6l4JYvq8Hc/WSc1qvc+9ON3deuRUc4
5XwTzESpBODwcWy+AywDPQs9fSxWHSt4IKm2m2NIfSbTBsEpZbA6tJFkuk/NYMxL
qVhf+jLIyHpsKFtSoLypGFS0BnP1f0GLDUmEDbriZ5wcsqb9CuJgIlKPj5JljZdJ
q+4TlhLGg3oKLxm/aQGK5eJmqs8qerdYG81Qm3beYRsStAdVGuZTGyKaVBZ5mDIc
apH0DLJlBDUv1jHyiZ2JEQ4Nnp34VX0aBMFLRmaJVEUozjCqSRCWSxJcumDrIYZK
yWlwBHZ+r3rJm+E2PW/AJoAQ3MKx8KsonAIkr5oOYyonwxvPyLBYKDel0Z8bLk/g
O5EXYL6cCNl5CQ1AFNOcSTNsdhC2rJo4yD2ggsmjlHs3ab8ngW/vcMGAqjlm/D9e
Z33eVbcBvA3WBTZQ6blM4JsWqj3/E0g8ut/Jbo4W+r/smHecLxAa4oD00YuvmMwe
AdBdllXTke0lpLCsIOPCwUh9kHFrhxW6ClYICfAemtwE3LqwhOqc5ZKBXip/H4gO
aFvBuuVjyKvrDFhYvmObQEzTTreXbs8NEHtW2KZEBf7qvq9nP3gpII8XjOY3Hi1T
3qe+GsppxtD/v+3SkdnJao+kYA5fWcuNZR4b4gFcflY8JbM+4wAZgDuvN01ONW5V
ox0nVIljedOlbXnaPfcnT2oc4bE/P+VDCs+qfCCxa2cY4rLb+MZltDvXuUcZ1EnY
YWOnEzUjA29e1A5fOAtWzMFzKHOw1hK9jRJNO9hNkukDJtGEdzMUAOpHETIttsGe
TA3gCdyb2p4fXuMBGnWbQR3s1URolgTjsUu8fcRh2yfFpprq8OMEg3o6xVMIAlmD
gFePSvDg96MJtf+SV6ngc0MZKnj8yUIeqshFVMu6LDMlsn6FZgA3+QyiQed5el0x
PaGQa53BPta9rXz71edlCPPezzYJyS8dkXD6QEIcf6aH6nOHFKS52ELGIomF2FfA
X2o2RLx2UtfiOV18xGifO6MSqLjiJ8BVdIUm/q/Pb6Tdine0onrxoAaE4jvtKWG1
h7mSxTW6mRGRNToRNEXl1fzSNkciMMwSqJTUxITloHYMqRu9fFrBf1cOz5T5/rIs
vQ8HlnsCznr5GFJrgWQjXeFiDpMrYoLDNCAMX0yXZ2oLOfOBI0stFf57xyovgLCC
Ye/JPhERdCDsI7e7/t+J239ht0nWpyVyApn+l2F97HUiQNOJvN4AprFNIVTYnLfB
AYtdtQY+DGWXvXa2ETDSsj86q3Z02rOUrYpZ0Sa8rYtcbNUzAFyuvLbvkhV1hmiM
hOQ/wkrr4lgSqUblkKf16Vr2c9b/WBAaY2AJeYa5zfjfWX1z1/Qf+KQm2D7d9Hb8
UlqluJP5VN6T6oq973qZj2AFkiVg7xnw6KMtNWbb4UmCJ3nS1a41ttFO5JfHo+ex
4C42nPj7+CtlrZpB6/ZgSebxL4RM2MnqdmmLtAgffI3d/qnJoFwU6GhsrVxD2qJW
0+SWLnWZfiZXx8BF/tOmnJIhQOWQjcmxoFOpDf3QGyT8ayZtWp5QWF2ssq4vsLk9
lM9qTIhOmecnzDiwD91ydX+YCiDPRldl+1ScUKmQ941qJcy7a4iuasCoCPmwp9vp
zFYrkgCgk4ccbgo3kNphCOelCrvdJqR9styTjT5J/LJbp0hwUlrm5cmvU6pVtEL/
tym+CiKoNJANkbWYLtLRH5McRM/wZF+2ar+BobatNvmK4mARnrgHXhO3XvmZZyDQ
jdVm6fX9/TCpx0Cg8nQWMLoBdlcRwS06AIFzqZR6jf/s9KaDOGk8yVPdZV/04ETX
+5AsAw0kERrfzJedsn05FKp2o0X9KScMEVpDgHz9zPshbIqcHXsMvJcXIU+1/6Y2
VFQoMlsEHWKMFpGaPEDtHreYgVO76Q8wG1gvGwE3SoOQiuYJ5INapELz/ieoVHj8
1AgsQ0v6/a/GA2mjhbUcvm0RuF7ZX1lN6IuvX4z0stCuE/D/J7xIMgspIbQq56By
fBswSc49xDu1JPq59PewmfV03daalq/BkLpWn+sUEpHpBcEO6DZd8L1xlBPXKdcH
VW/D7IuhDuiBsc3p8gadCZHLQA2oErku0uPF4FEkvC5zN6wcpJV5BstpbEnTnIWC
NHfLlNsZdoDPO0ZmjmRW1y6BGQYntdQzRngo76hFC2LnK5k4vbAZN0ujk9GCpe4U
XwBxt6/c9SGIuUcQ+O3UL2Ll/ZZaiBB1DQgLaIufr0O24gKzc4JXE7nkutqQM9xp
H8MSZO+dNXYrj1DYN1JKn5cSWbC4o0/GBwpbWhCTYwqEtrj85+CW3J+tKxwy35Ei
B1v//xCw+UNaLnkTOLNjJWdMbob0X3TB3UYZsy7w8PYU46vfuZ2ZpW0K7yFHTUxp
IsOfH2oRun5Utry+D0V90aPDitNLdMRiaykCkk55ZCUcTpdB85Rdl1m3UwChfT60
RWds+EbmngoXK/1bWJk8IYNgicb/YGv0j1FUswL1rtd8ZUcTEqUS5utOBfUt6KFx
9qB2dfRKRUfXEWt2BZ6gDVJqUZu/rStzcmR6GejyleFtccwL8hVEp24yBh2ficXd
ABPf9sq1W53g/qHv/TQj7VDTaAdDFVQvzr8aElousxSXL967k2S33eENl6N8xtr6
weRA14BXn/redKkF77mKX4QJG1bAFNITH2JxHRX61AbIqKHGyWXSUYhBVC2F92Ys
deAyOY9eU1LlEIi5kLjKKkUbsJgNl4JwhgQmNDWZz6WT4CZHAnSHf8juKXVFaqMI
eiJMNZb2dHzis9ILu0pRfskhzK/Rr4PmWjJtjmM0oYaChll6wgtEQj1PiWUYCroh
u49T5U9tTczmR5D6IFNSmtfjUv1TyBhV/w0mwhX5pqSdKZTdBd/JLvCcEnMifyFp
XlFzrNSMaUTmFw004M/JFEJW9Vbi+bZF5FbsicCdXKzYZRhmUX3dT38KcStGIN6Z
i0hgEQk4OnbDJfRHF/8BfwQe1JbAfyYT7tbupGmrhbSsP+E0ZhOFQGldiMtlqZMt
S+21z7yJXHfhh2DKSQ1IfwhvuLCf2mPrlYmSerOsagjlzAMEMD4gXGWapPK6Pxpo
s6bFlOQMe/FIRuCJKuXAw3bZO/wFBb5AAX62Q+3jKoUvKgbEhnSD6z41hkWh+Jmu
xfm6wfzCPqQHaaxIEKMwLIVMBYnvcALJ9Jax/SANalg8B49z24pr0a/0Zqwssphr
3rr6anX+JOKBqlyjN7jysmOCbYXIb3i4F66bcw2xBWKLAfLCuK5M48wzdnnlpeyL
ajNgFC5HEkoyhzp5QkphJJnlEoctjZv0gYUrdmORwT6dOpr+2ScbpGn1ugWWPm0T
ib6/pB6Ae3U11dZoYcPl724rHrAYWQK3niRzuPdRZL02wEjacvGPDKu1SxfSvC3q
38/vtPa/QD2S8GbIU0lBMztsZwKH3L7Kfl16UZZq6JSE8wB1rx4DKIcjuVYUQAQT
m/sRLUJjgVGVCRKFfT0+XAaEhNK1XkFWeX/HrfnO/VckCBmStgscj3gC6Hai9eZM
Oqp48PPTop9hT5wZoQBwwroBhCQjajKSMelm1MTkPBW5R/W7gBwSKmcJ2rcISv4Z
20HJfMuCzzRSrNd7J4Ov+Rni/rRWBdwMIxj3dqwAL6K+V8Uibn6ogYEaO1/sClQ/
/R/cBfMRGErszoQ7epsxBG9kTKNv6fDLhhqA5lT1Lo0tGPJIJFLUN9PKW3w0XNPF
3MRt4c8MyKQ14mrTrHpjAClqKVe2bIA7MAO0kSOeBFP4HBy25D3qT4StNphmqFxP
WTdKRKD1LXTkwcP+SE2rNy/S0xijuzi1gW0/Uv5IZq7d/pwz6Vhe5Aa7uGbqQTRe
LHR0M1d07F6xJ/pccYm4+nTGLxtEHHaD/WFlbq091/58Ulr81xmEeFouLBB6r70Y
XsNnqA6KZr3DioOAqf4XtKSQmtFMqhSYvS7ljVpw6Zv8ikB3kOH7y+M/idne74g8
7HWLp05rspJjHsUDfejHxXimG+3HO+d8nsbRouQiu3ZrpU36rKx3MOeT8WuZkT3U
9qJq+w0ANc2GUJrQ4iaYfT3f9CPvJZJ4rZYJ5d80JTbwYF7XAhtJBd5nl2bVeSaT
qZRL/6awX6aXRnNxFvej0eaZ084n5WrFWv3sQolq1HyTcsHYXe1mIb7Egx2YnleJ
Sn7m70yTFKd7ojawhnkguyZLtoIFKD1hWrwb3zaA6+UCiYulJDP153iZjRU5+/XY
K+bJTZOJv+QEXT+hWXMRAw++TnZ1j3BGitzegdDxK9LbZL62jFezE6pwvgIsI21T
PpAr4S3GNGldl3eCO5GRqR8ciFwWVRSy+CT0wulNPDNqbgABBVL8Uwib8sO5jWnO
ivUEUzfWFAd8ebDqMQPzsAkPqtfHXUwoE2eZrbtoxgewkZB1l6Tbe2eRaBnFH0yU
cqjghjob0zpfzvDz8+3+9+blrQ553GuMGZjH7PEfB2SCXM9SSK6A3fgUPU6k377N
uBWqQdRqadxgucgiA+9HXplN/OdyQnURqs5EtdKg+jxqSxibTUJoxqj8YAuFQP/P
B4MNqNyypB7Jzwo0mWfA3tM8+vglhwPlcuDGZxnbqj4cVlxdCS3z1vC3nOKpdSS1
1CV0XmGvrbPtar8rDDSaCXjFqGexA+svvbYSlh6q3o4uWu7tMAbGlHJ+qobP26td
VVJY7dbecmhMs+SgZj6O5Cu/2/MDOYkWR7XdMnCf5yB4Ye6VijwILPKi7fLfRU/8
f8f25TyyBQ12ojgLerU0SktwYi6Wb3tws6HJU00pbyUB01KPGwRkkPQkgK1r1MBI
3AVMcfEpfDX2soS+2JxdDzmJ2sJB3b0HwOBGuzuBopePtPLCKPCByeXTphcuVJqI
qKSUlXdMCm3I77DG46jY0rN8yc0d+3qthMDPimENdDc6Z/aUx8fqw5rVj7VCAGlH
x0n+NeG3RN64jReZnfuuUmYheke5amRfxtOuWeos7hXzWs7YIAIcvEPkFvX/+cuh
Mje13Tf/s28G/pDpzcstCUmcAKCVNhpG3OZOFFOCYCCsm2y4ohaHBnmMjZVlRYdu
2HB5BCcoN/yZMP8N9vVBtHioHDLUPOt4nSXk3sMpDTTGpa5CE35God1jXxS8o5JD
B7aFz2RsKUloQSKwau0GS32VcJ0BveM4mFpQ3SWEmE/BQ0/h//zi5VFGxYlWtV4X
u9TmgR/701yzY7OLP1N/dI4VSKYUF8dEjk83nQ6hpTAyqiITmOpWvpOO1VGHuP0W
00Oe7StAoSPQC1EF1snguiKojKP8TwZEzZSuSxQ+sBcRQcyzhDEla9zDsygIiAtN
a1jK0JPbmhU7hYojf4pu3479EafmyzQG3f42jeL7HvyuBL8RbiopSjK5szc5DJ/5
FMDpGSaT+2B3LcUsVQ/i+nkr4FalZ+77C5bAwj7jvWFUNQcuZS70Nb0ktXnEM/nd
KEKUm6H5FO8qmNV3duzefEB2PI2urp0r9TmhCSxGD3u43mFbxQVyFKOCxqziaLn/
WXelkVKFbnIv+vR9Byg/8fDj99Xn9EGcRXDSAZd1pvw1VjtQMENeY2oBhvYMGKnl
cv6kq+qL45KffxeLiaF+wizs5+DOPyCj3tN7Zyx4ymGRM1i+mGXkMusjXNEuCrWG
aapBB6ydaTKVIu572BZ7aV+fmbyx9F1v+RvAzUpbL/uzZTlocYlbIOaq1OsXKZMa
5e8xqMpZLWoEUnK61Tv6V1z52lblLGDx0TAfHol8O39Q99TNWQi/tb/L9ETpZ988
JC2MIKcCcnY3FGkuwCtbN51GJp4NsjsZRxtekPKax1meQtdJYqYM6z8Izl+FMCdy
sJi93ExTMc4VR667vw+BEymD32xyQ0T8OjbDqCfDDTc7YNIcU85VR+4E+CsKi6N2
vsG866bvMh038eJYm6KN5/HoeSrzhDsknRux1VHMUaKozYYvCNHzgVvJKfrJLWbG
H0s9zKOPEoPquuhflfKaEmmx/OYN3fNZKgcX7DRYe/HmGG4V5sFzdegOfGA+aTRu
rA/jDrO/lu78Uo4a47B3ZFrAhQclikHIO/S7uBa/qS91FZqQYsmaZG89fX5myGZa
TjCq4PBmogckjSyKyYZaUmNP/DB+Brgshmzh9x2Aq5NjIaqplswCrIawp69daGgR
YdCTWJQy4QqdCZ2mHwgz+871I4ZeYwAq1Nq42OvDrXuIkWHPqOl48tVVPKNIxokw
jPiNuVgE4K/DXBOoCRxVY56yZSrYEemNtQ9Dw9Oej/Eup89m+Df4cZ4Kf4xJZjIK
bUZMpCG35EzxJcAbP1xLUzPECjD1WVJRPMNIuRJFj5gYSCd076beXMpZIPKxb10k
fsFdhRzkthpe7mhn28JeF/vnBUp1A1uh8B89JYgkBAki0pegTrVIKAkrroHqD2eS
nxVrNSHxqxk6xkft5jQazDiQSNVGnEnxGqjUoAnaW7vn8vY8kVDRXZRTVn0/CRYW
/NudmHOlljgDvIffDN1zks0n8MRYzUqRgDwC1XmyDMLMsSeU3xECMP4f3Npebt05
Kt3sy7/z5DI/nmt3aRxPLgb9Y7CcQtiF/HcKSQiselGKek2WxoAhf4wN3dczfWmg
0rTDcMxK28P9LQ0eWTG+4mOHEf39lL7NHsN05sfNUch9J78EflKksO2YIe/iup3P
GyW29wvQCgegOqC+OJJg+HyWK3iFyXgvhTk+yUyYLbXuZR0nSRqyivsLZNhCYvBS
OqDVp+yj1fGQb8iPGyzhu6QSWj0gCgY4O7zEBjYXwRN3LtB9JjnWAln7/d8/PzeR
YicReQf27GUOdVgM8aznzJ11lzGo3+KizbBs8TVexNsUZIS5MSeWZKgSuU2l5G/c
N84cmZR8JjW/6wFgAiPm8fg+FYukWut+eY2Heuh9cy9ZUc+q6eKk3TP0+lqXdqbW
kNKXwjgmyzJL8B5Mzx82jzUijK8Od01MY2d5VG3zDxYEdccEM1jtmoS34DgVfk5w
oWfJvpFPTtc2VqfHio93JRNgCAwtB5KZ5u8Nm2jW+sZw4LOm/3YGoMhXoJzh2UYA
1JXT5YRcd3K5yegmznnAPIUvkpog+sQswWaGaEqilDTkn85kLEHRU4Rhjun2Sh9t
s7WwltQwYWckjfT7sYkfntDSsqMAZ92DtYsgczVHFy0x1fW1FkZjNqNVEi394/eA
4FYnyun1pmryqjxt/i0O4fiM9PeccPi/UsqCONO/riseWw9tPOTWYLSNcdV85BT9
fCTPBunyHEq3JFJWb7JmHvycVpmqRHSEvH77JlTilRT5oG+jP/AA9rgYzrZqsG+j
6OS1j1VoJT9Jt+pLqZkiNFDagIz+mxFPIW7jOapL7QeA31u42Jge0ogQX7dsCM3G
tmPfmY7cUatWWBYBwaxQ6Zj6VHVbsQtO017lggUdp5n7KqP0m6g/fOckLFPzNI8I
ioLD/amNRzojl7Hf+DB4Pjbwkak2o8OIg5uX1LN9Rlck5nBBswvgzNOFpfsyK7T7
XtRGXsVBxpFORmqRu+l1xtPpMXTwoVHhzbHHozM2M8a0CHLFzTfcceyP6pJXTwV2
bUAYR9vzwsr8PbXXygSk7AD+DR5X0/Tk21CBF6oPcrdS06e33FZcn2Cjn0iLTef9
39hasC5jDz/Io9H/qeDvLr6Ovy0/UzCniNxTMLor+gnPjJQcHEdym4vWIfMc8HVJ
ZBA9AGJhNemP51eMS6nFfP/MAaVdrw+GQIC78OBYAsfpMnKjAG4MtmHWi7ASnZ0a
oXm7XFsjlWPrD0WB/l3rietRY8N6EWsyVSxQi3llvQtiunVkPcItxAsQOg9rCjOX
Ek797oX4SonkuSkiqPapvZNn5Cdubt7mWBqj6GFodc5QBuowGy1vdh0ZFUSIzqHf
V0sVFMjcvmPDZRPVz8KrTMa45hfioMnoEC0/0CuSrjQHhgPFKA9CPL3oqO/oFkc7
mlfpPZ7Pl86lz29psBB1lEJDFLyPqyBJgWjy2z+IR2iXHRQQjVGiwADj79UQ9Dpi
Xwi4mxQJ8NV7rsyoiJxcRvsl65sQTVVdM3p1yoNuM/jtRZxBxCJUpBJnFUqdaR/Q
KgaXcZLlptEKH5BG7xvMFbw/GToqmZsJ4OHLwm/rLSJFxJeZCeLrL0mHjjNtV2dV
tLEF8rTgVkDtSjoQBDV3Qgj2iWzMA/NUMCDUTJylgQfbdo+AgxpH7eRFPafGz4g2
4R5/qJrE3vETdn9pebf7vERxmGrSHyWS8Fapk1IL73QNS0cKXikxG+MuHL7GAEaa
I2w6JADtT+MGUfu22dXxMBByNdYtCf8g0R+0Ms3ue/SCfudi5/ztbgqmV/wcV415
yFnwD1APr+gsHeJCLF5azNPXdrJ16ytQtoBrGXKca47+Dbj0kNoKsynjCWbxR8T/
xHSt/x3/bRkS2AttnguAwN8T8997YcxjTdoGihmUb9oRp4W5FGVjJN4unOll7iEX
hLOmuwKPSnVGjSFg7/fkaf3QtFblEsQX/FD9ecO5R4yNMNc3ZQ7IAP3RbEcA0eWL
yFhfrccuAADUBGwmraFMTBNPRDIJWsg+uGR43YFaMrJr0MCDiH56+sqilzDHbYwX
a79Zq3oDrLadxHQ0/O8h/lZy7KLvfzdBuuX9lpGymqU81qespIavJ3m085xe0fqD
FmslWSfSALjtroKuvHcq09PnmPdc9bAVZstQYxLKrw0fkSu1JFJp7ypnQeEyMnCr
lCdNvvihDqazyoUGdPW7GLRXbfQoSVprdR/w3nAvW9DlVqdrTk9LYiQYtA/xp3ob
iGkA0BnbCfZIsSgSbpbb9ZW2aQfaDwWSzsGQyAfnhrQtwJ/brnzaPjd+aNnULuG6
Q8hnzLT7iXUgZ3n788Xc8DBd6Ht9OQot6n6tjApap8DEuhVAJJBzj3Rddw6Noavl
irFucgfglPSTrEC42o3GWXHqSf1zT0bVGHXTEHtmjQXsYEfBa11YxsNO/zfuRiKF
xsV0qIWpEaYypt5dtiR+y6Qr7g/J0STKeXCWuArYJlFqfwdsrz5FGHfOxfO6IJcl
CWsqOqBC43Xw0to1rV7DtXbZ2EhijVUXyfO0guIAqN3vvqRksQuqdLghpYl8ecL1
Ue47xB56jt2glk64Dj9z8DCJzqdhjCZDB1gc9pYJC0ZhNy9ACebtz12e3rXe7TgV
tHJ2xoXDSB5iIM0qfwbeEayciHXKYnbBVUiCUGH/YKaeKfDWOtRKsCH2fMoxCgJZ
D9Id+hbWEAU3h/boZi4wP0C+JsS1YVqegG4ZqwRwdxk47Se/sCmPFFKH7CXiOgQi
dG9QkJWVvVPNsSXM/YKw/hz7ptbsO6YfGklrytNvE5bHQzD7GOl1yIPji76Ej3RF
wy0NfWiFzYgoqsvfVXlOxTaKKyefRmrF+QIr0jP2B/uIwrRFNl8aQZR/lCmPE+8G
kOq/keXlTkBpQcUDcuecQ/QcvUSOOTyOeLmr3wU5NiWhy53J5oymaeFUxoKfv0VV
bVEXGzeD14mp58qDtNtrESFAIunsp0vyxl5NHkS/Aa5aNdWM0kdQIxc41R9oXsRC
EATONI9oH0zLoVbOEVTeEaWE78o6AV4b8IZEByKA7MX7/47WuWfB7wfqPugwnXhI
OYoy0D6dyxRVRsvUAoqsP7HzisCc6DdugDfY/5iJ5DxXUgUyqVZTmwYDx+5wQ3c2
XsOskVbSIUE2jbPRRVA75XCAuV7yOy+iNGYc2ZlwX9aXL/xxs6r2tLrSnjbSYmEz
1yhpk0YvZfwBSgMl3gJI83ui7Qj/JMKkoAo0sIBYHwd9LVdpaVG+QN/5feyYvWIE
8Mmh2yB8vNtRQN+qf/8dqfARcdVDJPcwn9KxksXG+z0qgwIbgmFjT+5NusxAKs6a
5EFsS5F+8zQjrpVgpaooHwcGuAqiCcY+fcrNpqADD+NoUwIE2ZAyvaNKV43LYIi/
rD2i9a8aSwU9tWaxqhPA2dR4/ZLS2WhQxAwCfgOE2XFi8rC7Wmu3NG4oNEibTMlO
a1ZbvNlf8YrABe7PR0DmtMttLR3cjVwq+lVsw7K8pDAW3YtsxOSqlkJWj1s3MiLo
OTfoygsVo/CW+0sKS1SxnjzesD7F9H7I9b+tzdM+4S6g/Qv+5XBT4Tx5p+JO/XYe
wfmLlvbzFw1hdagrXqc4obDOoxNPKVwWx0iA6CCzts4xRAAJ/alsXIkrGMXfmnA5
POx6Xljuufn3vQSCK8AEmHoex1HUG7BrY7eOOCbEkr7zZXUS2slQfn6OWkq1JuOo
ngvDC0ss3aw1eJkG0uGvmxamXEWIRcH3Ob9kuokMMU+r3uySSOY7QnCtam3lRfO6
nbL5FjoUBZBo/v/Boh/gcEiFvOjFDR5QxlVzxCd70wIxC48ZJF3E76Rugg9VPeWh
uB8/wIJ4c/HdaZE0EWI4FTMyzQsbZhnKmPHBd7+wBwZMsm0a4Os/TzPxcCrG8DmY
/LAFS7VcloN0P0Ot6IXoT0gRwqMcff19PJW68mcty8ig1xBOXtKpYeeQ8OSZQK7S
L2RONDg0EB8FfsugqnKGOHWF87+5nCJvDxd1D1Pwv+tgVp5JYXG9egktqZSzi1ol
F/Yo05qVvF5eFKYXGPG1DyhdKGCqGI/7Bd/H7OKz15rMgQojMBTUW6hBpLBlHIHy
yKabrThCu4DTx6alqGNC1f6xSNkGIx41YyNrqf/rIP3Nlz4UVzOx1jKffJ3fexlS
0qXZ4fKhzZmJo/kV7XBpBeXewmH1JPtG6KALRhtdY8P7EF0IBUMzT9972DjKsH3r
0SN4Jtf07Cy4hnMgGAiMwD4qFGc5Di/WjoGFKjh36aiER7WYf5GGQMKZZRceibFT
eZRyuSzc/l3qx3LjeqbW/R8ElSgfvxs9W4JM9Jfw0KM4ayegecNAzSZEgt9C039o
Gc3FVnEAAXX7Bn/ClhXvF5aI5wNaI5gqY7QmloHvwn/KFjRebZTjPrJoBDKwew+S
8X+5vJz7mJKxFN8DB7eIRHr2ab4jNKOzzbWqGYTENl0oa1LdXNnkykR6zhnIrz9V
Wd7dkz4kXXoUuaonjWXZPcy5yn+R1YBzVQ5sso1sjFRY9XLWV0ZXTJU3fJI0ZjDf
uCjdYVe2jx6XbIT4Esy2goJxIRHGHbG1DAWlRpnh7JmZMMJigVYhGQg3LeV5iMik
/OXStiFO1qx3MZrMY+RxSkjbkYVo+hM2bKbowsUnouhQVk9ObV5LDwZsVHrxj+Ns
os+MM7BdKrksZb2RYJpFWfpi10BXmA9XB/kZyClFtzK4cCgHlox3AmieLl2J+f2m
HMIdQ+PlhrSb8GCyyOX6ddUQoBP8iDigvvzrQndn/aw9upxBEp36qzTJfcxx4Wbs
ZmqqDK/FwIP1maEAF4DGWewrOR0KqfEqHVmDJsbrlfmtjxcQ6LEk89h0Bh/xNBac
7s+KLp6u9Aux1FW/BXuSMpO05F83u7f00dBtsjo6PLC0iRtc973Wz+9c8S3+XAs4
BfXY7gvu9tkz9NplOwi9mn/huiNHMe8MVl5YJIsRW+WWWfH4yUCfa9RtjHRXywiP
0AgAfV/sm/S3xYB3JD6igcOg/BZr0qZyn/HyUQwM0EAk/5KldfIes4TVL/SW0A/q
i3NRdyGZBtaCIc1Azxd3D+cjZFj1ymhPticQ4zfHO/PuB5QuRIZDZ7q/7fzFC/Oc
F1JOa3DftsUVSbPRaUyFiM9OJrCaP7g7tm8plD4X72kpXzmxSmSl/I6b8SJmHYm5
uF1OychGU1DoAvltxPxFOJmfaKZZXjVRS6K8/rjSdIW/cF3p1eyAMmxbQq/kndZB
aF71aUFklQvrOYLvrsAtLLKoT+23mbop8cZLQk3Zgy91Y7GMghApTQiuSFB0RJ//
iQLw5iSIpWC9CvI+2M2/xTP8Ta7ljCBlkbf5EirEUBwV5ZcDj9wAwSmDos2sOxMu
k/xt7X6MzDwlY62Q4A4FYBiAwFlIMn12D6+GkJbT+vcwORZdD9BmutaGKPYysasL
kPr/Kh9z+4gWrQCAGNgmxUkslo/NlJgZDwebKlTgsOKfbOuht7+j+zTSd1vNYoxo
97LKuJutd7OkDExxkh7ubn3E8KdjhXn9EHe+8rEdFWiM98uT/X+Vd1vodmkP+Ec4
iJ/2RttNNn67DAv7Aus3GrnNTPSapey7qt/8BReG3bLnQYGialmaFaZa5Lib5BHm
GVE9fwwUwsOR8NvJrLGLTio5qe4Kl31SbE2uB+OvdcYg5Y3QnS5QJ+Bwuykev2R7
1nLw29KNC8Tq10HxTJfTMa9r2MAgydizg6wjIHgsmZrmUQs+zLYEJ/oC6ePDLv3g
mFy8+5UZ+3HgdjV0a0SFkmiK+grjgF49ngjkImxWMiE+BjY68ICXIPDyq/rL63AY
zqC6MCmea2Zv+ViBxen87uT4NVUcmNKUqyoP4uY5QJkZFUach69EPod7KWGlt1mS
RZEXIDEA76tvAm3wBQzBIhpLqCFle1E4XnX9JO9fShQvpKqda3ty1FGoLC/Tk45W
GWHjj+9hwcYa+zAUzcBQo6Blj/rZZUnrOBYqY2RhIV8uUD/X315o06KFC7+bZGH2
+fUwyPNG+yBgwHu2FQg1D+bKLLZI9EOCl/rR/EIkjcOgcXhh+/NkbafbZTt/dNjl
mTQ/FfYGx11xsh64T/BKjcrzQ5fBu4jX7kncSz24PwxfmbgtJy6ESw93ksRnE3fj
dbqxtSED7ncAq6I/gtSmFXuzFH1ktsQ3JjsmWui+ZKrIO6T4+w0pL2NYjBM3Gfae
e0ozV2kuIScF/bN2hCg3mxh7tBsJ7XyVTM8tH7aakID2Pm5VrEQqiBGRXCRQg3OU
4YlmAhIZ4eom8t5wd2IzLjcwTdY0rt5dNvPUUt5iz9oQIOHyw4NiMViZmv3uUmnF
NS1kYCOI3CnU51mBhtMd+3vApe64tleEaK9JRcvgE2mM7QruggWLAS40N/h1HRXM
52yL70hj1p7BhYWQlr7HcfvREpJkV7L2zwOfGs0tb1V8ZS95Tq94OYVWX0OcbrbD
SUkoxyzdUeVXEYXza49mddNhNYBorF9fuDKxFcR5PpLy5RJFeDXM8sgETIvYSqQM
oEdn78PAYe7O5S9/lr3FNFhZLCb8U8ztsHpXsloe+wSPhG3l8VLb4TGZ9TUbrkXY
lQxUjHa0BZ6ntsM4/OpMmg9ZBJIF45bWJBiV+WqiESXprNJrBln0wkrnPgHFmtCo
1SDgZydShnKSJX8BBagTKTel3Ad90NAlBb/GxfnZlY5Jf6rc+xs8qEIX03qztiGH
iKMN5pfGrVVo8cmUarBMGY3KAagq1AuNRWw0wBqFVZfmV88xbd2esK7Be94Qj7hC
YezO5cAy+vp+A5reRs+YfUZ3M37yyuK9UaGi9gKQngWbTbBILwu2J3shvrHCwPaC
fGwyx8IdmjQeAcv0Db1/mEOMkrt2I0QvDz7TOhIX/PHaOA64PS0PPxgSPaJXhxgj
4iRXpGdfxFZM8EwXwn2tovf+pPbRnTUzG1OLZZ1yOVYvcD+HqezoceFX+pCFgU6O
Xs/RY3TBeAthLUv3qfAScPuMBlL/WL6HZ2lkQVLeISkrB8CbIPTnpflWBwZqVKaO
ujy0rw8K6vd0uClKSaF1h5nS/PJVxtDN1OLVBl+gb9OHZqz2klXQRAkYSN2l2jxi
9HBpFxkGPOO9j7Xp6zJji9GZ3gv3bSruT0nqmbWefsWOSOV1ppiGWYkEO0vDH8Z0
yowlatUb324ztjGHVgpGsrFPkotoKQ8xPAplcqkg9kIrXYg6/EivpAoETWD0lEuR
zmgpJUlRe2ZmIbI4Nc5vmnNjYnnOM+nRSAyaqMwwy3KsAhseVlbwUkWcV9z4Qp+0
IzP0u4gUirxRqFz5bdngH8dWCAMwo0umxCprVaysaGiz4Swvq88hXAq+A314Xelg
ZcK4fdNPoaqYFRvBvKeCpQ6VWUdYUH1L8Xsf+L0uUTqUsHWLL6+yryEgFt/Go3FQ
rlsBjW0fjJZYY6pdjmDYDnsEfEMI7o7bm35eXop2Yq22GIG/jKkUvtRnMhSS17B7
xJmWsAcCOiLMmQJkq3V7Sjyts9+Jsg8BNOMRotJ0qPRAbyi4vlWDjQN+x1zhA43D
bzRfF8ktfMoV+qOnbX44IsfGncW5txXQXvikRro1dhVEp6dwE1vstdxE97jOiXuU
cMmDKe80GhMszpYEoMRaj2/Lgz+W5nUEZ10jK9rcH2zxklboFviVow9Ml6tEmF+g
zgDcTjLDMxltu2IAkdQ51xZB3ZqsmXZsbYbTWE23N+OuadNJmQ+lLQaomUWkf2bC
4jBRPPFCYg1IeVZhbvQ7GXwoaMQUXTb7sdrXKl4fr2S9Rmjdx8PiveLERaVlcfWv
74umCWJrNJlufI3rslbNRLsDXphuuM3YDrTTiwusgSE17EgGnN93yV4itopTvwSq
mzIpFxqI1lAqNgU3veuS16Oyb3KmOyYuogPCenipL8tdIXkSKwdPwmSOC36ZwqOT
Sdrxy/EN7eB0uxVCgmrWu72vcCu9phX+AGaQeY6W6GrcA6SCOUUJh1JcuVV9cKqm
vezqjzQEBEDMe573ovJyh70sMzNSI5+UV9jl5ep8Uj2kFHA9rgew1cQRLVfl9XXy
4hX/xKW0+SYZQtJNQ9167ko/RDT57IQ+FbMVfKOEWRW4mbcsKjO1ZImFFFau2M3I
K/qwLFyt9SB6Zni5mMot1g8uxDS+5FSQEa1GmEuITkbjt2fUIGJ4k4jIOnHzj4Tz
2h2wamSux4/ZjA0OzB2fDj2PsAe1WXj+p1hYNRSS1PdC1Zmss7M9PpglveRUfmzV
ZiHRVgRKUVFWWqpGXsSoyBToT+sCC45ji7HOHd5HhJl1b54G4rdX3uFqCSXUD9+W
gbg83+7jqmPIn0buRsnkfklNHIDjri4+6sRf1xWPkO9/kLl1N1sFZr4JS+Ya8Wd1
RZYzvujYnic0DrZTkoM7E8LPlxq3YDmSu4E2ixRb4Ih3fdHnRT018ilAKCT2NCHG
o/9E1BGXfzTXMd1vhYlSXyZxcjm7cYSsRUdWib3dVFph0ixwZafFzkBnFEHYs3Od
PTqpoeHebjXl0NpruTtA3eEJ2+XGmusARL093ftcRbCf3R5T0SW89brlWiS0bmaR
W5P3XZvEfBB7c0MISHXNz0XIchev1vTfF48sMVnF91SsJXMakCPM0IVf6WstYpWy
Yi3vtrvrrUBiulWa4jZLZzoRmdTXxG7YDTAy+weHwAoeMSjxG726su+1YyhwABu7
G6NkIyldHNfxHr/vIIRCsxr7LpDEjiVBHMAzl9qzwqF+nzcmEGcVdrlXzykohmKd
gJi3YmxL9gCCt3V1O6dVOCsf9mp4zZY2dD5nrWmCCo9PZ3Wjw5bFfwqKNtW3yR5m
4iEMjmctGcdtdRbyadSJZp16K9WMma2NKIkx9xb+aU6BxrdsPNJzqoJK376NG8H1
GKFB36jycxsTvHT0G1UQjKdKGML4lHrJlnE86++Uo5bYPbK/dhubT6fqrbRz8tXX
PHFW5Xqs/u7rr1KlA1zeXW2+vp5tENoyFS9qUbA7GKP32oD8+8OtgNNjANrfZrhN
yutO16Sveps2mFeqUpRbPkc9wTvvs53KXvTw1FirPCv0BpDZydBcBxwRAVbBgiaW
s1lMZl4D/TxGpeD9OR5qnF8FyEQ5LYHZCqqYhVv8ToG2sBWEXAoQFinEr0SaHci2
9e8ZCvu2Imz3e/ZBz6cB5Bh+mFV77QA/CujcQG4nwP5+RzsBpy48M62JCeNHQc5j
9p+nO+zuoj/eB6RgZL712LYNdxxAHhfxWMlTHm9wbSZgr9Ep/mVwCBctbFOfMtD0
e9iPEZzS0BMgB6H+nB1L+ynuS64XfX3uUf32HT7RIKSAKLkok08ay0lgeUKigmJK
iJDGQJ8cZ6dbfq/sb5UPGg/AFVFm7VQqPIPl07UxflymjQzRrbyTJ6Uv6rq/OMZY
q5a/fqhU5eXiLTp0FKsqX7I9soiGAEwTHd+RT9bkPa5kbCVhPYv4oJHQG96LAICr
/kMUpmOMWovaARM1G5eAgcAzvrEZ4xbpuQxjIp7FuUkBnNmGSvYRNOlthyV8wRJe
GDuH79Z5KOjLZlN7JYWJbvvueylCIb9PCZ2Ob2fS+2E5eULvRsa5Gq2HAA4ksBJL
Kkesyi6H4rvWOoc0qyqao9vhBID7nNlM+VE1iUeyqt66IevF+36lLVboCRHJ8IPP
dbjsvf7+4Lvtzl/olY3+leKpWxWCcODx8srwCUirZrB25/44vB8gLe3WotbZWdid
N3F7jy8MCdgCsvmZojHq+4+8e6ZElmuf4WcoLwvj3cTcNjsmA+gpLXseUnNim88c
nDnfl9CKZCXeBcylJuvx+S12o2paJZ2dZISBApioTwsWysO10M/JCpcUuBv6kkOQ
ziZL7XnxCQjZ8JgufHBzf7ylTbOAR+t0P8TKhbXd0fWiVplk+5QPZSAK1cFvx9uI
qGun5uljwegHcVtL8XDmky2sJY2itWfKXuSz52/g+SIM8B8+j5EKXolLRF+vQSwc
9XU08DsjjIRJTsxpEs0W2p1Dygizz2MiqruT/IlZp4qWdsNroSIqbhSU9E67boOt
HHUn8pDrFETxzYmFe+mqCjM3sUdI2jhAH3boqXCr6/Wl+jehDYAM4ZYl+3uB1gCG
cPBpvCTGRM3ZBvz1aqXmSyGT3WWSPNwFx1NvCe8ixqPP0J63jva5cDkvab387l1U
qM/P3P5iON6mAUB40jitWxk2PWBFNxBdSL7uKdc5c5MEY0gYhWOaKsL0kCxOUJOw
P36io8ezd0tqy20R6DU2rVnTIpkd2028qyRmNEIe/0y51IC0xqiB1CDLrmM4Nlad
j/Kl9SpDcDXOS8zWen/+8PQMTWZ+ZMOhaziOH6ngUE3gbtrEeRHzNtR7Y665Tauy
HGyA3Lulb6NZ6YL0KiWPY0DNCPc+sjkMTRI0ik65UK4bJ+ZjSTkudJw9Gfdns2WW
e/i6UsCFXQ1faUO40/W2c6se1/g6sK1rF/7RtGnEMlfdVrG68Gh0SY/eVzgMOoM1
GXk0uyEHjefooXnKTF7BBjRdio78JvRUun3s7ucc23qgI/1JEfci6VhSVtS9hm/N
tgBf33WxhVpYVN6DCMBll61uaSq6irtA+briBDWMStFxhL78nzmqNS/iwfQ1SwmV
Xpy1bMCgOP5ahTLNas/vdlRTLBpPn//6iiSGqygCi8p6f1OoYnG8y8MlSwIf0fEI
oo1qtRibGbYaWBjYkLIAcHvUw04zyNj1FrCEE+KKTxAVySzluV8kOdOSe4JIuQ27
VhXHXp4H4eoWM6lRtvOUT4Ku1+e1xOWVwwCNtz0R8xZqbSRbbb/8FjY35amVtVAX
pkX5LQ8q8to4NXgcNAfYkDnbeISLxpxYh42K25nFA8WFQK5VevJLCBKLlFo5gPoO
fBSIpQeIhkG5hfr5P7e5cFqInug5oZhR//a3ciKKCaqgW5/oXrTeVRB4SZ9aiqpD
pe1GToRnPhMSWlnZnrGgnrgtd1hfhi6AGli3246KxY0f5S7JSqOIBYNLUbhJW/E9
ohy7+YPJf8lRbN7FAQYDKaHK6P7JMlE4kyQkRhgY1Dq8Wj7MHpLo2z55EDuEWidi
pnIAbQeGIUPAwfwXRSD40I7rX6y9I7vpsRqcJYOwzkZo2hrEEpQc8XZLR7wQvPqO
8hgNl643FpLKdZ0wH7wkAnHPX8JCnLS8d11c2ulIeEIXEF+bWKDeNmBkGBcxywSA
bd/T64mb6YRyeG4Ws8Rw9FtOs78PcyuncyXXU5nluzTi/FdydpXikrNSVOV9quQ7
hAMYy0DO1X6KuuKZxzx13hSZRoeBh7V3SFuBkemH1Wac2yoJOlwrTsJpI8d7A0/Z
TdLKu2jTJZ/bZPALuOMSeUzoRiAwy+ze8OzOhi68lKYexsQ2w0Adm95xjxQvWz0X
VXLg+t9+20QAOilx7p+J3atJj7Ih8dXMIoT99/aZxdZcXTLqaJLsdGEahWdePoFW
tfnqO0v1kq0NN3jifFe0l+k/0r1FGZ5OotBtK0qgYT7IVWd1Kxgn9J0QW5t97H4I
iQ2ubYGJpsUZwWz9iHbZlFKzDVlEK3Q5rZ4JzgKzGSXA/HTzhZm9gLdsJoPGnjcQ
YYsVCc4QYgT9CLfwb4/by1vWy3U2c+36H7Ad+rbtTshr1P0bTMwFfXRor+gUrc8n
IHnSXpt8njHlwI7x0k5hfHBxt9ErlbjJFhCDKm1FT9WgpXKAAnl9fHf11BR4UQwI
YK4+rJGZmpCd+NSNlW4C3tsgfGtnQXQ2s7Gf40h7sNYZudsyaDLdU5Pj1EXAPBZt
zab7ACH+I/GDuN+jX0NriLOSrP/ifwzEEY1sCxYasr/kEgPmVdKMafwx9wT/Xzwv
IcboMuyTWU9wdmqVuBKge8KyjraVH8cxvB7TJ9ZK/wvnkUke+904boDHwe5SyZI8
ejGL/n1c2GN57/b1d1nvQVvaCBzoBpoaufCpJaYYjMStwpn2MDu2RTj9X98lYcPX
91pXjVI83TulfblA6kq/xM1qtn90gXh7axoCHBPcY4ZhJHUIw5s7RL+Q/TeaFAlq
A3wdOBm4ftdFuJc5McfTvJZIU/buQu6W1KtOS31n0rNZsfmE1bZLL7cTZCDBaLzq
hAtnTZsMH5B24p+sawMBcvi88hoBsi8UB07HyraeovNZWjq5T9uuCHA26Q8h8LRL
Q86pZTKa19LCsvUg3U0HFL07IkIFoL/csgXGNsYszMDgU37MzxhzkV35f6wXdHAP
bISAOqD3BEClhM+8yIJKvooLs9PlTxxcSu5y7jE7Jv/cqhwik1MMXyx/KbjLV9iN
6mTPSGuI+O53+cPihpDmMt25SNAdBh/lDa8HZY0/pwQOujIMrKrmSIjjF336xQvS
44YJj6sNWOgku1R2Ck9xDZ0XPvzG5MpCy+vBFYZaJECsdoAa4bgu1FBtOg7k6McS
fStfz43W/qtC7sgD5Z1j94RYyV+NWOKqXFcvA6/FXuxXmmwSaxBx3wqdJUpd0wKF
2AKPcfWdRy8eVQ09oiYZdiESyINuSISrcs5Cwxdb8+w4S2n8sIxGpKR6F6VVMHsR
TLyDWZ6UbzbOTZnGzPRxioSuVaE56gmoxjK+loUDTG6yTkpwF9R4Wlt6pUvj7K10
w/BY8bsEGXxg1ro8mdrVZpj1FQHE6QvmHitmVsChRih0AbyqSKZqTZpziH+vb41K
YzQ+X+fNHVkSI3WaKMeEVO5rS7iGUNisdf1Vk2185Jlzl68JJMpwEB7xQJq5GUFM
3GQ2L9Dsd+S/hTsCSoQnnPYdV89wz+BQcuOKyn0ezp8bNkaA6d1MF1jRH0Fc2t8F
boxcnNMxFf2Gh0iikS9ze7chMutRmkZkXPqj+BQsFJh2TKztkRks3Pd8iPpeZgBw
7OPBCf/umIRnfJhPvOPBV9BsqBk34Oj69BOiHd7OriJP0TtZSckN0GDVAfNkkfNk
DVXPV42ok1EY0/yNAq51qYs84CyVMZ/rFfbMqlDqCu280v+XTYFkJcTBkEpAGb0D
/YBxE5fXWFE0Yn5hmWx4Z9f+2WYlH3wbL0+1Cy0Ffps+nKajpfl1Lg34px79dExc
jBjuFxM9ckPxbuPogx4sAVq5uMqEaMa255W+Xk8K6GmL901NYiOeqB7JfCHLjCQE
uZ73HRRMGel2EGBtJM4Omqk/g1rFMGTH5ayUMI4ajmLD9pNjC+4Ej3I6HIDAMlH7
HKQtM380Ypkm4rfXfW2UYJDtvzbUBVZwZ7ytT8b2gAgU6ZFZLxCS+C2EccIBDtvi
I5h22yogTpQIgpPui2PlRiO9iSXKV2963mb+o6zft+8dw15+/CQvYQHxWLQP1YtE
N7SUYvUApoLyO+m76tbK9Igp4RKHF9VvMtzpMXa6GLguALEArnfhatAbXxfUxpO/
X+JXBmYtWy8jV/heGL9npRXOAvKesI3a/FLjEsLcDyVNxjIk7ydTsLjigI750YcO
8Za4vCOr30NdPMAxIEx72VA/QYYvHkgYFaaWJh9776DWEmhrMakCZezAx/2FTTZ0
VIbgp5JgBfpAtQYSolRbWp6x9Yz/sKU06LGrydpdhleAL1hF09S1MjupeYm+bBfa
DVsDAY/E0QLZlC/xrdow87ZXqxIJDn9OkJel0Tp2PLoHhm3zzPD+HaBuaOX/PwXA
P0IjQTXqskW96o8PISXCk28yMDImFX0SfbK+hZ41XfS4umJPQZuyRvRCgXe/xE5X
RrYoLtbAu94yKzuS8jR1ZPq/ug3QGRwvWapYLHjQx6CNPIHzBnZEix9YXIFoInDg
BueNL8379knt/EOfXTxhvwN4YfVX2YiTETcc1W5MVN3OVsWDmxwYQ+M8wFO6dlMN
cHPNldyW3KE+3XOMKXe4loimTw9V8bFKpwrW7qgdWjpD/A7HpwBcGAm/Q0D78wdz
110qdBRcJOq5N5eduauF9WjKnnZQGQ+somGGDKkicymCUDJSlLC5U0GgH/Nx7C8P
Zjib8HE8/sKH7+dhYb7GE+cZ/LUXndkxleJ0/ZBFXqu8pICBk2BttCVSGnniZnBh
M4CSpCfOqU4bS88GEMl7/c01AK6Rx2lRukJuE2sPN07+UO9Wid001tNCYU/vPoPM
8UEPOjAesuVbFlp7PzvsWx2TaSzsEylwfyiA95ly0U+8uVJEiAqTPzMB38W6gqT9
tCgYOzPjkZ3MklV0VzmahYx0h4fuYiKf1j73gAL3NkXg2ZY9V6igQx17z//WDfVC
3gVNvxn4Ko/FmBRs8bSM+Hk+tNryteu0u/dMsBcMn4rjeP0cNEayOzSE7tn4nbEQ
qXGaqotaMOMXEtPZlUyrzO0QZ+AGCjNWEUqzvjaJmEswYg91mhns5qvg7MOzZlDG
bNwqdGJl2HUFJki9bHSVcGi8/T7FW7UMUXFK10MIzMiOYTJJf2ub434Vr+D7/1V8
E1j3Zy3ei++vYTLSK4MIPwZgzWCXXnYUspBYO0jbgCkhh4240YfNh/SX21h+h2Xj
cDmp1JrMVqXxwxmmjSoCwlUB2fOW+DKcEfo4dz5UpUefGvyW3T/VzFAvd2tWztrJ
ED0hxzxNzzmY34c/Q1gc0Kv9hYmrrxUSGDfF5XKF8RzuBbM4zKUKQQmCmfz6WKfu
IUigmkoDR8pEnGamnMWpYDcn51v9T28SiI8o/0RrfoWPSNR+z6FRfV/WWOCNx60A
hE/qunCHUacQPk5cSiQC3Xr8U2QimnceOzS3EIppQnN32MmIkms2LpN8IPGcBswd
fAFvPVCe4SjpRAJdtoIhSvwbx9Cze39CE9ZbUYUgAr7+Tk8z2jedbHeN5feYE4HX
ZqqT6aKo98m+49QjRhGJLoe9LM3t+GWzm/RkSJ7WtahmCtEqqSwsoaZpLBogicgJ
CkvcY2LhvhqNKb3ude0Z76o7XYNQ2v3IF/83vayKJrI8bVGx9EnCGG7RyunEEk5d
2nkQVKCg5FU/Av+l6ITJPPK77s+UVpiDtxLsy/rIX5waWfvRUb8Uo4caoYnLmRl0
2ZUK3uTQ05g3H9qpp1FzjO+RAnHvO8+jlalHGwCaFmlE/5MTRN31LiXBQBGzrLs3
WxjVfEzUZ72s0MuadcHt4jxyxGch4V47F0WjavAz+Qn/rdDbRdx6a7S6W+CJWgZg
YqPB1rI7lgUG+9CnP+JFArFds28L9MifqH5k3ftWmL+XfWmU892A2HGjSSdyDjs+
rSfuUhzGBBb9Cxh3JUPNR4eaFzR5F+9/68NTPaykRyZrjOltj1fnyGhA1Rg1FR/l
weUqAfhy/EqV4iNAKhRpKJO/ZQMk4x3pH+bBdjlSPcRsX71w6xbiqvRlWDhOblTr
sPWmw4OAXlDYzzsiKF+/F/RD9UVKSCOrzpsjDV2kYhlSlBmoaCKZ9icbKz+PYExb
Ms+s2GY70T8SNGbMrd1sQ/5snn6c18IHyYZOJALmIhnswH7ssW46K2A8arEo2tvr
Cil3lgGM7ZyOnnmag5efmc1U398023ZStR+EIDSxdoDKgqxaYTIuuk0PqLbDC7HN
hs7j2OVEAtUERtpDl9F2AZq8SP+CJGF97UrHP7yCnDtyYrXTM3pR5SQ5G0Eah8En
hxIGDx/+Nz6Wqni91BII5632qhHuw8//eIeqARxInAtKUszH4Lw9xipjSflYRgG7
nUSk8+ByHQG9YgtQKshNtkng5SHSWa1Zp/3XH1C+mt+K9VK2kzK0tU4XcZlZ6jpO
EyatPMJ4bUAXEXX18wd5MdJ0ePpRK/ghuEJdLMVM4g7YJZ0oY9zgcelkfyNLWcF8
o3mNb19HKqrbXv0u9iM5csSP5Rqqh4qNXLrto5AU6usN5bzKqmDn+gF59xXLsdGq
P8WBERX0BqW+ZdDe8IcWQ2iF/fSQlBj4zgre11jv0VdM4T2BOVe5gSPVajjI5bGH
bc93mieVwrZAs93ZJ7Zb1CLhC0roho9DVwX4f31heLLAEVTGJHopR24AtULU/F4d
nNtfhoIGhFHI3L/LhnsjVcEyT+Ebv24nsMRA07HJ1wXGKraZRaWOEL3yi0zx7Hzp
CYIvjTV1MwLqkOrsB48TK7vxKuaKRyk5g4qRU0acRqvqD8Hw4IFIY8fCkkW+bnxq
iD2yI0pQ6KNcdgCWHRosnKhLA9K7tm24Lt/4KrC5VlrUKmatY3SJtXq19dp1U4lx
NvoNxmnTQW1kORkk4nLdZuN2TQSmA9ziJz+uZzJaAhtdek/BSTIZf6BmVe75vUU5
QXJgVkmpDMgeFmIw2tjuCbJ28EGthCEiEXlYH3WhAI2bu518p3TRqDx2MsZ4xj3k
FfjP7mFWwuUnAMRs/xtJGQafeWLrNF8r4L3+bg4lhiY9EqafwuMv0oaro46y297k
oQTfX/GTAlLYLftxrxCK9x5lF7beQHj4fOX56J9zWW9mfWlXLOddI/kFTKP5r1c1
N+SZvIbh6IVhqmmr/WY0VRo0uIAek1scSGlJL2sJWAk0g6p4/RnUGrjLSbYBm+QA
12XqANNKOZ7hxOtVBp7fuVXF3HYHTM0Sr2XPgMcA1quTW9+qEP6tA0hMVVvB3mSC
f+MiHl9Co3Sil7+LN3lhubcCpzVUOc9WRS6XAiFK7y24ambtQyIiF7jxIRjqk0Fu
3RmE/dSiR/BkEeBhY9Jhy4jj7IH82bUiOFX0+adikPP5+3O0Dy7NC2gNMEvZ3HWE
7nNvSnVd+FmGiOdwIsPxezFrh3SxlDIkbZNMxQe5vEGsfz7yjEyQN3vgPA4ujm5Y
ueLynyTlj7FOWI/pUC99peE3euFYaeSeaMwGrtJJaHiIEidkbOGuOhx1RWkKjFtF
pt8MnkOonNebD/Z8QAb0SzQjOtZAneX/4MnVb9G3THZD3qgbIJBYScYx8w35kozo
2DXgVbZPyJEjlnMwZIQXVD68esKzyX5/qVWv8c4w2nous8u1n1H8o7jMvIwgVpw0
J8lFpp3di7diCHF4hZTACvJhMcRzTVGwLXaQpudS8IM6v5/Xm6CDROc13pwXbC/w
eZcBmVSLnAO7djCy7v6jUuD4WRfhcLATGECbBCvjMUHcqgQP2GANgimFhoBqFV5e
qOJmxYPYvsnipJ1Vd7RNuF+8N5Qafw4NBKzES8lwb+duo38gelWGymn/qdkJsyCV
3ReuFDtDkhcXRYHVpLYCjBstevFv2vb94R9c3YFF9Kdo7XZLROIlVgntQ5fgOCq1
1AXulVoS748K1hEXYkFNKIF3/KaQHzZcRu6jCEamARc+iirTTpNlOMHh2OZd9hZG
zNXA8mBr4Fl2oJwzlEEUOC6OseMP2HfHfej0iVeemMUswUoGRPsRutWzZJ0UuDxL
2nB0NpmEciPwwxvbzQ0h1ATq2Ela8dd+UNagOvoJR9B7ZZgl01r3W+f4QcKZtf2t
N06Z0hcr5Py/66uGxt5pQNtuQyYCXizqSJCc4BmMnMOTm/lWolNdCNdBV+bL3HWR
ELYRQiR7jGZt9PjFrnTgDfO0u7Cqn9IXikFG+g+xhZ/tR5AzPqhbwx4Yk23FxXTN
Yw5J6u91fff10NUTxMwgbNLQ6pqiLcbaemlxd7CXV+ERw53qXjWEnif/I2iNsms6
b0vPdOZascXv7iKeO9N2dYW7TTVSapCt8dnOE3zkZP1y6zDc3+SKn4j3hRLpkb9w
M1JLuLNsBw7rWXdn1Uf/UA0wCnxrGVtbptKT4/0OCd3ylF7JlngmkyucSsVvOEQu
wn7f9ma2Hkt+7pw9BY6Rc56oTNPgpWBclShPn31JGyC/H7FuQovS5mnt/5VskhLW
uzxExL35+uShpQN8/I8M+FmZc010NDu7uvHwX8A4dcIoCJq6stu/uW7mYet6ajkO
fk0q5Z7Ym4tWPlgT8KQ6D24mDgKHOUX1jA+Pm2Snpn+caUTOQgqWEx8u650Dga8F
qvPorO/ugSwFrbkGhUTeg9MvXswCuwWGrYYhII98AkY2WzqOreq8FU9F4GPD8MK+
q76c1Ywv7yCK5wsCVEzTt+0lwKT37HOkjm48Cpy4NvmFDt480HCcJuFFMj8nPTdJ
OrHzhcgv0H8QuinxbpmLi+eVM2JeNsXOC4meCE5AGOTTnZboFY8RAwIKCnH+UKc5
b6t2XzQ+qei1QAnVie4vz/kfi+3K6UY2P/oy3QIqvFG+gFW+BdPwhxKkltibCuWr
HA+bJvodzPJaxhAu+FDAUu1Sz46nf0bUJWqMKkLQo9OZffvl0pV8aC7xAi6IqTGZ
Ys554P4p1wT/L/3V1X6ptuQu7g6hpTk7eJdyy4WiH2PIgN8PHwzFTZpWoHDqXZAq
6fKK2WiK49gZnjNic46gXtCsLiy3w4xjZZUggT+GwEqjmOFVpMKT2AwH4Gy0j1ck
dSmZJxmFYTIf4+7hCwTENcEtGnCYUFFRZRPS4rqCcJmAJAkD+qYZ8/xi4EqJ/Orr
EHCRfd1c1u7VDEOzbC2klWz1i2P8dyAqAJJETn2mlWNlEaK0xbE5hU7LgfRs8dK7
4wwopOUO+n2NLmSEfm8hQJO8uSm56PIgufOMTlLWg/HP358qtikT2rlriGord01i
Sa/7R5RO98NCVShlU1uiP6fsM7wdU4F3FSQ6dRymbVIdvc0CvjkF+SWFQiJ5+s7c
TWEDBSC2Qm0caeQR98qkeRjAKq6ee1FVOoGP8ObWbXlNFxz+OzJOlAcDLxwH/nNB
Su8+YD4EARU6yiTJ4JtzG/u1kMJmnC7e6lCTo1CZ65FbSsCnTPSlF3wtajnEZadn
hEAnhYDHg6ExcflsmEcBdBXmF28yYMRI79AoUZtm3u6Df6eHbMsUdWUiGD7+H+x4
vvjTA10urOnXOS9jnD9XAMWSlfCDAm6FLzTxMzQAfSmqTbGNsgYQfKnk98y/KOfB
kezslr+OniS52G0p0/T8Cn7FKuoNUnd9w2DQYlKbCYM7NsJ19bs/t/GFpAvk6jM3
2h3f2gCEuByJvwXyq0AFhh4XWtkJUg4zUqIg45EDym8re78F9EQHdB+K4MducxQN
flxPAxeRsY6GWcCjwsQhXc+TgtNsQ5cRkgp3bbNpgcJJIVIBfPWsK+VdJolAeSrY
dhcV7DbjjNmaOhoIjqS/NiIcLd7B98PCqickylLzQum0nP4CP7bJ14eQDcOQI5Yk
A8Y++ohVvpaBFDS0Mc+6vxM3dfZBr4ZvcZ0F/q8vd7oNVELtvsxRfM6k1ai6MVc8
fcPUmtFZRGXUuQ4R5qLitR+M7jIHoxgpmHSxvq3Wy1eQ272SVGcHtrX00vSjeiZj
l9NT6k/mHnywnAFuDQ0vcMGnWugFQ6mwRGb/1yMrj0FjsQ6CO5vI6MOK1fnle3bQ
8x+tVl51Y4vwcEbOekbyLJb7n9nyijgKL8OBJ6oCbr8xLcLwCXGR3VzFaKkm4qx3
dsYQfCZi5a5rzrPJudsbbf/yUjMoLcWF4ZVyhy8y2SEJp5nSx1xvIzBcDejHFLde
x7eAh2ysFJw0VQGwzQ0lJZPgCoYxXvk0EzBZUvO6Jg+fALDKbagGkO3AFzu4E+R2
DsElnzN0sdk+4tZ6vVc2TbGlaWlr2F5Zkn0lLgHWAowHcu7EDTe+0r0fpoJFFa3C
bYEW2YNzH3qcGrC8gDssFrxg+BdAHt8MOcilqPe3AOB8fnXRl2RE6k/M8087R0jj
bNjYwsfyiQoIX3QSm5wPK5f1fIlhIexcK9X+xF29IuIcFEl5CUqkMfT70KOgaunb
qFpiEiS16B94NwUMOo51YxZDGzTamdw/4irw6JnoTZtqXl18kkfTKJNJxzi5d0/8
3YiYFWeBkfUYLv8dAf99MFIIcBKzP2JUHHsIHedoEUfYEuwH9STQ716iNFq5fDtZ
hkSmqh/so9swB7500o0sPl/y47306Yt9DoV1n8qFkv7hHRtNY6lVSRV+cTxvQ8cm
ACs3A4SxmdXoB7bHL6Zb+EQHHYrLnyhgj9XU+C+9k0f2ancJ6hJEcJrEe3+RXp65
bPvRhUYliq1BxZ1andLO3zLZmx1qSOuG/0mjSRay4uz/Ci1CU2ijDZ7flTyLLHRI
MSUPrr9HWLUX5V91ay1dfYDRFNeQSKMG/I9jhYqLF/PNcRzoiUtSrgOext571Zf+
bmsMvua4RypnZGlutHKyBcP7FzjtVNhqEsyUQP4vV5bg4m+lp5VdozpWYPcb9sq9
WI+4YW9uiL+gcpjfSTi6r8ONvmuk0KC6hWUSQmrOcdKjL/RdLcbx/w35pitKNxQT
Dj1OHCWkRP9PBd79TF1bi8AnL9RTxKsy7FcdUptXSDTGLcww4HHykykg+KOFghRR
bKeQTK4WhQOceCRdmeQk1KaVphxBm5tSQJieuY7G4M4nwww8aLvlkWYKm8u53BuR
RJI3B6UDLk3xBeARONvmlOf6Rj//duWo4ugWhIqrHUBBdqMbso9fSd50pRGahqBZ
lRMiVnj+ECt6ME+M/9LT/XXv/8lCYcLE7zPlGfZ9R7DE6hC61fc4BVZTiatnmSdC
VoOTpszXzquK8K9BKD/OmB6r9hEyhZSDjHcR2QjG7ukUGuia3lW3FfvIDS6aWgTb
/QyZ4BT8E42+teiptAqCHfLh6mocciKdrLsFpGE4cV/3qhiwIY8IrBqj/CdoT7XS
BdKWObnd15EoqNA6AlDBQoHOhHuoGyzU756TCvSdj15d1zjwaFR6A10AjYjIX2KB
V3u7HRUY6fmvpkvvMxBtixYRB9g9cnRhM5kHIK0QI1MEuaDX78krH1kC5/io/kus
8TBAEYh0E+ShD68em+xQ8giyj+5ibWcYTuHLAcoZWWhb42jQYlmEpAFY+XV/luuQ
D8tYsxnwJiDkD21ktErqo/isyE8Ah8ey0/Atpl9C7GAGcz5J2nACuno2lElo4Q4O
DPtExmWOCUEmFg3LbE9i+aCoPcr2/5g10rD4B00EnhRFln2d6nEIEQUkZkf14FK3
fxJIdjEUVxQax6LDEQB7yX/V6aj32c1XVVPt3kWbzk90RZ8WUL4+tMyEu1wuvi9v
/qJKITaYf1bnco0ZRjqx3Je+BAMh/Pg+4WQE1lUYyYwK1inxpPxjTomFgYoRLEUv
Rl26qpkR6EqQmJkjbAhDsuLQUv9ucs2lTtNBjoLyxpO/GaXkX9q+DvI5gn7UP7An
m5bGHWRGvq4WbNBb1+MdAy62ZI+XYSap9vjGMzWDibe2u1wLSoNm/o3jb85pMujW
y5yY35L00/rOjyFPACTyEk9i/OOyHNUfVoCUEUVmZ+Q9E/jp2QlKoHWS1hCa1/Pj
rmDHjjJYH3SPI0VvvhxWzgDB713NtUXhi4EtiHXAT6Q9n3q9EerbU0EwsLkalg9W
6mXxD0CHL0xLXCFtXB6pq7qqVs4Pq1dp8qtrOrWn5v8oAStvOa1mtoVORyc/Ir8W
UvokpB6rKvxoMgttjbfz7/Qv8dpgbk8TwoLbPSJE6B6qJP1nhMFKdrEAUXPrbxsf
gXC7D5uGnE+vdSaL086vZESFCw5wfWW8UcmZmZ/O0XwIFWAbDjsoO0pp2cncA+t/
taKTTfTTIR5/EkMqSlnxrvYqG/U7c7U534Tf+szoycYS2YzSUUdYYm8QnrJ0BiYC
+nYhtbanI4Q/zpfxkiddgTAEsJnBzBz9t/WPVXSPsry3C/qccWfwDt/KNkD9fN5c
tntlZoxRf3h+nebalvODKYAlyyyMObWal0mdHKZHouebYpiU0Az7EqwZoca03yUa
U7XabfIyGuYZB7Uqb/obnMNQKJ3KvBlyj+9hA9LP8Htv2cNRero+KZ8JhUtwsXUq
Qpc/14TpqNde5BDhFXqzA4pGjpT4X/UA22Bz0cWqq2InFuvmPjiNyAXDjWIa+Mfb
MQJQtDB2EnfmOMnv7+bBUCgvf6Kbj76WzTbavpkKfB1I/jqfmOuARYmd+CM4GzX9
Tv9/4/iBBLk+quyPmovn5zpRfNhs47tziirw+RnQoViF6MG6scBf9VrH6PoxQLxc
9LdcxRGTacqyyaRU6kJBD/EMs9QkvzaDc1extoscY8GGihukOReuCqMqP+0sotaM
sNWblEQQUG/eB9SBWxPMCvVJs/8iUT4If8qRVTeFMlSt8MZagOFpvI6bTx9M+GkE
0++hecZ+s1Ix3Nm0tPAZw6+TlUqAJio9eA1/wLq/3Im0Aa4eOEh+C1PqHDet5rSj
iy4N6atxw8IP8E4Gyj+FHVCH68KywaSMu/UJ3Ens4BJ6NtTv9W9iPb5r5ssQh6wG
IQC0rfUk3cX67IdO9u2Nd1Sd/xxoCOSfnDOaL901WdC12Roi6PyKXuNjZtBJOcm7
py80zIGa9XMzE5Cosd/d9U9RwxRjz6tlWgOsKPl8No338jkb9Z74ZZV4MA+HF+Iw
l1ayfxIzOluFDFZsw2ARuzvu+aioxV+ACcECN4xiqM3sSY/bk+NVqaig8FcrzX3F
Vz+EvXMA3LP4UPGW9yY4Xl2qpGD/cgqpAB01SrqgcViOGsfPjBYW1so3XF9/ICWR
zabWmESMyA6V+DZcUyBPLWzIPwWfuMpkhc3eSLFYM//Rwhgh4AqpQTIaX4VseE06
cfpyglw++ES5X3u83MH/rmv+kdyH6USTCqouhkOEzgByEwePsatQaCpe3X0h47RX
eZrKZsFvyqH9NvAWOjMeICBT29F8RhxrSR3XKfHMP4+IuDC7zAlKK4ANcwV+Mf3R
dYb7MOkS6bd+kNiI0vj0LOEfk5xekyGpS/c24eYJBDRdiMNP0yl3W8cI0BTr+YWp
UL69DE3CB4KK/tqS0IGuAfhLOxXT+23EW/Axo/43klABtAGtSM+pk86upojuloVn
rK1j+Cii6/EUzZZ3SDm18yRoMip0cY0rp5tCqgsV1I2fm8u7YWbd+AzLhIVKgsBa
vvZFhJSUHJflhocjJMzpe9ENSId5Pp23mVHaBj4DgTZX0zslhZzXFKb9odVXCddm
VT31A1WVR1tV/x0h3D39pXPR9ILCpCwP1Mka3lgNpc8It9tQddNnDGaeBE3gJPGR
jk5y5UxGpUquYoXCbhoXNRi/iWrJKZ/Nzf0yC28fFwwLx1lQhDhMkPQnRY227DWC
z93leW9Jxx0zPfgKaFM7EW3JGKcecdixSAkZ2GRowNv1zTKgjK9MO+F07E1LT35J
RPtu3g1JW3vrvxQrVX7eSZXaLsL61/skxJ9YZtU4JtXXQAKV7Trw58lkU3cA/waq
9YTjH18QPTKgPDvDtSjNJrxf+4Mzii+Dl9GsJ8LDg3YLY88IsfY5D6VgfasZTc9A
rRsyg5wxBBj7u7ipIDkebxJ+sriMj8py1H0eJO17AXVbPl/qbHZ8+mbKyOdSdD7b
TfS9R9tiOIIocQWh03BW9dJAv8TOEIwc4bkCb9rFdRMrUsj21qSxoWTY8hzp2zV5
Y95vZnBUSwCIoABhaGSV8IjjCPojmmQAGkUjHUR4rg86qJa8HgOZ9Du+MuoqpOUw
8EHJPpfJ4GqXeHBQjtrBA14ievARiQPaVVjjPHbf3rg000LGx6AgRmT1px3NVLeq
oBSCcZE9kEyf5kcZlLX4rgu27Yx1J8I4qTodZ2pP+pPFwiviS9P3cnt2pX5z+GFz
6yhDg7NoEQ5KaMSC9AxZ+Ts1umk8OSuPgKyCP93Pf5fxS2RnfRPC9knNIHwPZ7q2
XtAakDgTvISWzafXkAZ2K6AGFlcoL2YyjOcHBQ6QSRtwsfR45LygziixK1Tc45PD
jGj3eZlLhtztWgIXlj7iMQACWJWJHt+Egj3HASoYZaJH6C4eFFACzgH5T+oqGKW0
MQ/hUW5VktohwBSKPHNgH1RMTGVr3y9Lifjk36SI5/DHKs1dG+1umsPcaL+P0qX3
0b3pEgI/mrOnv/r4kxZ2FDSFufLp8X+5ooAz2TfA4p5P82uj2lqXYxE4Vvdz80bc
4nmcUcsSWzsJPVMaXttW+ti5x19g7vDlR7ZFPwpxjgVZyORcemRCocV3Ie8y1Wv2
uTnIhtxHQG55T0FkGFi0efzIi3UQpQ+y9SlW7V1zg2Vwd/kInFxJlN0c0vybYWOl
me//aZGr0JWkmEsWrm70BQRvvN9/NWWX1BHk8hi/QgTQsTUup+J/uol7spf2VwHC
MDbfX2mbhc2jCwZTT3/duObT098ywra/Z6RPRkC/sqRq2NK9T3gSZA8wVj5hj+s4
wIbCcjrQ35h5j7wWd7WRFrG4yjzx5rX33dS9FGuFmw9vs7yFT6ul/5B8yQzDtGii
lllsMwDiPn3AKx6l46XVaNSUyPFDEuC1Bl84KPWxpnaf6Mz3/x/fGuC3owwxKY+P
5HPSbYCVN1brhOdve8+7f7dXuRCe60lET3nn14jE76AKCcc3U153SrgzQ+B1nEKW
qqWIz8AeztwMz73nf37Lis/lYnIqMctFay1clUcQDdAYoOWiaZ8xnEijcloQsuzt
fgudZ1bJgWQ2Jxfc8wBIjti3EKcJyh1zMqG6M1oOF4tkyTYG9YIW34fHZqI2v0z5
nAqHKtHgmu6DKUD7g8wEniTZ0aR9okaY1lVHfMPQN3Z0vGY0l1lhAPBdb+p3FnKa
EW4Fwpc0D8On4XgHTG5mccoDs65GDNBH+RE4Zq1hpS2/eXuPwAxk/8i9JVBVLhkh
cRf03tmH58RI2QhRVxYUTBOZMqAEROWt4BDod0GJIa1Fwn9E1Mp7ca4gH0j7UnoX
KoBjVXPuha/2Fyczxd6LJ6p6t4ii36PyrTzXTt/dj8yGDo0AnGfzFmbGJkWqLc+O
7nfj5o/ttrw+3maXvF8zyyjtgBhGwMfrnAlTZ9sYKK6e9Qlg3pWwpxDT5eOiZReP
d/ZDSFdmdb5bWpr5CiKvaXxQqkOjbc90doGbOVRkqMasY1TzLt+jiSTEED+oRwAt
L5iSuWM7k5K755N6B1UzXbWGJHsvQJ+Ao3UUyJyA/b3TZlYEwgdLKTjs6NV73bgM
HbGean1Cjc3qpKCpJD7YrrESLsu/PJiypr17uCXNs8eCG4uIA9IersG4CJScbjyd
TyvlwaT36QdKAxcHjxib6L/xu+lHax0FMCol914pBXdKn1NdfcyWlNSNHG95KkNO
nS7qoV3kAwgnOLA1St9I18C+2Evq+icySrZcDJ4cGwqn3YjR2qvAlXmatN7WY28D
c4UnPJ2n/g6bqZmNGY6a8RdH7zHmIsP80LRo8potnXgD8/LokMuM9oGV6Oqk41Mt
GhQWXGJs7RoyNDmZaYC+5RRrpz7uCUhYLIksg2OTTqnKCdmR6Mckg90lQiPG+zIB
8fFvawKhWkB4Vd8Vin4+To4UKRzEsbwsY/mAbT50BswnyPKMg4LAbXe88rBvcIck
xzYjxQ8owXRCEmWeA86AS6mtDigOpY7w7mLvmlHYk62hGtg7hxTzOPdTuIso8Rnj
mOUVBPa0yNcuTyETDhej+75uFRLMjBGgThD+61gBfnKPrSSZKYUl/L9+av7eu+uB
SkPZJOO2ze3EoVz6V7Pv1JIEa2kMd9+Co05YbQ6eOhbwLHpYsi/huinAEu9l/Ars
ZN7tfYsmnrtxIvpF22XIGnnS06yz4U8RhVPLdUSNvwZQudB2c02WktFtskGUCj+U
V/Rpw73D1nAF41SnLI2l7muChcpXLYoUUsokwFUvfmUw59hreJdXf/5nn29gA35g
DzMCdWN0raQX2Rg/CIQXHwIBXEKLdZv3/LFazhOmCKFLqarFmttpyf6NSJwUf92L
Pbr8LZ43wiOoZ0g4clvz3lOLIft+/T3KNqKs1cZ/4BABBfuLIfbSkrRlAW8rsLQo
Ii69sjOP/B9Fm93OSNtzqsrpwHr0WCpFnWlmze3EnwM8uxUn0T5Tygnp3Er0KkCu
TkHGDFmNp2PIP4WHlgeHP2Y8ef1n/qQ8DYNd3hVNfcv5Q7KVc8nZxUchbMrTvK6Q
MXAMrOJPUi8E7ML90e6+uZG18qW4/uS4qCDdcIPxl1KV5MSZUjweZynVWbpu4+kV
y01yIlifBQLdpMF5L9Pu91cRHLPjWydk1K8k7r4on0J0Xj2hLHFuqy7kdfth2Xfp
0HHSUvhx/2fKSjCSWxFpDIZVF3wC7XpgvjqpEcKaatT9K+TiyaHKrKlZJu1buMRe
O35wBTCY4efIj/Ee1CZGWZBvNnw2zKPhA0PuCRFm0rQ5MZh39pty2GQu7OdkM1ao
m+9ALYePIrxO6p/cq/0sp6fyORGEFUdwXJC2HfWpDvSL/aGPyF9djfQVhRKQB0D2
0M1TYSuLXIsQCb5NZVr+SFzw0C/l07/fIqgLgugLgPxtBDglUzJpQV+P3EfxXZul
OJafT99VSSBTbKp+586btCuh2bqTHAPaPEp5SlBd98ol1j90cEju5YHvMvWxpYm1
Mkf3Q1pSnrFo2FrZ544KAbL0LjHH1Vj0jrTtSrqWuoSU2dMnHj/noulOhSNiBuOt
keAyj3Y6NMRUJ0eb5tPRfCGFeitiyUpE0P9Sm3Ed/08HT5POvEWmNvmxY+2AuZKH
K9iUrxvHYV0s87lhaFRmZ4QEBcWlmB8UREISDINVbZgT/erzS2DoZbLTa6/Yp/ap
mGT6BTtIWJq8REHgTnFkfMMUoao6uRFrbtqKhsB9GNjcOwDcsRwgDvY6UmzJq3i0
1Wc9F1ZCoNuKgY4OqJI1ld81VwtgkXC1OntGn5+GebE8ZmbFW/XyIs7oVx9+pN5D
Bt42EffOgyMLoluR0i1tJXLlcVqUNm2QfWbOYtc49Eo11QVpZSnKhFo5qI5dwE3b
TwH69qvz0V5A4+/wd0LHA0gQ09/5rtfByiGjkvbQBkeON6VfjZMTu49REQtHFgsZ
voplz4/klcDbVgr/TW8HJYpV18GzXrf1zz10/NDvTHg7tnnAZfrwQHPH5RmTgKWI
pdTpMjCmPg6PiW/RTiREfzQXr4F+BNgmUdrCf44HbltrCV3se1c+FRWigdWyqKeE
sa0G3LutRKwtkkR31SKQwmqW1gvB88ZkJL0tNW+yJuB17y32ULtIigh13xinHhxV
3+edeEwFl506+QQfEbwN5k7sLH6zT/2uDrt0LeY4bu8Pg20Yvf7YN2QirQ23fln6
t/VROjLXZFWfeaYwt2+4PySzMhDqyKEOFVay3NvwIM1vQv2YjsmY1yaVNxkad7Nr
VNuwKLJ8NQeXRy+jXuFfVgptRNdV9yyUXdIUQAMyCIdIBYOrgzG1M8ewizNldbV8
HhDIuzHvXZQr5m457EP8e4zysoo43sPaOSO+7fQIdyZ9kinsl4uc4Uj4DYot3yYH
bib4oS729vFg2gCH/UfGsR2O91mYTI+FQDRlncxP0rse1MfQaanJeQWaNxY8+iIB
u2mXeZ0mspKUmVwUPweVU0yhPLHnjsNIsAk5fKCdmkUcDOzkACinyrck2vQLRKa7
FPs7pZu1yD+8pNgxc83vOkojQTlsYeeyU8xIpvaqAzNM43NIRTvMwzBEj98dA/B4
dUsoakRkkXbjbcpqo084L0WEdzXiOmPW32HELo0rOtE3Nsveohfrxqaq2ezu9tjx
KeJEEY1c2WE2dZoFnf+rg6COd3gRPOqp56hmGR70BwiBEr45oxuJ8ocQYvuLkAie
Yd0y43nRgOO5FfkPdpjwznOvNW2IbVJ3m3+D8BCbBz+1eZc57l2AOWzwbWSlzqPl
TJFiSHyS0a5eBXK1Xl98HO1usnYOoJXvvt9FV0YQUdyWzhqvJVJkGKrWXwAoZHq4
w0TbfykDfE5ATHdHHUiyyhmszIzNqVTkrKfQh2irhADvf8ZY/AExzQCIgh18YXAz
23O6+UcQb8qvaWphJJ5zfumS+qcYmMqbWCk7cIrxcXhNcUfYvu2M9y/qSoHVkgN3
JCxpZHK54ilQ8ICq6o53Glvo33iFSNlpZlotnmxwSuH9Xol9uNtCl11A26jGp5J5
TxU8AE4qYULhRBU48BAFqMsPX/dSJrHenmTimEWiJH6vD6JG6vXgTpy5JdAaCaP3
YCj4patVPazQPinh3LQRu9IPa21N1ClNf7CCIIiTgXRKms/RdWoKpKhZU/ndBfR8
TlwwCWGlIG7PFWcH/PCGDaokr9XQ+r43u05Wi2TJitANGwc5RP2lR65xxCM9Ho0k
d+JwPeChslbk8zHWL5bH7rn6yM5Evl+OJb0AIXQvndpoNLXGBm1iYjIvjuHzhNqL
G3LAU58mfMPhOT3tijhjky0RidtmI1HAAkc4+QUTB33GcM4eOnK8kuN/nQMBrckF
47ywOk4S6/rMnNpuS3wu2QfxfrK5uj49/ChdPjpEcWRhoRt/RdPTLYyUrKbu84Gx
Fx75Xl9Hagp6QJDq48zzovUK/2wOUOzyYIPc0XHc9Dwo22jf//7VfebEoNdfSkOJ
J+WxYpYSiCAQ0BE4jsQrXTa786KSFVlmDBX6JNHrxHFfcuG1VwUjc6aILIx+Xq2y
8b57KEe10WydqNTf7PTHuT7JyCQddg175j+e4T08GMHozmDWRB2VZaTT+5yi9NX4
Zz+r0hXrb23Dfo95adSF+60DW+zptDS9nAdFacyZhak300WxRoULPe8+/JnVBzP8
PWY9MPxqmPx3Dwr87/YN/slag7d3ZnUrtu4nGBEuZjKOrOPOcJJaI6qROL5xt873
cdp3gZaFTpPR/VH/YIiduT54715wGKRGTdwVAz7qLm2Qx9Z20wfqyIXKqD+4AFuc
MwebpWHcStSrPzcT4hl+HbKoFmOYIyPg85FA4KDlS2/dNKTzRrG+sj+NRwRsETSp
tAhFq6OUPjEs+1giSE5K1pJzGoWb9c48wJQDzTVw/u9g9XpyNrTR4sEz6PiEQ1FQ
/4uamH8HVhjuElZmrYL0qrF0AcumCCiVwmJW+p03k75K+uBfF+Jc9MoGWYjAF2Bv
5XX/WaYNzPFzWWThOqik/6RX/K65ERLV4dScVR1kDUZTzYlLBSwkUhWxm+HmW97/
0unuYrxZ5xr/FBQCLj/R+gzyDzGCKpRelmGuQlwbZKH4vzDpFslp86d3CaJ7csM8
PNeRBizk4UIKpjYI2Pni544Occ+djvNo05fR97dKWzOBaEhrLHXXeT2HyTFel+aR
bpJAVZFltXrgzMuZym4kXngKE/xxPcKvBCGymhmSDzCOh6xdkPw3wuh2qx9l1evP
AZNFrzgHgTQkN9W4jdZKHA9hPAUE60Kup6zkoaxNyqvn60dBT7/B+FnLkuOvg0Dr
xgrrfdzQJ6WSwYNBZcDbJE/lCXE+o0naaxoX8SOnZcEvzIQazr9LvipdQWFQyFC/
hBYxgsdgnjCeV3+ZHfPfkC14XyNjIl+WzC/zdNGSPqrOgjdh6FBTY2mJAO9szP7O
qCP/l5ob36x0ngW7praPqSNTXWun0e/w0IsIlHKYfcT8pSPHs+Se5xZsftKxtOKU
xyq06r0GvEnAJr5dLLkZlOhz9GMTBmwaTFm+nhbQIYdfqG7tLLjcDgqRSU+jq5sv
i9CE5sijWOu88KuXPq0zi9vMxxeuQA1rQ72/yWyajG3nb6aTUhGOLYkqO8PwbFYZ
PcI/U/DLwCTa0PjJdHDJtQdIsN4hk2OPhIC+E4/PgB9ggScQHG2I2YyhBV67VcAw
DC7+EW9jKFRdW1lnXf2mw/S3WgVy6rkBWsnKvSCfzYfCCRQcDubDvhbuY0Z/Wsgn
WP1xiOROTu+LfmGiMD4f4dF5R1Lgd0jkz4n9syzXJQei+YxhofOrQuKtMYpmg/Xu
CdOkRNfAZxC8r1cgO18m31AF/wgUC1vG6fSHqUpULBhG8Uosp7N2PyZgIq1P5IsP
6oe4pl7hlwFASu+NOQ+vTtdzX0LxAT+ZSVgTHsa03jieXM78H41eEcdbVyw0eNAn
owVvSLSNwh9uuogtamr44dKDrevXQ27IaKq48OlX8rXbzrvI6G36rRwjLjrlRcd7
M1kV9GMrh4+xu88oxZEUA9akjLmNu5Q1wEusZ0NZQEEfcCKtPaUuBaPDu0FEhr7y
LcRx07oTlOtzjygdKenUjmBhq1nBWZfeGTG5kzSL2scGi9g88uOdZRoyR/epJoB5
nFwhVhf+HS6F3hjQWzamYpgrdOb+myFG1ZwWMP+KxfKK8sxV+hiiO2ZdcyQcVBwz
uBlFsQXIC7Z3NF5vhUg8LhnsmJFyyyVRVq41DO5EhaFHJdIJ0MfyBAt38dzcD9yv
ifWd82+I+cGMlv+gQjFmUCZ8zAOU2CiLMLQnf4URePQ1VaOhhbiu5axupa3PXaCS
sVCe+HSGitrlyIQgACcJZUvEFwU5vpOkGlO8BJ2h/B25SZbAx0KqNw1TfMz0NBoP
IU14A6NuRcV3U8k7qxPP4Vx4+/LvFj7OdEVX/pOLyczHDD+GD2Qq3TsuMtg2TsT1
rsm6X1eTboc2hnMcOiCj8345eme6gyEjHJlVGj55OjbpHGnUhzN3mYVflK5eYujm
iVmIKr/agm+BdkL5Jzq8fqoBdstYYnyisYpKuAjfhrJ78e4B2s7l/UZoOOIqglRl
l190h0PgX0DdQkvoPPhVIh4gFEwqDsVzM9Jth6tGMr9LPtxazrfA+kJ0WPtuwb7g
pE3dUntqR6N+9UXsLcZqM5RYHtq3jJRX+T73FhtnmVJyg/l2zuENg9iM2sinlGrl
mgXRxicg/mMuNYR9Yh7SNmgEipUhNpqzkk6gWbjdCVy86ZKliUIamc0MQWapvMFO
CMmXjXdrqzRXacvuoRogZFQGAzUez9vIS/5PFeW6fypr/nHrcb2r0eOW/ddle0mV
Qb79u63LzVPDsT9k0CZVkmvc2zgfhDlIrQxU3GuUxElEGQhltHm5r0LJU3AJGhGV
DVayLBX3vQwwejNpIgBdcRB33B0/8+N/80uOG7kyj51dVD75SFTqeBVt6W7NNHMH
Lz5BvSX8kOHUN4hBadxeMAYW5SRnZraJ6IsJDwnZAv4PDeHygOH1IC/2jvLqe0xn
tehk1IIspBh/2X1RD0VIleDq0RJ/fODHg9fjP25MiwMaTDRElM0xi4bYt3P53uYo
KbW5uUOByeCOXAm66V4Mtyu6e6AX0lgIbCXPVkZcPYp92lzGuL+WnX7GGM3BWArl
qNZwTsOg0hnF4u39/FH1clRbbzZ7ezUsMoLAgI7F79M6/cC0zQIv26G8KyMwqFV8
qXa2z5OSe7nMRWHJbjOcDh+J6Nf1E6S9JUbttlcqIZV94ayOU60KSNUO9yuLwXVN
IkavZ73z1Xg3O13wyx/ttbqPOkKmk7Nx6XLGVaXv4wxrAaKnN3/C94DUq+aXfbiQ
N689B05oARL27cB0NtWJQV+7aInt1OxNuydum0uf5eoWUE9awsT1BZADk53RG6HK
Vjom41H6HLfQNf7wweQ2h5bqkD3ZkLdiJgq6y1n0flecr1sUlsLeJKKLhpZ7X0m0
8DV77hbnTE8Qur1qABz4Zsw8yXLaA/XhbWfm59eKGJxW0PnSKZtHjLbErYkhbE8o
tZBVuC0MJ3dzVqJeeHxJ+GuBQz/SU0jgTbD0xpV3AfzthuvJOA6LvqHHRgTkXVST
E3jh0zVaq0OsjWL1mKPVkQXt6obe55PsCdcSWr3qWSYYg9PMjjXUk1IiVUp1R3ln
P3j8LtX8a4+WoBezRXrx2On8qTqVF7CPNQLHf64NqtGbxDfzoldpGz2A0E3tAija
FNxWEWHFvVjEDF76Ayg6c4I2u7PBufHWZDWzD0b5MtObQEWt9M0aDmFhEsAiame4
aqSG+tYub2M0okfXH9W3QalxHiSXQx9hatmYwjpy47FmQ2XWhnhN4UbvZqPjn1Cy
3X4Hc5+Ui7BWZvz7IMkxE+Kx0PafeZ4GV63c3TAjVZ75c1u8Mm/o56/tEnLoi8q3
+ldnzeVtOX82zTTV3f7O9siN+ZPr/wKHjFhyT9oW/18zm0swNoew9VN5PR9Dle4T
LVdKAesAiRLs5YL0jwN0+4SdN6sXwdUgSCHpChQ01cm305kXguNrvPAKCSUJ5MCF
I9CzO+SovOjNh04HC48bA3Xrl4TsNEhSgYWWC6eWGnyg2Nl2OgStpgGGF5aI4U7C
whdecx5PgQjIypGUIHq9Av8iFsEol0kKbYfYrg1d5qWcI/7BK4rrPMr3THQXHynl
SkcTjuAJXtoIdR7iWllm8Seug/tnWUimMhX8Ohc2VkBDdf4REzM/JAqGkuqhBbeT
n9nuQ3J2c6KZ6x1GYYFSTv2H3nPxgLCI2DwumYvyreuPyb+GCYPIX6z9sUzW6wIY
BAhBhA1SKgTG8kCwHidw8ap3ePZmVmzYpQks3ef5zepVQLrlNTdAJGDEdRc2piu+
JyB15q7xd16ezYoLDmk9ksk6KnUzNs9B+p7KTO7vz6l7+tJpvhovD8oMHKcsQGTI
GJQSwWYHJEpMuXpOtjE9F7n1USRsDWL+9FxSKDSh2MGmLTADq5HN72ovquIVwVhZ
MncTBAknrwWSaplhyuDo0nduImf+BAuMPO37VLKJmPVzKlY0lUm2ROgi6MmEeeUs
C3TiDLyBxIDt8zphnQJ7cF5WBT2x/whv0uM/ljSPGA23ujT6MW4Doloj23da1EVZ
AcrubvH0C3e207V3CxeISpDsz3vYqdMbkJqFXNQu4lHhHu74/dc1fnkF4IJAYdCG
0vyb1fa5kTLnuWV0JHtpdsvjR+Gv+5NWvpSxua2F5aYOIJcX/kwZHZskSXT2P69s
9WARCRXRM/3zZNNWdf88nPs0Y8ZUT9mMSB+AlRtHmZOoVIVI8mkyegVCyBTpUYDc
cbRNi6pCqj/0f9cCKPu2OM/ciJ7xjSc2rD5y7vS6xGW/VaInFukX4EAau4C8VRrk
pg7LabSnuDNnfH5i9G35oYI5pZL0OwK3YaIBZUzJer4bjf0AKwWK3IYFfH1TC/xP
lJCAct4P+Q3+L0ABLF5NB9fa0Q72px/6xD8cuawnQ3iUX9ABiJ3ccHjixn7dHHLb
jf0S72hjgtJpn4fyB8ye1TwHT7nJvKONQ7yyGss8+ss1v35xs9E/h2QpRhl/u4Cp
2YmKbUURpNPfu0yeGXqeM1GNQZde4rqI9hcNILCjZ/on9bgiApSYSruTvEhSTycf
nhTLdVpWC3tw066zC/JvUWciKRSaViUJ7hm6ppEy5eGJ4wBg5AkfmCT1fLh/C7Qb
8WbnP444zKz00Y6rkQZFQD5k0jxl/FUoy+gZN5wnlzOuzZOm95yLedZqQ8TzC7ZV
Q//tD2yW88ZsIiQQJFfk1dn+449bk8SakpQPlqVLgna8LmivBV0roJn0ILM18RPm
D1yYmw/gxnTyoZeLxUQ+JSm9USK+MYqsictrIlSE9zcjnO7rM6Ef0sN4J07llqig
6bJp/0YUfqcALGbZR0MsOWXfxyppFcSEUCcvhGfRFT3m4YWaFWtV3ftytiUh0+8p
AV9Jaz+i2Iy7Uy+F7yh9MaPdvMWIl1zPw1Vz+ALsi0jjfmii6P3Z/8W/ahe3PNUl
6/hDKmc52E2l85TGEFXW4ErofJa7S5cZxxFyoTYwQLHXZ0o279fREKkDU3qSWvDE
GoCXTrIKuHMj0j+H2fjsLOS3nsTETzHf8BWxqKMsu6b2FxOH0uEGw5Qnqk2oUjCt
RHEmkTSJB5bwKS0x9EEsgmcR7sjyCTLs2iG1V2OmR1ICbpnLZ1P7cxBfSNecuFSi
ZcMYe6ChMWeFfFDYRQWkmnm5WzOwPFRfX7hfvQdkNgPGyO8PEkdQ42eQ1V3Acuvp
UOalGaZ8yoTh5Gq/rvjW9LXj6mlZE4IgNKCQXcL60cnpSGQ0L9Y7WdftYb3sDFhI
abTgEiEqUyYAqzvT1R0AmxNjry4DGIWLA0POZ/u6gt536S7k5goE6Uf2omQjvQsJ
/TBpDQayVgHgohl0t6OSH6eo2mtLERvlambPT8N39xiqTv3EIv9HNSK5/uxYHn1i
RLCuycvYvm2kKxCP1mM+nAcGDKlXdK+aepGfo8GmzxtXNWITrx9PVhbfajfmwY3n
tVZ8aXtdD4/Xl4dn9df2QAfezNheme62GOya1pgTYmpWTrZUD5pszMcDCXBbY9eu
zMRTaAFTt7aRDqPDNHBKp6OyxrV74e21qwbNxT6adkQqNRgDelBUiZ6p4CEG/F+K
YBKA+wnTabNA/A7KZgekLp36FP9SUP0SALAAQMGFWqosim4piIWL18rc9Twpfc34
/SsjOS/YSCb88EnqdBhCDzsLnU8Uz2I8fn5E+CFZDUC++CR66saaxsLnCeJzNiKr
RqS0anrBHaAVLS98qzwQXEOSXryTyCgdCJ8AoULgrLVbZi6Zk/SAsl4udbZiEypi
KIKr8STtvVxuqMPH1uep4bRwf6qCz1DL6x4c1lZf1qv7kBh/fegmMqFmicVmYTXI
fYtt4b7mf+Qh1ao9yF7cNZ+iGhSSGzFeaV3OcxWVeGVPgwuFtndjpZp9OsBtQtpI
CWRdBrfwn97stSQ4S9BFpQ+KIjQPDsL1rl3xnrya2rSvSkLyvWBJHmXCqHoAzcr4
V3zKKKWjlz5lsb9sIfe96esrhFpfVOtxhBm955G7OsKoMe2/KlqLTNXoTT1Dl/Uw
FPklXDxthURgKn42X8h35Uf5EgwVXHcl/SB78f8b2VqaFNN+cuG4PoKnu5TOEJyv
2fcmKF3fCYdtnNLkb9cjtyT7tQbb40Y3/asbqam94XsF9U2yy8xMdBnOXg6egEW8
1EEr1+8ONhbrIQURsZ5ph+Ez04Xwj6QZ5ItapnLzE4q41Hv08Xk2wENXZvmkznX+
LCz85BHNJLLXnqlKbyOmZ39NsQbjob6cJW2FWKeu3q/0QsG4Ke02MPdVCEReBXe6
GDztwkHN40QyeYiwa13CLZrzNjfBkyerTbpLaMxtxOjCjdl+cCNnl3Px8E/h8FI9
mFsuvhUYHQLZvNUvnQ9NPdf0ZweQqQJqb+x4mNdI+fXcGJrXwt58KMUivTX8LKo5
Hy/3vOsYAsndIl7CF3so8/gr7DdmN0PYWeinNliGiAopnQtFXCvBJlXa32D2wtrF
QpGl77V01jwqJkjX+jPxUOwZwPklUT1UHdwP7z+gq5rOW7W7pXqOi6wNAnVgDrSZ
JnDcl+G3ao4p1u+PoWuhgkI6OOEbpMpQ6nawFUH0Mbq5/c225kGQ6vU2kFNPieur
WfcdVggM2V9D6jEGiOELmX6oVuuP3cFqKldzburaG/vkd+fu7fzlfRSZii1kRf0O
nvmbF6mF7XEjkWQQjPJF/gIhQsgY6Ffmy9HLX/5lpE4yC1Uw+ak4jwnsUdwsmiuK
zKWUMzS7AqwMZKrLhLqUYi1jj+wDo4dGjd0TUZm+SFHXorEhTLFJW9oJnMMltR1J
N9j7POrMZC9qDTjSN9cF8a9gE0t8lbHC0dzrZY8dJXR90ATmfbg8I9feV4kt+0f8
re7k50Il+2pMYxDjH1wifq8y/NB586jg4mZSFiqS/0N/T82ZVLXnAh1bTtbvno+c
V6iZU4oOdgVsWCWMusTGKu5sCQLaCGDNJcHeJ8cnxSsupXf8BWXcuV19uresiV1g
taOt1fUDjjX1L/nSzcfoVDP43cq4gOscjLYRf8vCp0ci5j6Bdn9DfgsUBP3c9tki
IoOc8mW+U+YmqEmsDvezRI/FDxmWHVNZYMvNBzDf4n+6CE85Dtanp8esSCcwJK7x
u8Hio2IeRBMGeTdfzwmGubP/e9zB8it+lY1Jz+SZL7guc1G7o0Huo0VHCqonS0Fr
2ePN3ci4jr/T/NuOuFzNum8BQyxQlkP1TYnzFnqJzp4UnnhLXtp9KGqMKk4zlXcP
rO3wMajlgbOFe9+FFoELf/SKLLPjjraBRrzMaT1GofX7ye+Fb9m7eTLBtLboeyhJ
WCGpVQFneHEDHa23c8v09Spxzg2LMzdyzzq5qTvyXVrQIcj7nQOS+qU0UFUAhUJw
4dwaSHw1ivbIsCXO7S2CsI1UDL87JLij2riuFm1Q5nlJ2rxBuOTkC7QOhRnGWo+V
ka8WxP2lRNX8Fj4Gjwf5P+DW2s7+jE0CcJ4xxzsvnRR1Y3VQLR4Uuzj6bQ9jta73
QR0EENGGTcWp8VLfsolJOaWvyJO2watk7U6jH2R9SMMUyjltgc08PYPUunubMi1t
RZdsTMVePqB6kWZM48QWHVVSUMMxNQm0SuRLxj3hAcP7E82b62ibh8cfoxK7hECZ
FmA6mUnMB+Aul62yOflx/fHvU8Ij6T8m8mWsXu/q5Mmw2iw9DAPIZuUPOHv5ZAcm
c51TIlBPWZffm3kYHCeoEX2bWRNj6lK/MGdJHq/R1rOZlCN8hJBqFbujxF2MPl7o
CKOFtiT9VWetbn87w7XLDPw3l4thTZMQI6N4L/jR2J1IP8m8kUA5fM+fGdnz82xh
TyAliEhFU1T6Fz5JCLOZURZiPQLdHwLbSwADcLmlOXnB8TMmQiEQqpwvuo4UIouT
t3OM5jlVUNxGDgy13ik6GRcSPgtlIUdFr/SupqnHootPGCJtbVkWUWAuGJ91A15K
BHNNR46VGroyokJedVyAdtIcOxvLy431dhFIhJqeNGW3As4swFMKpiKEe6I3p/WM
KN/4jl1dq1wMSMZYlJE88r8W++Dh0ryEQ/2sAlDhISWz3ExiaxUqLzIN84f2+Aty
p5FCfhdOM9zB4m/HQaPkAko6Rt6Mllb+7K/+V8sT3sL6E9alc7v4Ok0Lb3sE1k2t
JmPiBP71OOPJ1fzijDICa4eHkrMQVjvL0VGMW5/mZk+B1844gFHdymouhLzCUe65
4kfUTHrhAa4ODNGYFYx9Gd/sf3ICS7SsVhdGeJmI0HCEdDweUifRCh8bX/e6qpEW
Opg3XDV1ZIWoIgJWppUbGJMWP/UD6K+1BU7Rpq5u98X6AUszFTIFj6A2BCV+b1bJ
R+R1C8/PsEIDenwfHVr+KHOaDIh7pLgq2uuPOXp2zQsddVIG1u7+ZAU/4H/wA1GX
J2CKTjs6x1EDyCaknGytXo51Bq4Evk8SUDxqgRIsCTjxo6T14wlo9OzYay5G40MX
anI+cR/2KykP6hBkQ41gO42Cd9NAafwf4wNrSCls6Vw+VZX9Mx8Yk/TfpHRQ0EB7
vKoJ0/CEU8zo2A/WT4bax6RDmdkdwaNGqEbJxtuheS7wNO1fNoMpIBnlWpc29TQW
YORhz4zRbcYghbu2O5m5pnW4OOpVuB6F4JzjGHubF/7A7uOK3zNuXbNZVo0i8MuP
lHmP0kX6VnQWcjoqw+Oj2dGrfOQUajphFZcBwfPgMxNZ/CQWz0PyeHnXMYxvHRQu
AJZfeMn847JPB0skBOWxexwnKpzplAq23hpaCx+v2Rh3BT6sROVDKhUgjfcYCxnr
T8QxMe+Adau94fL+XT+h7lLu6hwMe19tW5ZO68o74Thee8yHghZmim3kBnaEdRhF
DibZqA1pLJ4ZJNDZ2OiaJHL5ihUWc0bX5rPcrFR8/bdTngCjCXM3UAkMlqnqc81P
ZuMlhU9LZTpAvX8f4uKyAOJeThrWOwwPCxA620BFEpaPj7U3NqiMCCAWd2kBvxj/
v10G+4sKOLkm1wkRezVzhkURlcTQvOrToW3NYpasrsC/3EOt3pYo7kBCPwFvrQiP
JzmTDDtzS7aJIsvGmwsUQfLNStHW0y3TrhOVk/VAK862AOVS+fJDyEHvIuYFqLkb
luSG5h4S5KU3gKdsJmFd004lY540QZMlWe7GSDatbjEh++szUDrsGxcen7rI9xaZ
CYF08GRRTghsayVOkXVGVwfShftjqz8CcrUAOYSzpfhJhfvnPjYCTQDdq/N/md1F
3e6cCKkqC23yP2eUgVQQu9VmyWdf9n+95kIglsCChOegNNi2UugqowrmQVioPEg4
7fYznpVghskxSXaaTOVbz0eL0qkfGKy2qs6/XO6igcn/HXCmfm4fdZ+k4l7PaTsc
XhqiA6lcH1KbqTv2vGruSjlVxA6lI35in2FD7lkhEk2yU1bNyZa7jXVWaysjxiQf
KM91747dr/X7+4AbYCxQALTie/Wrbl2q7A/v7a5PZJ+G2Icd4csstwlyzfnNIghx
cJ7qKfWD0flPW13iYxkBItFBTO1JtOzQKlGFSx192Cz7UjZQ0eQ4wrf8/BxnTmH7
eLw05gH3AIVPtfmjnPuvHU8NlRe1+PmuqxZxZLRWmRrtM+3I6Brp7nD6UHx0gfAq
JO8BNhva78BgXPMtOUXWZpnWVYAA90Z5K4hzsfwOLQJSclPXg6ISY1UmYkz42hlO
kBZG4aGf7IqzZVKa8qlCA6DZi9YXgaVs/Xm0WSwpsTGU90Y8TKFlf3DBZTbSL9KU
r5vSjQcgNYFyAgqYfncXTj4feSNSaJKXBbtnjEYa5AgvJJZ6+imw1iwiHrYV/ZFf
6plED/P0aBizjINOTihScwmhXVrvtkSmmPlY8mzVx2jvf8kTj3t3TCjsXoLnid2I
ZV7uza0L2zSsVy6VDFN9YWl2eMYN4nwMX8OfhiH/cpG5THwk9Cgusq0gCa4M8471
pdhGU10FU8DBNNlmYWvQExCskV7EfhdScLcMXv4xteKdtZC22S9H8xbIu3UgxXmp
dHbEWCytxic38hco0ePHEXVZ8BCZqCQTbr18WNdRDfVH+ubZ/NymLnq6LKTjRBmk
IdWkWVqzjh++SBHUV8msc8kkiXF/WOHMdZtHOf1uT/gbNW7z2tgY1FWhCrLeQeQI
KG+SDOXWsSiooKOzW+rPUk589LQKb7Xcy35y1MHDZYUukAHizE5aWkvbYfPmA+a8
/8COGcqV4lZgWFfhDA1S52Tbui/ZB6G2SM2r0erq3ZuY+SEI09bIdDKiGnKl7QE2
WkOb9oUyJoNEqFdZ5e9VWXsLdN0ilJ1FYK+WTSlWejKLwRn2QyU7tzxmINm6JzT6
poPGW8hnN1cagIoHYBvvHy+aAoSFqwpifArtnGElUmRNQ4gUW/j4MA6k1gJ2aeW6
gNqkOTcPkV74xr656ei7vFzcTemvYNTTpj7REd6iKpwpMOPf2HWjGQKfNEaYaBO0
DXeVekFxJX5i8+qrhCsCjX/wYU6epvYpJNfOq47QCv1536takDjDyPSpnMIEt4u0
8kMXQkRqSo3+4lMWCOQxLoXvcm0iiMGXG0KDHHklynDnTGR774eY4f/F0JOFyRQK
133oxj/Y8JMVZ7DfZdKtp/VNBJ/mEUv9A6/6d+VnruWT68XVhn9oSyjQlHcDlSie
bbwwHvpGivhu3tiMyICzLLffQK65vtLaiUjLGb44t4EofNSg0fYknok/EQ+3wn/0
w+Br19evcnPYTrx6t9deAdWEKuLiMhjqKjbIJyPAu8v3Z0zw8hpTlh2WFBsC902L
QjwXEHVoF9ObqZUVbGUapT+1WjWc9BtGuPIRAlw+I8kPi+/Ng7a/C4SkSxZsgLXf
WjtwYomC37W6JZ8VxuWC3ZYPbZgqBbMsJcdElZ9TNHs+wOicfhkiLa0z7WT/TN4s
+ekI2/DsvVSW7lE0IfmjhkV/EesN6Kmob04qpGji1TQJYPtVQM6bGYLrtJIcIdie
GsT4t1mxh8AiQD1o2o7HW1ie21ngDwUYEYm9VzCQkmvSV+sBDp2Qq/jmsKEhigH6
Ywg3ofBVLV4XSX/foWR/XW8z1yYeLRimBigMck1Io7Lh7O8AJ0JSnlyLohRKlDzu
X9qbj+ZB4sT2bFMZRtUHvEbL84/eL0BsDAZirZxX4/V2cSqiKQ2DMa8RClTWgPCG
StA0TMXfRCLNir+IIoFrtpB/utwm81yfQQyFBMx3aMAMjd85mHmsLC3/ON/JWW7L
JX/IbBEjvaTzskGW0kHcA0kuHV2Bcr05JwO54tAzpal1HdYgkre5wGHZcTEkeEb7
GSoUzkDc3mJ4ddlAw7t9P2Y287IbmFSpK2/NmyI02u1zFR9RVKzg2GuNlop7caJ3
6N136F6Lkleokjxv4aTXR/4hTT610QqVjswq2//MwLAUlucczL9dFPbqV6PFk31Y
lfZkSa1+EwmzRCDjCRDbaIObdKMn+14/tzHm7Q5ezdPZj1EVyF9NQ1Tx7+y9du6D
L1G8ECl3ouihV9T2QJwmqB3bdBM6B/bTYVA4/APjmRMpD9lHEgKw7JzorlZf2Fv+
AOTEMmHCWlzfafizKDsLqYXs3+Yy1E/KRQA5qSSTLzeihNBX0YyNUEz1lkcAYtEu
ShVW+AdIwo7m0tudFW+SvrrAG5ZohvUjLbWbt0bkABngPfbrOpaT6EFXblzx4dQy
4eEMPcFwwju5697u07rbTHKF8IGwLsxG8TMl+o0H67jqrgEicxf6uDIvM/68GbTi
DT0gEB/zHO57xczY5ZI/lfqrnS6KLyNtceID1fIATrRK7Xq5m0PCS33R5Rg6IpVz
F3am+4nkLfAwYHDuX0LB9FFsDqre0t9fiZJUXCQNODOCk7rzSm6B/p36xtTl6trC
EULOGcfHl/RiHvsmfzGno8SQCq24plBNNIMwtA5M2RyqfIAP/AgnsYDRrvugJ1B0
mt3iLHSJ+ZoPV6Vtrd2gCzYmrk+Ii0CoS/l8nmB2PdcVl3FOEsdBWAnT+htNMsfW
/UciXtGpdEoAjne0MBKGRFJH+iXKnyw2aqa092RiOTXyASOHFuxyci2BUp19Ypwn
ZJc5OjksuIexntEPsalXqclCKgjEDfSJ3rEJ8kUbbIHA9wiLbBSIQXrvrJhlFpPc
YGrsKzlLn5gvUpwTSLWgZJkN5T3SfdHJEpzdUgnVuaSNhUD1uhdRro2S3HcJxldJ
U4MBGETeEJuTzYwTQ0SM7A8P4/NcPH8tgMk36BSPLST1Bh7HElU0VtHnnBSHhu/R
oCZtnrjzfS7rZohRwopokmflRi62eSjU2o0IYLo/DGlA/w0rSg2raPABEspgG2fG
RXQBY/Sl1ZrN5aWqW1sAdgDaO+Wc4qiucgy9P31O6gXSUN5f/UwwN8UQLuBDmC7C
zWKH2qE+lwssLTyzsYVkPP6OEpJjH+knLeW1nqdn5Wxo995rGBBKDGZPj1rH0tKW
LUqfzRdbOUJpokW9sM0uN8GAEEMee5r7Q/sye4Y859ZAz2PEL/0xiWQi92liyooK
/OdHFxEw/VjKkxaxZYyf+IoUIk6RuE8C24SZQcadG04gsKWjAn5MLUHVFxZAXjvh
1GuPPFul7zLjf7U1de6P5fHtsDjtbbsQ9m0lWPErg+0Y1QpC1Vwta/B5ZTKX4Vnb
UZH690zwo5CMa4giRKOhjVuVWtqXkrbZx+3Q0X/qo+GqguNIrVfTJar5vAVoFTMj
w/2JhQQ+0B5EMMZUFawOcLwUXpF8jmXae4wlp4PzLjRnWvRAYqIADBYGkL6QTKta
8TLMWHAbtpqJqK/JjFYV4GbOugjLltk4rOK9/gtWOSCxW5GTqrPOolIIBPqASYKZ
mRsRdhoh5SUcGXBhDWzjanF4oKQl1AXCcKEEWvy7S+s3q8MlJW8WMzQkS6yWSABn
zY0btrn6FtzFheYwF3KsjoKcpG19XJ0BddN/oeHuMzhjGuFxf0rGgXZ6PPja7aMq
cWvjfx/cAi9HDcJajRr70os9USwhRAg3Jb3RbuXTTfwOGmIi3q388ndy1gVFVmmh
ZFGlClsLlkloEmGvt2rQvAN1j9lzovnf299+AW8cBwLqTKrrseg63s42GMKzqJEj
PxWJcGo63zaRXwt53bFCyWN8raSkwQdsX3QsU+bzF+3/yL9fX20WLA91gjdk2/xz
SF8rG+SFDURBD2Eh+HGRws+wvJtwouLRwyE3wqlnKtA4jRDKaDrROvEB8+JrIoMK
t5gx03cEK2Prwis0/ktu9+8J1ZtUpDLXraIf29NagBSA01mz4hdTKatblteX2JYx
0d545h5qCqJGLpBhz753HC1iHSdBVjRSAR1HGfaJcKMPzaozfHSpSuA/pBENXlJV
HR7hDr/eKn3tFtofH5specgdNn2XK8xSY/TJyXtcY8ZuH0RXFasCHtq4tG53ioJk
uNV+pL4Kgmq/rWrac1hQD5Mg4115KBg9YNzJBWv8EA5ZW7E8ouzC5KLLKp/RQrwS
3HIGI32IR5HxEM/dhSpDFo8249PgBtJhQdtzxIj8LCYMzcr+bOAIiVxe5hB+tT20
OdFOBAlH/rYKxchBvCFto5tEp4/itAzQCXpy5RoJHGfkzB+3YTW7zmKEdhyYu1C0
4fHDQhPZglN7ocpBBWLFbu5hV1x/7D7EO9IcY4FKSlP9i+aIpO7MuvimaDtwQ+2G
MkbbUi82eQkrfdpcDo8S87C2hQJedxxGjLBJRLbN4xe530CpGo453XJn6Wg0Gi9V
mbWYnc4MqGZzDkFdNviR8HdUOc+IRfo0e8McMvjuEMaVeiCwNnF5RyzGE3SuLTD/
15ZfeOhsHXFVq7Nh/vJgso3wj9ffX9EzvGX+cgVcBdzMLwZ5X6jVXqyOEJUp78v9
KeHQg08XKzjjAnelLmOwYziYJN3jmWaQ/UKMDEvwf6UBP3LyPbxDuqxqLmjrKBEz
9kVxZs/bWFxP9v8cTvp8yLhobDLi4hCZhsVgrrZMTVBBh3cz+jmHt+KaJHbjfC3U
HL43eRxN3k3cW8u95HWYEqrb2rm8I0t6w6tqoKVwqiBNvLVCkhcgJ8FMcgDlig7K
qyHzmjm1MEFguFG6Yt1dn3UDq17xWwjb6zYEcAfOEovqzSd9G5DqEcbg0Laell8q
HH+GGB1jaLYcHxHT+fQz/0IkOoYI0eNmum9wMFGs+YTkuqtJSnhjbewevlfKpT3D
pTKfXM5fJGU4AZ55bgi87a4mHLWLI/LVtJXaFKJ4FpxxZvxuErtBpEOaz6yfyRtT
qB6EVklXvLwLyFIXTinCrvtSUWGBj08CwoQmxMj8kn6oCpRm0SmLd2mO07TCM6y2
fI2z7lnqqvPlgmHDPyaoSNH5mVzCx50o/daDmveIrhY7SvH7yasdaXkUPlmusp6d
eYSQNn/eJS+67l5qdDNg8PlS4RDw9s+l67e4iboVSzoW5HfSxk8Pk/xOnG9j2JcC
JXc3nevAQwV672j+3WuZ/ryV0OSZx/jfXt2KXg9p37zRgLtYZjPKieL+IjGTC7xD
FEEarg6QUTUjEX1GMNwPi0pnnOgw4zcMCBIH5tRVTOjE+Q6yORstC4Uv19UY8MiY
gtc89vCr0NAUs4tspEV0SVpkwbt9u2RwIMuJy++xgKKntZWL3lfvQgmtGfrxDkft
aSDlxpbNhX/EuL3CBs7XanZLDYDJL9AzJluYyxthFYnA/bsH7dMhtVffNwhWGOgF
K4ITKJC5H+zs3KbqQzmASQVZbCEPfupsKvl5qvNZS/Aqfjx0HBZDorqt4QlubJDR
h4fgppPZBfjTyLVT8vKzqlxTE5fmwZAdeaxZ/WoyMmc6UVmZ/73VU/IDl/8KRkWk
Tme+xlD2tYOOYzCgQnQz3LwYy77+69Q7JrLUby4e99ZynjGzeCRoJ1IlrLXhnoyL
7ALvWAUMsa7cwEFodI5EOn+qHf9trGVX+tnxPoA+fyWthy+2uOACBLbXFsfi9/Nv
NfJwvJ/uhAYBcVCBc+EUDCVx27rLYar9q6UrXBtBxkh6XYPSjTCCPGA4XQ6lrppj
pCtY/vkF3dtIgF3A6ffb7E39ONJLR8T9XQfZt3oz1djZ6WlVA2OeQi+YKBIRpoXC
J0KBpAdpC1zjaIyBWsXIMXRDFpDOuBG3uTwx+OgdM05SwbZ5zd2+GYhiyuERDhjD
sTDv10jyp88vmFth1vPSsk0/M5MSzSfbL7vPRtYweoQsTkeLm6o2WthXtjmzidrD
HPNXWDYqehMtYQYFvevfbZJGKvoHQSawOjodN0mXqPJRFhcwhzEhOCCLTm1Qg9Qv
LP3Ul8Bbu3pJM7vr8fNjFxq8RllAUxbgSNTy1B64e1riAleGtb17fOkCcQxVQJH9
d2+mzFco5YaXItMD8f/UOydduD1Qv8EMgeDv1slHnsZPdMN2Na//7fJQZZt2U77R
RQJrODGLsMLf4Qx1xpweXmVw+ah/3HUkae/dPdN4Yuw978/cgS28dW/Nhlkg4IJU
c96GtYG4oFE+NlY3nEfGyur0BCZFOIZezODeh3TS6MSshtOzXlv5q9Y2tS7929bt
xKKGUCQzEgYCM74BflQatIG0uP+JJ5UGz0k8lx7RRnyKmZi8zkwlJ8MMMC1B98ow
PBPR60Q5R8Hfq+P9pzjjSDLwHWHPuJ5JLGTDHbb10+bMfxvTot5k/qob0ADKXUg6
9PJxOlmjVkAhIogqX3vFKpC+1CLMhvfQsLV11IMoRdQs9tWEdYWd+19E0taayN6L
D0UwV1CQZoKuahxrrJqLXukdguXd/aXMeWL+ZFe9eB52WIdSxMtPGYmpmaE6Nl0b
QiMBbUVnb8mNzojy3jgKgF8VfdRA4z5J3yCty+bOBC0ZdkeeQhK+ReVRkjbOEGZO
/HwGYrWAFKUAu82ttQQtuGAZ7Q+N0mnJwjxByqr6ohlZixLbQrfshzMmsBPNVEwi
F1NTn5orhb8Lox9iYPPW2fYFJ3llZzhO+sM+CBgrlBNQJKE28JgHKK/3vNxUgEgz
nRV2miTCpmoO6a4b+I+fOepthoOylqjcI9TFEKG1XheethPiyM30fXKaTjy2Y4Mg
t+7HfKidZAsGZ04ZfpZJ/F2jMmZ7w9FHTrmhAoX+mVjrqfswUWorOw/Rvd/tPVL7
YkKsidaPJTA0eLTIlfWj2oIfiI/iJNQ5jqzJ000/3OKBtzQjZ5LevrkGGbFIQozA
iuPkkCymd+s9o67eHC78wCGZ1dbge+R2UW6iSMFB/WpjFCdwb2NSoQFi7Xd3YtmT
gH3RO/+p1SF9SYaKFZNJUMBr+90C8FEUEAlLxBUETlXdOTIXCmhkONy6DTQRO0td
q5RWtu3GKX3aKRZT+BwaQ5gelv+Hl5fY4zkBYHgJwtspxLVOTmTAS5HWYwalsbqF
qvB+dXnBULqSjZR8KGYiG0I4zKM5vYK+ABNMhTmmgyx5PuY0YLgT7a8RbIdOmoAL
SR46+v0wH9J3oB02IwuP4RMpvuj7MHLs2kuw8vfaDdxR4ipuc0iOxLp1Yyqv/g8X
0kWd2j6+ZPqDJ5qTztKbLRROXaxaMXD7/cuEZRSHVVe4UvAG/NTV2hNpGrsbPj6p
hkT98IXyAPdC0DGKgco9DYeGoaG4pQ7GW82OOV+J2ONDvy0CqSaJA6XkfOJH3hPa
hETp3ylFvvHG1sP32PC7NtM3JA1EnJajbOkF4j5L9To7U2dXd9JS0eydOlKFtF9A
1KsEjGP6etUmLd79SysDRIwCsy5huuTgAmNILPR8vEen11qZoS47fXqgOnAj5e5t
n3PntYmTgon+ZdYf3SjH2pfpwlJkTxg6fv/HWCjZ/tHV9dhCIWY2dvILuuiyZpsz
okQJGP27ZYVLAxHxJ9j0BSdHMfjF05ZuIDsoks3nwYMFbrTUbFvUkJpJ5mgy8qCD
Z0wInsuJzStMcIqmzrxdTY3RDqH+E7f5gOZ3PzUB/2gtmFV3+Ap5/9kMgP2pFeJ9
tlx/fcuNCt3NutTCUfFcEsyAHdnh30nss5wVds58+t/7HpGosuIcAGoDpLGNqBDX
8wJ64Bux16+iOTEY0MoBSdnNKwyWRg4SL3Bx16rOm9f6F/jCwm67eqjyRKz6PWWq
f3aCo/dgjRIW7JIslNNtAl6gZaGhFbGULMyfOlFc+sBXhaDIlq0MBlNgRs4aMi6W
MxUV3m2SKPz4ZsDygCr7JUOZHF4oE0SH3hkWO4NPsaYir92pd34wQQJNNsKSVzsn
sArIfkmXvjq1yR8H5YII2Khm+7ptjqJ8PS9fCPyOUt2NX81ZVPtl7sm2WSw1i9rj
ydZ30w/Vf0WZMziSuDMuEuvDSoOOcopHygc2UcLrEtt7IsRxQruufLjCVPesZy8p
h5qJLbpgcTIBrBJb0NIfoL4YYpXHAsZ7H+cQMQ3F/Ka1NllpwaLieuveuAq1cdxM
+ybF7UlcP//Xn9czzj1VpLgxQQmkFzMioZzohOH+zmR02DR7nvPbipQKruh+SMy5
YAwdrIqNqItlBTqmowMOpxRQ0XLPoBQExMCIwn2yRiDKRlOYL3pyt7EAkMfWGOPt
K18FPhoUTOhIchZZFQDE3eKhYqnf2epCMuOTjfOr1tOnh3BPsJZqv9dzes5n9UJ1
I6oHphfxniKEWe3yrmltBq8shGpp4f1KYMDsDpThW8jXc6LUcWLHYmelyPhI+iFj
JwH9Tj9UsIhB52+9pEtb88UvbN0iuHJAsaiIaAA3hUjtMsW+lta6DOzY4N4S9pcX
qpjdvotqw6R+tAPSNzUuqMrFgQ0wws+HkBX4DcnW3FvKiKyUhk8lCMRnOQIN8GSG
BEOUCoBP6AkqrOX+eA8nhUMc0YFw0TeI6nHOhSGEmojYK02tDWB2BTkRfxxUj3cg
Wdf0Fnm5y7RoZWzHqhcLr0SU47ciWQ9j3evcylvIx//0+fFL5brCGKvRU8/lqyA+
1VaL9bJflNj5rxTQBDD7P2wO+eQmm82FyeLUCXDIxGbhWxNgB2xAXbOI2Qcf+zKD
V6taQxxfyKWZM+Mat7nqLoTUWkGizpXiwU1WZnqeoNqqg4Oayh0mIThN4KavRU3n
GiIYILWuXYmcNoXI3DXmPf5VxPNptEzaDKRE8XVdovfh8LWHpoIk4phKjzKR2N4n
q/HDPvWd/Pkgu16mazNpKoFGeHzmw7ScImQCwjUd4QULJFPoeJP5g7EUDuEopXNA
B51cZxqqQvTMZj275RUx38DHLM6UanXIhdpUKCuByySy8vMhAhM8F7IQYc98Y1a9
pmBEQ1SELH8i1Vx6N0xjSwtvyatLjWPO/J55E5mVJri3fsLLIFe8SGiQJssIb99K
9WHeRH+3Yx0un3n0joahlWJ9UnQa5MEOTTojsz7v6h2dZ571xcsUuAxFLR3IEqyr
1LOjr/w8qujLQvX7JFEJdVz3yrWzbniGN/sdVHwoSLJ/hU3ygXci/Wo9Oku3eugq
1EM1KPxeC6O1t4xEER4LJ+QgCCEs2gisx4PZAolyUxdrYBZ7JXBDc7+l0Jt2Mzej
PYfJZ59JypRI/PhXHpY8h7QuwRQLspCexn+COXjjbq8ySfZmk/XmF5CLjXDCukzk
HbjxIq4vzYJxKrE6yeUwJ0YYQXLrOjAjljcoaqqhC7vNqDZNVbuFdjDz52x+TJzA
wDhMFKm4k5/YPQ36/d0nrkLtg1hDjnkvy3Be2liuPL8MYNZNdQLe+Nc8LO2xWeGr
3wl1r7CiZm2XADlbC4Yg+TBAgHnVWgrVsP+0HKz26xLCb5AQcHRKF6J+8Dl5Chia
xCG0lKLzgM7CL2wxdgabX/BQ6SXMDYy4WQ17UyaJso4jC2k2ihKhcXy/FZG1ySlf
3SLeXUr4sVWrYfSnxCX1XSVGk3QYfjlD/gvQopCRqxKALoDTfhK2f6thc1J9JGhX
qIRRRwtgboH13t/p3hkK0gTRFXs2Bu2cKZ9t/DgoLJdiJFr5biTWC2ASRTwHlzO+
GT7ga1kB2LcZWSFS4vEVmfnFRl8TQSkMsDxj5LzSPPDNyE9zALbENQqXh48M9Qqn
o7IeABfLVDL3Sue7A/p/rzhMbM8i7hR5dsIZQ1qdDLB2tvuyLwdA+hbZYXMDo3wN
kto4mgEs4mbPMSyY0tpCzgaMOji4XztFnbe1gxmAUZyfGJW+Hk3UZYiMvKoppUO4
82NuxrUgRFI2/GF2BDcFLpKT5x8XJza3KxIztSK+kRkSYrgBaK3PBx7J4DXWlqJm
WR4VxXF8QPr7g60JjwW4pv97m0LpHTbl6GWRdu6B9jYLa2+61pddue0eH4a0wzkh
srP1mjJGr1PxP7tF67K0XToJoJi6PpUjPUqe7in2xtjrPV9tk6hPo3N5LdSyy4Rg
Q/CYGmOQc0n707VTdNcAHK1tWUNY8LJuXoEz7X+RCNlrkxJgVNx6NBaUHnXcc07U
JHRC7wVqzGVhvaIdweyQ2LsJCLrZCsMEk+Xpn9Q8q4PPdxDcY0E7iBE6ShIjC6gu
wmhhdgA0VqWyEqQtxXnjSTyDC0NOdGUJlA5gtAnpdnOrHKwDYfKh+/m37o46Qm3B
VcPrqQXhRHllo4dVbpAHGIFPCE8fry5mWCxGbwL1L+qEpNwxH0Uvbg5WysDWKNYQ
0tQnKizK3SApX9S7RjLofgu6xl+2iGNFYGxeieXp8subirgktF1gDNaQ1LtdG9Ki
i1qCJv/ayH42cLyAeqQ1h7CG+ItII/7AlOkZyc7Mc+kBBXql31oh3bjPSxMRg6CV
l9aQNKvv7rjKe/ppKYDwM3scBLzJDrX1trUQTyjNQnO70YPsolNKRJEkGtwNp5pv
l4tCZqODai3504SL9rU66cQJ2cnojOQbUGJi7RTyj41FV4LwEL1tGZLHDQHhI9KI
YqCLyRqsSWTYsW0ij1O0ni1Fv8Bbn6LXnU6fa4P35InP6oboPrm2mRtG/S5p0Rk5
uXNzQWI7bEk7X6E0He4OvA2Mhy6NIobzL0o7wlJNUjJX6TBvivrbiMh4dxdcEI6b
2Vq+nGGOqpItuhC38AGG9YyefyhL1xlZdKnjwQ2MEpwXT8vZyJ+lW9M+ZXsDThLm
5ckZ5yX13Iuzp5SqRCjBLXo0DKiA0qVrUqmogLlBEJuss4pH8sl+cwpmjF7SLz71
+AQZvaOvutRg0+7S0omkP4L1cVSYFjFUnZB5Em0O57ySYFRwmINo2GXJULFUyCuo
ChTDXhuv9pbWXS0DYXQwWA4eGyHG0V05UB+A30g/zvqFgUVGW6II502lwV0gDfcB
JxYuzVnWBAnmoNfYnep8dv47pwzdKA2oQRBkgSVkMl013dHNf2fPSqjd/IRcmMCk
8ypavhBS/0Pk1ogbDNWOKaV19ici1tjvtFkY1gKzHYrNBG9XOsZ3UxZnJKxrVQXh
TT3xWwaZA0Hl5VoGs85b9zP44xh9yp7Ny4nAhON5lrqWaqTxPll4ozdyp5VEia0I
kb0cRDTB5k9XRX4A1yR47gxAusJIStsM65SAN6ClbTc6/wveKFi8P9FHo0203o9A
JlCGau/kp3aibvfA8aAGPGhcFlFgYKvZf+e6pKbMJfx88gpDvm84Tl0+Yemd28Bk
ok+MWOG0o9DtPqiN20ojmY20oXPkjK1XJ2wGO7fE3JRl2gWotZjaN++zkRoHNN2u
fIYpdX0oWCOElSCMd8+ZUCHglgpYyVrPbhDcvU7gnz5LPFUGOsQaCSzd/rtIhQxG
61WnUbrylRJRI/+AU2d+ftF8HKNPQvxFuXidftLPRu9GHfYTREuk7GeKjnGkECOa
hYbWV0gcZCv/6/OlxJaKO3rEC5KTmbY7b3TdqZbnYq+bDi+Y35t3AchKqdjR0H4K
GHYraInywRotw9J8NJjZQM8hKvKVt2Yf9iP1W7NefpUAbQ13rArc751RqsTV4AUU
WoDNEyJBuuftRsCGtCGpqfCXLG8OhK8k50mUijlgHqy1b9MplV12S/KCzJjEuWiy
BKdceD0QELx6vAgjr1ENVNG+8egLiVoSFQ5B3GLTc1q8l7MtLneC35aHC+9OrzZe
9mub3lCjaJrjnASsIktID0S0XznCtqXu41FKgowprjOJmJVVCpMkrPjIjQoZgkmq
aXpPVWpQizW67j/8MUoXn690hEWkQo421t1R0zZIUuxq+/H/gEJ1GiRPk8/1DhXx
iciI/aOJ7orJu27gVCie7woEUJ7KkY2wuX0cbK/ueKKukzx+VfZC4bdkb1rlKrst
3lmH2apjvAsJrsFQMk7NdL4Vj6Uhs8To973c3WVX7Cd4GGrxk7kPQws6kTWoZhvs
lCSaC67hibo0EmNxZGP/QFSkd9ZKeoCj7q0mzs0ZtakIdS1o/Xz+alFHOIm3AS5r
yY4BQ0uFEW0eH3ytseUllTMuTFzv7pBjLEKsGE3YIBjGHKvHO/qLxm5Rm6V4yPBZ
UvMUkmRpqe45WY6CU5lQzTqs7AcSgjTpVY5WFGm6Mv2j4MmbQxpV9iscQd+dswMx
2y2aahR60xrlp3IdvZPC8rEWfX1ofca83hbQhl/bm0PaJYaGuRMe2Xt2I4z+6aJ9
zwOeNxI3m3lShHkK5BJERhjkgJfGQycMPaCbpd2r4PBr1ISxDBhncu1CjU+/K3Hw
qClQGgnQWzFxwcX50I6DAWB/bxluXAqq20i0j7O5HxC2FSVaFQAF0wZWzYhftQqg
1TI4Vewyv+SV5w0+wMwvB7gcGa2Oo6vwtSygHpYmB6o3oUH/c1e46fGexqvlwAIC
k0NLIytK8/HVZmNLqNrL+UoEs1eWanHEqiGAH/Itfhr6lGKf3lYyWfpbd6MSGoiC
/yB+6FNz210kIHW7ylr5SJhv10bbM1hOoCx6Lngukh/7DDqfrxV51tY/fpgA4GqS
sOlR0B19w+NZFB+JFmlfMHugSmbkdKLUdOa3izdiJEzj723YnzQx2fmx+rqGCgwy
++L8BnRB6dpaQcYEdzFS2/eaGhSgSlZvlT9JZJz55nX/wP+8EXOfOhSJ6ErxmVkO
DW5ncFuST6SkwNPGJYpyHvladgCVRPPWWFMsXHTamCZ5RkUc81iIpQh1k3X/dcA2
agOGrCXYLKPt7ccW9q63rkBNalLnWJk6SxAfKiqCUIdv+VS+PdYreU6qMtBLAVN9
KwZwE5HiYwCik8hNycwBbofzVDRNz9vr+EsK5uNq2KJesb3yx3Z8BAP7eBONuD1C
ZW7NKXQi+Zu9f6vu0aCNOocOIBu5/Kg+vbud1/Wnupa8CCL/JxHycliKtcxkM5Ps
Obl7vnFMUGVsmB0fv4xY/RvHf3H20caWnT2vJmbzT2AjXjMOZPwi1JZxKWpAs8p+
GL+z/z+6Z7PHvx4Bd0Qu16ds8Gw3Qbkq5hz5zsIp1ShGZw0bMDurZIl8NzVAln98
IEM7WmvhZKNLXjKMTz8EImroDMWFgUfLNktZ9hSt4sJOWIGXIuEns7YQhsOVRREB
JgOMyx2ylikmU3IMjUh7dmT4EoxcSxbRED3Mvd3CH+o67/8WQKQMCKMHuXy4VTrQ
vlpoweVzETt9QveKyvGGOnPDkOavqmNiUNeAYsxj/1rBaTjLwmtqs3nla3ArgdJD
uOU1xK3nL3QGEwpdj7QfH2iLRGHsRMAdSRilKlOi1sISgzBhM3aetMLti7eHQTqR
5KNxA6M8tF96qMILbmNJ5AVcAVSJPqtRWlfpv/SXG0SRXn/LQXCQA89PPyB79B2T
YJuiVd/Ccrkj2kaTVtUu9H6G1CLReMKRlzskni94RSQLrWDTYy7zCdaHxtMiBwDh
++M5mdiX5mPNNln5DlikejS9FtSy3VP5jgRiY87f1q32s39hq3CBvL2vxs0UBlh7
yjlJ0KTNLrA244gnBwtlpxDOPhjJAh6wKoX89veyHj1iBOOe5MbccqxI2mB+GPdM
kP+ID6K50Hp519OXfm4XigxprY7NLqjulsl1P58geyWnJ0QgsvYxoRK7CkGeA6+6
jz8DTXUJh57awOO4mQvjxtZwykhVuFIe8LBjDaFmziyR6RySmSQQKc5u4dyVBGSH
+WypVQcP2JVWsJprf/kdLbmXSSWxvNba2CByZjIln3uxTdqwuP4pQXABYJN7ot/K
x89f5n0r11AA5Ew/70LsFpq9HDxxbGwai+9TKrOW5JtKBpU/F/MEBRwGpx2DpJj1
YlpDI2zq+xrE+w0bq+RifA4ERvyxGJxt7gKhu9TIecu6kv7GF6YkijGbrUpeVQQf
Th6QPnavII/MRmG0NvdUb0YBYa3LVPBktqhE0h6i+j+cmTgpHcVfxM+6/aLQ9EWw
CbqKhlf89b/7gKQl3yEpVbFJEo4p9m2NIjrlSQCb4bAaYkPWiGHcLTeo58Thb0sh
Om9+ffrD64fOYvEui3zJrs8byhj4Juz7BA2QgkFJB6KNA/aaOSYzoZlYw1Ki/j+n
d9sMrTLcby02qByIbutGnYTKq/SfEI3sZsO7A/P270MoXC/Ug4oTxaVQ3mchmZzc
4XzQtfx6mC0cj+W/3If86dyJs3MTqLhkD4xmho6I2Loh5lJMMJUQdyMsCmhzxW+i
HW0/qd/LmQUKFhU15AqUbzwL+TiHem4H5XA9RoNwRxG03NJZDvIoqmHS0b/+ly1Z
SbN6KX/AX81LuK7qbW5GgDrJ3LN2g11ZenvkJRuH0MQPDtef2e2maCU7rqNoxAqi
lVeZsv/QB1Q92eyUZcQKvlOKHcD3C2cCJ2XlSlac9Wrp3zMOBCji9qrhRnwPTaR5
fupD034aRL2c4kLXBR9WvjB7yEZDa8FQ8HZ+ptVcLXQxFU9DgZ1sXwwfgwNXTK7M
nk/zFW6bX++XWe6ZCC4SJKbro/rwyDd+3e5XOdUGtxm4N3pJCIvPV+0IQ6Dl6ZiC
Gi2NeCw2pTARySDEoJWKH6P9e7Dm2I6U8aZ7atfoBHbiprqP83+UGmVtGmc8kjiC
5xoYzVyGlipBH+j+tEXJfvh7C2H1FoacIWuEuznvWaQb8193b9UknAEGpwmagrTX
wOu53aoW4cVIHUDSOly4H1J5T6WYBEWaP1lLV+FbjPtxyAhdWYDI9dMuRrxOKd4A
12iG+mU8Mg9ROtNNwgMKlyQYx9P9BpJdN19wSSr/ASgJcict0cQ3DLxFMSyVvjoy
pYcKLGp2qEfwn+w67LKWBSPNCA1ZwoXO34GjUuHB+aok6CWrgpzOc6qNL0UGFbhE
5ULe5wGqMr2K10eBY0GajhOSD0b6XMKsqPpm5AOm1PGh7iYw/PmmmEYGnWXIed43
PBh5XETGdd9qNtLApO5nTQjcpZmjUVMBIgcdybX51LV1N5Oqbe8f2vbhuJHFQMkK
5I7U6pua+PF1jdT7ik/cpT0VY6LvxpfummP/8R6VRJNfmEh6KReqbQ9OR50IJBdi
wygEhPt0SuORuWml3c1KR/bOdAazKkhMwDAplO6NoRjl9tf/KilJn7+Mftzxocrs
WgrDoFk5cMbSR69MAI4gkthKmzFcvpVDgqSzE8/szdld5va3OtDUjnW4WIJl25k3
t5j7XP2fimtkfWlf2egCXiYUOvctQ1BNNmo56xfWx1dQmJ/J/wWxkE6YyfCrgh+5
jXxObbCRYaYlhGcagj1tL2gj6W3QdLH/AYy5AKjZTMT3/kcyD6ax+o+ucQiOQxfW
qcv86QtX2BCOoI3f3clzhrGzmAydI5BMWFRXXjKuCL3b1LdoII/uIBb6X1jRKpVJ
zGPWljgYro/+erR4zPFbaO2A9ggA5apqKlGOJg9e2ngm1PYAJniPIZXPLXF3MhSr
yjmLz2rKf8RVS2VmU4ZkWT66jSF0JMgzTwkFpPxWEvqXBuurJuviY+Ha//bISOi2
89eheKg5Zh5qtkf49jpoIgQw7GfPHSxrCQxeD8CgUwMMfPJUpP9GDbpEXLw5A3C1
cRmGLr1g0GOp3/otTdI0rNzpc/XdrKyt4mOgcMBAqAgvJpgZHjtOmdoWQ+RzSc0y
T6RG8rOzppZnMZnhClv6N5LaQyul0x+PUNhQDN1NrWYrMQch1ODzeBmEFKtNoPeH
pPdZJiUBCfDCvz/KkLKedHbJu5N6KjSAqeDGwhmrKm45s3b9v7c5uN8JAu5H7lg9
IM7aLF83BbgLKitggH/aCAWyxpNkjve8z6VzCgTAL1s5iLSzb6fgFhD8jI7Oxx24
TSrK7pm2bWaO50sTLUTsIUIebT2JC3laBtAD7VkBkM4BiMaZFiX50FFCBLpjDMoh
8l2QU74mgm9eaDvhPOIYiGc3hyVhHLr88uu+O/4b1TaVnIVgkbajdFEWPxmHmKmS
GLHj0Lw9nfPDUBJmvz/TBlUmP3an2B08iALWyrUF6zaVBDoBCAFicys/ytmTTgpz
0PP8BpqOHkmMde8AyDJk8ozEq8Zv4MmtpvUr4pzbZpa62MxU3W5nkG3jWm3hHpy5
5GxT3TYbOramAreVsK3vvTzTBGBrAYNUqFQt16LMmvRwJV2yX6F9aGL2LLtb7P8R
7BmqTb4auITch2chAGGrVTlaBwSejVw7euSgfc/VAlHNEL/d9zXCymm7/jSz3M9b
PBmO74Di5SC/TPMvf+3w16PlVW93Z6Fz85B+XjGplhupyplHiPBv8zQKmXx0eieW
xINbaBDQVY0Mi64faGqUk6T8A30kohZg9hpRzZZSxZCtF615+417nbIHaBhHlN+q
YcZwZNtQW99GOaunmg92hcnA93LlL7m7VVD87lehiiBx1HDre/M5E3bN96lfdLME
ETL1e158jticuqw2N5qcM975CGwk6x97cH04jlyjCc2HEbTckZtvRgS8G4lC9Q5g
rvVaS9gh+1HvWrskgJZHod72+VLRc3JwcraszUZopxleK5BqfFM9E/YIr8tEMfbX
OlxlEYNfCxy/yFl77tXxRDQ1T65AnYSzwjo/OBEXhfRBSPYHqM3RsEl0QN8g6eyM
+qlXq1ZjLiVtAym33Lk/fkn0uCwv+x+m1gQua7+qkrR0RlLJaY+kECozCb+GFyxi
bBdv2f4GSx0/pw1T1YrzNyjgxUcbulY2wEFBOTLyFSXoddJFQkPm1dswx3mFFLyB
TxJMN1UJa8AhWu6najeenElBuK87FmQYII7y+VXdvfemVryd5wcZnkNdvCo23YJ8
Pdml62ylaMx5ohdtIiM6HIq/cn64n971t2rB5Y+XgMzJpgQgQqIIx2Djk5MXyBDz
eoxOkIRuoh+14JruOWGS6C6WEckyCf7IOJRPaAlElBFD/yUVUZI4oOcONiDC5nYh
sZmcVGAOjhVRvSzRtKs1QzHDZqamZwrhSc5pY4asAZJbWWAiN85NvLicX2r//q+1
QJqaQzOvwayAgzeOpBacwXp7N5MV+ug1kg9moOMB4ovmCW/+r0bA99tccaOFYYno
HiK3WAh9RM4VTQH+8LceviPW2PMmRuAtB6++74E3pHjVVBmg03AsK/6WWtkRTaGF
xHyLmGKnubyZsPRfLhOkAFp8knw1AKlvfOaYNrgvukMus4VSHPxoUCUdl2F13kTm
dg7GExQRS4wM6Ix2RkE2U1mP8GKxJgM/ausGk1XPmIu9RphqWYHxI+JrJZQ1vfvk
ZQkgnTrTpVhkc6N569nFYQEh4hB1UwC8tRsnkNlVvajSA094qMlRWbSBazCun6bK
MOfgunTCIVRIRMCEvF0NQum9cnhBbUdZShcWneqgxNtY/Ov0a1axzngZfLNyukgi
+x6e41xrAi56kLIsOj3QQCPmvK9C7+Wn4qSGZWHnJU59q++IBOJBX+UJwiiQj9J4
Z9wTzgykvc6YyWW3pAjnJyINBB+xBdKpHDgZk251Uq/HZ4J6iAwXd8dilIC3ustr
ZtmxG+MbjF8Yvhij2DJPyJ9ckstddkZn0fhchtm+qSO6G7HC0AFuYwj0gI7v5TZz
EFoNrwHLq176X9cTnOSTTJV1ddErnncda+cOm2eIV5w1TUUI66LpVFP+XMDa3QlF
bRpaQFtYeUZMEh0Q5qE16inHhxaU2gynML8zhDZfFgIGeRerVduhZPDon0j0lAW1
f28jYhWsrd+ojxR+s1dAZB253B9DPKL00jnkPUTXc+/0zKi7DmoTKTg18Pkui1oE
2OnCa4hBSu4nN3mJqXpRo9fx7lMBGq1/PmRWZke2G9GymtGoHadfZ44ddDtbd74K
PBlDwAqVYu8t4EAen53GwtoEGe2icaOw+ItKOV+uqcIf4dhPMzDV+e9KaB+91qeo
D0LPFeRlQt/tKjQ1G2K2qzN7fSGEidX/vCfjh5EiHEEqc6x5xyCpfKWOwmtMa6lQ
maBwygbF4krW7/yM0ljMUTg6XywcDcOj3VPBUpufBdX13eB+scjXIz9MTOsZeCp1
6GbbUEvPLM4Yy4rlZNYCWf8jESFIaUDYmi6czrBV3kv61DNRVrOC2vGa6j5Bek0Q
EUSTQLFaiPAGojkl4mVT5yTNviUxelu3cWQXV1dlUY9cwc8aj0UFFn7bAYgujhU2
aE5OHRp3DF2S/diNLoc/80GeJbhzH+QXFh0aoZ6Wb4DCa1UdW05XPZcrIlb56ST/
B1vUTAUD3BgaoBP3SziQZtqqrg4j+QxC6nRwUkBnMnihSz+YtPR5l01LvueRGCgM
ovBheechVcLDl6N8fP4bnz+75WDj8Sn1brGwDGCO7ictlViuviDs98SNM6NbwITI
ij8+2X2oVF9QaaW0yyu/MIqN+zhBVrkNvMb6LOEnPngq/lghgdJMQwV5XFMTdOy6
jGSbgFSYtEZ/v8PCAssFNJNcBo51xHYHBxFMssU231+2zuk13IUpv1sUgP3xVFQI
iqR5PijYQ35V8fsih+ADqULsgCGwV8v1qQooU+iDV+c45HK1Su3qgt4J+RgLBDwT
MmoJKSgZX0UXMAu6yJOYXDSX0G+VcTQesoqSmsOeryW8B0x4EmnmSSGSVWZ8pCxq
m5J5GmWXBbPoRHizwiyOgNs5Q4GVfhLgt8XbJv87c/SakuELr48sx62gLA7h8QHa
88py3jIWK+75OqF1lytazna3PdtXXchAWoBByydQJv4YH1xGAS8nZM8dmlhksCn0
6lUiu0jEN591N8nGMZj2ADtHJZyymryJhEIP5fVZHkUxjcS/sAaYk/sFfKMSsz8W
GLGKf7haaI/TdUDN1bAjdKZI0uW/imKb5KnZ3pfFYMDjuqKWA1BoORvoRkiqhZ1K
WYhaZUx1+PBmC/S66bamL2RrE99Wd3TwCkp3U7htJwDwJc9JbD8GlZz4nSbHJWyj
wwJn5noXD4v7NGDn8H7N3ApuX9XMldz1sMbthCv1jp9NANToEMA6pR1eKB6O562Q
Cd/x2kvt6UKfV2rOnetoJ4ddxb89PomuufGX1sYAHgbQtJkXQHFWnA6asTACVU8u
qxm4UiNyCt7qYtOfWKc/rBH3XAtJLva9F3O/ppywjq0zY8aJDn8xw7sM1T8shEuz
qejQhI4YdfaBLadvDk4oYQXMC7PhY6OFlb42eR9yTGldlwOS6j8iTDDXpVML5i0a
BRFW9N1bo8jWucxBaHwhx+j1VOZCIS0lJ1zS36V5bC3amE7uI2rucGOgPi79lPpx
uarvZAsEm2ECIvPLumIkaqAtT+/cIrrCzASABpF6V0Xmhzzg0V2TbxE839ymCr0n
It/skv/TdvzsrR8p2gvb7l+NNPhcUSjERij8S5C2zkUalctNmNYWiNOydP3FWQEX
7Ux64Fi2LSPeUT+raVNbiOZRuPEn+IYC37SCnRLxO6DNQ+iInkUHgYSL62zsfw1+
bmudg/S38l7a/JrhRfAjZ7am/tkCWgxX5gIQLe5mIsnL+17tul4WHVJvi8+fMoKh
Mu1VEYAb1hwq4yx7C0XDdjN8Os1QKpSnNfB5aAyFoIAYWOTTAM2ZryHVj1KfELtf
HjlHENgxO+Ax9GQ2EEFlXGZBXBWn16J525y+HkhscdwhVKTKoRuHIqZBvk5WdYb5
utcKoeNvh5xbtKjY/GKcY0Y6oN+0lsmD07NwcyVfCfeUhDnigPDFVn8B9/ArYRuG
dcn5f+yi9PM6u+9KVRnqZb6Nel2Op1Ta0ml1Osc1voDQ53i7m6uJ8zQGj+E7MwZ2
zgbxmMzOUGpSu65XEYoB/2GZ8unqxOD7i2xV6OFoF0z1XBn1d4ljnSNbA/rH1Cjk
qMP7prGy6fdKnAz1YLcR8t79I3LgnPJPpNOR6xZAYuFc9ac7PYDCRu8zEK6Ppek3
Xs2uVk6vCe6zltVXOE+ewEWNhzUDdpgbq8rkC4eZiwwdP3SzGk79wbQK2bYRVdw2
qvp8fMyx+moJIH8hRG174WPZP0sRqDrd1CBqTESjw5WORTXuyGxPeML48kBldCq7
0AbReaxoJ9JNdwFjG0xp+Xp08FMvWVDa1509vBN8Khl1rDV3eT6TgKAaDn5ZmyDC
XEsvbYJiecHeNXV0RqahfMGdrR3wO3eDljlCtd6My+FTxBCmA8B8M1GKxPnVgbk1
uICSd1U4n4v1LlODBd5jKqTvdMSP/Gs8SR2brDeAAiTWt4FU4x1Azej6o70JcENp
WSwwtAWmBmkpIkflrSbb3Jp4+XeUXk51Uq1GN3NTWtFSjJJG4KHDRfRgBkSEPfJG
4o66qIzje+dXXZiM60vJWoMlADjuxpk6pnJhWylVha0UbPgFv4gNZDF/kKshIIrk
NoTgMFo8yOcERZ/UhTFcWYyQIVg1gfNFVxH/QJtVRy5259ZXvvKsXJdXv8CxNiHu
IyYgdoGejDxYlEDf9ykRTEaxFRpA/h2/hinHfbSLYjxIFEatRh3MF2aZdYwaXLFQ
1d/tOrpjv/O5DtiOOxwKxeSKUCJmVewb39/zN1yV57oOrnMkowyw7aOgYlgrpPxk
yRr6ELC0W6jeWnCskb/uqFiOQjU2EY0viTumi2y6X/UgPyV5p3LvNDTTL6P0alMZ
/dbZ9YPzX4st912ihb9m4nKsPcQUNESNvYWcvqbdtd4emR2dgrF0ocHpnsaaudSi
xemcDKN0GnS7Jn9FpxR4Be08T4kj4RRyYlradFUNfAzuoB0WEOpbDwYWKrh7uLv/
iy/eKw+lM810ITbyAbAU2vLou1xi0StKBIXnVj7bf0gZMJLTrFTHhjFRfdemh/qP
yz4yYKtsTY1BbihZe9U1XwElkZtc9UHw4D1PoN9RmFl5woyWo24+ivZcpLmn3PIe
PUVFzSKYwSzrERwt1fIhwr4XWpcXEiW4IG/Cdat+T1Jw23vqQ7LKlk3zqWkX3OwI
Wntil0X3OPeJSrKPc7BAydyRwoxIt4uGqzVira2WTB+d92Ic/WoQDWS9CG/e7tyZ
RBWMXSkI4tdKpsOaTFuiMGl+2cEt0fkzlKlqA4O7i2xywsw8Fw9awAmZU2DSs+B+
vEzdN8Ht1KJS2Ym8CRp3iI4reweCITcu4iCqXpcVtGWo5cQ6+0jN8vChQyW8rPby
x4rdf+ZanVJ5Jzs+Jtwso/nnZWjaO4DyhxYi1lVPqXyHJNRNtmDXi9HyppQfdGwn
2INKx/QBQ2EyZlALVmBR7mqd+o9ssCZBslrVtOE5aLcnOUO8bEYHr98vCCaKnaBK
NKFbENXX15IBDLiabdq3biWRkO3biAMmuLxSG9m0sGV141XaH5IWy+4yMreLsITF
nYWaiDuXk8mVklBQgv4ZK5bsBZSt1gwKAODs1Qp5sn0+61DVGvwOiFLg5ciQ3Yga
OoFu5kIPrHjerNngAtmpwIBRIQStgpv5DJUyQxG0vgsu1KK5T4T/TymsnDwJtZY9
MdQaPYSTVkLPJrNVYnPgt904PArNKLRH0M4GDmmKRIV4zBd35Ivpsy9Ufkt7lqHh
3YW/UCbKSG+qXLzmLsnXLi8injVSmE2gd4rsmy0BUhYtaVWXUmhJ1UJ8BVilwSYj
8mS0bP8fa3utOChiF+9O09zoBKafFO9CkQ6WIxe22citEPBCWv8p6mbI5Sq2EKiF
lu7SuM9o0TLqj6n/JpMdiheO3d1jp4yBzNgjYZHaTR30ZI3WoOR+53wFYfHt1Br0
bAccajbEHbJ8md7Bxnm3kciGyBY7Urvd94kkI3GczxpJm6qp12h5qt3iK1RSpeRK
Nhr1wuVxc1XkfPQMXbXdbPG2Wn1oEbfMBoqdPMz9CKbUXIKZsm53S2LuUEg1V0+P
9rHdvGAmtSVidP2rvHikqLbY9rE9rrlTsi+QPOzPsTQRZVxWE1w9ML/8qUAWyh58
qtkUnqlkhFDWIzLdsyFgd1KFTmeUdIdFpxt9ppJd9dSsmu1VwgaEW/a1sQ7gtpl8
JGxYAux9PiBA5wSVvVd8pdUFoS+NKgCydoGFY8u9rhzwkw1czzhZL9vcXVuur1/e
UVwZPikuKNKkNwtF7ati3J/1Bp3yqBvq+DUjHMAI/WR5rsyJbku9uJ16jqSqwrZQ
vrPSp2Uu/oyL2vQDmWMriZslXMSUOYoWzwPLcEGynBD/42HHUpJMOoC54ZAq0RYT
HjzAv8HL94pya3fY5m3cbMF5hAdjGm1Rf2G24sy3vJpS3HGPSib4CyTOBdxcoQEe
O/fvcsMJoXLfHGhxsioBQB35By8TRnf0Bgelx8lWndpoWgxoZDkVSmyFUB0T6qKH
RFh6BB1j2fgLLkBXOmFvfia73XsH4yGLa9EEzwuptjDiAJ/ZV1lcZ8QbahuZGUBl
2+il6oCBIrQkwjjuxmFPMAVIhi/N7QqJoiJMP3ZVl/VuadxZJe0PP7ZhL/jHJRFQ
Yarhrd+1Wsqzmp7o5PzSVXp7FuSjKSDxy+HlMmU5P+kRCqG7YGPh3YSSW1ssqFMo
5QHEU9wrVzg8eeWA68UwQxtsYlMi3E5z57n6lczGgFRBneljMlylEAKx1Yj4fQZS
cdT2EVHAIbkbQGQ/QO+lRcCxXDD7k1wP6MAGnOTsBTyzCja79UEjsW7+zCwUmom/
ZACGX5dkxmcSvlIfN71JrAk+R2lT0XnaVMfRCWK34hhe1pLd3FNhCUzW9kYGoFU9
NigxFEbiL4lQ4M5exYaeLHs55+HP9cFYC4HO7tUObbXd4NWYVrUE/ihP/g0ijpto
3kvQ91+sYMd/c0V6d5cUqRWjwmZqSpK6qI1gOqY58EnOtNwXmXnDFV/AZ1pBBg/J
FhuGJ3WEIOCcg/ApW7QqiYIEsKKP94sxVgYd1RxHELYoVh6JhrIgtnW2Gxd20svO
uze82dttPxnKKo4aj6Qcw/67Tfet0fxhh6sNhoUOkqnV3zbwvA6bdnNFV++GtiIP
Z6mXCNxiJkaduxUkJSUTQDbsqBEiK0yZH6P74hf4pyoaUnr8j2a3audd+Ruse7wZ
Jiafu2akvT84oonjGGpdbnC+lfyE3ZwdgJgUfgKLFzn1PBLnwcSRCfoyhXj6Ao5U
ae4rwdJxoIVRiNNIWVtflRYl/t3FoulDT7aEJ3Xf11ZqQlaRD3lZSqp7G0Bjj8AS
La0R+kVEz2JKgCsyRuiwYpiuGXhzCszgzdqOJSP2khBOFUg5xl2WoaR27JyuRE0T
tTYgVFhghIzPGQ5dwblE6t68jMiCYk964nsDCPMPy+FjsVrLMv97hEFu3MjPwf2a
PFJFFN3WVwrLMe1BmAH64rGyNziJuZeIfmAkMPQqOHnCEX3GxVuKkv4IoURjrm9f
NM9J2F86axz7CexCTSbNbviOoBoDVjXFQYGf6hK6Qqx11JimPxD50beimjWA+Fo9
q/uhuS3aVq5nvleKPOcR3m43hcJXa3oS6ullgDzeXuGXuyGRHdxs7KAjAryv4w1U
9U+Z6jVhX92x6lpr9UHC4JHItg0pp6C7p2xkPVPHzgRrr0rBIy8hx75fWZNezWpe
cJmPG9egwpvP+Js3a8jWxW6P6t9fmN0Ty7iPvJ9vT64t26aqwp29hTSBxG1KK/ZR
80b9onEXrlBF7yc8eRy0fwCMpUCsz7D5eyTNpNYx00fu4lK+H65NX45JbBoZb5/r
pA1q+Wwq8Xi7ArXG+wx3/8o8TOfo0LkyTBHECuvsAPGYORH6KhdHAVLM18B58mym
ZQxSnloK0VwEDnJN/Z7KrbgoV94Rxu/kC+B8e0ot/ytDeVW0VoLYJrXjMEt32WAC
oCctN7kAZijpUi7n/L03KRF3dQ3VR+tHT405AXHz8CyctC+Kpa8XegKpVdJWEObQ
bc8qbih6RpaNpNjZ7RqQZa1lny5DEgEvmcAnhISMb2bXgIFBUqpb0PLbjIx0Bvff
uusdEzA+99W6KiRZu3pSeg13gvT7Ef3q2/LsybBwfEM3Xac8STqxvihHTvp1WQ7k
3au1J/lQxhypHRy6x4ggYgkIYMrbjVWGhqaPsp/x6/fZqfdGEszH0cIRcXEX2yba
wp7Ekpeaz43x0VXZIJUYGou3zcbtuVI+/ooKavbs8eZpsSrLc7uXOWRauhwDs4z5
kNMLk+eGSkPVFFHcStlhu2jOU/mEBknCbfarYEg8L8gsxKk5bOXPrAtDepBYBgxJ
5zn3y5mdzGjrn7skcaW1ftiR6thOpaTgtdqSQRcfzXiYNhm9OY8SgMqR5GVM+Ouo
0C7lYfqCmwh+0dHR8xin1BblkO35e9ogFtfxg5IIuAYvwQSgwBW0GK17zuQZiaqb
bFBxFQLgYl5LYdZ2KB8DXhZh6yD47GtzMsx2LuUI7pKAIdkcNrvpXUKqk01xO4q6
NyuujK59sc7Mcu+y83nTaGeboVOIoZciZSHA4BXhaSMq5KWOZkl83uboBomir8Q0
WZXlnb5QtRgtkZ2YYXqF2kwkRnqzsT4N7yiN6blRUkZ3iLWGiLJ7TRz4hwvnXBlY
8iW55PPK3pSN0JpW3H0MPJr7AqFiIBUvImpQR5QwUqdmRNNdB8FdJNsmPtZaH4o5
7GhPy/mSOVuSgoWIpxRiZoKXy/OQhMGE5IX9RugL5wFZL47OYzVlQfB1J9OHCw1w
I2AYn00LWo0DTBGGLBujSemuF0gadjrO84g10iM1EndhLSWcYajb6JwzAP6XIpcQ
W9lX4mUhwyC94+SuitLof6/F0hbmM7gizG50FzZzrN68fbtWrPFr1puWo1b2W96X
8zKw14w8leEnxgUlU45Nzw3t7SBeAAjVLvkm0HAtH+4ccoqJxmmGvXGzBLKbxVCD
t+JrmD2l5XSRraIbPvdoAGAfa7TJ27QBvKMo7ZDw3GMBNpMoUnuHAwcwDR/rBAEt
CVsMInD+Tug1xkA1USFztYo2HQqqZXu4zyJK30cRgW3otu5WtOPaNrYbrzXNy3CT
PqKDZm15+cesrxYwq2IBDPyJjAHbx2SvVe6E4thFYgIJpsJTnLxsBAvj7luSMAqZ
EGSMd8/xaGtBglJU/PldBaGJHGW4Q7+xLELhLXTp7ggYKphqwLERm6Los6FnIpme
gsWcinhavsRtC8waJyaO4V/YMSiag4BVEXMqwyXgUIEHFdEnyr8w7XR0G9eF2Rry
RNWTCmilfxmWmzm2EZnvm7I/XKHVIT2k3k7Bih+rCHADC4Ef+9dy6vRjMiOaeQvd
gCc+k06BfS28xQTQLGIYzVIhak8iccU2BSaLmubNSNq1rj7yGUC7z6JtpjCnjRwV
BDdcjWgK557jpG5jW574zJMs6oUlsPIN+21StlhS60YWIgs0tT2+HAsTBP01v6zd
JIlr1lPdq96FRhDqEHeQzAjPwdcPW3POzxXeBl6mfzUGy5kwAQ7LLQqXvyG5m/Un
mi8hlTB65XVTaZJ6efQ3opfAtwhxKIA9uTnUXahVcdVcnPvASnCL68e9mREdYr75
tY1MY4Emfff6xwCoesFgWbDyvfAxXFwE14WJ0DkkXNkjhxVw21UgpvdBrfyqamxI
LYESipBFIqjPKHB/gKO7KRfnV2jbjdYft4YioxCZCIrIBzmgilzmJsoV77NSp5vR
bzNsoA/zC+Lm7Dqe7LYl9VpuBeRjaxs/kiFBvAAn9ydCSAChGdjPxxl3fs5Sm5VI
kG4EJ2Yrv3FT6kYGUvGl2xXkkB2buPOAJMZnoMPHLitNJ+aV0Dw8yNd/7jL+KiJr
SyLHqVnRbOYUBUbX5ExSU8pMqrk3DbytAE+g3d0cIOLUlntXkEgUUEyhB/c4h2Ie
UaZdj7U6OPql3/YxixOlLuu4zL/IQNKzZ4GUJhWliCVMnHgssANXNR+m2hEp2vTx
Ma1obOyY3PmHTYnYiq1e19BmRCmd9bjl7axJML1Z7nnAl+WlTZ11EDU95OaNEqwi
yfRVzfa4+LfjB61HkYtBRaWYAqZ/2dvUA7ArK1NnKp/rz3Kr1cYg8QL1HEnJGqk1
4mbusEeomIHG9IL4HQiTG0mdaEcWVR7gKypSbIrJmgcttUkDPKvPPk3m65E2QjJE
XRjO9FqtY2bb7US6UwnPpoI43xqf4UyMnov0jKoGXp/U2XdztQiB25hJv+n0ynRT
dWnSwPfAbUAnOzqihuwPFWd/qHkJNTdJPOqDI+XjtRIw1vZQ6t1+4u22NxhuEkgn
yF/tFOfF47ve3ibD7QmzKMdXGhyDDXrJEQG7rggt+nc8aJ6PeSRvxIyLq7oFBkux
dpAC9N4ePwStKItKLYZUWfpbMi49rpZ7E4IKUo232WNye0+fExFYnpGcOvNmveHL
aW8dvnckrkSN2nnByrGv0RZyVMHHAoQK1pysNY/joC3B/Y9miADDiqrlkV/kGBma
/S1tZWh6irsHVzRJg7vb0gRpgtBdGG+LX7emcTyB6a4UbnzYymwxaNMQlZyZzK5G
gfgBJQNQETLBIbyPhPewaAvCAEVGly9lYiYlnoo4pdKo7KKiUcjJtX+UfCwD4abW
A4tgbuKh2Xyl8zROMULNw6v4caor1CnQKbvvFzeFcVAoHqhhyFLLqPIislaUmWhv
wnJwCuTXFgLn2BKXJ1mzabqeYynRkYU4CYpyQ/kTmLau0cxTsUrvuy7khsCT5prr
l0Rxk+bZqsOTHbzJwrafeNLBjBV+ygeA/cxsvQYmr0qta9Jpvg7ZF1aypKe9vbwr
W8+o72xQrMofx1UHX+XxNVmHt7QitFCsZsEMs434s1O5QArvDr48rH6WrZC1641c
xQcYkxMf0eA+uHixqhASw/laxDXMd52ZIHE2qRlYQDCVoH6EHub3KQpAPWvy44Th
BwHQB15M9R94K3KFAsYcQ3g7iBI8IT7xhvxA7XA4BDR5ThvCuVURSYrhXym1j8ju
nLBPFKSZwjvzXHFH34gqi34jRpXT0PrzKoA7tlHq7zCwddz79+qXP2gMGoMKlqqT
tadilnt8kSgTr/Fpz8jizwtEelXc+aJtTOm2aD21445THY96O9Ozm6UYHmL2A3AL
3mjp03CBmfPqwAYS3qC2JvKBu0LWCsDTL84LpWRTfg2kD140K2gCGhl4mTN9CyMw
6rjWAjwOENQ98GpKeGQl96NNOSBDEGi3ppkJYn5HOVtfEVaeaklLpXDkWvLwM7zg
XBAsrieiZ6B/qAi+yXH0IApFUXFIQThW3H+ysRqwAg/wnP9q+SD8xoa6J9CEMIU4
G0GxbTd3dob2XzqHnrnemk2tjrPu60wV+4eItp5CtgC0PfCJptXy2o39Ee1xSUXz
vYKw+O2s0QH6qkMN+9co8YY7exNCv7MA8aY4l6vUnafrbIY0HXQ1yMhBr9mZpPSz
PGHN6Z5AimBhal6v8ROjJLMhl5m3lJZyPAK7L8W04sduuYDwq6IMGXmVsseC9hb8
uONXtsK8/BkvA+uPl0vNuV9ONrc/Wp3KslegAy7/k+kNlgay8suLMApB+Q/5QO1w
gIhHMwCl2j4CPkQ0h5rvD48ECUk+dqymlaSFTLTaBIeK2/5jFCqRwZj3cJe9jNC3
8lqZg0xehBIBCF/JYQBzRr5UT0q+mmSTnKtxxZXbUHsNkXTIFYapvYlITlZGzCTN
9GUMGybesuz9h0f/Yt+cimVcBfzqPaOQluDj5lvd/suOFAlWKzAWEPWSbebTGh48
jG5GUooMifu58FjOFUSoTfK7SlxNY8o7A55/kJUa2vchFGQfiN8rdABGi666czYm
WJsrgGHZ52HeIXgjinUAWa93azLAr5IZeP/wKQFh2yvdANRve6H1EoIl0QT9sfxq
ZW2OW+lLa8TYcSxT8f/pscH1G4AyZCm0VeIEyYV5LCxiBPYiyKGysmHu39iMyc+Y
HXfz4PqG3ZlkPhR2mm5s2b60C8hWNNUYS1BuiVwJpJgPoCGW3taC4w1rVF99a+Bl
bADsEmJtammbsIQxmZhtX851Yuu6CLOuAiow6Bvrd0UuFk/dFUGCRKFBtn18+18Y
SykYOvgGeSwSAl+mqZfytr3oXaENOfni22icfNjNntcLJttrQDffZpewxRBFgHkH
jXSjK/RJ2X/Csyq6eCq9mUEslKbTdVdeRsuANuZ35GR0vB/7X2TXDCx+5bzvsirM
m1IGhMUquRoL8KOU6SMJk/4+3rEbG4A0mA95gFLjpAOLIiqZYbQCceB6wPaKDoVy
udwisPXUhJeZJsrQPKiQxp7JSJR808iiJn0gPXVr6d4AVp/0DqHGmYfT4AZDFX1t
bZOBc4/q7//ura7syI7n5fSy4ayoUFPS0UskXZSLxe2qfFJp4BI1etLQbR3X0tJ5
rHGf6+o1GQuqrBnBV5kOM3TyOjFPiURQySOsEYOB2nxP6dIRMOp1sXhVLPV5ZPqj
RW8T4C7+vwHjz/FkxHQu5wPNu8cBEiarzRy4n/sh8tFTL8AtbDRs53dfPq6Kps8Y
btZDWuKvUD6fKVcrU6BDZEEOuAHbmECx/Ohn5ax1tw/C95Je2HNhJ/yYPWcsGK1C
gQuCPncPVE6QgSl7nXvE36IKhqRhI/8MbVqacQXdrYwCxjeSLdfQwfMyBeiBpZYX
HxzJdN2o3MbaB/W7xXQJTpTy/tQeYBy1UR3mQFlLCk3uF5zEUhxlcdjUaRkwNDEj
k0agTr/sFGeTrh42Vcfhr599z/NJ1/QwDX++2aQA6XOqZx1msRFGGNUk1DKq13Mg
u5nYoyGtXjpAOmvbE26gQgGClVilBrmQTzwi2wVjKqrsBKPkv1kCKOD1mtDfn2dh
M9FutaiylJ/MEMZdU7OAJ2iF5Y5V6bWX63QVFfiBhF8AsvWUJjUD24OdQuKiX4s8
J0wXuVJuw1u0itHIMZar+bJJUDOsa4LRP5FkzuUhQx79Rq/FqdrVq5oMsDetIA5d
xH1hLPf2WgHPTfFDPZxEtcq/9DzEnZwSFjfplxzDPiYCcIKeO0R+0RwK3w8Yjo/V
NhoV1GFguTgdRDPfjD3URBGZZIdB5MSsG1YkAJI4jq7/EOPjE1/frxv98o94KMkj
ZYatecqJpLUrwT9lnlWaiYO8xMTwj3Vg9HPEom3CFzWd/CCBgOnbOkcFmxM3j9fe
3K5pfXDdrDrguW0hkXHoT/TQz5p2rHVwGkULAuzgOB3vLTn5ja5TPrsEP1mcmdvv
+AKYdVY/DQfdcDs1Dag6NG58UKtM6PhNGy3bh9pT8KETsJ1Scse5v5XWF3EfpQHp
p7qWmU/18qryx08gkbbojK/vc/Ugi1YsKBAwljHDAxmfg1goc0nW0vm877lxNp/h
T2vgpEnanopbIhPomWvna5XUc628XYSH23NX7EfiwnUdhuzNpPylxQwouQ5/uBUw
X8FprpZDW/3Di2OWfI2TrBpnB7si0Q8M6kvkqOwRb7VzEpRkiZWjvRea8TygffQT
Cxh2uefMO9M7azBHdf5MjgKXXs/4HIKcQiOZe2noeBujmjamIZZd6Kt7XWIykIVJ
eNniBY5+kzZfBixYycKzXb7zxM9WCXbyuh7ftvm4VjB25VRL5xCxW2Ct4D9KN+ka
o2NhSs9FSq9sLybBH2QAUfK7dDqXz6aKBeZaGRyhbqPzUe1LUQuC121blAdAFLwz
WunWJ8X7FA1gBbkWYBT0DY+DFfPtDOXeR0T4tE50GuhBfGZqodC2WYGcdBf0NnXQ
fPlnmLcR7xnfTpSSQ6Z0+G9MnyWE583UhUuanbI15fY/g1B1tMQY64W+axeW+g5+
sHLPMm53oKdwAOZt1sTaetQmQM6sZjreJH7W7j2xtnp7jQ2Wjs5U4FSuB6E1kWDX
eLjFp7lPijEzLD+cW9+yvZy64BF4o2gsz67k/ohEgGRclnfqaygTxOAg7rUTHyq7
l4IZgijfQQkIIx3psTtViy+VcFJ69obLTaMBKtQgTuh0HGjkoI2fsJRfR/tDuJCQ
2Uj8EoxgMBjmcNuqOL+7J+ovnfhsrPTNWfjPmLw5DMA7OFjnXIxS//qw91FMjZkh
+/zkQyRxAARfxK87cQAlxHj5mVYL9VXIcECprQiZgtElvR/4GQ3vEc1UpsUOXVn9
OBKXcfBsUYqoWEFaUkfvQXB1NtTNzzYWGKLluP9VFO3hAPeTXo371NXmKUUHzKOx
ghvANisCvDdFTf3oY68dEsZ+uahc5x7bTb2ihQn+TIF6WcTJLQWXqim9zb1e1+8Y
XEhAHS/19pYItY8d9rS22Gl3ft9hWOMxfLS7CWl4xGWgvPy8gtuJmgQP7zXkW5Cl
zFZz1OZI9qtIMl62f7v967r+6YnfQ0SPvhuLOiCcLrhG/H9rmVkCoE7ZvEvmWwH2
I3byeidTiMy0Ell6ZgVvaJplJ5bqpwC+xVZf5lUPnYLkeHCc7Vb0LKvfurM70E3m
50OC4wH4Z/PdM7ml3Hz0FXyNVZawYt7u8b7Gdi1sSSfaGIwhKX01v4lHJ6lyeNyu
Ue6GpLEw+w9pLmNCUQ1CDAXP97yLOlM+EUYTdiB58aCScG/3oOwBgAoVrPuhOl/G
AqeV2ivqNDWTP+5n+YkGw8wQtbJMaFa9jJ92MZ+9f+tKD0Um55PzeUJhA5+3J5Vi
Lix68RB424YkFPz3FwTAafXk3m+r00QlYW5yXBcnq01YwRbQjPq6pDd50Bz/T1v6
UNHFycCpxqAVnni5RAqORg6Zwt6h2aWZytIZKen7xFAKokC3GDywkoVtnpEz9uN1
c8wqfaqeq0TK6TjP/zzMGoLlWDj/BNyAPs3UPxYf4vPfhrDDtttgYy/V1ArZG9sJ
ueBzaWjkt3UzaSBsxeaBSDL2ZxmTPh/k2Y0RvX4h8DTzXOtZXtpLbNTy4ThWD6nq
kgTTKptZLExhtjLHgY22suIqtpfjYIduL1gfHPLGzGw032EjjrTUhSeMdFytm+gr
DLf72qADkTpWD1gpgF/yrdo8AXD0RxwFqH4zP8XH13SjWmvenm054WCW0w2jZBcJ
CNKzm5wvmtkvkZbQnGi6rJ6u5968XLRhxj6d1HMm3V5ld7TfvDSoNNsIpxrUqyQH
M2tqqo/cAjzY3M4oZmkXb0rRTuO7l9yYUlzA0/thsyx6fXoGZSAigNldZzspOGXY
L/BWjuHZP5ND5dsBOV9MMTiMbSIQEFoFGH0VJS3UgMuWAKCtoTxa6heJVT87VFOk
RcteASfO7Cy2kSWCNdN+/jqOQJ+kbim7vdKjyVAxLJjWJnfvaazmXqAWLXseIlXM
O44nhxepMtnDmh9Xrm6Hm3Z6dpcw3eGAfiJvQB9WO/NKtlAIrAHI9p9szmzx7rLY
daREKtYmAfMf53UVwew6QDBpiMu1uzKptcB+GypDTJwVUgdEaU7DwMUtpRigK9Oe
WaGwOElwUhAQ2aPemk+2sGGsq0WzlB3XQywC9mIHz12gMKCb8xWC/b2jwMatLj4r
041hL6xf6BDblXruygZQ8rnajg9jRFZryiLozONHiPHBYGFC+Y/cic7uggJkO4VQ
cHkL372Zr+DqDM3dylBQQLbWafLOQ7Dgp7dPjnFdDdTlTzQirOSbOWI7weW/i0Do
kexTp1fKgOBG/lsFyGJxuuI383xi7Psz3g2SE4pD2Sl8B/VZ377DULHqo04XZj36
tJn+1D5AaiHMvR6y8Lsix+Pe1GFVvQsbDY+t6hh12SSk8uAfQ234GJ908ePGw9a3
RO/PZrWXrFpkMwSDEa2uWn28CtYLh7hCQ6AsUtjibzNT7gh29nqY1SKTP2nyjlGe
hLITqixpBeQV0ECmcq8qyD41zZ58U7eB41YXSUIVdWD189g6cPkEFR2Kt+bznG6y
LZRcGbacAQW236H4Kf93RVZx1m8GiwzroY+21ICLofy0Eq3Txpo01vpx8aSFYo5d
L3nn0bl87ty4idb5AZE4ckBZvfiWn00AqFNDQLTY8FyUkzJYPGWZlVk2nZnFBxHJ
qoDAChwZb2FohoGSuC3Eg2iXiAFMV0rjEEbpDWBsl1sgdVgbkSHhUhUVLs8sjVWL
3L1wosnGYtT2737QkP84DyYZEQRJl9AeSn0kkndP5SYSXcFLUMiiRGd/q++mz927
3rxsICax7xID6/qpL1/ZSUWEsKaenfcKOLDxmMd8LhbMqTworleUCS6JJ6ZmqkRj
1tbq8/hmB7n1Htyye0iVFCtH0cCPmJX7BiGp04QBYJ+nttmXK9xfwLxn5v5FsjRb
w+gHabR0pN/ICPfx2fu1mPkPee7mptOqcgKTLpfykl3PJDV1wQfWNLxrO+VZMazs
tdpwxsh8WUMRX9lIUKDznCQdii0eTpygMbnY8RjjdGJh6b1iCTdPx1d8oJPdfStj
S9oSaEjVGEUFasqsOsgW2eNkCWWt6VALpUhVYimoy6bwP8lLpxp8wGylHXltCj8I
o5f/fFbfqY21B6ovsr114cT9EnbWaHTN/cepvA5pixAw22eUoLrowwTW5dv8xyOu
B5H/Wi/UMm/QFZcMDA9LvU6mCBl9aHvtmMSuXabC9PRXbSKidD65JhhCqyGmWv6D
rCTJd62UfR5RGGY0RJBQqSvKiwrOcoY2Zr+0bHoAds8QIqMAz1fiOqOHPDIenAta
/2yDeD7FtmYcCzQk77kWSeJHK3PBRaO7uEwkc0Xct089aBnxMWRIrqCOMmMWcZDz
/END+RyUuPzudQcMB3OD/Yq7t/XCCuFUe9a+lDC0E4Jffe+gDNeWvOWFOVDiUSWk
RsajJwZR/Pa81Qkqush9H8Mjb+nYK+EYazfUnRYuNus/JoKMOvAY4XJPVwyJ/10a
GzDLsrLLrNtrRX5TsYk9AobdMRiN+ZI9YU0ko5OgVvc5N7w3gLkzZZV/E6pTj5xO
I/LXLh/tDoTgLKIdtLMulSiMxf9sP0BzMINMMkNTrQejj95+AlgdicSDRszBSpjo
OjMe12wv2Usk+hs6rLc0d28LW4s0CNp/oS8vJSUlArxVnEupe++U66O6l8wQs4Kd
OXLknV4D3PWZMvlR7bipiCm7AjnYsCuN6R1HkygJonajN2ofiAMJntAzpUlScBkL
8KB2JA9kZ7oGX1JObuAvUjgf9nngH+s80Z3SI32EYlI6N+/IRkizWS6HCQzebEhw
NWrPmoDPVrTy6jDnAgHVFTVbAhJknFtvDc9ShcDbblYSuhb3z6WVUYrGTSJZdq3G
elM47o3ixz/HTEB/hRuzmHl7QSqmOwlzm6xlePQdCk3nBzrOhJ/IyNmj13aomgtU
nZPB3lABkpk44kZgZvCxKH5dodtvhopGx/b8vvmRbwiRA0lOP+VUSSLFH6b+k+tJ
cySN0sIrKJkBIROxM0PTsf/OMmJif1TpXi0C85/XBDvvlwMT1XTeT5mVzknclZv3
RvJVfcEuH7mXzscY45na77tU1VXns/tq1D4Bvns+tdDRk5YSY6J7yf7g4BSKVdRp
NuhxNMd1OL+ylZ7nGznxTolUpvHy1OO7ZzdyaYIjgAoiiXmhqE+Mc+3f34EP5qz0
BrDIfiy1hbU4A8p2z7AAyJzD0u9TM8fNgmz+3FjolMi8DtfWRSHv6hpz4j+4SIfg
jXP8oFgQZ+bxNhJOelIWaleFznkYS8BYkWpbdvF3eoL88JW1fmiwYln4GIpT8kEL
zP8H+pVk2S5jHRoCOBMJaIzPlP4Tu8XrxwMII/sQVWuZZswm9djwqAeZuGuI5zCR
CdcZ6MMarN2NL+pcfsN3mIBcTgG73+OMk9EvAUOU1qaVhv5GCPSLvJkvGLqKjbk4
sp4fTaQleVnjL98A+VoA4OIdRY8YlBx81mcijFslhMJkVlMO/xLKU+9YVM7j3yaT
N7gYM5MPV09oShSifMgQB3UzjCO0q+qMeAHRDOtaUWQ5xcKlth+ViF4SoybKgIni
xKkBtzYEgrDRXgn6EM27e6PXXcM2EiyuRhnudD6TcuIzwxvTqdjaBV1TaGmBwNsy
POSEgR4UF7CWi/sxpxWTCNgdLodS/lGC/zBDPBgZppXm5mz1YfkrAttbNrw7EYCP
YDUk4w9f4fSBNFwj5WzUPuR8pBnYNVUauL2Kja01GRStCFzfOmWumvDiu+0hjbY3
Iw3G8HpzNryDlxqBQS5G4CkjQg8SdgFmTVX9ggSzBSSewP1Wdv4UlPPaSBm/9uyp
n0radUO1fma1kbrjaDzlY1e9aTkYlVFMtKm94Ft52Fqu8cdBSIuQOZVnBsvTJ5Bp
R9DfPjQvLOyP0qyoNKmKTP/C+WjdpXggy6oRmuBvwEl1xgz5qIqf2zgNNsxvCIMP
AdoXhRN86ccM3ttZFrdh3fJIpfjH56N4ZtcgckEM4IvX/5Gv9+uW27z+bsmLiUN6
BvHmri6loywBCWE9s1nudQOM92X484szbWdRoZAYMxxZixvhHYkcLETwBgAOprub
u0PydC33YRqtXpQn+HkVBRD3cHL31j1iTKMVaS6PFLtyX2V9S9AmqN1mbAtX+V15
P2HgegwkzC+g2oj2MOg5eHU0hFDvCMlC9QsoebQuCLl2QnDVqXQajw6iPkJjl4zN
dzJO+JaofJhhWJYh2Pd5gdgheBwqqL+uBdQ6nMyK7lF5bZLuA8NQIeduZ23B63Sk
A87n/qHIfYv+zU5AB+Aq8z/Juj5BwUe5WyrkMsKhKn//clcIC7hrvQGGtfS7+aJg
pYmi2viNlKB2UQ2enHkvi6QaDVfz457aR/z1Mf6mRBSgOCi+Qtrns2jRJNGqrXyz
STHE/R43W3Se8Swxv+sY6qbgoApVFuW9KM6H/rVE84Oxk1f9AnL+1HzklP1EfjC0
ANQcPQ3+BX8E8zZzW5bHYyX1MT1pc4calmgEgcyNWumqvwIQltI24FPFjGPBI8ul
1bVPqj4JrHoPirwu8uR3e9b/3kljFU8aJf0uUe8X8b9mdgnkAzaU3lW7NhKCNSXI
0jSJBBDfI7W0345VfX2LdIZiBc1+yjNtQ8p7iZUm6Yx+YyVqJjfI+npyaBsZ7leI
FLa3TfR7AatTX1XMQINx5RduPDjMRTjN+awA+mLObRoCcTTFEa4nRsNMalh8awfL
N0hVGeQDl1xtImrstAPv406oqlRn6kFEKhKEULbCH39Br6VzV4IK1kD01DwXCDoE
0nUrxlfM0IaIBakshUzG12NT+/D6jqyAdhuIDxjY1Lsr0whVnWZfCgRf6RddVcET
fR4OKO70Fl5u/V87ZKG2RjSlqQsufif5hFSUbnYjEVVxzGQt8+PPv5F6vLgisl3r
39PzVWOgRnaMXnNVVmZzrSsBO2U2qfr2b6FDGYCTAFTF5aF80iyASd+bhE6mw9pd
2uuM/8V0Xrokr7NoZZKIRcf6NM2inOXGbiSYda74BJVktM3ACVprKpkTmGnJ94/8
rG8aLs9HoGqOXChWI9vNhsJlBlyZu+l292XQypj2bIOMoKJvQHfgyUf6o93rl2ak
Fws+CPXP68Cr1iBNZ0xNyfhfhwKdzy8O3VuaWzyIwV5r15b1PzktJKPvvPKmWMdW
K0+oNpRuI0t+MASBbMp5HLlyuqYenJViqkrJXrfSFoZXwQb8SFC20cHzCIvCqwwc
ht0nkaDiznFKBYlHQBGh9GG7esRyumuXGkQeX+hpPlkzzxICukTOAFHbdZeVHHMy
fBjYsYavFkc57VHh8PO20bFjtevxdyEu0nIAQDiBhCfUwjbrIPGLCwmpxBEEkp+6
herZqYYMld/yhwWbRUnijL2AQ5V+r9Yyl3GjDhYhdzDgAspHnPYFrRR10oxGa9YN
2wLxeGzs0ZmAnXzzN8z8o4ksmpQifUH2wIBgkA+ck4v/83LVkB7KZ6XRgHOXaFGU
1ll275rrs56jpYIrgr4vLnXNLhNWgSkctQ9Wb5TEgAtt4hrPw+HohPnhkWAgBO+Y
CzknVvdQOF0/BxfLdT3hQ2z44Vj1yPE5IIKgw6vCvdFfBqQwmkswm5DIf4uSKmgH
UoSHYnQtNKEtQYQ3SqgYWEnwzDSNKhu88u2dE4nKdgA1TX7h5t+2H3ytDMJNy3zM
KCxQqheYIwKH2PuyLoqIMnCSgkCaCNt/JAnSL7/onIIsTDcmmTD9gB+iS1a/b2pc
P/Aj6+v6i/SQbLHnxiC2mnFL37t2VLgr4Rh4gjAFuqlRqH0VqHPRXtHWQDwXUZbr
d25huXSr3LXEWoNBFEn3y2/IDDMZXLwH4F1S/4InmqicrkKiMsTb1xV8U6pFgLNS
UrVGk0C3k/2lFdKC8NSWYaYa1s3Q4tAdH87ATCSJ2/pXTwDzMBSmrVLBQA1b2ssx
dcEG5yCXTmAzN7wNeC2g0kE8qoSOIt1+J9wKcrtWJ+kO3GYZHkiT/9rXeDREOY66
8HqM/7PZZ9yaQnk/HS/GhS0L5W/lZSzE0HZGAfOT8Hti9H7jcXXKMH/der5qNBRX
zeiO9hcnNh9q2EYf748kwAlsFPb1mYSzKzYzsOlEOFtAZhRuaTNrOdZNadLvpuFW
CFTN/dZ/WAmGIoLDREJTrBtR1W2qr9+7ktrP6KCaDM8WWG/IttY+nROHGWMxTwTX
qCrMKGcEEcNHA7dvfo6C1lnI4ZNY571gSiaqjPa8Qf5EnEkuchAA1jHCI/wTwZuJ
Vjf61+s9HmKh+4ZhS6ujV9am/W5I1u9b2lV3KBg6eRa7UGbItYTVSjVK6OLNfAmJ
rRKCkTqdzn+KEpRdNBXgt+8uK/nmUVyEgTRf5MYDnj1X6RbVcT5V/guPkJRNflpe
a8wh2Gmv2PZcYFeB/eMYcXmJPV0nNdTt422XbxEBcxlNBeLiUtYSqgUPSNRN3MXQ
rX2V6cZ2QGMRqjqH1Xc3FL4O4ratp3Ppd40MBl+NmlPzYJSD5RjqIUhDD1zEwsxC
wsxFDyY/z6MzqqlvP6VCHfJhbnvc7r6xqwOY7LOpiTKJhthOEwMIqEeFP7QmndlR
t5eeiHAON5qsSavgOO7nU2BmLtA7EWF+hH4maBdhQWoskW7N+soHmocn8ggmEspV
ZaWRgwY5jryGtb4HtebAc3iPniRa9H7RBqhCYFIjvXDWOfegGvg5bMk/pYrzD2cX
DiVAIco+pzKF6uxp07gzpxs5y0YKbk8Qc1Eh/hgZyVx+Il5oodEALmHSp5eze3Ci
Cm3fR74sBUrbVuddnQQV92pifqXGjXzTtn9co48uSgLKRjbsHqUqNzstRP7kVhL4
GujicH9zjgzxdnaJ/Rc8hAzuZaemr/XIr4x34RB041fWJZL09UpbIWVbiDby7xOe
bpIikdbNc+hkNqAklOKzRNuNRomoV0uihLENhmLhYHFnEQSyVH0jemAs9Ka1L06x
P1XMTe6HMOVYVNU7Gs8ZAOM3uowiDj0m5IoJ4jeczQXkOhMN/ShoI1+plIu3WoqM
J5PofGbdyjf28Spj89JoSHfFDroMb93BoyNLMQVsnbf6/P0s65tZafpj2l/QPgt1
qYTCVgtwkhH225QFEBnTtEro9jLHRUh4ezAj4x/lmKbwIdHxyE3HpBHZsRhITwKq
vQvQ62uq6WF+HuFVM7V/neIyTcbwS9+nNGj+hw7oXWYF4iwBVpyTfcdfZgocuY3r
KPpAsi1h1nhBmduJoqzRsJkj10LPHTH7xe1bJxeKbDXzT72kFzf4HoyqTJaA81yy
hRWosSMDniPUzh22IywK5m79pK2DoeL7F48114kU8dbIJRrQwpGIotHb3k88bKT1
C/K1Ijrqoiul0xtlgqQ0Z7M1dYuVct4vTaiiNYR8u5ee9RETh4SSK+nTqB4oTWMI
btRuRuVc3x/0sNDJMJjNGCdpSB2KtnArEUT/vz30hqUcgKml9meH4410iCH5/kop
LYItgoEzlM/HatXB2lrp2/aLHqDBnozU9NuiAQM6wzgARRhF0q2l1Zf9VqwbOc2A
LqcGXlX7W4QTNKOh60WjKr9SffWJu+K5RenrpETVCaHebHg0YoeV2LySN7HfStz3
gqPXHKEjhro3paVmXSX7IxVFGYZ2WHwNPNuud6B5qQSNavdQs2qABvcRs/gt6xZo
9MnyM/KdDHSC3PQt1/8ZvZmSXEfkN20CXqax+aH5u6h2krw3XZGUD/Ss2v57GtA0
KxvKF3JzfRoaEnoTXKz1oM92Ia7e0MRErAoXFYLVDg0ic/s6YKyERRkn+pHAIHtK
Awb8HMTSg6ATnox/GIZveQoISUOzE7uzgSks05TBzUKEONmqozxkovVuZhewJHy/
PYx8IYIhKEeRmn5n2Be+AdtFQkibtah99WAEoldzHy2WnzYhNdUQYGsGY9TTS1J4
+vl13Rh4gmB+ssvY8nW2uvO2rB0tMzjbl30EWd7/lgBuiIG/1I4qrWDFlk5NII7t
9dDMNsIsTjZgznywaH3M4Rjwf1bkKAC8seJT7qLxhAyc8moQJ1SadWXeJsFtqRbW
Dw5ggG89Teg3ByNZMuhWw6JRZTPKVxsouVTGbK9kTn4kI0em6dbxNSUad9ZcwXWl
PIHiK1piA9rhviZizDcGlPibbcnx44CZ3BbCfohFtjbBUVZL3i7YF2Wqix5l3O9q
0+E6rMzDxwR0eG6f2a1u+je4/2i4XfEovteuSUAj3SHU/ICzgAmlteJjmuteYhE3
0aKFmpypj4Q0MzIlwfPLlyfrmotzACZ4RSH47THG7D2hNB3vbHj6/4k1I/Rrt3r6
09IqdppvDu3Y7ghabQNVt02Qub3h64vu25wlMiKeUfQIjCEDAQeSkRNr9W0782u5
2ErGxlyVqNGl/5F+ew61NHxt4ynBFRJyzK1L6lmbWoR0nCuGk3MIZGqcqRMqCiGC
SLGpV7GNgbSVWOWKrkAvhQcmuKT0e5wkCrNADKXgYZjauerKtFbedNqTUJ5v72Gp
7Our20jTtJxbt+ZKhRmW/i1fAINqKgCxw2Mmoie1BLqWGxMVNv19ir/m3r/XLipZ
lFAXQNllhObM8Kh2wsWkxONXWAgw9eKhFDVlR2IHjClB0dDb5yqI4cwn2abj3ZkN
mfai8EFDqXKoJ/vxd94qeG6kvUCkmcVMV+Kl53nP6nrWg1rIMiTi4F7RqHNYgwBd
KBRrWQ53wE8yLmwJs5HKD1RCJYH3B6qsCCJyRPN2VuSHTOb8jfd1dPjWegQv7xgP
Zq0Jtu83RcgFRCyuusU4mUTP9BiDybaWpJLSS2qp7DESOLjOqXxVzFSJwGw28Sll
r0wBYLbHTfbEIxGV4c1IZ4KrtHRgFst5+CZgUxdvYVnID/4yWkKjaDvaHpgqECHh
jGIl4mVE8ub4cok697wlvVm+U24M1jLkq/3LJEqcpigake9SdPcKQ6hbUW/pBqex
ygSPs8ZxFIAKR6flGafVGsBaHzQgVhKlcDYrWNk7NKMd1drOyj72Oomm4xvKUzQ4
pt/xnibUWjDTzBN2mgMPMVnhmol48IrMZp3B4DGnY6hMrmSMbGY+qlcKM5zdfkmp
8ElN+teRgEyhDkcIrr0yb4/0JTLMqsdiD5Q0lTnhQA/njm8/KxCJsVSFZTtvavCh
oTmpcibZBC2tQPJUHEzow5wWOvVEbyjA+D9u1rmJ2CJNrPI0e/iwG8IvdYxSkXIy
buVHPwLX9KWMnrdCalszTr6lwwovBTDdPT9FjNjI5CE6nWoU+v2noLrh43HU1yG4
StvGAUJYa789Y+SENc65yVKoKThe0OYDLHnJw+mhyowR+OFIzDhooqxAdEfe1y+Q
P2mrzDBGP1Qx9gRUhhC0IWAc5esGKKzymk+Zjf52EF0XZX7r8w5HViSLh2OO5349
8dfNgKbKdljrtztB6yw5blffywq04lJaJQqVWQnfWxASBfZ8zSGJeCEcLSnJ7vO4
xysrkiEXYQ+QP7qING7u+RPkZjgszT/vsRaSW+SO0lXxywhw6dQsfZ8UmVcHkjye
4Hou1ZQdWSXMin34Kq5zQrbGGbfa036AWweF6ZAtAGrhVNUKSG5IOKTNI89w9Zz+
5f8cJHNAyW581TZGU54QyVn067ewgemYJfRvbfVp4YSiEp+7T+1FIsbPylJIy/fk
oPvVp5Tiqmp2OJFA7g5hTWWaqh8jMA/VlR60dUTZCH7hfZg8JWLPzMZEBVxntW5a
4AJyRDDkv/gZ762eJldItlrQm93pgOPIWdBl05RNXTSJOCko1wDatb3iixciX9I9
TEmUPRLRfK1XBmMLQCuSTtuKmaIx0g1jmTHP8HGKIkI+2Czx5Uo3jUDrIzh2inmR
gSQrCFjdirnZMWIjDmMkQLky/B5y8jmwtkx6hRpmzH5NdgzYlJitJ4VlWCe51AYO
zxZik+HzPm0SVxkEcvtSesfunchxuiXmb3oTZXDNrLA9UT56e2FBerBL3O3wU3ud
ZCzjVZFIC6v+HzFYY+Y2zQbZYSZ99ulVJ++pWKKSRpOHzwnybLlOV8b69LF/pEYo
xQpVcXG7yyppesw6ABcs8CTaYU1/5Qc354tifc0pn7imRD0nFNHYe0YokKX/p9gn
RRfcSVd/wX0sg+V1TayNjLUg5jFwASzLDMG3heW2OfM2/FjZD/hxAZy/qnN2fLoe
WAEQwByjQ11kBFFKYdn/m25AfEhDe1+Hk6VtnCMJVg4JdZ/CIEUri/jqhajxwC45
jlY4cgzdhr0s6rajTiZrXsjORRZh56RF1vsjmrQMi6thku00SMfb4FDWmnW/odMp
CxhEjwyvm6Ux9awNJA3d3ghlakIjg/wKh/Ql705vin46Mck0RPQm/hSJRB1nGfHm
9JDrobtz/BXiH08rqyDyB6YZ/sJhp9pz6PKJhHdF1VieyWNWVbfN83E5COi5gJZW
9kws4DKvxgfmXGkHWssvgqe/OTDZ7VswtKVHZCdCzCGfgxdh+MKjaYxbj2cEDBVP
vdXREQYtb8zs6V6RcEjbYWv/2skPiT4WM4t4k6AFgdnG/4wpo66z8D3WOQPJXP7/
prJqK2IltD5CjpMuuZq9RS+5SUDOYrM7fAz7FKXErRQ9cnSIB35foPAfs0QvZoud
SwnqVI5MDNhlU1Iiz6iPN04vgVIHxG5+V0wwa0MaXnWcvutOQ+hrtVJwxgwrbtjK
WLcS+8/hXkNunH+vbTktAzTvAy0k/bZe18XXc/g3/LF9Nzgj74Hs11gro1kdHhbk
IvDQyfOVtVpZk+61N/wS2N09vrW78xoF5ow+MaCXrfDZ1vYNg6+Sv89MuE/SJdIV
/UJvOTOEuv6dEH/M3Kt/6KZL/ngqhu+Vzz50GpZvo2NhH0rSh/tvsHkZmfblLWxA
ggmLZm3taNuzWvZDddM9q145whn6hl3iB3heo8Xndb+gCmBxUB4lDjkNYDrfxMsP
xvF2PHBfri91/8ShYNFOGpIlbATSesXM9m07trIxV5oCHGdpcGEv8rBzykqulJ1o
D3bRW9qBsQDYsG6ucssdcgBm05wTc5e0WUMlSYIvs6JTm47SxKkvCrLJiV3Bxm+E
S3800hF8J4GnVKQq/EeH40m5hoWz18SShBEAThuZIoxI40tjfj2VOGUHkxCYGTDw
NWGYQRSGBaTYtZTVyFcBZEwCOVCUUJNBnWrz6GQpwDb0KMfSdaZXT+8IJ0R6VDW+
osCb5Pg/C+uensGXas/7RS29vjsUCyPa7OdpSeWP4i3SyIkADZTnBiEyHv1nTmF0
tn5aOOLZpPQdDfbYMM6x6XAe1L2ckqQ2dlrRocp+aXACcoTpcp0/iFLiOI7qnaa1
0S9ITWoHVN4tl9h7KkvzmMX7ATm2Ut8+mfjcXl5Nh9bwkt5dmB5FSousOLmUlZN4
aJxpJ3r+d3eqrwbyzPIXNec5tmUZUf5FTn5IEQxD82fan0mGeYbLDHUVIUaB9F71
uGZPASNpnVlwvzKSiFhOjLdTS+9zobm9h88TI33LI3zKHhxDvA2wH65yDCQqZ3yD
4w5r8mCLTlNInutLPt2jO0O9XofWXaOVwYaC1bIv225FFYee5YFjgIbaZYpaqbln
Zs/CwfIv2Xf9xLeLTx0gDmo4HsH4QVVoY/O6oyQvp1U/9A88NxxWhN29wROLYG3r
MDueapGbM13i48De1PoEPlfbj5Na2Kl+HPFCs+vnZzJsoMikWkNqpqa1ggjHFCh2
hbc5uegP18IaauXRopLjLBR/QOtlGribecD3crQ1AZuthliDThFUbSL7BBUvbOti
fJp3aAmqK0QC3tVDGHPb5dn2aDYvkLHbmxxWVtbgnW6+eIrdZwhGERjFBk0gi52e
lSwKCs0exe9BThO9ibV6eOnO5SNv+yR9dw93JJeAtXqdQh8hZQGfeYmluT6oCkVD
i97z76/RqmhxkvsX6tRx7tdUIHQvTiGHVbpbq4P7Nnh4sVU8DLtm8/gCQmiTwr8D
jWb+NIK/KhNGq6YnOzzmAUiDKGbIHXfoyi9ofHjOTwIOKXlkez3viPdqSLybCCGX
rzD/x2i0c220mz+4SvuREC7x/fvsj2plEiE6aYIKR3+cM4xfedrmvBMHU28bmYDI
3dNeoCtXpaEsYuQfY0uPONfaEbpJI9737tk/qwFz08TwI4BJU6qwUU5nRKuknsCp
kw/YrR42gNtkU4xflCV6WwRvPKCrUlg6ZumyjLkyfARWfNba8PpmDddBfBXb5d1Z
6Ql2C3M613W686gK/ZgN/xQwhnJILJlCzd4LtzhnKxUvL0YcWgdI9LI8/uecSL2q
HTrKSH32hPkgqU7ANhIub9KOFlG6q85NUGw5sh9lElR1KcVZ5iGeDqKcnnv3hRp9
6dYNEZUZKNyVB6u3NlGB1slVDP60giGcY+OpWPcBFBnoSr4GGOl797f3tVMBh3VX
32+62sBwtOxurNXTg3GzRtWecXwfpXGEkDITlh3WYoy+uzh6oOhtu0mTuvimhfdg
MHAFk+7WzFSsDqKVYToaXSB3TWCcwQ5waBKqU5dtT/sTwnos3w0TXoMi2Jbs3Miz
ZiDEVfOIioOsb/o2zWeHJKfyKbOAHHMUppDRa84ivzJg3VWG0q6vYbo9gUyhD0sn
IwA/1qx3TmW39zqVgemMwnWyVWBqqEOEq0tp2MRHQjYhUnTnJ09YQQTKYTJrSXLH
Azyyr1OWo6lWs8PD7Wxc61AxPn8oIi1tpLEQJTw83cI+0lrfjHYPG+ZNpVzBem7X
oh8hGHJK52k8FVmvQ++Wt9iYth5AvYzn++ay7UQy57fn05MqU8zgEiyiIwNvrRTm
3m4OlLoylPVI41zW2TQcdyJPeoWC7ukRHA0hJmFYsaziGpJo7F/NShsEpBbx4QP8
ZMm+uZHVG0sjKP63/QrD8/mODt+c13Up6/JvwfuJeMQFkzx/2FILUeYhInLjgHlB
E2Bg+ObdlHROopWiH4DwJpfc9JLbqgSmPUOoo+nVr/9hbixdPpQxYmxxzn++KxPw
Cfkp5bolF7OYYgHkbZIIUi95p2yS4/W0NaOtbfm4ssnoUr5If2APny8jrqy3KmN3
5HAIooBBFBZs++k2stALE2vmcTzR9aNdswbVGr7eqh/sBG1rrQMZ2CdziJJ3ptsG
cxBsABDC3uTQBq2TISd0SFjDyfavT+S6Ibzb+6HB1zjY3T6wjbrJETXzqSkG6ju/
PoT4JV6BUwsYdSbasih7CvcJIOqBb9m7kX1ZUeqErZdg5a7kOhr9sUPXBmgulHsL
JavX9YgaC9kOLaK1XTFk7rznVcsood+yq8zRLSJPd8hMPvXp/QKSOfeM5PVnQ73d
FwSXFcF7RKf7VjYBvxOlSOL7Z2Xn/yoKVzTB0bCtd/wdRERV+OVfaezdpNRPhrko
XEbdFHas6DWUEJWUoeYQ8DCa5fr5QqEoknhbPC/jR4fWaU3gzwF6dKLtx3KfHl2X
6h5tWAarbLAId3nU5/LRfyjpOf6G8F4W8pxpGRPZopTaN9KcLS/o/ioiCGrMt72K
/GBgMItdfUyiolW1IkqVDP8Q1x1FeRfi7kQCiiDsA5yvvC8hMZDS0cDwMgit1a7p
o45fwvC/QyYR4/frp8C6Mq2WFexEP+D2MH2UGzvJob4ZhnD5pq54zbSMSgdPPDf0
F9KOGfGVeFiCvzwFBo3PfX9GR+gGFfM4LoQdTF7vHFuNJ6O/7YjdvzL0ocGwHQ6Z
dOA6lr2s8C2EHxDsmXIkOtZO2jiGL1HSHqWeGTdTgggVxsriuFsvmfY7FhrDAOIv
NQpOlkCSeo83m5NESs7FmIz7XdHyLDzFuYf7brCeAe18JfQ8HUWRajoKXdo5w2kN
3aJ8P82iuR9NJUJRO5amStrIASaaJ8vvFUP2iQ8WHux2/tCcVpB6uK+QpatcxK1J
s1ijp2APwspyHFi2gbE7mALsneweX0JDx0fTzTuEybYZB5+bA85x4rriQGPPNaC8
fMswML13c/Kra5kqqIl7B8LC/gmK+wHJxJkT4NtSOA8KLWUqD7LSCuRImwoRz0ga
W3PcgHn9wz1DEarOBAQ8vAA1cf0sNcxnT9tsNhfZeSq8uUWJakeCz13rAUFw2pCj
vELPSZ7GPF7ugraJGpzhSZ5S5edNWu4Ckrxban40q2rjwJADLXjrpvz5L6m6fGfz
zO1ycfKDWyoOPZBZFcuGvC7UVq2Dr2n8F9X1GuKEB10xKXh7zhIN4Xw3JBajDqU3
+tSbZS77hCz+WGgy7mWsGmR5z3C7mCkCv3UoagOxKWMS7nzd9NaQi/dT/gMxKTG8
SYepALga2iULg4EYXFZe4Rw77BN+Y6TGFXZrIAfzTBjwaN1SJB/p2d6EZl97XvDJ
sW4N+Baes0hr8Qz4zTM5N3lF09QRJmwX5CiOr5nlq30r1+ewuYNi9df82YEEZ5cz
WIbiuQj1+DaxGM5jEg5Ot62SI4Z1BKqfFpiYUABph6+jeoP3xzvOAjGKiKjT4Tk2
Lt6cH6sC2mWz3R1Bw4Xi23/1rkEalofFpU1rkHrg4N4wy9fudqX0tFVcPRVC2YHa
MtwUqfw9cmLAmjmK/Nfn7hOVtkBnhc6s8Uz1sxhPirJGfRhDtocoL1wlOTN3dgk9
cI0SzCKXOCMFUU9gHWJhsAttvsnxRBt79zJwwKVw66p1iuQaWZ5j3W7fZDjElkTQ
oZ1V3mKgEn4uiBPPITV3Bsg3vLhjOqxghP5/vPPok/t9lT62fbFnza2TVqlQXIv1
1xeIProTQpvcKbwactTF0AyMR9lSMN1SCZgcU0XEmHNYVoObBIXWEgxGZCTjlKrw
Ma/phDagiRZ4sGtrhlDHBl2DinwqO6vjwp8bCgtSglwCdNte4t7nbXCQQkWf+ko4
JJaI9WOnz54oYrz743pRaE5K3APRZcOKHRuJHr1UVdjkmGZxcrUkqbmUsLtGHqDP
a34urgTn3x6K+A9lgrrz8yZYEcLeP8MN3oMA2am12WVJ0mr0TTQCYQBjZo9mARKs
095xABtQkc7gQ3wSWNmmic2hdRVYgA3FJqkI8JJHMmdFt5/syDosRbRqId/slwPX
K0aAgbcdZG4pQW99vQeAYtG0tpza6mJXfGcAxGeU11peuhnlYoTRYxiLn6j1gFTo
pbRQF/UgA0NaHSFSPPAN9NldEnekcxq2g0PLWo1/mW64z32Z8a2TMuRMc2YLv4DK
AgO5CcU+ZeH/03ZFzm1A5BcewjOGNekiUaJJ85CBmT97UUyqLyCibvwi2mt0DM4C
FdLEPSy5ozMo12F32KbCWenbnvkCvXJNLTNatAyn11NfOF0fGZnsI8m3Csi3JisU
LOBraRjBcg7YNNzk5L0xK2daVEli0hn6eLqMOALZT7FbcDtCNiCSwAcl/7jESwg7
vkIhLYaBRdK8Gt0R9d3CfqPJYAj38r+Ips9+ypHwUf0Uh7xuvLXBEVHDo4Ef3AXe
lVBeJTwjgaDwKDBaWOG5WbbzjbGEjZCKRtRA15VL2DwIkracDRO5umWQ5WW+If9O
VawkexsBS/lV6i9RFVAAV/AsUAYmnF5d63RAPC8cWg8DkXBuzwEp9IKyciP6uAS4
5cbyaNujQFJjV8mIJJoU1o0blGQ7J5SnEnBPR1Ik6hiyndWpUAijFZLeraPmmYRG
PkffIIad+R+s/sdd/TeV2Y+QtVFHiZiIMtTpE6nnLgoZ1ajX1K8A/Go74SFyhALA
gTXgvYQrSYTlnBZtEssl58IuM3w1Cl9DGd+p12nOfnXQpQhrmZ30qNZcISzTOFSb
m3/GLvuowp2HYcotmT1MWokIhaJoOV8KN9h7LCMBy3LYCzqRJ9e3/8NjtNCbSQhf
gL6P3grDzCMRroOiFjaTGtWc3Jql1KmItEvHiGcPK43NujpYKTkEt8oHVqRO8fre
wYstnNMLqbI+8BHgYFPo+TzutsPxd71/w7zr3Jf1n+HVBIPMmEkW4bVL9emPQSlN
8dXUhKfo3VDlCsNFSlu18Mrr/6p/d5EBHmFKLF0dTDMyPVECx5JuCnDXGvNCMZn9
jXC0GNny9Wz8S3TqZl2mxEd1EmeV3joBBmVQTFO9ESQObhIiN4piVpuFY+M/HeD2
7vkyEHV6Z6mtGY8reaNydw5pXo/Y70Wa1dhLzU6HlQ4m3bkV4hWWZCe5aUyU1Rbq
fr5zFQryCX8uWn0ZpzI0yCslArFGPQQxSs6HfzBF+5UtYNNRzpaGhRyl7Vy3+9Xw
lWY3kTWkG6j1qlxYMUQ1kQyQao/zzp8Lk9sh0MiG9p9mJPNpDoBbLpC7wGZVCNDC
s4GcQJegJyDZDoZbhwJfOXW0qJz43by5CiAmlG+Eq5Z8oBps+TOEKYAhyitVq4+W
Ej/AABEcp/vDu4GmQ+Bkd2BSHP5T00lURWWDpgROU2IC6sMRDX0/tqNshLeHEo/b
OJ5QMPRK+I2jJjPLXq5pXzDqtUOeX4VnINnkqR9dr7LkU06VnZQDvQ0n4orFZxsS
ddkJCVdK7v3uZuRLdYt3eGu0owy515nePWql4Aoh1P6P7LfY+XbvNGrMsdTcz1gP
i8+IMu2dlo3SyLrjjT1Fgu28TFJlKlkcIMuG67MRr7cCoiIqXf57pf+WpP4wWHB6
/Y8WvpymYY/FmhkNVTB//9293EuXK9APPHsdY3Vkpw2nprecIcB8WcS5uJ0knwR7
LGKSTs6haT2r4IsCUiguw+Z/zSCLyktSxKzvylN7O+yNxtlEXiAQ0YZpNA5rj1rM
Rh5JVMV1RwuAhLlBsf+r0CQ+UWT6u+EwH2uWtBAjKPyS7ZevDF9JEXIhPiH4tDfV
GsJgfrphOgbuL729gvbZYOvaDSlyw/nx1406fW1BqMtaRvKufpzhmdwwCULirINF
td1+jQVrn/F3Cq0e0gL61PJxziLYh8aZZRcS7Sqnbbya6OXfSKCTvkLagWDv5IUb
MSZVA4/stFUyHhOM72AyaLDcoUuOAypZVIanOl4u6LQnQRtbNWLokV6IhMiFKrNU
kOEe1UwSxym9c9StRY5Qn6kaHnkw0zffaKb8DPXFm/UA6QGw3VhKbMFREVb1aXb/
FPGl3SQYGeOMvCCZJ/WaTzM3n9m12j9Fmc4L08kVvY4ZYJDd6nyj3EEnKv/Tpt4/
aRIBPpUBx6RUkI36wuyiFnCvcq2SqMcMkqESDIEz4sQSrAKXNszgLofS7bQPU71+
Gfzrh4QnVoeflq4LjuqgGMdIok5ql3BLUxGD2wDCVoZsd269dhSlQEGw0GhRTJKZ
osGCDZ9nTzzDrJHP/+lrKjDGmRfSK298Y/fFTp/sZAp8GMXPVU8GI4PhfNsnT1vP
z8xBOSaloeIapS7q+/UTXtmv7CpgrVsxMcNjWSlkXXSK3Jp16Pq2j+yQrKEA8Lgm
s1LHtjwTmkanmckfUf12hEXqlp3dTpXMU98SejHP4y+sqiYjhChKSrm0SMuUKhdq
z7h8qXVF51Jhx+gVOt14o7Bn/3mbLShyvjOA/zAyHbvkZbscaz1ubfxJg7XBOKgv
CPzB8eE/gQ6bLRqUMKuoN1pn1/+cu9afIjT0NbYlfyLpCS2dU8EraOcUQGh9qm0A
CIJQhFM5ilikpay9YeHVIHH23xXz/aMLo/3hPtyiaucvWwr7qEyLZgV0e+RDd7fc
SF/2kY87wUk+05aiH8p/xqmMM2D1SEVe9ZTIt6ErTA6CVbDbllSRzKff495/2/Nd
y0u6tQSCl+no4XHI7h/Z5A7iXpxKM82omHGLC4JHsJd8ypZIUC2Him4/oOtOiqNP
RHFyAj8YTnzKx4u1x2lFhcYTRgdVAASrnLZlzz7qyk263BqTSCh+zb0V6H8WP769
+mZj7RNvQtNM8Obi3u4N2BqNstufxKLMcy2jb4LECkmvqr8VJhDgxInlvSb0EM9O
T0qxUHxpOBYn1SvSFiwNMHarhvYFPRfMjEiYEkJ09lzGy5gEzowej0uK9hweoImU
1d2pIwX6DP3Pyzbt241IGNIC/u5K/lt49mx48iNrLjiZUjZyVGIl2UAjQnCdmxae
yLCGcSyAAscODKUazAWTmBE1JFv/Pq/A3QFQZ/rm7VqPrvfZUuxblF6mK+GXmtAX
RJ+MyowsoxtiRBGwUzhMfF7m6HYH6kcH9WG74Tr9q48yNADNFTV1Yg8pWCqk3bzw
QiIW14p8emNFqp/WlpX346yAa8d+eYazn5rZbPfPzTjYAWm291Kf+JlyANHaogsh
ViapfXW0Y61T36vLye1ANF2CBYFMrB+fzmmDrY/PFDpshf9plRJDx9UpvAQ1Cmq+
VxwFOP8v8t13R6fOreBFG7xlaJbhuP+rBn12TBHEx5n8/o4Vft6uBbTAmYGwJVV3
5Dj+gRgxJ5x3G4CTagG36wZKXNz+oZkVf9ljkuSvE3Gnnk9UW3Zdj1KS9BXteorD
7gKn/Su6O89noKvVkqt/pFag0BJ92DCZn1HCM71kEyeUb6q3ZUPiDVCOBq2Qrzxf
CVTgWck6CelKXbPywIDzHkmFz6uoW+UVE7VdAbmpglk+12VdHHudqBB+MBRKLOvS
npqdlzZMKZEXlGxBzwpSPmVK4kRHJDpEwteEi4DCyL/u2Xv7llN+GbDQ01e2M6tu
bu6zbpvOs9HzFShxz8XnhC8lA1FcUta4SqknqR4awGcF9G7SZLRluodB4IYyjLUS
raD9G63L5ffM9IKSp4ZRfOjJijMmmn+vNGZ/81QPbGERdMbexVPQdsbED6u0y8Re
0ZmHzyUPm28pdGz4F9yr67bx5qjxYuTElpvkO5m8VwmBAjnidf0zdCukvIWeGM3g
CNn1f3BzZ9FyAfsiHruK2EAiNPj1ROCiYk94e0Xuu1nROp5Xmi3jiP10sdIDeL2q
f4VNLeWdz5pVdlRP7LiVl8uVEpyJS2A98bpRzWca4xv3ntR/Rfqs8TbjG6oYoMKP
kDqg1D22PRqjhvVyB7gl3DE9MO86YdQrQOyEZ0I5WFmpezOPeGE0s1zTJaHKrisg
l0hmWIPu/L4/z/j/DKAhjfu72r92gunzmg/g0ulyRK7HCHHfBpV7XuxpI/ssCzom
qTIsAwBzmue+b6RkuX0yxvqPqfM55B27bDBueD53taUgRvY8VGOULBexyXOy2xwE
gK6KJADqbmcCLrKdLnklCccTvnecrMSgxePKiCDE0i+uBeKSQXFyamasHXqF1m6X
KvMKiXdEqnGGhgeN1HOuTvWiEOqTmYYf8smwiwgGodrYvwmFt34u0KRMU5HktRmT
YyhPRJWvEn+GJJPXfPDdBS5m1XH8A++d904Lz5uODlGDqXh5mzPT0v/GFDdgLn64
55Lu069QfJ0XhSyMTjCOCkc3LxL+zqTu70I+8SSEXGpaXZP3Oo2/aLdyZEODkXTs
GxVr+Yh/Lo84c3gEiBGvbf9xD6Aj7zvy1aCxX3nnZin/l81ZKYunjgY+DNQsbvjP
Yt6qebpt9UQDhjy9+wpsuyJ1DF3df3cnDvJh0K3lyVuFMpGcW6mS1rkmOr0EgNxF
TfeAf7VXdjJBvznxGHyDTw33tRC7Jz/D+2hR5qdEGpzisnaDMNDKrpA9gC5fvePv
8K8ME+KyQaxfz+9h0UD8+9h7cuFa6Fi4smD2Yw8UZgpOmh5B6HPyF/PIeYpcF+Kb
dghbNUhWs4hAhqGVTZJiqaF5Bj1Kub2zzUOdZFt93Qt3EJ8nXfVvtEcfQw18mIMp
mHC+YdeJzthr0D2HdtOZq7/1rHlgws6zdb/f4fqUsbh6wpnCLD5UeKM5t+UNSLf3
b3d3crFs6gwXOrKjmh1cKDIj4832faI9sk3TFFnlr3XqPJ6QAQ9ZVvjJvV6mLvEl
ufyeZ0Gc6UPzy1lJH/uWijsu4OJiS/5E2v4XU01mEdGrK5V2aiHPDMOyFmqe2eGC
m/F11HaSN8687fVuqCYWv9jk4E+H33IFDGjZrYC5dK+0+uRGjTfFA+8cUDaiZ+CI
zh2A8qtJG3P8Y8JCm3aQe18usf4HyRANHNIb5JiVKtJl3hUsKIWqfnvRAETc3sbP
xPx4ApmK+1XuXt+/G1RxLdxt99HRf9MOfPtY5sGaJ9pFToss0Ln13UDn0zv2d9Hl
TG/+tE6LLrLM3jdxXRn+d7h/stMI4iyM15Ev3u6eyJ3Nf52Gjl1cqkOjFLnSUDPH
SuwxYFdy1Y+8Aeho0OeRK+uV5Su5wNTs1NnoqIT030OK+m9m2RPKzp4XWmS9s+QK
CDOCbvPfiUJHt2sa+NfIHWJh4iV3foc0hheKz5eqmS1t+1U7DlCYgK/ZxyVmAij0
d+mzxeRTlH6N6T2dLNu/l7FIDF+SrMZlXvozdOU+ikblZmH8WAWZ9ntUHOIxA85W
j00te8cuqE9dftWMWzfzWr9ehz0enihbiYIxR5zgYzlm2imk7ifV5b8J8pAERcow
Pa6NL0hAiSngQKXy1qM4qGMX6rCXGWVMh0c1WA3dkhFbg3SbvBKgmgPoJYnSenii
hxXbRSgS0TKcnyV4YrsMVxV6HVLJSFJa3pH3fmwTjxoXmLOb03QeKwtRwgdtOuFm
esrmkXMO5Cac0b+bzgzsTN+fFG5JxzpOGVoi5esalyTzWjxZJLdWLexDo0Q39+P3
JTzD71qJuNrp+jWSzGgaAujF8Wi0cZWXgzpV+U2vn/ipWdYmKNJZ+ssjhRMkqs/7
OAvKI+cBWdCIxrnzfHGdUKZdDTXJyr9A4PNgI/f4TzwaR9aFDQWD0YPlks5dwO+v
x4SPNdLfj1cG+W6jv9+FkiYqd9JgZiiVoDfOSCE7COQtbDxOj2hp65oFSHCwK9Bi
p5sy/JHgbd7OcoSdDSVqgjvPleJH8ob80sUIUUTFgWMssf0eUBII6cmLWbWFVXhZ
GsbFgulhC69AUWPSps3cmjkxglX6L33C8l4Dt7YVKVD7qYnxeRX2fwq3V92/miOS
TI7ksamq7LU4VZpRzUP1wtq4shmPUz2yepC5w3LnolMDDY6fUOPG3wiqWtmFJkK6
oDP/FuWx1hFbdb5KLqZaFoqVgAde9aLHEqhEiKeDiDyKsgiApwWgNW4czSgJ8Cqk
I6zA5QkedNuA9qEKNlL+s92PxaoFDwsUA98cCAYdsBGjEH9g2VYqT3wHvJMbXFWF
M2+bwX3WWtcSttHnbS7NEILlxPyPSF9JdDp+I83sGNKs47FcnVHXzV2El3s6l9IC
T4klF1s6IbX8zx7YgUKQ6z+YiogS+UUPKzt9RjkKIk1VApEByeOp5SBTiK5UOfHv
45XYixT8UQNCZLFY6RSvFgdEgz978dTb2iyGTwxH4soPOagwOCA2mK3TZNrfGgGc
DyvImc8QQGryU+dTzmnpiqHgGfBBgpqY/DQBr9KSAF7oqb2JnF4xbaHUoh7fdmJ3
AbywdgBZcZM6c1ju6HV7dg8JKn7fhGKlRukFbV3bBuW8vJpI9iVBW7K9WVZrWMUs
cn25YB7HQcrYfuYBO+2tQ7K8ZYFuk1cIWIfZXFcg+04bmrTdZwX+Se1xPMgNLXpW
OvtpQaFcGgAbvw71beAvJdmniwARyo29hQPH9rEacSAVSQHk7E3gUd2hiAacJFiu
hQymIZjjqXv1N+AL4yBa0nMmZnftly1ci5iPegTgWWpP7/7UGl0qz/p+Appq4QNG
RKX/DSdZ+GMYck+P2ylQGPrhWoNEHPUR55fTC2pTO3vU1VkIWEdStfgRyK5sBmiU
JP6kTBM36gjSVO2Azfla8uSVTbIrD6SzWPy+bzgn9ljU2ERHxl9Lk19TFhh70geM
UXz2oGYWgwNg6jRvPWrFm4ySxGoiMeUEe6ajlB1UFX1oLrOiA4TZSxP6+nW5F26L
GD87zxXVwqFz8TMCxlzyuoFu4vEyZI1iVnCXrnRSfCI4RskwrSJalDJ/OeBVYuRL
1JHlmFzocivWNNEDHc4F2N/TPCZMOEEJlzLxldMW36AfJT7vKbY4yEKGnyqjA1ZV
C/nv5Yr5Aa+/pQUQFhCqniQaDj3O5PStnpjdd1C43uDXsVyzLEGsJwdB4NiMR0Wc
0awkr0rVjoLPZ/v7ArnwOvAY7GOSeqEm8Pb+QE3MEC/DtZPNaMhTiZaDGgdePYz7
z88uCbm7QyqVkgqN0sbXp31OLXaaYLzg3Q2rK0EbbDhFIzhWbdYjS8C6DEqe2U4E
kReZQEzrJqOqByp8dIULiP2jEw88XV1PXNHqRhybSMndsh0aqBhcE1Lpkm+zkmA+
sg/2v+BYuxU4GV2bLMoycpSqexW5W3EYfyEsb7ZU17z+IMk/gphiYcPP8pn2/3NU
csffpSvL+9u0bbXB6hud3m4n2K7f8PYFoe96BjKjuoIxP3R4pz8jxNzDKXGEjibg
p728kTFvHKI7Lu4G08yraBSmUqh/Bvoo5ymWkwL/mb/NUyurWSM+fnojeH/T5pZ3
OjU2M7H/PC2qOcZUcNjJIo+hFj7HdPedpMJMb1tnewYmKYyNIfNYmfINpyfZLFvn
vwKRFru6kySY5jOfx0JaPGeVWAzwYU5645chtG+ikYTpOyI+Ok62ppyPqxXCCXu3
7MtzwehY8/2Lz+BclCYPkIk7ItB2aRtfLMLfMeP7mTW5dGqkH9dPlAP/WoS9Kg+j
b9yvnQR9dN6IDjRZyl+NJa6OZjgzfxY0IszYBX6DduP1ixisCF+lhKHBr725uHR6
4CpNl8WsR6Dm8PN45J8vLwyqt2fWjIRbiunZ/rLJfFrHx/slgPFNjOrDqinChqrH
CdcRWW+98O+CjEikayC9jqmk55MkDCEfQ9fqgENBPxfBftRk+JrieHtBXxDeWWJr
6VDD3Oqw68C9yTFhmNoTAOyyStaFZHwz8AK/YjWsExqaZo6lFse6jpG6uGRbZCs0
/6EhVGlIhr0Jeea+jDIGMuAyu2jC3pqlw99dyGEYLb63QekKSuAfigxWmZjZGlZj
7EW+BMnytw6vHSKd2KBuJ8Bwlk903LspseCil45F5nDJP2mXlbjMzCEV09yaQm1W
MYqcCN++XSIYAvrXn0J7lDGptU1MvhGRBcVKDagTLpvf+fe1gXq3gLiaHoz2FpVj
wVZXMoMwVZ/IyYvleIYVdqm3jRGFHnE3DJk8sJBR51x9gxo6c+I7OaW4GdslnMQq
MajCir4j8u9zM+82QOFHmslV1mTMVBtuciOR+ywgeHw4BIzHXe8FTFn0BCwGGlJ0
rsPEj1mQjJF8Flrs4Ly9Mi8yYBDcZBJeJZEo8lphJ0RVv48SQfPAJLhdRDOABrs9
eLaLNeQkbWvPZU6cC3t828Guocb+qEbeMfUQDKCR6RqdGTPsFmTgGTEgwqWUKqwK
iNmpZkDyOTUE0jehqsAIqZK5RCAGTN+a55/xCUw8HWVH5mhzBcLJ/20qtHc487by
6kkAkNmAk4pySaaSRMGt1b1tFbaGE381BKuTkN2OQT+cX2pPHmGHbhBhjPxntXr4
L8F5GjUhHDKmat4DXv5VuBaz/EFOmIuL6Z2EGBtPSDqqz9o87e0YW4P4/sAFkrNC
/mapWvrshsmOvXd+lXsJX1p9ru1Vg/T6JkTxNP5U9cS9ZSPHyjKA/AfER9bzIEhR
ULWeqer040+NMyr4KwJ2mtiP7B2hnnJw0IpPzl5SHR1loTcyY+OJZtmLK1XCzN2Q
MbXJABxfaUJMiQ0zhj8wFHN+V0l5Q2FamcCmHeHst89ADE+3+zLGfMpAT4va7bZL
P1zacb2rNymAi/R71+lixGEhk8bjTBaHtQ2acOgBSqRN3GbpT4eD/2I8gcr3Pw6W
qNFPhZ/KU31Y7Ojitbd0e7dC1JRbEG6vNqfm8Tqt0JSEI5E9T+foh5tOt4deJQYb
XOTTl7qzrTEqoAHlEYJ3O7yb2mgOphBlonYIO90E3AZwIVjhQFUuzSImVb1bLXPa
P0GL+nMW4ocjB6iW9umaiQLhu4n/lvAmzTS3Y4knIOgNcjH3NKNGAZoTeXHv+AsX
kYGhERHVomeM3qJl+7NcWhFX1WVP005FPYcSFZFjGqQgbYvLX69O5ZYbXqrQMuRH
aOE+LDZIHtlXg/KzD+dHxj143v/R4JxciNiejlOOjwQOQvoseIOFvnrsCqfw6Gwh
7clF9NRcdyOnSRJWtRiu3Eia1JSnGgrDJs9SEr45iOQgr3ZCyw6GE2bM7iFx309k
yaAEoc6yb1MarMwiIafeMTOzOu1sSGprlp31EhD4ipBHv9PaOzjK+5j5uwGV1KBu
bDvyXgt3bxcpOr1WxOWDxddrhQjfp6FKnFocGghs4+trEKVdlKLkkVbAVvDELzkp
fmjm9pT/SMJaP+GwmtEg79Nf+SyPGtYLqkwJcjkeo5SvWoAZfKHqR+d020K2+KX9
YG6IK78fzTCrV/E037YBcjRzMM92Gi7i4gDy15bm7Kl+vSY+VyNPFUZsZZX0Z8Cq
bLwcSuy0Hw5JJD5aSGNeEdK1wqP6iy4BybJJ4WM6LzrR0JN+vuKLFJhCs+A193lw
vy7i1fNI+OXgGH0u1RFXzPqFSqetcSqOR36ufwm6o+QKYfWtej3J6K3RaGSlyp9W
LhB33+absjRFlFMXx7HtkrNiAlz8j+1sizCt4Jy30G0XY/Dj6CY3i9at1Pb9E6oL
eSgSi4QunCXHrxJyVU0fuNPc/k1oYaml4alptHanIQBPjmFD05znsRLxNJ9+29kQ
+RdfbBnDMp4EJjh6XTPz7C7PoQj3HcXE1KSFphbfc+qYfUXAdqt5svd1hxZhZZ+M
NXLudEb6L27kD/12LLj/73xW4u8bzb8WYvdxgWNuo456NrH4xof0IhwEWfAXPWio
oxk91fcRp9FDvPgbm/hHDTrqetGd8ucR9c0b1kfzI4vnuNMbyx6GkJ4afaX9WK16
SPzI0hFBeNQLGJGo7DXleseyw77hUkQ61t1mkC3mxWctHfya/6T3/5SvLTc0iBpT
7fHAH16ikAwHzKP3hrSygxuqdG9BO8K03MPjd1ZBL2N4L/22hLmJfaS6lkWQpBTW
Dm4EgR8KKg0t8jXXOngpQn7fadD6/Ch8//vt+omnkxDBDjKfuAieBQ75ps6DkwWt
Z8w4NoZc2BtWYCr7C5QjhDsDQSjfOlcEfLKaiaUOP8u7jt7jm8sw9cwl7vska5TW
iHdA85AIO5IIrAvVPcUlRaKSikpMdWisnFhVOIWyUPwOh2FDf79PcLcpha7Rsqun
05sw59w+znoPYDJAUlN7WgjOQz0TQcNBur46LrR37DWq16VNXipb1woivz8h30y/
/7+VdYiTkQ1GTJUiWq3CcXaLACsbcQgVvsOS//0DCzFldrxYfvui+r3mSXYUT6aR
opv/WKxX3ZX66Er5fgj/4kLXk+Ikua6y1nF7AZqogsWefOYapal4CmY8HqSTBW9F
pt8q3CUTiULSTlU7gQkMu+5P3YsF5etnq9LwOfwixb6caJYavtuZmJQQXfajbEhu
I7tfsnfLmRoz+YQUmd4/V88vXhKWmVppPrxufjrAANm54PJnapKCs7mcYkT4vs+Y
OYlLvLarwseMOBRS4Y0H61oDIlQamHIhw57Gts9OTrN/Eeiti3wMJR3Y0f6tbgAb
duMroG35jneIRKd0JUX3Py8cT80AERmTrqKqULdxYfvaRixDhNNJN4zQIF5V63dk
c+dcrOzR9icrt60WQ1MwQC8CCKtrNVTEEbSGeYbS4DJgxZggJsvCyPHP46DivyRT
EOT82RJweJ6q1QequZOq86jg+kiWZcqEr5fxhJJRB1tRVZTkP6OSk4Gr3eLz7A7M
8ujpaCZlP95e0piboNDwdklPt2j6LVdmAcbXffs7qIX9eCY34i6KOIlswo8Gkqrk
f0KmWx7e5bl/qTllB/8h5EaF66QJJoymNauvOzy/qb0ToCmDkVGS7uVOcKLenFrY
M9BUDewytHFDLtpRCbA1WN1dHZcTd7lLuy3yqHW4BGmNDZF69kAEdKWcmIiqQgRP
0Me2R3epmhKFdeOjxpzau8E2H3cOrav/1hqtuVF7muHHQt0TPaY0VYurdakCBbIq
zPwM5w2JQMPNvoQ9TlAbAm5fG1M1nYjC02j/V5+8eJv6gqAaFD/jfCaym02b4cP9
S74ZNNKyc1JeHefLlDsGywfsskFI8JiyM7ax7jPUMOUL2S27D4HrVGuPMyJBQ89H
AGdtId/wk+qcRx5pDush/fALDRu6TxQv92zZVjh4cRdQIZfD41xZdoUkxLdfdEcc
Xqoc6JEg+AqDUSj3Xs7EiFklOUApaIDF2o3E+0+POm0eINngNXQjqImqBDQ/L+Vm
6rg1OtRjTfXUsKPi4KcypyeEIHhX4kOvWuA0+hxkF37DLYdfv7wHrN/FDdpsX54n
3QZsrhW/LBB2BV3PD6PrJfmzdqopzmebgW1b8pIiHUkPLsVXtAG8H1EQOKVNNn5O
M1E8/qPSwkfxDX07B+NM6jOnMjGkZxFASIbcfWwtGhB3FOFb/EFYvpTNfvsgw4G4
7pxg48HA0XzNBVAAfBYZaVTdzGTCM0eSHLD0Tua+cdCHwE45Yi8bUbC0IZ5L0fJz
rPUeLcvjSb/horVRxTL9M9anJxZXL+OQXFyDRP/8mDnFKN1Nb+9FWTWjwJxQP0T8
uwk5CwtZgpiFW7yGpjzC6ZmygbAfx5LCm7ApOpY6Ya17vP8u7Vlz3eb3Wn2CGjrO
lJFZekqqxFhluuT+0IeN3CIAmDt/uXDQQDqocrxCCuLtmDsPjDDbrMD/F5QDQTrA
z3EWaMpb1/qRK3J8bkhHANr0zOiLrpxp3BBmizYI8VEghFqXDRUl2RyKDuAE3DkQ
MfQYndOWZHc/h55UkuZoiJsiIgFbRdJxsO1kAoAH/wNW57+ZRWA/CRijfOC7pZm3
nZwrZI7Ahtlk2bPY7vX8uGKcSSQxZQgqYLyeBOpBldT8vUyxam+2BjapzwudNXnM
KN55JnSZy+QEQ50HPJ265q9BpM467W2VJtOZrvG9f37pcp6dlOYv9yE4dMUUCz0D
N+bNQZThE5i9TnjKTSW4MiydHJtQ94sAp6YRtgWiUqLKutXbNDzj3CnP+E/NJJYp
kAo/RHaKIP5bnuWzGBEOLDPpXbNlCAinepAxA4B7FahJ6M9lNAVMOtrTVBO47djn
Z358bjpBtjlJWnXH2pVFe6rySZgupN+mGpTP9qn1QBIV9Oft+2mRGX+iBd3aZ5Aa
ZtdK4UyxC9DJrZyK3kTLj/TRA/ZXw06wPUvQ1TC+K4ehKLYpRFpbQyx4WKeO8ZDp
rStSOH9oRQhKNwlqlu5jvC4wcgOgLJFG45qnSOwapL0zjrUxK0AJlDWAHOf49IOG
lhOS+Q5vVmlMXWmvOx7wocj16oTKEM+9C6BbXnjEGINksn7RvYOldh+agQXoraZG
7k74aWESNMTnP4RqjDbzt9XrNRwc2DgQwQVUFCXUN9sikMZmWcPC/oiKxUaBo1FH
xfNFOqzgeCg97NOTPO00YlSgSi/SKwP15zIUtej4XQVAKSI24yV/NpIBc52vBmCF
A8VqdfSIYArTqRk7P1pN0f4wV7RBDfnJfWuN3PxlKaMsL5DEbg+vMrg+ykaGCxHU
KVgOYB4gBeSZY3BWXrQoxsOCx0kFWa9aoJmM7gh/sZ7C7U8RsmwiFUCVdbWGouTm
swX72Ip2ZgXMHbf38TO2oNtc5GOb9uGh/kLt9CyBo0lWjlJP8U8BEG6+Ef5hkUFl
3Fm6iV0n2YgHmcNxc9OwdOPYoo+DFyyUCoyHtNocNn6gLOh98kM62FqV8OAKiZWO
G+ZtvR/+brCfTLZdjEKViP+nCZrV5S1h3GXpShhZTzQ8Jo/7SKxDqNsJe9n6Dos9
a6lqKMjgLYqUCW+rXKY5fDAIqMlBC1ojWdVo3Z0h8I/meJLPYEX0PO2uupiY/4/H
TbD9I3WF/oZ8Oqy4d2YTmqa5+xc4f9ZRp8DUB6eLsaYWLcrD3kM+S4CI6biG8E8W
N42vWGJct9rYFnJ/mg7rPtYLJPROJ9bsTPJgXTEVa7LU0MvFFhcO+R5QdWmstQe8
qLPM2EsOuQZHNfWhRxL054i5jWVw2XvFgVtDSVLsqYB/K/ZQN0rMkhXIJYg/TStd
MPh7iKYBuQXs9Ejqk0eDxXQxvZ0kwt5DYCgVbDZzubShdlXH09nfD2WkvUO+xkOx
iJlEsT87p5RQXsueiHg2GoujO+NWIIY4ZFEsVYPn2XtNS+EDqJ6A63UlTDcrCRyM
YETo0MG4HrGK/TMTCbEOpQkdAKHvUXfI0wg2nY1AvNlO7c3s/wZ4wbMJlCvoX6PS
X4w+Jz0tBwSBwUjoVHnBijE/i1D9lMHo0nw2v3wt64xiVipwfhDKU8cfEvIbaKwM
dfkeX4fMpbn3TsknPZVzZ+izkiFdPVZtV8jGWssBaJAOpm2Wf25U23jijWZIBljR
GQVD90dHH7UkaK96wJJoSfKOus5xK9tu8hSwpl/sMADva27DypX46XNU3s6TYzqr
Tv2uZTlHKTQKAkeuRE6rrstuG29N3HuWt9NiPD9uVUZZTSWQmrxCvFvpDo6+CsSP
cWENrkrL2Zz8RCiLGGsN2JcFwDN4fAyRDxX/Ud8JmsdBwLKDE6lDSqFTBSTdk+z2
jCqtTC8dhzF8TZEfV0Jh6yBEEASgcyFq2FZ4BHw6hj2PURgvOkinaIkRZYBAWjHF
HWepgPeKNBR5IppcrLmO/Qv0Av/5QWvjO4IWcHVwYWqlfQNzBoF2ybfP8Rao+XAp
p7SErI+8+5ExiK68OqIexognWPV0H9YHmyc9zSHR4TCrTnJk7seF2V3O+ztTZrjN
CAeiZ/DLBFcnL6krHY2i4+eOlxahbx0F+zDUWLW1CZIvz/UAzGyUq54xSwhn/AvK
U1FfFHiVC9/0RPvm8ROVV5l0bfExnBsE9gbPJp/18tA/TkTsU9gIetQy3m3GzpDq
73XETs+koAO+JGf0pTykEPuWm00fRDHT7sC56gSsWIbx009u2tYMiV1xpASDLboS
KtfigpUuBkyVLev5De3YkhVkri4gc7ENOdeBRqjxSjlokmy1bHZ7Mc3Slq1qgHxW
yLW3EhAdZw1JmVSsnJGiB18pHqEFq4bsk733Mwf0f18R/NuylAWuqKeLMdFMSA3Q
bckgq+472853aPAQ+Rf0vK76FRfCBpp+3AkTYY2/f/+ZJvLhIOTWHXAQEcn3hI3T
39D3lx232xwffkDe9N+sZd6Z3jnMlYPqH8yb692bgDe1qdpeVTjaVv+jegnDxqOJ
2pztVTOguO9Z/VHVRSuH13a2X3JuGma048G6wtCNdXWY3tub4Gg9u0x/i3wg02xO
kYP+o/+Ilmw94nI5YoWEFe2M2O2ODzpQuoGRGXTYPasAX9zxEUQj+zX4hjNKJqDX
0F6A8h/cu3mdlvS4R0Nrv/y/GGYR3HQhe/gOEONDWndQAXv8cb/EULv2mkA9zxcb
5H9uK8WDWpTT+nhI5xSNOL6Twc3Mg1ZBkgvPJyK1JbT5RYz1TSPY88tsrc70k/vs
uBHW1NaMZ8owPqw+P7PYwzuFYxDAmcV0GcMTlbZWevlXhx7Nk9PkX5ivMX53gLDa
JhxfYswl72O24AGLjP03Z1QJvnX3SjJEvXgRn0nWT5SuaOE5rlrS2GAHIlO7bYnl
2BrsvoJZtEZS9hzL98e32xFU9wKs6TZIxXYsntWBEqFqC5Kd5EsIk5NNXEDcw0F6
dmvzUregFSHe5ikepwNP8KeZWdY/HVM+Nu/xaWqn9gUDNUKgRPKp1M1eLZSyAJrs
DuDycbF2r1ZwUasLNWeCDt1bYkigTCQy731Rqc8d+7dOFvqxPGzK06+eH5/0Eq/+
YNnfARuM3cvQ5ljiK6EtZjDSvvR/BLbLBnluonnvgUVH09UdTGX6rnlyit/yRYI2
4Re5JQ7mAWUpn7qKLZ3jkUl7We7ruN4dUCeXuvc8jjB5Nnpf6F7J/USh8j6scpmC
6v+HuNnla0JqrxBrcK7ZjrsJY6/9LrEU2q/3JaL15PbT3OjeSFNnbTb5EkBOiQTi
cH8NIKN66enp9wTSvY/A9euGHeJxOYZAVADaG94BRxlyNHfTUWia69aNzJ/3LND3
z/k6D5C8URdjRDSFI6hrrwlE2usLB1WfeKg2I/O2VGIm6TlOiLdySeeSljl+tcDP
+g3I2u7dR0Ib2c4zr0wz9ZU3cJu3y4MuXy4OWPLd3VSR90MpXgXqmwc46xK6JC1x
8AHvHFqZuEEAKW28G2f+QEZ+SJ+KWzCVW1rSLDGTEWgaagwICb5ohNGRG/BWJAwH
0g4SdQZecSCVEoMem8ElO7Bn6iwZgnIzLhjpvrUfAc98t+15nmynNjREhkZf+k+w
IxfnV8pYeK453rCqF0hjlAomB2SgGff0b0PqF6zZ5PShF6pXu7brOFJYi+bABrlC
8vSdiNeXHb2dZuL/3ILK6o+ViZdok6eeH0chc9D2y54h1WxuqGQOR+PnEAIbBCqb
c+0PBfNaY/+gtBRlpHvDKSq2u+/NJ1pRuZPTxm2uOmZuCBZ3DZkbb2pJszzLQfHT
nQ/8cDN5/+sGiKRz0Ojn03ZlwdpsvgRMvXBNrp1MvWoas2GDNSSufBKPMpJ3Bz5K
M5jw/dH4LHhnt0G4uAwpaPsfkWWZIo09DstvckkUTnNEqal0y4bK7IfCsGwvcQGJ
T4g+nQONLbgLAuDZI5i+L9fG7I9jpJTuRQvUugiCSRVJeDP9AuWJUgqjiFxBTI+3
NCUvArnT64G98whnXZI3ApzwufHsHQDg+02kpXjC8h/SMp9oLmR8KFeE42p02j3z
nfgnOOiHy1EilrQV3PmXgrpYWbphVtpCLHNfjHGXDUbZLzavPicjt9sMGigoeXNV
W1xuY+ZvNcYkjAjMdoykXYLsGcB/BfnP119AgydRyzTcvdnUPeCpM3kO3VRJuE/X
/F9E2g+qci6g6lDrENnbdjUdR9MtWJ9o9zdFjcFPc+6ZNwDvkoch9grzbsZxORmH
uA96nzeJyrs1dIiUErYd69Ns5IMrZJ4haZmoNv6/03PX4AYtfsRNLQcLveucGTq/
CtIysKOgj/0SWU4OLmZFDttU8rmJ2pKjjaCpw23KWfEOXYjyQQ1WayiX1Bk1hhSo
tAy71xlDW1vyZPBoZryffQ0H5/FTiczL55R9o6FWOVIQIndWzSumgwEYwhYHp5tH
k36LAwJF5o35K2eVzHQa5RRZkaOkEHGVpeNq9cJ3tmRL5ogUM9Ph6KeHZ6ndhol/
/w9j/YmsTDDUwKiWw7LJDNqoyzWLTgt2f6KTVUTkfjUqOXUS5NKmqu2V5CQsGIqL
1VtGG1bjCzu2hs4Uyye+ZV7Klpjvh+68FiOYYeitTdTs9gjl/IsG/JKxDtSQtBnl
eXArCEAAqy+iX87AWtDUySevX1Y88uuPP6vC3pcjqGfIVpOOOVSB4hMo49gN6pf3
cXJGZnZoi6xjaoiByte/w1oJP1iX/pdm0zuiz6AhWsvsz387csX6EGrc2F0fjqvH
q+52KLFSzaRBlo7H/aL7mQl56a6C4pC6HRK3jWsVNIMi4oOeAi/uSLTUK8+OPgaP
miB3uScGko0RhulFI/34+eVO/su8/qQUZNoaPdv9/cHDuox70yenZ2iByCmXHIw8
tAgDI2otgThgO0TgneBCiYvMY03LLuJ6ob2z4C6Hf1hfgyrJbNi0Y3AxyiZTsjnR
FkyrR2K4f/md1AZxDLcSbbKnrhCb0CdtEs4QRNoKcULK+cgTSFBiIfGjDJ+mxy9A
tuka95nvxzN1OsS4X2kjnH8EbYrS+Zu+mrN6mHXnByrkn0dCdW4sX2hNgBY5/Bzy
QnqW6v230V8zFV2pEPYNvnO/JiLIcc3EP7ZBZOi+k9+9EL3K7QjBOldh3XEekdeh
NTrXqrX+9OUEIxHvAdQxB9OcwVErxJLPbbG25VhlIyIIaKWqjGJu7hmXYn7pDHcA
yKm3sPJuVZKWC/RPVCxb7WZ+rJzZ9JBfl7KMFJXyb6fZem6sriCgZDN597z0Of/f
pw/27sOYylqD1BozTQVm17/XRhVEF3z9vg7JKDigBE4wxDIt7ftKS7wu78JoM/4Q
hCZ7Cod4HgapuToDyoGJZe4ubPUP2aSbBBdMC2mfz19hKdPO6eCDQD8x1+cX//qK
XEzQwgonI+JFyQy9BgciLGJgPrZtFCYYVhVyba+WXxU9Y7ojw77XSP8hCtYs3/68
s6DJM8wsXaXk8en6YLMOiUH2y6QFCDt+9MgdbqEi7wu2J0/W285JA6yXZbU6MXLf
P+BNhn1WFObx1pBlFdsx8FxhQL783TPIkVq25ywbIyMPHyEq2Jy9j2e/i2UceMqK
gVsympaw2HXoy3XYRO3h6GORggoEn5X40vWPbzpyZTEp66HNG/yEYyjTLiNEOrZo
R/axyrX1ARh9/PyVF+xwe93Dr2ZEfjJq5rWNF7qzrRpQ38p55yfjJ40tbVeNiyhS
bYj11Wy3/issgr4SeHxqX4xfwtvxKGO1tO1Ek7NaXzbjo5aGlvj+x69o/3mR2RqX
neu/3GPSkc/bw/si5idwi1uNrq67hp1Lz0oA0f92hJJ7zBH0Y6R8/87JK1AsoaXJ
ZlYvwwE/XYRRW57YAHQRZrMqIlIuSh2wiV1Wgzj+YeZ9+TSj1gBt9jFg0UdBhrIg
FWMOM8XqhL9xpX2doicVg56oA9oz0k964SLKRW4igJ6teiUQ1MWqq22F2y9QHpfM
wIe1TMuRv9dZ/4FE2vhpqPwMpgfsGt0pjw+c1ZEw2ZfmFhwB8bC0H38ma1GSbhBs
jgIkHzooFRkiFXiWLorLEbcnzWU7ZY9mr7aHdJ2SI5tRXBZ7dJSWi6DKeNbJ+Pf9
1sWJB4ZCynZEjTYIfi7iORRx4vs8MrMUfbGyTIqDPcrLUWEeBu/ksHQgeV2y8oeM
lQaI/4VrPCNDypt/5y2MSJgOTOGW3lEg5l/z1QnXvy9LVq9QuZeCR5Z7vPwobXwL
7R1pwB/FZiuh+jGXytBpE8VdCnZQizuVbLQmSCzzBGLc3lM7RXTO4pBa4Kjgedh5
S4Zede55grx74XxB+AebdQVyD+SZhcOyKmrfjFUFuD3WRRTsg3H5uWUevlxFpk/1
mfHB9b/dlNfBQfnBRqyI1d68pi10uOlwK8QqPpHZ/p5YgMMda5TandG1UkfAQpXh
Pm1VzaYjewtUcCgyBfkNVwCdJVlmsp9miBF6pbZj/Xpl2D9ffBKl5aSCksr/4Lwv
p/+oPLgstNBb53fm5IT4a/br7ghQX2AegWPQUNDecn6lEf2zkSjW5sLmERkBeI6K
soJn+/c86ChQeQiVxhofT9frhcKwUyvBVaoBGkrWrfg/TThLzxevuVVPj5cR6/p0
wE97avWwG8y3jtDXntNTMsDmcubBeBp2UiWb/0E9ckdUtrGdZ5SxbBmcfHpXZ1xm
28CL1IRw/TkjTmnwxMGigbHgvEAzQQbu4ndOyZNlxTPtaHHW1tDjgiM1YufYDtQD
sg5yHOsRHdnd9Y2dt0dhTe5cVhKSkcGZ4NfTd7uyfpMzlNkZ9yiu7SATyOLwrRmB
kkDwq7kkIAvV8C8lM82vP/N6adO/Kc/C3zV+jI3nUj46RfVxM7Lu6nbkAVFoyzmM
Bg/7RgxOlsR7Rlam45PMWjS9Vh4PLEGYuQRp60X7DFFhcKXv2vVUezcalPfQK98p
qRqfBBh7VWFI7XVMxzdtzXi8OxDQ2evLrSrnFjjZaPSlScOprz6b1qq0l0Yucrs6
22TYaXjpYD11qTln+/OZBt3oQpbZMIoIDAqAZutWvaSrYgI2GPJ0MgIJmZ/llsZ0
In/iKIkkIgfGMQNohKAN5Z75RcYkEmzsF27GHzN9xPNfUFppXf6dbD9uEenoEriK
ePd9WzJZYk7uYLvEqPg/+ltU/UjvlhxQCsYDezBElrIMcjGfb8kXNo4d80mLXtG4
6uCW1a321VwYC4Z/Qd9PDrrAaFlgswKwfqYHcVbZZ8vnMurNh9P2Y//IcPh7qK7e
bb52iubNFmg1Efz6qimWsSemdD3U8X3AgwDSRZkN8ZaOJpxKNCBJsfzcJLVPUP8q
ETYmbG5fpRRqMxyKm+IQQwef7EmgKNaU7dtp50DkND0+JRvi3wi18nwPhKNdZO/C
UOvlzLe40+WeklX9nxxRvmiEq4FNg5lLGWCcgW+menSFcJjHPfSJNvfn8FxC0ax1
/QqLKftcnEiMTWRF/PXMYycWZ5T6W5AqtDQscSLNo4s1PixodRp8KcLcpEX0oPE5
mcA5PhHZ3RgG0t/vmYTFTQ00sZ6Kb5pISvU+tV2MqwD50uAAg+oV/RjwZswbiqsm
gp432NEDSb01o16SZr6P9iHW5fJ2JXd2QpLRMKrKgmJnpNcfkNY2G4iVk5+rM3jE
va721vuutcEZPWuLG5w1LPWe7iSiEu9ZJPFHITcXouhEbXM2N9fjfGKWVMEwcDdU
NiDl69xL9XT3Q4cLanJblyo1hYteWWuGq3ytOPctY6w5G2ZyWJvXZqjTdmh7OUr2
1O/jTRzJIniHQ66UuvqgwQUft7aSKrlYtQ4CztMxjSTbrl8xJxJSn379h8EdXIr6
SRSFAXPCEx88IkW9rJrjoOz4wg8qkfBpwc4FJ6M4MOShj5Ws/t62w5fH1Z0LInwh
w9z6w2owUBzFEcDeg/IAQTpgNb7Ify5TdIhPC40tk0J0vSL9Q57Hq880FilIyJyb
1GLdZ0l9dmX0KerrMQkveUPWg5eduFEWIXhOyLCRdaI5EvpbZTjoEd1Mv0SJTL6g
w2u4sa/QTPg6Z8uVyrBcMn9Vns+TIe8MtcQM3lVVl4iKGiCgFzgwPq20asGBQweY
hbWBz3G6LH0JD+gSe69XvUSZrY4Gc1QUcw0qPblZWeOI+CzMZd7t7tde4VEZrnad
WjxfbG60Sj5P00ZoszNotnSUlsQF7N2N1XhgEHGtEtnmj+JiJoYCY/hpAAhlPFLV
NC9cq8ToW5QcRV8sxDhVoXlBdifMlfSmYlGNg+4lx5DhhJLXvJouB1W107snS1gx
idKEe3CI04Gmhd8xpxQ3A+3LTEIlW2k/DpSkl/ZYtIEmBm6XJuxQF8cYpjDdykzt
D6LRne+SHW292gMjGcHeXzx5f1OEzLVpU0mBCa0hRbc1GVXBrrqwSPMo3NWslZlA
RSoF6yz9Sz50cz4g3O7bCDV7DHOa3KjZy2dynKskQ3ssmMqXgEy8Pf9+EapfYixT
3R88+UhB6xKsLo/vFCuL1grk2tvbp90Hjb+F09oMxaScopHyhqveN6x6mfjS13NT
slNJ2t4lHmkEi+yFUUG1luMbtu5LkTDU8PtvqSoZJxbc2JWmqnkktkJD2TvkSW7z
fssyc/0iZpNjBa0ZF+tK2a+kYeMalBcPMHNHFvqYh/SGNf6aU4xodStSjXxaz0Bv
a/2mXdThcWnhy6BXQSkcNES7i/Vx0hogS/pqownR09nC/59oYfwefISghQJl1lPt
IqFuIghwu5ZmglzUlK0iFNEEmZ2IjauyB/e7osZZHYPFNydjl28anMkxPin5qyI+
/IPyhRXSIwzS9tWxu5wWMaKj3FVp0oXw3FMACIZOxQURBhW7xRK7hQx9UHvRkBIv
qFtB57mQMB2UiZWYsdVN7mblMv3+8FBttQVucL1NS6+J5xdYbNG5bkDRoji+09lk
oZhhax2K3I0TGO6o1Q1rP1Yu0v9tWaQX1NnOxhLTQU0f0iy/BVRivMFOOLQL9a9C
T68xgq0EkwMswlB8HEde7DW+SGdM9RWVVtFOXymQ8c+2Rh1EUGxLkIz1CGjLLKq8
bvyTSIk+f4b76eySUwed579ZS3yS+rlWx73NaDpw1jTRUuD6Z0N2X4pj3UuXruFk
iqp8sNM3xpwO+RwqL3gQrSDk/f83boQ8VGPLhSvP6jddurDyXA/9Jz5uD2qc63y8
FsgEFyFu8h2uF51O3XQmPcs3ekxF6fnDoYlpXeGVo/xl9lFB1cxwllpgWw2hoRyk
ivKPjvxOmssiKDMUAJJsgn8b4k4zvI49K427K1SkoyMhugdOe9vbsRoq5OMjEkFp
KjXnYEW5obGnyvMiFEwuqaf9TjuuXIQR1cxOHojblir4JCFcgcfQBJksXiwL0l1r
63cXCciDI/UBQI0RlP50lk9V9MDt1Z5PlhIbBcpgv8ADo6jZEou7o69SIqjN0K/B
DL3dn+O/GHIO+gRywsog0bvQOu2u8S4C7rr2LnA7PDUeBf4QWi/0burO4QogVIu3
Sp8ftnrTPaqngBhUgAGAnXz7LDerDUHQ6WoxVcoxHpv+QcLtuiONTPx3ybS4dbEs
2NHwo78ADzY80TYYl2X8w/JxRkhTV3Pdr3HvLbERucQ5RstGXDN2cGKF5p1VTn29
AjryO8eC3mcvdF4g5pS+dk8cIm787KpCiWrCJWWX2aBrIJ34HVGWD1QjW6y/W2K1
EzgGZSyDGOjZsvz6+zRiA6QOIE0MqTbHeoAS4zMqarhy7WnckFQ2KiXCUEKBOh0e
Uuu/wKd3tgTGBfqDzsc2UqVcr/owoH3M0ZP0Vcr78aJNyIMbdCszuT6uRCj5dJrc
yGNlm8zI2jEiOH3VRhZo4pZuO/FSGhrieLH9dobLB2Ppikt/IX8z5kueroHF3Al9
4fQG1vtA1JBdnp9EBG4Trt4TOZb1wbqKsuxyOQX0SVr+GNwQ/nCNExx9s0tF7pNr
h+7OI9ZZZvaVrmKelhSaniT+vg4VLEu4u3wdHw6pZNf1Il2IrnEzXMKPoRw4Q5e2
5k/NKiDw/StDaPEOCIL8HihEEoQdnINX2bf8jpRhGNbZ5ChabY6P+6h5zGYSgjjF
9A3wm9aR/0Pz3yUMNfJfMzWwjYY51/sJ5Srky3hW5snu4lsfpdMlSL+hVjBlmfKv
dlPUM+CSOem05aulseZeyn+xEkVWCiwsoMnFk6uJXS1dtmXNqssifibBjhaqnvja
nDZYMdVPkDafMcyq7P1KpYGUD4D6fYToxw0jQxiEX5TOatHxgfgi7MCIz9trmDnz
YmhC18+E2uLIRkTbChOowbWTr4VoI3h4bsaLy4IS88JjVm+93WsetKYTxwmBjZzR
mwFhEba7cBduj+4QjgdKVGK49NAVojRHf1YFJ9bxrBv53cWgdY5dFf41zEpC7un8
sVIaaJYIxSe2maIsn544xmvkN5JFOjxxNV0PTaZreAJTCvnoG7ZXTqw0lInCJXF+
Kye+gyYjDHFDwJoGQtaOa9TrRdpd43umFZBq29YC/wr/6fpr+jpIoG1ZL4Ca6L5q
Sm9vV5AVPKwM1h5T6tATPEKssd+bdj4Aht/0BNBpozOQZxtqIergIVMdPG+rCzlh
JgF6c4L+wapU9AmRqjEGayb97y/6ylcYGYqG9nJ7qqTEf0a49d8ZvRlCLOWMLjXH
QJWen+oDmqK0YDLTi0bw5DJVpowR1FIX9EePqJD2y6KBvBp3jVU2ZCTBjGnk1TzF
B8jzPXt2RBNvYRExMPeNInCWi65RTkKWplVN5Ps9M4ZES6wbofXP90xs8GVy7QZ+
ZFgxWejpEnt63ovaew9EhjN5rvqk7o3wqhZUzuiCNldVCtSapHWvcA0/jsb+RiQN
+CUxchZXGWJF/Us8ykzq1IpoSGz8pdPxElMYDu+6nED5zMIou4U/dEdEZVJV3GNN
nMvUTMK/f/guWxztjGHVkiUUq1FfWXfRM9ga1khjo6FkVx9REBP8JN0MzxTvDaCi
PVNXSeCnyoJILUx4VrZ3lqnJi+WF8c71BDJZKRb+lwghz8MH6xM8DA2zERwj2KuY
LL5g5gjW45EUZJVlgWw7yDWYlM7M+NS5rwsSCqaZ0bP533kgUodgLxz6dIuNPFN9
wD57dhVX8vLNN6MH4lBUn/elF3UfK9+FUuougR1n/KE8n7hvMB6GDKY7/Z+pIo8O
icbPuYsH6VThsZqP7m2wMqMqKgne22PaofBjNyhFSfZTXT9ZlZFPfFvz+YgfeD4T
vURy8BF9B3dWEaeomxi3KUoQUhJ0gRyNiCao8+DpPuWU4+glJfhza2yUyHcKlIlB
aoIV4TMHl3K+UqvE5EkV6wsFfHcpPucyLmM3fMtggamTXSSITwOJzpvD64j6FZ7J
yF8l5pMe6MrZ8gf7OFHCRsupOuj7VJl0G6J7IqeolzDMHsVN8iX9FzPRf/moIRsF
GbacjnhNTMrPxq+PxqyWb97mMooGcbp5TU6AYD7vWwhpQcNSFqRyf9rEGoYym5Zu
ISE0ZRYZTPtUHJoVEoNi4qbkXMRdRZAeAYgco9sg2V9IUT2KbOkQ1l9td0Cd+k93
kAJGlx3ThuffYQDJp4zxFK3qrw3Leo5MGp/kds2QSguqD+iyOKoja+dMaL34h5SE
GWklGyV62bp/co+MeUig2MRB2v+1Nq+FIdq/IUVoJ1hjkhgy5Pun1uZf8nTjL5Bq
sxGxvQ0penBYqXrmMfzZOLjbtkW68ORxw1hvDN9AhaNgb885bgBIy4khiMbOjCUb
KPbVfM2OEiYqEZFrAJ+0LvN5t7i5yEXzrP+Afe0UFOrmTV+dWdKma5QELng04mRW
ihSGURhAlcuu5b0aDPJZ1vaxgwG9o2i+vji+nfTcr0NskULn+Vt5k5EAMnP/PX6R
wYS0PBz9DG0VQ/q/kj5Njbm1iY6HGFonA04wCK3aSI7zYiI3D5XbkYnfnCWOE8IX
uKRGJmLBPGah79N+xONRZ5ajmyVP0C1Pv4vNxzq4Z6BMq6iEIDTem34JHhgQmXTB
Cs3tV03UTeUdpFvsIuyNOCkfgdKVmSB4PhTpHDc+GWodruHCsN0lEGn+JXKXpVaS
rvyeq820AMga7AolvuJEBurtLV9up4RjP0TKr4AsjQbcQmqMtVejvaOZU7KMkbbd
GH287CXubgqNCHM/BMW5IaX95SWSBBh73bwrw+Rjbs1DjWWSPvWLA7IEyT8ICcM/
/uhjhywI4ieHdftwi2txwK9bF/n0QltB/8H/rN5oHH7UV6lXEjoHwEWvstAoysDu
O+Eodx6vAixDYp9S8c47qe6DJs0rK0eBB17w1zi0rGpSaVDUia6LBribxbbfLHys
fY0ltgDxXujrK5q+NKoREh0lqoWzrTqnO5Ttrr3plqUBfkd7BvRFv4UF1mUf0mIR
Jo4Xcma5OXrvW+gk0sPmVWxGjD01qdT6KefUsIARe9SIuet3HyRQtAoMcMvJgV60
eXSd/6ibt6OrcuhlgYKMRdqRAB6IVg7GpO0s0sfJnlL4TNU1ROkIq/3NsmhuevX2
9CsI2w5NJXqds3sW0F5BgClU303r8i1A6pqdNT3lF9MyOm7H4Xw2xsZNRbO/fayI
HGyW/i1yrHfgD5HecQ+PKmjF5wnh2Gm7i9Ex0yEzCP4nqUl17wnqsOUSh32G5T+p
iItQJpzeUE6enlIVzMQX0tpBPLVKkabTopQYAF+guSM2dtOd3pC0zLnuwTaYVGJt
7/xUiYGbiKDzpp/gp8iB47ucI72p1GOzp8OMdd11WTFV1CEna8FNZfEILaBkZ5Os
dRVqiboxLcyNLZPeZjl0tFmYxr7QkqANhYKAjpKprgyVMn20DQ4RjHPbPMlD9Ah7
mV6ywCkMqB3VZ4OPq8+PmDGx7TVz8XXbche2ckVmTwnaqr768kjeXhGio4SbTDMW
YcFfmU4JZegll4CUP+qdFEQD3wSdmINZfiL0mJomF1ZeMSTBvsm+9/P0/g1VJbUO
P2/5JNXl4HyzUjBvW/RB4xkq8MqOIUWR3vKydpvm0HKVDV4l5i0N6AEB2fgCqq17
DF7MkJ5fYNIpj5EKe3XPxNixK9bHp0tkkGwGjQ8J20oG0aOtxWP3InIIYDRKf1Pz
e8E33uXjRK11GaaFkvL058PYVgfjppBoZKUquM7eiEvbG/Vlhi+vzSanZu04/HWZ
TXAQHNaelHWrK+546bNiknZkyORr99Tl3eiYaAvUeyaLhKaD//3xrzaiUXg/A4G9
0pgrQuZYwbZlIJ1tGZ2La8Xsi6BeDHTJhakClP/mF8onNpap0NJFMVu08cz7OZG2
zOcPN96wE+4qK5RiN+Ase5hDo0g/ZJzpHakP1re5pJmvBjqfu+NATJLuGFv2Mvlg
lOsIfiGH/B7vzCoDQaKYaT7vPfUtjels9i7kxUMzR+aAduFZ3xltPVNJ0EIwQHED
s/uc7K7sHFy80RiJ/BvHjBJW3H3XtugdWxTEunlwQ0r7EizFVa6ZrIXnAHxmb9P7
FmdaVZ7xtXXNhLGAWVWnGCyvCakieLQ5vhrqsh00HCeYalZbs2heGyAq4Vl6eanv
xYFUICHOcRZ+htT2LmGg8n3GPjo13prORxzhvO8ekcHCZgGrd+FiHf0j9oDOEcEv
iwf7G0UPmrknsbse3unjg288qEpLGt4sdnaY0YLkcbhjZPAzfdYhXwbIPCogPQ+7
WmBucJjmPKdnRN2+l5kLVdGizBKM6/7Sm/r2mB+fAxzjz99bmTlEuajMo0WSGioL
asMs4vLlztFc5p7N6YTuUUDiyRAZ7UYfCsTwTxC9QhMLxgxtQkLP0h/2JqzQB3n8
lahdwFOmKMEWkNLM4eM3Jvs4wA7X1GwPdNKPw3i4aIeYgg3tHNTGLVDeaeZUQrED
lrurUACDwg+12xPLP6vCHLwf8+9WhCmjWTQu9RV28MIcBr5dDxTMWkOFuxFO+MfH
e/JFNrfFe6zrqVt/gaAY/aDKxRpfk4doKpzyo2BqpcbG9hv7gy5epJ6fPEHc/Gcu
VLuO16WAhz6R3vQthY+gXdnMMsnzlW5NDpQjPtsOdzn5CnTeXwcIiygvwDjx9GSH
N9lEeekjrrVVgn8jwFB/ILjrzvmxTbTXdalEJfoPm4O5yDKDZ49WSSlj6HZJ4pYr
11ppPmZTpsgCGIevpW+g7+wGMietbQ1S7kqB1SlXGc7/g2mhs7SFUNfiHaHO8HtX
MJYQk2rhWUhBr4PCxjtk8t7thoj0n5TovsDvcUWtecbqtziFP8SwfTgzuolxo2r6
0TRoOYkkvafN7yiar+zKeau497ZXCQP12dms6UN7xnIx3f3MMtmvtltrd3DU5AWB
YwMawOP6y2IpbCHDqDQxj+90ERhiO+D4bXK75HZlHIafXUoD/MUVHL6jUnVsWpQ7
vzbhHF9HYUQ0Nd5qs7wvlK4YfnMhj885d93YQxvzbf0z9VDGSFXIXtQoloOh1LzR
RV3hROMYcO7LPoQGbkKXW8sWbMQ6ZO77xzMvLetOBEqwsYoLHbvI0zstM8iYFip5
dA7RVgg+BEYdw4wN9qmwPonIrjJQgTBJVlsukfQQ8gspQ+fLvUgXQ62lZezvB8lk
zkPb+7xcT+KFPOi3Gyppx6gZm6bTmM/cfJSVIJ6IW0vkn88GQrrOna1ilolflOzQ
2QPqf9NgY3jz8TaEqhkJwuUkizNXm/CtrHsRNa6qV2iPgY9vymBSjXTTIdDeUwBd
gc5TIvwtbD6wPIrWZSw2KNpXdUIz0oTzmYbR5xmsUVewaiknXYmtgum36/hAT082
hTCWO3qH6Z0hiXnaNcKSVVWMPknIrlFGOz85GKIdHbTuyaNtjCVgz0YS1na0FOsc
fv3G4gF2oMJaElALH1IdYfDkT04xuBbx2yTPUocxnL3bgMnr4tDs5QpzSitXjKHf
cWWwl67j7UrULa9F4WDQ2ORPPr+sNn68ZdPSHRQG9LC6aNPi9+/D8INgo1mJNqaN
8tcKa5Y4ensDwzvex9YL/3jGEJ2heLCeg2BYWzZySdJTyY7LaV2wedbLX+M1detX
KKhtNLun7saIZBgtsI16ORP3PyeI0LlQJ37p7KZn0PJVMZA4HpKlJ16s+lZHt+Fu
JJzGOK+q9VH97fW6kWSRlvzRNpWBhSej9iWDk+lV5k2S90VxKlGdEGkAn9qAdSHR
18Y94kdvzcgNv/To2Fzawk9oJtsrYr/lNdOI4EnE9dwap04iHw07V/rvrE+D+5yP
LZWTpdQEAkjDH1P33o1TUxKAPrcVjtN40Gt3FTdCJiXKU2qmGUvHIswPQ+yM0kzn
m7dEDNemcimilOdeL+/BmbBDuify+Ksu/t8Nu5Bry+NFul9vd7IYcE14u2fdBMJB
qAgM7/lI5VcLxY6kPyBqr+YLGAc/s6tGLVnH3KwFxW1N5ECfr0RmFKNxbk1qo9FJ
WQ0IWiQJkM4JuDAy1syiCnacB55xnEHcwBsZ1vIzyF6MVuAs7laOSrUHPID2TdJr
KeTvap3g9zeYl0rKSe7LiKenK5C5t5YexypLuiNX6+YvIe8tpvgtvQb8DVTSJ+ji
NYee2v57J7qAtGNYjdrMzWlY4yy/DzTQbOgM214zdlUtkDB8KRqzi60pMvB1EWob
lVPsQMvOBF3FpzTHaMe0DgXJU/1tA2RU/PZh06FyOBvoZrbGEG4cFOS9p9HDC5Cj
dlY+k/ja3VwbWBt84cS4K/pwLeq+hqYTLT7Rhdx8fv1rSoL/QwzD1UwrZNRHiTyM
c9p9dRZoIxg2ZD5rK6+69uia2tvVVefGpnHv1vDyb4kkny/StpWv20jhiOgVPLwt
8WGtAQQ9BBlNmDsq9HUwE5C7rTzIRg3GA22eCWjZWJSqU+i5UHT/059gSxK15Bwi
eQXwI6GDUHr1pXyvXA8sSa/cFDO4j5Hg+Z+kGNd9473QR6BNbaodsZUvmC1EXhnf
IcntQ16ZOM2oEri19e5vy7+YVgtF3XZfwMtHQ8t2Y7diFnKrF9Os6kR6DPj5HcOR
aBmqI2M5DcfNui0L5Iy072WrdCILwh3OsKoyT729r+nWaswliP2qBy7bpI9hKEQx
EG+Xe08HBxJIHmLUrAaK7NWd8qQU1ntVxlfPXtaj3Jd8/P5SMvAYfJBDgj87RY/n
ZiNimPEZCjD4PtIO1V3VDvlnPgN+aHKs7P/MwsLLQQJ/RbY657oIcvOdh920RniV
5HzKqDOdW/pIMw5WAeBZmEFKsuD6WYdyDSwka9UkZjNJ15P1k+R/wc07/OCf3i7Y
CPsDkTdjNY+nYdztZ/yt4uFFnIOEiP56Fn8sXpe2x5d+vQa6SipesQmWjOzJaIje
YL7BMoxcC+Hcx1DhvzgTmVVXXIpRwiihv7swp7iE38kdA0w2XU/5sUkauaJi8lZ3
AL3xXm7haDhZlklt7cKcHHBo/L1T5ENGRee7kJr13eNu6Ojb5akZhhpKb7BREAhp
A9W+hOwgwr9R4Z3QAEX0AOF0b9V6bXsK4VKmP1jfzN2FErshUHSxm5+aNyccvYIs
CiVaE5u0zw02MPwNVjvXll46NLkPXZXjFhF5nLSGdnPgfON5g0cLJN7ARLaJ1/tc
peU8ADWO81ydqz+jetkoKsz0Xx4nTB4QvDt0Nw1i7lxjzh5FQiV6MKLrwouV1WEZ
wm8KNAFAw9I41+oYuJUwFSJ6aRKtpFFxlQc2qsN6Y2XDvX4HLu5mbN03BofZnTzy
D7k3Je3jUe9Dr7hnCd8ZZ8nzSiP4hAYxsqg7F/k0L/uIt1aW3GwPHyBfxbo2guEW
mhJmnWeG+0X5Vpbrql/2c2lEi9pNQZG5jHT083WLLVpUD46sGYhpAGCE1s4/f3LA
mDNY/QDn0zNSiQzNf7135QG+AuRmDtiHbzqdaRGeaLnHQg73xDIOb0XHN6mhDx++
EkxrmfpamrofO/NRaHioNGv+wQhaogKvIzgBRltWmWmq9X+sXULfNsd5602fIvgU
mXd9lFX/KxCG8HXhYUSAC2K92ZVLj5qVn82idkocdofxHq+pxstflM0/p6jf8I+2
7opYUF+R2lZF0/Fy3CQhVypj9xBZztTaTASL6RD5WD29Uh13wZUrqCwqPQn5KcJT
yy1pKv56e7gohL4djxuzxZ5GQhG8jtVxN40XwaGqtV/ePM11fz9iTK61zYfCrjvY
6zoY6y7PKLN2lucRj4GJKLhTXmnLuLr+A75RcLK7bWmIJ1yerbWhpHI0J37f69jR
osFlxpTNIvvjlvIPKR4eHdVf0nCeTHXeQcntLM+Zxrnh8xZLpFRd2TOpGwYd5+80
CGaHTmBx4UbJd857JnadGp6PL/MzoTfrubT0txqAqmgIjkqaxDInqpqS2siD1ro/
UIP+ufW850Lv0qdhoXfLIjdXl+l7VaEjQL7x+FU4OCXiMCN/BTBvcH88lDEh6kTM
hyP8A537zSAWTHgvvvrNXMs8J1Ghvxvxp3M63hGnssrvZUBdckELuraaDGO9A7rW
AtWcM6zY7I+wZgNGC5kp5YxOXv7TJvHzwAQ6bBNBNEtGqGVyiAtXBXMksEULRLos
Lj3Ce30dAnIJZEULag2fVJVQBa3N1Ey5GLB6n1u/88e/dtQfDLsnn+NHNzzOTENT
/h2gYtNp9EAYKBFterKQPwKkNVzzt4nP4rzhD/xCveeJItOJKdX/+phqg4XM/AwS
qdn5qBOp0tU2fnk82GH10/0Vcvh1ujppq/deU9xcGa7YppMBuQ5H8eueG2MIYybI
xsVOeAQ62H1Sp1K5FwLir2/fc7k5EhauH7VhlKnQDLZ9Ck8OnNu0Pbn7z73RmObe
5u2INxVwBWRHhUYVhwR3JcLuOXdPuwOJwZzKk3zXY/SeGTy4ulrjoPmGnuPfgSiu
n69S25e+mRJEC4bGwCorOADJZhwHYvOdB8E7eFfDmVowl4gP4Zwkgq4M6DHY1CtB
XG9vkVORMPsql+RNXFaQuW8zfKSXSITwJgnFd93FvG2CbDPsXbKK20NFxoAtWirF
hDrdMy9gkmLnoNmj3aNlBm2zDYy76PYF5c5ryzFADvxDxDzuB3Iyti7qaxgf9A4z
dmfqzCG68RLS4sLFS7sEv2Vs+s0WwSd6at4cLWMPpQfeqU0Mvsh+KH7z+pVNbstc
SORnVO66WU1LSt0dXT67UCGCeqZtxDf6Z+jkJcOVlPNrodR6QNVIr8rhYPX+Myfo
rGQyYkQQFj74PzxTWd6Su6x9xNFJDyd/Ankqg80kE9RJOZIXZK9s81httF0o9ypc
DHlquLnjMhjqJUNKDhkAlvBw6MJKIHaABAsWB6K+UtA3Xzi266MkW5YhurNiO2gv
H4p4jr1wQ3Ly68RXyPILuUqt1l1a2bHBBxnnxFljc3ZGwtnHQT6AzCF1jHDgPAlL
5TBTSpYFmi0wn1GfQRxGC6rerJKs526XtJDOlDLSzwHiAmoWBtsn0bfhYzJ5S9S8
YjGmTDDFW3ooeFuZVCJAFRApXxyvyxyS4W+/1nkpm3jVQZW9YjKWhCQ3iDwJk8sk
7QHV+8+/zxbgrBLKi5bm62ffnRU0Kek0lVJ3n9GM6cPTwlsUvQ6PXiwCxfPjo1Va
Lf94sYOnZRAdWTztgoiNM7eH7vK118HGM3sIKpKpgaqNIvRqOFtd/BOBFjBq8CNa
LcJCx6u4yG+r8K+4+TD2AduXh182eKzaIK+L5/tpIBsoQ/I/9TJG/XXBJVWmW0jg
FvyGV2WP4cDDK8tQ8E3iNyv5a8U3lqH7S3xNhFy8DK4/m+KBd1UF+ZRWPF1o9ir5
lxYoX86VOtoSGoFa8rCz2VRrTUXIdk1vAlVFrlTrUbuy3K0mC2ra+ttTTw/kSeg+
zwKbRzT8/dAT3SZVwZeSq/85AY20sULlJ4hGd9doRCze4mhQk+AKRdugbG4rTw3z
zkmhELUGA42ettu/odtfxQ5aztg3mUSSaGKfKdAj7uKAYfVQSjkcmjbjEyigwyj8
5e+2p55GY1ZCsK9oSblwgfR6oUmF7fYrlLPUiBPXcwz7fmPi8YHkIg3Tor3yX1Hb
4IIVeZojT6oZJIiUoIJQzaWDqk5SSMw3wcFEPva4cYhWFAVZjEGgYrEStU967ucT
q4iFSXcstS1sjmMBORymoKvuEh4IZPjQsMvPRnhVqzsnQAdgjUrs62FqjCtZIu5H
RrivBvFmACwdZdgy1erHFF8njUb+9rCH9NhZZPQueg/CEUmdb9QX+/m75dk0PGSL
gJEly4AR0gvri+wuGUeLnVlMVvT77rHAekCOKw2bQv2mOXr86ssNZuwxtV+jGoZW
jXv5Qt0trVeo62iaS4yVgpqMxyZZiNhNAAIGTJlzkOkJdxnhcT+/0CDKLjhbGreh
91/j8h1GVd/471OwpLgEWVi7qNCojmrCNp/ldGP7RXbsuMJZrUYysRvrypxeQ66c
0fQRYQjEdi4EdREVWO4rW4Ds/luqLB04GfjWFu1glKxs26Mdg70qx3wWht5vYZxo
WYJSXinxo9XfkHJaQcbjiHi4pqKZRf6S321hB1yS3r6GMGIT4CaUoed6MD46oyso
AZF7uX3uFNbmRrFVwiTqdVJDIp+WSGZU1wFixWJj2vSO/9vkEpNbENLu4VbbctcQ
53cITqa7EOmkjKSsY2T0I11+w5IMKXnd0RbB2B1K3fi2uzVq/DOwjUUELhDjeN0M
karUDIqqmvt7/O+Chedsz9eJrbJl3LDx5T0HQfYKkef9Rh7sHkXDFousb6z8B8iU
6QoBv/M3FgUhF8ygoDpfIzyxzcxSBOB3K6trnw8u7yubrwVK+q/CU7eKTz0TqTft
AqFdmv1docgzBsIqBcLw+ulCvBhv0GGVldy/0BCdnIBXqZSBn4SWb/dpjHfjtgi1
tVw7ApOnXS7gmd4CtkdekX+3NlrccteAZI0aP99qAM3RHK+K1OJZSfuNTPDHY8pY
5kWfQ9PxCTTN8tcwQVfCRVUy4lCIqyNYj6pOKppIiOLy7se7axxv2UDu4z44YPnx
i2eJag3uXOtv4msAuW8Vfy2HXzqCpfj37kAFUbxnzm44mWuekDJFPgpYfrIT/NJq
1o5FL28qA4ypU8mf2YdgokEwXBwsdHIkq8AI1sghKIlNYItGim+j1hm82cRumZ2p
qKbNqgyEw7xyH4RM8j4OYfOFLKPl8QV1JeRaRFKaphoinzRF7Lk6LPoUwrppf2Jc
oteyszq1+wvKYXjergyVUtEo+0kIIWlXyh/zbhFdraw9Xm4Wj+XjF56oz8JBr0iB
k0pulhCrdTRLEpyvTQI2ggTtVmCvqFetK9iHd9goHca7Ahv7BlplndqG9JZUwBs5
rS5lFT0fJW9xOREUKEqQbDZeMvAkjKyiGz4BA1UGQLVirsA3LY+SR4a9Hsmureo1
jHteLpnDp7XudaxxPQWBn0GXxI8pIPSNTUtrnoL2lL5xqEsDOuCPpx05ZhnNswY5
98TzXZ0hrWyrNWqBvfee395eGmIshDFT6owa8ShWjv2Z9CDJeR/UVlhMqtRNgMZB
1QA7L3FY2weDHiBNX2GUB7GeSQSw7RmsHmm7b11++k/EMSal3dN/homG45ZMCDxO
QXNP7vyccyYjwYR4USqtAkQYUcnTsOugLrpKnpO7J9gfEpD07RC25piFI3cc3aeK
/3Q7FA4pjMKxbm50OZT7qPtAcHP0pqobdMf03TNa+KeVTcDKdtRYcTGwzmrrNfC8
XDxavdAY7fXYN/rqAzaws3QjChkEoVjlj+TGGYkMKxldDsZcxbBZjN6pZqsFdanf
KKPmRvBT8uIwte82210iFmR8WFUv35+dCmQj723TZLFbwIs0wJQnE9XOYlfZwGnY
xbUocD1kK9DYDk+82XAOc2whukSBsyaMEcQvJOZrx0RqBz5x/in3Fx233ruFdn17
ctuwwkN8UGdGMytX1fP4JAik1xAuD39YeuGGVDCdGN2eIzvtD+omSygcWm+g2bfU
ASUPx2Uih6AP+jEomc1P9C99XUyfvspSNwVGBhqjTbXY4rLCOXLCl/hvCedFDmcZ
Ams+hjD8NsKq8SkZJRfxZz0lvINh0HWBrTggbHnDx6JdCq+gnpQdzcaubF5dUCvq
ZnpI64VfO+A5IyEbL1xNEKo1U6Urj3fceUdXGSxtVsf/JhzBWgsWmABODDM6BGtA
zs2dDOIiePeNEBRKv4+VE+yANXe4P+fipWt1hlMoEZTHA87Q0ADL7ZzhL52j4flw
e2XaAspEPLWPyAamf+YNqlYCO/h67XLdBnjmRWZkskeNzOMCpOI/Hm/yOxKDAXhE
GxoK1kbYUP5/SvhQpx1JQ/5X2mtTp6UlxVvg/N6hH9v+aVXbybCR1Ty8dxjEzdcG
E7tAtf8H+27N7V/DdFqbQsYiO30Kwha/bTz6BbtRvftQQt2u1zUcT7Oyxb8sr7lF
7R8sSVxL376IFSCJfwIZVpgNMQmRIJiSkNdC42XQbMEQHLaiyClI+vZegQiooCYB
49ZQoXL0gIYX3pNCVAJgYgIN3TIcxI28E3vVFQSsHNlQx1rMpA9ZKNm9qzdDPAMI
OeZjxgLjz2NP22XghnM+noW3otEcVqrDeyQ/UPLiFxjDwOHUa5EWlW9SxHuMElhC
U0EaTaJCAjWJ4APKnFqLlxSo977xK6bUnWAXhKZ2Uuk6UA0PnID74BoUnVjt1Gzs
IikW5FMMeJRKVjjC0OHhdCR7B/0/fhXzoh8kaXV7Aigi6rwLROh7M6CIfWlGkq85
g4eujkoBbhvMYzpR44ah0c1ox0HYJstwKlrVKGj6dufRtI5mXrBYYVDCn3RZz8lM
pNwU4mF3SzpQg/Pk39nAh/Vl7VCgLe7x19wF594af3M0tp9sbW6TxsvfpVqmzmuA
IDFfUgTn+tALaAqYtjjLAYJvP8lNgjcVik24WhbipYKvisc3Jx3C+nywVDZsBd8M
CnSi87qDIAD0tRRR0Xg8jeXb5qzlxaOA+SdkH6fIjwN7wovM0iRSrmPEieFpRtuB
3WQBItW4DU2QOoAURj+nulmT0+oGXIIB59y4O+iGxtsBigwP53DhEQb0Ix2hif8M
6KgeTkN6Cezc/EHUVhVKcH88uzrSBZcqC0LabjHBPOaA74afYOM7nkhUFOTeJ4ED
onKnTWULMMwbUnym8DzX2c7OkCtZMELLkbNuW33+0pqRxPGEadcfX30YLfpbQIRn
vBsffbGKvTi+0cr3nV8pvrcI5ZRbLepKOaOZNGuIjIuOWf6kED4D0gEv8C185WRk
VBhMtCNiM4uf6I8FzMPeswgVPVN6TgmM25oiwHhgZVLYxlTWFXWitX+0FOJ0hQoE
MN8i5x9j1e9QeVErWIjOZygMVDomNz6SPEj49PVAA/E9TW1K9dYT1EQNdonLcy1i
oe/dc7Pvs35eNC+KAMXy+zT62SfRsLXfqmmjGVfqdButKcwuvofXGH17AskTG+ml
T8sM6OvEPMaKvYYYwTt0y/VQ82TvzwbVbEPWoUHnZwXCOI7mZi7pu4aOSCYK8Or4
lgG5/aUu1VjPbUplotea4yHUxWqWyh9yxDWfiHNTK1UcDZE3Svb1xuXEjoQD4m9c
5Ue65xuCuzNRc2HxgSpLeong7BSaDFl8+mtiox5sTnpf/X8wTwil3CRPc0Hin+wO
ql05MO2t3ix9on0xWjqHkEAvrHF4nTTADL7LGL7O/YBybnXZbb9DiZn42l/10qDW
hbbtruwrKLeQEMi3bdV4AhE6F90/5jUTFiaNTYsle/LRQNH8TfLx7c9KjEWOvWhE
NM6qa50tiw7rrZhVUifXWkNnEgYa53PzqVC6jMFkxcivrcbmfyyEwMzKOfWn95/3
9Ui4GN/2Nh+GcdpHjmWwv+TxF6xXdg6hGFTHSL4HfgTQpg8N9nTRZn6xMaNBx+9f
/gEaS0UfQPSC1hfFAt18fcbbDC7kN8J9pPpiFoKn5uFJ4iQ/jdIACT4twlj+xXfP
88znQMES6UDmi1MvnLPGTdTJumyc4V/mUeL52J5x9YcmKmRYFaA/jR+zHqyCCpPv
W1PeJmlntybbIGywo1naT7kMmdbmREqSExFwipDiQGmL7hjRA1WtOQMqb8dTUZAD
9uaIH2R1osb6q6wok+bolOW+VCjKLLJSm7Fw2VRT2g1gAZUJ0hdRJB+6WpNYwrr6
FWc+wATQ+Aiq7/loO7OJCn5iyobjIIUAufrsyZHx4VnkkZsRJaeGSXXSlXfT6n72
PeMMH9rmMpTkljwqkNKKnqnoBct7IcUuaaz6luMTo49/SaspNCDs7yU1m5wwoDWw
AvlUnXsdushjaLY4H2NhFZ3N6CTqBcaw9eD7lxdH85CAdWoCOS9zVQmSnmDQ9JjB
HjWvuSwVc6tBq6xms2yBFM7ikf8qITndUCOdr/szBkcUWSZCAEg6HJsg6NCfVYLP
V7Eupf8pLuN4QI8idqmgnuHCa7YeZSSo8CPzFhC+aBE3SIMTG1HzA7FD6zWjXMii
PwR6WjBKWrAnLhhrLyi1xTimDzk1+D5RJ0vTjG0vmQAzyN2LV7Cq7OFWtJnGjdUB
UPkPLkbfsJ4sA3pXA3Rb4hGODREWG7xD38LRRuImjkWziV53RkaN6NeINsXHSw5x
p+B+O2km1KPZtsYqj59midZ/zRw2uZKN7ruiIa2zXNXnkjwCnjg7FSFsjw2kbK62
Li4n+pNulw8DpZdCjIRp9qcBBiwYTBYcftckaRm99gDS3nfCcuWNKxlp3GCPBmZw
snaaR/boaEYUFbbN+jOyCSheqFRjmsKMIHODFmytmqUAm0AHkp64wIFiwSjyF4Hk
tuXye+DvOQmIeEH+wg+UG4KIE4rOC5Fkxd8FwWd2lCjtWcGVzy2hP1ajhZcsNcyB
zCe0i4enZsxMejWu5NJ6SH/W/RSL6YqzuCE40XnMqVyIwlcloxpXWRGx06t/q/oO
Ussle42TNi9n0Zj1fEtnQtBFec6jCM+pPm/oy+nAEcTj32RYXPCDbCAqwcAFI4QK
0ei180/6jJqI/dEsfKdHy5+aa/F+SMdvCJCqaB9E2FJryF8t6lGebldPvJ5Dc6yl
QU8mvn4MhL8mdY1FS8a9ufRCro7mhNgDyRe7zEXFnh2YaApYeunI271wYB/pe+Vh
5ZzoQ+8Gyy9u2jfulbJeCddnBYZMJC0Cvnhts1OICUdvzRf84sM3bNfqAmTu8oCO
hb8vSWacm0f0VaN8xexP+02jwaxKRFkCEpOfFpYjIR/8LGoAiowYtDe6NrsCubVk
qEBW97B2uPbeocY0KhlbI9rF8/D5UTrLlsaKsLNkGmj9bhAnxZWKNAaqbl4m1lFl
/tCXsQ/N0Po4sxgoWki4JOSapGRyWlLVK4ZPGeW/2aHGn1wCyDzHnptxhF7UmXG7
dbgSV4MObwQlKk0yD8sDpLg2/jB3cQsGjfeqqT8VxP0EpLa5GV757tra5Zt3UTWT
q+HASbgMxAYr3jK06kI33+1TNUw9qxcGzl2/Q5L794fQB+00VTkvR3SBtQS8ghX7
Pur5s5DbrTraqd/2D32x040k3nLck5RUiEQDcwQJu7N4bmMWb4wTjd6OVToO8qmB
uZuxivwJ+ta7ePAtStMAO04KpEAXz5IWb4uyZ7zCxwI7L0RiRIHs+Gff3YmoJMW4
kiCnblTww50Zp2BBOtb9VCsWwDqUVCwrlU7mJDBCeBC30yEVwa4+Xjw3CfkwvjKc
PQaQW4yYB2QY5MronKENZFCau1LFgal0XWnANXNEv3g21MUGf1LbSnNy3/KecDsc
fmlzMGjQSCVow+sWjBx8SF8uK3Oy0prIu58yA9u6qGkLowjmiIZp0tJJQ+KLBXhV
DUcv+R4ru6asCWnPVahR18JdC2yLGZHjx9Z4fDlTe5l2YEbZG2/Ee6d9pbeHqXO6
PGMZfQeeBTIc8WxkDCFzUQRwXRFo367iITrZ8JboejsInnhyait0x5qUqAWXpU6K
lO0r/SXaCRl4pWyvtNUGWCPfDb6reTDlNrdICZCKd2ZwQtk2rONMQ8+wQvVAOY8m
VpJ8kB764o8tQ/aHXd6zNhkqeiq5aIBOmkIDRMC4PMGAwqP44CgHyLd8RsXHh0km
Skzk8/o5tTFBTxOjlcelG1FnJP/LouDQPP6uIt8Y5rjNceeAkRwYxDBEurmaNIAA
oBY5dDzh/2kNs1guxRI+KVCzhWDyMisShRjEpZ47Kc/w3igHCiq8PofVueYL08F3
NtRMLDss/f8Ci+xnjU67QmBvo+S6dfs/PvWTdNV7VcSNCRhUAdVKVFA27ptf8Quj
f/G4nmR6OXNJa2RecyOrXJn8QPWmLZbp+ojLInYZfqZ3s7trmbu+IeF9mmIyjV8m
SliiBxhuhSMNFjoN4HCpY1zRmjRahsauqRvaLXLoPQdaIiEBCZ03rV8BJylnKHBg
xpZlWbD2msrkycMuFhYicRDI5otRdcZpYp4RLtAuiWqctHpLvpC5lSpNU2cYaPAS
O/dX1AEWXtCi1sog/38ugXn9Jyi1LTlbJ/l/tw8Z6Gs3ZB/BgVGDZXklwyUYr3ao
kcqQ9IBnOhChWE1TNb3P9k72F4thEKIn+nWDjuiokgQMWOQdug89qy5VpjeXHA8p
RXxQJMGnCu7T6wj1MeApsRQWjppCPhRM+nv9HM8kpgQo8mHoNknHogdL4j/IbLtM
sC+GwjFVELIgsiZu/vmXhjp4BJ5EUk5Wk3CX+l0dr60qjfaupQO4Eu6/BziQxsHB
kcoko2LTHjGnpbV7LKG5eANsOhDRfhAulkKH/pd53aAY3vgU5OnDv/pc4R9wqEYv
9WwVSOL1BvSZqWCXRxaY6z81FNIvENq87cvrM8UUmWht11R2JdMqdwmXcT+PiRBw
Qgn+cVCy+3E6cojmqwqQ2xTVqiuLjrXKJMd1vGdrL41sh8G0ArZoGvUWIK6V3APO
AZmjt4RmqSbZB9jMnQOdMEY4KWGPVG6P8mijNz45BLrXUvn7Livm1VdDPOL9CvnE
hwmWfSIY/JWVPkaXnJG1RDnHs8wfzLLZ04c+Teo4dg8e+Fv4AITHoRG/2/1se7lO
cEu5yKgSWeQDON6nEDz7QRp3GtJQq6uQ0eYJSdkgNffB6a/ognDGkP6tHFML/1NQ
6OLD30e37/plMbhgd2OHCztM+pAgSK6RhYIMRoKvcvCtrmcFuODbBW4gtJCfn2mk
AI285zhrzpQ1DrEKVoGVqEuzX8e+uOdOxqikYsB87cF7S1Vj3iquXS5Ffy5yBgf2
e+EKzZQnmgV6uWACUIebl4AM6mAFHTo5wK9kBmh5E0SbIZY82a9szsbTMRcS7EGa
KXY9GNxZI2gJlVNpFJUS5XFzTOF2KyUtNq4GC8NtJvSt6+8aQByN3TbpxRcxons5
OVR63MmyBXtvWVzsAVRUMugnEsVzKZ0bWbmEmYotsF3iwV6TbKiqRIsPX38zUJsb
6qmBghvisCOOBO9hIrZLeMxLJuHkGheK79+6UYkbl6O8QQt9rkTedFrzb1dROZ+/
OOivJeEJw84VtzsSS6i/YzNEZUOGycDK2pREwO4Lx9vJM7HaKJzlNoR/aR6wRVRM
2dJ4eOzmy7unG30d5TcYYyniK6BfYhXNqSKlrGGrHgLv4dpHUzoeXMLVdflQP62t
r9KNkwWJzYgblf3wNXigP7Rt0wqJszHBn5EHbtP3qD0NFBSmfAptvkbCBIXfuJlM
cCRnNVOwm3GcpBMCKyeSgilZrgu84UNhnLmenEiKHYxeYrv/l4N5aNdD8UajaFvu
yCkMOEarYtYN2ItXD1aTAMrCnvROi2jTwHsi1p64te+WrJFmK9uu+zZbLPuP8l4L
4fqB8YO9SD8HUwdJjAyMf0pCzV2pCcy6thjDr+MX6/0G3wfH+JFkI9PU0TPAqicv
vEY9DvyaExEk6hYMuBTEmDK7mkJtSjFEycZqd+5IpkC3Lq3AgAN8lNpje6Xs8249
PWZmmf4j0SazTQHFMQi3/u/H6FS3raBedi69lPsi1Rhhcb6E/L9MsJ1nxmEJprFr
OfODbbcs4os2kdP82E9pJ2gHKkzJZ6fpoTo7UYeUC+S3niVblxc3L5s3PJAT2vfv
2jlp8LwukFr9z3gLE56sAPJDekcwyL5IaaSArpTQ3vv7KuvxNKmmu+nXk/s01LTa
PPZeZ5CZrQvLudKh920MVjkAadgKZiyJlOdzMqIl1PbFUgy5bZrUm/0pH+QivRh/
QwWH1iuq2bxeXuRuJ3+KtMRJVz8V6T8M3cwfQ77OBOhflbqOGsDkD6hHCRXe7IdW
gOH4d6F3NECElxoTQAOczS9PA6wPfcgn5inFT/OgPVvDuGceJWRuBVZSNGW5dlrn
aQD6CB2aWcDy9dEFAG6+2EVB+/ATfrIzGhB8sqQSrzATsfSSkv6KEnH/lJKcjYpR
aFDQlsSxmSZ0YxfwiSLRdpBgLkinooPoM3yYL15uqjIgFTcED7UMI2YnZg1pMcWG
uJliYp5luQzXGDSD/f8KUlgQsnCtAtCLWZ23H22G+BjzAWxmHFwQNTh3coQae587
Z+1MlDjiIMJRT11NeJepYWjnWJLw1Lpq19btzFaF0kWVtp9qEqnXnlZULFzLMErf
UAMH3+x2yAQIlhrvr6KgTdljAtCIZjMn7VzS2oy7OJcw/20pISUxtoko6IbZB/ok
yn5Ca2meUFP2aWQwQIXtLtFYEB6JUifjdFT+X7SbdUk2BSJ0RTd4P8RMBlCvMbaT
7jLnTohxXPvguMINp8Pz8qvyw5pQ6dUNGdGKvstBpZBqNoJ4aUtCPEPkIEQ0eaow
g+sMoRTunyuIuJCOGqbPBczf58VudMb8Zbrn9xBvThRk0ChPnStED0Qw+C6t1CGx
+bq690ROhCckWAx4qUs8JVCK2rAvTg8e6uxxMwwovebx+ttxlpsjWlheKLkfrnYv
U2KMuDdL0ry95Yq8firpDnwAal/gZU39k4jFho/FFVNEvkTz5xqrYwUl6i7DEGe4
c9leYgLMAiTEOag9zHoXO9/ZUJK4K+VU89ZTTI1OkFqoY54LNXI0qyR6bbO2AK+0
8PHdVl8vNyznT5X54Jrhb4PhSz21iRoccQVLrttxMCvxME3ceQbtcbHjWU5mofDc
y1a+BYvP1Iz2xTYUTfsQMlvRPl10NGfzerzRwb5ZfPdzCB+h/XhCJAkFOsBDj1Y1
bwBk+qhgARe2a9ZIr5XdoIMBGgW67eT9JR/FGjqb0Wb0O/7e2oLwEenmaOPxWqwR
uq/1XOI9TZnyXd/iVWZ2HBdcTqOhngW4HZvZ0UaMphdrTtfWYtRsah+qU9/tnUq2
mM5v09PMltleFcGhAogjmQuqiQIoaLzALr4P3t1NcfmGvajv5muNKyaJobkPVW47
LK/YjeSVngfnNm3Ic2jvoo/WgkC59CC/rVLZRFdxQxESq6Y34XMlunfykqxny4CG
ez31ptl4APot4YzDvCHz6p4OevSXQgx0eTIklJN6Z78z+9K2LrUO8EX5uXqogOXO
9bJp88YkB2u567fr2Qx/s1oWbMYX93/rLFrj5ZE3utmJDeaSIPwBLdVnRy/3zvNH
i4yqD1GP5bbs+KWmddsN03mLXQI7wLDA5exBJmyNQwlMm5FD/Z7N4+Jm2Ey60IT8
cUa08dixjkOh1r//kwrsufY2NtOeHigsQRVp9zquQ/dLbS3yUm+H68cYI+peSw29
DSFJn4ZPc2zQgc2mGuwYHzY0VvLjMzK019QTgl8wIztf6m0yhxssnnrwFubdZy63
f5128GGk62WJ//Qo94OstvHrMBZZ4xw3xGgjCwWr5fMSe8eCV9tuOzB7MP0CjzXG
lxWEgWtiLNhCt+5kQuhQOALWOlW4ievmygV36382b8JazxtXeedBKzswbELEcEF4
uKuF+LyqeZzENEE89x/tBND6nGO8XgTr0BKF2mWoo9qITn0Q7I+xNJ968FztqGlC
o30n94pxk21xp5XqXFBilv+JGojwdkTGiqCLQzuBmY8SwMzI24HLDCxR3LRZro6h
8uw7TSi6txJpulzH4xPbKfsElkYivBLNy7cLYgoFsRz0Xopeuf65VXB9+aF6WfzU
oLLyMOGYZoeXP+SX5WWF1U9fGPQU3K4TWt22FoCRibOMVahfEcB4qoFDX3n1L7CV
tY15hCCnuFLIRc3O9ckGCYedyHtApuupG60gD2H3pb4CG3U6970KdoVhLxKZ8JRw
s404Zov0ktNVfp9TidlEm/eqrQAvVkG/FzOkuHzykH12DQXiCa8dvQpJkWxxY7jo
VXMd+CYYYvLjoTM33JuutDm1WP5v6xPrGx30YebU3sdOuZUxj7Sj6A2zQpk0UXeK
6fgmT0hxaQfndoAzZp5C7M+Iaxg/Rp434lBUKmCGEpGvxAEAL0japsL7IT2UN4gm
58K55plTw/YtYNFKKaSpHDU//JI/HVDr5etGbmLh5yUhfQNMmgf74F4OnsxNu6d7
2BDyEYoYrDDwO8exqyRsL3R53kilzuaOPgWuWYkLwLw6P824H03apv4a61XgXiGb
FBRmNjPdLdLXZsl8TmMxzXJ9cIHDu1Q8IYbf3I2XMebBehjBl3aXEWPEJMxNnpcZ
GmOD1cLudUKoAR7eRyeSv0Jr/px0zDLL9n+OhGLwYyk3b6Q1iJbMt+jaxK5UWjPr
apo+v82vgiNn3Y1psgqHzk5BEM1HqJKgONxDWHWnyG4sa/99CmWlO3U9sUTWAWnX
aQsC+Yra2UDbTqjn+TSZIxT5VplIDXAWN6+5ebVl2j74tYxX5cEKsQ5c4UAZT6Ec
zh3vsTnrLixZz1yxrVAtYbp94BHNZ5ZWbFHUH0Q39xVJ2Egp9c0TojTTDMbLjbsI
bgCAK8R+rpus0vypFeQ+Iz1kmB4fLPcZP8t9KAc1O4SdWQYJFXbhRELgGqruXyMk
FyMi+GRXscK43bg0cleoMsCxa5YOa+3Df93GayZhiFBr3k/Pbg5dqhWTLhRvWqPN
kxA658fiBlavRUF39+DIwk53YEmv5QVCu/NkROrcmmT3jrGOOmZIK1XiKqC5O9tP
oXW1Rt9Zn7AA8HhPICXDBHs6GoYVNRpGFEidIjNv6ChP8X4wPHcpwY+IENR0cm/r
402Z8AUEarK4TWZilI9sekRq2gWksHfv5yLELFAuSaHTHWWXVmQK/fcL9xhJ2bki
GDhWWVJ6qnd4vSpYE5GdQIzTSk5KZuFU2DDv+lK23+ZavPeaioc21kHe9Px0uSdU
iyqojiYxOiaSeYPsSZRISRE8m3kMOjBhVvSRHHpizon3h7ODQ6ILLapVo6T7G/zP
qRqtv9oB7/japmXA/icJ13dSkGfBjV8mjMKkMy7OmVs3tKgrM6O4eBjXuM5xk4QW
Y5LndOkbDIIbN/ooQXoimTpw/EYUI4PacS8OYmf1Bdovj/WZcHSwb/PQ5UY39nh8
L9u1/EjntHduSue8phvca4+KwkNRLpOnXTxn/+wo+oYiyMpYDroczczGoWF3pm5w
LZvuODcuA4XpvrdRA9FmVs1HfP11pkEBohHnMC0yy6lIzNgRtIQX7unwLEIva28S
ERxcOKKJ4oVJbX10SH1iLLoB8ZVk66QlB14UVx+Y8sZr2LuHB+eWYA4iALy9NQrJ
B9zyfncBExZLyDV3zAlzfCH2K9y4AGXR0oTleOWPzYf9L5FVaTew6Yl9IRA13SX+
nUbK8oo8IJ9QaE7dgzKMrDndD5h62MS/wZ+qx5GTDKIpdR4MEcHUpO6Cws2te5xe
YrWmvGOT5IlrLqST567rkOEHtztQ6F/vOCQMTp2fjTk5xuDo7HBT4Q4JZdyXrEQs
5yV/TdHE5t53Z8Lyq1MVOErlUfBQ8EymXClHTdZXJz+luJvIPG16vUp87MAAPZDz
ALRZYAXyAymxnauZ5TmNz81faqifywxFZJXY133cGIUdPVknj/XXKJbJHEB/XlER
m0RXcBE38Ba48R3e+rfv6jSSCoC4DE61ukLETmBZDVbMa1+YNxoOwjVMMnAUsugt
rSzJUZYzxi+EJHGAd0Q+F6Ktsc5J3EQ72px0f6Csm/x3jA+Jci3gi7XqO8vVCc3D
ACJ+LtNhkg08zhEF8lvg0j53japFP4TCrije6DeL1FvNMx+H/NoSDYoiQAVmOP5+
xW9ShT8bQaaRxL+yU20xtT/w5A8upaGEbipYLUzHuQGjP3P5viw/yXt6w4HcySe5
y+gttf8/TOrnyFA5CLJNk2xqFhRSJ6zOR3gKGea8XFoSGstMdfhilfTTT/6FQ5Ig
F2HUZWLJog7VBi8TGFMEWY24bdFyFHpDH1ZSoddAnfL7mSRai/8qzZyfpm5m8r3N
OENxHoS555H3dj3C/K0zA7mcHnpSN09Huz1DFr37b3cqs2Nx13cWoiT+euG9f/ln
HyCJBdiy66UusrrDgAUQ2PFcv/nZ4LHTBJJv1L+8SDGw/Ju0EE0S1HtlQiqTGGpQ
UpxlA+xNHUG6G2FNAmqED5reOqpas3yoLY+muFq18XFguLiaDECybbe+D4RBMiSj
MfwPCgWAyWSNDGPTqmPqw9xVQ1fxp2R6IRtKx3+3HlgmZUQyaHx4fL1V0d2bIBJj
A5ktdrKRRnWWKloOH+mbpyzX3NsaB2K7GmU2AG04UUikTFSB3mNEWf3S1Fprdse3
lTU3W83COemx96kKMd6gdVhkB++VL4njTBQSaUMQxC+E5oHcwWdytPgPo2rD0gUw
UDUdr/N074ryh5XYcIcwFoYtG08N/MvHPoxR/eEdHZ1JViB6IHoCZZzMtnYJZ+Z4
lZqdNDU8wbunEOXiJyXSaUmgkp/CtFiTYsPwzRyGJYGS9Cp3w22KD+QmHr5PWZwB
MDudeBr0XAb3Ywt7DnawNvsUHAopVAYcx2Wpz1Xs+QHIMW4SOIndk/gXqY22qja0
ooXCuPluQAmFsE2ckbM6kbnIIZdJn4Qoghd6vN541S53dCr3Ff7jN1NkYyg9UNG7
M8hmZRGxWFG3He8FxVIQ/mDm+y6ZwI09bZr4IgTvbkWEVs7mFcZR3OeoVzSJj0ba
nvedbiPdBvMfVIdGo5CKSXvysl5wUefql5ns9yIVyexwFHvVJrBEt6BfRCpJ4QMZ
ZZpMHfo840j2wkBN49otVgNVOBvEtFq9h73DqycrxxgSzO7Da5G9tpqB0SpP3zAu
o9v7qZdwd61UFOKlKws274qo6Ycqx/Tq9AEoVjgB8GZYTaFLZ5LFP8gpigfBOt3d
4B+ShjpDFDO5kSiOuyKVt7TSKgZsRplWo4M2bMC5iRO2wkUg84bX4PhYbxIdDozt
hQlpzFYg9HZTIqCtEmjfcIT9pcp5nKLkpQONr85PLAJ2J6K2La9aDn3LUnKD7Tak
5wp1F7b5o2ZmCr+vGHRAYisKzMg6QYGlz3NAUoZIwuacPD/JeipKNo60hxhbtuIC
Ha6dI2GCZ1mh2KYM8eQX7OIjd/PFN6xmcyd2blNtVzVLSdseXkf4GD6Dxq+I23nw
XUKzBABBgpv6xL9VVryWsS/RCQZr1Bz1tcYv/3Mq71/hVw48cw9iT44NHWwcs2Qs
DI60Cc2vrnkHHkWQ6qjr3tD+/q+2mlqymgqi5bHoeJCG5FjeXhfeMyGAnK5aYN73
aIzwbAoHzgD7e884lau13EhLRc4p8+6I/TzszPZDUjiUThC2Ee7tpp3KQBi7rb4I
1n/bHvdSqzKB9EB/dAF/YBI1dko2KAdPwXPEfABj6gEMwHADw7ZxAIkFQXXLSwhH
dksUk/BYHhP+kTchH+rBk/vaTGLeJ2Ww1nl+7yQhyrYPEy8Q9css5bPVaLm/hsf6
cQ9t7rMFZocF94kjZN2PekXxXLvexBUFA62b/AZRHQXXc1kJ4TwdKmE4ygK3ZlhW
qQ65+SXZ5Nf0c2Cf49n3OeFcMaf3nn/2RudvRUgE/3UU1TpFP/FPJhhOhX0TqHMf
dEYFLol9fjHYBb+Qu302GjMe/5aOtwpOmOJT6XPLjjJVLzM+MsJkbFSivJOszUNw
8DxYWN0uhtl1BdSe0quo8QHiOjv/alJrhUHJ1LufQfE5Z/gI64hjOnJtPfBTEggl
/ZLdLWonXUowUGoEeiS4uaNpu6pAhoynngoPBbxnUbh9E1wzkR935CmJWTCXTG/X
OmdT1+zS6Uj0HY6UhSiWWm+BYe8lbebfh0VcL/VQpviPvpUSb10FNP9eTOBCX+Z6
RMAds7/jtAwglnQTzupZfvmyDn7kQP/bCKTpkuPYiCGnz/FaP4NVURk6OM2rp802
BzsCKJeSuVOQoBJ851OyhEqrOW01o1IOJ+9b52uxU5D7omKVO1XcqOwii3LHi3jC
OvdQlKpXcMgiDX0pc0xYsxAb3OFR2VasCN6Ley/FQYGTZXO6h0XSexrFmq3SuPgo
I8GvprNbpSUv/tT0n89Q2d2FnZk28a3l2R8ODEcS4IHWMcVlocc77uB7H1ZoV/ZR
U8A2UzgRcmVM+Wm8dz9tJmrCctbNkFQvxNA3Q3Hi4r/0KCcFGa1vsmWiHnx2Z6ZK
C8iG5MLx2silVfKE35erlbLdJhTw4gRuX2VUvrECPeYlAm3mIC/HVx01sFJO3Jpo
QqsEmVkZ6D2GUlh0T6j03UFkGgOmsnJXFAJ+GgTGhy8O/cRWkf4dgHCOwXhrpfN0
H7LleR2OJs6GJxOL0yiUzbRHDOXFbYCwjk+SRo+iTzI3VwCkRyEmZxd1JUpjWg5A
9SrHD1Eq95ANFSldHcogx+/SxPg8rAKjLCgtAndf9XoE8breNnsVuO346Kt6/Qv1
j2kBZ7dOgNrZ02gS+T7MItjDJDCZMcJI7gSA5cSAIcJheYVcqFkuiJBV0JLh5Z+T
j+a6zosS7MY1pvai5q2EUO3+IKmZ1Y7LZP9Ib5Jx7U0yUs4MrPFIKJHojUGHaT28
UHKlXZU9vxGHMEOZchYylYmL2gvL9rr1JqFTJPy0wKMOmGpe6BwJGR9Zfwn5/bm9
+FgE28bCaORRydG2YeaXboJwionurShaxhfiQ4w95AWyA5gA5jGEBv3t+QXlivZ5
fTsAcCyrMptGpjwtVD8Nmlmt9wlXdxQ/0L4fce9Cdp4SfeXgic7kWTZlqGSnpl0O
gieaRH1jOgPMe2bjxotM0Ms1FNBYT7gTg+3NjI0NMoV79pNyVsMt1YJZaKfZ38bI
JuqeaY9Woo6zEepErOcvFytEjZLVqeYyA5sA4tCpGpdVTYVaUBalWp5Av32lsN5W
l5gD1EpwBy9E71ITZKrQsQ97tWIhavrYtn2/G1C4jEEFWtw54LpjQTf+/gYa0Gki
63M30u53HUmcq9PZwre2krrTf42fr9AGEOY5ynYA8++gFvrV8Ks+6nKXP6w2rce7
GKgTQ36xypnWK9/qb7woJoZ+8F3ZfPOq1cCDyG922THzJpyEyKFFfV+dIuxvyesp
5UlLSLP/yMYW8caBFAVmGrcpvGGW6fru1Y8/SOHkI/gvJ6G5m7lEyjgH0lNkY2gR
Ye1WSJeZLxKIQMZZspbsUj338/6i+Rst/tm4LwzI0G6HhIXfccLQVUAPHwS8kUJi
fQdJD9j4rEiv8z7DyhfpuhRZLPR78qMtA2b3hD/jHh6vdJxFmqjD1numat595WU3
se3JEs5G7tYLQkb5xXyJcmNBJrPZRhec8YcCtR3lModh0Ud+4EE8lyoOpuCCocQQ
/Q7DbBdSO2T3gOsJ2FoMuj/3LCWMMJ8ipOy5vYs+i91MHseWKvNz6fqJjbbyDscD
atmlTs0niEubojj/I0OEQMfOpUj97DRsQWhoJ8qlmFHDgYN7CqKymP87RpOXaOeH
YO4H3QQWKd8wiPUI3WWC89oS+elELIVgETAVJ5Ut/+0cp2D0GsQL5Ky5r39VFlU2
460ToPT5rnesL2qS8CfZrxUeIov6FOM7cKK/FcvXmSzKi5nH/nACmfmQreU54/b2
c9Ufd7z0Ixuso5PZCLmopgZK/ovZgVKu24GS4FIA4nKAa8jwKw/s1XBpfUtUieP1
kGeLaIzzOoNQatXztlsfzWZ86AYaozqIUU5eeOSjSv86y4gYNxopsqkw8HKqgZBt
jkiwvDGLH7uxuZDNb0XIJYLdVUB/qPeOR/SeOX5Qlg8kjYyu0k/9na+542JreuTG
YoLBl1yQWrZ2x3fTfTdwe/UK0DDpd5GqbMKEkL6GWB3K/S+mDn9Imc9QEM25cN3m
Q48rig4SnUaloOmEpRl5w2r7/a3BRez/vp3vpw+0UWiA9Bo0TUvJ5kv7Kb2uQpqx
n+3LCzvHSNe/OtAYSeluhJ8iskjjv1NhF8iiTHiai/Q6cCmICk1iIzsruv/33WYq
3qO8sNhEnhZzz69FJXyPwiv4G76UE6QZh4G2JlKvdNChw/LkuHa/A3udb9pBK8HC
GuONA+OLdbv4fLG1cAVDMuZaCSZIyHGN37mIZ0I28kKaNA5wC4tSAOry/e8u7Toz
6PHreP2z+pY6iX4PHfYJykwiK5//shhNpJc3gnMp2mEiy1wnJex5N7z/GntozBsb
KB+nKIw6lYDM947Y3MFc1fv6jKEvQchOA5zRbUVOu9dcZmU9RWjRCmD2YDl7U5Qp
5kyGZXkCBtn/CNarpWjNGCu8F0Mv8uF2/wR7sQo61r29DCPcbLOgB7B5o5+hkivl
/XxGxt9LjrPm5Y6ukcqrOrUxslAUgOd04H4fTlgtW5Yhr51u8lVOMctSmTti80DB
xgmGkv1s4WATz4+pI6g2Tn3hUTDBmqByv77KwhmK8xsC8NUgbW6V7xQo62O2ExEf
3Q0IKN+NvG9cswvBbdyWbGaGF+dzVBG6B8I+sYt3m0T+wCf/aBD6Bm/e2NAQFxXx
4vCKzssoA71r2m0IbJc+K7UdL/0QeNUzz/l5kue3E+LXqDIsoQ3PQln4EmCTB4rU
d4hO8BXpAWcvHS+6AAmyOWQgqo95haJ5Q5p7OUZPZ9TaDKYLPl//RNlkAg8z6P+B
SkN4Uq7sdkc4RUNDH9i8BHe/zfnQEY6kMjjXz9zl+yn4Y7urfEzf1FmFIElSlUqO
YlPueaa/nKGEH/tapfZwMZuMqh/ClbbVjMhDHdrbvUGcx2qH8V2QEybxeITh8eHF
JUBv+XiR89+ct26tUxxlKP0T/pS3BNPbEeCc+BDUC0MabUoNsl8WVb0YGMmE3mwi
liQSn0SMva96SP/CNmzHfi5AUQm1qlvMMYpKRUxCVRG8T+m2rj/SqzM/jWk+PzN6
087fLR2pmwg4XBuQ4jecgYUSmPLYNcrF8pQqBKPYhlSMhpZD5x3qViTKd5LE0dpO
G8ontwIa+FkJ+90F6oPyJMvC9Um8E/r+qFXCBLkd7Bx23N31O/UeZ4MOE1EaYE79
E3Y1wepYQiLmWSVjCcGEZ7Me+9zEPOAldcyBypOCvVjBRmLICvTukqkOG8cfva1n
OJRcb+mqBjS9jMeRQ0y2YI32blcDuvAL+dBJhWQvCUxlyCOFbu1A7MXgJxK2KyqZ
Vw8aM9fkntTF8/lMhaMVAq9caT0CQ5EC7aucRiUTOU5XAHE6XK6Pz95NpZCMhNE3
OY3vB2H/qVg3Me7zrtTsvMPq8N9P4dT2cY87HaWwEW8ULHlQTHDUryt7Rfw89RvX
sqj1kFHAtWsnR9QMqCNTprTOnUNlZSK3N/tvigL0LkPi9deLPJfgNfXiv+WQGNtN
k9+P0S+8JaCYTPwFUnH0YUWjQAQ5UaONkFTOSGkbZAOU32Ec/9ffSmzHBuZsPDj7
cA5GohqqwMBq1cJERbP9JbgE0oJEugGL4vF8Ozd92hkDQUELX4DsRlwOQAN326ys
5r58C027RFkOFHnqbqcg3BIn3wsWu3MsMyqw3F17FPeQbyjclrzpm63cgO5DrF23
jRQvnZbwI0kDhXqa6XveqjUFOtd77SM3dAvhIawZ8lZm6wLcxd5vZZB6DJpWkCEt
2RS92Y+Nolg4RMiwVTofJxrr6woXFL3x85eDoola7GesIHzreMaD9Ip5a8Y2fkFX
D8N/ruWGHqpNhq5z+OVKkEaJjmMo3e4YGmmcJz+5jiv9W42sAIJK/HWjuDBMJrtR
XwSLJaBT9D/oF7Jze4osofZKxWJ1jkqCJXAqp0B/XjIsbVlpStFFYWGfv+/DiNgG
c++lNr3smfYNUGha4Wg3E6b5ipcJrn8m1dudG672aD6qUes58yPZsJV/oMztRmQx
+ztizQj17gfb6DrPC2P7ijrwoNwTGhqlS9OZAYfdi8C23MLSIQ3FPbcanIKyiK8A
Dlpqy5SQlWueC5Y8pkTiko2vDn+XlBQGM3pIjBLlEFbPLS8SplSof6acFTIGIfpE
NBRVIFP21kaEm9HvB2NIyQkVB47JdvTuk3WOjJLG1trjz1qlVxUKEx83XgTtAIG1
oR1z8UFe6lbmnO9yugbvFXPUaWcIZWOcJdmQDdakb2BZeHR+zuabUrmPrAac2WAt
ZreFYB/gCuqSbelfwuArTvbyvdHotLh5VM+T3IzcujklAci1y5y6QPdxN79U2hW/
p7+N3PL9HNeZ/b5pyTnTbidBokL/TrVpCOvip6eaMWdouaBGvWzod5siGrs9M1QE
udznnMO+4n4wF53hNYhl7av1E4kqMuDSjvUXZ6PuXyoeIFSd+CH9vohVBxe7nOYf
Ieei2E6rvDWZAi8kch0Y/FTwFcIZGUqdaodjI2r/oBiIoyO/4npqX5ivgarI/Qss
JcU63sULuz2d8TzTBzse+2zy8et2rDEjL6sCsPntnTOUi9K5ohFjCMUdZR12SD3H
8N7ufe3Bf3YZR5X0jhB1KBin0gsa9Iaetm02NeZlANBMe/kDm5sDmxgEb1g77lAM
Ga4MrUkHKOMXfrBdp1xija5oTJbSeyiCSbQ+MtW9MpXwW7Jp2XBenHyleBNHGder
OIwWHboY8BQGZccZMrapE9iq5PLdlPWRFix6NOgnElBnttp+h2WdfbfzCkTzqlbY
5c5HpnVPjQF9zZvURXIK6NcxcMF2TnmZz82nMw45Cs1kxCQmTxPx2cp2XZzuXpsl
M96KmwpUOrEAv3ESjwOfzMqXZBr7NDuzJB0Bv6pAHYgNUenjRETZONi0SR8glHD0
489yZI1Nm+FMZU14bEEYhaHPoL0fAvWGTsF9DpPaYrWmmiftQSGwYqgy5/c63u85
wsRUyr75kixVu80SvfyXSlptIS6yx/OxfaW25GufXz60D9u68GiY+Ndnz+1lja9X
ADdh2suBUw1UnsPTcOAnfcXldOzyGGplntmatPcgxA8Uy32eW7LXbXbFv5HOR79r
tfPDqXyX3hoGHv24eNLCKygdhDHN3Y4H7w47f1N541YhxsB2842NX5LownPuux80
ySocIdWGWgY2pVpzBlaRU8HyrrfKBf4Bal/zNTtsIbpt69q7j8G5oDCRTloih38G
ZwuwGUU05nK99YRBvXN4qLykkLVGwBq+prwd8k3YJtlBFcgJcCFKBnDaL08lblKu
dhifor93C/cfwVss6K2BX3qJFNkLN2ThNctJLmktk+ZQF69ZS+shr+Xiwj1U0fbV
6CXCGwj9nlqXMAS4Xq7kOp6LrRJ2Iq13nbaV3PEx0nyckdZSOFdeiYZREJe7Vw0p
QQqtPjaAfhby0eN87+rY69rBxwSJT+Os9kZ2hkhG7vjU6sF+IDRJnifri8m+o5pZ
MBdoYr/6ZxAA1KJqz17nvaRD05Eb6V+8iHJdVumS7I3uhpSlRePrTeJmxQgOzX8y
fm9ccFZhP2sep+4XobCRxt2t/k7NvfXh0e4H2gmMARvFCUz9BI+5R25Xbbd6g4XM
u+e/YoWa5v22sj5RYSPwDkzTdRX3Ei7RLcQ68kqah71at4qoOJ9bquCh5tXegtDB
c+UtVkSNGXlvLZXWeohARVp9x2SG4erFOycMGliz8tGQ39IHWav9dj2EOovt3uLx
164KBaFkJRT4gA7YUaJE2xiobJ5Id/fKRALx7ULA7NV1goLDSCh1iOfLxHTRlaUg
jnNVB82wimAVKt7Oka+bbMPaQuT3XkCwf1StPjuL3W7UvSVhhN87JI4ZUWisIvBO
RCjsSbjK3mdTXN4dxQaXS8MJu0h3RdSwTJ/N4MDKOoD73uxizq5tRJZsIJ109zov
TXCEclU/5aNZV/Hi3fdkMrUEGrmBlCrGfV50bvTGP0l7AWjhWm9ZpMOGZ+EQGObC
plc5nCGzWcdBEiI+edRQfKfPtVIo4rQsEXxnGKpMlWRkWhxn9m5yC7ygthYcQ1GO
N1jPFqvHDv6bCO8NkEGfGo5c/r16NZ28Xkq1974OskJQCyi8rbudwxkzRJkLtYmv
QW3zgDbIjU7ONwRof1Jt3VxtzG4V4FXQYHpWL5W9D0IeYV7+YkwTrXSG0SAjeaOA
QWptYxfogVQzfwX+7kS45FfO0H+JReSnXz2YqgsS0mNwvOE6nT3QACDSbLT34UVJ
BnWgvmqG9GnSBjd2rg6ev7AdoysgHgPlCf/P3zAbg016SM4S+tI9HeRLikuWwsiX
KJdUCyDTsCkH4nBoog/5bB5UEWKDOTxoIf3uuv8B7XiXaRaRKbGx/PK0LVG2vVjn
vS1OBd4UfzUTDzns0rU4xsxeddkVioCwFVdPemIRx5QzHSbjGeLGPm3MXnURY0Bn
neytEBq5NFhvrBZRSsyG3QT71KHZIvW8Cp1T6riLRFr54q9xBFEcuCITy5AR1VME
1SwGuv0fdcK9sf0qSkRmTw3DlfDVKOYHaIMYn+DINvBCQVYv2tdXURkpkkAxUcw/
OT5mx+FsEpq65zHvGncABQfeWng/HJ8ceXV2o67dQJZGz+mT3mOwzdFUKY5lPhp2
NMsUYk+TvCEbxtPtCFqS5LUJdAuBXNKgEajb5Xnbt7mc0mQbeuX1GhCoTHp2lZzq
hQrwe6VeQ6DMmUm9ohcPf9iEej6/QLLzvpsDg7ubn8SAloiTjGfO661j+6DthKMU
Cl0T1DbI4cNQIp/E6o8OYQGQJ/XgvzG7AGgDRqvm+cK45waq5R5/jLT9MZRgSnsL
8oh4Qif4Pv3d/1vAQ2eBAeABKb6peASbuTBkKKs5FrIpXsZWe3UvyML8TRIeSpUE
B6IquCpbAEFnCnwIbzI+rMi8cYpnsu6S9N+fL3xwWW9E0YtLqJ0HiIO/5u36rqm9
p8CnltEuONkvKTKCJ0+9ZbS+s+RansUdNKZGa/AoLhSaNhAttFezcBaEu1O3Ya+H
571KInS8NV8rNdZgf5yt9kbj/ZuyBKtuzf5s3gDS595uD4UYJxgA0Qj3klQqQaCZ
LGV4J/NJAqkrxVFsS3FFhtPo35GftSrHNa7N1A2zDpJF7NCQ9tILR33rj0zRArwn
3+t7v0QpI+Zxoo+BjUM4K6JbTC0Uq+wWM9QZVlSkP6yr8zmVAuaVVH04QaluK2HU
0FA1pEGFq/ylTYHtJLSqw/WwSVAat9KoWBiPOwoRMVZ1JrXoonGpet0ndbxmgRKr
xG1HM4vfzoEtCgmuunD17qgxGSxfFO7Ox63M61WdMzXBRhLAoktYK9wCq/xAwn9C
leRo62TkEK/ZhgBS+l4JGDLA6e/E8wwU+ipFfTgv9Yhil9+cQaxk8ZhW+mLxJxm0
FM4CsfLiv1msYkz43+GkGiXb2rVT6Y+FmQ0FDAjYmEdBORCLf4XdkMEpk0wLhZhh
w8rTp7eiXNC95gCxDjBnF9tQW4KCKLCS78XiK59KwGtRYbfuK5EVbqgnLe7hihCR
6q8gxBILq/ylnitIZoAkphDQAGmQfsentC8ImkqJelVK+tnVo/XbSx5KSFCDJ8KJ
rCX8XYUxurAXcVJI1pxeXxublkrCXoMkhBFfn6Z1rSCY4tCLkCIDhyaOJ7Zghjwu
317y8sgZKTLGRsWJFv2iGiYSWqTDYkeWVoF/EwDQisz0dRDz7EDbvkUaqWJW8wMo
SSHMU8cGg5QF/7Rr/0G+RAWo/cEVFv/jKGaW3xtVj/U2NUFIoREEPYKLHTBpcSxo
LK+bNrCjX+WLMsEXrC8kU6vx+LmrhfA15YwV8/sC/zBePQYr73w0KTr9vpk3KyAR
caeoVRPhDO90KlVz4nfLCrmFZ0/vAJablM0tFGSgOxbyZmCPnyXFUY/7iLwywe02
T+kYvUIdY3NzzuUXejZIVYlfnwKp4+NxyQ+w++2uXdEeaglrM9XmqN5WcwMJsGV0
ozBdwGpxEPTGFxR8pkfmWy3zvIkiNxGkP8BYl3iBA5n++kqpty0fk9F/W1t2BJUX
9R5KYZfFBivP9Gi4HKlv2mllFl47PKAQgNJWKtXA2ANeXskPCNIx38MKHAXFzmly
OY0RQyBfdR9hb2j6rdhPLSyO155Ns++rx9cM0A7O4ZDappu+xvPsUM/6lBAZ+xJT
VErwv513Pmc4Zhj2roJ9Slw6NVuuvzK75AlBRZ4SecMQGIXx12/gt7WVL09ZojaE
hMF1L9mz4iDL478+yWlp+aOvXdhZkziyvmEeGxAJGcOBFbnIx9DL9b/C2XuJyN3R
1Q/oBct92jL5jasUAHFaUqcSras0NuCNkuSME0MolbSv3htF92qN/tEqO/u+WU++
rQEXfSiJ4hZmNWaGKFYkrkw2Ug/5kpjqVpy9qoMduJHbbOehI2PfU9+DuR0kN6pp
G2fGr9xTsFX1aBcLJmFG3hnR05lXJjbjutlGESGABnLJiPw1gbraSSkRtEUTZ0Um
PKyzTxpINSFgwMeHtrwobCVDEWD2M01pGZWDAi+ycKxjfZP4jnCV6HrS2tqjuvzb
9HGTH+HpdBKnwtyC4LL1brkP6xUiH9S6uaSx8IRspTVm24eLTfVTpHH7iwzfd7NG
eiljnhOf8xq33OAJcnpu3fgyk8zVM8j5CB8+ZPjErHsqXRqCZV+Ns0LODSLOO5AZ
xfV4DkNXXZtogQ+FhHYARpfBtYtfDSU83XHCrV+eTu/i8yqTo37+L2sCGKweOJ/X
zKt33hB6QJ/AEyiWfNU+E39/0VfnvNKyFXEsb+hWcgxCTUo+E9tr4rbrHPJTvVCH
wrPUjhkjqbIxH51sGKOwJ6ec6+lvCGbThwzyV61digVhlpuSMv6WrHF0WPcynx1H
0gbAkjQTlRf44qpM5cnq868I7PSgPKPXVzdee9PrxPIBSN0NdTTFCA28H8PC4A7X
Mlkgh4i7/eXQI1V96cTX1xQkwZGVJP4qlsnYzCcmYV7n0mxjaaRXhKgfCLdWtIJV
kigyyk4gcNUWsVOzL46Dj2hpr5WhWmzkv/p+WY25PbOl2pPkqQtK8cdblWMF4/xN
XQFjDQ2mLMCwDWKsuuC1LtEfDkQunwLJ1KJytEBc0RQuWRMowS6qPL1Ts5Mq/DLa
EI7O5Ny1Eg/G7UHH1gdGMv96luCjY9nGuUJRNkyLwBqCQ2rPbnbVgpnJFeo1W+rP
dguayufD0JEkl7/pIthF9CmGDtW+NdesmTEQ9ccsdcj8b7nW2iWCbHzGRmnCZ7D+
65HsVcDZz6HhAPolhTnTDULKLxL9u00GB3t9zyNU7iG6/ld+wT8Ny433YG4XjZkL
Oxm88n9CW6Zn0fQqQUUp2o+BGZHmoOjATducrrjr2lHcJZBk0NOIvMjqJP1W8ndF
fTrHzBWa/hFKcwpUi3S8T37hZv08Tp9syXD1qs0lE4dG8/BqyKg97ITeW19NrWTa
KbBnK/XY+nON9MW2MNxCBJZeIlF0JGh9WrNnOI1N6lhZZ7EhYd8jEFvunbBBHbq7
1WZDXrNMH2aZuFGxqTjCmToqRypbEWHJRw3n2+ajOZxX3oCfe3+OAEY05aG3rKhR
2nq/MR9EtRPNWUgtnc9omjvqH1vBuouNEO/SaLKlmPdX83TpXvuw5roO5uv15U1E
jwDbD0pkdSOWAHtWNj2JrC2pU58KLELErV00X6jZ9B1IdT2HGPnphSfwjPZSjuFu
aE2ljjQh8BCfWVGQJcxaax4nLic373WWJ2Qsgv7IYD6rkXS4fgP0ytu2LNe+ezIF
ClMM2H/XPn8g1Vvg35u8pnkUnn6d06hb49ZclRRuGt2VvvGQLkTEpuEWkQmHexUG
9U2wPHHKrejrQRSW7ia/YQMoggF2tC5umDUV537lu/RpmrKfq0GsvhHTFUhorgRK
LIlyX7s28ea05COPq0Hp4lur5CnJ4Kmnwgi2F6EHI0q9TrJe6bGtg2s1BoIJcRM4
O70ArjdDKt7pBhwLPM4QYswS/4J6zgcAztAluweufDMjCbb10pMVzdEDJUSqIxSZ
C23va/54Jq0UEJgePVmtC7dL+oaIvvoASTt4td9eaPQ8LxSerN9HEY4TzrNs8aGp
pvBo4DyCrtEOwbNEdQ+gESeRRBrx7mTs7xmuzKi2JTWJsSD1+53XNGRmgNwk+ZQ5
RCZ5Yu97muMomeG9f5GSD27FrtP1Vh6LBJjjPMA7XBsqQKGvwYA69ezFGgI/zfBu
SssrCGXWxOY27G0ZBFyhOBxzPgerZy9jsIe8LBDI1aJlQARxFJar7Uxyj6so8/JM
IsYKT2u/zIC3i7uNvXgI9rp3LeU7yYdL4FRUoFiBC7eo8Nzr7wOb9sJ/NDNnaMoY
FEI3nN/MmtSASFBvr0BRgLfJ4lGc6Vord6uDK4X6fas3W07C4wQQ5bnSsKEQah0t
kgpeJWn2zMZMDcJ+tlFS3jy/n8V2C1WD+jt4iQPBT2vcm9yGYu4PYBpqQPkJiccl
SfDEAd2BDYHXdpPNy+KoqoGtWukzNMyKvCfMZCrh+bpygGv31yJ7p8hNJHq6BlOh
FFnOVx6fZTRaFbztr9AH5p3SXtmG3zpAj9LLG/MjKUWDwW9zyv01ghh2CJkUhAAm
xLafRXOuRFQ/PK7PrhB528YSwjtG6zXUOVqVXUTVdnxSvAXcnsxCr4ydIAEkjcGf
Ut1F6mtfOpeMSuT6SxLy6A4u3uVCtveAlXtB+U28AEBL8AhFDJMJm/qAF7i7VAkn
colj5FetuyA04ZeoUgzOwMxP5Aztf5tjUQGvGqO9ovEP5dKJsLn4DRp/qttTLSah
NHa4FFypdPcdpwH0rLIDHUOzriNdsIe5uKIMlEpK3gi4TnRmbPgWirJRHDN/PIzj
6p/tQFInzUMCT8zfI2t6t3j4EVPKIQHH+LgGFAF9yuymsVKfkzosS0NvQmPBsNph
K+NEgZaDh2RmDs6QwhS5sTznvXGQZEGgjh1ZMjQxGTY3TpdotLNW5qkAd60j55wG
HPMcozyiq7ON8ReFOrvgM/tFQ5CyyMBzn/jF6nJhAGvu8pxe23ItnbHLRjAJudJ7
+ukaeZx+Pu8aAnG59Z3JcU4FxLSUggfdIb+0wVRGXGU5oCMin3X7mv4WNHmlAkdO
5QSIf+SytC95ienKS3fgibafAdYISMOKMLEZGAuT7jJnlyViztKQCDGD2lNRHT6l
4cmLv6tNNR+fIAKu/QAu2Z5E/L5KTJQGDcmT0ZTIpV9dFf05zults2fg5oi1opHO
ggQg2sXaSrpWXRPZ/3e+kG26F40LxRfwLKA64m6amBGegyBuvjgr64cJuiTm+CH4
HhkH52G06AojFpevTW+E+CDAfGtfz05oDFGF+D18oQtpvI7N86eUslfIZCdwWRHd
3lIX/Nv4inxhsYO6H7cwZ03IzvvoeNCtITf/t5T8Ue3BK6lpptMiubGqHhew9dyB
cVLM+YJScv5wZJ7ZmjD8aqafMQQk4wrNhGtbzYck/ET5SQt7eGCMT0FtkZcIbx3I
w7e7aRJfCVkKu+hEZ84N/cMUB1BAM4z1pr+ar7HtEs2piTYFpJ2x7OESNUR3ZOBI
fMxra68/y51JaWlHXYkz8Alh3vaRY4dAULYnLQbULZUXqc6JupFnli3oM8lIwYLu
k2TwCuFCIHexLpTKkbxQ4fijgXgMYPqHuaizkSwo+10jlwiOQWjCJORlRXLNVVyA
Gl2xsL82VBsf6FFdUu8zq/If4nbUfqpb7engD4mWXjGQL5o7x6yHeYNaQmIwqe1/
SdfeCwSlktIMPGsYko9oXTmXzFXRU37R4d1WXHUt0YkWjju4e48A/DtRMdkmNcDk
EfqzPFKwCCoT4Hw4SbkXvNdI4KCvM4pbe/2iL0HEVarmeU2XECl3THcvRQGJqZFP
DPkYQVo/G1YnRe21CHtEQKgR9FkXVYFhw4GJ9rShmfKrPKEuoRct22l1QJaT+U2Y
gYnVBZjxCHumNvZ2vV6jH9VtYCVqwn+xBCHSQ8vQcKJyl/CfzWRCRVwBQRJyn+k5
yx2wihS8skZFzOAZ/RUDQe6tw4dN5/vGHSSCkme0kWapd2Axa3EanqNe9KUIYsc/
JQjMy+2orN0e6kGqslOTk7OQZqI2NVjNJBE+DNgmGkmzNvHbsjfYFhhv5w8lfCUa
I1W4ovyZ3nhTq4h+dCto0rgbFO0i36ym1lQA7umbvdTpwzPF2Sp0yZEuMAISjFn/
mcl8c6Tsx/Gf/Lv+UD1u8EX7WiwtDNmBv4j3FoFpB3Ha3dFCp6r4MniawBGajYxc
/bYdB6TBfc/lxW3ANA0gyJzaXbQtaad10sE3ocHHC7ty0YtgRue8w09azkk2eq/0
k3vnYiGZNBrG88bzsZuks3d+wEwu49/wJzVsO/CIBaAOdn2/x3fGMgMGmgEg2idP
1kz24yfF38gdYS6ZNYL9Qs+TFXah6dBRvTGVTbVBcQice1alE33uBgJQ4pqRv3wO
sGrRbPRg7DFtYn8vRC73oQwj4+aFaG/aqW/KprbquZqULRsjbtv4DLBbmQpMyY8o
P6YJFvdk6udfs17Byv8CIFCNbqvwUQzhh67a0Flz0t0O8rUOl+4gXAtG317YzhUc
CzjBAx1EZAiTpwcQKd7IVmVAs3V8UlM/CspZNaP3lJM9lW5sx5/9r1yZe05MFZp/
P7luDIdDTUwXN5plenyMyu4/EA1nEC1xcdUix9ovEE7sVAftHVHp9lPxxdEY/ocC
Tn4sCWIh8oL1PzjXtJWMmgcbwbH1fVLGH9Ldzb9AR2d/DZr1dCnxGWfROe/MU7DV
2aiAyZt0Wwe0rMrOTThrMVsLkYVaunAUwUfS8X77oHeVnaxwEGk4mFWFyT6ygEWD
ZhS8Twnrn9hVM8bAOf7HfUxs2TPLBZnqVnVFcjUDU7KlYtbMuLVphxk7fLGEsiJY
OSygk04VpFmz44zO0OytakHhuzxrw7RCpD29uPxQWgZtfyiYIk9QJEM0TtiuE0+u
l1I9ANU3LpY7JLWjdtu5+b0XjVjHd44AevGZdPc5XKDAi7p4oocmUAjJrC+cmIz3
3no7SxB9dFEzHT5A/eDPJAT1yssmFuKTG+hV13zxFb6h5FQB3YBMGjUzvO1sM0sd
47tfC9gk8Ywfhpb7nqTAjjUue/9nNmaMtlWE5NE5P5rlD4CSRKBoxoz7NtUHbp81
yxB6jUMzX3MjtcbSo1Ns7Mrr66H7YGfTeCxgClRmDJaz9VdBxNfjDkv+nK7u8gTi
KasfRHqwAz+KMSFzgETuImJylxIOkQFBwndDfzDVa0zJzuov3HuOgrONXhAxIKkA
M1QGfYo5q5iBva+10PM12FTfwBuL3RMWRUf8x/oG0/QnkeIb2vzsH/Q8W3MHUF2g
aPJCT6k9xL5CXS3tEktOsX3Djd271caMyjIaekxzXu8yiV7j1w3mavHkHis+sYhu
FuOCppzk7NB1Co7qfDqGyJnwG1IKdVEkiUeR5QnYtDOIC7Ypks7b3TAfyJweVM/O
jT331Lh7Zes3GUrWvoPVpBobS7230fYqPJgjbCxwN62O8VwpddotlNsXy/SD95u4
EUQPjkllHAP5YXeXVgYixzWDMva6QWNyfl/uwVkBhFtD/rNhvUHooBntK2UsB8jF
U0WjodET5vSUOxN5+vVDm2YyLNb3QvyKlOiy7Tggeohy4dwswHwkXaDwjtfBc4ES
WXE4ETWV+qVgVBk0OJMqBtGWjSzzXJIJ2yLiMQ4PQWbScwkzWf6VMpopkkN9MxYb
FEeiIge34YS9GTUUty0riJrOEL2HEOYrxWlRE68DQNlUtvPExQ5oAsddR1q/6W1g
SyjBlEHQZ+cxY0HPlVvV3CpKTb7VBHzky73k1ZBwjmeiR6vIk23N1I4mfNTvpv/h
GtfuleVOA1Bj6rcyfHMf0mSZusegBQvIyYq/GGOoeil6bbHpA0z8dxmdDthQM7FF
160YeNIa4gpVo8qYTPi8FBWxlb/hKIdRIRGwQLn8Z3DpGvGaG7zM2NygkfoO9Aui
CsmqcR92B9sT5Z5pNDujDAyLfHFSq5Cn/NX/xM9+cByk8LazpakwpppWbtSE1HNT
RJ/omZiJ8LathDFzt6dGW2dGbUB6mAfGPcu5QpAe4POCubAOCPJ/DPNEQxsjwlng
GL8L0rzMaf9AYyVmD6k2mA0jqYY+U5UPoRso31PVAlrGqgp4qSdnwyIw/Xg9A9aA
McgRFqhFapRTc3qfiNANObumDziav5NpDTEPajqdToDfYlxalEPwO1bcH+mdXrHR
7FdOFNMYXO4aS+buDnfwOZ5AKvpWlYecfD11K9ZbW/MzkaJGDtp3LJXTSFIr+oGZ
7C55rzGk/YVAJiw5bDCVjtfilR0TOqnnRS34E1jy18QT745oLkWtCoY0ExSwHThx
2bc70M3zB1KO9tI2DQ/gw7aAKr8dKvYUdhk2J6JBVPAvUgAfmAaXMMEw7mJ5c2xT
QDMjvLqmxuLeBqNm/dc+JFudHtnx8cEv/+b4Cp2JyzkHYPgmOHzTdhV/ZCMHtE/+
H4XtS14ll+wUE55ioaw7bD70k+ME4UzPz46I9XSJvhDlXSy17IDXsWTWlpG4xBTn
iiV5gYf7bNKL+QbXHDfeNj+7Js/qKqitHHOMnfHGvhSnSsmgDGPAbooLcpuTjZjj
M3xziPw4P4COoXZg1LvJsRFuawqt17DbCe3qGL7WEyiSVE2xsNb1sbOcfWt2qbYO
vDAnn2P5f6i5WuKqq67DwAkae+n+M3IATBPSM6j2ewrgnouBjhEeuNsqK93qpKqH
YALFIRVgKSOy2qKWSuwtInZWbymiFv2me5agkKB/q1T0TCdkkhkP9YWIZJ9ldpYO
eb7uGmJ3cdY9t+in7Bz7r9uVx3lbxC+jh9mZd2cjP20V0KY/RHCB6nwatcV6bFOM
kan0xovHLAcsvuR2q7Ras1MaxcwEralbAgt3j+t1MVeomCUH5IX4mAhtLVh/63nL
QJWuemsJh1/2suoNr0Pe+myp5BxeQWlWf0E5vHsma0KImP+QEeXSlH8Pf8G1vuA0
6v7Yo7laIuABR61g3LogrPh1eSB98ywFRK6MzJB8fhM4fvPFfHt1RCkmMXqWYkuu
n5NOoDRTIKNroll8ywncK4olNntyceLNaa4dVq9enJuiKZ/ZrSL+qH2P5f0RpCXx
mtyE+DFQmZC+rPFOHYlIgOQjK0SpmLRXBlqCpNZPITq8vxNtz7khiEVk3JRRrf9q
pcTJbRfq47jC0j1/9V1zXD629ghVPArOcjiV74504efzvds993pLcOapOjieP1cZ
jFP3DdtV27JMLbGGL0ekPhKOuA/zWfMN1Mv16jm/W8gmooFLfzPxRwIUrAZ2au2i
JNrpZ2c3C99DHFaalPm5VBdq76isuOEV6o2NJI0LH2KVbp6owvnabyiKmur0cEG9
DSWm5hasUhoQRlDVdYkRMZtGvDBtkHILT0wmumScg5er60UMojl0JfWuEmez0l7C
VOzpYloPsj5IuxsCx7ZK4JB58mAL+on12QYU5jJp45paaoODViCqWok8LfZx5SCV
zSVHBom1W0B+9ew2zQDUPAz65O+qrYyW4JRSZwCScgxF1S+oYMWmNMp52y6LUo5t
VnOhjEF45PzQbRoRdR73bP3ZJLy6meVM/1l7sIQZ5jEW+wlhJx77yT2kW/KGPup8
bErrhbxkIGYEXJyCgN8NihM9aVyQhAEPHU8ubSdbXlB0EN4iyG3ln9cIPvO4p719
+kPskqJnkJnmYjhCU3tHWtlcybd+MvPRm//xi3x54FYMMrc9hZDnlzlJSDaLkPZP
jG2zfTrxtuy0t2cpDkgOTRI6aKo820Ak+P1I2LelKt0OjOtKb6m15N7o1173YOD5
/1cCukoJwiZqq/dFf1j2Goc98fqf7LY3a0uuoPqvqTyThPU2ReknOBuy5M25AAsa
DNKf7rTBUUgP6e8TAPJOOMl/4gYHZreWCTU9bRVC5JpXGr7D2GXYompjqRCUSndS
av8T2qHLRiCzboWrT+bWBohqySe516VXQD/+4If4T/Wg/Z6V9i+tzn1mgPMdYPLn
qF4WRjPmAnNA0B79eNWXp/NysPqBcxkDLe+bpbTOQ3k6t/z5BVvMTOhg5JG2x7qZ
ZVUi6AvXzv0RAyNc6Fg6TY6Z7L5zn/1j60ylPDgoDWjWHorF8wX+GRjrtgDNgAo+
3aOUBMong6zdzSwJJvre74VmOIGrGo/G+HN+vMonaqFAhqvZUU/YPV0xRplYdjcY
FDUjWlIzqv/tYSGGMDIG0LqmJ9+qEmjnE12Xz2RwG2ZVoMLrPSwVsRpd78Jh9euO
DMk+QQXlazTFffv1LkGK+UVyYCKmMSdQwn/s4A11nymRufsu/B6Orgy+hOI/zOEw
YvwIy03LqEhYb3Xmewq0OvnoUdDnekwzqS8CbLDZltADDr1ezyly2OilZ2TfXVVW
sEm5QPi7l8d0VPb6k2Le36x7LDv7yb2YQ6FvXCmUmf7uuJe7haF6RR9I5qbDSI2n
0EmNU+FtdxgZGMdR0FNSaKGrW5qxZGZI5/N3PQazcLagnNXw1KgEDj/rDv3BgrLK
NWANdHMH3ncFMEBsNUs8YUR9l5b5gwr7Yu1jdBfsbPtkVHRtlPO9qZANGTqULGeK
RYoATsXLtPsNnFmKb8NVqTuV5Lanxs/HlFOggyUCqcOtC4BnJ224TOMF/zAR4MX0
UCxAF14/tqZfeXa1brO5sH+fJIM5o/+EoahMHctS+BCDg4esIFEqNwhfkk7pr2Xm
feFOdKuRGnyYlN/SaL+Kq27qBUMNIGW+Vq7f6ZycwBrYKI4E92Oy3qjmi74Yb+0i
1F39LwPJ4/47Hz1tZs02C2vvxRJbBU8oAr5uK8azv2e0oxtEROyzSWuKxGlW0vmZ
hq4ISxF6seQENiT+k+0HnoWd7D7szghjZaWBMtO8DyRG5fHL7OfBvuW9DLubZlmX
QsMJPvBLqAMvY/srm1Um0wnTdqtR9gctbQ/Y2yfCChN20w6ny/EaN7Z+SBubbHHM
Lluqh3l+jdvw91ohIXkARdc2snlRGACWwlsrqDecZD2Yo4CSrnBFC5aq825FayFZ
yyOHGU64GA84ynHXeU5iYF3fjgpT/n0S7j80wBoAFh5Izl6vTNsY5Cd+TaLjWGGs
cjptU77KnqDcSGLZ+MvttX8iHu12TydiC78qWHFDZdVFApsF9uLl1rIPf+YyzK4C
ZRpkfcuCZe5PMN+RVxPx28g7rNYUDfYAJEK6dfSc4vLRTr0lvvo6WkP+rYjEFnUW
9EX47UkxOa9rbRnMXW92q/UpWvA2EaN6ZtrwGmoieoYu/k9vtFZ6CkLwtpv19xB9
enQ9wv0QURcVT3SQ0XDacQUkzJQwJvUAKEBuEMB4Nsvheq6kRnKFaE6o24apu8sM
owXKX0o3ccDIi2lYDp9bEbLXQ3+gzWKJJd/ohHsOuf9+hdsEOlkEdgrsZHdoiENr
tQzAQ7nQ/6DKQaixDvTbBnO/OZ7mHO3Qe8TC+pZr12+x6XaT6COJK67IKCiWhmkQ
+EYgSZLP8kP7eW2cy2Zy0IG15l1BeJmoW92E6+Q1mvcPElGiR7a3Xn/Ofqp1/0EZ
gb/5rH+M78EW46+CBM7HVf4nvHfC6x8EFN6VpmWu4HKRc8VFdnxwhTwLz/2GJfqp
fG86JGU+S0kJFRWbTMgq4V56DVCznIsn1vCAX/4nVhcUv201QBQnlyQ96zb8sKTo
QCU5BmIVKsv16L1cKp5JqHNwU+yoWRQYyJupOyck43bbc0+w9Rii+Fifc8rl0ReW
TjtViz9AAmEBb4kSRxwV+ypR+CUM4j0MDdMU/nGHLEA7MxL5gR/+AotBiAGH7fYD
ZkKFCdI6sPZ2BvMMnHMceNv41be3NK44tbFLdTJB1JOED/5O0q2ggFqdV6jzLYHp
Enlk78V8ATQyY51p0DvVf2zaEd0jrf/iR78EeZYvrztzF2HVZ779eA1oMfa5/11D
gf2TpagZ6ud0G1jGRv9tmCdlpE/qIa5Q0BMzM6WJj6Wm0Rzfz1fVNYI6BJdBq/KG
zG9d4DdpARiuTxbhMp5o4aauwFyLbFQM4e3klUSJnd0Swo4DFLDSSKXVDOq8QrhC
UrVUc3Zmpdg+o75AmlXaOvth0mE8vA4E9+EHL7S9Id4fO1niN2IaAXL6Ql+YQEx3
Fkd4HO0ltSOGt/0Zki9zOs/7Rj7xCVVWwDS9gw4zuEvJFwD/hAV5apC0VHyxfNan
eQ9p9xdfKn+9HrAHIBRw762YPi/wDL+tj9issYcEzBpodWx5EnEUytl/lSde8HRB
R7IWtNPRKQD0cwyR0QGDl0QBFbnq0YatR1WOQKnLmYp7Ry5z3SV+t6+ZB5FOYF0w
NAnknCI0c8C/CBD/bCyKyIRGuyB16Sl8luKIArWtCY0yYO5YjvS0WOvWEWRUs1ey
5L5OrI5p6C49aD67c9UJMIMlmll7pysjattp2SxOp3+b7lzz39c4cxJX+bZvMGkM
nTSgLFOx9XXIeZR0x2TH9vB2UzY6iqeGEN4U5ZSq/H90Ur+ETBVvW7B1CvgeqzvW
lMbRWM97WewKWISvFlMynqqtivc41YO7HMaWcQbMqgW5rOwr5F61UaoSS4hebjyu
aB7HRlz5KGgdxFD+IQ01xhFjoI6VV/5AWq3Nf21iOhm7s6by3ij0SrbT1RglRZgv
e1Ro6KejUVPQagTmNVj9F3LsDVVaN7AUriQSqb97hdtbiFNmuEbU9DmXADD/wI/a
o2rg4YNENdO3OU088ix7hcsxhBx+NGynlKhmGeoOogp2JgPDuIKcv95M4zrz5+93
eNXVBTwSX6dJEs4u41eEUTQkZTJMi2n4fk6KgE5F7gy8Q023hkrWcvuR1DTufa/j
YMEW2hAM6HhfBQuX1maMUSMpKRD7pdmdefG1TeiV53UUPq8fwZ8sW0DXpNUVoOi9
iafkkrdcNif3zw7ZZnPDIqA0FHDiKl97+lWp/CdcqhZmEEjJnDZVC5thxOKQgDTg
J/Jevsnp88NmLa4j/kr7ESMuWYge9EeSgvuQBcO3DTdibeXe2RYvu+x9+kHJTiLR
Nb4EfYZhFd4KVj5elax0z9WKzmuMToLvBT6qNxjUU5YAna0spPZwQ0be5xDFf2RE
mb8McqWHqGt6Lx7AmLa6N4cmyLkbQeIfywDE7LdbgjgAbS9RtpJP5xbHn7owKWdF
xt2C8E5Ykx/OAovTJoe+7HycFxHPZnjHcdgGkzAt8/64PI9fDSdYXzIwchdjAioD
+5J7tH1HLk2IDmGLar26z3sMh7LXi8pmXP3tk4w1NklMiMNxGcaGr5MARKFBMqir
6X61QI53M3HpkOIhKFSAkqep5T0CHugVHokV+O4ilDeGHAMgTd6hvBsHkhGc8UB0
D9yyRIy3EfBzMEGFwqZZ6igvlWM1XAbVmtA3Xq0Ow7/lcpggACxJ8WsN6jSRXTzO
kbWl9QBFk7YHnXy5hmAEzqjj7xjD1q1jh+c337WVBWjdQoVZ/3d9HH1XRkiIXxDX
Mtse2bYI7Kd6yPYF1eYxqWE7UiuDDj37fhLZM1GjyHNbnQRFqB4P4DJU5Kwt3XT3
d9OP8jumu9mV2BpqbXzbKXZ4tLrA1Gqsj0idei2mSLvyQuYIEQyYYiFzPCbpXxwH
3VaA0uRM+btkLPmS152t2jDIXeWI28qxOr6pF16S/gtVtMFAt2Bvr7/mdVz7PlVD
99QrvHX11QZ5Nf6xl/btrRWr+DnVkedOhbQbtrwrGQE85uIzhsRDdklvB1pgrhH/
x+ECT2awNvWTbP563j259zNVk4gYQwZ9Z5H8P2/YADlmdJrmKB8ARk51fXh7izsU
d0zatnbRDqU2TPVJpe1qHnApEMKBZTnCYkII3jeetdZBOohC7rR0P8xg7w5zwEfH
jwSCj4VeQN/xLspoE2ZXaLn1rN1J/Q41aNdS1TwDR820T1idF5sIiba8VtzoBZyi
AwWGuAb+lsqdLwGVDZ4ta5exSS3sl8Y0Uxz9FcLo26f4svVxSCDvAUgmikh+D3/d
Bl+jyUmIQpi5eofFe2PNtC7GXSD/Sv2T0TW4rSd/DgJdvQ44oeeORoOtyDL4SkXK
kVodT/ec1R+QAXTDCbDNnQcZ3bRaRhhzlIrFz7o+LJ32BFNTdm1tPL5UV5yZcazT
5/PuzYedb1AkpzZN0/36/xjUQmsVI6QCj0f/gZZKE5GTvPNrsTwNHqN5AGVzpM2l
gJbkzw48Mug5+hE4k4f2DA+y7aNgXc3jHcSa4CyS0lC4NK5DN4NE6TWqYYTk1f2S
yYCIGRZK+qanEX5FHX8bKXdVS43bKr7woTcKee8fszIYCAvdNQyurX/RgAd2Ld70
LgeKAwxnxguZfOQq2LvMkttHPyJkgwOPIKNtKx9Ah+//wl3bN2T//dqsHQkNqzSr
We3GVFLZlzQELaEBH/f6nVF9rQxWjD3egwDyCgsIqM+LVg8P2CfJfSowwlc5Qm54
QC3jpIrgM7XqJABZCILSr1Ea2l7eIIc+3Wjmxwzp02ODTUTatcnMnar6BH70eP7J
BjV+GQakR74n1IhPJ7oeqVKv+1IG8sjSLNXYE3FtjUZJZEhSX8EeHHLNOTbVpLtA
6VUPNiNxzMQhsL+CIBad/pdWrgn2ZntA9vpejhn1SGlwMM/pbHdyRfI6QLfnnVjB
+r2aG/QRRVFjR47fZKetxSt6vNOsPq4OojdNcuuT1FgQFrVGtziK+aBa4KTg6bW7
Ucrt1b1xEE8UvOPXeMQltovmNE8NGZrCF3q6iy5CqPkvX1zlQhcaUbsnV5WzxMUT
CBqZH7UJknpikXxI6kfwHl7Jwn0r4agtzWPBNTR2wx0QBAkT3wU+Fa5xCA2JresE
Pl6DIb5NDZIm/K8uB4DsFWObhihwEC7BK6qflZBFjGvia+AiiSXA2Nz7a7ak7ymp
Yy7mHX80nNjwFMWimLRbyuPOkF8EkOMyqOfQ1DOHrRAq3JypYTitP9qh7lve5NcJ
aZxNz3ItpVinK3E/RpnxJZAvkJ2haRYkLP5rU8/n68RutyZgTOTr1vao0gCtrICh
q3At0S8o4tI3ldMOQZWNi7YuzgSapWiUH6oMvKaF02gI5MO/Us/e1h/sMECXaE1I
qXhC4hYjc+BYB3AqwPf8QO9hOq6QSrtQMjimSOxlzjZGomajAQVyM9Er7QslZiHv
wKPoibS6ABHUrWhNNVBMTMBZfsYQD+Z9KX6oTIVqS9UkCeXlkX+7EPI++3tOCvoo
XK8StyRC1Xw338PQ5KVPHf5yGGXdxZXCxpEgCB9Tihp2U2yKwSNj4QWPpOuXzJT4
afuoQwESo4oLT97wua/UarGaa7vmfMMw+AianXjRDa4tyynzY6ibE5MgOwWXy/Qn
0DsAzwU9RHAE7XsmL/T0Oyg2E0lHlv5v2cAO+Bv6Cfl56YF9SoJHWQbdtwxGZTaG
ld3+VGKudh1W+lwmxGdiOa3y3WZ/l9tu2XXbkwEuyLPQOfskOU+IDnnt917QZwZP
YKxKrYqLakSxb4ULpwCmzUZUHLn3OZWLeYStPxM3ucghh+k2oDxtA4qHWTDxhPLg
R6kF0AzBk/j9NiwMyRd6vBsYebk5yh7jidb9W4udJLFWjqclsAlwrmkmJTA/TcpR
j4yIh8HDOS6LsIQGnNQkygjezQ8f/GWYw+IkKwyeWB0jnyAzSR9V+3Q+EgkQnU+j
up61R/Ngj63EysuuJ0ViESD3I0kHfNfx9dE8HwwdPvW5uvZVZO08tsPFl4r2TSmd
+BWxTmBlKjzyZqUNmww0o5ynLWuiJxM/qeYGjrBv7rp0AWGvQIzCA+Pfz1BKxpLd
JYCe5cXb1jjz+CyBUORlHXap7VzwALuKAYDIvfu/tuy2VQfg6+QQq7fbcPikPCRR
cLR19T0wp+vfrN8UIAt0oEQMSoXHTgiHPLaxU4ieAILi1PMauHWlGTldUqtd4v5V
Yg5ZxBUTC8XZBxW+INpUKKKbSNm6Zn6pxVWcuKuB4sDb0xGmott3RAmBuLXxhTnk
Yymtkfy2/Hje0EJsx3OWL+Ml/7QLaBugR5zgRiSSYpFaPnjDwvXp03GWxqxZElA5
tlqvICsyaWGtuoPpis63OE4lYKiJSDVoZeN3ic3K7zXn090tmSEFFNcDClR4HnyV
sEJfxbUBEG7rm/9uIAPbLpCwjHm3o+XA0zp8DzFwGpbRldSF+Os97IR1yZewBrFy
ATXPF4Ez9zo2sYeo11d2G2ygS/xQ+6NQLz4sdL9PfSoas2/kJt9j2XMjX7JUCnsT
c4spkbE/rrbd/Fxb9Oa8JAxGMNiFNMOkB6w+EfHFxaipDPV9fJkgxEBtFGxMyemW
XwaqlSqU9nn9wczB7HpHhbFZmWWvlpSciQkraJGABhaoHY+qsaU3d1t8PJoFeVPQ
42aEBosE2t2QRcvsAoIcd9bvLil8zaFY4LLqpWXaW+wdCGbp822ldzSv6LyO5ODo
e+3BDMudP9OzCrL1pEIPF9GdJqfwyU1DXROLSqh8cDpBS1T94bb0FBD7oTWzdOcD
hOE3ScP31x1Covzx8Zzf0VFx3rMKviyjs5u5rtj2WXJb3Y/0DsiTeBPcTtPqaTVz
rrxwPz3cjCFknMNmc16/Bnphe4AGxsJ5M6xp7uzyjwq7OdeVv5Dffico1lZtjyKV
ci3+n1mB8UzKhtwXvuoutzMciYMWqyl8MSPWSEgW+1w6MMJzu8XGLjH+cNWcqB34
eBbWuTHc9W0n9zUDcKlv/9PbiwDA9gegJHJQDrNNBLhEnf2sSJWz85/KjLH7biBp
EPvxG1yjrI+kxpSG9/YB2NTPYRdVBIurizv+IF4yw7q0F1AU5yYscM/NG86GjD75
MwDwtp/x29ZDbbWa/jXeGZo/VTG6Wy33KeiqUBxdomQkK+Z67iVNXEvVUV0LRvOi
V+UsbGQmpxIRi63+jRHrEfAnyGVk+nEm6DOgKUi1iv78jTa3373BSm50re8V/CCE
h73K/ikTZxnZ/RpiLJMHP5Mgq5s2yJnk9Czabm0AQffsANf3ronKX3rtCrS36hV2
u0gMLWPzLOfV/lkQzuMMMARKJfC4A5hgBBt/e/yNMt9g9Z6WsEbYih3cAKyIndKk
FN7+gZbaArDp4zGYIhoQhGU24R3bf3eyNBnOUHQNnu5sd+eyw/OrhzuxapVTcCPd
jbQVJKO18TLJVJenyiBhVVsqJG3TGMwRK5y/A+CP8C8u00nv2KRWhC0vLuMkYL7j
XnECgLC1Ffgv0UWJm+BzIuFXftd3lCwKd6BttNFIeUPJiqoZRCVYanyvCqGnqpRC
Kc7H/mso5iEcn2zrHkYIsZt2jdyM7+bvx12SfQIaE4P8/eACatAL6h7QJ6a7R8S6
S5WDshXhncyab1Ba8j0W60pYQ8D6TVAzYOWL5vteUvYU3Q8smFKpmN2EUFvcbWDe
DN7S93b8DMnHR74fgw1vvFv5xclOYfA7Erry2IrjfK7Hf0Jsd1JsovtCX/rWubus
0CxtHjx+xetNrzspN9ljkfsGnxhc+j0mjRA+lIcuMhxniJXLkWnz/179COKmn41d
aPQ8P8/NPkgYSGhSRPCnixUamhcODcFLjIWXma4MW2ZqJ6gWVeuMVz2u5mdOStMH
MjlwbXnm+ox+Xj1RjvQdJYUaF4ls049KI4lgEZPx91eDfPK7H0E+HtmqWdjqj7kJ
NlO0pR9+jRyesOP8S1NgSER1jGVziQME+KSrgQcHfG66bTIayj6Y4rmfbazWdpb3
4LByuksu+zPAGHW5wV23oz8AOvazaBmXlQc3MaCJ5ahg6tga0Pude/n9MhHZakxD
GSEne84btR5pVqxki1pz/k7ArID2TabkQwPfpHdGGNY/xfYZnOx+4S32IizFUDZv
ZfXIG+iUNUG+H2B6GAIfTCMa9kpEuUfies4OdPsfJOnalJ5AWA8OpgHUFrVSzKv3
OAZmxQ9LXBjPLD5iIgt+QwqrNgiJCE95hxIvrSmnLxeQYmAkORLFJW4awZGhZjPU
nzzNr0CN/nzCzV+GiF12xcdLGsr0FTJzoBLKWiZv+Vsg5Tn5pfenKXFE2umu0ke1
6fz+MRWrtccYYYLcg9/m7+uczAYt8HTACGz956P6ssdttjRRAAw5BhsQt+seIRxv
UssiqMIA3qUZokojWvJ7VNqV/T/ggynKKpqrFQnoP2YEX7d53BacMpRw7lwv6O1m
LpoYkNw2h+scV+qILaVdIqyXYsSejkIf+dDPmw3Al/0U/GvnAKCRvupmzVArt/vL
+chAJkuKmlNdl0q3fpWavLZyyhx6eykC/Lk1PY/W46ev1vOw7uezYpXC0DxXalc8
NMe3nIx9OzX9y9YxiHAFuYMYvwMII/4a+EnmSSas4VggY3XB1RJGeS1fCsIOpCQb
1kUH3Goqe0mU36VJ76nHu2zdl7WnP81/c6kdKTwwIELNb7nF1LGGUgs23s2dIsPC
U/q6gG4yoIP5ouQIitkt48437Ia43+7q8QR2BjbVBRfQKe2iH9slMyNMShDIrAj1
UaVqq+6gEt7Lff/4iB6WASmn3xAcj0hBQ7SCSYVTh6PCGmIW+7JCNdm5ZTuqHXLz
AbztrorLeXeTwqgNh5gHvUAQa4E1uhu8I41uU7c9+Xv3Ocmh46jU7eRbAqlpNJvt
JY36qKoEV4a+B8FKXcJ99IdyL1lRPKaU9tPqKIdDJ4xah2MSVI7xs21Xt89i/Xa2
dvoWwxdM0peJSUltWdKHZjtYQcE8RDP6Jfzc4PHOHjA49MsasTkTMCn55b3o8+d4
OU5c9HgQ3A7hDeICsTEjTTwpPKLoAH6zz3XjxZpldYEGaq8JON1IPzv0e5uHv7Lm
BxFsWm4TmMQdYTGwGGv062ys5XVXlcchppksr1Nj1nXxCmrTKZTHc9NrNI23KJEx
yLBczPZgLNeVj0CrjXYzv8DvRPfyhxUuwft1TESClI4tat7odD1+Q3+wW/Gu24s0
0CUlFCgaFUGuexxDSnrSlRSxVWkercV4o4suTC2koP7nUj2NjRQp1i/BWwSWrQRI
wyOrOFDklvTY/ssUsA25WLMVGWAszlfj0UTp/DGrRJ4TC/g5whE5gQJrtBLfOPzE
eOAichWt8GMY43ZcT8IFEPRmeyUm7HwPp0V09whAnMSKptWT4NYPORO0Kt1tStBq
/Qjrx2JwiPWwigVKHcvwcmmFhFqJpjYV3OLERUXeaWPH+ambORrtLwisAAmXm5f+
sjRpRC0lHKLB0mmWy3repmLDYfaod94vXwolbw0WXGJiWb3lx0LCnk5GdXSPSLJl
+B9AR+J4b/j5H4noo5D3flJX1yYjBIm7sUqkqL69y0OCO6uQL+uYIpB6z7Vuovid
1oeUb4liot6ZTmowrXu7g4ztuxZstG0eTB3RcThxFn7G4IH2U8BCAWiqD7RZyUlp
oLUCqoweVDCdK1No4YawlzyBhFtdCTiKrLOOA4vU1GOQk2QzuTuxkBS3xj+bIna+
+aUjD8wSfc+jHnsIUZuO2t3sErTSIDm9V5zWYmN8WoijWEdiLdDswUE1AMB1PpAE
axHwyGbtXRiLzwqm2BOXW+DCoG8BfZqsHm5+dfbbl/Hf2Y7KJ2b76q4gW2LXdvvF
9M6X1BsXZz1fkVyD0hwOWdKnT1pQtFu++vsub/UritmrqBV9iG+zdPpQ33p8k+Vh
uk5b+0jX7z7QbP7Lj1y8dM9Z4Av0qKbxYNCbVzn2jTqoSA9vWQl5GGt3ru2I1fBd
U0Gbm8o2Nu3vfRoaRDKy8OHns8T1QaxxalaMDdUIwTA09kpwrFQH4zpnBLC7JKbR
sqrCjBlBhYlmwdqGugodR1g0nqEUoAbQfH4fnHQdspzCuNEY5MQi9SDxg01TfWaw
4tmV3YG0t+QoXiYhonrNLm0uoNubh4qvQCHrlERHts2xwKLN9Us77L7OOjKEu9Wt
Eu5osrdBtec7Ae3AlRzBtM9rUibQCBVHTG7tUmTMutI3DP2YdLxvIiYtj+PO8bPr
YhB+KiqOPLcaoYXNPd/H2x0QBRnQLFvI04ad5cmzbjhfoJ1t6AEyTtLoO/qffbLc
43BGIUrz0T8EywRgpbbAddfH/6C6kjtiFanmtNgdXuXzfpfKfNH9F1ZUYXj/1cD1
qHH7mS4Z/q5mb+JFnkQNv0tardFQRCmEr336uTwtLlPrxTjZnoYtB3OvHNAVElxW
fAH2Z0HpEa0CRnsaYTfjqEqWAztGZGKXBrr9jOMwsAQcE23xy4xlZgeAYFEyGz3H
iBszwl0jjY+mlXxlIZNL92+y+ZG7wSRR/nn77yw2r+0vnTWmzf/ZcGIOQVQmFI3b
0k2Cj0hxzfzAY0v+grz6Oh6Z1kBBqfWxj3WhKMW23pE2yfNVTFMojqd9/w/O9dpW
fCig+1Abavj5/qucJrsDetU5tv+L33jll8fnz0/WftBGn47j6tWIrM2jb9fZrkcD
KTou0p5/iEUWI7sAfcA81o9aP+O1V+pV1bcCCZUoabA+r2hTnD1x1XYvCMZprpds
LRJtQ2B6E5lz1WdUnSxiizawt9bS4Js5iSX2Fg7oWnQrstji7cWuQYjVcxnaztvA
Kzz3riA0PEzzigpcvtpAtoCkHOufFRL9keUitHgJcjx/tfJdTfaDr8jqDUH0tp6g
ByMsEtI2mE8nxHBa5gfpQdObHNvPWIRyYVNyOvt01uaZtDJp3/SQlk7X2U0Br5AN
SToMLJRLw9LCqEIkvK9AtmtrS2ar6EAIelhmyFGoT1YXbm5X97rC1hi6ml1Jh8NQ
nyMH7Lzb+3ICVbejdOWEXdDPzeE2lsUePbl461ZL9+TwNziLo+8GXaaUbsxBTpys
KGMiICOkQ+Vqff7oTGV6sDHNnvQoV1FZXfc/JejbthNnZAYKLlRRZCT3KcN/PAwE
2TBvOat6egbzIBCkGkYu6Hr+1+NyCB6YCs8rf+AJ/ASdrRxEf9yhea5+JjebeXZ/
sraZkxovYSUIZ+N9K16pTLc4faiCI4qn2iv8HJRiSKfCWcP/IWp0Pe1ZEaO8Y0jR
x8geSxGWPS1E89UDWJo8lYg6bS17hpFtj14831FJOmYcQQPdHWxxpF97ZFuXv7D5
IWSKWKUzQWWR7hlcz4O1sP9Qy7+7s2Osy9xhGiO46pKm8LXGD6UICuWc2COIJ62n
l0c2dG93o4y+sMOMZhrSQT5xBiSSItiHa1+qJhcBYNH/gaCk2XQrzAR8EmhPpZv/
XwNL4GVzUpTORZR90ZsZQGxShsRXf5jtfFKL+svtOs/yNF4MZKsebh6VNX1LyeVr
prOJJDDGwEniu62v2mTJnH/W9HpLILYprKqK+le0FBGur+ce6ZgFYOLIVUcaMTVv
2sAUUzEOPRUPCJCs2sey+9JDhIZ9oIeZ8uYVwS5+gmdKxMe/zV43R2EuBykVA5cP
djca6uC+UCUoCRa6an43SYE+JY5o6H3ef/HFtohKKXFdLXbyF4ZHKE3Cu5Lt8nCg
hEg8Hbw+5C4D2cRskKVpkbQy+vx9Dh2OmfJ9HmL9K+GoFVJJDKqtkrVtzsWwWfzL
VcwQkFpaMy9XKQqUdM56hb1NpeVjDFDBBNvs1JBZLSbB5//aJPlll5ULACRQ2ehh
mpWKQYSa4rlNb6RRkRsO19LjrtDtVEHrM4haaZr0YTiJl9zxvhtAhgxdAlAVYka7
vAXy3JhrYBM3X/akzEyYUED2gaYBgddz+SbhRecYZK858Ib1T7x+LqfXi2roEAuR
4ovAgLLLkfidMWqybB7pSfQIsxtmS7lBE5dSfXbq7/WRGpX/61xKNVyPp5cMy8nr
8+3XcqbHC5wX+9vhSscI6hkYn8d3pqaF3npmudfppilm8c1BABZ/oHRKHlockYYJ
wJMvR6h5ejc3mUy694EOM2msiO4q1SrRjG0XD7tDa86mfZ/pd03VKo5XsfyyYQQ1
iNLOfN1wvgWnyEBD0rxlKU4edOUGT4ObmeVC1bMAPtH7lW76ZPlAqJ2aLvrOu9eS
PYV468K8AuPIZifs/Nbejy0AGdrGU289LgoX+ZhbXGURsncen4hBv1W/COq7KyEC
DJlIsKtgOAioig0jPsNs3D+S2PklEuvQFyI9t1u2UnEuekNhgZNvyKuqt3wvTen9
s74HBof+ShMboUW6cwN4RLEMOp0WnYTOmPWOxestQ0c35oMjPRv5XzD7WKMvsBpz
5GuZv6Api7joByObdBzyZVpoR1zAg1UlCBoqc+SylTPGFk+cuW9K82CrF0d6iadW
b1MmadV6G3sa03B2sfA5D6D/dxn7l/tzcIQpAGV+BaH/08+ht5XOHf2XXKJfw18b
JMFKzt7nSIRUdup+ZS4AgFwRHJtjLf/80RMV+FMPops6FPhBOPPjKCPpd2O2VszD
0ChVSCkGZCv8Ya4bCGLnjIKz9tz8WfwRqjzyBkoIHGtbuKi16XYNc3NHskx/TK6V
v9aVt5XJE4S84YgTpqqymMnE1qdbllUabUCYUs12nzRlazR2l5SqQChqibARmrpW
PEu8Ks0SxkIxiyBWX9aoJNUuHKo3TJv06AIocYVOeWO1y+Pzv2y8X82e0yzax/AL
gxscpQ6IdF+gAgAx791hLmvNg6ln7UxuDQBoYje4WYN7Xtf3Hxp6pkm/ttX19W/u
SUurmARqr8u7WGm0DvrRrh5wdsAgIMFik0eB/ubYH8RgZc1pIvyt1xzHaxRVrH70
Sf7IRBeUE2VUUKrSmONsShMJELKyO8/cne5nMAoJiBMQyc8g8yM53BE2/GPyk7sF
zy3wpIW4luiEhZOarWbNIDc5p319DKPwpJVEw0IyhonIpKRh6YoFG+ELp70DuPZg
S/A3sZMGEM7/QH56fiVBX5YRExA8wC+vrWBblJBcatlC7o/+wsDqmxcwylHZUm6i
AVlIXqlHXB+bz5tWtMK02DVhwXoqiVAp70KJnWk8Sprc7SWCwc/BVsZbthbnNYn7
62VgcVQ3AvcocHw1VH7S0s/FyG+RZmy12e8D5dBtO7jeyOYBThEO/44pJ8It1vCM
DNdxg5wb3VLdm2j4+7Eqi+7f1eb+R8JUh7CB3GoTMaNvpJ1rXH2bJAh13L0QI7wC
c2UC1XJqgjRYvdkBgcuWg11ho06oZxQRiXI3rHRWmJnEMvn/vSm+ruS5xP/3tO+T
TMyFPf0bDHGUNUbTU8r5VocLe8iXxULYBP9BEeMkoRsOQK1GJK8FgPNyffaHswJn
oqbCCdwUo6I2pqtMgzEKpxiX9zfQP22wc5GXuy3K314RJ1dxC5aEfDv94vSBkmtb
3UmdGg8R33uNrUePy0dY18PCNPBn+4n1dExwBQSXvFaIGfBkgwh19UlMFpEjDnAi
u3VD/GDhUbWFq1IYbKCfKWri/BqHkqnWAjIqWM9pO5iVO8vDhWbBgJui0Sp7IPXM
3wE73kcmrrmJSOV0ydH/9lxVItnnPvY39tFDCDuLnDLpIpJotSpcNx6NIq5ghTyr
RfSqYfG9t0v2hxpzYZvr5Q77uwA1FjgfGdCZs+QUz2O1sU5JVAKYnbYkY99O5bIx
pC9/Z8U1CdWsXWzwciKXRP9Nr8j4R5Qo6HGKckHNfF1RmnKz1V1RQ9rjgeNPLLAS
5W5xXBElkfr/fuMk9MaSH9/jEfm8PsXxe2SfucA+50eko8PXw3sGel7NjQ1oQT1f
4iwyzbGtuaoksSW/Qj7l895C48dc+igtV+eGYvvmwze16EeHcm/kNCEtSvb6AD5G
rVJCxFyPH5ymuhwwcGJGTDVp63uHW3+I09wuoOQqvM3bsGri6OCELAZ7PLeQEcbQ
HtMXJN28CtwnHDAxJATgNMGsRtPdIKTw348p4RSkkh1hiRFBfbmdlBri0qUxMF5P
l96s1PfPXyc9FM1AKX8NWA+emqIbdMEbYlRvE7v3W3KDr3fIPGM4SQ2aJSJXc5fP
TkKoPuKyC65x0KGgEU3OKJB8B1432tIR0RcLk38caxY+yBED5ME6R2aawSw2N5na
EPlQS7x+WmjJ+GEf+h7t5i4A7buWQvjiHNK1jvFaUurGmJKRlQhRWn6mhcr1s9Xr
Di+aHvi+RO7/ED4Yu2dN/wvlsMUdfDhOcNL+0jXJV2X5VIDv9tbo+ca8uorGNgF3
loV7oVOE2QttPxzuwh0IVfkihLK8z2E+7n3DRnqAuT3HPHs3DKWB3COq9H10chA3
VO+I/B/rTgMAYaq4C+zf33EuBOTg0ihaHWPyyo8/LYqMZ0f6b6+XYjoSkM77bZrq
jxefpyBON+wZVSyCKODN/YYZhjByIU620/X0BllNLhQVoa7+BOWau+vUXnOKwpF9
OkBZdFvSyDHK7JH5FeLRpEaTzggfgcAvfPKoHDCNxkv38r/ob9nU6xGRh5R+lELf
hGLF8RwCgq5pPckVI0m07hUdch3fmluRBQfmFTbNjLOqtwRjLk99ELTbq1+vEgVa
FIKfgMnMO68gN4oJtTM26OgKS+fxsV4Glt1iYDzLVKE39pciPwp7mQ7m2rrLlJJF
RDJ7ehNzHDVIgBoxGxsHmIkId50r7o4W+RyRr3ogzwZ4+ZIkpVw4fLIwLmbtrZ5D
1+EJNhcEgFko3M+XSd8gjk+fWBedcGBltn6KMP8P2sNx8TJvYw5lvRtZbO+YlNTj
FKH9baMJ2YUKdl26dBYMt1CRQHwzuI1KcDh6JGx0ZYxYqNfnxEsblVQf7tHor0HG
YL+oqz9CKFDdgAaziIODouLRiN/WZXCSUs4PhWgy/skWDdAQGqg30lu54aYEiNC7
gLMRBvjrakTfDab8vlTMci3zIwhJcMtV70iiUhOOdJgnJJ5JRiP3AE1847lc7cml
qmlSlTSU7ukJQIDlzooqU47+UYd8jd7iZiyKPuVb6x09xe7sC7eJ6flQo1VUK+AG
ZYPTCv0zvdSw90tho0F0bdHjziwmy4i4xN/Fw9M18biMHGseFzPPM3Lj6EBi3WrF
+lYJa42RtfYWN/ev4dVboq+/RbLvOaETMA51DZrRUKW65lMzFbreTyG4S/T9VZ2w
3jI1XVAnwNrtInfrSOKTfQ2m+r/EN1UA9ztq0STR1oXKLj0SlldUV8LsUm58PkKI
8mo1a5IW5PHukJoYa7urs4QQMGxWysgsOZoE9aBFVq9P0uHrCumOyoUdZCbKaWP/
3lV8GhMdwjZTujV36SJ9Eb8yEb5kfAKoP8/xxTxq6dk4nC25q/41rhx9a0jq1E4v
rM9LnmhOyT2V6Gn7aP+BTHL9a9W/j4y0d1zZ8BZF/4E/kyRRHpWg+Cd1+Ku+YHrT
4KBj/jCPyoumQIjjm8p50yxmydLpGbHzfnUwHvhkCoVXiG1PwsXupgDp2IjUOaFu
FlFlvTlG45p0DvZgFh4buUgx8SBhTKmh6Pm01YHBCQfXauRgbyh7cnkwLBsf9usl
dwyUzpJyEYgRWizHNf3oLWxY5pDwUwqDPqFqAS7ntxIqf+DYE0+NysLELztUBmcQ
DdgOieZFPDFRm9HxApsJSOuShrQ26LUkJ/ronYkLQjGa+BwS01rT/+usd2R5ejHM
Zxb9BBLK3w5cWi+ITFfUib+Lmyi69bUtNXWXyQZwtQkbKIfjygiUJrWMDsijB9Wy
AQu0qlh3QkZ1WJNjzreS/Mw3r/dN7WCSW9ovt7h33YDmeMCuuOXdO9dppRg0v6pe
FbWZkw06axYT4D6qATdroerUUdFU4aXqtiVuLRgBlBnUVkq9onSq6Agi+ALOb6c+
RqfX7YV0tG86kF/798f6RJJmq+O7aM9o1jZxbR9eN9dQhkrRNu4u4K8XoiE0BhJV
vA3PGRSf6EtCtcere/CgbbpTKSdBfTcUm8IvrFF8nEZomkQKI0sdDdI/b+CSGBFu
I17OPCUlWU8i0cVTDl7l11+ic3AZFixXpiDUJ5z5jzn+mLa/GkRuMSNJYVAIdcaM
nm/0hoFJd7u2mvRPv+xk32pgw2lUEsNYTCwvgr2cYgNkRg+8CfEj+kd3ULZO7p9a
c4fKfFN4ay4aEW5aCM1F+V6IqPZuzbjbkDXWD+PxNAbKgoyof2QfC+H4az+FWrLL
k6dqmQLJUfHf2CYpywmIXWJk4AuNDqrM+XFJVU2fpLYnnNw1z73duqYTVHjG3/VV
LBGAoFUZuKSy4g5V7URTnun628kjYMqdsk1Zgsc56h2sSdv+MMoMMJNyGLSHJ7QN
rW8yQrgYQqY49e9FJY9hVCD96sfXNr8T/UbGQIiokUA6CvqdXINmeQWMWLAEO0CU
7G2YVbXLKUjrdmb9HmAA7eoI5oRlEJW3M7bJKrUW7EiftdkHQIR0MQXEwGw7bPGc
873vyArTB5Nbsm0AkYVW8a013eUHkw2q7lbGqYA2KwT6ZOaQp+GT0GH1eZvHps9O
x5sFwYA/IF4FxKn4Uupx6O76qDR4Cj0s3a+XhpZFp6tUdZt+1BkqgFlXi1beaTol
0EUeYjhOBNT6MkPr7AE8Jk44eLQ74CcTWBd65Ro+Pc9R25SxvBNhwrLJV+cgyzv7
6ryYkvSbAdnpRssR4MGpivSwd/xyLZ+HmQpmpq5jh9GdXecVYUp+PR64LrxRKwED
dU64KwvDJ6NfWNkxn8mZrZF03nPpj8LJxpEASkCAGqtivUNmNBPwtGWYQFCNwXs6
5yiFzSOQ76/iM1plP1nifVIFxQN0qU9mLT/EIgETdXacO8DXK5d5XARYL4XNC0Go
GUFd9bYYh7XfVntTkX3wyQQWTgUTIGkfz7OpPVR9lzMinK09NsFr90FmZfskSrEw
76atqayBrtV4Z8JLChUpeBWIDa6jY0wEhki9/WWIAtMK8Flv3VlKIChdF58hkzDr
VvQ6Du8h/Jg8BQf1t6BzoP7MTBiROzvcSghYHv4Np2DT36UI1uRic0kQcJinVL4A
asJi/ggCA/i8xYrs3nULVc+x4bpnLaqzKrDxsGy4F7npMA4gfHMLAGeJeeKzcVgF
6UB0PTBnytIFdrmYCVuMSsXpGhvUkfcFidrFAzHw73EgYgPfDThpChJ55L+LOi08
MxJ2zLIka/3qA8HQ+Ml2OR+wSSMYu4Gc8UY7FuhyWsmJ5gmVONiNLL/ABR/54SDs
vAAfMmKZtj0cM+Z7o1wJ+QH1RFZg+N47xvx6uUaPImXhbyUpkI22fma+4GYCEVvm
H5jy+2YyBYmOVAp0UYa3QfUeXYgtbXSBAaSKoEGYmNtO5T5Q1PXJ/fiiG6GIabnz
QjQ01HPAFHBDxf08bDtSnOEi8zIIJHajypbtItwsLdaI9qqbx9nksUhL69/h2YsO
bwNWaIfj7PkfN4S8UdL0x8DzCoE9xYdaL1f5yTAhwt0H8x2KAliiAj1N6kGY4/2p
3JdyVTqTK6e5KpoAYGiebG4Dz7dtBiJuy8QpJw9nrP2N/KWMt+uPzFRO4y+zSLLd
K4PhZvBZNbM3KNC++GZ1Mer27jp7eSrr1ZHUnhzPUylpFmtVqeOjeYn9mIdCnBtj
SqVPq3KPp25MbfB8AUMw87VhQ2Q8CELJwt3FbLSw8Ae7xi4efae7LJMdmPg9d/UA
cyEjnx1LYQ7eX2vmaa2eQmTvHHJeyUSPYI7w13SEMhTKQ2jXbnUnhkGj9oaba6Lq
0mCDua65xchIuvrPmmjJE9hq09Ga2o6UbE+yWbKfVNjrbvTt7gDrrAxwlb+Bfvg/
HV2zJ/7BfjZv5ZvjfpxcGPcqJu0YOWzmmGk9r08GvfOs2M3WZvpxX0Zu8slMNoJ/
n7H2XOIGBtXb/QjdQ7fPrtcI1VHyBKuIqpsneWSOJAqNnLSS09aF8dVt3ecHrAib
Oa35xcUJhb0RghgbBgsVN5r6WX9tT2HsVnEx7jJwEPvvJfkJS7zwVKwcJgRJSnwQ
bXIH/MdsTNQnIxHzWoU/U2I5NNN8/ThflXW/JgNvTRi+kF2TcmPRYG085zb3NY+e
5+4EKDOK9yCbjiuF2LI/5/9/B5IXcnpNmGxSXrB7htyE9mCfpMk7eeXMHCEjDEKy
dflTJS7fut5KJY2H3Hl3DHrocj7lnKf02Kf7VDvJzLI55qthhLgB49nOpn4DYXg3
9zZXmvSn3f+DA3WWEivTjBIc4wN45jr0CTJ0i5PIA4QrEarVz34biIRP7YeHhJuz
bZPfO3LOnoiMQ0M+opeb7QY6RzEeYPeBayO3v1cfBdN5q3pTQLd/IrimZOCN23mK
3jVuYP65FjTEDw0cq2IMdVN/eYJJ1c/iD6+24z+9WZOfzVjCh5WySjo4AtiA9lmP
1/AWHvMXnGQVMG+fjFEzPM0xhGcW+6sM1LwSQ7Lm/ogfBmh/HpBXCCf3MyGshUyS
/f57n70NLO57mqbBh0biB/cu6USTYlXqC1PrpnWJ8FLhmdOB7MJ+Lll7cJn9U3Tm
185kO1zpi5uIb/A+mbtPE4GTYfNZ7t3UN3iSKPdrUIc1OHQugFMRTy+mnX9AP5Gk
hYUKwNTs6xtc9qrJmbwFSMoqzHHGtap+GRgv4Wrl+7jEGnwIz5BhBMdGeZ3f6heQ
W5n4NLrJ5MiENZcIvugaldiCQqf8JjsSqyKsqF3Tf01KkZ1VOLv8T/NCq7BD98jR
ZVDOarqLlVEZx1hxjc+RY7BF1lnJ2slAh/Fv75BA5Dp/9I1KF7njGbVw2lzrr0Ge
2SiEDvtrWY4NCb/lNkVhBvG8qsLH5rXO4513lnXQboGAcIyPu5zVozUnvAnek1Jw
dc0rs9tyPgfyeJWbk9Cv840GW4le34Z13yma0OJxAzYFbLVu2dflynvzvppVPHPY
MR7HH8zJoRimrKShEOFldB4BDeuXzFaqX8YxGngnn1JI8GvBcThJC1oAQCO5R4Hx
KHJc4vxpuuOd902nQmSATN/5uF2X670ypIEk4jdu6nCmRIUWYnUTwBLMJCOf57Jq
svAWbQv3mMerA0m+Oatk48YXgrGbDaErjfYhp6SU2/QEA5ct3OqAWseDohQ5KZYl
ulVaGH0zoS42kX639Dir9hNNr7WimoYOioFP0lQkS/aWpel2buRDUFmcZtbbjGtk
hVIEkr584AtwANRt2eYCGLwG3ovcpAIhix0i4jamCcc2keaNU8MXfY1HDA3k7Ksd
XdHzX7nPzGVvqXEvrjnqdFxarbJCXSvIpOe5osBfXb1h+7M0VwE8zBks2DX3yCwa
vtMc0RpS8Bf28NB3M4dGTgO/1vBnBeBWro6qb8K/0cnC2y3Ic2lX4oDa7bwlAfQI
R5gy5reXmZk9dRS9bcgn31qH3LjNKXKqmi4yqWvM0mkXjT1zmPrcYkSXTPZR/INt
hyNVN+cUN5KIWKzLZZz6IPbaumH0+g6m76eFUQlfenmL+Cq4YPPxriWCJIA4X9xw
GGu6s7MrgQhQBf/bBOoMjq+joa+bfoJsiRuRcBPJvsg6ponNrwrp55FM90SPeG17
kkH/jv2scnCSqLxNMlSXDif74YUL+VCK6C+clt2/hVDcXO1IZR8g75vpfe2suLAF
tXa8L70mFF0IxunNmLxKN/ZDugTlfgUfqb+yKNvt/WIXo+MyWr+rDgroOTcqjTZV
JjAaAvGdiwTe6CRKdEsvhcIi9g8hL2UOuItB6z4nPho/CX/M45NIeLWdRMK9mR5o
e3ezrQPllP2PSyAsCbicn1xkCZNa3OkMz4gAgzu8wp0jUtszXsqZAX+9mvvlE50k
+zBXI0weDCHuSYKeVey82jXOObiNFdbLOVmkSqyj86sygtEt6QT1e/Jrg6Z/WfB0
SPSCmEVwtgbM880DNHj9wLNTgEu9yC49KfPnJz+z4JmBiSdCloIgKktjYfNepQez
Xhdd61jMOTDaqRpzEFh4usc3drwSRV2fiRhkl3uKdPh6EMH7oGFLW/nr7DGyiya7
TF41dAg0401xB9Q4yVvTGCQ7K9F5Ggf/XwyXCCXIOCTGCTUFcKRZN5X+2RDEd+pv
PElPk7UJXoQKcfLPKOYTPHmFkkR6d4TuQNCkl805m8dYjrh6eXZVehHQri2E5kzR
nsRDbD1oywyMDEG+rDQwyVjZBsylP61zOJeHppbeHV98kFeiQCOwUpkxOCRMBDMu
38keqZHw+Vv/00zPxCAsv7q5BqTyRlzLBUDByb4kh/fNM+nAUYkKR7mD8CaPgV3E
p1ZQE+dPlEeLf9O9j/yFFI8OQdAKY2e+06E8Wi0rEd9SXiu3/J/FX0pq2T44rLgX
NmnGdUR4DPG8rW14zk9fnbcJIHR0iDACoHrPAgepwue5kImt0khCy0XrDXduJ7SQ
gQ/JfDovHYYurKPEpK7ph6Y/WUYU81IYqtY3XvYgvaYpf//U/foBeyEGRAm9DoqU
06XLEHof1XimzQp2u1k2/gYkU2P+0AbEln61g4aMewMq06KGg+dcq85vm0Z9x2xb
dOweGTXTVgQL4j71y7P5Lu5X5Nt9J9dip6HWYmIK5/gO9l93RYx6rUeFNFp9id7Y
kaMB450VpWCBizvuoxbPf3KvaDQgTqh/EyLcROmiCxp/iYwUuFkwn28ukzeL8xf3
Ih7h9YxHZHq0MNk+keTFCd6mwzlJav/CJ8PDOyJFnDizJmDmMJPvyNY/SYr3hm8S
Kyl7gTE8nIa5tSVWL/p6Ds+nTeSS+S3tMh6i4mPk0JXFpPLQSXvVWBGbP90vT3AS
ajO1zW1Zas00VP3UI6/hPnNDuP7vtJHAirzvARCvlJzqt5R/ZjK1L2SLh3Nrv+Rd
4+HzQ7sLZL5IIxOwUZ3ddpDVqyQOQhDcw2EPjGPUr2Hu246h8k2YyF5V3oduqm5H
2VuUGAyqGpRsDLI3LtGe2hE1nrBSX4ARqHAJ4Luh4EUerEPxGp8xvTr0QrvOvy0z
NbmBgaUQrj/5iARAWjJbt/30BuSiRrYI184Ok++19WkRi63yO+GwD2D5h2ycQur7
o4OMv4B49sPRdviI8ZWfp+4+ebjZe6oj/PEUsytTtDKXVyoKcwpZNUfMFz49qcAf
0jV4yytw+ZFriFvbfC5AvYGmc511kzyXNdAW9/uDwJfr2ON55/SaxjOzM7MVAKPY
U85CZLWCUVxv+OjLe3S8IzK+wkxXwtqu1ZNCagoJyRqv+OVmum3mS+CDBigrihoJ
05/21AYZQzHvYiIKV7DFzkir8jH0zeV5hU/nxIQ5cx4B7KgGXOe+F2H9tMS3013C
qZ1wJzXxTNut6d5vv170JzfOkb2/Aw3d//AOCvNPpl6q/Em/J8k2ZOcCcd82p5NK
fNHf/+GYmu8rERCx2TwNp7w/2oBH0oJGdbIRaz+5M0EOm7N1Cl90AuRmRRjzj23W
qu94j/bXFFhcQwJyVC1J5+3WYl/iDfGs0isvuOwt/w7dZ10h2L33VSfIdmECwKZI
Rqtv9E2kS9dgRHJ2fniBvFYp6B8tSSVAmeCAPmI2dGl25lNHm6jHb6U8WnNG7tYU
tTBWpv7Fx7+LdLVwPBI8ZyPfOy5PWUzsP5EslhJ9aPrpzuYPlqENV9VbadwgWmik
pSiwMhMJx7LUlw+tLKJK2o80tjGCjIwau9lsMMiO7Uj3KkBL0X5wMDzfuektSVkM
v7HRxN9bYqarQjK8vdQ+mpDlvdTlBebKv4cFnoyaSVbh4fkA2fTcKogNbCQVimM7
N6FO16437tPIXmXebsphjeuAk8cJWQWHM4Wb4NgF3YBzw81jWJG5DaBwwrA/UkHQ
14yrhiRWFrQqs7cyZdIAfbNaf6uC5mviUefU2iNXE5/WL9otiigz7oGANbz0i6UZ
sRbD7AGwzoaHG2sE+1DQA0X08HFZMiczgoBd9as9HX/HQg0XQuFcPqEHlS5vemzZ
SNzyrhS+bzSEdhC3MEZuOoaH7cdAPQpZ7kGMCAvT73GnHf9nvdePyt+jrt6tqLkq
guMYzWXNkamJhXRjzVgvpYU5BXs0S6FTOwbmCfvOKeDneTttKnny0dTC+JTC7MGy
yirXhyrrfQiQIof8Iy3gB6BZpiVvac6gf8XMa35rVF6EvVQ1gikePojAgRpsAT36
iVLJY7NIVmMGqUfz6gqMezpEJp3I2V65SynGnZ0gr7tK732tzSwFeJHCO0T8zTmh
gzXWPRcI4M5TbOkpnuteKQivmmGq3UA0hp7cWq9rfDf9yORZBv5Jmx5qLKJW1k+b
WkaeF9ZuUM2xD+wkK/Pl3Jr4lf5I6HkMidcJDAD5OK5fqGRZucs5lbKteYPAQbaT
uiDSaidPb+h2NeZmN1sUlIfp7M+SD5TrHDFOz8/DrE0bkcAh6pCe4FassqUiCWFq
gAnyJ1yItOn2Y1mqdnqHqeyw+Zk3jkAPR/ngRXCSJRfl7KOxNzE3h8GPqlg6wjj4
dIu6jaPGBH2cEqNaHIm3KPgb1NAmjajS/cfOidu3+rFnLRKl96sEEuY9y4g84csM
yNOpNeOzg6Q+x5Uz0p+9M2bi6UsF/qX25iw0G9BecqU0/OndDQlWBWdoKvzr28RW
ax6FUp24H/yqTq6OXtHjoD3f3KWQ6GfVrUbaXDk1nkSmIqfBlyOKwAqihnkfRD9Z
3d9cgxiPI1R2kXgONLOGdnlIUOixqk6qxF1EyQ6jG1tQDa93AIJHMWYbHxLfLYK/
kyHqWmPpdjiF7oahlWWgh3vOaQpVGrxmrVCCBiZe1jzDLOUv441y6N9x9rcICB/a
GNgkDOwftJGcOarHM4s/4qYiSZ9uj4Vltspof5jY8GvaqeIzMt29qse5OlEKO0Vu
TN5F6heM7nJbF/+mX5IEtqyKihghqOgWRzFR3tb55vomugxyCFs+R3/DScpMJQLO
fFoj4JKj9hgTOYbyHcYze1EGjIdVNXHpn7Q33T2TIN7Kp5VoNm2lTCnHGZF4QcVp
XrlBiGlVejkofHP5yHJdchx5sygS7wfcF8mzCQrJFqkufEVx8PnL0X3vacPydhcj
zTow7nSIae7Ucd4AL8s5o5B6Tv0iBwKVXfj67HJJS6nZba2LF+aDVd0138T2eMAL
tWL5WwTSHoYZKDi33CdbVGb78/52g6MgzyJv0oBwRQE/AK+ld2Ei3Z1J6Vu+zCtW
PiRNEmiSfR/7lxf26k1yNRmM7PHG3FbHCMx52CKrtL7P6IE7pUaOaYJ9By4ZMyGK
BBdaLx1+v92OHLzdcdRO7pYt9RZ5AhmKkRA/Gtz1OMo/RkM4uj1tEUepDmWldZss
ODueRXx9F8KZOOH4WEOze2m0q34kNMNsR8pBKWNx6M04MjvCPNkhbqjsIQ+B922W
WroLuD5HEsJsYU814Gimex79ksTvN136pCZUU/4sxlf09slAos3pVGyLBJoKfesw
jJDEoinD8nVDLO286l2L69ckEJTYQTH+jFbyHQjcYOIxLGUvn4zeE3Dt8yvlPNn4
DWUUr7nlRy+XmwYn6v45wl9uSQdOmLyoFso5VvRhRyFJAy0M7HknZKcLcfdcioHD
766/QEs9YCFKe1j7lY5+01GBnwN3EnoC2B75MOOHG8oz4TbMsSEFD7jsAXd8D6Rl
yDAiyt45bL0RPo4y6WYuvWlGTKzC78tHC74QB0F0mTpPbowU5U0PWvnOyyXiSWGl
fn5rZR59K6AsqaN1Dn8fYMkjkfv9ovWESjs1o9nUqr0UKRJzz1N+OU7WM1h0le8b
cfwb+e4D6/WPPcXiGoSHpiaXXftd4KRNJPQ72Z3nrHktwP0tod5wmWCcpxcDhaoM
dsVaxHooBeK91IKpeH+E0e3lWwstT9BiaAn4wxqxdDytRJhCfgrROh6aZE3UrHd9
Uo/BdwKNG1JUjpYr42CIt2jIkklmQNIoEkj/iBQBY6nqxqhJVUK7MvsWBv1/92ms
92axYxDsNpFCPxfqQ6i5PbZMWOemWyIXU/T+oifnEknyA0JN3xlwLxbjnxgD+wom
SVxoBw7G4E+3EwsEJn5UnabdgAA5s2mQaQ4oaZKLwjtI0jzDXGp8JOrmbWEeQ0MY
dAR9z9ogHKlrPddwvJo+bl5Yg7fUHDyK2dRmuPnX+VGqnqRZOM4STD0/iIT8N5+U
yerc5/FkFuGWPYCPQcsJIx78vqdAIpf7Bpe6JidhEqbZozqAw2rCtmnxA6VFpjAG
dq62QJHXDHJtobR123+mwoYAKRIaBOpxyTxyLKOgFGjRkp+17r2mBxXIJV+jM82F
hlk7iplJqcRzFV1YQCZV2u4ARSCdGWHP1VbQ9JYehLWnIAzAa7mLMrXKFF0iHjuC
WAtZFGM3qBx1y8jmhE9VIlkHY3YUz/GF0SVZ3j96uQ5ujD8l5WB6M4ECXhSO9q57
CV17TDEJDaMl/jS+gvQetrzAVcoUdfLL5We6Cgu5pfP4W9twOXRwHlxSF+kD05sS
TjYoFtcxFJeqBBxBkS6JkfaqoNpjuWn3sbLkbRro9K4P92DaLJZG2uH0h44Kbc1t
DyZ9vDnCKel+mv7BFkcQyAx4XAGSJHDP9ZvEbFN4j12suciYCpuj50t9/ocuW0JV
NeRnPZV7cERh5jfoKzsKnoFJyI9BXXphI4r0zon+QJn6piBh/lwoDBkBl/ZsPTGr
tJKVeX4hMEtbv37PggYebV4WsL7ojunA0p3at40DwXO5wyFoFgwEhPqHY8hO2kz4
VJIW4qeJhpJsNehBVKGsLCFErqXPcBLfK7xFUSTIZ9QSfW8Gv7GHhdFAKXtPs+Qh
eqY/TF7udaZhl3rLHNEj15OJ1Aswzutj1tgnYUgZenwTNRxxAUB/F8BHjwvwVHaJ
bIGcjZEsUkeVV4sow4NL7FAq/+3/JAJkZXDZxX0RdbVUZE2U/2IgdTRS0SAzZprs
eeQmMC/OqLW+YWw6clNKrHEysl1I8VG2mnBWW0S1idjhW/gTdAH8rEzyRXn85JtQ
NFSfhD3iVHoJZT554xreJJIt0LovvVHqxk8K7OkKKxoyrd3NQkEGrbpr5siQU+96
K4+WLLIJU1MV0Ckvp/RehCN1/BU0yK/Q+nVl7NW5WTWzIIhqz363SgSggV4dTz9g
R+IYdv0eT8QotebzxRqm8Stne1un6060475QTejI6ytMyteXRVTOipZTUN2NAZeK
I3gGD7j5VeGwrZsl3gGsZMIcw0/lkyic2GMqCwsnT4jV3s7i/frnAJ2ZldTbCmXl
lkcaOjY+Q50NUnfm024Xgh/KEHCjhpy+MuqZBDBnZ1clN0gDiyK7GT6zf1yVBJlj
eLtSCau+J4Nrvk5oybLEOPKC+W4JCmgCTqWdcFm6ORuC2VQCWWXtth6Rw4uCbDWv
Mofw4CiQsuW160FCZmzBkajvRmu161NyO9BaCY5XiGsoBJFXkah7X4T5FlWhAiqY
/pVoDEhu12b0ODHVWB1ON77sR76dyIdkYiIj0sAz35L8YFDi1iHKo+NxDYPCzaEq
V1XknS8RDtM7xEgCML2nKY0RpOiTYvi2hwDOcn1G+6+0SWzuCNqX1nTTTyD4+Lpq
uWUqAJqT1u3FHNP0DpZ/oiDoEacIXFZj39N0uts04ZvjTp29u3m4RS/CcUYY++/8
fJAEoV/UKIhgX9CGk9zaOy4ErFbWlHUnt5/NhPvN7Q/RF6SDTGgsQ32u8BnFdrgf
vYsF8xksHxjiUlNLgRe9P7U8cixf9uHp/quzd0tBEM/rpkKPIBvJyJ/axWsQu0wI
iwJqLUN0+wB1T2A2F33LVmk4M+nu8yjfbbkhbkv4FB0SP5hlRcI5mUAcYjlzRrUP
sIgwYwiKQYH22Pd4eB7DSxnWTM7Xq3bTBpVd+5KGzldr06tUwkMUmjPW8CMAr+K5
o9Csoz4VqNm2Dkfzd0N3FLeFqp1wkyqiobtng41OQf+tRVC2hWrP/cGsQpyH/q8g
/5rNfyfVoxGcuJok/85b3VMT+QDd1+NjRiMnMqsWNUm40dQjRyrPY7xXnk9QlLvz
+H+CwTPWRVfOsXYnbBtmf5J3Np0kAqjobn9WdU1T2FVuVq2ALIB6mB+ZMsCQbM+R
nbSeyh6Kiy2NpVsuCmGF7NAqAT6yQuU/wFNSv1BIlgiFubgBK3o/np9lNsISEbal
6bYXK8DR3X5xnnw6JQTG1dryV9wzcr8pC3ePoMeL/Z5dzpiiweThAm4j04mvgVan
nJyzxNisZ12dN95V49/1gNBqPUie/41PD+gqOE9PJRzDeq51eHjYOeEGcuTSJHSr
ImVnN/NWPJkWHWZjDDdYqGZISh+kPbejFFCGkX5Xuwi74yI20k9SqvccLjP68P+W
IQe0QwhHC4xDNgWkW5xvUDAheRWNj5rHuZD1YcvnKSJ6qsLaBbpoKTwUl/AFKwwO
TQLlXdNvzN2VPT+cUjjulvLvoxopcp1S+3pVGMAkiyauuZXYPyr4eDqVYd7y5vXq
fAxHYYNKsafOv3FIXL+Mc1rtE8tbBLkf1atu5G+JBKtW2Mszv4AKWbeWXE+BiLM3
xbbjmVs75h9F6yFtBLZ0p+d3Vf6cEMuE/kH6QfS7o4gjmiLlQxX9muSXAL2IGuAh
MQGhS29EFJ6RApEmrTZJUrFMBGSWn/lfVLpJXRVl97wxyCiRlEehx14lUNq4Z8cx
+mjk6xzScnMKYido8IAQRTIP6m9QsYLcAVJib/+YhqXjNvJt6zWKfvk3p8gQMqmO
hXlhwMwzhtM+nCJonwsq8p5aGmszP4FyVTqK25nWJznu1mqPwV6l3p3GgJ5QBIMo
3UB4bXMvn38cbmkL5u5aBWBrLrYBOBXOKZ1s1pfHbDMYvJZh8CGzeP+5p0pJI6qu
Hm40uqN2/GVB2Q6nar1jlu6yNck6NPaBJPYrAbfc6u8LEW3fY+eC/VkkwcBdNVCF
QomDqNdZV2+Iza4iprUs67Rzq/bc1QZrfdsz02HDjmVRzVfHtKhUZiHRZwIocwi6
nKqT59IonyZkOdi0+xPGOy94Pr/UES6tK6yu1usV456RjiOhJFMKmpMTohFxOjcg
ROI/yLDmtbt23m4MKjW8bnUWrCxA/T0IWGkWCMBnevL0MbSw+yxr5hpPbd1HFZut
LuBFuduSUCEjdci5B+NcvqyAhxHOsDLQbBG7HUC4MSejpI4JXz4aALy+2Yn1KU7I
O0alTT2sPwwy+Bynuttt85eTuTCeGaQJQtFpEkJlARksrD4X4IWtSuV9EeX6ApXY
i05E+QJgIShRNbeZRbXwyOrH0z55dnSi8QbO+AWlyLY0m6H7yl81B2C1PWz8CwSU
kCdC9+zE5bpyFUA7jA3Btiq/qGeuzEdHaLxLMaTrs6NAwDVoqSohcjXynbfMpXxH
A7d4QQz0LDq2RPlUZ4ZqHOl2v8QoLFhEMv8bFafVkaSuxxaL9FIb/U4xzB+zALd/
j6FC5aWEpMvK3J6LxmVPHe2Sh8lxNj31fEefctphLhcwWsAchv3uDl6vEHM+Yf92
AOL1A9vXP0tUsjHxrfWNC9yQUVMACQsJnw7L0YxMiRNVZu22Si0WaLQWKkrxC45m
0HK3VN0tVfsZwBbNHRTPtu5L45xiz36KoofbOO+htWMwD82wW1O/IjdnZ3fjLvoC
CicSvA683Fn/6XaZAI/9+eLM+OolYTi8OSJR35WxyBmcHVgjKPu2syvWOnfUkjvQ
/c1PRiQiRy73JHEGdAWPW2wxhu38bsr2IonW1PK5SIJYnzdGPtyvCmsSv8gHNEBo
oUx7taXPyQO7XwdlCOcdEtfI5keDC6OE36ZUbuu+Vvt6PhXvYWX7qmeCmuBkDiN8
ALvPY7eoL+y9lQvrMN2QGBEi6i33VHrvX2XlWU8lWQuynZNvUHyflbUgwD7eFvn8
rMTBTPOwNSAUAII3f9W28ztNZRxcUONVsv5zwWl2yOfvEe41FCJ17YA57sGeZ/Yp
lJZ9CA6gcNQBlB09sJ6ZRsqYxGdlD4r+V58QpyReWYZYl2LFw5U+qJoUdvYjWVQy
/B/uJLqTbANhxDVMCo482QfYc2iRPCxCMaiKK5dRyklHtpfFOkmaF1rlmKSV4esc
iclmRCrJkbmsgrQjAgWI1oAt8Q89xzdu0PvpqJAxhLF8ojUxi9xBANyeN435UuqB
AgJRLQW37MaWnCG8TRCJ/IuD/vIQ4mUn2VjjR7UJgqj5OqUiC0SPW5P4bF0jTUtv
iIpwnWH3BnICGQOe5cA67wkgQO+qxyTM9K2JFrbL3Kuio7H1nbJvRUFA2braZn+o
fXL6kSsSpw9vOC57qCdgr8IOM+xry8rZdi6OzJFodHXDZPb+HOY3XquhcydOevLj
AdQVnIjimdUZp6vHRJTVPeEBxJ5P2OmyIMAGuxJemIac7WJ/OtzVxG6Rmq8C3hb1
98RG7jAemJrPQ5pMzDw7v8NDJ1K6PnOLNafR2RVmlsJ01CqR2eutjHPAKHvpZWod
Yuo0cDqZPtULkgmmKMKKEraGMefGLKR9F63PuXQLGbcWffVBn84cjhifBp1rc5CW
sgYFkf9n0nTOZDy04QHBvbE6RlKIr7JYqwy7sAQ5n4UPCxWWCt43cr3nb0Z79N76
RESqTuVAh8CT9tEZbniUTeIxTbnZpbeHNgqXc7CTU8k0qCS06VPVcBvWfIJ3eqTV
tZqwAhqPuv59fq+TRC/mBIdddIYkpWDZSZVxGgusnklpGmatPvyACw2wbBJ4MAGC
Zg7aXyXdvabY0ysI+/IsAnSF4DHyv7W+4AvXhOugfqHmlO84napgTJH/d2h/9kY9
knZmJR9Zo6dgxYmBV7EDojj4g9QNx776F3OeNbGbCTV1AtPyGer1NUfwIH6fvtfI
SeVXpfr3+23nphPbp4V2YMqABvFNAc/nM75VefbtmEO/7Ta5QIHre6jhWq7TM1vc
oQeivXzYFQJk31D++nQO4HDmg3sEyW7N4W4Xo5daJi4hQfvU319hchfKX8GBdQzE
x1MGvFN2UwtMOOByL/lM6RW3ppmvjICdQB+j9EPNJ42HfEMY9htjiNKZXjA0J/q/
oMipp9y1g7cUwT/ALdh9KOsqU5LPbXpd+LBLok1bPzc0WhMS4fiH8Hm382SK356F
1S8gxGLhAF/7QY9huofV9E2Zofl0ckz24LVtXXInjGc2D4BTSwoKEUVH4h+MntKd
gduSQ/L1UGevDPHpgOG+zYoNNXgsMJnSM0N8lFxUfHfz80oJWjKhurs4XRNNIkpB
2Z7u6BGNCq4Uf35nvKb/FwrXGqU77KitlDVIstwLxPzynlU5m0YeBGUC0j6yy16n
+EX1tDnEvgDmd0AZ0o/U7M8KR6F7hoUSd5Gz+Zxo+4Flv5J3MfxlxhQhUKRFmc61
c1uFK0CcA0PLZKgDoWCJF6jJrWbmC9XJfegeNF4gP9/YR+XQtiHz6J0C69hLpt2O
xcBMCcCqfSqNiGt+oWchc7dAA4uj4+BKxlRe6MYo97F41JuFQTzX0VKLuQ2hrkut
hymJCdYPH6tN3yBEN3mvONMeNdY702RjW/qwVnGELBVpLtZ9QC5f6nPKr/96ns/P
8QRAdTnudiBWBuOSKfDvUL+cJm5p443EtQgXPkYw80q6pCVoxoA9nTXd6gxcXsWA
Bh/RbpM08FralD8Rg5kr9X1G1afMH5ouD37ewgTJZJJiFYyC1mX3I40lABHOj/xB
BTnXqMQPFtXomlqPyATCeS4LlemTnQGGlhAEk++LvSEECaNRefNPhvm4mbfyW9mF
+UG5QRRo1XEpevJdktwZ5v5eFBeZrw+pEraOOxovKmTjMFFUD2nfCFiBPyurl4mP
Vv55ayZ8QGPVTublAD9pSNUE+6o6kgwo3FyjKIs7mkIt0OXzm+KGJWS7f3G92bkX
245jLkGI5/JKSD+AhuRXvO6BwlvUa/z5q5EyO/FVMSR1hQIiodCwa3f8yDGanTbX
tDkFAIGQnIS0xYdOFB89ebYtCu3RTjtiFtZC/JwA8dpFojsQrYWsMkYr974aekoU
OyfX8VbIuOL6bIoS5uyg4h4Inw7SEYEhxMg3mwJF7Je5jr1rxQ4iz76xDwrh6iyh
1JVfLVoiaYDKXscVOsKfOMBQus3eJzVwJ8pGhJTQgAfVUr7vHyEZL1PFoW+SGTwc
XyvcY2gl5CdxWvAiUNCGS0w+CHI1sMj/pkPnHcHrlfjh/9vvbiIhioCafExV/FS4
7x0WI6fW0NDCFfmKZu3Ze5iffmmNkoJd/d6pDGltqQBCrScaoM6Oj93elmNQ3/Jx
hNucJjbUWvTQ6+tA66wvzv860dLJ4mrwog6rGrZnv6uQx/XASP4O9zfVTU4YdTwt
khCVe/ww5QRFzzt6TqXk65N60e3O9cQt3vMLbVSw9ZWJ0Io7TLqhYSgItZTtqHDF
XOxjKOWXZdFUjNBtbaZZnO3IQkwDNetGREJuxtvZRBt2gcPV5zswCklbrmZdedPp
NH/TkxXR/HBxQwOIU06dgLm5qVhdyPGL8R9DgdJ9ZewkpTJc6+VbjXVXrBs66Rbk
kTZ/LvG3bCyLYdOsHf/8r/oYbmHJkIB81sqxg8QtLGk/8QKvbNTixiW0kZ/7gkxO
rPFRRP8xiF09AsN0x5trPMkbWD34JC1SMFCt8wW7+RUUcI6DYLE4p2y9Be/136YY
gRitRb5WH7Gv7zV3Uktd0tkzCAyWR+1b8EQKs4ssusKTaj4CbYb/lDDvZJlkYl28
sEV4uovBUci68pgmSa1evefDvjIMMOvVdUVrUcTMgrnCspBs727p+E3hpbkAHA2M
Q+tJcv0XiAuWMmgkkBvqlBx/YUGxZIHGg1u+dFOjch+w1RMm3gcg1+XSHk8dD4lB
uk3l3YPPl2xs+GiLHjW0OXotDcFGl1ya01OME2i8xfZcAsLVJMMN9mXWop3y5fpZ
H1LZpPgJze9hOABx7tEXHzBA99i8SEgvDAkIBqx8Rr7hTdco3c7KupcJJ9LJ1tkh
HuRFhe+NncpyP9sbHDSU2wswdcwKGgW30KvXMjQzG5V+AJdx0cFUSOydDf0yJqET
ZEbJQl3Do0NlHAdUbPOeIZ7Hbsy2mj62d0+2vYtyKCFJfUI/Thea7AFprX6HRnWj
8h+uomk9rw/W6sVT1TOrlSgskXauEJgqNo2ya3PfZyuZGTHuAWwGiF+uYM4YRzvs
L8/TruxZXYDVbFfqqnTh3VWBd+lA4XTnFF0Fru/i9+/DaCbfUwnDt7oVb9B0ePw0
lbaj4dqCruMK4TAvIa5xSYzKNNevh3KQy0uqEZ3cEiP958bh6f0MqGi0+zJ0/CKY
Sob2mdT5euIDkUXtJW36zJLobwuKFKNWTXxUz4cZzqqDsyx8byb7xPKjQDap5LDF
LFuNOQ0mXtpDcHG0Vl6tG062khi21+kMI4CZEHWVeHt5d6Y60pY2uNnSjG7w00nh
W8A1CCLDIQKJLE5og/kV9JCShapZtwXBH2VgMIxdwWJNPIOaxFw/KEBmjPBq0O6Z
RLOSgW1QCqVcgHsv7JKT2w2uybQLKVlUbciBxvrIGwiB3o/Bw+7Uza5utwYSd8MW
Xl49wakDKYEk1Ur7N1nI3ZX160uXOA8l7GduoEGWnxZd+wtIHwoULXXh93m9FsW6
sBckMSks2hXkFGx1VZXq+j2S6tTKE/ygukeklhtTsD9nC2DiPtALqWJnz0f+WG0o
gvlk18MzWhTfcOT4Mk5r6VUZg51gkcxCt0vV9PMVsMEqvd0m8oygBg1gLXnBctON
/HwfC6xKUSfaVWTi6kv+Ka+UnftTxn8f9v3GgFrS1upkagCAGTJ0db3s2O3s3fzI
uLlN42nhK6CioyoCTt9laLyri/e9NpOnP/zaFo4kNvgraruS2IxNAAvbI6gkIHfB
bq8Zvy/M6V4F1iUwdpUyOpoll//RdRyHwMl+Cpw3R8fFM3QIEJ7VvL8ujgpwxGV3
o+Fvl8zxroNV9hB82sAQCGFz+BRihs05Qj8tUVqasb1GL6P5tpB185nlbLNASkWx
aMJR1KOHvy/kR27zjEwZZtEBqJwCiKQV8ntZe2NFrg7UvQCA5sa2BabId9kSfedq
RTucUe3PHKXrB7iuA86u2IM0bTh03s38YC95W3swMXqMrlj2tt84KB7Q+0RdyU+v
kqgRcehcdQZcYdHPSrltUOoGKPtflyZaIJz8uEVWCwmFXE//jzs+1fBxe0izRo4a
9zt4RqDWfmHKng5iPamHyfFKFYgiFZ6wF81Shf0mvmC1sHPm9qZKAPP+1y9A/cof
buiUncmYAfu0OhMkLo0AtEMArN9T50d0ppLTkUYaVBHBAk7BYPNhwfML1t0ygVP3
ZFNQvHEN6p3sGQ069QnHItA9L+UfOVDgPTcpuK/aHDs7XbKQJ6LS39mk97rONuSd
4BWRI1342DFzBYEYNz7zFJL1hM9Wo+uaW0a+XxmvdI8DlppkcxGPTDWtF0siAhFq
0A0LqDTGtwZ0BTUHn7MzjqHpisEqVxP017b+vwrOotsOBgpqF9+Ptj1meBEiTqzy
OsWkFZIw850wMyLTHbiWP1H5INOTK2BToZE9yHS2woAj6skWZInaC/b+0OxrsdTP
L27OE/HB5dWxzTVt0Z8GssiWcMpLE2G8GKzQ78EZ1G3fN238xIo3ljq9AiZ531Io
evp679tytXGONXK/vJELv3EUx3wFLr8dVjWzCE2lPykqOvoF9A3GCFAv60fL3gBH
o0BtVa+JEftEXZEBIHXa2dt+qSaPTiniercgshl97yq+W+izL/WCFDsYpuuySlD/
Far76Uj9kwhv4uSfNj3MXG6YaSErEpki2MBSiYwFOuXcQ89y3f4stvSszm0gAq1N
lrhN66wxvMs6I10r6I84+EVBbufzE888lpIzNGBJDESrvIu7IAIx8dToZLXhx/yJ
g1O6zWqndtgrioFpSgCRFwwt0MYzlw7+I8Gy4WYAGdPJnEo5uDDd7Ps/11ccHE4b
1MxwdCEFdW1KhhfoZxRsQ5kAuCnMGWD+hUA1vijt5OzkZvk7l+HtOkhmt31Ac9QO
tXLBwBP9af77el77hijMBPW2fFzaODukyHi2FwY8lYXzPRwuvIxVwml7zAaW/a1A
biwOlUoCQoj2EdpFOt/0WVci1tp9g5qoX7yvpQAb9MvAxw0cr+qLM1Zf6OYGxRTP
duDXtBjcwCI8sLgNCXTMsZ7Z5Uk6nfdjKQbmek36QUuUYqBp+djz4JmN+PBrHvf4
VMwqFQpKwIOu4swyAgcjdf5Hbkzc3lxElCsspHFV5NPHg9suBPRikfym/BQrklbo
ccMZO1W1TrTjX7zveofuQGm45yzdT0rVUb0eGQkZJrAO1zP0fsQtbbsJutq/gsJA
IvuO1xpL0IQQctDzH18vt1UWLxUEnP8fmbw0ELgm9Ygh66S+7hVAWj+oHkJslTNv
YOn9ol/Kzmoq0EyZ9s3Am41unSv1esyrrDx0nG3fY2e1q+Jsa2K3xhfXm6VDzpVa
3m+G9GLLW3i9PtXbIqPBGUYyjRejvDasQ11HTnzq72sZON2L+33KatVp7ktsXXs0
VjPl4H1nhsJYA/qwn0QVKCv9sCnvKTKkCwJE9kfdGZ+e02T5hOwKMnCbkg+Kv5bN
eqwTU9tzSfp95R1XpQGIrt02u2QBmqKBVdKz/6ySjYmMDiWYRNcwITc/eaeA2pNf
Ch/h5sC//haysMqFqAe9UuVaGFKgKNHgVCu7YoZVYPSswfsi/xVolMfnUBDzWaPF
oU+dGqZEWejnFZwBzyuaDCG/gjqcCHDYjAcI5xWG4aqGCgyg3NNO5tBQCevXoJNh
VCWOqfO0VJaXYoidwmflIurcQRuqFZZttiFXhrqZ3/AE6SQwnuFqavsrX1h8ZNq/
3JS1B+zAYYvShn59uu7RaVd8fmhZ7fRAOGBUiyxT0agbpTxi0A9rX3geNk8fNmm7
gnZzetR6L/jYBmYw/654BdOkKe4DTB88oqtUQ3busMbdUvuza+cV08WrR44XVqIq
LQMjnaxgjSgm8lrmzIZjIgHFk8sR+M0nLqGx0UMxdgcTi+0mf4KocyO4A0WNhGhG
OA1xDeqFscmwSBBtjGklpNXntcrEvAaS96QRQra0LP1732s/ux8ArQUviW57RFS/
ao9GDLixPC4q3juScXLPXZhfjlPsk7hMIuSF5EhLrwJOGw/B808hsYijS82hRU5F
UgcremqK9awJQRtGCsKmNHBP9ctOTVl/PXrPu95KYnG+bglXZG+/ka5A7G3iMpJ0
tJ9Nm9LS88W+67hwxDb0EKyjEzFkP2zhrPLRJ31vaDsaxeEllZKoWRx2dqCVbCA/
zsq53AQ8In7C3kYt1NKXs3zUtzohZpJ0MK02W3ZzhqiuVhASZRE/RqYi8SNbDpvk
qf+ovhfG+ZvFgFZ6MWoIizwD3MDzLHVB2wPMP1UY4YtyhzdIBHJjoS8Vxclbjkiv
Q3LOg/oqrK7Vbg3JK+wMolN5dlDJ/IalcWnj8YwxQCH2bdxdUdAHN3YLRj+bzgvd
U4RYkmiZwjV085QRCGETNqMnS+8olTCnPoMTq5+WwDX+9z2Uwv0+Qln5yGGZ4edS
Tm73rnKfBPo3w361JhRni8lAwF+g5ySA1utgMgMdA2DjMb1E/PMCfVvoOdVbhDF2
RYy1wIgwkterrliyuTwSjwgeSXPyXIPKCR07XZnyQqVu8n96h36F5BlJiL5+G53T
SbdDgx7Dtz5auL42N+TCqL343njnnfLvOd4MYOaBMEMoHKyCjfbX0/8ossQfoOa3
IDNukyrhrjRPpvgif3/iquxd6ylHY8uzyFr71xv/BJFou4sjTFm67tD3/gHOcZxP
WqLhqIYsMx29FYbJ/VBd1vmGo0uE8axbz8OFl8xpQSs2rxES0CO5/aKTB+siCdAx
QKC6b201vT+G1MuHPfDS2hu6rCmi9G/ku0vM3hPgnGzQk4QunNKZbe4qfLBlrE/Z
mhQEa7gK9y1u/Kd+qdwqaXaLhG/99/Xuje50VCQUlE9gP5sUPblQyDl5h5htaVQa
gp1QHbZDxrpijImz34C5XD0YupU2KJcT/Amc6uIdTg6I6PHpdsWpH0o3f1gY0e08
NrrfqhsVDsurTG1IVMIqUREuYOxtfZbrt6wks81Ge+1gBwljPBqi6W/td0tcuBk8
1pHHXfo+FQbDD8yh1NMrS/arAibcv7eRHEkOgN5J93kGt0BxgsEbLXxRtgJlvRDB
EhllhRJHbqTZ7kiQ1gZCI8rzhRWSWSlBZOt/gHaiPxaxRRXNSLLxxmOX24LZbnnF
0PfbzbBK7/vl3k+Bs/i1lfri1IlfL2rhatixS3JoBFv7gPTND/QXi9+l+/BCjfQ/
EFUT3VxvWWh/a0CR6xmAnTCN1NLItcxKKwKoOysES+JQx4wYNHlFuvOZyAwMu+3E
yIwW486JkEFEY37CbApttM/YvLKxsGcy5J8I6JZTdwuS1SUqRTYHgrGHyWfNX86u
P5D65bdhxdtjSj2CfWDQTBLn0TTV/B4DDvDLD+LigoC0MyK/PPmVBSJhnX2rHl3A
Wp3H6L6a4Qv8HoFpTL/HzCDUh8TcVdo7eBb5eiWL4NH8hZJ+Dt2OTCMSWpnW9b9i
INLK1tWyn2g17CigKqawOVcznV+zLIfcQcXuupvGU1UjtaomOAEtjPaVxHIc279F
VX1gSOwXjMOwuEKb199uKkDSzPhcE9H8p2HTKJr9qVEhshgeeO+wufdyOHYgC1+X
XD6/207EOy1CNEXZshOHYRaHpTECgz3oQP160n6XS1m94lkxDmvbPYGxRw8lo4pD
H3iVtSMfisEM4KssrEMC/bV45JZkZulDfWHOOA+0qlj0n/guRpU23o4pRe8eBL04
YuucCPa1vN51/M/qYRFl/Q14p/d76XVKjF8nQh/KYkrCU+IldRp+4ldNw39MiEbV
xlW4BiD51lCxYKTGpYXwvHL3qjxQAvKe1V4aokf3Q2CoMAvdLw9yutFDdvVhXHNI
aXzncRDYjjokBxbHWUlygyu0nkPySWhHrVFKat5MzzUbCMjmiHYPNpZagkRqCHUW
F4T0VDknuzlQ0aGBcY4j1VgzA2F6LhZ+IMMBJkeUnnThCfk/874soaipzf/3XBkc
iSg8NYcVHGY205EOu4czKdBNNXtW/SKCI8hsWpdeVymaHUjDlPWbAfH151J3Oqpw
wWURyGCIuDoYtcleiNCX/7IWZkWN66JWXZ9RF0y8ifI3kLrNqECiKJLIBx8jV6nr
6z/fRU5Bh+REEMZDZEnJYFobVOJQG/sHUePJNKWinqPSfFyHNaA99TwT2cB68b/1
4ESB4TdCoIY9jPb5f/rvZYQjlhJt3x2Lp2OlVat+peKihYhDu5Ify15Ffbdo4xK+
NM+mTWxu0bLygcsM4YszrFVa8Fr2669xT3pcuQfoO3++OdgSokdIIZxMczDS9R7e
cV2gTz7otLb3hLZDid29cKzKFm3iGIR9p7w6sjglJ8vpmK8Ut4al9X4JNui/anAI
ct0Luj2keplQ59mwMe/f1PIHG0vYFF6fXbrEKU1u4457ZEQaIWiJTHYlpgx13Jsq
ORNHi5zC0lZk+yD4HkEkgBLHPznzQwBd8n0sqh1SGtrmEC2CdT9NwV5JuTFthl7a
9JKbajrhXnlh+h446Ej/IAObQ2kP6AgAhp1wZsn6QIIPU8SOyNQdNqA+5PWocTsi
sfghBaIualSshz085AHMQTUTLFh0Cqk0Ov0yD3xOMnrq1pCQ5GIFAFrt5lExlmT/
F2YuH7J7wfydJLgfrhPNajgWcwbGXNk24mPyrqmtp5VcjV5nYWvFbxu5PIgmTjcJ
jbakE8UqVqC56kJ86x6kzEdpmCAJTwcpZEhxLGRD27vSdyUI0oHKGjIbYNGrqZxw
EU1rX/buSR0x7MY6pr9tiDEWIgmg0MzYcDCxzxzSSNy1QqnNNqeNLGVqy/fF0ims
eF+IfzzQonOtBvwpDA49FNCynFH5JRbPT6oBAnBgFoBcBQhbh3Atjw7Ubn5pKpjS
EZhr9yqzNS54XfOdTwHHtcGAvD7izAdMvPizy6oXyCNVOfwp14AduF6xhaH2rhC7
ua152aIU9jvHR+nuW5mEqP4gbb29mvlqLrME+/jCS5NYmtnHXGweexWFHGMRRkaK
RssrMx1CHnk0aEd29eDehtqk+ehEqnUoXfi6s2OvE2NkHIHHAhQuql1TTL+kjCn9
hlgfV/L1gAjhhHA3lEZ3E2iolxKT7KCW8Np6iQc/Smk6PjqJpuNMT++djI0wpJdS
G/TIX25+glZgbw4LPkWq2tLEd5wo6Pg/jHQ2eSpQ7Z1KA4q/Muen6d1xFstv4DII
FgkZSm2s6hrxfME1YUBXU4aikn+NDNcr7ERZqb+WDSmM+qboWOm4Oyc03XDCTNcK
n6hR3Md/odXrUfM8zsU6LEfWPD7TK7OuiYHiHqD7pJ0Oyd+qzIyueifOt4ZBMFBW
j1dCB5Dne/rORpFFeRcroaxAFA5x0eJ/EVGCLUdo1qyb6jrhdQcwppj+9wvEaki6
E0nf1nyQEjHJAPJkYG3yM8rIWbJqcy4dbwlj5kMbHOd0XuvEYRmhmQNG2o7VSxVA
luXAuZLFkWa9GOSggAMk/hq/HX/qNMo4/+/pzetYBikUzat0PI8ZaVCurZtR0Ixm
Md4S2hfgJr5S+oQCJMp++NuUp707TjY1nJWWIjncI2sc72FhTpG1cFH0UTGp/Mf3
TMYa6tATiUxr6n1h/6tMaESSXJVIvgfYpBlco6NngMXV+xYo8MEdoJCUEW0rXOXg
08/ww4brL9ZkFFwHYOh2uW2ZP2e5CjdadjmrcTzQLzRjfvpju6taf2WM4y3ZHaXv
ht+SqQ4fGILWZS9ZPNsDIBRTs9hUxQIg6SZtGwXlH52Jy/cBmkK/USGh1/ooSs33
v1F6ZLXDiawZ4ykanpkXj1tA4/7EF+HX3K5koMPqmbehmRnHld6YImNWwP1nztCE
52SHDQDbno7g+iFyAEdHvo4k/SplebpkLj5QEAmN6asLp8rbbtX9TD2q/vvbzAZD
P4uTaklEnQln+kjBEuc8p+H9jJB6ZMs4Yhawt0KebS68HHleyo3PbFuSI5VtRn30
bJ+VaHgzLqSci4muHBIUxhl/CSp3GG/73yqJpKVyJT0OdsPOLj6cQMaZpZzpEPqT
K+iYapQZ3n4BiiOEJNODN7tSuuXrYU2WwP4x6ztwvbX5AhIKmWNwPAPK8/JcbO/H
Cic426c7Ek7WxgG0e22LmkudfjzPJ+OF6F9jcpIbE+XLgDozZbsUjVKNFjXgQz7P
p8yKzpg5hCKYIYtOEUoXynAjcwofiTZtpQLuvb2YuBPykYtVYqoLEbNC8/eJRs9q
5Lzpdvqsr8YVNzIEDzJtnZSPU1SxwAwnM4cdm5AABN5MCTLQGojJAS4nz6oCyCKE
L1jxaKTBfFtHpVq8i9pyzrPZg+6igxGUn57+E1pQIQZ/mlY+yynYrCZJqM0y1OQ6
0zPg6gFAReDBSKN3cvl1cjsbTJRmUQzsBrJ/gxbOV+fY88ewTUiCOeVBwsoahU4i
Yd4WZb3MgEwj/6qSaKRQMVO3kiQ6gILoLIbkW34H63YhIem6gRuRSDS70dcTlmfp
scga3qNQfSn2zjMuLIy3qUjURkfIvOg9M9bMQJGQyuRTLv3VClsTie+MKNyHBr1C
BqqzFWfPHu5e7U6+Shjkjgjop17iV5jMpE28KWaUCYpRMk7Itelcp9F8FQ+2TmRg
C+dHjN18IWv9WbIX7jCSbBKVwXsG6OahiyUhYFaL2G2o0FO5xw5zSIurF4YTTCve
uplHrdxNIvoiSlKTJo/a3WjlnStwoPlz/1zhHJv5SCMVeF+4Z1NPyiO9UEJDmDAo
H/5Yfz09L20v9H57Am/ASHRzHIJKV3uV3bR/EQ8XQR06NggzNPFNVF46KbCAa6Sr
Q3Ef5YhRqLpavRYyfjWGoTJFWeBefmzAVZXk9j3juHIqxFGRCyEdHgOVZLCwjtUs
Hh0xgrmC1bO/PzUHjRBIRR6YTWFFtLszj6eQ0gT4h8uEC4Jlyw4HJ2QXfT+jL6rA
E/tFg/yBIIJWEaIEebkC8/sqGkB8JVpQKzk+t0nxoeUtZC8v2Uhvrhhy2UkynMa4
q82axgRcoq0gTLl5+t2l5ue6rsGFsF4ZgF+7obzcD/FtLx8SMeZwuZfHD3upIGB9
Ss5p0kx0xA+PjXX6L2M6IUI/owl/Sse98vHLQMhZrzEV+OWVoGPAICvNn8OnG/6v
G7rNzG7ZhgWgZAZ0nLsqsh294MvZ3KGL3dmT66V3QT9WYai8/91utYYRPMnq+Dl0
IKCtOBV9pDIL3O4FkaLJ2UjHtwBP680ibCQ8OonE2rYJJtFOR3tnaNbBYQ0JqB1b
Ff4i3Iw5yhSU9EBWtwMKw7Ld0Z0FQWqq5Z6QzqbRXVJEHCfRuGYlbqKWPJMEqDpR
OnbCTYEXC+5Hm6CN7yMl6/WzfKYRYXp1uxlP5T6M+4l6ZWh7Aor4FWwPNmHvQ2f5
afI5orgciLfG6/ojhgT82etCD4pNvN4FViRYnt06jQ0HMd3xbMvLMaagPjWwRXkc
yluQCc4rDlErG6F7k7nGl+T/sirUYjBmfGPsMxs0l0uOrZ6S+ssmsG690lj3AvoE
3933/6xgaa0D+2RY70IWR6pN9MY36FxOQeLAVu3KbIMzzfPKxkvKnFddsBXeTxJ4
CSKSpTtV35NBUMUmgbLsO0AtYVWslJpc/2QUb22lrgSrCrh7X3kxRq2SJ2ffTXBX
C6UsATchswEGoStF7OSsjRBVoncdBQy03X3Nqo3zpip3+7s0OCUkiZzVA/5+jzJ3
BhH5N6I8vG6vaujUr/dqNQs32pinKkRfDiVdl5uLOjSWl1ERNEHWU+yH/BBQlu+9
nj+Lw1viaqUfmdUXFlST6xHPTKgRgXEznIRIDDSh8dL393f5B1RI9tYCGaDXjV91
h3Taa8SuUhtFOEYa66KhcBsxKtos+nkYSJyAGswgzVrWEewzARgIw66kXWeqAUBU
2tfceVZLpL5wP67Jhvv60BWGRBrqQCL5AwyOTbh4WV3z/UHMqZmemLxtYl4NE6Ew
xxqxhRvEiyGVXAtAFz26r2UI3rCCIDr8wDSA6IWbQVRqKneMlsl8g8b/G1SQ35zA
fMCNhDs+cxm80HWHpTz4pf1hBw+Yh9lhD/EUNOu9TmNIqSgoCelwD486lAzsyQVH
64NP+8R+9y5lOLt6Qb2Y6s/YJx9rDT+9/3TkWRY/OAD0Q6zZ8Wp0DFXXrXOu9ssE
h2YGNBCQqsmSq1/CF8zhBBa56rjeE0G99B9lpQAqJ5ky8wuL/IjM5th3fRC7/3Nf
5A1rORiruH80c0nCkrEglXvvQpal34LEXmGh4HuPxMcsqnontu8eCKO7WFW5Zjrt
9P804Wil8iY9nHyDurhFmbLKwnfe7HjLqk7uT7tjls8LRaRyp0U99Tpymcvl+Lw7
u47GVifFYCwT1/WEl+y+iRRRBR8zfJT6NzdUlPETpQY9p0jKyr9rWWCUTtnauDBB
sH9hAXFp/1lPFyQ/DTYaUBAUX0hOYYOiaSy3y2OmFGyWnGYkEX/C58xsmHcJyiyB
P4h9jobljb4YvFqLTLLH0bpBCLeQTA2AlK8sxoyJu201+nfCYODqEMABuuO90Tdc
zZ5/uMaSIiM0ez7ZeuVBLYXAby0zZnWb/c+Mn9khNvafzzIqHdYQ4d1MapLP58AC
82+ilYUDxS1sNKFxRy+gPYQtrM/ebcmsMYfUttUmGVJmF+zoe92Y6m8ocX1G2/6P
kafnRR6cTyviAfUdS/8ZqDRanoi7rKIjK/yUM83ZosS7FzkunlnzE/jhGL8pIwUF
qqRoUOnrNqYstoF9FYgSu0pXw4AdOJj8RVcugZEPRSrA7ddJ1+sY3RLpVKHdTrpm
hzFvdz/KKc3Wohh57Hln6JaqStfHeyAkGXFZyZe73+jMWDNorYCaMnSDHmK+Xdma
QNfuunGQcZq4d4h69zG5cUphae89Q4qICAOJxI0VjE5iLCBy1ImsemaVgQjGgDix
DdcNmPEaGnOGC28UdhTdc2YovWME0AsTAwUxKJIC5qeaiHG4xOulIV5s4JDOKzNT
Gml+whYxllbHU5fjFhU9K8oa6tPZ/OmJBWvfElnezeFGmGBxC4+c2NWjM5lYmOXX
AesYWgb+GiyDuKq6qikEdsk/VhBiZFmOWcfhMoATBqTpuJFlKfn9aCRmR1tVzv9e
ISqFvpIQiVvIg1gq4I8ZdGhcRnRPTDjRmd+pt0ZkxTpXdsxyZdrJwcd2z9MVqsyO
qasJtDJ0Ynzh3xyVR4+M4JFzJIqXvuUXG3rRsk4/ZvjQm5RxvMu7QpUG1pG1zGF5
fD3ReiSWov/pyhUzbZ7h+TvfAoN6TsYfynCvS2TkqG0PMlDLMZuPmgAk7kB461J1
c5R/K2txpx0Zz4hvQNLqW8NzD5a/2j6AsRjsTpNgg7+K4JcdisPnCYvOruxhzTac
UBQ28KVW/9yQis36SgGrgWxyXpzq0w9mgLIFYsxNvYZQdgBGMb4y0+an0EAdSbK4
NKVCgphv4lrH+xmCj65tAKGRWkIdsiO0pVQC6ogZU0tupd5Wvt62pUh3yQTYbMM+
kTQ7Oja9jTKep5FhlnPrwFBlNYQIag+zDuJbGTWOFip6TnPspzpFf5VJ41zCI2Ez
CvjsG5SYcOwm4Ekj9aS9Ja7y5VM+N1OVRSPIDYkZc+QUc+2Z+s4Ss7ccaJx11tOo
g3Ztxg5CTA1928Ywlc8bXr3PREO6YEap1qmSVKR8w0ZeM3TXQygy8oYXc5xvTCeI
wf5KgPzpL8Q5dZ4PIVqYo9fHfCC2bLVtyOKs1gK+UC4YCWfYOXV/veV3rdAlNt1T
CZGzlMasi7DT5x5vbMGQJ+BZFxzq7u00mMl6Ck+sR5pYoq1OxLwUAQJMAlGSug4e
rsKJomgnKK4XhT10MLKUEl8mzMdz0Mob6GOjlZShJV+3BksPyeiwZaaejX6mBtDz
6vDHDWCHYQLBKoSNJQh4da2ohXinF43yEurD+eINuZkOfWQk96BqxWRMysiv/Nmi
j8rg6s/VsMpvY0wqBxsjGeMQ8vqQgB9hTXiNseNO6H5D8oVPhdzSkCwC6t7Qiu/f
eMifpfleOWrNNF7mYYb6Y0DJ5khiXriCeGgTnS1OKZcFsGUmHCpYJMQ+wJW+Lz/Y
cawsDL80VlNl4fcg61EZ2FqjFrkl/7oE3BNy31t7aNsiNzVuh3epFbTylv/0O0Eh
i1IG2x6YgR369HHbX7uwwk1UrGnPvYHj+BFxMbFzBa8krXvzH3qhRNHrYcPIzJmS
5lG1ou1HSnfBfBDYV2ewxO0fl056BeT1xtL4EReiyKTC2L+fRAbJ6V5mb/TfwUeR
B5/Djx+V2aU457dG//3LMq3eMI97rQqJLsgZXqeSb+lK0Pn5XWTicYp4A7nZB3xM
fQOi6gWkH3bwfyfrIoYyoAaEB2dfpU9LoO+/UBLbVYUpqdgh/oDsUGZ9sCs98ZGb
SPdQ6vwl71AlDoaOTnteBzkzphnzZ8X8ba1CSg2f6/erUG3yusUjTR0EjyzOUTOK
gYcqJnBiKJE0bPMTzi2dQULtKbBMq0aL8v8Zqabpy4cT+WqPNe4x/JCBngMmb4RH
H3JDl1l8zfmqXHrp19a7/84Ga4I5J2wgZExZ9zMSyJz2VzcZl2mWUQjib1CJ/YC3
PAsNf/0JdCyenJX4I3kKUXqvbSnqf9kg5Cogp0im8pcyWuAYWOo2xHbzJ6OZWwfu
sMvY8b7O2hlcw66PzqTQWP3117l9qn8DSD9CaisRZXKxFtdBOPlTUAYGVq/O9lbd
+2STgmApibDf0wMHSMFlS5HUJu2t9ngxSV2C79J3tWDn7axoPV2KSCxTKp+97bRf
itwAm4/SgKU9LDQrMArlPKspU1VWK4wZJemr0poR2PWah9Vxt+esVJY2A2RzDw2K
XqmYAccno2wcR5UwyawZgKS4BD2ijwehiyWHzCBT+3DbPjfmdOYqS4it3vqhW/dz
OP823AUGZqUtniSggCU67XsqG+hBXE5fBTDa6XqmlXsV+rJb3ZAp6KkHr9nYK8FO
Tr4fHH1kk/tu8Nvhc5FkeRp2439ScPAV/CycGYhy5I+rBXsASP0hoyA5RJKcGVrt
repNGvs6LinWWruxO44szaD21xiLKYlULX9atNUgd7BjinWk7lKHFOAd6i4cGWwW
WZ3s1PyI1OdxbhyQP35jzqpOf/5KBL0tYL5RActxz/v/R4ojhsK7IOFPt/JmaIte
UigopjdP2LgEWhd06jU/0wrdE3iSam2gBd8Qa/peggsKtS7izK8jO88dYRJ0hyZP
OcowxvF9kUD8iJ1fgqfeSOu+gifC7jVUkxR/KU/e2Bu+GbED8LfYKDpZnWdsOyl4
bWJ84Q/B+d577a25HVjPeC+5d3+MGZYSLhB9byjl+1FXmuGs+d8+KX51/4ICEB84
rYQovBfWFmNZm2s50m77fMo8rHkJSgfn9zaika6v4VTTDv18v2UMTRjYWpeOquD9
H5IsxPkguWnrIXthR4MpsGPtHG55NjtrMoqhUGutojiOkOuykRh5fKh+n6MJ5l/x
2IMIM9aRwoP6Qc1BLeSZPjXCWHtGGMikB3i/BJpPF1j459lm8V10sNAtmQak7dgo
aB6SU1El1DUzwpodPhWccJEuo+d2OkPY8Hqk6h4K5/qdHDmQqq6Am5LNGjgvmG2l
9M7p+kuBz0fgEtiqchoCWVm/lMSnWQU5pV0OPGSsnQFmMqmdLRyvcq6GLJGYg+It
dvDkuEUPnE6PBVbkMERSyAYRd5bn6pbM9fMX/q+MwLIsUdVGFJDA3hGptCiwMkwT
0n4/0tsU8RAX2amtSxoBJ9uBXL9Y/Hp8eIbjgOLfmNn+zMwccCHFzycn2UmchbdN
jysSkUX7d0r2Dw98p4FgPIvCTdaZNRD9aQac/C740uyxVrSLBSBlaBHfo9dd3xPP
NO2p6sF0cS5SY6XwbmbjPg+RFpTjqSyjkdJf9pWO7zR/Ow1Eg8MI9gHEE8eIKzDA
iiPNDsXzlGjSuv1jGP8i5FnHd7Io//38//8oknWvDixwxPV1sn2keymHZratvuGN
eNewyU7rLLikpsqoJUzJNUojtZ4171BpZMti9qgipGv/1SVHo5j7/wUek7AklYz3
Z67zxCwv5aR3LuQLi2hI2VLoGfmOFVk9NITDu7v0bYa0HeFJnaurN0OgBlMjZKTY
AilNMH7qSSJoNnY0eafLivQ4uJQP1UnUX0VqVsNKkT8851k6x0h0NOuRZ0fY9D80
no/kmbKpJxVWFO/aswkfZBO8tlTN0tM8SVjhDh8iDPU8vDfZGAZ4q7rP1933cYJ6
yStfjfLVfxPk0Nfj62GgRjRtHgOj+n/HACZnpWEA0XntYIldOd87Yg0eYnHGtGdk
j/MXSDTekEfJAS8CeLQNcF9498rv9PISCpTaI+3cUF0yA6xAEJ389f3XhIakr4Mu
s7hcVW9X2bv/Zw+xKpTffspKrsPevBPi64xAVcwgyYTNVATjUkKp1eduQ8rJehUa
YMxwM/287Rp39i+u8QmxpH+iNR1rEwLwYI/Y9Vdq9GQgBhJt/gElckEDUIB1NoVu
/ewg8/MsS+Hcw8m5XBC/Q/xBd7MSu6hn3HzvPi8q8n2FRnk1Kd5f/bhq9PcoI7p2
VAAIIOxMF+TuE67s9WkNFZdelGSCQ+KpT0+MmptY2ID7fsyWIORCipLhekveyUml
uv7mi3BpYpwQIxfMqDNmE6oL3vtQh7Q6wYrMw+anGuWN8w9Q9W45FIB2BBn+RsRM
7B3ZGwCjWK7+NknxV4Bm6xoDNGvXAyAimmg8Lpt0qLCzEIpAp/GTetUU7kgNKD2A
NBj/ZvggQJuKthHqK87iM2zr9xcjyPvClBo/26Nl/XecrHyFx20YfROuUcsH4L/f
U7L94rmOeJPkxHf3b9wsIPptkwXDlyAXcvdJqBIns737l2XeocfnPxM1+yqxH3Bx
bB5UQdmq0gIlHe3RtEEEzYZS4odPzk6Xx2Dq1mQRyjDiQ3s9AA37Dj0Z7PwYvk5F
Y1Y67ugb416uGQSBDJCz1edGnrbIdSxrPzxfo5aKyJB1PivTLe/awI9tNk0/7ir2
m6wtYeXl/hSVovSWVF8loTn52SVfCTvoFLRX5g4qanZIcJ2dCCXjz8EEx1P+M7M6
idAgMkPPqTsue5JUBqZkh2YsPK13rpvPEucq8WMPC6AUiAnhAjtAqkjSb1xcAh5D
rZoOpPRTX1YVawZ+EDejtBLBgjXCFNysaZPZDTliRgWHkPqucZFlbaHBUf64mCSg
ViPqPD7ddgqqx6IJbvCnYvHsKQKk9694B2jaMmOJBeTrH4kisnBT1WMn+BIZlXfZ
cReo1KOwoddZ9IH5vC2lG3miwxLIRIN0he48DZ1FwfCJ581+0vl8boHd8fFH8hsD
7hcmMCsY0ODNDdoo3vpDx/dooMK3Ogtvb8qpK+JW/9v5QRpuxhg+Isc7z3SSW0PV
DauO6ujDlzb+ZjuFSt1Rg/WEnbfIsFc8PE1JsrwTL28JISfsJYUl+OyDPNqiudx+
k8l3o7KuYVZSWMwJl7bZxaGcXwRyATRk7mcJzQJheMxmWaMM+2SbPEdz/Zm8Dgfz
dSfUlFKsRNwwCgvyLyCJqWsqZ6P6SOYJw1QkRtxXkAy65p87c3zf3jndnPOMSH9B
EN6Vj+9LPIPuasuWvRrKDtv1iZXmpjI07eVLXQZNsdT+gh/vOBwkVMwOnb9Cmdh+
/c/6e8JMg6jvqj236bI3mSYGp2wg2P0LUveNTNuNxkIyqIuFBcmnRqhmAo1jgESD
VNni054qX4eUx4RlWSZrfTEvBioOeGr9+E4fLDrOZ2anY5ZO5xuLxGnKhhePffNo
0EUlxvGPRpwiMpH9kyXvZFv+C3/qFccuf1/jua9n10w/t39mT5kZr1MQvIKliNMq
4xInS53x87PXv59lu61dareYdL1efAc1DsYxVtBEcci8BDMQNvaqmtRJLNRwO0ns
RB0ULWMBD04zGP6NYuTjPQSOgDdAhQU+ylt8udwAHAplEnArR2JgfhlcSBoVhDVM
uiOY0XSQvcNlHpxkTzhc3pQeK7Wd3fUz/E4udSeMFL90UtPGV0qhXbdFzwQ7ExA/
CxBdZqwPthAAgB0eIeYB20IxeU8WaoPV6yQa5dSJpmJg7uJDplKXltwlu1H/VROu
zgm2jjHBSiShSe8Ia+U3KE3hSBbOxqXulsf8hk5T+Bu/6EXrJYzAtajz5B+TRGtd
qk95pp+zhzNsXjGX0cLbNFxZLdCsFjjE5h3KPNKeRToX8oujxFABYcaIBVBOExvQ
xrKLdjB8LEWSNFL7PAk9qsXtrZdpqS1gWnAy8Wu7LikcZC1NhZFruzuEi8OP2epF
fDIZlfyy1hBVJwvXf1rRwfNN6qXKffg70pXsEKLykvDZhzEuo01Qx1PnWHhKGgHf
NVP2cjMZMgxOrBYfe71hW4XH0q8zX5CveP9eVsJwHjC6R8bxu0SAEgFmntPvxO7S
1txj2nrZIipwUDTj2Gw8BE0p+iwahfIoy5zVx5uFBRFysxrsPFAVtQcxFNaVg/Hi
86ZUCIcxzTXRKayMdkTrJSZvFrgFQBs28hfjdvor36lYGZwEe7JbTwadfL/E/3+k
5H7d2mAsd4CTFiKru8iZRgZdQOu9J4Z5zir6rZEXj6Oo8eqi58hP0x8FlTJpnnmG
sAIjlZ3GlCUrSPwdMIOodKhw2Rq9Jy0bL2ZyzFygUD2lScKd8Z9SmcBiJldRxZgk
tK9xMASlCcOwmenOrZx5EGXdihKxJJX7Q1gTjMy3LcpcivhDdnNYspHWKnJRpCG3
QliCUXMWF1HOdAiyCHtPiuRVLJdhjPop4xZsgvhQJN7PLaFLE5CXQDvdzkJH3LOe
1gaCD28GmNZ4pkN+LKgspkhxFSHdeHjSo5XH+ie1L0MHvXOYEiha7uDJNlpeNgfq
NNMaey3qPS2F8Ha7i/jbFDKacLJC1Ntc5HdVyiIuzwUnxWeBzak1iPwuaoBEMvJT
zeug7TyxmHjfmfMWOuKuLrb9aTWeVP22hvdp9zrQbrbT0PDbsOY2H0j6XV4XX8T+
b/39JJvdbA65f4MzeloTorj/mlcVFy+FOtEOvKiXT8475ITvLwLSgWfhJ8GJo+2p
r6m8xUXSFgBB4lgJokMfxh6q9Dtk4IRWB//hMWmhYegJ3nCQNg4Ydg8JR6vgElDR
rRNNB3oMWOZT+Lv4qPCpJZsxxpGMrfxc+5O2Jw2C/m+xInI2VAqNg2t5qEnq5Ssi
IHktpV3Lsvtv7GaoQoYUCAZX5zhwfPXcuhqSfyA8kip/j/iYuPB45JwyART9ikN3
aQ2yo5JqhNNdPdq9O97IbixZsJ/eog2u9rq4/VoaXqd6Ko/lqi5AxIrCeIY9hkT9
S8UXWk+hkpf8E8Hr50/lByWWcKy/boXEL440p9D4AFbg1Bl0Qwv3z4TOTPOSPe41
7O0e8j30X8X7JMqCni3gThi/MoAfIwBJv2+0DfvaFDNUB6WkeuU0usmqdxuOT+RD
qHJ6WJ4vSyAYZsndeCWa1kl/uw2V4T7DP2eWUez/8MIPVo5Bj4PcVBjI0AH+m0CO
H6kDmfI3l/afB7Xh8rKB6KSHrlPbuE9ebIvOLdd+n+5/YQGB1fbOrQL500zOkgji
m2Rz1dlIGvCEj6r971FJdTDWJ1B0QFDg+QLrHMD4wtU/Ro0PNCZol4w1163Xvk6/
tYIknjMKDGj+ledEPMYpSc77vmu2kGKqIk8AP11BgCWnosqy4/dmxITkF6RMixmi
o7gy5ULeMbQmq8MXdv4zw9eJVYDGuKVJ8F5oINtW9PMmfA4WxFnLuzL2Eob6zuXZ
e6Pa58F4KBcNS5r721jlxPlGVakRS9fbRD7QV3fQkd+EyTq1GGS3mwGQP0AvZGKI
sC5rbKkAHPoQHK8/TFUJD0Nx3kOivDEmttrSY6apneZN9uszhBFVGi1HwoVnQqTu
MV6UHrXpcq8XZ77VHS4XCMne538ZOxI+GruVdQjp0KOPK1999O3HOwmrcecS/JhO
Zq9JCUbOxoq/EUyZqlDfjeUBfsY9htch08kfGExClkhL0B7ZQWhBnO51JkS64//C
YeE2UYc4C0yWy7XgzmFJyIfR7OlquqxJo2X/p7PGi6hUopP/VRYbSNZ0tSzQPOQh
ElexlEWdNncoIOC6nzUAdPavQeKAKeA7rKFFpRQXa7+CinwevCoRBPOp7nfoHbA3
xvrbUjVLEP5r43rPje9AY69ClyrRA6z5v+ZJt/NaqIWP/ergyHhU/6wN+0dovg5g
fE1tniNe0dCdtzjNHLoeIrJXpn+qPduxdE6HTAIhRF1dtvcKd83GNAB4IUO85zHP
ENjR2bYTufYLqgewNRS5ujobhYU2DCtGimIzvI8HLcSKhLFfpFYfSvskS/WhvUFL
e4b/e6EArr1OvkxlsT2rPwmjbugfGUWSzJKfa4gKpJS3EEpJPw2rpj1ozNeH7+3D
VygdZ0YUXmGUuQj3QmehPkbR5L40ydJ7/vBV2oCt2OUbqu/Bw04EYiVs72LT+HIS
RNR2O60TvSBMXFX9OfGIO4mr7lijd5husUVhUxlws0hnK9Au5SMbGVQFqXYnBoxq
K+baNDRjFW4rTTC/OwG2do19ryXEEs0EPxp7x20uaK8T44PlwEmXyFQKTj+yuY1X
9ufUL0abNAWIaSs01xelWFCUEykBxyE8yb0KWSd+VLZCstHdTw5AIg/OxQyXU1sy
iY0/J0roY7luV5BI0TeYrd1NPIDxSO9eAELYG4s2yrIPuYQ90IwJe6fkcjvKhPxr
Jk27w3CL5zmEgWGun4GROTZgeBHNOcWvsnNdSQMcA/d2BDhjd0jJ6JVuhYZYku5T
w22iMIggAwe/c+mmxC+y4bWwSzeTJBrNDDj+oV6kKCdls43xNXsEFZGuw7AD076R
k4tvNSPglUZ2pRIcpqxNvL2EQ3hHdHWhD7gBFUALDzteujtQ3NDB2U0uSZDafJCG
3gM8Lg6juDaDcktL8VfXg3+5dVIJvaNnLX+Q7xFgZGDrYKCEkmLChBhyntjDjxkJ
04lkgGjGGF+AuUeP1ZlvrSqZsPQ9gdj8m1t0kLT6spOQocySLXw/hZug3u3GQHOH
ncPonKvV/V5iw68S5iGXUMqpfBxglI1qiekrnqdd0E3wUdhmN2HvkAylVWyf0axH
mtLDGWsO9ZFMs1jcVe2heV6Du10uDBn75suXWMjb60Z8JdM/+onKuKsWZmlklqaI
ydudkTRzKuhcdhY5RnoMYCkLHHDww7zu3XhtLfq5AiP+HS5RXVHhttEPGUZ8ld3d
ivDCOgRD5373pdKTtSa5FcD9ySxs5aHgsBTTpPLYMwXWdyCsMosedPqkKzEiNZqe
UjCYQTxNC4r8c4xC2kwrm025pOtNrgRWGCI1vBTeNXmhYDwdhqHRoLdR9gG0E7uv
tM1qT/guu8LCbqYjKKYvvQ1+y4ialF7Twwe153tWe8vb55Fn61ANBsrv/Ao623fq
7pvGQzPqilShc0hD+P7MGwtcXOqTd1Trxq8fvJ91oo3RvJEbW2alNxfS0srB8iKu
CdszO22ClePTSMr+6hXd7UM0EBgVKU8nq/xZIZZGsdGxXInWpeMnvdnVBWhnKkwO
Ojhg0t3MH3G6cZuR9WxZrxGJHK/rlNP/ssWMiGzUtKBvFhjdf6qR8heItmeTluAN
y0z968amZbbWlhun/6khQAMHyVSgSMimdj3VPrcI5QLphqfpFyWPjcoOlAWTO3wN
DyUf2ThjnT0kDfq68o6R3aqFmoAgpAO3xEwJQli7pSVp0dAVPWx7s9HX9kj10qte
hvEf5fDDq32LnqJxzEKiV6ByQtg4w67XjYghiIQBKKLM4FpbYLIp00Psw818BhPC
xNfm9PnrGk6Fkdvzo7veX61oqJsO5YAefbcWwSageVq2VpdhKG74QtUpDv35Mhub
T+1yjkp0M7ayCg941SAPfgxgTx1pCRERuaKklMnRc+FjhG7gmLfYob6tIviE6teu
GTfnfdFFNZRzBivNe3oku7mSZwTAGltocofA47Bs7Hn6+V5ma+VM81aSWNHOPewl
+/tXD24h8d64vN/KAQMMTmUGjm0mjGXAf1kIfOjBy8YN2uRX9T9HGGTOgrpHtK3d
+GNPkVHc/c5nI8qizuitGc6qONJCxOcTWk4T3yensyAEy8F2PVDcZUGl/UmtSTYc
mBhWr+8rpYtyJsJFhljaAyCdJjxXcSIe2KGB/wp7+Cj0KPN11r2wwvmikthPid/O
RU/jEQ0Vtz3qDjL8S2KC21M3s/wkInnoS5dxgcNbf4RQ6qaotAhSYp7S9wnHI/dK
vBVECbrABH11gCLlrHi0GtEZb5vpspRuqinszBeOhZ2YJU+Kbs6MXFCBdWhG/W7P
mHtiTotEzYx+0pyWcKiMl1b1n9sh7Swh0Mn8g8XKm0TXRtx6K1MSEPEvgwpAF+7l
piMCBRouVBPFdgLJVycB4n5bdiUxHIjDjvjsPRABgvO9D+ZpbOLUVZFvN/S/lxwN
eahHmEuhSwpOTLxnhHN4ERBxkIkD4IizjnoUg0RSRwmBPMHyrvAobwLF98i9t4Ws
xYk+fW8lLp7MRCAPtgS8bEPFJCWxybvud0rNJO7A8JgB85P4ERVN6BJOJg3DPTdd
+9anChD++68a+yjNxdYBg71KYb90xwggp0zqJdln6XUTz/Ym3+Isal08F4Vqulmz
wNGYUqnhye8Zml6FKxsYC4rYd2bJlWegUBEbpUci8t+oj0MWMqojZhHrWliD93Nl
IzggLh91UoVGg76M0MW5FUqlxw4dVmqFwp6Cdm4UyqSANyj1LjnB8nV52KFYn9Tw
XaYivPhsIiCcdMKM5TTxr0QA56ZmXONhOytbO7RD1r5EFESt6f7VQ0YY4xSDNjFI
137Lj+FuPqJXM5f5an35SMReXpygXrAnKnVVCwYtGUatnI/af1tK4+5GKMftqmNv
w6FwyNhRcQBFFipQQE0fJhzgWGtN4IRUFSGt4J2G15430tuqWpRGCVc6ogX59XVx
oBq7SpmzznK0jx45RmYLAW2pL4rLs41WvOC1+Su1YfhvALDGvwydT6Bs/w7nrTD/
pRYAteejJxE2R3SWQ+Lie/6b08Gwl7WqXZDozBttI+F36KqcxjjAuyGrJH46Cs8X
X4z69X9e5P1MRyVgIhFn43DIwJICR74SQ/00/uy5aDbCvxXDcBD+vtMgMVC2fwM0
4wcTNTCg/q/glNEvWKVA1W5u4oq7hWbHynqrUfcm9AE+3MzH2VzHaANJQDOcby/y
7xuJ0OtX5Yg0BWHx1t6EShgncnQTFv9i+o1AB7bFmSQfdtwlLTBd8H4JxSXRa/XL
nefHRGniJ31wVsvxdKKjL6xNuUGJxEe44foQFl7mbyiEdNiqtASFZGkeV33GBtU4
YQ2qO1iM/TzEIICb84h+ORpyCAHIqgUwyfzm6ZlqoTltAGPyrQotGSAzqgjP3EAE
t8RB3hAsqzg4dfgVHsBz5B2RW4muS9L6b7UgugTIojHdZkqsw1DCBE92/iUQoTlI
2D17A023zn2xclu2k06xK3R4FmKEFr6H5m6LKUwSKquuZVdEKUcp0Qmiclb7UF8q
/rT7dsqjhyG4VYQIhDY6W1GaJnWDsJGVk+6/GTx5KXOLl5ohiW51ut0BMFkRgyRU
MYEaqovZxDlRUruTL5NywDxqvCTcJ6HyicZT3S6oYMErFUbiXFzoKIyfG7ZpD5H6
R/HUNsBBpH2KTGgIBNMGgi+wfZmbowlwh7SBGkwxxhT01levzW2MSBoclZXat3dy
V7hkjDh994y/8vPmqTlGl8+1HlHLUKIM37ngIPX33IYPwQ354pdF+q2WXYoJwr4a
AhGyUS2eDEkoyqlZVZvgozCOmRnVjKh9Pnk75HWCSyJznqmmjdM/3yRrxc6YIYiN
i8JSfnufreIF/HSQqK2wipBZ2MdSuSDnA0wCPT2xPxwpAGUUA/qUJ/lZJxT+X016
I/A/76ZCd1Aft2hT24PheJPM76a2DwbhjWiBeUmF629jgOH1KK0VU1F3ZvQIrDFC
R/JIWfHhZ2UltZHWSxxgQtfQmiRfTZFZbhsHdzoBSDhR8pC0NHisNO2ot4USiKMx
U03rrqCw8RqZZ1k9LTaakWXz2mP7b4AuWtVkhU514miPb+sWemKXKNiB+pT4X/pM
zhyR4Q1OyiKTWo+inthHSLZHzsO2bEGF9w8Ir1zwje0Zia4KMmt8cbPGIumXUZCf
+6E9oz4Wo/nVbQzguy0Ln4FGpUnby3I3e+tc1/vuJ1zoyxGzJPGFZpSB0nBD1hRh
HA0cMKNba//CzDHhOqiL7YoOW43PTTmyClWhRaukIbxmWiHp7dN5qD5sGIg8fVHt
II6xuqysshv9IRM3zNArugBkyq/0GtssKBZ/6vrLlaKzomqlPIetERodh3AjNytk
dfD40EV+xDCYTKDmW3G/6/wE6hkrKlynKJKQW16itjMu26kxIM2UbarIOCd8a6Ug
E/UlDRi/9V1sTsa3jP9HLYHUeiSSwvY6YPjruZsco5TcQzMtjE8gA4JSPdVNALPf
HHzu+Aoeg3nIHaAB9vr7ywziBPPm3IL4UR47FdXPGHXubePBiQPUCn/mLbnSZAcm
i6qblOuyO2Wct2ypYVwMe/VWJShZq/2hbjZm0TD+cZRNgHFUNo1v6MSosI3r3Wmj
uxRO20v2kdiwB5xgphcsfzkJkkmTAve+sIGwaGEW9L2TplnaxLKEERQtIbpsLTXX
83yBu0Oi48QOb5qhXkN5f8LVrnp50ubq+FqMs1ijUMTWKrdBkGfY3TBdk0uRiZ0A
cOBNIU3FUfjHXRjy2/MU4AdlW5s+du4vsZcfKSe5++UL9J1qtdBzZFE5WdrmUhyR
NPYaVeV1t4yLOtBmtv3BBjoEh0GOPZFASCczIj5qy8irsvPA9IWQq8u7EZcanSyt
M2VoQM9QMkWBDZiUsh9LTr0+5RxKLdQCZBbPvZvq0Ex49NsUA1ksaVod+GaeO4a3
Mzptj8zTGhFgXHzXW6snopzZLtQtIh4GOhpUPhzv0z3JHaQjBsTEl+eTbNRHnk/w
oLKsGj93btNEs78wy1XItoRSUzKQlSvK1ShDsDV8lQkjysFcNjN9O5Qdc+nfTGAk
0uMpH1RaaVwf8r6ixfsi53D4RF4lZUIFMmY4F80mtwVxmibcqYK4eUWLPLe4aZey
EUTfTD5KaoO6KE7S0shR2mUP0vAiMfj9OipDlEJmKhm1PUAHaRS1YwKvpgwv8eJl
IcabdRHx0G+C19p4xX+q1qi1ahzocOWscgXORWInMu9tNQPy/1lYyud2SXC0qWwz
Mp3HMvEvl1gDEcD02Xon+4GbpTjhMHcq75xA/yJW8nRik1rYjIfRTAgYhSXoSXik
/UqSxgWZLycH5Nm0knyTCMqCkHvFlx8/aA+TO8zOSB2Qu70XOFwleoznVmeSIWhV
udErIW28OXCexPBQymJbam5T35sXsgJysXvjfkZEwotMj8aXO7CynNRqV0ttNOGI
sJ8ryoKAz/nf9S4bNK0GksIQpEZe5z4LTNd2RS3xkIp65y60T1cm0C9cSntYGDgn
cnOh3AWwG7IncVIBgtdRNizvOZKmx6oQyaxgVXYOb2tpAUxJYxyw/gg1P2MHWmbA
Y+5YIq7wj/Y0Gezbf9FIlDAaQnZWEkgzeJjqDfyxZSzkZYmMgoAV3x4FO38aBbHm
NUZGaciXuLJuoSZv19DJCZWixMIUoy0UAIccAnabqk7hDYoMzf34KrR08I409kac
WuIXOYIjr3dT4EesCndnbAH68t7NKuF6IsNz93qdQRKaf59afk7oCdBdgVHUAVE8
nRJaIGCdUbnw8bc76WFELbjDDEdq53qNpXJnbhhoha9I8BLWg/NwQGjfRcn2PhhA
+iiFiFmVTTuX0I139fjcAhujIC1R1A5e+T3uARslxElT0MRCU4tSyMLuwWCeAo8J
KsV5l2dO2phrHCIhQ9bE1EE7qpvEMGUgmyrJo9MXQqTFpNa9CEUeNP8/v+jKvX5O
tFZ1zHLS52uS+93XjDWWlCTFr2yHjTDa6wQfPlyJ12FOL6IF7c4/NaaOdcKNW21G
n5yD9K89StXxhShsnW+NsUtprg2K9sPb42I6OpFqE/LjcVIP3AT2+y3umFZ/90ET
9Bn3lkv7YyKfFGn6MfWz6iyGPfOauuad1eiyL+aFvPpRsWskBvTVLhbBtuuKfbdJ
ePvGAzYi+Udo2ISwaiqJS/rt/JhgfOoEezpn0R8Y+docNofGoygyYen4zQesP4/7
efPFc0DT3P/I9fGbyDy5N1U1c3hSw+8HMM4+Pv1fjhVC65FmHa4D1cGo+6HkAj5U
ABxGp2/myQ0wjnBR93XRUVMrsh+BkwE3z1VLeK3nprRNXueMnyAKxKTYPNaXlAip
fl8eI8CCq80f37VQ5ucW/wHkinZQ60fhiJ/4LDCEYDqLio8h3cHAcYh7H23QjViv
wwj8ISV07Pv/zFqeG5F4eCW5T3LQV61M7YD9bpkKrfkQtfQAOrZCXcEFDkAdYksz
Ojn0D3X5NViFOsgyVE4xDXnJobSjVwT9V96GxwKzTCJ1bK445Lx/eyVfZtm6LLlR
Shj78WJeaReORspTivq1Sxy1zzggui6+EzkXL52KRBVtIi7Yimg8AJK2cEqf0DuC
VYVpUNxVL0IJTLHLAAehigWTaO9e31j7zmhxKFIjDLHqBNfmtT9aY9FYcnTGt2zc
6+orw77vZuIbX21fuPvaX4K12F2yaszdH2U6iDO0N/d83A5rxxICUm1w4e5+TSzD
iouqjWYXG0FjZG1Ww2uEOOHG/AhDv3ryh2qKdYf0mUsLAu0Sul/7WOXwiI/QJGtb
hPnlU+Eh1Z0a+AyBLEgHusmejnWK7Z7eK342Bzl9n9MqtZ2dYF+vU2RA1vnpJDi4
2uSJorFJG7NLxiVnHwgBaIiPQD5p2+ExR+s5/erdrqOz+rXV7Xxx3Qr7HTICGjx1
RZxbuTF/Kuo6ZS5b1z5SfeDd0OeVtFp3/4Wn9aiKkuXFT0Mw5zg8L+KDBrFvj+8D
pfIYDZBfO0tFsYlpNCcKKpF+4IeHlzdfBJbiQwkmNE+342p2qbrcyUpICal/A5eT
1n2GydQiN1f9/SR6YT+zipJddu8RZJ403EKXibhTeiP+SPUw2UWE6SqwF6tHf8r5
pa1S56iRp8u7AjAifseeedjSJ8YA4iVA4TwWczgxVUmQ35OCpqDGq/8UQRCdm0iL
FXcgOPRVpNIlu/oRE1soOcs8XneWkpHd5MbtlodhYi7gU9ECJSayIiqtubU02pss
sKBhzRRfX80Kp9CmtfLIcXwwF+r4QNfHE13Dz2DT/5pTNwtckG4h45uOzw8oImyl
KI+mGJf0mNL6q2HfbQDMZsQWxZfg7lh6H90205zKdV+AARlFOCA/fJt6QYnxcHga
o4RAJr2PJ3PrINc5MJVdp9R4o4OG9i0+ZKXk/opsrgLLcmEFKvRUrX3S76zTR3GY
SJN7+hGO03YyCXSKVLPl6Vzxw5SHpvjUbWAoSksRxnQ7EoiuL1IPnr/KoQgPsbej
2P9GsKoKQZoNQHXl70A3sxhNwt51Z4P6J+8/7ajRUJOrDRaPnAOmVP4/lUpJle4a
ItC57IbIX6RArSzWYIuU1yuztupIqGGGaG2xKWdqz1HeXQ0L0pMLRFRwadv5IPkw
Sk1/j8MAaBhXYaLTLGjG9gJlppaIqmjAc7ETGdQcoHGRD/VNQfPds0lVEObgUyhy
D6a4g3PRUQQCBsXmBMvmBXw60iYdok0LdxVc5bQGQg3PDwezbPI3IIfbtYUv57YG
jbGZdbIMDFA1WqZkaK0m97NmEBEUvrCEJHgxiQHU2QGY+jf9p7OKQjvcxYphZgQB
v4D6nHE7M9dFij8dKjnw+dw3DUh5NCbJNXbIeUGSuP5fj/TzCyXfYSGbXYDEzn62
wU2WwtCSZLQYTqSDi13WPLnAzOo1VakvzvmIrsENROWB3wqQ9XkadtqClCA5KOUo
UmnrJr37YMR1Ab3h6DxX8SRKEdQ9jvsSqlrmDHjazhRPt79Q6MiKPVYg6Jj4tFCj
Da8c8pApuIVhV+w0oVaMADmRWzHR2Rt6tFUmD7AJJaIXlgc7q/m+9Zk+m+qZ5+r/
fAnP36kmX7IqgvrveISgiGxxx5Ayphms7YFoQljtKOWEziXnb0uQI+ZXQnArQmuL
GtETeCmeO/VVZsquf9Zj6GB+W7Me2dIO+U8OVRntb9JXo3o+ikKz7i9eXiXT5ktv
WE5C++dWWzOPPTMPHk38iReCCSMuuETgUPB4aJFEkUJAQPuAWhvB7GC+mUqUokb6
4TTh8waG165iA/SQZm7mmgFWyal0mddPXMKgQ3fboz2qUuuvSA1ypXLEWqxNMZEP
xx5euQsKu76NqnK/wN+13mFQJhEg5PVIEu+ujBBaifsAD0WKWCwFtn3qTHuyPDzO
k8dCpOIQCyOh40JSLbdcJY6v/7Bd6WOTG0KhyOsg8Da2/yaN3ElreZS4CdawobO4
VBKoMB9R7RK7xLRwTpYMkgtUtplnZRtw2VHSs0bCxEuooJuRZNFFWiTKU1ApIPgn
dv9pWaJekzZvOLXi7ktQTj6KuBmgnisjaRBYMK/+4DDQZfDX0znnmIilE/+WDgJn
m05DkaHId47muFRBaXPOVO3X9u8NwGaWAauHhW1BNLrno3aXrPFGa7s22VEUyg/y
zi9u3EyBkj3dWXlj9qDa5KIDFoiHjFEJax0sfNlk+b0QuWhGqpalAGjUuoH7D3f8
AeHoWHzY1z2SkMEsVKikKQho15MwWKlDS3s4bexmyjkfb66sSdZGO+xckvRqKaRn
BsQ5g54UJe7T91T7lodqmnXUmBf5iOXUP9SzZgmfIc+ZvE21ygCVABG3hN0m+kNO
ocxzdoX6+VBs0o3sZAg4VZzaC+BbcbWbPWfxbrR4hI+m4WN7DslnB2p9wvXSAfnX
X8WIVPKfbjIf0BhXSM4yxpbSHxILP1pkJfwIyj6VaZQmP4aCbPoMSRUvk2ENA276
0HJ97JU7brlObNiiH7/BJWA4QLYPgtdUOr0m5/XM8hYglAAVVfJLT7o6CXi6buMc
6FexFJE1tq7B5+atz2SbqEyEnRIa4H52VebDzltjLroSkQF5fJLnoiJx60AgCXtY
m3cuzkTpgZO35oW8pqFBOuRVBt6wMAaJ58vFKpJWweyEBp1EuXMRhhpubd/z+H3T
HmjvQUiZi8teeax2L0p3luTUW+C7C7XDxOU5Toim3t4IaMwGwBft85eLAXTLSK+s
CK5t8ayYka9L2TAz640Mm1Dgj1mVNF+7NXYYd09fnUCrPvVrDoWvUIlH95f0XZ5h
O/BNeeCM9aAQ3rt5IjdIKmWHaj3Mtp7baFSBuiP4wjXGe7jeAZErKOsR7D5vY8ed
VhcwxQ72+fFA4MM7FF9MshJjUK4tyc+BwPbyKBOJGg8cQs/Mj7MXFtj/w0FqpN8X
CmPCCdCmnIBjtamoXXuX0+jaFe1z8tls58P09Pb3ux4K9oMbfejlIevFmWKdepzl
SAbALXyRdVNXED76y9SYcRRdogh8U6FXD4/vMtK6qeA+M8q+gIrqxz4+Op0Ccysx
xBTinpiGZN9Ez581sGOeZ50ptocryuoya6AmYhggmuw2pOZrsAD23aUkEmRDwYpz
C04KgGUUuZPdV+0Br/0phdD/N9Ltrzk1v0XF7v41osYPwXKAqgluZ6up3E7iFzRj
rUwRag3fUiKzJ5D/kuYjFLgjH0+1wXzr0SiCMk7k9h0640FVVzNyHD4y0olL1eVj
7zBKscgU7Q2wldr1Gw3cxTAbZHDtxa/dHYYn+Wieg4NRlyei5Jr2Lyc7DHdqYGxU
iV+daPN03qNJP23jXsd4RsR9JCps4poU6dJ8nlUHD0IisxWYvw6WCB7q/veQU490
i9MSnPzOLN192izRpRIq8a7DfEkTMsQKknefePZhxheB93mpfP2pEek8WMMIw9iA
GekqqRHfHo9EeOgDUkuDZquLCHkv1iUh420W0j9UUNAyNEooQZOUD34ZiB5W434R
3waN4p1W3sD4gvgtKV8Yb7NXPQYXwzYzI80AwuIdHwHh2zsO2axJi/iIrSJfcK75
jv9dkDxnhN41OC9pFQAHuRP+NAmpu6RnZKZlytlSMlXZn87DiZQZBHbIxRCw3D6a
q4o/LcjT6ILciqGtyiCoMban9SS1jy2fohAWRIp9THINh/5ufsSJ99o4BHTYxMlJ
u9QwRx1HhDctlq6U3a8d/ucmJnQDv4Lt/AjhuK2On4rV6EUgkIrBx5NV/KikRyCk
LFHUeut2VFPo+wWEXgrvbm4GcVhRJgFCy1lswPojisoMqA380c/xx+E+qTg8tivq
GBicjwDaBWs+o+VzsvWMrGK9VmvVc/xYEs021hIj+EMuTL4ZRIPy04wT2ya7kHjM
nF+e7kvTNFc0lllF/Ha3nGw4GgSH7Xmjn78E1nw6608//pdjo3ZujtIe/KBUGA37
DBN9EuZU3GajtXLJX0qy4X4kV1tIF6XefqScPifeGbqnhivB7Dt3RaUZ0BuqywWo
e6VWJT8YAPyEm4jGBywrwZDVBraMzwXgzsCBc4b9tZB5aS25m/9wQQrSUaDqqfyk
CLFnRJOSmXY16WkLNTSnJHo2KWOlVuJ/uO60Sbi5JOLpU3MwuaCZrF1MyGfyjnkR
XecNRN02M3vWWN1gfKkUU1lEj/LO3HEkswu137lMRLoGiuz1vHzzSGOnXCOw/ZL0
TW+UhulZ29Ay073SdTXlq1zrKDE3vdlCgg0KAs4AAnk1hYDkJkP3LYIavvt/oPH3
vYTgzTU7hVPvrlfNLE/OlYCxZZIAaAk12nWE0H+r9fYi+8qGxApqDeQV6hZILS7R
1iRMUIm7iMf4zsvWvejONsxHiN8nD5K2bH3gQfjk9Kl6+S0CJVKuGmY06CENFSXI
UECyit1nr4jTeujmp40geZUpRKOL6WE1L1J8wCbs0pRBKifq9g7JB0UkoqNzLc2g
hjHaZxZDH91oYFWyeeYYx+YCtO9FC/NPHZbHJAeWpHm9Vs7QQImo4mczQHl4wkt7
VfX6xkj4j9ZpYoOeXOOQxR6qOD4o7XzO2i6vUCw65V6WBG0d+oETyzEJ9lsTyxqY
ZDncz/Ln/cqgqiccpl60MT4Xaegx9CB2o7MBw7uNYFYkasLNDgMgCFxLZoVHrn95
cd2PlfaYl6fwk4ORHRBpt7oTgbZRecLmi2RsIYTw8zsok6SvuZQrR9FDZRfeEOdD
uWcKFXUB57JM1QrWODDMzxU49ojemLCidl5JIpmaOKePNwOUENNRhobSjibSaPDt
Wn0RfpYDhVV/u9fobUOAinOoVavT3dBA4Lm+5IHJo9ee8mks8/v5xhNQgCBpUaaM
nlTdMAd8BAiFIVGHbKW2F/VtamPrSl1Zlv9exxTcmP2f/kWtFdct0x+xf21GXBOL
gOcw46jpyIhxLh2iw81HTt5Qex35lkg33tjH5JYtUXOJh5J0WeUrxcAwlMZ6gKX0
XIrbsWklW0UVTY/Fm6Qpw499s0j2tpX1/mEUJPbrrFtrIbcWV/JhVA5HZl+qdRLz
+q3EWD6vqhRM+eFbRnnPuCg4IzKFTAgCVIL6HGSkVbtQ4V7Osh8LTUj5GMzcwrCz
LfwspUDyz5697faBMGVwMu6jdMENwIkyFG4/IXgU1PZe0uTBvbcdHlN2IWo5wcdO
K5MewRtF2XSIFU1Rn8o2UMFJcy0FVfkgwu8xcrBsYlpp7cnOKoS2F+1eg9Os82B7
DUUlzKf/G743YfR6+XL7uIF0xnDV7qUovyJj6+0n6QLjyTFWz/925ITW7t6nOYbL
sfce20zBnfi4RsxXAzUuDWYc2OGQn38QNURYeZQaHVpgqsbxf2R3ZAgDsn6LsXAS
wlJTcb2YFtKclXQqFRxrLf/CNYaENfTUycCGIZEg0BSDzY0JvxEf9GpWcO+DTINs
2iemXg/ah9ZX4F78+SA02SlUiOFhIxMpWix4C72/LlaRm8Abzi50kRhzPcrldV0Y
z1UWMqUTouuqq5GIap4OKKQwNLtZyBvuoNXS8D8SFfMbP+oHa9aryz4bdY0bKjDc
zdCofgJRvIErp+CGGmVBLjykw6Ske7WN9nG09miqS7HV5C/BJGBXSq/VQu+g5vQ7
RCRO+xMvkviEjsWp6tVpBCcEWyUYa18xOCCCeBfSywxf7OnfoQwuPXGccmXxNtoS
e8nKx7nQMUq4bGTgiZxxzYdmrJU3PI2dMmev7CXwjKYTS4dLAST2ZQBc2ZBOICli
Ydi+wI2qMYaOB6wI/ZbxyKY9B/RkOxtusyTLb3r2XBQyq0Wfxe0I0kk8B+Vu1Cv2
PAplW1HHTX3i7osZF16AvmB3iR9loZG0k6Ey+BDxCN0jekuAClsckjd167Y5+TM1
WMqZmW5pwDAIiGNo16BTSKvArQrg6TUyjQx+AKDebjR47I9x21RHRob+VeqFAEwK
U7oPwya5XdE9is2xtustoEEdMyygFp6SIifykAsRK9PZ7LtOh5FJPbdV0snjUTaR
G5KlBdFztBt/oN+n2l+9ZtafpUaREvvPpV5QJotA00i1essQaLXWffP4tX3BOE0B
rxeSotQWQeSu8SsE7cE5tn3uLAW9XJZUtagh8Rkn4QfzF+YnhBh/8oCCAZwkVhs2
V0g++dzHui7ny+K6aaD5fbOGs3XKbmsZDY3NN7sHsfyD0rHyPpsTbMWBKZZEFXhl
iQPDXvHUu1U4m9P6tWrskDpvGvNAQ7WipX8I34oxTp3H7A0QW47OdeN2DDjWP9lF
9AYEsv1SpTh/dUtYYtlMkyL4yPaUW5CSm6tXJLd18WFT8mBbaCw8Iv4wRgJY4g7A
C60ripe4LeY3mS2zUZKx0mvTgacxBGrAOYIXaVns8RJqawx8YbOPr5nccEbzurEy
rJYjzJmTDR779Pm5RwD2FxxH08kORccmykdvpsWmC3IozYE3hEvAVuMUg8pgonGW
Rp9S+Qx8BRdsew6Ab9Le3U9DYZ1uxvwrHsRHhwN8vLVp+eG/vggBcDlNblVjI3rh
b9ZodJ0j3hgV+0DFhII5Hy5lqtxjkwOzwz9zDeQRzcMMudfD8Dn+eC+DKqRXJ0tl
bAcwR49IqXu3NMMqAU0dcn6ZQxPiZJ+AOJLpb33kY1ksrCk2ny7nr22CMBAi5JEg
IGCV5wUvSJnZoWjPNChQjmW1kEPrz2BV2ESsW7CNCmvuCedQJZtxTCrNoXa8xGKl
9AOaCFJ0STcuE7slnMznRMQRlkUsTAif4ooHUTkV5bh0DejjnL6Ls+2aooYtPb6P
lXxY6BjK4hoEz4Ut1CLs8az3GKp3eF8omf/Q1NDgD/uo8di5N3mAuW9/WeD+7QTF
ekhrOo1jC3pZE75Gl39CbDkDTexyy4lWgWogBTlF/HrvfE3l26Qe4THdESZQ9oU9
s6e8RSc+VGr49vbES2LwdYjBbzDi0aLwuhvSflTiMouqJ9VF52g4aIHbbZdTsXcI
izUlVhM8kBm63dXRa7kFNl35VWDbvqeBhFZEvPmpqrK8N6roMRHZlYlDyENW2U/4
69xopT1Ludm9uelTr4i+FmLrMzFqQoD7RxiM58tgBlUovJpl5HFWMDYYQHppLVbE
+OuTlSynARY1qg08hV3QyOiaRzzv488viPmL1IOrnM7OlRUaVpN2t5Imn+fGE9z6
U/1b/gyeiS1CCAr2Jfhfyeg6TfrCGjr2nWQ7X8APCSkBRRQ3/EY3GB30Gtq2+mP2
tj6qcQ9L1ZasF3UK2f5VSMDGw6ZyPt9UMSLoVhkk+obxqm/MtNWpP3/Qn9gWdZWi
UKFbDzOAzSPMUZ+hLubr14FCAzLkRrcjJxrO9mYW4+Rk31C2SiPdjP1g+Zn3niOv
1j5Kn8J5Dza8bGwSaJKdeTLq2MK35wt9yzbawg+ep56QZFefk7HWniHV0iJmNpPy
h9uvtZhY646lE89Vc6b6NhsmwMBNwhYwzRxN/msOwHW4Yp6mX94/VLjn4nMib3zi
DahZgPuouU5PZeroimivgfFPNErg87WxjpzJS5IjMFtChpzlHzq7nSWyV31yJIW2
E6oyNYMThlCA9hO012d8koV8npgkDR4Ix6QULgWavwZHo0FMWYZPgptNIhsrglF/
y3jBGQ0EUvIgZENwybNDuz+FC5DxCxZlrelml+qzJXWNir2/9cwTx4/6i/9/IKmV
ShKzUs/xwsAxNwpRQbNvju88ahWzXo2ju5y1/gSTPI4a8uvPHtUZnTAqHpy3zr28
t4fsFrrUuyk4cJAHM96DFIIvLtKb/MbBxyKjdActRloDaTS98pl6MLLRmmNAvyhP
/Z3gUNRI0IfS1rndo6NcpbUWo21zTj3AYggqQVpjNkzCcDbHhmZGaidM6ZoaZae5
xzPC36u0bYxU/kTxZUoDgDvzyX0rvHpzZ5KSLGOQ4fheup/673eyZdYysLZW8YD9
Qhg+ArrHoi1mEQfkCn7HjhPzXBpmDszfu2JsEOTHGwnP8ohGcMBz0N120lNnU6cO
qF2gwPAq0iJEIABDTNvBB8ZVyUkYLWop9TZ4gvgv6ByuCYMb+K9LdKLGPfxN9L0D
PevX2dHVPF5ijrll18WPcLAJokLivsLqS3ew7ISqrNZvtrcqUP0fXTw4bAbOHOIL
6ALpbvGHgt+0BkQIdm8a/+1LXUaK4+nnPIs1SaLwsmO8UTaWSvndR7mqmL5X0iBl
j/Ls7M4komCwd3Q9k2d1zUvLkIvIBxFadUkJA/DsjdSHTmP0An8b1O/vEXp+A04a
m4+4ObiKgDQ45FHQN8NGZjpaSHfesuxg+1synqXwnoJU1PDrw/CbBLAIG577Tspn
UhkqQf61eFNTvBtAb8KCmRxsexHBAUi7JR5tBTmln3JAg2fWbr4gVSCr6/lRo9Bp
CCMVgYF+TVRguyiOOpFzh27gN/ecWq4u2VyaGjLL4nMHONKUE0XI/Q8DSRXhkwK3
X4N2ywOkE3RJyioC0eEprAP2clxa/cOya/Eru64joZ0EKoH5OAflz466XAKeu75Q
Vkk8qvRvtASqZ0ux+HXceUS0q3ZXEDGJf80Kj+98o+H5bPwH92W01bUKTMigldrI
ury+cYzx37wiQBVn/RgXL4vIdoOiW1yTYm/GnpND3QlerNYwrREsQIb07oK1h9XE
/Mjf1Xi75tyJE+GKh9YhosNqkQIe8em3zau2IR9VdjP2Liac3Av7s7/e9nD9Gc8g
tFBiK2JxzujViaGsKX/OfitJtQ6mHgqdlR9NV0FCaU18N6chJYMu+0mIFqkrpHAZ
ChiQwJ3L2edmlwqnhuppdmVXq9e39nX1N9GN6fH06sc/6l7DdModmQg1WMijxLLV
2Kd7h7Fr/P+YYK2ZFEKHcbMkPevvwH6BzW2J5TcHwI14jdw7QmBWlBfs+wAtZmg9
cRuLw9Eqc+Aw1+W6z+CbhGysKiSSHEyUbsUTeeEyf2x5B85bhjmJUid5WYsS3x22
m+gaq+f/vpLZ6EgU6+0Qn3amM9yi9A9GoSW08/ANflEdBM4jCw+IT0B9lEv7vLPx
EiPQJY98E35Zqmd23jk52fhuG3+hcA3TIR0lcMWkWsmAJRKpaXlhYlxPcurAs00U
yYcMb2rMMBzhCvNopm7Ks/Zlp4dHAj9r2PEhceSi295QE3Olo6wQQWxnY7J7FlpA
0fXu3m6pQ6I0K/GYSb9fawGL1air4Q4liqtVnaiY/2QFqsiNtFjXuFQs0758gTzt
n0mJ/VYy7Wa7RGc0guJAYZTBwufFrA5r6MOUhPbi0inTFpumnYYxD+Crsi0i2Orr
K6o1RrfEDELORZOTm47ySo3FhidNb9arDswPhcGYobiSIGvUtExsyXk46eJo9Gtp
cnkvej5kNx6xT4+Ty//nc5rzHoswtQ9RIJKM9JazNnyzuzrZtcdX779cnxc9iVIN
wp/87maIzODACpU0QMRswbgRQCqyxZ/tbLd3vqcn0pl8087QiGQR5KmG4k/mrLRM
ntpJ7L2UekRSRtQE+AxHudKBOIfMjbiBYTAO5AANIcNs+YJnMT+91nDeZ0LwxSSj
LYa7kwML7f8EmnMUSqb8elfn6vx1lbSuUjdXlhGRX6rgevOLBTKWH10jIX2Jb+4R
KD8HHqN9s8g+aNWU3eBg5/4ZRqVUnWQSKXFtCMQCTtjG4FFXmE5asESgGvBfQo0d
MFhSVWR4GlLwHXawSHxbz6A9/DB9vYZ2HWybpa+MxhBt/YSY0IbWmCYQuEizokch
Ig6eAD7dEocE2XmS3ogkvWGFn9YLZ0RberGuFtiJvOOeVLdXAyH3MpgeqhrUg5Zi
v5D6Q05pe1J7c3FBTZOkheMO3CvXdudR0iSUQ+WEUe57loY97OJXp7IHAFGL6RRb
UpmLK7Mmss9kU45r+R0nxbq1lmy6qjsIH1IINkrhHEbGKxhF5aKDsvfkzHghvKAj
EZfzr/C7OnJUvFwy8Pd/4kvGW9XIofhZE8pUzvnsfujEB9IxS+3TIwluogy3ftlK
g8IKcSGOvCVO4cZVzMNoE1ZjPZR4Q+laAAtCiz6+KlIG7G+auaY94qJrsQxc7FOR
IFECb4KCkPV8eM4iQvqWlNvEsId/dt1yZXrrTJZgsGYpZ2JMOBDgID2UqKjeEhs+
fQELgb1iL5XliOABL3S+IeHdCVDJMvfRw5FpEhLXNPjXqq+c92tHEQsCqNX08rl1
cOM/BGFT55NH8MCvgOGr2M4QDJh9WjQBdnWIrxuwgkW9KJwSVsi60E4Eyz8JSp5y
mTZU7zAY9/JfxYSJkhtiLoe6PeZOp+RMj+ZiRKMuatjLUDUMmeyqLQnmuSlSQS/d
D4CyEGxicY5TBj0H2bAQyBqeua58Li3jLqMrphWtghiMw97ZsM4FvUStNMY1tLN2
o7pVZX83qfymhLtuZfapany6Jsau7PkDPBGOzrq3V9xeMKPKs5AAHuo3S9orMYJ/
LOgxJlWLWkYn3Tx/V5hkUrz+Ne0YVF3GuwjIiMedFXmn9BwstwU2NlHcyK8wzPGY
WBrZyVltc3+qv7n6b/bGnXCrm2O87anuk0Ejwnu/+Ft5FC6L95xydw+t5YmOBbry
UaG1GNDlG8Tv7F9Eu0orQM7F+B2Sp17i02dKPNEgh9Hpy87IWCE+9C+4RsnpDBKl
b5sTjER9JeEZm0/F3rxRkaW126gvVa7wq4r+d9ST+bqExJRGjiJwxvGKV0IRc3uT
6ertMoMQjycVzAOshNTJOLZXKe5IC8CTFQl9fnKF57/8TlrPA4YsCyWQ/Qbg2Cba
K0/EzLqKVYGCuH+sq/xCzBSXJteVWOn8TIsh6nXXeb1JG190HiUwfVX2H/P2bbLr
/cOoncUg2lEmrrDEAniP/tJOYSWtnH4vj2ChQnlDttVJUhwzenw2FqGQ0H/dFreg
Izscbm9UGmvBFWUQH18DEK8nTGBYYmaj5urY5tDySrdi2NFQQmhxWVfXELjXSxl6
FyHC2vHb1On38WrJO/00X9CtWY4GnI1mdfZwWo1+WvkM/vasqUDcTnaxXVQZpfqF
PUKj3NA58W1FqRO6E58i5dgJtgGOq92V4eVlVU1y9RPTMc1CDQXKgE9X9ugUSSVg
3T7MVAbmSGNuqBpUz5c/zKV26IDQPduI5L+POTHWAXIXxuTRLgthz5qhjRq7CGdQ
SJ2/wmFA5PlLmdd/LI55OFqp2NLEauADLjjMPw80s1ze3AORONox4nR+X4TcNA0W
KUqxGWFhsITtxRr5AEa5tD1w4uYGyOygH4iW4j84bh1tvDanrorWeApaSFykCTWY
s3DHT8xjIrXsA6HhRXEuvHImWmU4MZd9PkrnVG32d4JCBYysWQmc2iZsi6ScNL/p
cSTZ6Nsa7oyoMreJUgnRIyyR0KqYe/4TEtO8+YT/xoER/ibgODtQNaL5NTx+je0r
aAp5X2yLsuZvmYpxWQ4y+x4JljRcXaMJJ0b4k+C7FFFE7mp+ClsGoZI/DUNIB0x/
xFKsBP6jQ76t3pl8U0MyewVUrT81zZnV4RXhQrZKeisZr3jsMI5+1219Gzi0NhpL
INQQiLMZudQgIG/JZpkoj3C4cPiJNiS3/BioFEv89PC5s+BBxINGI80PMoGDfiN1
bZilXkHXQIIpKZqR+xMLO7oM8AggqUsFi8pX9KyyGfr3T2ZVel/DeKdRX4T/FVsD
li06EKUSPLccra9AIL/7csur6eQ5dGOwgjIgcUWrtA0fjTOXveFz74f4C44fLtTB
34Jr1yNULzKtw73TXK8pFadcpy66EPlZPbUPqmdBmqR+Rhn20JkQPiHSMKCvAIS1
GvlGcOuSRVDYFuodzqhWq3bcJuQKaIpVKlyJdkyeneT0uOWP/XSAF8LGOY4tHiJv
uRM0wkRN58TnrdNfBUuNnIsvmFQYFXrtJoiPea2Fv4oX3rSu9s/6ft6E/ylpRdz3
Z85cdyJwqqaCUiTH59WiMGO5Q0ylKsOWnF7FJwKIbXt9avPyysu6SAhUy+sG+KRq
U2sxZbEazhHcu3FychQoTw+nzh2FJeZINVqEswX2dF7fbCoMVa8i6LZnqVQNKYXB
/Zk1meEyOcJTM6lL/M0vqPsAQyWR6xg6Id5AEXo/Wf2At7IYndvQUeSZPfV9N5dJ
q4AYjEY2nST7dM5Zeser96Z1v2+SJ3ZPl8lk9D+FC21c0lj7kbQbZvUysQZmrZp7
Qjeh2E5TpacOvrI8ck9FgN2/74q7aGmfCdCAh/gf07AD0ftOTZlv7cNIRqa39GAv
OmPltMGvKJYKei5mes7s4W7DzEIICTPSXpjauV56yJOE8fPbJ2stLX5mc6W4yDe3
JSvD9I8AyoyRRjLQnqVkYoqfx9LIny1yC/ncsC6hjvZm7zSEWcwQC6YVuHKsk9qY
LqRq6VPCDLLDCxcL8We/YHjVMuSLLPCGXKEgAABbLNePF+Rq+pVH/nwZT0jkdoee
M+aj9P2Gcakvct+D2sh5cTdIu5Rjzo1yhRIsSq/rDQXn5LQjNKHyDDftRLzF88U+
2yS1oD3n09M1NC/r1gkb3GjXkjXmnIx0Ft2/ELuN2lq4cvOsqdhhIy5smU9yVBbi
2hu0SpYPsZJV0r/t2DoG0LeChH+c9LIxd68Ien6+R9NNni6mjkgmFjp2IlV+iOYq
8pDpsFxzPU+TjNVG32q49RHuh9iqHJgYBPX5u6AZUofJec/AZRwSDBhqeRSG2Zzg
9Mc6acdRbMc3Q/wdn8AW9gHwV/z/UVbLhT7yubo7DtlTENEGx8VW4vE04bxrY+Id
vMu4/DODUlpuxV/CZO2LJrceuGPBGGXzVemZ5SJiQ7tbk3n776dsBWKAmLDslrcZ
3xRupzL6kCy9cklGpwiCPrMCKUwsCO1/V9SmjLNKunVNG9pt5XBQFcZ1whhneHV1
sUNbw61kQ8mWLSlhq08KuGawA1FJzYn/TzbIkYg9OzQEboBP+axTg9clZ1f0pMo9
Dcnmp1Gaciu+3jK5m5CnF2wSWyt4EyJlYswaDcG6+jG8XLjNB8xSUGmjCA5jkJi9
4oZhC7T5tOyfhrZ+taz5aMc2v4XlWoIgEHXhBNZRA3DS+HBikQLOOaZwoM/OGy6k
I/2qC8V28ZLQyqH556YVJDYi5zBJSVAmg3w6p0X2Lq9tZ4i9MisX/Wm8/te2Zi5U
5CBuLFDJbq7fyttNYF0jGy64iNLNvA342GqzkAxITCkz2rPDqvZulqGCHa58wPrI
oao/qAtGCci7FSQFK6ghgmUesA3lK+rGOapF5GqhtQ7wOQoExfK3yxQ0aw+5Ikot
nG9B0Ja5YST95uSZAJwxVCogUtAzl9M6GK9AmMCapYuCJCil/9VTVxeAdnb9Kx88
jiOb99hzo1ALSgy50fnBRtl4b7B9LbDyG0v8HJzxS5NOOAIBj05+lSaNBv+0mZnm
J+pTz58klAQF+thLZN73xsFwJNws6UxaoMWSXfNAYn8nsacCAA3GriRY+7773rMo
s2joEbQeHV1Du+m1Ro4qwTzGLMC4KBf85Om97/oUVSqfShIbUP5e6qo9zpF4vUxc
MVWde55ToSqppFUJLWNr9oVb0hylZubemyWtIh4o7pYZCHjR0KQZTpKonyTARyIe
5Lg/h9fYYQTCKVObG84A629daMbS4TUfs2hi3M/Q7Vzqo7bci0bcubW7gmuVCHph
eUPF6x+vIOrVcFduSXo30GLvz0HjSsS3CPHXGA9zAlq2lCgHo6kNCG+jHNKgGLF2
QFrQNfF1sVQkwjtltD1O9poq91QQLR91FxA7Ud+J24lJKcAiX1Ij/ndy0UfnqA9i
deX5+XegYfu9kj+msf8PFaski42V5xtnFI4GNpMp3+ZS2UU1lekWeSZJUQ/XwhZq
mA0ll9kpnpahpHSbdJFw0koDqag/HBeKlgISuwwtWwByKSusXutZ+TrcsQmMVYqt
Brz+9tEZvnZdnM5e2SYZNbRVpeqBZQ1f41lgAUZOm35aDPECwgOdCeUWiAaioLTT
m9czWUcuyM8185KiIevFWMYvrsS3sYgFsD4eSvGmPPJbn0K7/9Q9hyQPjTaGVONo
xcE4eX6kxS1v1whmdnPRS39Mb3FHMDLTCVPbyL+DOvT/QMcS2lLedt48AcunaTYf
oKZuyY5q6kqh1pvIGddzKQuFBT91FuOT8xr1/oNW0SEwKbuWnKuQXtmmCN3zqd6+
sYpKVPc4nnGElxJd7h5I3w7AQYS+cUm2V+5fAeJZkE1hfHYWee8l1Vnp3Ckoi7uw
A+47+fmlys4yZ9IMjCe6nLZP02rmzaezlXNunjYYw46vMYdkxmhJKbG8f27NXiCC
O5RjKr3PnC/+6I07E8VOG+zk7BSzUvb3Zmb0ePukVFUm3Sj72CS5d6E+T/Hm3Xbu
SNK2GSkzAycOTAaqHz/ThbfAT/vOoEiThTz36W0ki8jDyvm5eQKiFIJL07GRjUu0
LR6iS1decKM4YXYK7ftBC3OvlfVRleJa64GCUoCva5HgpCSnHZD74b6WsbIAlzeQ
S1thE4QrDoXHq+PJVrN7w6MIMmDRrUJ2pMu7QLWr0S6zSpiCxJoWpz49V968yL9z
f+PkIFpa5y+9Jhfw4BCpMj49wroctmZW0DSsZ9OpfIwZsQRFjiAis1vCZmfrew/N
ZIRUpnLnMhaAsx8CPueAepf0VEd0TqBOyAubauzIykuAw+tQ23BDj4DCmG/slCjf
+qTI9wTl2lr2/VLJMp/m6kVCsBkMbhLCe5ZD85ZHPhxmcSLV4rIysI8Qg+LOngen
nPkg6OO1jzaIThxBNxNSbH2yHrkfFtdwk2sMjQCKDD+PcS2E2WjLn60ulPzxq9zi
nMYQsrhW9Ep5vU0pCoojkaGaBTgWaqLDmSkSWr9H+DNA5z4DTwmBL2ScxGlVTPRC
f2esS1JcrLwMUQqcE4f55yjFeS57fmlvhIAKDnWBLVV4AR+J6vSwDI+Q28Mj5VrO
+5HQqmPrxKI6xx9FMEhtKsUi4CIQbrXp3QoZMFG+XSBuigRVpLcj6mXPvUYuySaA
3GlRI3m87h+q4JN64W4f9w/4NAUb2UGatA74t3KwHPl2QUhF2po/MDKL2+8QCNqL
rI3/haoXSChlIqAwm3Of56ucehNRHCAqUCOaeiIqk+kMIRe4+2BoIcRS6R0dJbb3
r6aNjvEtEhJgSBOcDZ2ilTi7ipzyd3Hl8tgQq1Y+BlhRPUX98zCfn34zKKZwWP7M
qn1IVsmtIPMSfr8JX6XANBwEH371KvlZ/gAtb3CzY5c8dk4M9VgZ+YPoo6VBevI8
QXy/tgAiXE7lT8C5KgjZIjf0DhF+EHEPkyvhgnspWQCzTmwQjiZoYo8MSC3f2PfR
vIkoucgQQ5mwGj2xw5R2nJg62ILztzDPd4kuRw+u/c4LTJdk5MagPUIQgs7RSuyX
jM+n7UIPLcIC2Zk6/eRNLIfTa3IfK/AHhjTP5AWR9CKpnF5gJZztUMw74O/zDNuO
c8NZqtZk9h335hW9VVu1+QeTiaxSx8cwAOH6gRISDixSEIKSKWpn1/rZdi9y8TjM
sS4HpLT2CvXd8eoG2FGK1x4YiUGdqzX8dD54AfuRIqlsi7XJ7p8F1jJZTjFOn3jI
p4GibqIeUN1VUgMBKZRoihVYk3SLOX/VqZoRzDqDSS5yd97CFr/XGmGrXbt4EZLo
yC5sPhbTzBrQr9SkD1R6zqCXeqYwl4NB7zVC39hdz7KJDrNebD4k8xiBWUDuINfv
gknqpOfz0HU6Y1lCEZJ7IsmzFBg5N3YmSTu1Yxhq6c/PGxsOOORSLScWCEnJc2Xw
Y2deScoqod/w6dTFJ0wWzjrDQ62AoT94+LFs202YeAVb3mv1lXtwYQE3vXTCXIQt
o0naIi7Kd4/9/QOTv6oMTParjTp3cgGL7s96bMtReoLIUYmDUEaFKOWjItbAdJHW
z6ZHzQdIKn5EzIPC1sB0QsV0zuCQs2BNBCm6Ws79Aa//D/sBXR/nmt32r1uDh1z0
b8QAFnoQShEmxnpaHFJf+lrFEdcIieZR/gG76Hp3wmWavMEKWy6fhRNKr9DhVqMe
1bgD1ISTC28d5F/ARP0bEbU98bsRg9CVFtzTEPjmlVRCoh6xKulz2UgHilQL9oEj
ALVi5lIz9tG748JkjggoAtRcWCh5sSP9PXU29ZMtyoRsfKR7WKPspI//JyG/IwnB
Gu8paHufwEJZSNAOxm69ikYcRtZeJ6D8UqK8olUojA8Bm9FozfwRLiBAaPLXC7BW
n176Ka3Us6IxYQovp0Co+cnaUvbQjsELsHDqllIjtvJywLdsIYQvlHD7TzJtKLxM
YRwutaO/GjoGkdcoI0/CjFncHrfwlaWuIpN/JDv//0cuqlDswLRRhylilO5PqN8K
ki52o8xv/vwOmirtiaad2EToko51TuGUp0qXcJ9W4h1aAHO3vrKg1YxmNNoozump
vSrb1bSRN8Yb0Qa39rEREEOQwXb0wYOqMvhovIuv7ParVJoSHEP8vLUbX4nGlM10
twcfykYO1+y44lewfECtDI3CZLl5OdQLmpLiNfd9M9nV7M1ctO0YDfnf7NqxVLx0
AORlZFhsr5WUbtPO7yaoDZdQNPADS7HnjLfor4inSIPeXjGWY22fzMEJBWYw/Ybm
pWvfBir/Bfkj357S7htz5PS/u9svGGVmWNWL8iW4PBbZdGbF7fw14EZEgEv6kxnc
Bia4MT/8z96SKx040kRMODpW/owyJV+rbf4lQgbGYbZIzL+f6b/4AzoL7UFZlfA0
8iOR6YsgVrhssBXu9cwE+qGHMNEwI3KqoWS5FOQh+rOIZE9SqjTaWiCQn5lqMRU/
IbMwH0fnW1eVmsHYcF0sB6nhhhADDJRdA2byq7P2E+jQHvcUVMdNkGeXIQ/sLMat
4QOzn340oKIWEXrtXNhKurgqmi2zLZoTp8WClTz+Oe6EbGy+qZ687gsvTS5F9XTp
fKAjxNE4ouYAMj+Ea8LvNLDPd2xCM9gy65RYC9NsF8YtqT81OR4j4GpwyY1mGEcV
aWA0diOI3yC2RjwzAVxuR6QdFdWxMqpoeQjmsoavJhiCTs5MMDFIrsdcjT4bx0So
mpwaqRUCKeSi4vlwhKVWXngrdkFUosis2dOsxkl48epuesgP2isV43ggy9ZjNrwZ
ls3bNrzi4n3pyZdyBhLDgN+s7c13WzPViPhsG5xXIyLvp9Gzl9nvwxyMVdfwOnbW
E1FmqhtWQNV4D+R+ZAT4FSIMTruV3wlEP7yz5L/rsGn9n2OKL90sazwyZkLJM99b
wwX30KW1NWJnezb/LDq1s7ujH6Kp260quLAJTY2zGQTyxS71T6uO2LYrzoaFpS+o
Vk+nQYx0FR5ds1jeZb+r7UBPNDmsjVtjAi+7x55Dbs7ho5g48iVSNLzBPfIFTDpV
DWpj4oIevrMY4kYgtdV3impZpMkzOZCznvYvnJVXBpdItn21arGsQeHPjt3rKu/q
XKwnO5olzt4N2sj3MCjuJk50pk3FwD+ddcYlIZkcfmNUSJCh/8rb/i660F/rEj23
uZvpfozgiQd1OIlp15TNGFcHDZ+nYC+GycDgLc+h4LPfqX7bXd8s9Ed5JSltc172
xnOSiI12By+Bp4CDQwVyYWTj2IBQdpY/G4VRmQ8RvwsDXuQRyuJioN1eFTwYxTpl
gUdHhzvnUeXjihbT3C173Hj7DzOlcIhcgFhzFphacRr49IjBV+WcDKYMmOqVWU2l
LWhNS9YJSqhc5sYx3mMcX0bl8+KUULzZDZ2Q3mrBuxEo2+kPN+EvObnkVE1E7F6/
gFjrWK/oQUpcfuai5vGBpWeQRXYbrV780f+QENOZut3VSl0y1QYA2ENXpyF95zG1
j9NpNqlCYnSvylBLZzHnn49jpY9ppdaToRQY7qtjRW4ceWDm8LR8+mShR7RIrPFE
GCg7uRq6sIVnB3FldwrJEjMVC0Cgazo13ivOWjCft8SEJpNaiH/JIn42lCSXCD3/
43qriW5Lj7ASHlSzPfWHxGOCiFeOVq9+ho9nNrw1taG6SPIjxsKbqRiTTQJ431UU
Q0hNLqSDML/HfDlpz2aIhqL4sOU8hqlXsM3fbLGLFEK6xfHNYowfiPTHhlj5OzFf
s9j/VybEehlfzJWWPnNujKp17cYWwu4SVYljGBqarAmoFJTJFabiu9lWJrMZBKcq
6suiw3NpXsY6FOpuXx3e2brCCSi2JDA69S2MHNRJmzzr2cjx4VBxlwqzHoIh7rXL
QChBxhV5Sby9Uxj0ElREZ9b7bD67tPeSM6N4ucprCKZoxvISEx+2kyYEH2KdheiQ
P2Q2GGwbVCwKiA1+K+rPyKgNCluX0u0+d94Cn0hehkenywsK1XaD3VUK9k8R+WJL
UbXzWenGmDW0jFUCptqhr40hOxK2JDixNMDEYy/qYWnHAu+ORtSW+zn0sEiAlQUw
w5gC05kj39Biecrkc0LyhfiKbCmUTh1NKPB0RN4jvcpyXlPlDjTTDtR/u8RB+2zX
7HxfPsNGpSNXAP5/F7xohywTSNwvCIR4ufl9GUi1aoRyxn7v9z5WIugIkEkOB4TU
kMzn4YieADb7kwvQ3B7s4CvB+FeiX4SD7P3jd84RFYQ4isFdUBrek9mlhItB1RDM
4HCyAfBkE9CxBLsYzAb34RGE3xAjrbGdxuderB+sz/TwV2T+T2oosU/Hnov2/XEo
EIXfmTfW2ekaqEQtUEnP/PM901jnkUmePqHp7CmoPBwFg0Z3OQtJLoqQr29Xq6V/
7VQ4wZ8BUbgTVwD7o7LjvQihWHYoQtUqrXTBN5bYLOqPXfaDb97jn+Ap06uLUJ2n
+6vEPHEfSpGC0b8Y+aDOGgroJZagjEXfgNp1yarQxYwKCxgAr89fJgQteZK+THFB
fRQ65Cs8RzTHtrxGfpBjY+J51lYKncb6kTEBHLuDeaL2xPQyhgSeeE+eMijoq4cN
BsqAyqHNOc3z45Gc+vb2V4aaDfJ1TxARWlq96xXMqNV/Nqb2SJBufv5afP0UVyny
IAoJAWGGIGX4VSmibN78bLjjfcNVvNLlG7WHAq/YeU70DE7JIt4OiAMI8rM0setB
EWru5SkTvJvqgDGgsk9xGnrnyRhXkhdQDqTL1IAYoxPC/vkxkUsSK6ap9elRkoB5
4yYmKHOyamsNjwEmIiB5iNemCUyQWBx7DdQF89eE3wFb06q9Wu5S8fUvLZrlfocR
lfc/GoAL1hjaFlF1urrqdGQaP791p8GSSXzlWToI1bPaifFBL3TpFAIR21bJsS4i
MeU2Sh0WWjb7nu4PlryCCRhkm9IpzoHNN6l136OTRUK26HtBbxNUReD6AelX1XyP
KpVezI+dBLN2IxTBWwl0LjpR2P5ec/bEsXLWiyO7u3hLapCzAhfxzY3P0JHeLocX
DSHvnORe5439OX7PwzDnr6tJlJQT6pC5uXVGAdSYloauIhVJ2fD3W23ajLvmeI5V
oLIY57nKfmx0rYZW8CJWGMGGP08DczZ8q6ejYT2y+Jv6V1QK5G73Xf6KpUXe/qxV
2aJeHDeFeSKIj/gCZjOTScEQxtF0V5kfTb7fBTmB+Trx0hXru51fwhIlVUtxu1tL
AYdfzL7x5HFrzqh/Yh7Tvj9BmZp3+Q+4XVWiwQ4IbpNNqjY7jjMTUXSnNMJnLIwp
PdmNv+WHSgrYDsU2+cfJWCsZJKmuwjTwZLT4vfwyeHkUr/O0yQ60DCyBoa4wZvRp
WuefXgF+AfyTuVU8aYcUJBWEPU12pm7j3DnpdPfsnrsUsyyckpR7TDuF0Z6IZY64
gIbGMsNlfrwoYzlRZAERDfTm5b26v6O3BTZ2nsKhOQypBq95+JMbfgId07vmf6Ft
NBhK0L0oOA/9j1pvpPjvBAo3UEoQnXirWGNoQzQN7KciQEgMWZGTTs4dvxZFcAbl
s4zR+UoRmSQisy7BjbAaKtPUNBO8rnXcrvYdzYzXWFZ/0qIyojGznSdIRj7MULhk
DUuHsdGPKk6DCSVmxCHdvWIwc4JDXQqkMsxycE1HbxqhGVjTTwwXA/33Y/Oml7xL
pXqVQhhSsfTzTHA96RpLMZgFELu3bkCZFKajGrVWkf6AU74X7JTrbZrN/d3zC3SB
7cjdw8TCaoCKUYJkWcnxMsJSkw7K67wCvN2cl5atfo0jYJOa5NcFALoqIATLj2dS
/3d8sHUwNayivWHGIv2ASnLtPdS6zEepzlfTZGilb7blZaorfhFxHQl/gOT+rQlD
AhDOxrA51v3w9gG0S5gatpJC7l3Lal/rMsx6fdEHxHTzkMI/a0ljM+IcGNf10PtA
y5AxE2k29GkTSMPqMLe8b0HvQrTCA1ZSDcUsdeY0ke2ERgPXSbE5//oBdBg59pN7
wlITusnzAZ7m7i9/CAZRhx/SlU+4BYJ1ho0nFbii05Ndgn+qx8mJAz+pyzwmIIVZ
pB8j5SFb4A+IIKWa2XadOHrLB9Fu+vU2R0xt6Uce3/xR2sF+TxiiJCPVK8SsYmgj
7GhXIOLl3cP03dMDSHhNkSgUcMRboYOQu4W7OpyO81DMNG0K6GsFlkM2XZuADcAE
dwpjVZmloe7ep3MvcGEOr16+yaXz7pZlzEHAyzJVDciuQJGLLQxvSoJIBwPJl6DH
KO6IUO+kshsVDtAr2q7KAWKUG6XfBqSzyZI0gsgTuvXF1riMLUCcIDfhFEKxXB1U
Rc3x/Tz81R6Q+YQoTSowU7yC7/qni4zEdYiLp5+BbMnStMj5OuZPxMyDPdz5BFXi
s+e2wdIgZ68ngHi3pogRC3AcGqKoDRo0oS4EWIHC01z17mxjcn6qm8xyZX4pFq8n
wl0TdVUKQxgRInxsU4JZ0h0DFBxvzuOc5V315ABx2lAyac0wFLRuXbKnH4jz1wp9
sbb4uHC3ZBUgZqHXN4F1gyKPtQ7vuFc3DLK/NKDP7RLmIvXtJxNSDivPf4YcXoYB
UJuz8HD8FjZDevwPD4g3LHgYzOuhStX1RuRzDrlyiKs5Idxk2AfhvHQ1+C+omQMb
SVJ9opKJLr1xdzyO3i+qcDZkv5H35Q0UHGY0Ua3e/QR3M1kQ5NYsJfneJPo7LmQX
G05GngosEh4HNLihjs07pxgbPjTt70ePjErRhlDhwVlMZ1qoMQtkP61vOVFfgDIO
tPt9lpv4n9cg5qcoQQuamxRPHp1FLRFKaG5EcR/v75QTDN3SXWAz5NV/gfR5sBja
qcteEyWnRcHf9TpNwkKTOg/H1zEJyLoM5oZY8iZxwLw2WF3cNOLI5dWaJ7fr/i/D
tyfL242w5AYyf0whrvv2MTEiOnHz07aQ/PPmMwmilhCgC5zTB6y38MTPxAMkp1KM
/FSRufHMhI2FmZCvGQdDMNVObvXpv+9O34wmg3DoXt/wVSqfwDATUQ3nunlYF7gE
0A7QUAkTCZI43HrvpNQt4xVrQid4sSUDVMYiCL5d1JTwAnQ81bAe9GX19Sj1wKZz
7ZOSktH/PAxJA2k2FsePx0OYU9QICz/w0RjbkuVZXabNheeRUmemKCQPWNLNysBU
uegRKOqPRtxt+5rQ2RjeK3aXo3w+ZzcIciLfoqYhbMOzGMWhEHPPy143nvy6mN0k
MhykNMqLm3RoyWCvud9M9RkA71ZBNegdmqx/oVgtyIuRfWP4ZgH4YJoUh3PZAHKi
d0psO7w1my3zOnKsf/FS/XHXSInn3m1RKKMo9SnbMyv/cg3jreu6mi0EACiT9NNd
O6NIGvIbLYF5SgXlOUx84uHqswjYYUF7kGQKiKgPflS0zc0sGvvR3aIR83gcML+F
ETi1yUjii1JsSchlWXcBoSAtx5fJW08ele6mNWQiTwsSd60sJH/VyMHXgZC2ENbj
1gDociNgR3cDo8Gqmv0aBVbYhy7eBot9zusZ5XSgN57xbFxZswJ/GsJIMxx/w5DZ
VCZ2Vj/GJzYXXrR4FKnVeD1DhFB0p0oSuTmhVopFI+iA3u9GQc2kIrHR9+GqfOVs
oPOHTvazxU3RcIJ8B6spd4XYPgrh1PLd+BwVWIfXNZkb+x0CW1OmGVRryJrZNXRy
JO7PLyNkpaJ6OhOxjaeXEz6ZPc1FyL9QKz3SSVCaAtcho5Z04Ej2z7JbRHFVwE9R
I+x/PNHOhLhA+ZhpumMAkVuE9uhfHagAGihO0e6828XRnsFoU3Pw+wdxcm4pYV0S
ThkS+CE3RB/MYOEb9JF3ucb2GWkvJ8qwFtVQMvjHFWqkPh+0cJRawCrdFgiQhMr6
PHS1a5Vx/pjzcAiNfBYPGK0lkm0uuNibC81MnYMx2QVnF2Qgn+bpgPFULnq0whTa
/alQYnV0thjLsunz4jaMuQ1SnE6VYmnMvdqaHQO5orSRvwN5armmuw55/b8tgUf0
6tJSd7rXwtQEHjiFyJsDxV2/RpDtFt7ruOdNXf6n0keua/NeLtQipF6E3oNsIBMM
mzCTZe6vR5W2QLUUD4VK/D+v0iayTkQ1I46MLLf6H4rjuzaqLmp++3myGs/BhEIt
MITnVFRWVPAJZIOu4WIt4W46II9YoB/ri0GU1Fct8ePpw6Kl4/dn6GFxS3+QCsxw
Q2q9Jn8h+cy6x7lXAP4G/llYGrNAXbbibXNFqPxMtCxhbMsx9R9znJCaeWTTUgbw
c2VBHvMcu1xM5sVqiD+8GbzClzZITKoKFbTMPoCzvoJ9HSiMXmjFNWbk+aJAgA80
wMpBbkGPuc6EeXnP7Yo3CB6aZ9yVUddml/4UHB0DHKacYXjwemZjmDlkoRgATTIB
yXjlYpLnOBrAfhaRzniF7ESg0J1PiM5lXW2vguTnIHepJ4hT3k9hc+hbeY7y3dWz
4SdXyAvv6Zurp9yyrA9yfqdf0EtfX1MoJsdFH3fqbU/mY1+5iTnd32Xdcvv7all0
lX5i0A+YPsNQmq04xygFPT92l2a6QTyHSr1eV2C8gTYWWp/KdlvJx6Fgr0Qzr2+5
T7ubBZ7+vbXBPH5Mld7TEu0n2FKCm/c3k02zIvqQutblOsOl0MFYxF+MKPs3r/kb
NG20p6914Ap6X5rddp3rrHVk2OiuHgWHgWXhh6vTLq4JcP/3Z8pKe2YlDNMj6G7I
8gOlhn5Xq/3JwlzpJyvvPYcyDMSltvWw70PnxnxRnXOvvOBoVIccXgOZyq4R29ik
r5MeBVfSu6Zeh0o8sCGrcjK7hIuv08dZdsTHAV5aJSNI/nzG2udQbMg1H/ftz0se
xmvScbiCHMxMGwSU4TvmMWkvQoYuPD7m4LpJQDBWf+NGB+2t2Ls1GRLqEZ4w6RaT
yjeH4X8w6lwG3/11oSu1SdQnUZA+Zdij5rB3Gpa5PUApPhA24qXSw8+XJRwaio1p
MSWOIFYnAMssTB99dkpwzrBibkwAw1NdOTC5dkR5+DaVR5YcfcbSALko4XsAmmYd
tHnOAFBqWsChi9oeI61a1q/JS9c5Hbix++0bW7Dt8puApbzH/iXvOexSs1mIzokk
5rI5n5FVwc956FJ1cF7SNdYRH4KfTrEZAiM3S43in4dvxfycQ1qBMBaCnhz0aicc
YDr2RDfqG3x2/4VvjEUXAk062QoGm8hPAtgdbq1TIzfcC1Igu/00Ge/ghMTIZZET
KSAfX4f7ED0Rs67bOCsV8qz90p1mnTHF6fLQYAutWJlUjBf2zmh4+y8JUUg/Xo3T
JjRtrjCDf9+0CLCoVbqWkgg0G0xdO+R3l6Sq+oCt6Y72AyjdrEah4Pvf9tG75RZB
1nM4ng1fHnjkBTp6o2r/7NGqw9CjiNEDd4Ru/GbPnR06Zc2MQMMUZnJPIqQU+u9k
s4Vxpldeg9NVemd2P1byojmnKcIuQYmgho2eXGFuS48647ctvfgr+paCBdnVoPK6
pZcqvz1RxceVYXOhOLHIgd0sHaWlCF/sgA9uBbESerC27tgT9qiIzmprhOL6fSNe
yGC7GrqIbTUXReM3DOI+1WWz8/YTakhePQgaEtZs9w1FXovsOIDXPS+nFJAF8YqJ
gO33PVdMkEbJE60MuNGQE3oaUpg5rHf6KQwju6Ro1Z6KGXJcQdWNs+PcJx9MZcU6
sb31W2oQ7kepIShcfrUt0hB7mX3HPCe48Pl3ShoXPEu8xfZT/fGMxdHln68SxAtz
oqR5p26tyvHMIvoIAfSeqgmsJZmVTJC3iZNSeMth1CXH7CSYxxCszTPKq1vDlV8d
A8ndpmhH6UjMpGYKzbVKZXOlO4TBoklPa5/buVwoDGh1oMxS4S6t333IZTm1FsAM
aKCxpF0YlndQzz3bkrzZUhxDKOXcjKWnEMi8+TdDr1SdX3GSY3XtLqTTD+eKUauP
Vh8NbLKE/5K9k7z9kCBytj/ux4YYlcjDL13AslxRBIu1hEwIPegkCd+tz134WQt9
HDqg11i+IdYaTTx5kLKB0t0XYfiI0Uq9Y/DYO8Bi37JX8OXjalk3T01FIGd1udwJ
KGW+WvWJAK4Bv4rbdgnSomUrqWV2KPyNem4DF6CkMu0qSyfgC3DfxSA0LXHws3mZ
0M6JGUOawORJ4KO56gGxphD4HsD7A9XH5oZ8ZqOtmC5z8Z4iRrR+jeB6+zcWqj8b
Hn88D1OwP15UdhYVO4CHLJWdpc6QEn/oZP4xGV0nUL9UnKRs/HM1O2alV+M0mz+E
40iVr8/oCZK47qUMKHd56yLyKaZ/aGa6UhLrm3p6GcVW7IldeZ6iuylvLyMUzJZJ
p5co3YOBrSUePMeugJLKD5Uv/wAjeRf9kLzGa6McbWBDQrcDx18SboBNpeR6t2nJ
GkpgA4GtLIEmhc+m5XRhExEX9W7gOTYMXQVmZX37IsWSyCC/CQNok1BXgjZcr0JY
GMAAoX1wVqZ0SEt18U7Zh5lkkjYhB0EFcbmxdIWN5XZ0O2a0sFSYoaPGX0YUc80N
B+2IXdH0FdrHp2HWJOstoaJrEFtzKe0g9lZ+C+e8XTkE2K5loswSqxe/XbAh+hTA
Gt4OnVI2/ezPQP0IdR27aRbtLM7QrtYsSvgKC4uJflZMH+pGRNupKeuodMKMO66P
JWSDGwIqopXUcGGYaEBJlRCfg9240FMSHu81jKTP/KHNIYyOwAec7xP48DGhuWm8
TYX2N7uho0Z+Zz0oD0MviUDPZmb7kumBfF81GV99brH5zIT0ile+4+jcPjYkfOY1
EEfjs15bzrLS+manbQ7nXEnWCpbFRieDh5VLpG+M+L5KNkqDnQAWQ7u6mJCva8sv
VD9GAoyUaWWf9StHKd6sI16mAwWBG1O8kLHeEcUOmpWr0L1bTFnr32hDIhriHc9C
EXZzLiUZprGQhAtw78+rz8fUdLUSIjZSaiugYnbfid6yLux0pTRdhVmm5quA3pwQ
TYer/GuvE1g5Z48cnD/T128SqUimVGwpAHEeuhOKsGZeVJfdE9Q7svzvRwH/0F2S
8WvC3GuKwfo7BjPqP2g75lacW74Hyl/SEOTy4dFwwFEBVCwfbhWW8Nyt0QDxY65C
0ApOFUzAhrqwubtmJliOpkl5t8TQNpvWR4l+1eNpRav+xvuh6gmGLN7SbL/a5aZM
NK+BRPkb//RXVlEejpwGaoarARnZRCJ9s2RjxXxkiIyXYkoFkdIlz6fodi10psZf
dt/UCGsGXYQdM01ZwmrXxLrkXzI0O+pP5+hrVwOMrxoJPaOJiXseWYoo3SZX3cxr
eL1hroIQ8Q+Vx+tRfGUi6PepIns9LzCx/y6L1hWoSJCcyPr3bZXEiyEV8XlaJ6pv
btfqAopg6JJJZIA8DE1ZcPqduUcGp+0uq8QVmv6Y++odC2ClmTSPJin1S3j1eCjn
zF+gBazsRWPFbMspWlY9NDcaE6QjPYzELUGM2bb1aeFkJqGu/lPevgFu1iNDDrHh
yAm/qW1FlKK9SJcng/hTVEwhoGnZ81z/x00Dnyz8XphWLpgO4vzhAtrVuMRUxk4s
bKnyDtbsBwoNvT4GzVYMeI0ypXUkkumoBgQMe0HFFyo4F8JRvspDgtaStmeOicmu
zBmzP4gHmhiTR4EcH5e4ncqrXWiMabKymX6acIFa7y/yAbQPYc1VVK97wep4B+m1
BQ7y+j9o7LN+tY8Cg9w9ZC/5Uc6pSCbckOyUYgaMJ4hFrsVVPmpZl+jNqAVl/OXF
rq+N2s0l/5d5KcHMgpz+y/vzT7C2eK3ZKhBv+NAMn9qfOHj+NiYSEf8gJSARXhQ4
F1j9qRFlawlnrx79jlErVG8FnoY1BLzqWI2c+xu0QEsP7bujpBHn4QkQxPaXmIX5
+R3+ejFtbcsCpSPzX9oK8kajUPKDbG1GFcSqys/MrFR9ERa1c4N8rSWNXEUjz60y
YziWeHLBvuatEleXpBsCUuEsYZ7nAk9jDw3mp5M51TgUB9herlPAasoxcBq13xVA
fen58y07ZpDK1SRbtFPrNh0M12qvRl9OXTlfAQqhUOZ0TMU6O5HIQ1Oz/GVUwH6X
i63lQ/6CqQ9b/DtlAZpK6cui2THeA3EDLg2yxzbe9m07WahiuUc/Uq7Xypl0fZBk
iYXVMqBiB+uhIW2z3Txp1LxryshGCrQWaLSFelc1QqeKxvCSgmhyCdGaJUQyATCr
Cmc0nSDsYUSja9l9kylWMD3lqCrLn8BWW3H8BAGXdsYZ6oHd5877nY5yN9hSSkBf
EibSt5i4beDEZn+R/AUWy1/VIQvTEkVOb4BV0IbCiG/yQe1hRgTrzfix9z+Jl2ny
aGeKcNVUySulx8ZE8Oq0u165HRYYO6KOPj7p+k2SaX4VrAotMVU0wUwLsnWFfsYe
02e9ahtyiQwuFH6/cLAzhToS0JeHVTuXbvfbFlYGsTQnqxhSZuj3MeYV/VnR/qbg
ycyr/qw6W4zqH8zKNfhoP4j+7abH5fMGkS56kE1odeSKuOphyTZR8idepWobv7fg
7ia5m2vxCy33NsiCzzys/bsPIrx6yl1SsSTGDTNaQVDInA2iD8usy4Trx4lceYqE
K6DBDcxBYrUDueao54wwWqM0AlbiPceZAUDz8d/MR4oQ+GUKWUzad74LJ+8pB4zr
ZGf7qFf+Nee8esio79o3sam7J8i8CHgoO19jv6XGX3FflRdes/JkimiB1AjKunrR
xWczyLbFXHSyeJs+ANMY1wr8++FzPSkrVg/q0nOxj4xD4cqV/b6+kk0dzuuOp3hr
+cet5NNoyN6SO2jwvpg30exyN/YI3l6r1EGS7Bvq0cZMLPvJLb9QEI0huoGcIokS
DiwuHTNwrwze0YHnQ4EFTe4c4LfsM72FcY55SXPcsWn6/Ay7Wta4l2+s37ZGEw7A
7K7qPAVWphwe+OXyy6B8Uc5C069iFAEdZs6K0JpKoVirL+IheJGvqF425i0h28R+
5BN482qMXXkLTqounjZjXQkXTRWSRfh1g7RShGrQsNfyfWEOrKj2btjmcxv/l5o8
BdxDRJrx+NWFyQQ+MZXgLgvhMNdOvuZuz/k64v1KnMFDBdDzTXSAcy+VMJ3KjB31
VL4Zrr0E3jRTQ2dzQXqOvPZ4SH9lKYUYxKqkplaJQmxDOdUhGDtK+WRQmste4fDq
a8MzOfmR/tnH6uXLZ8SIoCMCYUaiQodQbmo8FVe4nlpYs1T1SqPv9c9rCxZKwga4
3bFPovc0VWdgLNvuIqQZQyE4pIOR4/YF//gktiPZX2zELhzKdc+RGVZIKFJQtabH
w/uXwJ7s2qu0hufT5EtR2b4WJZNiuuAd/S77iKOzSHbq1SCm62cEPM7V0UHfbYUq
LiXG5wAJnE9pnrtvtAAiufSvKx7BO/E7i+AHh9iYdFXPyiRKXFATY8uv3nxHQwr8
kAiek2NwItSNfaLyfA7z8780t1rVn8J7Z9le0ad8MDXbvi8ENLWYgyUJrA9z2n8j
HfZsvO0FgToobBcXRS5+0XJcNSjV8+38uzsz+EUxrbUWL52b3QY+zu/P4IhvEciJ
gdEMq34Ze1fHFnRlu56CAJTpJDosyq1q6RAGPWsbLPV/zzkwSz/cpSBbbxiI6iWU
Gt02jb/PLRQyTVqkn1gJUtJXbV+WbOiENrxvavOG+GkQ0shYuyWelSyjWusGz7kv
RBSSZOYMEoh+1e2oTI04iY5vcr0f8CiL2zcUBxP4LhnekxJJo8PlmoTaEeHOIsBk
1JNrxiIwHQtv7u2q2Qd2wzVHsPmmQ1vYpTkegKIaN/1aHzKs/0JqOVygWufUK2AE
REsKdx6Ov0vfOmNZDaQYgENrjUCN+Xr3TGIPBbJIRG1X8kuwNhShZZ2pqw+hjTsw
skvbYFkqqc+AMshdoWI7KVoVC4Zr04wm9jW5+Pt2rH01JoICcSytxPEUe/fgog8l
sC1SO+Gbzu6dkX1Xa6iGn0eRnYxtunotpP+84BafXD2TRBDAeO68TqnT8tFp/c7j
Gk5gnp4UD6rLkGGBqo74YKt5tq6NDY5lZJKkAfogduAPzlqRuWRHpgEaS2DtwBp+
nddAvP5uNPjzj/go0Cmj3zv27ioNBgovOVTTJkWTmXelsiHhPAYVZknbzl5osWxn
avCTocTOzdiwRMDPqHXQzs8KIe+abkmYcrJcXM8yxKfmDvh9JQV4wqPvl0OK7lEe
eYVjxzgOhpfgVeTp7FPzqIUAs+xvYiXoLVfwM7xJu0+/vPSvu0TDxJpxiYe/mEGg
25NUIteo4w9E3EPLWapQk6/1ITJAtV5iRODua2D7kneAiTrL4GyXgaKpGzNtzBl/
urLkM42RdnSxVt8u9MulxZIVNxNl9JryXwm3wZzU6pi0oyLxGpO8oHofTqEmUoxS
AI6xUqP2UKSP294LaT7Z29xOFmWw1MZ2+KokxoQcDJtKjiL5qXZ/IwKmu/r988Wa
aC20XyAa75RL0UWSuYvxvaunFQ4dtk8joGyz+OdCxedsaaAw8veIrCFjAceMCt1m
AvU7CXRlKidTxpX+hyGFGgN5BboYl4MtDHmt093ejzCHtXStsE5WWwKyzu3hTKAu
ds67A5+bki9jP0L9sZSVXdbjOXgMf2R6Zn9NiNct7MHf3qLkXAvEAfLI+9k954UR
sWBSUg27VF7CWzGkoX9be7Vfb3h6eyFsNSwv3yORHGnZI09prM4ItNSuZKtOUvjZ
VfNspsXvPeD9USmqGZpZqjcENRuofw2EjeHmoSBSDnaGzggNgY1iK/4+fZOecpZX
HQmBoxt20rqxjBoIYdRODGRxf3ZaqRhHPN3TFzcAYwZnSAI8QU04XxlnzjmXnqtF
/qwMVDxaQrIFxnWGdtnf6/vroic5PEXEsja51uOFdD0owQIKheniwnuQF6V73f5h
1K+domJzj0Jh1JhEBcRE6eyNE/IjC+5pbJ2BDS/6S3sXvIzl8CeaIHEZMmaMhRhl
fWfQGFIrJxpacSc6U62fMJIhn46zCkjCZGANu8+GMv5o5YXJlsJ0GVGzwsfimGA8
wvPGbQZp8yN3dszCL/ZDc3uL/d9wc4Pmh7lSFtYK4evwzORR9NGTBmb1GNBrXK+g
8MWE+c2f3QpNVrGmteiytxI8QQlMHRPW5Gt9kQimti0fQz9FgqqTYGELHwQgSJSd
Wp/SiciMDB4s69kEmlLmQqxvAyzPw7C4M8tsg6R1nJFOMZKI2MQovakDxt3N4uj3
EcAELvgSLmOnM+zd6tt7Damv8ItqXS/Ncx9Q4Nc0Ay4pUTwctnReZyB1BGkCWcMT
nDN4H3i5t41bjaE8hRH7RGaCw15GiCr6hnamtlnsV0tF2C9j/8wRGwhknZ8wm1uJ
jhUlzVHnSY0rU8xjqe4+K/5lrzPd6A+uJsej6t01uqJqGRSu9cKNMf6eL841p3P/
Oew5UbD6GUy2y8nEOPlycvtFSsVFyTlai1BpnyKfpvV0BdE0anXVxnrH2GgYMMkR
gJ+sEI7IY1xXrcjFVNmJTcvqUd6Gx2Y26D8rJo7rWQUcQn3TQaStPHi3jFuqgXzU
2+o15GvHFekeMTfR82O+hax3sYxypGH2yiQLp11z0sBIeN5+iesYNqD+BOytywwe
rlGYJ2H3wRgMFUqYn7Ltxk+HFXUa5dMOmmDWFGfDsOrTI5jf2yWFAh/GOgUJSCfS
/cSeTunepPo+IGPYCsWifqKPAQKpjBh0PY+i54xwCHhpUvE6qX0p2FNb6o7qKMUG
G2pkWefMMLbsLee/6ztzy6aP+xtITifFaJ8KZxMAyqyjnN0YFpS9DhgTr5s8NnpO
zjcMR/xt4gD0/eUxm8VKdciezGJjTvFjdy9Uo+w727BSXfOLzL/uIKokoiMxmFIu
j1rQ3qWW2OeQU4teUwmqEL6SWv+dEY/V3LpmlQkeQi93CEbmbAkL7gsvN3wnCkBX
AAE4zhOw3BKZkIYdytgQSANvWeE5F83Vk6S6jBhMkJB7Q4GCoWpy18znupJfz7Q/
MiEDyHf7hx9bxWP+u1Q+uObgJ26Hj2+OhGF66Kspx5tLjsEN8qyg+0S544r1lQ2H
WN+hU0ukYzK2NrC0kkM8W5N/cX0uEqjTaTtT5A/DDDhoHDKDgrQetnxNKuUzgP/i
wyD4Fv9qKlXmr3zz30PV6dv6YDNjTHThlWzPJImVOKQbTDHKajxBb7Yv/6z9iHQd
GGohgweeybUL/e/6ELRzANKuRKpOUmWdaUYvZwmK/gmJCSvIAX3fLp9IZy92G7s5
RglRmdOEirhsMj4egSQ/3nCPCMbcnSHaVZL0eMhP2PSuxdDE/ymyCI8ttVd0wxnE
Y707rYnNSkFKDtcLp7zikD/XUH7FDp/Fbw6BCklD03zUYke+aIv655MsN2oCvyvS
BluoMgNdfF98//DTeXXh8DoUbGo6V6nzMg+0QqfPoeUI2zEMRFR+OqNfugFN+luG
oUvUrhrHgYYagGK/C4/kM+HleIkYMP0/Kf8uKhrINutAAyMT/gYOfw/I8Cly4VWr
KCMD23CY2Q2TJXj1kNWty1vffTdil2Q64G0yvAFe+2Rmzjucr+mnrBIIAOfnZDPp
wteWNsW5rfDYo5462NIuihtl0vMJx1bKJGm8AQP3sqWii/cRhfvRx75SzXj1Madg
+BEx+BwupFRoRNe0ASme9Zd79zFzSqWV3FCdbjJ5HzSNCwwe0iiitYwGc9Q1FbYF
wvocDd7/0ppZToRk5mGYYP87x0bAQlxyfBmW07As/gLNXbk7hJJgqm2MdSST9lKv
N+vauEDizKRPXFD+v56iRo4Xy41Uum7VNOkyMBYuLdIdHCbPUy4ma+9ymatk5YfX
bcv6AbtsYnXcloEvk8lTtCEQgP6Pdg6OAxOamPwvze3eDAPU7zT9BSZ1+ZwIDAfE
nZ1SF5C1cFiMBkvPVp/rRotTmG3hVTrstbsZkBABqdeGQrIzwu5s9dQIWOKZl89s
lfOZCZmDjXOXe/HzsS2j869V6SsAdUzLcG4U9IPDfYXaoQqxUwBBYPCtLIuka2W0
AHSIVkg4XAuAoHQVWMexOcnS6wKkPye6czus0fabVWzcxlbgWstdAxW2BrPgJ7Qx
sAkssVmC53AOv7TM6eCweW/UjwFbQKGWNQKtvCXqPm/usj7Z5TXsZ8AtjSRmXXet
oXzNqJvBy02SX5fEopK3wLQlybQZYB30+XatU9KlBEh1oMQ8EFRJr8+BMcISB3T8
aevCRJix0MY3ElhW9TI2a0VtUzVCiNbBPbX3TeFP5lRds9fzNeVTiFFcpQity8cR
XrIbM7DRU0Ak6QTIYQD0ssRxoQJvCFxw31WyY1JFSBjNLjd8eVHX/5TDhz6ShGwJ
DqBTYq5MOkNqzO+hrPcs9AMSoUDfPPhg4SFKfo3wU6I2bl0CWgrQQ9gD8QPhBG4B
nWvf1nz+5gaWxxi6J66l8iveFKJs4mElMeM/gfZrNCYR1JZ+6eJpuePOMw4vYj/m
Nup2AOYnfbmTefdKKqBv8gACKhZQLMws7w6UOUfr6wtYBCn2CbUxKOdlVeQWI4ke
VHRmimZI3dy0ttxAPi8JfcI7AWs6mlJcvBG1+/8D0vtRFE+sMXV0EqPdhXI59OPD
w7isl8rxSrMIKVpMxB8LsisGfGpp0sBsS/LdUN/Y9YtcDHU281ZUv5CItP++dMbT
an2+DLKCfsbn8l89/qqwCsEuasEf/s5pzAKaUx0ihBpw8m6NCodvpr1j8mgLrmf7
7jvlA25B+9ISDldFwyZkGuzz1SnpYR06fQERM4o+0LFWh0JcAbbj799kLSvrR90D
hxVLkkBR230PXaC40ND3aA94x4ZA4Si4rj2osVHVjmGjRdcxOc3nuWoZV7ZW453E
1SYi4MxbvyILF8bhBZ6Jkx5r7gBgoJC0hg3haO66bVe5/PApNulzmcpzd1GSP2fm
ZrEQmlecgppqdgEDmIcbk+IHTJTSRIednyZJWhAPuVqzMlhh7PkNAVgGl4blFSVb
AdiIeaxpKm/cNeaxdWsp90hrIy+9bYG6bFVkV5iLeP2gk5CLiKQ1/RP9kMkBx12w
UszO9EJ9HwmTMfJXNBx6zFvMx62PoRQC6pfMZ80hszWNTgoehSNrqDkB0+gQakOP
8bBQwN11H+9/XkZh9ECxvKA/Oy9lEJxqd8PniHDNEBo5jrYIEJEoWl9uS/tNF+4g
7HU67mZMDAHbwN2xXoRzHyFPz0AHrQas9eqpzt2wo7lY2G6fxQkiifiA4mhcw6Lg
w6v4giv8VBzBr4LlMOpCdSWImk3T9eZC7TvaRcdzrBa2nY20h4jBkFmKze0cYavn
tP1Te8f4lPkMDPZ7tYWI+r0pimrGNynbfwVlB03hfe2MjUtZubcGYKMZ0XehTaoy
WB8yrqqnesEEy4QPtZ5gZ26QRYCJA6apPxzo2gNfRFIuo17pYerJISRWey5TejFU
vVrPeQ3fJtmG8Z+8JZPtJK9cZUYyg9KRMsnyq6wnAtfXizJDKjGR7DmkR8szmcV0
vwIjF8N4SggHVHk/92Jm8VuPqAUPH6gyn1O+z8oO+rjN3eLHq6023gs95dfhfcAR
TrDB2jsnQ1gjekDnDx8N/8XzVzbaXS3kwPqjy0ZCactP3ZtGZUqebewnUNqTjURT
9/mEbaN2VLfIG1F3t+vP0qvRrvXWG8JGKn3dMeL+HMQ/5GL7Xa0SzExFqtUn8gub
/+PrqnHsxLoVJdR0cq5ZQyhQJOgvBeA4jS29TPvln2JDx0c66Z9/hdNFXhdYy+3G
Co/nJXs8Gm29qlZ0rSPtYaz/nIfRFe0uXwei2RUU02xu0fdmUhM3yoF5akXpxj7D
L9L+fIObk+SZrDyVsa2qM0M9n7+WnC1rPuAy2I/JAb9OwBlRbjHMoLh8J3GbQtWA
9ZGeuMz57RPxTOxkqbg2gQ0gEN1kQtlerSdAxas68P1igOeTSY00/6LJX2fmEYQC
/UR5PdHkqbNITrgF1tIRhxSQGRP1TpkjRzkqhbD2aAUD//rDL4xFkP+MD7oW7fiR
unWV67/4eglgElZXUquqPX1R+y8E6OB3MfJRXVJQj2rRptMcpxqQiDBQQOx8pQJB
TZ4Nq//BHLK0sIqRTQ2PC5vxRO7MaGJM++5O+sUMSv0ywrrindRQRExUe3rqbtA6
3nLXX/Tw7T+oCuyxpEfHMi6F/PERWW37dMOPWjTyb1YwHcqtLHrtBM6w97laKkqt
BmZlyaoMi1eTa2bmcCI9HcmbbQT1sL4MSpcLbyj+9tvSUbd+Wp46hF0+fg5Pz8tU
mmFrZ74pzeIbt4wX31fUePmnOi5/CXJ7dOti2J1TpwvmIDcx9kxp6SkGQfRj2oFz
yHtlpkqOt18cwyHHJEIjDtTZreJwZAX9oTYkZDF2Oubr7JcuFqlHsxLx8LV1f6nN
Qcmxm/lLcDS/q2Jh+Fzi2Ofjaqvu4gPY3QztHy7gFxxVnycHGnbLjNkNxZ8u8O8p
1MptvqHV1zlQkmhl7eL7HeZDWl9M8aNBLKIjGSncy0dntCc5swxBHaRurXCQaxng
kaVv317zDjFuUymF0T3b5eF2V9/O4Z3H5WNK+XVuwJRifo+tO0GhTQF0M/kMcvj/
cB1l7y4p1QKrKuu/Q7t1C0IiIZeigUT1uKcpAHq2xNUUWkawwmK28njTRF1UedyG
J8EBQAqSJoxgGaVkuz5ZzDPI7eBkWbg+IiaeQmXBtO2XO5mIGzB7DsNvRaKR9BNL
vRw8U3uStSh3xwrTwD78v1loQwW8N/IdOEQ7sUjfYxTtnjmnVlqLSlC6CrSSBWbk
n8je/W/24eto3QXLLItQX17BhKFR1mZRNWYaFQPJhPtwMjqKlsmfsa9WfL6aVDkJ
CblLaRNlf1dP6MTx/ppoahTtn7WIprWf6HOg1ns5PXGXqWco56jIVJIZlQUHoRPW
4Ge/k1kCX7nqT6ltvfRMF7tu+QZnjdcBNdxzlpI2T9vEdEnp3QLQdgJPeMG6ObYB
hlk+xsdwzmo7JcPUuPwK7/8q5Uc89NnYWbvrFEcw8OHzNOgeL1zLl4WbIff5YGjy
q/QD5jKXmHwMEDKsjGN+8Kj/ot+2LibBr4QYGVLQDJjTgh95I7HaFzgxyUBzsnck
HUXe9y9Uin992SFCi3gi5oyGUADUHShEuuxE8WvnD5OdSan6h4SK0OZqRrUa19OJ
2P/nhVE3d+zvDUa0YyHaZm+MMx8g50hCmpP28xHD9DhYYMVklMxztuay1kOASv2L
46qQBwkicGkwGZFW3RWK7iGal8y8QTugd/psQFs0AZD3XIGCpeVYXZY6dzdDF4SQ
zM0MnNQGbS/ZsNrMrKyzzx2FiOnXLflQPL7srmMAxUutX8jKo33E4sJlfFBXDt3V
yOcz6+2N5ECJUtFG4Aty8HnYk4atPAMcgNZwd9TwYWbxXzzGZo/aHRVKRPYq8E0i
qMVr4gQ33cCP01Cozy+lh4aUJ7D6GMMmqOV4GzSuzqQLP9X/DasWT9Yp44a4fwdQ
Sqy+JGQ2bri9GtrlLNDDvT/1Ow/5llzLPO1mKEhxvozjhFxgVLrrdYfMUOK/pNqv
Kw52hmSpQFpfPnWk35UYFkwsJH49sMNzaEUW3Dy/XbthR1JI30EQUBnehoqmMbRJ
b9xZs0FN0Sh/O9BaUucZfSaw1chiWRLqJmHOLA1vqSRpAX4BRnWmwMRDJ2k606WV
3aGYPZfh263Dj55jdAKbwqoEbnKJEPCw8mSm4DntlB8ex1v4467clrM8yMrISYh9
KvNRcWXaCw2ARrtA19w86JbbTolEy5CJdNVhGqlhnvkVwtADn1JhGkLMLYpwoAmX
mc5BEO1T8epAhMDWIMfz1cfUNvNHvy/I1IA9xoDVG/m5OSoEl0MlDqLk/d/D7hif
du4LCSXLMLIpHdy8VPIs0DD4XN77DmgItFuusk1CZvYf5co8nVGsn24SvVhrMVya
wOzQcpdb0O4syIlM1buj8utyAEzIgysTEM+U2BF3E1C0EHTdD7+f3MDdH4VICwNh
0EA5Ow0TtQU8IAJ7L/VMhSc8QF4vAGXum3q4Podw5u/AoDmQsERZ84t4qTivR842
p4xHZIRiyZZYfllefezwmlR5Rb534HECTWbmygnQHdY4wz91ZByVFLaBO3S72enS
jKxXN35zURwsTlzcS+EVhUGAmcI1WMouFsdNUyi1elN1Ktfk1iFO8gUjQn/YeUe9
nlu28Ft8aojDKGKZhFkdp03/N5iVnzzIQ1J66R2AMUJSinQnTaw9/VJpNWLiEbli
TXsajE92Vjhbh+HdZHn+Oaw0K2f3LZWfJY/1KSBnDplFkNHYc0JB1pTsGha0xhPg
qlJ27Br98WmjBI/2SqidTDZS10LeI/t22JHARKcOKrVbR8PLcDmNeMA4MBzw5eQ9
d/4IUWrVY901j9TRxikjcF4/frG7rNf5mifXLsVlUuD4g+Eii88PzLZGqXeF5TmP
Q71TULb0u83z/p2mcWWWIyH7a3u0qlxSuCqQGwfg6kVA5gQQsDjhNVPjkSBddoAs
a+uGff1LxMSjlMOMyTPgSKZh2qZnzYN7yPJ7KAakSuYJisJm/lxHFD7vf5Ens4PU
DAZrfhfLbh5iG8knZbS6LwdFy5eWRF1dyC0TnMlBSdP0YbB2LRBgt+wm7kB9FOqS
asrm94DvMg6WMClWAMD0EHu4P8W5Lfuf9WCpUny3N+H9ZJgVFJsXC9ow0uzNjF2o
fkNkAm6MuRxHFZMwvAiDHLHBZpCxNGTaPfZBOnZwdwem5FEEJVpnyMrvc9BrFX0B
JqxdC3GFJl/GPayHqgxdqMH5Z1MJkRICDGeCspRljdNL1lUk3BxS4QOkbMhg1YJH
A8TQYnZoJkGZ789smpULQrF6zAwNIFqF/JumB6oehsFLOteve/DvmwCYNtg9I3jy
gbmMsQFW9WBDXSNa1gOxp/UCoz3tMj7zdHLGVXCpBHB/RcG6veVXzMjpkLFy8Amm
SLewyvW/mALdcE+y93UUhIuL+EwSl3dvOZK5j/krrBmSKPeTl2GLGrt5C71J0Vmh
DrQ6L1uv8Wlfxo7gU6Tux3SYn+10KmJW72cyZVTiYu13tWRj+EO7JFNRzExoiZUU
Wg1eLB0SW+LcGz5UyeS6XxeXbuSyThOGeQZ9OKesVDjtG/q4sWobWn3bGwZFTqok
30bKCxFW7TLsyZyaMOWyjSJzToQYfyOafQvELTPL4pAXE8uh6A+znmCaxqrvSDlA
ROp94QjV4X65//tbktmho3LW62FnnmfXTbIEycgdgV1Z4+NnjSII8GJFywZF5xJC
67B1TfWdapmpYySxcBmfIKlAQ/rLCMfAibC6RFCCwVJqkotq2AOfyA14SH10krsh
fOjCy0MP1pcjISY0x5uLCWpC+pmj5ewjHJzLd0OL6LLoj/aLU8moCyWbyKXor+AC
codARbtzgk5COiI3dHP1wFTHj4BHw2mgd3ipZAWKamEt4ohETGXVDmfSO+zG1ycP
LNRv3CPgGb9/gxoy93DRr69Rvn6Y83lZoTCGOUl1ZXRqxTqsSOe0s6orT3BZgSXc
rw8GMmIeIIBmSyA8dSn1IDlMFCf8M0GjcwN+BLLNl5MGMbicmZU7DHiOiecSBeOf
gNUHYS4hY+OVt1kUpDDRawoLDgF4B8bqJcXaR42j+UloysvaEatPZtuVMcuPP5q1
hOsTQ8f2khVh/e9HlTFAe1AeOTi4QDDyiOc/eupE+63/txhF6FdulgVrVFBiXZ/d
6zIpcAwxiAsvJLLKsYKtSUNkxv9T3g7G2kbs0e5uPMe9VC2/u4hdLAaZRv9UTF4F
SIcAlP5te0IR0JNSF04lVeu/b90rwwORsFRG2CtwEG0FutpwyhxFlsjL25fAgTyH
lNTjj5IuhCacvwFBv0vci07XSY0e/qhXHB8/d2lQQ5qdzt/jK8xdwS5nnMSfNrIS
PrdtbLbGB430C/65DWjtuoO0ruPtUDZSIV0WdXnK0idh4TwNeltI1TjCjwBSBVRK
p6KM06GO22ZSa/ODMCeq4/0xAOKuyVWZ5M1bO3Cfm2Q1VmwSZDecZt77ntBl+RNc
0C3qUSb6Ke+1Bq+QyTf17Uac1IrIVPFtT1jIdlruZZSNmAcmD5HoleNEOGVdpmGH
nOJNAjKEVVNcxtPZYF0weJY3SW+TY5Xn92dbEV14YhS+guh5pwUIkgWi/E1nkeEN
tSq9N2Tq6f9tLmBuLD2ByNkgLYkFP+z7CL8Sr9fNihnD1JLUazqCn3Kv0twR69EH
5I4xIiqS7QM784iM5stJmpRvlvDGTRIK/r+yhb1JxeDdSXf1VRnxz4TaCtWt+56T
TumkRjYj+7elDSEWigOrgcvDsJE8SPnCkCmx+1IvQabMhKmwA3YB5exx8wQa+tdN
vv8/6J/2E+v+jxzEBgXit4gLzfqxol4lSLQFj5GUNClKAXYOit71DeKFWMa984dr
N4NZxoM27MWLsFTV/oKt3T/JKZMnFl887X/i93o0GwyB/rPHNOFoYsY9E15y9Fvs
YXFpnFUgmSjz8jReQ52jcNh0+LxOctq8XsHfHjGWflDJmpAdYKFaKuJuAZceBvbV
B/uVSNx7sE5wnJD/8vr35/7TEW1xai9oZktDqF2erb602eOEA28XzFlrwHMdNcZP
1QIu0u6w2gF9D6HqLzDQwiDJTEJvTqW8edvGU/97floDuQvha29pjOOWcYi8fF1V
btyze39K7X5SfzHiIJf0104BkywVtCyJk2GuW944Dzv1FuG3nRORyXfb76DFRrm8
XXWqO/hLaXCHkDQ4wYwgUN2EGhK0HdZ/L+P9uROsqA2xP2rGfVhvv1FyEr8tkC6T
0s57LRW5muogWB3+DKRNKZxQ51IP0pCmzi1toKH3Vzk902EaWcplL0zMXzyIlc/n
LhELhMmG9B0gvSPY71T5BY9GwmaoESYG1ymPwKbn77gm6g6iDqfRF6YVp6ZTTN1t
YyLy8XmZTuHDyZJmKdw2mAA5GtDYtdWdlyhGrrAewCm58ddWgkxNe/pLdqkDsPTU
q/DdsV0rRogqdfzMJ4Z1kDPVLn1DYI88iKS4+pybj7KPSoMn/BK2zk9QNygHyVML
K6Q8tGJSw4XDFqb1b+3FV3XvObdE72gfgcPH/T5p7zMcN/7idktYKDwCgh2X/YcP
M9BXH8KisXi1yld6Wx3IJcCXYzhYMSxLnvRmqsZUFKWKWBQyGFuKZgkk2ZRU9isO
+Ynhn0+tG6hG5AiRdMV/BMmwXTWELCJT/dDvOzAnKfE6He1w4FnRkaMeyBO/oZX1
4Pkx8Yi4TpgIGY3/8tKoMfQyWYusVxB/JuCHjGw2TdltNjcrQr0QFyVNADj8T9GE
gW3hZnYHGinin+H9a7yyhR+gtepcANHeQES5U8C0t1zggRd0fr4VFmoY6Sk1th26
LDRxQ99KvCzlR9BZ9k71BM5Lb/IiC8zJmfc7UHAUuBWbtvZrAe5QItTNuV+UG4lt
Do+agMBu+N3RwkNBC3p4TRwk0VpUofImEcPT9VgRIyz5IdMdjAckryl8M2LGQRIl
k48q3zP63PJO7jC3qDjcliN/vZk1eSuzUKzAQbBYQ/VRGLWf41GqWuogB1vNKLap
JFCzIRcZgefzy2jxtxmP2Gg+LjUUjLV/0V8JRdnbjlipCPuhlRRvfpv/UHwPxoLl
JRm2SlQZIcAiU2iLdVnkUZ3f2UwgGhbf5d8Yf+FKqSJ1QQTHYcaW/wE+v0NxLGq2
JCo6XiXqDZf7S2HOh2zq1HdAmddAILPs2jj7R2wZJLOGvRWCR2B/MaiKAMmIY4SA
X7f9y2x5QCFutckeIed6Hzv3OI7/3K2VZd86aBKHwPKocJfC9cFKVoi00y4xtay3
N4SOT6mPR/LjErGtxwfoFKs7hKQqko4HCkren41n2/pLClWop71KGIcPreX/7EZa
y9//4dKvZZtozrnefIY9iS5pBhqTsUYPI/gXl6xaKxDqfn0pCcTPd5gc/EFkIkWw
k9rzwy//TyWPSlWn4E0uzCMIT8EIpUCglFheOxw2nyFXTw5amHpiPQ0r9UeWtzTN
oGajEbwCc99Tqbo5rY1xRmde2CWvE/2UJiP2DUcEUi5kDyzCprGgDbFHG6hFDW8Q
m3sF9916g/ZdmABHoJsddcwxJIvW0UFPvHwLGBFBPtW2hgXcMccVsRCZMd2SY7zu
MgsgOzpsWRpVaebv8VsgkmQohgg8hbgQImHfKfxdUqntspA0rVeWNcZpMGx2tIqX
/gZkhKRMfBWIYLtBd6X19vTZgePULi6syYKukOavGwmAd98I3QkUoFCbV/72CQ9n
TJJ3yhk7XJ16HZd0D709sofpLLCKxzdyxFIbx0CGyT+2xtWiIq7lXmPBlFnXTu25
sVftPLJzl/+yQ865/XKgSMuuFKC4XKumNgNNqpDgCoetiPFxg/7Iw7C5zSWYuOuh
TLUkMdW98zZlkOY0+toK7DUR9Rxbt0iVocZOpl8o6bgLAs1CuLGY5C/rJv8aj2T1
+IH71S6qekYd7zev0j+e6Y2qYD1SufaMJmIfi727Vuf88Rzy/i/g+UnULLpFR2bD
9eJiknHMiZQSNuEr0DsFQkHaX1Vr6dWWPI50TEftJWCJPY5r1SlZuSJ2T8g17ojM
QCOoBV9qWAcclccrZ4crFtaodku1+DX5gkR3xwb6m92AMq0AR06jwWjRhskCKDvs
fBwD7FlW2047wDRVnBkGGGQZqQl6XDn/Rhz8I2o4/4APTGih54XdE6W6JjzvyALQ
5qQuQ0l+HHgDEN38I35KpvZK++pm8xGHvM/NzxHrhRe8PpllptJuCfIw+BIUlpcN
SGm+w62MTBAallN5DzbenXlSjd+MWBqLDZ1I149nT6e+cCgltrKg0zRLzspPJkZV
MuXztLVabJrTEPvEXA3sLhG1Sk00vfcqg0fPpIh8l7/j+ag/HBlkVjksPPahavFk
gTiEiZOIvhuB3wtcJ1d7GUf/0MQCk0YofVmRuII4xDtGUVODrxS38Zrxk3C9hzge
JJOJwhy2OGuYOEpzIi00F8M72P7Tzvx7Up8RLuH7BrnKfP8G5GqNvB3dwE/HDx7o
WPNzeEUu/vWIqHGHIDfrLqqONrtxOmNHFuR/TpggA3OSOzEC76d4260pi+0VWWY9
Nc/J2gLbfql3O7cKvC3GFIe/YGlRpIS3UEfw7VoTOrdeL/CNQ6gBpn/xKwGtNETd
3k2QXmiU6EQZr3zuj2oIf5Oy5iyWRgEk0YUQjKtWyEKUbUFWnKvjvlJxa8ycuUIL
xE8kJnCR0WGJh3TeCcfqktmi0cbJ2TYwD3HYRjF/WV6Xu7FnxyheDtN3GdhJtAYs
F9gDx7fMDdE7Fau/mJyajdQdmAmOrDb3b2as920l2aJkTzNh9RJEAjJHL6tJ+VdU
OWCZH38xFcbXuLUrKpwzGMCiNud7U97lTlryofnzI2hpj2/t53DOh3POKAnKuVL8
ftWwMpM1AkpY2veGntotW56P2srOrkX1g/TfLL8Y3yvIWhjcw5vqtW2CbxgurfUf
BA945/HHHQEfeWXQTUdkfMwHHtjXOhlzeZcHv1k9Rc3A/ODLPD37n3ileOX3zFJ3
t/pO3AQoTYlC4eZV2CohWWlyLzEXs1zvea65nX196xOaFGyPHYH+Kl4MQbW8gxnd
lIsmi6NzZz/gxjYHRVw4QEoa9S/ILzOcdXnbBdHD4kz10u2sUlixjk1y5FO1u4mv
jAuV6Falp/Jh9HozW6IW90r/tTNIgQoh891fUBA6nc4WzWVn8ZOkZshU31lFM8oh
dP040k+HNgZ4wTFxyR1NcfqZ3DYGZ1IcVLzpLowWyo9T8D4DXCJlCFDQvhUef5lB
mDsI8VlRSu6K2iZcIESb08wX+9ZXhg+ckKwFVAaTH2piffXSHZgCFSD19WDan043
hSjbv8CIpGYAZtTxmhasF037o/cxEuifpSilbqaE8wjoDvbt9hk/TR4Kqq7RDM1D
IpS2G394WZXsTZVU00D6IRQu5si2m8dP+/bHvdRUzdJvwFa4YeuqvaveN/5nij9+
FFwfOWsl1XjhBBHiRPQBuKwfy/2ZZW5WL9aH/1s/afaFkFSw8u6TkOy3bK44CKkj
39rWbUo9qZn6jIE5iJkr4NBM6bTroUJQClYUwAVnPGXfjmuIKEUcCtRC6x3CX6B4
AsGEbwYdE298mY6bZ7yt7YbfL1byiZLl6JDJLWKWJJn46b2f8Izy7RXMPU1TmgrA
hzI+RbuVFJrZbNfsFFefOChPH03FMqDK6kWZZiuBI0q6Hs4GrIQUda+ozRN3pnHb
UPP+oUqUu3jNck/33rxd1DMilhKw+kVop9JPofg13IVmW5kSEHI9xZF59ab9QAn7
bMk1PZc1Ckc9vD3W8iqMsAlN5HptUuOftMscRasBaHGegHB5vWkYWRjaKqnD+v3j
oZGFsikySENPISUkTXiUNLK26E8DfSFgZ+5J1iywf7FRXDP7rH90uK/R3EJt62v9
vqq1zKh2W53L4A1wSpS1TE/6nJS7sqLO0/amL0+FH/UYHStWu3IZ2zU0ljA49slc
ln5WFRjuP5bGXUAcPxDSI0GTg9+bs89Ik5dHaYOQ3RXW/Oqy4HIE635+DHWy0iOt
Bth/rm2iXdHVen517ZA94In7rJBqXTBDIPP9hRjcpCryvkSE/oRWACd8k3sCGERY
M2n5gGgD3GC0pm5uMofCAEhMxBetnKEgw/xzISGySdsbAhuqzj7SHoHJNN+PSaiy
YpDWQ3q8wfG2Af51TIY5dWhuowNZido0yYA8TnVTNacTVUPUotvd0cw5GdN+0lIt
DUKmIyOk0wmMg3MTg58/rJ2MnxnZe/fVg467g0o4wS77XnPeDwulcAEkuRgmUPXA
tq6xOvteqTfq2GUw1T1BR4bgbxXjWw978gP8SNrXhdgbH/xlB9H5w482IRgENbFe
JvA4VouV4GH3UA8GekJGuRvbgyEpl5B4iVReRcxSYYCrXzpUbo2+X8YTBwepQh1Q
0r4tK3Dqzuf+p1EucvA09/OdniZ1edfpNmqAJLQRNMI22p6g/36NO+ZpUQD/vV8W
NgII2EWXOw8vDhOlo6wqFZQRf5iZjoELd1jq2YienbhfkpiAKUnqtbjbTd+ELn09
q5pYjJzlaOgtuvUfu6wyy72zi4f/w3k3vSqsbq9wJEyZjSBH1wFXWwtqUpijOvjn
KvY2xIKDX0I3nCWeppM66BaQEowV3+77z4UMKiEK7i1Z5lhCPNFDRmV6izGsuy4s
+0VoTQybOZ2yMDXoTsD2pGsvTU6CPP+92qeFBMwTtjVW3Ujl0PazzIfRou8xGDDK
JJPjXI7xCgQ7tjouMf1A7pvaAKN831rsZVnv3AiHc8AC6lkRQ+GOYqO4MyFPY62D
BJ6qXV+TUxP82WHf6i+SoOMAbofzPL4Ng2KvnyaTtN+zAqv5ll9g32E7JGXA5bEI
Xa4YUVe1ysxgEX+BTpHVfwWLZuxuzVKBJjn5h8GIV9RXXYa0xsDzTi4RdlUqYsGR
ddrMXdUmYnH9RgYNNNSiPH/Q+bZq3EfFF9M1ttlM0C+q4u4Tp/QT3zzqEgY0RWec
lCDvM3ocwPFt2st+TZzFVu+eL9qz3SkU7QpkqtdyjBpP0zziW5pJVlni4QpCo1jz
OOHOhVkH7sgJyjo3U8Jrwyl3m8CJe9bDa7K+l92/Z4TLdGyBIySq+kl1A75WkSwV
dxvCnLIiyA5ItmzDYB743VAGbIn5JTFGd1buFQ2TcfPHScf1IcVxaMEzSWu9/Hij
6WBEJs4bdQHzsAS2HyDSaV56kNEAPUncR+vzajei3QKjOQZXRtHy6l6qWczYlLOP
uaOPFCRvZ0uwV8f6zEN0tyR3/srGBZZj7TRYpkRsy8nMo0RBh6PFyRP6JQvmjZ2T
xyfQWEIm/G094vMpTWq4HTVelNI7rTkISvxTdgpnnKugOY3k9VnNMcoqOirGqQw0
rPio3w/mvYUxyPfpaco/lnczw67L5U6/Oa4xODUJQyh1H3PoCrOEfGo71jnMXcPU
Jm0K5F/Q8S7tibgb2ZMn/bl23Yq36nUaEORsTgml+uYhvZod5YkPU3pqsFSZAe83
LZpB+ug1pA5q+0U0X7DjYltW6/5blqKN5rmOnpdcrwAZnSG05CVVy1RnkQSmmGCO
J18arcOZaYz4cFpOChq7ZVxJRwCVQWzfMvwsGSNawSdarPGWxDeuhvNYRzF4HOK+
jWouhYZTz6OLvu1Z/mJB3KWWhUeyJCKyGkDaL/GZXr7d3vLMwMj7W+y2qgFNwoaE
KheLkRdMmFCHZ/v78wz37qYUA1ONr4Nu4v94lb3HDML3wvBAkURfm1ef/Pq4hIgn
C/g78wwAE5J41nexnZY+Muhi8VPy0WVKy1uvFY6z+N97Wjub1ZHIHy9sLJEvowS9
atnLGk9mGAZ55SFSaadrJnFi8VXZ1yXfxFaCxU9gVmidHoRmcj+aUocYoQg7nGau
VjRQmZgjtnz95WWeT0XyShsfqA1+CJQRgmdoB1MUPTLDF8rCzMQvlVE3drNwJb6t
ywJ0zHOd6F+kNZQh1u8VcxkrlqlGeq4K1060s2mcr79k6EPLoYlPm1vsBfjJg94S
GOP9mSOyI/qsybcrsiVzJlgBCiiuveUdN35AvXmUncfoqTojcUXLze1LJuxH3zr0
wrvHZ+HzGYaXuuuO4Rf66w0w42o2Tp7BSQA9UA2zfabq5Sz1IHnvmwAkMfTf4Cm3
MrLSplVn2Z/BC73ePzO1QGztQ93MBA1r9ktnCR2alRN+uqrj8jXTlr90Om4JH6u9
9IOGC5F5GZNvr5OLmRkVeCgTn+yn9m0vwVYbEG6qz50gknRz7sLGDdgV3DNv2V6T
Feq4TpHvba5gEj28ktcivQhLqfE3UGeCudsh4kHUc+E2arvxGMfy9UomZvqd4Tix
+WlLokSGYd50IaTOGtsvvrdd41zNlIwik1qCdIwarQO5two4D2k9lcKfsN4lilGG
OOQBebTo9t60hrIDccxNBzQ4gR0XJo5I4ydyMGE28gexWsDVyWStCd4bvKbt0ZEU
vnmxabHW0gfOcrVmn3LRVtrAbBuXV7EBRFWZNbiR94xyXRv6lBlLUIMXJueGNjHb
Aaxv9z0+VNSw+bTrf9RBzBYaWss5kWOvY+5xxce4m2f3vMOzySgmGUpy6A9Q4AoK
poILHxSFvBmQeF3QVfESyR17o0pcJP2R+lUAypkfyK3G06abs6RRA8YopQ8XNwZE
h6KZdZXRN02Ql0saRPzdNlYj0ZUMOfumuaSGQn9jqhzPr/UH9cc8J3uKN19m3uwB
jGoVrnyEnddVYB3nvzlFSmwjkrdRB57tWF2TOt3cM/0v5OvjLJm1k/viQ9t0U49m
lvue8YfnB/4/Ce0KWuyPIbdE6vGNHAPqbaTCJvgtNJ1RDd0XSLr7TbPdSP0pWV7s
n7BBUyUf1BuKXi/hQb8TwapQKhajTfdUqeCRloLtXrezMgcjVUSDRTxQF3uhyz6P
FyHozYhafYlsJHDCKn5RBK5pHzMugD6uMVeejGhYSb+pb52hSN0mr/wjnw7ujbBJ
ekTztIax2wLBbA/oT1GWeqlk0DiouCktAIkjyFfMQ1I+/6XCi2iXfho0HQea2YJY
n+7XeyUUhuUC36g0t7IwrB6QZVVHQSjBilp3q+KYR3LAlQdN35K9/8IMe6y/pX2D
Uo9zLhS/uCliGVjx5lJvfRra6sktq+/qiE9sZm3pdAAevCIs+UTEy9biCa0TJthU
4otK/nakBE/dsAW9ltEBJEDjJ6EY4MB9kYfmxChfU8OqpJj6sIzTFYxVegQd3o0Z
TtV/buj/sCzO463sAL8RfEC0xYMkCqnSFQ+JCe9D6d7a7AHjs1m3wDDeND+NQyJy
Q3ApY2/0QzdU4FOtVWfG6u0UuQr5SJB2o5c2cMw6FHgMGDIV/6MpQxe/n3+FtwLa
YKxl9GxXhRkP8j2sVdeHcfp66veVPY98SeGKSRd5duzfD7x0+1wTievroHFMHEcW
an3W8rB9uV3nA1+aSm08UEnrrcvZ1Bu1QvjAikZUqsEL4Sbf2fX1EB0UFWfOLlMM
JU9kiBiehifosUz1GhEIC0tKJTK1+7AamarEXVZdz6gv4oPQeARVtNIgbHhXHhDD
O51kq696aV5QJTQRduzuiGrM7LfR8KUgSd/+VJ7rWLBvf/OfKvdzacMOCExR9BYT
tduSckXK3eWSRsX81NhciWN+YD9VB8H7RmWOk7vxrd0lwP6B9EzxL4kpQVxDOrcy
cdYEfMm5KEp856h7glz9b0v2UkN8lfb3vML+BGJOzrdgve180JEclZuS5K9Wt7xp
liQ4WcND/WZnCcFALtMoZ4DWaCyQknT4Y0l06NtYKiU+DOivCZhwwhcwpBazA4b0
SC7d3uPuHsa3Z+twHheoJr9oC38LFe4vAWZXq1V7XZGBoqdUC8UUZry9JibtakW/
cEai6vB5OYT9kgDKFj8TGXUNV9JpXJMQa/5ATZD1CtxKEDx81K2JJdXV699R+KYC
Tx7Pxnos+3SIap02krCnkkf8mWNJVnTRksCa+Lzitgzo/qZEtO/Rno1WiaDjTH+n
uTGon/e6Im8w8qp9w5J4Qexbw6fj9M7otOEt8atDX+vkyIppR7+BgaGBvZvONqWF
/Lw3LBrSXN8VxJW7FCatIFNQePwQQ1Bd7oh5qSNyRrJSm6Y5rwHzSjMAUffmddW3
N5FrWK9sjc4Pccxx+l8tY2k0+QTr/UfhuLZCcZLSqRv7PSsouH1FL58lEaitBVLa
/fhJlWqfYgkNNtuzg2lr6N24Fypdvob4Op89EcSsdH9Ovp7lHON+51Ab7DngbcK8
2xlsGQZ6FvlrwfHYlJHiGiJIplaFqpa4KFkq6GvvcZCnf8yJZs6UR8n4OE69YFle
Y3mV80GnYbhwdsYsjI7CJmNjt49KoCUnmnG9QA0TivBIWz1iDaL9YWSJCCFfUFT7
vl8oQ8OBWxKHH8jneaxdy78uQ6JheEenroNv5aYtE97ThTLCcbX/cnDfsv9gRJXH
HRQ/yhuTfoOE1mbMiOgIarvVqpq6lAi/VU2d/vbjgQQ7oLBrGGAJz+xXGZ+TXioZ
YGyjQlQM0D3mIkgiZ3CdTEUh4h80FGMT9ucWJo9sWWEiW1wNKAmvpC97bkLpqQbI
sKjnDuLhIcvZhkil5VQh3U85OA9klX3OuqrWIA67JnDneOiA6SZzH4a93L2ALNh4
xmYZDd5ivbllr+nXgEJIQebuk8kxnWuUqLy5c4+b5xXPhpLw4CB8H4mcA4DYL4Gy
SfilSlHcIYo2jTC7N4c+xwC6xIcAow981WGyPdTrtZ3htRkTpxfSPiSrfY9e6d8B
gOSVlWqvGty4r+s+4gpi0x95NgdfhIjWcyb5GAoBm2jxYs1jOjWj47bU7oDnZ0TP
mWFhnuNeAAviAw1qU/YHJ/SlWMRjH1LslslJMbWXlVYCAARD8SRm9JCB+46TA7RD
zEaKCNY85dPvIT6rg8/dFo2uaXd85agPl3ATiVQh4ZR9IJlOB99rOmivYbGfepGF
/GPglvsYTsv4VRQhIcm6NiyEm6JZ52jH3XifEjwFJPq0BUjTrgQUC1dHIRXHdDyH
/t33HWzt5cNDHZQV7McH1TWB+acrmjpbXjLyfCbYcExbCyHYP7YlI9r64YtaKBAq
EtkTdQDz+ORZ6rbxj05qldv9Wfn/NUMsvVtGXM52Jnmx+imo9V7Qai4s22G+ltns
Th5QaOMMUgNtSJ8EaTbmujmcxCluAw2+VrCwmWX0FU3XQxtTtPjHi9ZqTvAW61Cn
SBD/uiwV8IGce9b4pW53PBoyOpra++WoB1wvo3UUfkzfYobNifaMjVToxRzn/rvo
va2zHsS7xyWzrl247jsQv1VVuJGwtPh7ve6hD5qFTnfSarUh6HEHB0OLyUt8Fdoh
CJH1gZX0NV4AcCM69BVq1epEsj6sWvVrHG+xVv6zXWAnO21FHeQ4MS9tkkj+aPsr
4SIqVzrDFz8B2bD368N47Wh07bKG3nn/HCwtT9H4+0K5SzvZSdRbI0k+lLCdG+ij
w1+sBpV46A0kQ5SA4cMeUYlC022KNIknpqLKgpN/0h6scnEgXt0MzVh1AzF7rpR3
pbe0q132ImqckzpeXnXsiEScwUzRTTMuH7tiSZxReaAy9R+qyA+rYC8k9p1U+ueE
izloDlICzclW+OWakpMMrXmAbPnVUoRtOX8uXEJX717F9CysQr8nbyvNsBl/JJDw
lfTpS/UDO7H26DOP2XcL5bqSvvtoOuf0RB9rEj8JFOGsWW1oQb7dqvX72CIGP9Vz
KWi/oEG3kV+9NZnUgE9MbWnN92EhNdDQ0mBosWqpDxJ5X6XAfCS8+ZgYgrlz+Czj
G7hfNKLGZ3osU2jbYfBkNSKgkkYIdJLDDA91KPrVIbhd0vcRVW8N8bTJkLC1zVVl
S72bvS9ApkLd/76tmXN82NTRx0XuziTggtbn4DinTTE/vg9Q3xt6mLMyDn8dDcCA
xNRIWV4vUzCUAnV+t/Mmh8vLOEzGdZOi1e8ey3U+PdJJwfmpQUFXR6FUzJ9jOlvD
do6OYrL030VjlLDxWZyYBYQZL9HEHHFZpISVO0iC5WfmlH14KjDrpACdXvAJCA5r
0f5BFBXBMh/K1SC4EEj9H6AhmrvL1ZuKiWRe4HT5I4NOZMOo0luLeJKjM8AFXtrU
S/K8r8+Cl4FyZzcIW/1J0VGXgxSqfD1Yz6hx9+yEgYmPPuTGrzwi411SvyofcLI9
R/Aq4oMHnHEa/Tc9ndFkEu3Sv8rY7X7Kx/lCKB477wuxQ1t5igzRvUB1CnfLavdb
gHPWWhn3a+jpAZYA3DTzxbwf45gs445sai/xyE9xtAJj5uubXUFiYUBBNFmfksFi
L3uuMFd7oRH77EYJfCQhK/e6DiXqP3VSNXAO493fcPIO3bbpGXHQYbXWfrIntbsG
uTu+fmGcrlOtGoJzT1vloNrPg+A3XVC3hKwOqoV3fUXa2+SAIeWxirWRsDeVTpZq
7ZAh90IwQYsgyXvSYu5ymo1nY7uimtOQH5q0ZF4uo9gl0zVzy11U9Mhzpmu7IfQo
2EOzoWQhapv5Sl906d7lQsMSQ69nm3LA1sBI138wxEolEKyupuo6nE1eELUvGpji
Bd/ZQNfSJmgbaTnJUeqFw0vXj+uQrAqvMbnaYldwocskGPL4ILIQPRrStVf4KWee
Wk9jsTBLbawWQvlnc/AUINSAq3BVxwMigBwcJjkLA8APY/981rllMyjihHLF6w8Z
QAaqaPiljoEsWvNIjWC29PDNFcTlsNe5PIRiZDneP3Zc6DoOe29Ts5RzOw2pH6hQ
r1boIQs3S5ZiMRNyf8A4HenMFi5on/TQZb19TQpg+ruKX0zOg7qwQx+O66tKcJB/
YMWyUZwTZ1bRmlrPaTUGWF6aeL4DB4KmUrgHU7xKsua6BlqMEp5NWXpTXsuoKkpC
jFYct1jqifQkjHxknYAJ9kj7sl3gzHE6IW1G0NMEAdJxXJ5a1sZrFpGahKy5LMOm
XUq1ivBLmEq9fZcLrwisP82yj+FGFFLbDNyBsvJ+bKXTyFtVlZ0ViOYdtIrHP7b0
Mt/eyxGMA9imA1uprTgqDe11svsT+r348fMJBgOK8ux8+JVPSuzQjlyiiPmvSl1G
Pw9uAXnAzu7lsl5tMbJxUsN6LeMD2iC9G1SPNyck1iHtIK9SP8tU5s0MOL1+Aab2
RzniewVPh/8BmtRb4L45CeP4OupHY586A9uoXSJk4rhyO8A1BN5U/g/OU7C9KNJB
SFYEt4tzHeiv0XGIpDIh4gmpUUDwxpxEwND7WnTHK+7BV+Bk0gSh3fYiPtSzN4rB
Gbf4mP8XMgxaA8h+41Q5qt7VwZZ+IkJq1wOF7mX1JvY8PiemC8qSD/Sf5mnDtzr+
0Gx4EiBo5dvWdkFPkB4ERW2nz+YQVZHzviYYqlV7KHTjXYLR5pM5BoWQ6UAqM+j0
yqnGj9458NrzItphey/wqKOJE5jJhrfCbF7EdyasNR/o6mV3otVkGZMmgMVtZyLz
reHULdmYtX5TJjZsgGPrho8+YaKcpQdaXgcJwuabk8xPrw1suebpGXww46XMU1E3
VOtwiQZl0L8C3UlabePpD6h5jkVNmfPFCVmsAyqTrUNvwJ7/PZYsBVkz5WeJUvH4
kTmczxmcRdnQ3q8sKkHwP0q/WQDql47412RiJdRcJxyppKyo/XZKdVZqQUD1OOAB
Hu0k02Z09UxmeQpVe4mMcV9ypxuP/Xv4KvHtmBj1dXsuXTNmsJQnJGK/CjAF+mLj
Jehtb1f18qyy+z4oVTEcOAPRghr3TusXmburmQIH/tKxoALsgBiRvhYPgwwN3AsC
wbGc1gWc63vehAzAONXWvFXokl5wwz6dRhpaz795xaN55ymCTbCffZajtiqWayf3
11I1g3uJWeNK1BTsAPQvdnpnILnuan6QcndC/rT0e5jPXs+PF7C9joaeoBYZ204J
NFNohUMTHrFVwN/9QbBvnvTt8xwsJtCgDuc3/wv+OvuXUgtv7x0SvTVxxneETBFb
DcCJLgz1szF3VeTYRoDm6ep96LMV5LeOPdvhGS+S85/KDwylVIDn+jUdQE0t74Xj
KWaW9wMSVsE5bUT3TPjj3pO4gnIG49p5wPBFWc29mKKckBi6LDbsRIB59eKQeeS2
Q46mvLYYGFSYKgnYr/21cM6CNXbhiXH15rjzFvgEx9e+Ym7nQa4MzKltGsThtssa
TXXuof5GXMYYlsI2j6L8mSosjwmt39PUU48t9ABdWGMXifN+oPmmmgs3yru+89kJ
iGlQDPVDcxYAgZFuUIRPfolmTCO8fTRS5HD4k9etCw4GqVl5O29Q7UEoQFacVHYe
kZY4u85GHj3aNfmGZarQws9vYaylXAidPgmqvyckXgzIdq2n1LA0CdSjKuK0ywGD
meaVlfcDJQJ7yTYg1wbsA7CGmoSOt3T5GIRs8JipaSbEWtrHuoE5Vk2HhDUTMwaZ
bIi0Upof9SMnUIBRBh+u57lLhVMIG2FoFgdmuuAh07mLgsFBiRPnD2Pz6AI7Uj2f
4z76lRLcLmye2yaR/6hmvUuAuzoi6dnTaHtC8C/EzedtNrVxu7Xp+EjMJVDPTQkR
BKsmxpZJEn1LcfnOTBm4NtaeaLySQtBAB8E2HfBXBD7tJl+VjVFTKSbRiuhkpORx
VOvwBOiTlY8bZbRwzuEterCAl8h3GZyNwhT6RhBDDA6SC1yRBO9wYznSmV72NX19
nkJHxFwrnK527GMTC5PYxjtEfBnpUoPzS1tb4aCTV/1gUcbuOOZ1kc0T8laxKvzm
b6P3K3dJehe2UStVcXugDoR2k/NqImCFYYKsQU9EzE6r5WRQ9V1H3qfQcSr7jNil
L/lHKG04g012ibpTX+uqIN9EVYfUJC4BPMKeo94Mv1x4HOZ/RECCdA+rsZIAOE0n
k6Gi64Jp0vVxpdNG8WTY7D92gHjYDaaB7Q2zioRwhkQqV0nfYtjlGWIDErY+StOZ
yb3jORLaO+87jRzrxLchXeM6xqzxejwnPTuCOPdaABS42BNV/N1FCluXA42Ps/xz
qwJmG2i/gYcVvOVij2e45Kza5nPIoZqfClOEE2inxCJuQc9x+wILeeayiBOmklQd
LIutzH59P+lya0TwwBmkoMOA4m9/vu89m2XzhSokXZBAm1EXhavUtWTDZ5HsiW9h
CQRK+CHLrSDZpkcDUHguajlNKFZxDyv1BWHljhPXK7JjNTQtIrWZoyouDaK6Qrwh
Yie5vl6QsdEbITBsCIsz46DkYsps7SIPnetdJOGsk35QP+tvJTkTt5s9Zntb2V+t
5gSMs13QVruGbycSyAuWOYVs9u/ti5exRO79EbG3UfL84BQzoYbytayfbkLM+C36
qAJ9MolCYIbQpz45ZlvNDfzf5UnzXz9UVNW9qwZeDWyWx1CrI8vDv2zCYIP1UESW
Tu13ou+DDZgbQkNJprLrUoMTJ+OZZTAIpeEEVH3Jyyg9bd9h3hTjgo48xM4zEuW/
0SPPScPmdqwdBgmlHfUBUTm0Hmv52L5K39TlOubcNOueVqjW3pOMSoJB6+GwMY8S
i0QMmdMHr++rMheSnFFghOx0VrhHX+2dmH97z5aMoVUqcKAQlGYBPQG/mhl4fUiv
fV0P5/xbVj2Ogc0ny/DOgiTfqFPIY2bCZSyemZEAR9ZZjtiEyfe/hLd3ZtFCuiFK
rUB2dgu06WXtuskO3BZeGmJcb7FuwDSLDiWvKtsgRFARE8Y4+twWmuVgE8E0fT9v
N3RKlZoCTmuNvcCjRPgEH0mN1iH6UvUUv0h6mLDOwSHkOQerRoAcpavMalZYlqKC
v2ZPY/LJjd4RCmuvtpCLNC+DF2Pl3XOmt9Rb02XxEhj2F8wIP4rtS08X3EVMAAMM
bmnt1RGnZS6reny3UsnXB0/F0w0yMo2MYVPnJnLt94LJkR8CBeyxygFTlhXQSQeo
YCSax0oPUocKupnABLRLpuFt2TfAavfM2f/G6QEhXKmnaQ4PKMPIMzKf+BgWr9bJ
9hLExDHJOkNxRwVbJFQF2/o6P94IA3s5LjkUjbo7QM1BpFomcFBmnbTVWL4EogK1
fdmT/kJyBPsEcIcifEj4DyySUsmliNkGBB27pLk/n1oX/bJHKfQGKeEaXEbxsIiK
upizV47HxEz5FX0Z9DWLH3YC1M6bn9xKn/t3fjWn/Q3b8EzHywVaUNPAPqrQHAIn
/FHTXj721cgbpkht/G38VJbj97V65r4dWW6KoHsR4sK9mZu/wQfTmGi4rQ0g76nZ
ImuorwFUvdmSWEMAH1/nOrRLyPk3mL/VbY9rmt9spT+OmuH5RFq3DRFhbUWiKZpc
DZxEJIa0q5+HSOdhOryJhJvt260xgQQ8Al6YPusfI8dfi2ETIevOwS1fhMrWr/OF
4/nXhaWmnY26ESJh+t5sw+HbDRrikPKZ5Zgwg7MnTSNYkav4qJ0z12HwDeWmrDqB
A9loqdsxgXU7NXZgwWbdY+IuVEtffuVaF5yjiEIwiS/t50mEbzMxbfdlJpDubiOM
FAri0m1vdshh8dbJcVUGQUSS96q+rZ4MrYuqdW5wRJMoKE8VF/UyQBwOqfDiGmt5
FAVwCQzaZ1rQo3uMe4GbAEWZJIclpKsm1VrP7YsRvVWXm5cvAPChBMEUutz32t1D
gWIV9GUzJRzMLrQZAMh0nfd7MysUaHtcOZUH4eBKsJj3P4ca8nk3ttCeoHgs8QG/
QUaOCIj9Zm72Lo1dzwS6u30afHtATxx3h4EWQKPGyO8p/E20w2gWILFovYdm/ava
Ze9pWLfcJYcUqYvDu9VD5U0Sdt0WYO+nJNFbq0QgGHiMITZBkhZ6SUAoKmiSi6YA
3FQyokcCjp6lPiNdepTPdVWUPSqumJjVs5EmZ/iPZ0i6lfE8jCY+6ovXu2BA/eL8
aEYo8LU5NneOu9GoTXN7a4bJqGaG889C78gn9tT8GUEKKsqieZ+IToTSOR/lRdDZ
Wwa4Scjf9UZo8AklhwCmp59sZBCzEVJaN8oXhNTQ6/cYImC6FqLdLjRqPNYb0Q+T
OxdG6amwiVb3EPKpxVL2L2GdnoSAzZ5/eUqgedWnuPnZVSKj1Qy0nN3uqcutbcxs
wC9hLToB1i1jxFUow4jY69ZEvxeTlppPhoyachY5wgpuwOyqwlwdkRBMd4S/Xz00
jHLVRWAf+bFh9QaW7xfvgWRAakZ0N5jjGL36+TmoNXHcyOAGUtHPt3s7CMussfom
4l5lgAE0RUPLt7u2VluczCIKTWy3vGbzYfEyBAC7ECQiaseBpYdIMryH5BbmsMih
+AfQbXo4QfAWTwAd9FuNN0fYaRbLTR8PxfL2H+kUy6O9qCOVzGxgjv0mfXlAm8N6
IJYvmq0iKMtqV5nmFEtDMPo4CuiKithp9os1ExybDgam6s1FfF7WT8B2mmegE6jQ
+Zp7SFlh5XvoJ99dlEyB0arwdB3Pk4v82gThFAY+74Fj58Pq5iRvajT68X3TNRQQ
fcxyzhvpJYE3qqMEiFHGonsePnXtK0HjEEo52fpNwHsI9/N3VI/1CrR9n6Plqu0D
spAhn5ksNkW0yiKWaL75naokE42cHEp+gyzuyqaJCAgwUdSQlXhTNYIajnctpNwu
sCbVp7UzuKVLgyhkobQwhZ+uk7DP7LAS4rhH/tFdJcZ7a46u9hDS6MpSL3AW/kuP
yUQ4peWJq8uB589b7Ms1te9uULNFSbjRrElAWRB0GH8Mnk+aWNt76aWeF7xHiRzx
AD36nbNTAVbxN4fm0z6BS5Tjh/B667f/Ur/WNQgtqZ/haq0zA2z/xgj5r+/2QvFB
bWWj0qJeZpwD8zlYdzx8WeCZJMTpsc2NREXFadh0lafGMLLDLNW1fCCJx1A9nExV
1ZBzMid5A9v+4x+y2IammspLCUM6fk4DmnqyWCti/IMGJ7R1VlOFXeiQ1W5+q6pi
RGZsByHkM9PRTPZoppoNSEEcQdGOf2vTzzQNxilhdTRiK5ww/NP+U0Cnn1Tw27R/
gfgQz1tG7osqe7MACYZnV1TAsoeJSShm6ShiqzS0SsizOHQByInNRmVbJnEf0wGF
5J294GQKwrm4/IW85Dkv1a/IIGyYl61COmPdm7Gker1fmiRLbf+qk1RerdAtvPPR
c6B2Gg3LFKHiRSMCTCKYqZ1YhNzIDw2qLHzVZoAOALb30YmZ1TBl2iB3L/xONDvN
eYbp4jVHelGAu7oNOmAMQ2MClq6o+yFsjB9ixoBG2NRoCgUh4WHzAiJaG1M7Tvmt
ar1SIJlkR3Tcid6RA01jruq6VfSnPs27jZqTKO50YORo7ARyS+oOAtUoTr+hABZl
Rjes9dsEBWAGdPW7JUBrGi5S+LHf4CadVrs2BK84wBfryhMCrnFauEZ1bBKHMyjo
oFDaXFNcAMtZULgkKK4JU/hQx0UQWEre57sbS4EN0j8J5ADcQUCzFMdQJNoWzouJ
ZvGHgpiJV/LqWME72BBMBsJE2j4D1BDH9ierBY9YKnaq/rbxkGTkje1QeWVwUooV
LRpyi9Uj5C0xkv1ZgMZasd2SyrnF/YK12pcZNI+sXTLgWiDNpm6m9EfXe7D7KLJB
YCl+noXBDxSNl+CYub8+6MHAJK1uSbO8XA6ZI8wBZcoEjKYBHgxg7zijk4SC8fsY
tF02EV6k011IygGbpMh+6TK1QzDArm63z1L2XP/Are8hJBYWjBrZPTSGN2L6PWTl
CvgV2HAB+iyPg9uE5pBwKfzJe7M8X+zVYYSpWPKlMWYkhEvYBHL7bQdEV0niiXI+
XXtV7hrLu7IBE8DHeQy9T0sZfpTI7kG2jzgFjXMbIn4VhrnQl2uu2dy5aGRTA0c8
z9qmn/WSmumFxrmJvpAjtuZsmN4gkp12ewEHaND8CVblQvty2y9QWAvaH9J+hOsm
XfYzJiWtzif7nTA94rCF1eIh7FwtA8SP3aWzKT8K2wapl8YOimM0RPmLX/9Nl3XW
GtcXtUfmkyuZQBp0TPQQ+cPcmEod6PCSunZjU42oHzilEl7an+zf1UsjwOAH/IsA
82b7FLS8HS2JmsMCAVOPy20hnzl4H6bRyUGiTRgc/65not3j47VFll2QopTTWbgT
5GtYf/lBvq+kY/y9qpJCdYcK0T1XS0YtlNI7Ya6LT5KdYqVx2qWr+jFvk+ORxo5Z
cJpoUoDgZtmidEbaCdkZDV6EnKXWpxYbFAdV4GPftCPRUFJnHyplL8pI4/1LQOUc
BTi20REEdFHReCobWjYC3rLn3DrMXBlKhMSEoLKdhp0p4x5PgYPp+bQ6US1gjfWu
DXnkEMr3eZVUttAu5TzoWiW81ZzCe9LpKIRp7jf6n2/UfDLBacUwXSyExRqGYm8m
OLDawqhPZ+zQacEpw1l17eigssnNeSLvlDFhuCH/W8HflHUi6JG9zJlOMByz2zMP
rcU1xC7gBEbxbsLSeGL1wEeJyunB4CakJKQwWL3SSGm+lF0InSDSopum0/BL/ohu
JyIDg5ffspfprdq1sqErDo8LfIB6aSplpsQr74ernUNfKF17YkwePWq6kHsGZC7z
LqOMfxBfWQcoWE+M0o0alRFVr+kWGdvPt2QGP0Hx3JNUs5quxBktCIKoqLBXz/uG
NrrIVgc8+/s9ZrbbpfZnPEe5+19VSSTSkeDU+jRmrUgfMUIdjc72HsRHCRbQNn5L
f2vbe0J4D5fwXpkysNsRWPJgSIGwvjMTSX8aVHFAcU9cY+bZsU9QO1uf5vQKzHYx
saSW1xd9yVJfLKOS+0a27xh2MD5Do1cvNFdNEazn/K/dNJb1yeWrg5Y+iCFhZOF4
fkUM0LuksUgMybxU10NOoZyd9pCq96oiAGQ7OigAvcV3rrazGbqcE4HtfKrjNo7A
CxBRJK7zBOlY0JO547aV+LMEHcF8cunNe4zBSwFBO5ummbmSmIuF8XECLEgEJz2s
fLrINRjoeCPonDf30XsVGAbYrUPi/k7t9+tSHKGHvTR+A6JtPKplpp+PkDJtk+h1
ccEerEP9mG7ZimZztFS02civPYIxA4nwH43N9yYz3iiOHfE75+3mDfToKn0zZQVd
EduZWZtseQU3JEdFBh2tFqIiJqZdi9jphwyd6+zlQ8mdphvrigWq2W+yW68Ik6y2
F37I+fzig9AhBIWhByJEriluHTmYn7lZ6LNgXG29Nnl8chrE9Ftr+wq2WZuKaSG+
H4WEon2eW5mRq/toFIhQc2QMJpnNFubFHLzEeyPhIO+qKZ52pdQU1PXAXNH5EdCu
bjsTnrhR06pI7GxMc7wDII6X//p6gwCKT52Lbv5vtOTLkxnLhPxrlSemBOZA6d6+
hbEo9Z51jvxiBhENxpzfcUpvfmK/cCTfOIgq9K1VGktOeXNPcc4Axg7QLyMQXFkK
4cm0z4jJzAfZPNoOP8zcr2L+YR4FCsLT8yDfuoZZC6IYU0361OjjLgF+NFh2589u
UqHf2t8E6WsbnY6WCToYtIgL5YdlW3Ev65hQmt63Ig4YNhXtUo6f9+bVLDM0e2W3
Ct/Cdej7JbwmaTSYvZLGC+5VIdBqlRZeKhetSdkckp5CS/55tGdsbUpWxKyk/+aP
H/rUCjFonIQcl+IZeDn2NHjmaji5nZNHULljjgC08m6UfzINxIP/Q9szgJB52DEW
PqA8gM9/wwVyUDcsPDQ5TWtGdqq1u5pIWkEpbckPr3CT7OUt7vz57P5x+SgRoB+U
t4c/eO6UdgIhXiCiYHQOuj02sJnpmLiFAuwCtCpmHTvHCV+dTa7R8+MQCIjvfEPR
FPaaR8ucYe9owK8xnXnDzkbKVQ26V2Z2GdvNTzqmchsHTaSkp8xvfKuPnt9bbM6g
eyzLgShNDDLVz3tFoEXIRXzrH8/Kq1Wccyd3O9MH3aY3NK6Js1pSm1IaNBInMcOl
KuBfJVxGENL5r8sp1LYN7b7mJ22dIRx+mt/V8AkPPrJz6RHPUZrwsZRlW9qH17LH
YUWq9FPHuYRAI8ojgg2+HWQlFniK/RJ8X09t+IjGr57nCl8GgJRla4vRkn8a2HuC
s9j3tlW+YQevymzuK9es/O9+qmcYsl3rXtjH4jQpWRT5Q4D+z+NM5YVrt7VLD7gS
59ERgfJ30JoBhXp6EBab6UkgyzRPcpjXpXXPcW+40ByLLUmeHw6syRKxDxzJjbzV
W2S/T83+DPG/bTwIa74FSahdSUa9Eiy8fO+sa9IAm/ePkQmDHVklqyF5oTzo7wdC
fmRC7hGghVNRQ14A+Cbjb49IYlpmOliispORafmGmrNJLqDAc7On6KGBAfZuxmis
BsNqA3KQ68qP+I44eArPiTm1NXlFA1YvOxLtRULf+rD4heWU8+Hh38lAzaceU5V3
fuGG12BbX8G5cUqNbq6VDFZuZ6Mr3FW7VAS5BvkhudLZelaMpn6Sqx1Fh1mpSXHs
zD7mqHXwJI1yCN7tsbJIgUDcs/wdZ/XXDu4mV/y+/tkhnu83iOX/9ab6qqiX7Yd2
x16/N/vHc0g8xt1+Jh50B4tigoRZvSNfJyNchB94Cj11V3PQviS85YD5CnLAQbm/
PvRiAjsj8xDHEY+9Dm84xsKuE3rp5eo4aRzdX4R/1FyXOlKEpcAVgF1JCvh89bhR
44K/+vAFpzC8FU0ZEpoMVzYonRUx1CRxCU1N0D8rq8BRB9UvO2gp7+UhWsVH70ef
MFAIPOoPK/aI90Le0OF9tsrZ1JqJ3nPQdSr4+mVIQ1pBOYFFbgKdOWBNCBws11Qp
ULm4y0VNwTl5/ChXp6O/2zQpJX1rrtXEoDbdUnsZHequ83EEprZ0Y+peD4vX0Wq+
OWcrkw6c+IRCAtF7uq0zLWhpSwjH2CeSswD3WgjgJrjgxtc2BMUMFwUqFtKaFJRG
5CqfqxpKwaiEj4odkacVgYXGYpwicKrw79pwP56JBwea0D6MBiOw+7mn1uL7zvWa
MKn3Xvu8tjHCNTo9CSxnhCQPTLEk2GY3XsgNkXFqKt0D3lawAbZiaqRdz4f77Lcg
uA4godhw+nNxaUm2jHaU/ijDD8EwgInDCtkCOLkTCVCb9SQqXFtTCEzioF21xWP4
RC41dO6TEd5XF8z41GmF8N5R1R+2Vfjy4tpXnJnTpt9MYZ8xFhP8O3hx4AzEy2T1
g8zgcH8LIAqKKQaQssqeVLq1G4MAFeSawEdvXOH1MmfD1xpvSjv5wiCPR7ytw688
ofhKQmLbA/7R6aTZ00QKJ7poXD15kLvMKZSmVFI4roQZN+nIZegj3Apq4mUDhzDJ
gCt6XQOKmRFZPtwysvH7izjE3a2eMglku4S2YgnMS1J9b37PwG816LdgnEBXY0wH
0rz7aSyfjHkFIZ74eJhadfa46fWdR9Ahuw3NqopIrX/UcmWTGPpLnzH+07lVFR5k
eeWcv3lNdSj9r5wiXHELWPOu8UVVD8alo3MYsFG4iIwUhqH3EdhWir1mHHt4i+kE
Obalm/n8SHvCji68ly0j4erp5YCpPJ87DDM3oCf8Hvu+O9zX0bDUM7T6nGYC2uMp
KxOkl4vcsZ3tFGe7ou3sS1uRi7wK4znmiD+ryjfAO8ljR+SdiY1cU47bmcADH0dP
O4NPcaImIHGkF2CMZObiK05aigp0dqzJrXM7QvBFEmNW2lMdQ6sy8YtKkM1fa8ad
YTLcGiBQ6GvWmUOkTYyGBSgqxqrz2UsAqysur9NrTcocrA4+yBKu1WdUwidr24AR
Id8a3m5vkbW1EqVX4/rieflTEQ/bH4fDa780B/PXSnFzHz0mIKVN55Ie8MGSz/tC
mYdaiYcCKNaVznbUy3Mr11OtHQGbydUb1MKtamPFmYa3XOXyFt1cHz0hJ5HoBWAP
vHihT5ZiJfEHRyXLjOU7a/Q40OJGNNEcVGLIqKfpsxnkADliS5cgHbxQzg2wYIZS
+HzJGYbCKvs3wZOpI7sAFxdBvtcIxl+FP+2d/827nLUlx+R0FEbqbMpirBjdYC5m
C47+EsPe8mrELkSsbcnx5Y8rdzS8oDXDfJ9KIqoN5BWCOWfgYJjKVOojidQKxt91
V2pG2p/0jsWRET8x/ZUfAYnXDq18GEgvSka++mvNf6gBajAfSfb2ZL5+xn4PHqJh
YqQS/cB6iSPnBpUJO1j6gxFIM1hPlURrBoUi3+zOWlFL1WAz1DkWOYTSbHVuvA4E
gdjj2WjOtvfLXjexwcZttfcAttItUZwz50L3WtSMOkddS/9oOfR0KImhV2T574a3
9h8HMEOaA+QmWPKC937K8shMz/IY5Ka/jIVikdD7+Xfs6nBD2FWHvteacfoAhdJa
JDhg3f7M7/y4prhWFrW1H8IGryBtFR+3U4esTHe6TCd+0cMmq11edHdO9m1OwKgB
USkHhvwVquNFYKXDBq1TN+5wPUq0IaqdIjwwYZN7gp1gvqDHsQOwLyNS7GBVEAhs
pF6nDkC40WWQWDqUxyv+64GYTxyqLCTHyJtFlFLTGev2GgDs6HMrY+uxoXYTG7Qm
Wq4xcbfPSY8bZ2Cl2j0IMxvGnzJU7G8NjcmkxhugHxSELXR69rct/GbjoyDNngRO
gaVZFJGRZ6IiMdW1lxrUM+pAq/ykZwvO8fv5vrpmcacrWguNi10eUzGnAF3SjPla
VHBzDKcm1kfBaAHtmiIMo+bRsKPipc5VHcp0T6hYmui1/ms9iarU8kRzp6zdkGKn
LIySIpcf8JXnLWvdcqKm6nOTgy0YpV/2ouP6wNyYBYYSj8lyln9ktprSn82jOyss
JZ7XnTboeGOu4yQxkfsQ1pYDbPHobYkl1bvhTIb1aXVw/LS9qJdA2TztPzuYUmna
Ner7wBalKdYL977De41HzctunMuJDGuw6ZlVKW7LamAGw+3vd5wi7MNVLz94N1Ra
w0/5actWuw1AMmqSjKQT6fkaSF3HTfJDEpY59IgOj0E8BEtnfC3+lrgmjTBIoNA7
+464syWqOI5WEbsrqn1Zeyz1exIR9UI9HdSCEVe/twTqFeR1ak9EKIW+AtJ8rklc
Es8Mat8VUYP75dQwLSoGsjFHcZCJujKQdNcr3vEOJHpNjLp1ark/n3rz6vJ1IuFP
ov/o7Dw04ziZm6U+DjK65BPtjDwgArBvStwyOUVQXL6nS5ZswWJTCUDotVxBAmnp
9VTM73ZIl3M4+KqBMFupWJOuX+MH9AaM/OvYD//qPePI0VrOx/6CtazVQH7W9WME
ulM8c0iTY5I3+BB/YTfdpTSlFqojHR1//fwG+S8C4t6Sn3BqNjarvO7H9z2LxUTP
PBdA60WCF99i0Laao5Tidx4Tk2qNlUlZeYQvsd2CqtwmWLP5z7CX/TQ71Uh2TAJz
y5auC+TRulXzaHPj2xwXFJSfXtwG+IjVbGhfysa38SMXbIX545hSnBNTmoF02SB+
EAGQLxjlDoaJ1PRgvjZsiOAHUw2rkBjyhKHk7nEvmfzAZyHH7aqlFchNJ9O2nMl5
b8G0GArDtLX0AgCFT0x6ImdsRYWxJINosq44UlBbtTx8ciWXymADDqN/R+G1Be7R
YKyzqVK6P0h+eSLng2RWGXTj2EjeeMrljmm49sKLNJSZzaWV1Op58Jtchu7+JAs1
NvgGNu9nPzAFOKXEpCQI72B7j3iF7XqdO9xvkoUzBtcyeaRWrgIDX/+K+w/5ZLKc
csU/DBj6YsJaq8WR2TQ7z49k5M40I3UTsoE19Q3PaRN+WQgDJk7pYQxfimM+taUp
/QHhmR2Idd1M/0HKZyZ9ieYznF5+TAe/MfLF7iV8uPdRmN2X817YV2dWehXPdLyE
mx0Fmf5n9lDgKdq1+ADdOqNhBRuN5bE1bmvCso/IrND3oB0LwrZMYygcpq3WIngV
cWn+5OzLXqp/BTSVY3CBjBBFzIBaVJDCpjSzQZO+KzgOgDZqPR8iefEvd2sC17IE
0lE6kK0AfaZJ+GGbt4jmAfNqN9QjzdYcFxM1ImXN7WBx4a4bJ8RudmO5avKaT5VU
kj5SEx2PRYLEnXDHk5VlPXahsSshBDjyqTZjFJotyPFCHikf8DJiEjv90v5M73MX
I98A9JFrVz7kvFxflFNzsULlSKDYeDU+ZCKnr+OsWSyB3kvImWmOdkW5afkqOOc3
Sl1SK1zKrYE0l+a5Hn/yCpKdkrhSIMlP1oWaAYaBHhK+tRhuAFyLngiw9kptF7lv
lI6S38E5n5UwjaJfqwjx+Yt2yvW731qC+qObgMc71kAWKwUyR5Mu8ODVJR4xPPJ+
+4v4pCwJtuiLE848C6BQUIpFsS5wmoRv1UapvvpjsinVbfZISkCsksG6HbdzO5m1
GOXN9AY46ZHyEqcWJIOMt1zJimRiiqbp0aS1xV33Gg3DMjCHmjQKDUfkcRd6/Dvw
oTLmyciHu6V114ogR8EnvckceHuZzTEPZeo/hxkeQhLST8t88ivArYhqGeX17EcY
8egXzMqHk2xchVcVR7rmiAsUXDnl1F5XkNF1S3Qr7NY6AbyyLYXseDS61tspXI1C
dZagH/6Mz9vumjN/XXf+DwE2hjeit7/qKzjhnZw+UemfBGxs2JJxPVNhFIWBYA96
Oj3GKEuW9weqGi1625Z1QDxyiTQtz3872GT9tG9RWsMGrtDrnzf+pTH0IKpegCn/
B8dAZXF1N9HPdYQOwqBgynTosqKyWscCehCI4x4kSdMPV82DKkz+BTog8SvJJ/No
SvIoHlEgXhGSSFkZhXFUNThYmTyWHqickMSZqUO+gMSai+bl8mPqoxHPIk/jTOdj
ffb/4qkb2bR+OfDtfUKgH9HzSizMRSTTvGS2rU/0QdJikk2G1qYipBvviEVrSvG4
8LIUSysUmUC2DMcz3omLkXKqIkIh90rmmdveKhN+5VyYw652wd/olO9Bs4zLZjQo
LzZafHpvPNCxeOq8BUu2N3lTDfLYfCsxpiZ/Gm4I75XvztVbyGU/Ewu8MnhLZ8gF
z8+AwUqfmoM9yUshl1fFnUvSc/II174HGT2CAJtwpd6qDY6u6893dFArjaErLU71
+XzsQ+SJ900bWxHGnFKD88s3HgFb6y2Zq2BcIVzHbKYsejGOMStKRb3a4zEWz49v
SG/SdQB3MLo0YOhuwhmlXeLokw00o/Cey7XTGVomwbKq/gMDyktJ52+HCtYCJgx2
laoJT6kQB0UkUA9CzxDe5Il5ycKZ2WJ3gI1dhowfUiJolR8lJJFIughZhBymGx00
9+Rg9AZhIyCJ0+VOxIHlhQGHjcn1QGbrAglQ6pN+kEm88Qpce8dGPZxsM6y/o5dw
HIfubHNUN1eBVs85wNx78/3WK16fgBBYv66+HkmbCtt6Vn7NpnRHGU3j+g/DeZbr
vG54kktRW/d3j2UYeatLWybNVi6hl6nR4Ehk3AuI5Qega3B4l/266hgOGggBS8mK
YocKaqhXvMQjwRyhkioVXTvYpNY30JxhyIn7X8rVpGCWj75iDTnrdrB3E/nZgVgH
lRfoezjo+ZPpvwqaWMkK9MtZyCsz2en8zQ/vIvbuJVgyVexnEzsGqAoFp/BOcfGy
e6NTt/eK9sWuD93v0xbjcjoOIzWbiID9WbxkbhRId9vzPRSW5aXRUJ0NDnB446Uf
gf3TQtfBsk08QL2o5Nk73xVxx+hgi6cKDxH6ydeSqU58LASBBJcNRv/n73/iWyM6
JkGulm02TyXaXqg5fQqOPcQ8g3wcu00m4p31qFT65kr3F7RxxGFbQF3KxdxyIdGO
DbWoWa+FJHlL/pQKTmm35MiWt7sqyyF2LoyTpfnleV+vo76DWCxRDYtnaoN53ZJ4
VtRfQgsT0/uDqirxJZTjwFedyDPW66Qj7J+umMHhxkmC6bn1IpTD1lmY98cNmW2O
hlKH4USrW8OMlLkrUUoelQUjDRBVRt+Spf+6EIBw3+skOTSgqbY+Jg2dc+GeqGNv
9+J7OA66CNqOL3QIszvGeHu6g6uS8uS4WogTGTW8qCo14qWifU+y79GsgrquK57Q
k8kRfIz94oANgILPoOkZ6NstXjQlNXdevj+hU/ZKnezXG77AOwQQ43E+dLMhCiWk
ZlHLIeIYyskNFjBWasI1tBBbtPh2+MotT7UVMH2hQ0mRl1dCmDLSvBzkVsWZmN2G
1yKhGnDFJhsSmhcWzzrVUphqvWfrYkB6KNMdhKO0KVj1ALniEtuOxClgxdF4HjEI
027B29kcLGm71P2uAxKcDHztFLMHaKe9DcmgPZCLV4urH4WyiWIz4OVxwydVfLnJ
NGV4QycDNuxsRPq0yW4dAixL16Omp2fsmKjwd5cYOVzybANvoEt5Eu5kY5PLHHSV
iTSoOUY14Dsj4dyqO6w8leiJ60jkO61HphesCrD3Iapb+ZxwUXTn7u1mkZhM9WRG
LVtxH3Qimnxw6mXg88S6GwEG9tzSqEQx7At1vR6dijGIes5GJfXOjsjMbs7dW+Z2
Ww2i24Ib7jEBx/wxTv8s+w1LZy+s552f/hQHrorhzeXWligDmD5EHsURnY9Ejzk4
WwYjNI/qNL4gsmoEHUpWQGwwjo6TzrIfM9BVjRV7bR+nk03LJ550jH8A60cjR6/J
uZpUY9AASaiFXMPa3zSSIw3q/K3BDhNNz1D44H3Y3sBqxCmitiobgE70Tx2IV1yo
wPVfR9hMb5P8lo6Y6+CSj06BkIfM3cjE0L3dCQJb0D5gp69hcH159RFy+DAJ2O1p
fIO2l8BeRkHfby1WmTK9LTAebFHQ2+g0mVrLfcy7HtNofpVjVZFK0sOQzI6skAGH
3mfltbrqSbnBLg06iKqZuMU5SldvPWDyUOvhEaZ/a1ECI6LSGUuCcTUvWjwK7C1/
s7nsZOl+wuuZUATFmzGY/MH/ZY5X+ttqN7ltHN96+YJwCVt8NSOPqDpNW5ppwPau
z7CC962FRPGypd7US2sHOwYuSEWOny9jWqcx+XJ/tAHR3IS8dCrlHWWXB7pmNO/l
RhFu8iP90wt3y3hkjV0LLMIv8b7qhf4Sc6k9yEd2bTN4hBgA52q0wJ3GiwlF/69B
KXU1zp5Oc0sbNukrSliacRuftBI9JoXMwFrpYyTws9tkWHUyZoZ8sLKBAIiAlbGT
UAEzziatgOX05vtqnRs9tWo4UXTQ6bwhj8QqSPhE8z8oIN4rhDrXo0RfyCekMvtT
uDzetc1RYUJp+9wEoaqSoDdPl1OmwPubtAv9e27b8kV/sfd0w8XNSRhCc1uZBhDB
Xoa78jiglN8KB6gOPCYlfUeArKZxCgY8bYExWtRXGr/ABEiPnNSV3vrlel8edyC5
O/Ajz/lO07UXfegJQNPB+VGA9unaoW5ch3wqkx9UptIxvHtHNN3/0fM8tHRiqrPx
vbhk0RQw8aGOBd3c+mOtcdv+KWo2+0xtSGcwFE6w0oWJqsRBDPL2i6shykK+//Cs
9TSTCMWeIDBGpdr1JNYhHiM0c+v3il6hJDCwfA5YO2GajGq41V1TsUcm9D5/e1hr
PSHdzumnnIT0ed+MOR8RwbX6G4YYTQL7cMxnmhoQ2ABoExezK4EV9gfsNhDMKlUa
US0rqooeRgt3WBymKLarPVMT1j+TQ1Yv7jRgrQz2vTp5BqGCEsTL9pZzZ/OFAX9r
PHMauDikfYBKP7IS0txfVYIHrszK8wTDlAu8k+mWlJtslB8lOHm47m3dY0P5mKJV
34Pa3BgwpXccKgE/fGH0S81HZ4I8g8L38xSJJsZQBSSj5TXUAeD6TtINIO3H/cIa
dwkL2CBkvJEFCQ0UOFMSt+/mvH19az5Zg3TnQGmQNgWt7np51xJqqxiuamh1Oz2o
8HbFMLmq15nJU21HHQ1LfzMchJB8ZMJ/6GPPIBSjvd9YCStFiwrW6d0xhUe9jVA4
TctK3X670HooKOfFKSNCh5macbd7rCINPdsDbR3p+lk9E+ippUWarmKix9SFr+/D
QW9EI7pWCWLnvfrGhl1hrbs4V19R3oBFAlCv2Rfa8vbOO6TM/LJkmfMhmrCN96pC
JbHs00iNJOMK64mnjl3ucdfcvguhL7lxF+KEyIHOCM94496fSdNdVaOhPwOqRCg4
EzWdDwIRBIAn6mTsMur9XSMaYnCNv+MI++8e+7nsVAC4A+mt3vO7k9vcSvUkKxl2
KNnXUMrD/bmr6UmVIHVCRZy1s5ti5gGPnS/kbS81TaomIwdAySh8sYGsytve/HtE
h74H+LlfKHkgG8LJV3PohYiBJg0jtkWMTA9J+G6Cb3X/N7pEE9I9FI1hWwLQMsBi
IRvrQhKRvRy5M7RO5/pqj8x91GRYWGvycofqwtWEgVoGCEet3j1MKyxum9WS1iF7
UBExdxMkzgZAOjvJnoMxGMe4CEMaNCJ9NbpTrqmBsJHQrG38f//pA/x/CqCcP/u7
7CIBcaBbUEVh+aqL3/RdD5h/eOSneMOY3oq0hZUHSnaHvmNvdp9+YexFAFmvh8wf
/MyKjTVExEg0hgYvk58PTEBp9iwATP0++88MTtGGVP40uGUXUkDaiVINPtDEwFg8
FH5ECAsmeI2/UJNSBqqf70RcX6m/9bqdBXZFSLKlFhE4Mne6Zxqr2GworsE28nj4
+h6FMjz7mqGiJA3LSKzNLlLj74/1tL3d5dpZ1IAiVaqXUMSdzvL1/tJFcdWtyW7T
DYMGO+6KjCbUx4vt4wXVt7rFUWOEV0cPuRPoB5uAgBlYX4sd+dO4/Z0NA+4TFC8i
A4JwwB3aOvQia5RSv3MleLnFmgl77ekjgKVWEkHb6UiKaYz9w5RFYWykxZmG895A
92N54vuqMvQhpeQSdveI/NYEYtaXDYzdEZ3WMYQH4xZNjwzoWyYsdZI7KHoT5WRI
TMrZe/yj/G2lTuiT8+kzuiObMS6rjTAopG0miX1JS4+L3Yle5ahTDhh8bwG/j2RV
1wHtcO1fIJ9an4M/UTVuI7qWX/dX9jCiLetfs25UDO7BewA4us7c7hli+wPCo7aa
qpbEE1KRwM/Q4ufdmIlgv49RIZASD0TP1gJa8/QNkqtHfdUQTdCHkZFcVxL253be
Xw5FSs9ehnpL2qyx6EJQ9AcZkJo7QkxncJJ+VdTucj1zrfuwG6mnvztLYdutTM4Y
RYdJjbYafIflgQCXZJcxOLOIVy3hevQf3oWjLAcAUlwAm7g6Tk+okf/WTpYxqCki
2fbR/WiTMxj236MnmX3sjCv7CC6W3XU8vF+vCIANv1woTZzBfpJC0DMLEoEgWD+h
nvu50UESscqonpc1bg+e1aOYqv8wm/vJuowGh1MOkuup5soGLI6HkH9p5LqQ9UZW
1AbFIlQ3yzuY0wVwBjWBPVzlJf5x+wshYRykfILAT4rLY1rMqgrRataox5Yyci8V
31Hc82r/un7BgDoVaemmdT+xod8hV+Ue6nERZvXg0iW8EhcXsnjW9rWQ+MtPTTIi
wjtMt+CwHIvQCv8gYCqo7PVvtBNgGAymfcGWENWsuX6Gf24crF3QGq5+YfJR4pE3
EjFvKu/e+FWa4qOEqZeGkFTyGiKTi2PQVI13oOvtOa8HZwuaosBQZTwPFTB/r80S
J/JGl2miJbnGpwVp4XojrIo7GQAfUWRpkG1aDOzUsd6bItKc6bFTbiCkTRvKjZa5
TnGju0AbGuQ7Dy2AjKDF54s6cgi1PdLjpQhrMM0V5joe8BespCMOLXB4bv53Xni5
LUKApttlv7T2si6p/A7dBIltLoUOyxrwrhMwfmkWLXqvueJ1aj7RQih+tW9TbO4m
oCPxCUDHCyfm9dt0CRHTynUdMIZzQrI921Mrg4XhwWv/0irtfwgbKJo+M1q1x7sl
sMStyGrnyJfy5L/b/tgCh+RupNtumRbrrwiOk72xbg0SCI8hCbottGzGRpGQpGmN
eA29oV9x2cHLpRWTIm8Ggng/XoOfId2rHuP13fje+4f5QWhzjmWN4E9akP4X8/9C
JuKMMghJw7VY4aXwHRozY9VKluF2JiTf63ifHCf3gPwfNHm1oqpzz007R4IT7e93
YIkcfnOg9jzOcRCzu+KuouopSa8ilgGiHaqHX40XIDv46Cum8KAITa92XHgyTH44
jDqye8E8hh4Z0SjeD0iey8ukmBNvqbOJOatpmsuGlJ7kVleWRrr+5H4wbimm+UVx
TdDEdkbu/jkBHXhYQ1FbnVdCxvrpomqlL3wh2OqdiPU8kHy/+7gl3ySzQWKQZ1lY
UZdMmVicB8SwQVwQwCryQg1e5JE5mOR6i5GHbOSt83ih32NlAv2IoUuiPl2dlhUE
lJ3I4jYS33+pqgqfNwaRsE5AT0tGLCFvNfCk6PiwppIrhtKYPHw0Sn1/QmcSIHjQ
HSe0c/Bzn8E7nAnTaVofafkK3SBsRVnQHqJvOsIB3FJBtFIzwIQKtmJMbPg7gpT3
p4PLW+ZySKxKW2dRxDxlVvrEbdpIf6iIAGg9nH5tyGcJwdgVtYq+FxZ9gAusnSMg
h4Ximh44M/PEBlqo2+m7DkKtFMB5P9/TnQXkKSiSW7pSD+txaL6pvo2VGl6NfBbn
oKQ+lOyEKZiU5Qz9wVRSHmGHYqkwcSAH7/919FTvoxalOpZsZMaEyvmP0wv/YkfU
ej3YT1IHbkVLEZ+rquxlsFUPzeq5F8UIv2uhYvVwjAZV1lYfvGEeuILyUwb9APhx
f4hJdUhswWR9uk3whq8Mkfg5ssQgr2ngphH0IkBW793KWDLN31cQkVsP8NAiRbE0
+ah0f4ErdBlMWyr47VTU/Qft1V1wjEBknlAWilHhGwbNUgwhhYGH2bzs8KSYlaFO
WmRf9qsEwYGRH1lowLb1WFOOuuGxABXnfaqJmpsNnMkUeErfxMK606OdKgWJwTiX
4tXBc43FBJ8gvdeqHTY9RO4p2KrdXEXihadaVZLHP7txd9OnboJUpX6eF5hpvoet
QF60a1sZU8ivcRtdDfrob2DnUOyoYMCiNfmC0ONxpPA4rE7hkYWFPkokD8HGkH5z
xF63ZBnFO5jiKLNfFM6KnNP698FOghrqvcUIZEKtvcbziiirVGv3jhnDxt65yXki
yfZN+R7JAvwuc1rV8jk+Kr48WrBMoAeRvuCkNwgAKdgRx/NF76OswLCYpfu051KQ
hjvSxfZjuMg2aQwiDotlmP/8XrgiFp2S+JD3Th9/RtNxC11HQSd57IWvEUqoCXu9
jvZ4ehxKYkwaLH9EAmRBVX2dopnNJiwGP9KsZwrVVynooLNDVgwo7jitZaak3hc7
+Me1fT12Er8bjBFZXQTYl7JgzdqY5G34BTOfNSh7tx+USfJ8Cq7Pj0eJnVJzrQ0v
YK78gmgoBZRl63NAM25VVnTBoGhv5RzRzM5gSZ2winWnlZsdI+IKBsy42fnMir2t
eHP5EhI1XBNccNY2eq3ECdnjOQ9tnESUjblxXSkgAJr2aWmVbLbr+uszGru9T6vM
fmhuawwcdTgD7/RxLyWrw5Naa7JMQUpBvABt5+ZgLxhoQQzknlbqlmO36i55lEi6
tph14SJACzp1KXKZ7cw6iT+QxrBvq/7lTFsUp0EjD828GDCm/qmc3Rv1TWbmVKfN
brS4eGsRlg+/Ds6OXq78oZZkCvsnM5hQRPQlR2zG1bGpcBL1VwX42AV1UEIlODA0
WwXGZroZ443Hyh/cUiWlM+NGGYF2ze99Jo5ZvYFwS5tpDG0DiM6y9LswKnEQITN2
mzxLDjTTI0pnf4Auxw6Zbynl3xcbOUc0j89nA5n5/W93JuvhpkjK7oq/Hv5eEPhd
tA87lwPlZopDtKMXNZhG9iyRRHwzMWkZki9Bs1XfLRVNASTOKBtfJrTYo4sydPL7
XqFZrXSpm4kov+gLwhpKBh89MIy3BzFIbxNc1O3WMqTGnIene+MxBfWjhdcbRZDe
Vf9n+qYS5wKsNa49FcBpRcrAnmLwrHEPGoknAtiAwaDJhkOOY19Hc2WmCL/P0bsC
Rf+1CrDGqzcvN9UmE4GtiSEnscPV6NhBLRjBcRBrBz4Qpvph4KfZyeLIh0DceRo2
/JTUAfMOagYIRrb+j4LyqWvUe0Zsy3xw6BMlBEhgo2NiACfj5PjSA9IEUMF7xNgS
VEFnRb8dJ1wfQ1wjRhG71dxwrTvNALj6VOAW6UOYgfvMrn3UPEJl6MReeQj3hAGu
HehiMl3hYQTV8d+XD4r56aiO3dZ7dOAJxE+NiIoq4GdpBsZAB8f+wEbiSATyspwX
SUb2POmDEnKVGZcmucsmEA7A9CuENAlLKh5xZdKxiwrcCO2QGhtSWuOA3haP5hoT
zj+t1zeqw5ECafqnz+GjDQ/8t03vQY5bHBcTgxohQnm1uinI6yTPLa2o6yahPdTR
0yF+gBeJlkzm3c02Yc9D15rj2iLSHoeb8xaoIw5KrC053VOLLqNtle9ugsgsb0lk
vynjzdww8MBmbJgiQviDF/Eq8kbgv9uyfjF4rZZAn+KKaVxM7q7aZ6Lj1ZqbOjk4
fc4j3fdIHiOVgGkez3d38FQtEw0NFbcQEYgt9eioHn9p7deT+WL4GFq9joAvgiaQ
fhyHGUXeIuEaSmNeRworF/E9oaqLybnIOgHhBNVdwSOHG08vuZSb7EHlSyrFSmVF
jCyXH5SDAoX74+/C5M4UCMikPrADWdHyvLLCXn86vM/UWi6HhRDoqzXNa83XjxaY
grVVY1VyxkaQAtxk472AbdsHMfo7CNka39GHSU752TaTeGgjUfbklbW4yKQJOOe8
0Qw6PTBSVEhxAWsgKzlz/9cZ1GbLKd2/f9L33SNWAuQY3O0+N0yjY8bLjStwBknI
dQKhi8PsiwW8K4nW+/294aE0fkztt2P3PDkBUkUoMd0iZT+b366LG4hdRBxlrRzl
T+iUxMhExaK1Vjp1xMHlEHedUhxhQQX1P9A5VgYZ51ev2DmCVanQgIfQwzrzSWur
owTM6hi8o2P5W1RzQCxjAyM+x/xFatZSuvy3JLu2Cf3eepjjKpJaRZbBRm6OdP2m
HeY367k60JP83RDvSIilIB8b7zIzByTm29zpyyBKXGcljtabG3nB7Ibo6k0PRu/k
lMAWJw3jhHIUgqHa8xTRHjgjwy1QSoDtrBrL4u2mYewFYVOiLUUqCVX6x3zCVXWg
66yfj6AenXSS9+/6jH4zO6NQLzoecx+4xzVehbIpeIvCwPp/wrfHJF1JHNIIiZbM
tQ6n5SO/zis31pfZO2pG3IZ/d7NlivzHCCLvguN318tLRRqFgttrQ9fOP5MUXgF3
TQA6go3id/WOSnJZHA3DYTYIelVA3RxTVbaZE7c4xa1nMWM0gcX3mwxHZqCR15xk
nR5wB/qoKuon08CyHm6oA3IttC+RjMZgCG63saOtcvwW3iVqxgI5IYScTD7cJj+f
xm849b6Z1znENXocp6c3pn21N/C2f+fzkNBvu7y28ssfCiK93+Rucn2ckNZcBm43
yfkmwBmiqMDkUIRL+YAIUk/EwvYXSLI81Nkh1+493UlOPTde5Ct04G/YZFXWoBGK
8kpdQ2x4B7H97LtL5w/M0f+55NbMoQN900rBjkGcnuPtllP3xPJeFuC2Ww0YDCKM
xDn5fKM9IHIFCCic8YVQzRXicNMJb3c+xasA+lksJDXK7tcJBQYsg8bFCzar90Qr
ngs6vm0NcXTgaQYHuU8vmQkqozkgZ6Iotuwcz+6n7Z4xOkgRE1j7ZFaIR+V1r8VJ
Uso0mazBNDnVE2FdAt44/yUVPF6IT20WnXB9xsJrn2hmjq6jD0dr+yj7CAQTRnVE
k+a/ObShewgBBoJRkKezxyiRVvBvyyo6zycEAQPEJ/J6+LwAK398P30WiGLOI5dA
gMPnzXlXe1HWBeu8sWPaplMRq9hOsH4BgIJQDR0lc/FEbFktHkhE2kCqneEX6rCn
hcnfL8s9kPqxl+Q966wSxwAglgIAsO9rgClbuRsuaMc94w5zFQ2S0nwAEO2y2inP
TxMy8z2hCk7Hg+neAKrZ0khR43wkjTwev8YxjX0dNlqGVAr7mIe2kVefeHIymiJ+
x5hefCdxtfVBeLdKCaoGAf0Gaj8Ka2NFQKIwG/SAWMIOMWd5SSh/jF/hAsJ5B4Fy
ljdaCpi/DaZZVPzvWUzorO4dKbPxSMnTwTcqRBO6ipU2HZ7TLbvq1siZFueR1vAW
h16T85ksSbZv63tyhH/U0c0xZgNLbta9R5EzHv9/JBDOdonl9tzZGBBhFQ+QdI+2
w+njUWsfia0RGsGw/436beivVBPJ1xnPBN32bDKdkfD256uApr8ucIOks/ak17iU
xJviDn98tbWbYpld87arv7UPhmT4z3SOJ0mtZLEK+JQJXvw0tecglC7XqdvscjIZ
7+7Rn6AroBBkpetG6+7GiQS20MgWN+Nc0FUUGBssWoP2WWWkAjoR27j0qBgeT0RS
zoOcRk6362kkwbHTuT4pDjYpkW5R/CAMfmLF31iaF7ckV2cBJD1Ty+NST7Z+xjPX
/MjEHbslKbe0xwGZAggLmEjSU9mRgtNgDwxOiJl9ksvINp7FWpXBUd+4qRRDh0SF
S8paydaqwwmhsRgpSoqr+UiXn+QWUiOFt0dh3hrAyFU4Rq9FONmljKF9gat15X2d
z5F/c0oO48H+UvgXJcgP9hZKPzgQChR2revpQvNOqWn5CrdYI4jC9vTwZsxuXlgl
EWQyyOmd6tAobVGQWPV569lVmn4UYxoVfZK/HNoxvJWtFIdhwsj8p56ze4z6whaA
i3TO5+D0a+Lw+0o46Ggyk5sEwQci0eagG0jRFk48Tmt7f0tqOMuntqU68b3v+TYg
XwQyKaobDbotNuaBDbcPnvjwXLkQEl/oI0b9RY22s9/phTpaaEvz9igLm2XUzSXW
H8wFFCYUjhuv4f2VSPLhaoqEsAEnFQwzZI0qJ7y5y7woJQSocrTfK9uRGM8TA6MQ
yX+vyuNOt/zZ3wwQkjqZaeAiOVjt5P0KwuMDCKkNF2vLKqwk5nm6mjgMpcR085Rv
rIVi0u92xt8dnOhog51R0tenyt2v3F2Yl7HPwiesmyusCl+neZ8h/xlpc2yBf0SU
DEpXFpm2w1l7n7NvbSlqdp/wg89jJp+a7CESarJoFztPqK+RGRzZwkxRQiWp1sNs
XDK6HQNYNJKcu1RfjcCvcclLnlua5W52BiawzpN4BWg+VItOc+VD9mr1nqXMPURM
9c1z/tIyFJBLL1/D+YeCrXaNiXBDX5hUxVc4e//6g/1NZFaj6vqLMgOZ6EKErkkI
9O427bGos/+UDSuuD51MuoMYwd9V/rosmvtprLsCvw/RFjfefk6dEtcGdvn0uFU7
fHlUcPqzjtZ0q4YZiq8Z0FgtNJtJgwe4W5khKTYZnNq/XZjkdZXPUq5cBSFKsl66
MajedgdVTr7NSJL/N5JLrahiOY5NWfHvepgE/Tg1EisjIVlFcstH6vsfFy2XUnZL
9yxivlJuA1xx9iD+L3e8wIV84sdoTwT6J9WuidfCgx8oX5MRH30sdRKm6GP2HqVm
ZmpuMhKBsgsy1MfT1IE51DdAIayuuhCEfeNMcAfSPp2izqq2isJLT7UGbIka1hg8
1vqlO+5Z9G43cYqW5OLClDofN2HQ4I3x3Ck0nUJ6X1MP78BNbL7Ne6kcx7dQI4Rs
bbdKUxNChIr+FWuRxPBkFBEx0Ia/+WJNPpQiaXgT9fOOdNJjtcUU+4YGF6f+CPOu
+ZRy0Fbxrbpf/fE88JJ5unjkqfqxwEAFPrVVnjP9SSH7iSqsa7bBNuAQZ61sIk0x
fcHjtf6a8HjSYrdJmH3o8H7a8W0DgBu6EYBSeR+AZFInmtGN7qEdNzF7RrWr4NiC
Cv7srnTMevNVhLpxs0azN6EpYl8XIPxGnCYsrluIwpJP+3QvT//ckXs1TGByQ3AX
7vWn+J+3lASefe0l2V/UERnKJd4HmH5Nc6HTtE2BbXgzYRYFvwv/DYk9uKYZWsUr
HIZ9fzx+NMX2ReEr1hEilOWuQnpJXwq2MxD48e5RtROai0N3Uj73qznQPEMWuhU5
BGDnLLio8dqanSMH51MaTpqh4obcPVJuvh53EHx6HH3wemOBd4ryRqj6Edoe41sw
k5u2NZYhCnvEvZG5LSWlSq8zMVaWOyF6BYvTzuhVtkVIc062zJAo6cDF748hZ6o+
sVVTFIoC32RE+F1lSiGm7figk28fzNdHy25i34ngseT8M+irToKCWvb8vk8r14OY
KwIU/xbxClrm/LFXdARBXRWcUspFmVxC+pnlRLZrXjFgIxvFcrSdG0Cj/vlBGd8b
l0V97mOWvbprZerHlflIXt68IXvU1i+/tQoSukQtzvaMSjoKUmcE7Bvn2QGs+0Th
IiEgAD2c7S7wI91MQCh3F8LLp7s3uZPV8pk5Jx3pyTsuBdGTZtD8lTpA9FBsl/P0
7ECBHE+ZJyn3VF6eJvax1d1QIIwaK69+BB5XE90tErT0noWgbA1mm8O8U4MhKDEP
6q7fpRzgOzCgoSLSwt9SQhjl0HQmFtt00pb3b+yGNDYJ0UWg1vsbGj23dlotGxrg
7cpbcqc9S8uQkL/AESD70R1WYgcpQiVCfBMVkcW02dGffgdpeI/mT1GOukJBbJLP
3zGOIgkd5Z0UWyktB3cBAi9AcOW2EP6Wg3s36js07Q2BgfK34E3NUZV0K8qfjDLZ
WJACRBO2S016CuZ4Q8t9x35iH77PyJ4JvbOeeSBU9lhOxhoC9nEKM1D3F51cS824
ix/Pa94JJLRdRYj4EFppzm0IBi3lHHzyznRbfbAGrsoP/B2CxK4YsEz/F9grakg3
LEVpfcS4ohlal9/kW22ZbVDgeDFw+MBlFDli42wABonPopfXvIk4BKrCKy1RWa01
1IIEXUOuOgeEYrahsRfp54B2mJZTQ4SdftLW3wtSg6iP25oj55g7kaBW0x2qmWqJ
+OrOmHMAHaiCabkehwreMsQY7dHb0eju2vZtqsrYGJJo+P9EHP0GVQU7z3IHpeNX
0t4pCZ4UemTAZXPYwU+1nvuuNc4QGNOHzM32cV+WzMrJVH8jePxzQwq0HRAj2und
ZxyMw9s2D2qMCF7EA59ab9erBJqXNfOpUTtp40qNT7GKUbYcAF00jLftue3cTD+Z
2GTEtbAIC6OHxLV/+WrKd24gj/as+ZLm/Gdgm8rX0Fee+Y5U2Dxo/z0bE7ULzVp8
Gymv2tk2JY9YEiUQae0hKR64aqHddgb+X/fst7u0PmZm2qhE6OvZeA3Y5z/CJXmH
2gvswrHW7IXeooV9u0HBb1/LIFIfPJIdqltNed40e9xJPh3ZldHK9HMo5nisncnK
uGRvTQN2tfLCH5B7QNiX86EFG4ShoDqaDjGudJG3G+/6H5A2GSTsntXWB/q5Br7l
VBiB6XvsCB2RTxyW8XsRfWieHS+qLTFgOpAlRKo2OLZfExR96IltS180VIaliXfs
xVVE2CFL7BYP9QnzoQkQ2W1D1YXUXzP4uGf/zBf4BLnjtBi5LeoeNaPUiI7qcK+6
b9krec5nY29n4SLa0ao4dG+/JQfluJrxlVUJNZ4LtFY+6zAljCxrQXko/AkoJQWQ
Ds8HfNamk2hGrk7JxN9wcX/Oq8/S6iXOlWFvma0WBvRsNbhWhTFGFU2m9p77pyuf
uq7HcldJkqnZgjguDQI6/i6M/lUtZUvFcXu8Ir7TWH9UY48mBMGSOfJ2yFocPI+Y
LAZO82snQkxOzVKGe3cfoyL+K5wKPN7HwunbM1R7DrX19bxnu37EBXNFCX6Ded19
14PsXyqMgTplONHkHLHTMOpqHKqDawtO9+mmamhIwhI3VTsVxsrdgSNyKSdT94+c
Bs1JnIWzRqUJynbpKD/PH6cbKZo+4R1Q7N3lvVajwacIDOlTkqnguGWvArNnjjJK
Fu4bytDNFTdASs7ZpU6maBRVE1nVFIUFuP9rZ4rppN6IjFcaCRt5CDztt0/ftXTL
DBeUsY1522Atfaxgvz/mHLEaV56P5bCrOB/26x3mQ3Lnat/ypwlygdcEtRzN3H0e
a6XXeb1kNwM7Vb6UlSUH9J8UeQUhug+nz2AT1NUTylFOjQOp14NjNKbabDilF/1A
cCyK5PlNhiSNGOC4yJ6HxSJ2oNuXadLLgv3uH3TC/xWedkBlUgnvK9B9dzPixEQf
qlhrVaw32s194hKNAQJcUViF0KY0QxE2C90JlvHO0DfaMOQtNH9Tr76l3cPBCFys
ECqqWNNE2EZtqicgtTv8GIblhlxdsIIkNvyY7AQ57u0sOh2ayoBVBO0x+b+p1dYN
VQed0OTkr4Nchzvk4L56ikIpOLmP3MJADOWLKTaw1HISeo7axotJKV+agWRJp0Km
omWpKUlIEkBhv+sW+SLITMeWmf16+5nyaEK0sBEqWmAVqhR7pyOD4hA6tk2tGeat
0OrdrZEB+b8tNp7b/uVeCDL4QeB0RylM4OJxI4jT2p18rx6ktsR5gGhiVUnjftp6
+XGCWMLjQbVspQiQeb6Oj5Bpc4yfQ12iNycu4JTOdirOOQwXyHfShv2iHt+eWGyy
AiDaxaj6drDxiVqr6LB1uD/KPp2A8xgvXmy4iLVNRCGlulyWrS1fymTMu97+7TRC
6PQjKKIlkD8HDktUk1+XJPMYdTbXm7koQKQGl+wMKMWPMFc6ho419o1m5yhbigym
ZDfdctivlbk//ta4QOOVJ5+PGKvC9vw24yTLqH4hs9joG5Qi2qmyah3I7ek4czrl
uqGbUczGWJWxEGKSaNU60CnArYZx3um4zfXRfmP63VPLS38vSgjUXHLj8TOAchbR
6IaRvKjjCrPfws1rUfCDmLhd286WPjqq88D2PmJJm/BsBtC92wap0wRN6VvIsOzW
mlynmqodRNboMMyjOwbNm37ytxjn3rOVallE2I/+ZyPh/CxkvodSD1aJ/s8muUkk
EQdVWV6tg8qRINX7gGdTSDQwx0jdErXK7idTLwBEXU42wA8s04cXTQJSWLSlz5dE
Ia1PgfepBMYlu3Cuv1N88h31hSgXgJOUxs3JN53/e70O7Iku+Y9J6fH5kNBNlZ3P
NkHTP3JEsH68lhJSQSVMSbdg3uU/gWaBPr/6/cdDxg7FZpbcIOa8e0QPDfjHwMiy
xe3WLNV5g1DxleTVtmUp1bc/fHXTlHtnnlWYRrz9T9qxkad53RCNNorIr++jBXQ5
RgypXfOLaDzxoaiduorz2wTI85bY5Zqi5sX5I67VMfSEUFQotSfpf3/I/qS0yGHz
BgcDIcsVXssbEYKCEoQWJ9ck63ZhqKtT6lzY5Y9hkTEYrsLuVnQJNMMloGHvMDnp
f6Ok+Xkpvm8xmkPVNwdseiguwRmH+lCnnlnhI3qGkk3InxlYg7lBygWPQo2By9RW
oLyR+YtmVfR7q/KRsRQMUHNNpQk7shAmHYsCD83WHOce5mbGZFaZMRbQWbnvhrFM
qOuMkCnkCtIs/l3yKYCdkIK6NfCz3OI35Pt6SbqgS1bxmBMp0cXUQAGwLbchkBrh
uhvD26Q7R3Bv4CnCFSW+KnIZ642GSfxIlU1S4PsJYLm6J2eSPuvp8Sc7Gk/at5sY
AlEubQPTinsY1Xde7maDFKmujv5x/LSgBCdTL9VlfnUTAq2sVkwPu/1w8LqsT3sv
8D0wR5/tTtsdALre2GkiqWEwtAdK1hhsW/izSxI8xaZxNeWx5uWzVHIuWF0PnR7A
jneCFN2DlE1aQ31AIn0pMQS4ViJdQZUbd1QgphehSWXFyOtRzQJGU74fg7v4Fs6G
Mt7vWC9pPKY6gySsBSyqJSBbP79YhlY/HD9BwspCrFHXeTNpLvqRFoSMXxO43HPS
HTW/3oAQ12OfA7YzCplwcJMBaWdbG9wgiT7tYtiQLZmm71RAxa+Tiz0jZRKgRbhu
IxDHLpuBBKU19K3PYOqIL2KANpACnuRiqH+W6fLCeAyQ6BxnhizjpG7RJfyg2to1
WIcHAL1no+cHP0B0JKpst3yTr+oaqm7gQ0bl09w1yBGnlH3LRCqvK39pcaEVUDTv
i7Q3Dt+VNL5Qwhw7PYRPOPpww1Q/0cgQIDpTnpqVIuovMlLAH5x+xV1/kgnYhiqb
dx460WiiZBgR3SWb0OAjWB/ps38Zrbn6E1XCDTlEfbnTIX7T/0G9Z1BQ6kKVLQ3P
Vs/t/dlpgc9QUJsTXZWtoJZNClp3k5hqiYE5CT99e42v25pJbcDpB+lG0xQEMzsc
SGj+EfAll+hXgDTjC0OAm95G8/9V/Y8M1bLivqTpmgPSzcjUYPLdvRm0KBNOhFGQ
MXw5YQWe5BILM23guNu3dpaF2F/aEgxUCToa1qMzSrIFW46DNUN4FoYFEZD5T07g
kMTR5yP+ltPWADl28dkRpDY7b1RUi0fO+dBXOAhiYeh+TfqS/4AHkob5Dopym8A7
BK4squ1GjCmuiJaZsYS8MaOl9WncTXAkBMYc8xF720njPPLbx1ftvCyqlHvfO6Xj
CPP4MO5mkPB7b0xHOI9k39qOjnQM8f9xADvfv3KNio2xDdijWi3WIVT2SIy6FkMy
aZy9gANiWWWnDZ+mL+j51rLyFGJq8hn7fxL+waTGbF3/3A+91hTm1k3ZBqiBczq1
Q3kORK0kch5Gro/JyzjFVi0h49DScwjBEjFcvQ9Jg4GIqljlZKJXopWU7kzl5BEM
g6WfcNBtPP9/dW+gn380UYCuFAVURedYhacF9I9Ojx2ov8oe+JeOm+wTrbMEUmxP
C+nKuK+pMEO0Rl/47EIJzrffKOiRCnPiR3xD8zjIN7+yTZneQOadnKdEr4Sm4hkn
gnIU8y72eQ2AnMzpmPY0mjP2l+U5AYirI60oeuidvFew2lUROAt4kO0nzKneqJvB
XsSQAwffRl1qvYrskbowJ5eBMSX+0vIpESspLDyZwQ7OtU/VyuzcPqkVb8b7BhKE
wMqpdFLd6G2OQi+bFupr9RZ6NcYD7NvzkL9z7RW+q3bV859c8Q0FVv4dh8zKLdYJ
qmftgbnTW/VTgpNqjq1e5JnGKfmwvZOM8KOxjftboQAsCXZ7ecxMbO2qTYwv2rwU
zrYlRz5d8jfvI55B+YtgHUu4XX3QxiFPyDvzWR1LCrFM+bhB1IVu7cbPIQtwUT3O
Ge+m5Jvv30qEOpB6lhL07frBdOxlwfCygpL/pMcohpR5CfLYQWqp5XoLjfRXaqIo
MyETDjd8a6w5zBZA6EWBe6SusjTwPbne7f/iPzYMV/ZJCTxAmCov2Oqwpn2g6w0+
WcAqNFvGQuNM6XLlDWYOe+ELj5n+A3VmNq1tfeTdzg2P+MDcDTZdKSEDbp/Tyx9p
/jT62/S/7Cw3WhXqa327ABwMA63rlXDzOFRKlpopDzIJkmJ8a2OHM0mJPyGb9eL+
KaUEw4P3FSNfbWIz/cdqMTrRu7GlcN8728SPHV2IJW5JpubQo0QstkfjBQ9gwiy5
D9cudgfdItihuySVxqrA8KSs9FNb4xqmTVaLUDbmpJCENs77wpdxpcV4War70B2v
ifilrCfaQJzQ1u356c2+iSzYa9UdfTQsEYcvk9hDJyw0kFB1g3yWnbo7S2jH/9gu
jqkaX3tpZ1+t3DXsHSY/hx7rkznTna9ni34B6twR0U9mIjIglSnvZ63yu3JU84hW
T0aXl86TT97msB/2ldyGKO0TXJVtU67sQtfZKSHwlgeiSIyh/IKqkK4FC5Xaxy5c
5hP8gM0KU997uZ6d8mlcmeZfG+Y3S8/mU/NV2ECnqbEC/79k0A/7zb2RPwQAAkNa
S3fXi82UoyP+dTdB+rbF11DNBIWFta1Iemtu1qk1VWbYjw7JLBNikkXQMHc3Dct2
I2NG+R+qRwpdoXKGTAgBDOFtFSe5lJ2WhzWM77tumH/KyNC0nbVNewm0OHUMJ0JI
Tda77YqrZmwFmBQEJHoP+juFcExcEqdWsldWN0av2UPJnG+V5jA1A8Z9cJRD4dcC
sf354pxla65kdsDskGSP9VM4hQc1pKEjUAXbF/G6eRGxF7bNFJvr+EHmKWq7h35Q
3iqDpFDlVv2NOJ6VrvFQkSTxZDSDkNJL9sKd2P6kPLL0TsghcWDDTQUqaSoh5c6I
P+2m3NL9r66qhHSJnCzoDeSOimzGzAapErPN2yVcNPhVBgbAykkmKv5mg2W5WaYR
T+i3wUGVMDvqDdWDa0v33FFPQRqvxdbUfuUp88BAHestAOIJSoisVClVlJ6LmaYm
i8KO3t45Kq+2kHLV+7Mrc7hkaFJGs/yoyjY9cyzMHYKqc3lAtvzY8kMarwYYPh8m
YV/y/mh+Nc3VSg89a4ryYzXjbkCRdWZgggBYl1SBoDKifLgwgfQ9HRUBo5av1pRU
a0vkcCzvLBMSILu/Zo8kwsvfEWmgAuTKH/DdVC51vF7hohgblcGe8A2wy9fevN30
gnjiU5sjHcfiDc28S+Tc/DZ5gWc9LcGHH5Q2H2ecsXVKFlF2pPvak4umkl+cTDgd
1re1uCkua07Nb/iZw6iolCqxuLfep6Ibfr7ALSrbS/26g3Pp793gC4PI3rYE6/ep
ZPmwuVI/kGLRtMfaHi8ENtUizWdRJaO2CQukYXcJWQ+7N4YkaWAEjiC8cjNiL0IU
CYD6gxrU/KjV/2T1m0eeHS2gZ3Q0YU7He2bQSfZltWPxY3BGW5BBbm2TirDp6Kws
/l+a+52JIA2zdER21Cy25kw8OBA137nTekhQ8VCLjgq7RtOW05BLiwf7LjlCKa+O
YpPT387fQcuVB7HplBe0KP2xUAhQdghTmWT7UH8RDceqNYA2rI6nRF2+uFSFej8t
+/8TZULJBiNodjD0fHrnRkVogBNmoLiR7dZXXZsc3rUcImqS0454k80Gm8YKv5t/
yy3k8pSSQl9f7RZ7jv0AqCBMu8pUaMvfkNkHokeMG05XV86wpX3tinb7XA20GpWM
g7hOAos/48UaRSnRxYWTcu6166cmGNxUFY6cU2UvHXtIke/f0Xt4hwnezld8rrTi
YkaSgaR7N62kVlrmgxbRfjcZzu2yc/1aBligye/duYHxl097jrd2DZpu4vYzX6/M
d+1H/DnuTnhQnR5gjdetnNg0xAYkiSCK7np9nh2voxeU4G9d9ntQ+V+FqXjJ0hTk
8Ejtwi0sFWK+HMusHR88bl/1G6icOgzbc2W8JtbRmsxuSLF0K1tkj7IwcEnfsgJE
mDi0tIaixJtM6x9x79DCB8hRwwmoW5bw5rGK4X/n31CrltN7FWpm6T8a0+9XICFT
PkI1W7H8b5v0dCPlgKslPz+6lxFsZsHZRp/mJfvvuM0MDutC8UswvUeZPIlPq403
cUCXCfPTyHSbtfKleZ9w6ZVjKm6JYsSp5k4TbGg7A+8Mxla/Vvz5gbIK81RiJ14e
JnO5mEOGHTUWaJbvNcMgubBGFf59jJTHTYgqjxVs+dN5vUzSsaTx4SnGRFrDQoDs
uad5XHESUf5j9nCeqhAEdv45XgaTcxawEpTmWsTECzH1Ap9TVCYK1iEOlExLcx9C
mrt5lgsTrIrrQOuKlRrdBgNO5uLOkYBWgFeH5QklxWozWEyVHaU2MzZPVcOhSB8E
do++mInhFjdW+Y/kk2/x769/TZ0lqJ2GQ+GgRHoO4W0ouDRv6NXLWBBQppc10zpU
rBZXJ6yE2S4pARv99+bTyKNhQHnfjhVsm2BzEhlnkZppyyfSk4PEm6dUK5kPD9Sj
adhN6YhT87/ltkHHbdwpqGQWljoVWhFXCeRnVjtaLhgasKP9pcB0zVmwi9xT8M03
NchXEMX14aw9tPNBrFCKfwk8vcq6gbdoFgZsRI/Z7loyXVZXzAZBlVMMRW1AsWqk
IeJJwhU4MDhtRHlDfMRhrqM74n6V6ZBu6PqssfoDTlZ1ZAk/IUKq6tRXUPHt227B
6o7gSa9rjkU3cco4D3BJrAmK6OfAxkMCmAvNq6/Dd0OxvxMyCUl6bTW27WRe6tFs
X+1OtFOlBiJ/SnccdMs2x75ZMp95xvqIOaIL9KuUmRWAkQOzUqHn5LTH4qo0lmZB
puefnlAuSDXkIdNT1obfAQJGgWxmyYQLOQmQ7zoiUVCn7WfXbEJy6byd2k6yRsh2
iYbk+4Aa3KBegYQq9CVwD6I5OoZtzjVnNXBIbZfszAZjvLz0LcjVJKJYZ6KuRfan
UbD8ILQE8VhHp26LKOX7X4ZZmJh404fuZCAt6N+U83H/tWPZQoFG4JxZhbruqlln
WL2v7J1scFI5kZUIWzZGoATmulP2tFy5ST5nL0f1WZV/+BJvA+iugykKP+9ZdeCQ
ye3WnT98sA2G5XmZeUzZELe8b32UcSZeJqenXs75bs9uWqUObWATHP2CJq5uAO5c
9/5EWaIVn4b1lR7Qm6jGtexOo5pV78cq9Lp7m357bmQWYsf+bP2X/it49lqgwPBz
A4EpNDVBSwNN0In42ECagFwZLidKvqbEwVlivG6sry0qPT30UhCXQswX3oLrL1nU
FA5uLwIzcJi5GH4aaOo00zJpayBFzYq6UFPi14K6RF9Mxw0gBL6JDnxktNE6vntv
bchg8UsF/yH0g5WLUf27mQERBfclqOfuinSKKepjVnBhnNe1+EL8iAIHawvlyDRo
lcxuVvgTFE92NH+VBd4oQd9YtS7Xg91s5EfTXkE3gzI8wU09Icl3zy8141NQwe1P
UWM+3lX4hH5jbet8UqVVTgdHENX2xWs/9QfozrtUQi7fW7UW4er2xnB+9nMhi97+
T2X2ppYQkt2EaIf0CnnFyAxCSzdfGsHfjD1SdSsp+ZwploNIBSrnKZemVsi2s56J
bBle2RQuTGYtdrr597rA9A5TN8C2wlPkGnsrFtS07s7vfOVmfCICS+ftiFFfwSj0
XU6QZ/VwBMHgLlQvMq69ZH59p4IHt6KJtKrzLRb85DunbwlmSfM+WIKbBKbH30rt
TLe76rlYifCPlReRPTF34dXUx0tTKfAbXjubgj3gtMJG75EvWsemZaTenG7plOtL
tyeA4wgWAHb29F2r6TfUIKQtKjsT0gkDIpdlYDS/ICRX2W7z1Ie+yQ7e3vmLy3AO
80wCgOj/3C85/zP8ER7V696BLEszjQyRpiqIUUCk748MGywK7r5+mWVDgCtVJScz
gQyKxnkfhnjRppw4YZW2zKDfgKLcQLa1ITarSP/OwC1Q41zLAvSP0VYTKM0vRD7s
SsUInWHE0vnXMSB4k6QDRVBXDxW4WnvK2FP0I6RxgHQKxogqnKdijI+/AqgvDUQG
Q9LSJya/yg/OqOdzFW59ATO/YZne5gM5CPTmNHhghp5ATgpPej5qqgax5MwmAv2s
CYN+V9Mw80+R/uJVhJNW/wMQQIq9eP1rhGcTGPC0ND2r0iYhbnDHEvlt4C2LkNhI
aA28DxPWn36VRsSLO23Mpf9iKxh0i0Uh99OrZZXXIJuTgL62QQV4mzWxf1Xp4raT
huPJUTxJFTW7mRXzi7Ps4XLdHio2gekPnapv78hGRvuXlrugzi8rQeSqMlPrd2A5
Mr4jKGDfZ8WjiiVg0Mm2upuDwT5PRMSdnM5QTmggJQdy1WZ2RGB9M7/FWsVtB3fN
my34tGjiIHNKz956AvYx8i0JyILCVea5wOclEkB/eBXnrtMAA2jQTPmiIEQUbYca
0QHA2gmQbbrq1OSK8pACuhmD1U/abACmGHp6LRm0XouLBDoVAEi4LkSGHWHqgQFU
DPdR5UD+OYTY++Y+A5jw1D3q6UALqxZTFHaWYtUw0vfIHzgPKw3mKh15DpJYYmIj
Z+X9ySc8yGzjweKCMtYd3cnEj+J1smC/4R3/53zs2UtrCcNUwVkG2bDVH5RcmzVe
q+8fq06IBsxXfFvVFKKGMFEMdmBnJfDUwe797uYU7dPvPmi9bSdviUYOHBWJdB7O
KdxPPZ4i1fV7yoOcum3lbP5Kbh/r80iRUd/77csUeblBMmJsa0xAWRAYuhLcabID
wVyvYxjZ69Z9N+vZ7A1MyiZGL6Ci4r/ukenqUSb+dW3A42qhpULG6YRiibXE4RyD
LQKD/vcHbgzXdg0yhcp0L6dqjdWnCmfLNjdqSePFumoezedquePnHeNJ1yErllHg
ndOTKkzE9BFLc0hOGINdcbNsyZlXlmAG3RpCUlxnQg0fh266BS+tZbksAOjV2nqw
M3qoo0NDsSSsUUjFQeeAw8RpQFoBduPRCvxcyf9MNxFWPqB05hZGGVwp22RGo5Jt
l+5KB8g6MMPUmf3/ExgsMHZMsMxYn7joKnpOUClZIOGAhrWrw9eBqs7JungVizbK
x5nLffOb34DEocobXu54tSZpfyDczEbZl2jqQLZeLUdZsduluzW2u/mbrQ2iQEKF
av6Ad3VSWX/wIn3t31AxQy+hO7u5wk4l6fSxMVPwu+vLfyU6EZBfABiMCMNXqGwk
immDp8rnE4sNPee+ipUShFFuHfiAaNbd1vKRpXY8l+LK78onkRZgFPtvhltcxZXe
w6edCI/nhgAJ0y5+jgqOdG2t3oZI8rcoZOiidnmJcFhYFHPKNIqg5snyTmGrUaDA
kUmpNPCOrlZ7xm41jOscc8wC6I01z9spfvAa0KkOpzGKQBRist6F2r/Z7gXu2j7X
236Qr3TyfbOVnFL2/4zIqTzSCBwYodqEJ4MlxdW3pb2OYklhxwfFyj2kjBxL/ih8
HCpYyspALQosRXHCGSM801dddGdonLoTKhXCrWpMZfrgwpU1xM2LEYyAlANWan61
AnSYEGk9usM80Cq1TgPebH7l+XbZUh/Jp41RsF8ZrXCaUJcHm344Sa1CpGTqdTX9
EppGjXtEhgY1g9H6e+FLAkpolZlnSjOWDjmr36YmExxx21A/84KBxDDOiPcST8sY
ySuPsszkq67UB63VNyOQ5tntpHWiY0NK+c6t0Zhuija2fMn2/pVhvnl+r+J8q8Q9
Hc0Maj86FgH4HQlM7Pgrp8UVVLkHSWmkdA3cSQASv1MY2HEjGuzWqwHBKLufWvVS
JjthzmmyvIxm84hUcY/XHkY0cVV+m/TLY7fBx1+8cCpw0jtDUWFG9xILwHiR7dwi
VgeFrpBi3lfs6E4FB5BolvU3Bsz/Q+ZkZSELODOkoltOazTAkND/oHLyBEXs8lq1
GUjgl+bvXOzwpe4EnCKNaM5twebz+0eHDpNj4yHMhK7POzxPdQoH2rWWfxyoeADy
xyG6HJ3cfvsiqhCofcSoC48lljFAoOhJJ8anDRxu3YH57J3wjO/y/f2k+Z8SUJGM
Uw3lMD8szySP8hzHO2mZd8QCzg5oixdl1lnCTx6sU47OOrqFfW7HvURaRQX7coVR
Qo3aucIJOk9rqKta+hleW4fauJeOOOoLVXRvvz4bmizUzfeoWfkW68IBYOydDwPo
CeCdrZ7j9ijCkp7h64C369BCNleGBkq/0V4si3Y64NWKxxyL7q8A912KOHje3M8o
vw8FdaVx0mYCj2BUknIx9j4TjigympzjMxSR493S+xJB3PVVH9uQGQJK1EsDvAIi
mfXlMnCBppVABZ4WoIDkkL0AzK0NI9bZY48RFfsV54D7LE+1wRC8MSnNOoCAIGdl
GJ6LimLSl7Jy0XMpXctTZdP657wGGpFrvOAfdARUb/ngV7vH6XpjqOArytAl8oaa
BDhyH7a17sjLBk/Sx4VyNS2fUd0H/GcuVLeyfetMyAWu/Hk1AKVTwA+D9MqC9v9O
p82Yi0QFqjvN8TE4U1Vhv68y5M2/CSfAS69/WLg+hZJdBge8S9k46ieBmmYcLZNH
risDT3Q3TPEs59k2AWGyZPjobXXETaeUP+v4PRufKDXDl4aMwq/vQxfRe41cmFHK
Y/n+kwsIdGW7/mReRDgketNx5a8LRS7PEYIompgivwAEY39UwT1EbCNZkyOWOytu
gWlTDJqTVAI15MOK/trpaj44+yv3iVvzVaHKNSZ2fL7I3M96/5WzxEevyqVXMcDJ
95KtTIqTBfQeHaY/LtCgulE065zk3hAIgJ0cMaZMdhUPVC2ytbdgQmXncaY/LVx2
W1zyZSAK+ExCNXMj/eNr/ZTaCzM2kpWNzYHPSzNlYbeWn0m732mpHbv8Xejl7XRb
diY7I/6OTCfUIz6AmYg7H5QgUN47YUy11LstPe9rO7rXxcYCovKYfWgj3jCIqBln
FYvFb7Ns1B3cXF6hKRy2/uOaBojLl5VezCE011T206gohaFO8mr+pRTBZZetQdeN
JYw6HLNtKOI6kE+giJGy/j9FF24ur+8nJj1uUx5IHyyqfHcb2juIbQo4vF5/qRkB
9RQ1k733FmvMHD9Kr6Z/S+4hhEU00QX9pASeLrVcwDBHg6is279h9WaqcJEXK0Wb
Z6yEafTCae23jhF0lgPfpheq4BMHcfk7r4h8f71dl9u7GoAPGp6Aso+jVpZ4hsXd
xcb2v7UUuhRYtrUxIKF8f5uyrpePrnJep/IysN1Y4txfVFokHHSDuYQmhWUZErMv
hGQGDKF0PNuu7Zcg9U//HNZ0NtWVEskA1Jjk+zU6wpxjF9E1InugxwYty9aaDg5a
yWLyD2JEJ+ZucT6vB3L7xo1plJ49kVTaRg/XSXZV0jYtuSN/MtUBGwrrnMe5X8n4
lzDbn8VOkL/vx3j4renFVNmuqRdxZdUXsbXtZVVOmDbG04QlDkhF6Cd6iwpmXS8s
PwTrk5m3zjhtBQ2TFveyJAbcAPOkftRmE6p2GVp5sfJBrM5XHGP8qChYQHMZzYCZ
LRaBRSf2Z3EsqYQWecp/RUZnk6hiZka9I/Vs+jVoyya7qsqX7MaLdpZHkgcADrXg
dj5kjUW8JafWjHCaDpPq/Lbr8ZH+m4bUzjC3EV8n317ZdZAtnd6gsvmKSVeAu1AU
9OEzZN/NHWut49MVQH4lqxJZBANlfp5sOaj96dqx9hK0qboJ1Kwm2JuS8zdD3a9/
s5T+RNWgHtDYeZXZ6DQo9YfMTc/7q9Nt18iRFL6WZVqugcCvadCZv4UScEEuOBGL
ZWA3Hp3rryWveqHC+c6TQIfOvBlnax9aN7GVNe2G0IulHrv6TwBSX+AKWwLAyGIL
9SVo+mKIo3PNbrt+ZWnnCC3VEUD02BAu+NwPGWtb/MKKZYtJcXywG9mzYHvlH6fG
JHZ5jxU+PXR4GlkyxktvITpWoSprCLHKyLD5DbjtwsLMc/ITerd5VUBiK9TMWuq1
8DQINYGddQmh/U11TWtUM1m6vC75WVDqmxSyS/uGfvGlDf8vZeaIOVBLTNErqBH6
j5rbbFvmnorQRWhvFIVo2KlmMI8RsFPIHY0tbG7ef509UN5ReElYCAPQiknhrFc+
Mm0h2quoWV6HeMox9yPtmxB5qEFollluYOEZPhSiz3JEfgyAuKktu9xuadG6C5M6
C7Q14AOxvfHPut9FbSw6j5/mz7hQhoP9NRxhD8CFGYUMhEZOHW4Czb1FyD29E87a
Z4omS6+YKZhwUdmNZT9nZlG8CmLD+Zf079rwrho2dBLcE0n4SiJI7d743YLK3lRZ
KG0XaIDYHGEakZhA8ejjBy6o70U/2sLo9xDkVgkY36NOugmTI9kvq9qf65mojAGV
9NRdwPg2Pa/RhNyuaeQofcXlsy9xfk+tN0ybm+1OZx8XifxKGf+qHksvTvIhzyk7
O91HIAc16clVZo3FozbIWVi+IJ0qCr1hTNWJQwpGLCrbWEj9AtnVmVTO7Ne5BiVe
sy19kB+RUqtwNW0sDKTSflsDOG4lKknXu6iYu/mjylSlF3uSfnlHxiNrnppvLtZP
9WX/gvYhU4IzasCs/J8Tevmj4dnYKlb3L5E0XxrfXnLjSOY6eECn2G3hxPcO84kR
6gCMEXBAiO3deMiffpyPe+Q/IiL4yZEnqWNCmD3A6mD9NkvPy+VTLhSqRCGqMp1W
EdpXScqVIjSq7922ms5bXo2Rx58XjhncbJ0vGrC6kw7LQOdYxMK6Z6u5/NJFN7Ub
bmpt/GxVeVGdVSuh2CuuKjjBWv9BWfmMnTpOpsBcfydVU1Vp3W9F7izxvW4MTXGG
UhU6ZaKzHXmS4J+gGFh61lgirvKUQVKLMNHl8QnA0u3A1V3OgXyBOSFY6hP93jaZ
BIcIeUxqyaKWFJbShUd2sepi61ovLy57ghaTQdjBdQfLLEHLgQnqkNjmggDXZEKw
ZljALitAL7l/OJHnBUaMlbhL6a1wbFNWHkRq1v6bLpD3bqtS1vGCQ29xcuQpMuk9
VsgnfmCCVu68RU0juYsn5i9ZscOLpSOepcMR32X+cEoGYMCW73eEav3F5GN1V56c
iZRf0XVjkWBhkJYt0sGy7jttLc8xQe4X+7P7PtU/IBe0tq85ahJHTK7xVjsYO1/N
DK6WheitM+2nZQxPPggbPDNYW0h+oARAXAosG0YCAdk8pLOOKJuMcHwOHGa4CitK
Xa2cniyoFmIgTxbp2Ml3re1zyMRdd9hD9vW9ZZ+l3jHUJ2QuaOhRmBex4GRWYuLA
Trhzct/JB5qNQkEEwpUcjKSGW52Rv/4C1Lj/M5mC4sOCUrrnbhOs+cWRKtJdPXnp
0pULfRyiy9hHwDBhsF7AgWB0BU3hPWidqyRv/ksxEZQsNwVPE74wlh5ie63T6AY2
Bc4byKnLVrjmYw182l8T81OJ4vfo2IpC5zgnPcOG/laxgLxl2I9wzvquJzxDDkSk
Q7cUrL4iBSxDqThl22hZCpjMWQeW+alOYmRGZvl366SV902GY5zuLUaA8rum848F
U3Amxj7bf7WNJrjvtshiTgkdZyOza6MS0g84b9+VY0IEeTxZRhWacP9PDPsgYXiB
3vuBU2zbEf72+Iwt4g4cj4AotKTouesijx3ghmLUoOhx2n5q9MV4shoSVtCFmXzB
KcMeXE8nN6VPBrNpHZC3IFyZH+mRERr2uTB9loV2/fORaDVStFeq/Vy7DwNyDNbz
GoZ9bRxJv6p2F+Sfg7x/75T6llF80BWkg4xBCxzP+FZBDLKJIs5UjyT7zqwpWwDI
LELtCs7Lm8/48PPb+EvmPuCdd1z/5WRpnYFPmcy2LC3v5Qun2e5HsJg4IJGdU2g/
ArqgkMa23DDNzRC7evyZ9jL0TLJ2fFc3gxRjk1bdZ3k3/PnJU7iLmG5NSfzHsCWF
WpjPxUt3cU8jCs72RRQxY4UODFUJ4oDqVGyGh7R+iSxy2jmmW/WYPVjjqm9HcfZF
cN6Uywg5tRZoMyYTeiw4hhktZ7I3WwltckzBDub8HxMdqOr3d28QYIcCBT0t0H/b
eWJ1ZwPOHGaNoJoDKaAZ2e1V68x8cg9qrO6GWmL90KFI4MsbVNudqBdcNqwWrHUo
fSKNzO7RxiBTRoEdP8xX/H9qxK/IOJOsZn2RtEhqkEDaTpx4SykFvws7MPBcyvwl
7bRM8OBR+xRhY5oLLIv3PP0xFAimrxs8bhmnlt528Bs6PKwydBIFW7Kx+C7SYYr/
N22ICqCEp5qqK55UIGZhHy61RCA26CNm79+NtpaeGtnNo8pCWN4Ba2someKVSpFl
VPMhN65QcX+Ouemw2eQ6U7+nOjnMp+KNUvc8c3Hyi/2OnbiF0wsbdhoHECD4gFrF
iXfqWNDEoGs3Jr5qZauUbaOJ5qGWBGBNTCHujvRwERgTIwJtAth65gCleUAzqoZ0
F22R95+LVg1Nns4yhlQKZpkUFB6La117WhaimInay94rSWC2FDRa8HHm2K7J+jLg
9vVMRiHXf8GLTUx7QYYZOeGxaHW9ObGjB5aRaQeQe86L8aoI5krIkF2ml8V6hieK
4DbGR9GLUmQMjQ80qBtwgMU/UWsnAzHrohU/mqISNT3qjLJZF47rdfqjA266F9FM
vykvJ4btCC/6uBVjCBQJhxO1kVVh3Uf4QdR05AFmuBX9L7nYIsotwDgTmCHdla4c
yuaaYb+Hsgn0SjwwY1aexnvdq+NIi+Uj0LW0EGr8eLurRjkDXxUPRisZZsJ+Vg5q
C9AdhpaxkFJwC8OXjfbeRx7WMZwrtnxb1V6KUPoxMI59Xem/iuBs71Veu2gZ1Sby
gOWBCUjDOXEE/kjrx9CSs4FO5iD8T93CY6mX9MbRLFQKqUj2UbSrs9q/7if5x3Vv
JnegFZETF94bFR3azK+thbA3H/LgKqlaKaOfUXvMrGtfoO+JeHG47ReheaHuZRWF
3ZCNbx8o21tvBzTmP9Z1x/fhFFyi8CrvGLYSz+rlsxKPY4iiw+gRcWSlqtGoh5/9
CyxztcLiGz068igo+ZzX/AWtzCpykITTxCw+NVSWr23A8HLFr9nXVNFWdOoYmr2w
5GiyjRj/mx1gA0y8P2L237P3YFlFqkgp2BIi5InPKp6H+EAS0gQbqai/Hsbg+A38
TOBMfrv9bK89y037n2EMYDlpTfPZctgYjK5Tg7oBdyfbtZI+jV8RF+f09fG1fdoN
moY8qsFh6OYpCtqAFpDNRMTqt3O/GonazDKRii1FnW3Op8vUMO5E+NxuXXiajz4C
jo0lGZE90ylmg/XRgbl8QBLl+AT+F4P1tQE+2aj7MrxTIXN3Eip2o1Mp+dP/puwC
UALSXdSpL1TT4AcrMT/K/yassyyz3Hr6fDOOF4r82L6jnNwSxuvXrHZqr6qkO7H4
JqTSkupyft9CeGPaxNCto1l4Ds6+2CJeuNGEl7FLiuuqakwjDCcejNoZ7qr2Ahpo
QEdYukBog8ApqtyoazAIj9MOq4CHgZmyHLovTrP6gAwvCbCOwHIL8nd6QseSP+f8
p2BFT9N33Z5hxX1TF8oYgOyKexuw2We6QcPMDZctA4nLN18tuWzhHR5epPVyvgdo
r6xxkl1A4rBoTy86qI1PF0VKv6K/t/VzXBART2aYXgRpVHTJDeTAwGvIstcMxprM
+GNEqTRe1XdobY4r0XcMEaTsLrNGfA83rhNrDnQUeB3APM+mbeC8WlhX7uhYcAEI
yBUZkJyb4+ZXSKPEv+ZA1WQ5cbJxCttmN8JfsjnD58obUTzLzYEjwplOhn6WJSzC
ofGrb2SqPJEejMSGUBDlEcl8cCXs8iJrnKuLi9MAME2qrgpar2kKpn/5TjPjv65E
cPailV9sy/Rupl/63noEOWClSl1AeAUy6U/8Fsl3T7LRR/S6S7N38XXnbHcXXd7k
uNzv27AWPR9yB/Bzq1ymw8BsNQa9wZLVe+8jWCwtsVa2iZ1w0BXhYh/8APxjxGJl
Dx7ChkyuVawl7habcMaKco9p+e3P9hynkMcz1A3UvZ6+6Oq8mFv6YL/BioRihXvv
Mf1OwiZzrT/ixwq5wmnuAhBbE18yBjYcPuspSgwbw1xkVPiwe+tlNtJYnzCSe221
GWKp/Q9CmWCiivH9AkP40SjmVzk/QzEicc7BYzxm3psFYUX0hYZIxezJxl95JQaz
hrEvjkywbpcBBqJdGilb9MzBU4yn9oRnqR4vbOYm75nwmE7zyNHOJTJNRm/9UiA7
/51+w/XdavKYCMT5D2DE02LBUEBedy5a9mjgxns3OH1ZWqGhBuCqCwqHKWpKJwNN
uu3IJEBI/YciyeA2Oegu2sLUEZV4J9H1CrJPd+3xFFtIKHIj/SCeUhwX1ke9l92J
pafMLkrD5AiB68bf1wnm017trwNihlKqarFlTKDYgQx4K6aQDCvTn21b0U+4gW7l
YHPsiUgGNP+RLEk6gdN85SyMGufBUv6fdJuExkOXD8TlPQLMUFFdV67IGbstZRSA
AJ6/BmN5ZdbLSXNy45wApdFo8CkuRTA09LiA2VfyCJsOQ367MJ8IaPQyv2pUO+xK
vQKtlUTT2DheVTrIrxJ8DiSw0FtgtndT6X2jfoNh/vdrAU4psR8k8lxnPIgMjORR
NHmnLUHk4S2qQWn6bjpqIxrKP3OswFUBBhNG6huUmv6poRwtsjNiYiuuffDcWxCa
JVMc91ZlKDPoPJCwRPLZR55ZWeJtCS9AhnqL1srY0t6x3qC2GjngLLCvZDwbe600
/XsvvwWcEEzc1vKc1QfJRXzq9jx8EWSFfDIoNWOC79sDXpEmAxCAXo19UgY2Hmd6
8FMgQ9mHUqrNJ+Gm77Hb87jBfWQid3MKqkMf5FHXvghi5DG6aHDDg7dVfe8EADRM
4+Z9z9/UzLQajjr+ze8De4bI/sns08gpA0hTWrB68v2uAPnZX6ozHd0zugwEfsUt
uzycXHcpY/vep0Bt/b+rbG+zSJIulvKI5Vg8kdE0v59equRs7meTCTrm8nlR4Ubs
ZhRV+UPWW/Yfmx6jd1zBFwgCeNuKC0gunYzQlmTV6sLfsnkCGFg+tPedCzer6ZO4
pP/Qq7p5nDBOi28CYyoINLBy+u39At8JwPkTjSctXOUtf6TcbFb6Ow906uhAbKPF
y/mi5YkHnlSw23BI0TjTwaBuUCAk4S7FEtfBKVRd0Gh5eLiQ5D0jn6YIN70wpx+5
adDry5J7WtxwEyuS8vBj1qkUE0outeuAxublUhltogNh0niyCMA12+e3o0AjzWKZ
ia4zvkG94XP4pY3QqVPz8egNRGPqVFbw87ulT+oWl8/JzaRUtGwGG+Hecb0359qr
4XOzvE+umrOQjB8NFMIPfLKNc3W4ZY5LVO6RmpGdxDQHGqyWu7QMcsmLLIrAx3mA
iyq4HykN1JBWzk7VYLz5zbObWgEfHgH2j9wP/DN5fjT3Km8cYMjUg/mmSf9vJIji
G46gjz7lSdDyef8LP4hK7+Tc/4513wfuj0LKyd1rQrx6125Fvv/j1yeuXWnM6JSS
iUQVzz4IZnBYO1HLge8bqXk947Ntij/h0UZsBodfKz6y5KZuLPv8CPGF1VAuIDn6
clDshtUp3tBdb/nf+kkXPrb/orbji9P7UlL6JpYNROm2yCg8UhxuasT99FgJfMQw
GlLjw1omzwjKMaBGf8dD2W6UCbGEjSFTG5F9dLzGJkM3KA3NqjKi9PBcIzOSA0w/
9/pdJ3QyRUVIVyHqE5CZDH8bbaJ9WXCX60FIXdDVgXz8sUINB5xvCemtwILSZhJK
zyeeksonWhLuJ5KDbbK4Ncb3uwlLibf/VV8Zyc3/7wZNiL3ZfgpmGF+P/PluTDkh
TeGPJNfkfS31cUsiO7/iVlONC/iDKB04buRyA1DoFyjHv+MJLkijAhwUt0Zadt4k
9ZKwA9bfgu7NLYjD1vWJSrcaT4soKXlFry8qKrvGffHyytDqoaKMQRIkCICghAmr
LUICGtpevTI13tiXoXQNdIjsvEtTEQ8QNvZX8LtgjQ2S1Lti5T+CEm/FfFDHEW/g
TTk0j4eqFQ5203tnS/0oeWQJ7NiBo8hpTSSSSnimpRjGsn4p0Z4K4tdTC9HJlAuo
QGb0OwlArCGbX398ENefnkf8+u37n52eWNzg7N7erQJhV9GR7knQZ/wbCOCNZvod
hG4Pd5puKrW86krPQ8AOK5J95QQ7MpTtjSKdGXxe0ixdesjvjBPffyQQihLQM7BS
4wwaHvv+9nVPasSRbS3OFSibyfQEmccduSd6CoCkLjiYzXoxxtegvyJWhcRvjcio
5cXC70sobWdnCWyzA/wc2hqeF3fT85G+DYC9Kns5dt3vKZz0Q78OJoCEvdJFfjDE
KrO53mGpIQ727J+iH05b1ioTYW1pC7iMXECHOJZU8K6V0FuuNzbac5mORpAnUHds
ZhMgiifF4UcTYJB+GESkypmQnOU7J3qvl2X+H+kz4gjKWKjt/PklxAisgbuxUiMS
Vmm+mpS5KzSxANSYnZ1pPAKnaJJocOrT7lON9zW3xlIYR9VLxsxT0vpJQflnHGq+
46eH3XHTa4bs719+Dqw8NtlmUE5jRfw6TNHJQU22RaibHthV7x2ZjPDAf4YIB37N
7Ng1w0VUH7PPNSqw1PZiHVWdwbPYgnmRC0xSrBeOt6QHZKhnb+rdgetaarMh/CWn
rOItGLW3OvtvC3AOEEFoT1Lu9oSvlkmNjww8KrCclf0TTPoGLYkH5lDjfbrL0+24
BoUtinQCV6yEuDOeL7PaDLltSchMevbtqNIsV1iAFjmgaLcz0fL9/CuiaEHniJDc
xD2Lx2eBEKFT3N1el7T58w02b7qcdZh9EGqVsbpWXz5PLjle5wVZrKqt8zRGjim6
UVfBrSfqZOlKgS5ltP1Lhm9jZ5qgdjuD3b8R22GuRoHZ9EbaC3RiTDXcX/QyETeP
ftUwy5+TZo+s0WZO1MCT4AEIyMRX3wWeGlan6rK954NbRym6a8sBVR2Whjgwh8zJ
YJWbDygbTU3PpG/ClKnQ0tArI76iYLyhuYJh/u3MroYkXAXEdAIQEyajg7HyFMrG
JUq3OeGCW1SeoyPMNipqDvxmiyOHQT2DYvy4fCGDWdipljFFC0SUW6wVxJzk5lVu
20yuavgPk5xYpx9b27D7vg/bRGhaXExhVsqTKgJvc7HUOLuL5V/5GUt00bzjbg0f
MtocjkhC92YBMy/Q8W7FNQkzWHYCwLS5ZP4Jy8OIjiAAgWOGIFp+uwkbw4Br6RtW
HK0hqE++tX6iuA4kIEjKKMnevJ+xBFWhpla2oA5a6eZEhgUf1diHeycOxCeocRrY
wFIbHhKilu20xREt4zTHz/WjfJh/+miDJOHoAhKAsOaXNGXM8wMXHRCz2LiBN3lU
b8z26D77jqoH0jwHxQ8JLwsr6VK4vz6nasFJQAYFKayzLUiIDvKUxsyoey75S2RK
ogrF6i+OH80GxyFGkyebJL/SsXLevH4u+xrL55BIeDHPrdCInGE/Ouaay4ZuhHSs
OAWC7NmNTHLo1bIIsV4o6/5N7N0UM6p+w/Nn7+wbsnRzx7NHf4rK0g3JobyiGJde
6FsJK+2R7YAwiwucX1cNW95UWX8H147l/vTtR1SC/iWCPkOE0pngI1CEFUvXPirg
ARhnqWtumTSl9uaDqg8scWUfuvBlca7/nPVuwEfXBnQ8MOWWdrZ6OOHBdrNuvlKz
0UITgE8p3WshVudC3qYu4jzdRQXYZUEVRBixCGrhHNlaPfQlH+goRI9acfByIHMh
NDQ1N+atamFNyR9/+u09mgZBPL0ly4+ZVIk1nE+YPT6fb1nS+ouTqIyG7k+Bv8J6
PE5x6E/SLl4UpRW7D/e8icBLI+ioRwqc5GPFuxq6ut+21PFBUtFcHbmpr2xCHgG4
hdTjC9viw58+bpSKYzQIo7DYu/uG39aEmdHMDiBb0277rsvPeFWgPjkBtVme2vEC
RQMGNi20cQYkSfZha8e53fLV1re7GhWUhOSF7WuE2NpVhaFnULw4zcuOEpJSpLhA
OG3vtxUqqH/YZKjWTsrAVSmd3gf/MRCPwWVpRO+O67XwMn0Z78iXcs5Nw8PNhtoU
wJsc7jC60o4KbjVohYQZpIFHuYlLCa7EqoTTYPiRaMfQnSRHhGErKZ4sqK3IOOs5
H6lg8rb4/1O1RW4NtH4FLRM5bLHc523c7P/TCXy+p5P7rnzO5TLHIac69GFMOYfC
eyMryj18ZaDMtj5G7esakcSq3uwrurffwsMxVjTTUy/ui2fed0zbGIK+d6mu+nUC
4kSvG/oh05m7bbiTPcxbhTBQ+ozhvGL7GJTYlY7ZAyzc5VzYBJJdwJCg0DKJOubD
FUFIULtVusre7jtCSnXbuxQq0AXHfY0ustqaYcaWDD3wHo3FJ0zlOvkOGyrKBb14
iNAxF+oSDj1LtempAw3Yt0z3tZ4NACypORPsXB1a+QnuSpdves/aYo8f0HD1W+4E
c72JHCx6XbaU9qCT2MbdrDndLbFyu0ECJalJ6nIl3EUZpwkYPyAXs45Qpr3doXMr
Z2qzPVYlVMSevxynPBsLxlLf6B9rdQvFfqesL7uL3gcqo/V/wmusvDP2tpKSetu2
Lx789rCi4dDyIR1G4Mf7e/mo3bmNElrswBcHlIJvt1gNUck4VA5+JiOVp8XGvZft
GZRKZh1K403albslyIHAMUnvjgUwh8HS+PfwzUJQsVUQdDq6AmOAtXL10MqNxj0c
Rk+I/Xu0Q/hsj6tj+nuv261e5+B+us91VTKW6fl58cllKedzEDBoRs0X+J2u5xXE
dI5qBcXDuSLAFj7BghRVvUtmU3Y4fsiF3xyAGVwlD7LETQ0DNJWfHswv/JgS5sZK
RHdP3AjVQH5rm67AiUUyYOovBdtGwaCso0D8lT6a3wje0GPn6soYWYc5QdY9OfTA
oyjUHuAerTKtAoNFdpsKyihCmALXq8ZjC3a+URCdikQiHr3XlwRZei4WBtdzqoP7
JMRMCMGTTyvszALwULqxo4IXclYspmLp69/RPZsDET1aGIZjPRn5K5LEp891FZkb
nLAIcrUp6hxAI/jWS9LArjjxLVwokuAYbKH26FfCi/nRLw0CBnVkpt1xlVYXchsZ
Wi61wgrmlDxru3DKO2vk1D6RwSzhIuPmyb3+AuWAKKSdAblLlTKiCiLBkUgeX8/v
NCKR4SDbgUQ3VuEYcZK3iuWgPaxLOiZB2es7uTtK0t8NIDAB9PoZJkI9SDj7zS7D
x2D0KIhrHOGwmnB6wjMlKaiMq7MJvvzxlg3X10xzwhMs+VB5ZgGaku4hedO1lHFy
2WDoq7ONySO0a+W61ZpD9eDL+BvS/tOvyo1grjmDlHP7/uXKmNVEXrx1Z6VtuoCk
6iiZpyLxHQew0vjZfuLZVDX0Z9Yumh3ck4T8NR/S1vkuMS2U6QvSgHBvZLG12I+b
g/DvP8OkWj8p/UjlG7GnJCHkD4v4gZ/ihpnWp0zf2gsFfTu1wF4cxCXU7BBltYeo
F4dW5pqdjASOcgQeBy/NvLBCaaKPxspvLkA3hPQgyCvS4tdILy6857ipuHuI/aWN
TIKhXvRY7aqtJqtqVj83MiAM7/MasDpW64pzuDl+UahDpcucqKni/wBxEZCRktFC
lGttvOelDi75LQ15Ciuu7kOJKATYKZ/mtV/jHYDfErK4xtXN8Vdt2UplNv7jekZP
uzl3Si08k4BWDUN8cJJFG6j0cpu9vL/GkCV9ofRzHnLmCXlljYJc839uG35CEKNh
UdsLxWaBdwBs7Q2HIOLXpbXDT5mJTy4RFmzx3blHApLy/X30U/TTgBISU2KJ4K+y
iwshZ11v60aauUTvikbPgDCJC0UdZYImcmz8lLqq9mXkPtBxuSmepmuabgsvM1vs
jEOh+TtNmmAPVUB5doJuXIHqIW7qB+sqfsWkV4GRw0K3tm5e2rq0fl5CBGRdpNZU
QcWYL4e2VV6SngJFbAvUvuqXAKVUwNP5+b9cp47KVPm8WRzHZGG/CwXpjCb91EG4
fmGgJsazjTf3EFIeMtx22k6C4D0Qx0P5ll9ANC5GAJJUgFjQy2Q2payMz2NTY3VK
4WYlaX9/OHjhUHoiQDDOp++rPFWxoTuAQ/hkSaYOuow+W6AmpPrV+V5EGLvxG+cd
HKIPPwoTo3PB6/D+Xf66bkyrnJi3Xx7qFLZ9VS1K+8ahMVde1z/guJ83GthWHTSl
83Hr8bjKjTR8mLzmDYNhSHWgNqaAil67qxTDe+M6FBeIvWlc7uNE7buMu/62X332
EMziObdO1BiuhwBo6W3rv2s1noNjj97cSwnup58bRym+v+ScVZ/7wYYxnLxtqudY
mlkiTjrgL3cRwSjhnL9X5EXY8F98w04P8Sg+5d0TaiBq8XWc/UydjAf7GgbniiuQ
d7N4bvyQS+OxEwrnzaqTyzWLxyTiZUmiQ5Q+OsN26lzkWVBz9tJ3QZlTbzslj8MB
g/J3/2L6FZJ3u50Q9YJ+eYsMkqoo4UgXAg+9KJQdGwkE8FwICKVECD7xVTuhjmMX
AtimEtpNyrdto217pR8lT2aNie4HvGH9W77HXpdhiwIK0cZxtPNqhxiRWG4vu+jj
O5ZeNdKQ1ltKY/FcWciSNEVDP/z+7mag2F8/JkUvN7JWRss+XVBLzvi/4WeAXFhF
h/P8qfLVT4N4x0scfZOuptzP+3dKptK4oVEqVxE6PVANipSa5+5Qyx7SFS2gmxLt
18+LhSS+ShMFTaz5NFxwAYxgdzh0UyAndr5nV+xQD8dLYV0SCp6S/PGS41VFNWmD
D4FA4H4gieK8PKKAviMOfIz4jE9MrHccCAuan4tIk2IzuUiTM1RdhZdjbxq7nIq7
rwSlQmsMqI7eeU0QiamDvZUTu4WZypA6WFA7NvFcvGpZLcvc86sOvi34ojuxbOFs
0uaxoemVUP3Rz9uwmEG3tvUTF3FKSECq2BRpiJZrhfT531x3e4gj9J93D1mkXByW
RCkifoiaXgdTRvuyGYS4qpiLt00aj64FKBuSteaYL4qbBUXgHtqSIU3CGSfeyYMP
IEaEYUmZogbPGXKFdlrtXTFLYb3NEvM1AOSJwKVT0jRMkmP7YExh4bhudUExnAKo
Ydcl+23hLvqI1sx+72U/+pnsGJtf+jien+nPTNY6QlYtS/5oQLDdBf3Nto+/r/Bv
HqbZ+Wfkcv4J+aeDQ8mDW4A1D4X9qPcL3z+he3df5SiKc9RSzVaWzGAGCHEKyaG2
cD3IfYIF3K1nr7SY3r/7rz+q3IAc+OHv9Zx17NPzVemkLj6gQDrbScx2gEhRed7U
880A8SpIRKra5Sly72e8Y7FXcQwF3+eNa0uWjVih9IDveg+u/bim3P2CZsxHGx8+
qbMLFlxIe1y41NBqLLkRsNMtouVx3B2itc/uyLSsUFcGbqIIR/HaBkhip7jb1At9
qYXwiXwR9PtEGISjjyP1Zf2pqC/lFsE8chi+8csRRiVDhc/NczWdG7nUvIywoQJT
3w4SUXnvwB0M/QWJXywmHRsTboeBVtNVZ37RU+lUOVBPx6T0EOUlLC8nQIoWvqzN
+GgbGYlCWgF2bElPWl4mSY2fmpkDFIyGBzTBpenHsW/iQR1WX8VTzP6b10DQAYYa
H0J9W+zGmsI70tKaGzmJQjNDgJOgez9AvPrA2mUAFg16dM5U0UgEj5T3SsP+b2YN
GbFox/Vveox5U6lzcYnxRMFhfUATXqzONyl5cGD1gvrkpIoTBaBxvaENRsZ70oWy
LS9BIsyJilste6GfrCtbo6OihJsQ9fwokGSwAMtSZ8lvgtOcrXlzY/u8Qv0ocTsj
XVjxc2efRd9u4NAU0E+l9f9dZY88ulb07LIZYS1i/7sd1g+gYGKYiNRaOQwL84ik
ednC6UlTWlkFvZzno1n4GYsydUCoRv4VRHqJiZNT+QSh0WS6PzkAHl3EBoeweb6n
qrHMDn21kiFff1Ig9qoHWebdbckskIpTk9WL/57IBDHp+0fYJu//YA8QGht3Kpsi
oo6sliM60hPojkWyhP0IN7IFgTdoIMyYaUl2gdTd7N6vb9gzST9FpXL0kMKxfSjE
Fe6fdBpp4dHT/LAovocRv+PGxOZNxIZv5NyP6S6ihStOycGBLBz+MoVfzGc8cnr4
VA4G51xXYxipQsa6D9v6acr/z7wg8AG0OJUtAOSDpHi6dF18Fr/NA2o5VuEdv3cw
bb9pTQvFZy97XpgtLrlQ86ykYURfBDSqFq8AOc2XhnIN/BDrzHJN5IkJyZitbkQ0
3J509ZZhD0EAcIcFWm7NZhxefCW1zUBG7CUrI8yPf3VSOqQ97hZAn+JPuAZ2FM/r
Y/e13nMVSJxebDr2uwzCZvaLuF9Ou9ACo+e/Aw+Xzix8PT1T7cT81QjYFBs0kIDO
XhnX3o+e9cGBmrYgnNsp9Z6pHkCuW2kVxSwDI1g4ukF69teQGmROeyaRH1AKJm0H
FX+FogGavf61CKwVg3WeouUUx1vtLmrmke3R+Gav9mimamEcBrLc86x7JIPVtMqV
ErjWKJO5bfuWJybgSCEskCAO8dTjK5UqnK43dfK35DvKwWPoKIDkvFNybHcJaTK+
+Y1XPHxFUHY7Yq5YtCafJaEQT9D7/MTGNEc3yEsBAETQT4YEmb6qeZHWTiKN7Ubc
RApUCmC+Fp53ay2flNpBHHgWVMfMcfR81QABIArn/6t6+DR1ULgAlwTEAuiVBJyE
VOoxuZkVGUfPGeUpKnV8xZhgBHS5xNe1YENbKton2+cMJkJ/qESeWlDa3vGSMrMe
wYH/9ARtap8GOddXS2gaMEj3L0D4iTyNv5DbKBQsln4663AeQaKoFUFUWQo4pZBQ
OjHJFVi8mLniYnDCbCfWReCVme0qV23aFMV5UIUzyKZdBMmnGIYvqV0PwFz9eIGs
u1Ra5QZm2AkFo0bBildJ6j+UED1EpG8UwMgJfLxfOkWn1HP36OvO/5K69sdhhB+E
RNavnoc63rFbC2Z9Gs4stQh+aVLNvVS7Isr+S86y6CmUA7NaS7CqwwBcgLPLOCT3
DdOwOvbGk4IKzre31If8KBq7dqHYpS549gtsj8Z39y4Pz6QEBTNvakivyrAOOAtT
y0tLZQD5JN16x3zw49NUn/UACZr3gcmN3bWb7enwBDXgzRdeuMuemUBPN3yFkLbw
MEXNxBKYSvSv+vycspLCLmXHdWpUtiQM8/qMK/Bi1zQ8JOu1889jsXiriRn1HT0L
O15hXc4nlZlwHbDekt2HcqfeErEVDBAzeqGoWEVaHFLZoHcBB6sYJk38n6jMd8YS
lGgdEDsSisJmQANLCG6a5rf+1BFpJxcAF6ehZUFt2/FXPkLTUCbqsxMRmnbXeh/W
vnCPDpikJMJkOCQVPFW/8ThopZIRWema6w4TQVxe9dONrK84a4DcQYEUaIotkXUf
4P0tiOhBfq8rz9mm9bKDXCxTQK8FMRqD/ta3hnfN48a+1GnfBPgd2M+7v6K/6rzn
q4YFE0G5o2KAZhOsx03eCr0rFriiCVhuNlUPV1Cmg2XG05lpQwZl7B1iQqJM4Hyt
Es6h/tKkfMAQDyAd30fLNYVYYrhBEcW2rpO5mLwC6iyYddKNw2uP4otG/Orio6fs
NN34v2c8jVF7aeiWsSrwLrHzuTwcVFdkKsf0RRV4V54wtKN1OFa4bVcQ1PpbmnWH
H9eTppQulRX5//huqZcy65LEn80XRKIkE2bEuIYyqd196X33ORJMjMkM+vJoKDRp
Rg8tTklGgXdgPuCgwFZTluTFnYe26PZWv++8f/Fr3cTLEXa58TtQDBqkCgVPBkc0
QSY6bhN2bbY8bzsflnBkDkn1oQBjbOMqCbcZf0lzcIWz9wOITWRHiKHNdOafW5dH
vrtQNe9ImvyweENZzlPZeJeslesjeDGdjwddiR1JA+iTPwBckX8qNZuZit3QTCmn
Qss3Dwmxq3BrdWLVSjfM6kg8ybY40Aa2b4l7XLKQQJEtpjwlYSrfGnDfdAcBx58i
zSPNwBKz9x9ArTuZifAUE2oGnxQoTtmIZ7T96UmbAG27/U/xNymUu4UlBLqF6X0G
563BjOKYU/mqCjF5moV4Hb5fb+UNXRboupUO3Wt9N+NAKLTHR3MBHK+omloftbGX
RoSnTRfR5UD/tE6iuR3BV3b3Lw9pKaCNDn5SZHe/TqULk1T95tUnuZ/UM3OVqJhH
gTc0/f/38zGibTQIzHnZ7yDNH16wupNrxdN5mrpzXxWmFPAKwYvqdNXoApG1oGZg
o9/CjyXF/Tkpc8R7DAqeE0iqBLOVeP2MyVo4Ed4M6tMaeWSKGze3gI3MiuMRTc4q
XewW3DPc4T124L7JQoRA7F0BbvZGJ2usSbhtwMteRlBYwE0yVpBkLwGTEFO7o3Xu
8NkFqHwNjNNCttFUD9V4Iw66EINrPidluZlucUq4L4fS0wlbh50Qv4siLiFgKJ+g
8bwHKlSRAyzsjNBBauES8V3QXU+p8Gei2kFgoE1RxHcal89zJRGAVdTaKkENsELf
o3PJWFom80lDNh0vIHOBdUWd9vXLALic71Cq8DcmnUaG7J8ohQgv1hWEOID+WaAQ
nbAvXvn6HhwnAa6hEAYhBDxfYny/59UKIQWPoehWBI1H1w/fMzVVYQ8NLsyOJN37
OV3fSTfcy8Njj+36ijBIH0RNQRSNTBixatEuqs1WkMBCRopw/m0rJg7U2VDgOsHw
nHLLSrWYa2/stJOGHSdtEdozmaBogLkWby+Mh7vilCZJCDPORdRCC0TsOC0LNhd4
EDgjoIqRaaj9yUNEIZDN/OOL5UENai7d0DK7VjQxYSfTctVzwF1NfNSLKI+1wZ+8
fBYiHdfcymRZzYKI3z3pqQqIXjqCj4sNKmvxkIkktGVOUJUsdX9IZkuKABsEH+N0
tde/KTWt4W8UK/1qqj/7TiC7NCpY6VS+VJnnL25t7YCTMzJpyr+OLz0aLXJgCcot
m3UimlluZcsHiSGfhXFEbuVhhCM/fXtU/JMMFC36OIBGCI5be8MOuKdw6GGupl2K
AlLAp+sijHu78m1RRfEY9UrrwZ07vuTQ5lijG7QTH9yLE7n3iYQJte2jO6SiehzL
FZovNi/g57MVkwxKFGVbMGx4hW/ax9pN5PE9z7jZNELYtLRb1MvbHMxQzeciK/TA
supHB9FNcPY6nLL1Og0p7IHQPj2ngerpnzafc7W1V+MIBRtoTaEjm7UwVfYol049
IFIFMKnbnvqGY0MvKd93m7hGbF4u6XbuGeJ/E8RMaiQXSzCwT3yyt+Md5jdICbmi
pIbHvmsyPNplHcfwZ+qMRBb8J6SkZFWfiRrTtQYU1oX/62BARDRJOYmy1B7H5oGs
fgtcWQ2UYcO8erXSsWRAHpvhvsNQz7ZIqQutpR4HNGRC/L3zpnhJCyqOMF1ZuDNJ
ZdmffzE8dhuNOHdqSAU8sFIpqQgRSHzEpasn0awkDEtoJ9/aJihfcP6MxmBU6bm2
7kuSVkMZOk3Bv0Sx7zhicUGtXoNP9luFXjtXP0YX0DG8WSwlAvGKogHTK78nUx9S
hfuZFa2uxLES04iikxnZ3//Rt0iJRLWJKalbkpgm9rMNAC8AeR3vHIyfI4AwQFmF
xweGYBcYHV2Lm78qyaufwrBMYPwJgIijxX3/g91zDmSIsyHjvkuciCbH4AKMBd8K
VxfnbnIdSEfrNlLgBOkzMr1uIv/1B0QXwwPLcS2jbTVbjQtUk762YWH03h+PBaJw
pwApSEX/FtpLXUnEx2oHprMPJI/6NH/HAxVH6J9r+QSWcER3+veTJf2o69Aamh1p
6I04nsXGxLymcoy3R7w5RRM5o+ERYm31C2ox+g4Sl8OfrX+Dz2e51nk3On4fuUC5
AqGjBlw92ZDceJkcO/frFDCEOr9BYq7eqi6G65P1jTjTOjEupcNzfKsqiJBF+EqA
54FXDqkpHXn61L3Cpx/xW7uKbBwuWqX+AY5o2wZHqIEGNuSoiNf7v7f3co0Cqijw
vC+RIWiYlScoXBiOKovk9VttgHbxQagQCHR6/kJDYVIiXcHS+BQOV55qmNa5CAPG
cg3R+y0Rl9V9sr+qmNzvlvT/6l1ihJbxWg0RQyx4g7M+0FKU4ALYdCgurvB/+WtR
4dbTkAXyIaLRjMaBm4W6sYEs2fTCoLrD7beaxJuP5jLO/yZ59MurUtD2HijEHvmW
xvRJ6oL9Iw7vKs+JekSegYrl8c6zKdUGSolZF7oHiFOiTl8VV+Khk5ZBCxIHRyWH
1liqZo3HZF9OvwEIPbW9LvA7z0C5oSIQRT641YtuVBE9LchVFA/bLE6o/YE+y3iX
Zb26CSKjxYo8aZT41bWDEHKHbUs+WhTMZ/+7dOGnxlXKcAnJYuwQxCKPb4Ayyz41
wsY62rn8Ko/8pTKCMQLgOy2lCnZHfJ3Ap7aCwzmX0dW61IUQcZ7aHKVZCMlNB3iK
v32J1YkbHHxLFFHd/vLBayf/+10stLrZWOLxKMseoukai1OFdxxtASwBQD5dKg1U
vYstvGnA+1ut+T6dx9eTtreFXyNtDpR3wVk/K7dXA1ZHc43Y1O4zUs7+zhz4Ugk0
C+pmw5/lwZ6ewdjTx95rV8lb6IF/6mZfKJwthZT3XpTA2FwZZibwNcCdk4TftaW5
fugTG+PI1dPv7TtZiHxHr+p/IH1ucXHc4LNJvn/s8+ZGhWW8bwiPo3NaVPIqqG3T
3c4pYQbD6Fsk7UByvMEVkMs2KFRmi5rnE0DJv+pk8O2yIHluIi3a7mqFPQghKBUD
df1vvau8VtdxBTEH0YrCrDoEvR499tormee/fo29CIim/0ENYKigSsPsZf9qylpE
oA2GdQH4jRYoRCQpdhjZNZ7ymoeTf3CFTBvKoUjwza9sWXimbu9/c/6Q6aDXAOjM
olr95UmNt8pA2Opir8tFnJYHVtOLfjU0I9G62FsEYUd7wdTKR/cSEDgXrugKQcsz
Ej7HmkVAQIAdRaO53W6Vv/iuG0z7KEzONxbyKJCm9AWO80Rbe6cphEVQkZhOwuda
kByVYiQS3IpHCbhJ7UhC9qVr1kis5Ikgn+LFeJmWT7QMWXTVtix5P2JmzPeKeCTw
vIpdM/yV/r/RpfnGbPd/YKmg8RPzogmS0mDFxC7FvULEMMIdIcVSpVkHCA23mBfB
ZglB3phXMY/hjF+9tYzBFJMcD8sYccB3XLEHYoQJZDEMEp1QerDY2mOq1iahOu7S
QrNqdkcqYfKhbrOZ9Yqmgsi/g8QgxbQMD7lcjBHZAn+Q38WTbeGhR/q+hv1ngtMv
u+8Mp9VJZkc8urhZv2HYSoNPte0oZtxnqJEgFfekd6HSsT0Tj/7aynqqQPJMSuF/
6/BdGgjj63Ga4SZdL9KpE3gSiBCm4mQvHiXPwNP+mIy/I5fX8vsyA1ZYK6SlX/Ok
VOZqWGXte+ezo4X8PntqJhbdzIt5FWrit9Sk+F12ZMbRjRIh0B3ypaTqR7LVJiqw
35ZVSbdRmuvh1vrrakIC8wgdQdmuNliF3NfGNDf/LnWnVZ9EPnM9y5fmL0GxnVAM
vHlUCBRkAwB7gSoAxY3rmtKsDUnAHLiMCqTbHNKkhWfnj4L0/qUT9vYD7s4YDOoh
LQb85jf6WEs8hs06vYL1Lzuwt4nRxTnnYRat5PeVq+4//LSHS/xmtp8tpQPP9PUh
9ymXS8ZWp44to9rM1fB0sgYaihvpVl7AvwSyYbL2Ihq7epyAKwO2JwgjOqm9yjA3
RApD/a0ZRms+/8DBdmFWoNa3OpqBtHfROD8ZGTeHm4dQQZDqUpJf6A0YmZO9yEcy
4pJrWxJDYT5G/QduzC1ByCWdlP4k38u8jPiEiwgkUyPI2yPC6YKcqDkb3h7W7aTC
fAEWul0ddfVmYN25zPAXpgXfUgXeVVst2WGf5W7xX07guBLG/RFG5as8Mha/2m4U
I17rs2/JACDoZI2SX/0o3t1dB3spVcgSBoJJmmTey2YIoMy9goTpYzCSKtOlvG+L
Pr+PER3AiiOuxjSy4O6bhSgPLMsckbYO7lnMK9wht/9E7YSx261q5lCbm8KhHbl9
YNSRUUusrJG2TfMIGduHNwZsAL/cExhaBt3C3dqIHCIS8rVedi3JCfx4mwIYQnK7
H+dLcISK7Nw6YKlxAkFX+9AXhHX6OE9SPNMLpWTiOh8cbu7juPodoA5q5UZNIycb
vHQp1yvPGe+OO6qyJSXUBGPU7lTSpwTlxv6oxELtc58CkEJ9IhkZjz7MpsTeukXQ
71Y+lNer6sWSDM+e6p3iDwEbdPmiTRdkwhXwRB+zEXIuKntXYBjtWneCe/VjScLV
s8xJeq60Rk22kyPR08ur34Fpu91Qr4P+/0kPOjt3lIiONswI2Y/b/Mug3fgx05Cn
9js4l/sqvdM19WEMa03+9Xdz9FepsIDIdX8SRl78hH1zpRzAWDnEL5nYBtQd+dAD
vlZEcwjNctXbeiQFhQxjRjV/waXbFUYT8N1pacKGPRbWib8O+jVHj1Xj503ymgl7
h24CNksMH56xSjMpvJtGd7oCLEWjyeZ1I2OiaHIM48tcIFPJLuLutNPGLkgWE1ai
OpavtzNXZ3B09iwd6x9qMxiUAfsBTJqcWMe7Sxojl0q1fOEg3yevwzRHty08hKVz
ncIGYt/vW6xX0LUz8ZdKx64hfR99bhq7tTP+eXZLeBV+HIzdihnEPks6EjAO2GB7
zYEket02wqZD0xUI2dzXzbMX1cv7vWyznNI+y1KAgw6FXmcIxJ1E9NpKBEqqEWQ1
MsSSR2TEiiCDhMC7R4CkSb1kMxDj0eNYpWqpHfDBx09NJgYnsDxvI2+EkO/VMpQG
B1+MkDo6D9opqxpYs7mTVCJEhXjdFbX/tfKhj345o6D5aGnZhu5UUPoOWkUGx5ni
7IMabNTxkU+YWbWP8iY+ahiXnGKF/TUaL6S3ZZuidcsFGSPnLrw4XTfIxrxitdLV
K7Mfa8DcQmGIQ3n1DZdv1oUclQnSqgKxClHV2/5AF9LKZSalRsDlmL8SX8bP++YL
eUn/DsRgFzp0PPRjitW5uoHF3re2wT6YjOsY1TLbwV2on9XzyVfwYjOCidclZv2X
k9w2L0NMlZsUfqdRYVl0pzmkGYvwrXjmc4IsBQjM1yPcK5aLZzwmBloqkGOednns
aSuo5nWrM+FeHbzf2PAnCv6iMRQAKpwLWtGOjFjQ15pZMdxXQAxWH1//b5f0IzoO
Q4axksdkhKbODLSabyTSAJ9FIZKENiN4d8UVGqpaIz8nXSKUTawCsotUCDdGr6Nf
XTFxiVg0p3+cPPGtgn0m97btZyOc6VD1fM19277mhLqqH/UJAcwjPfdcfSyS/ZrC
VgwN5DiR0UxFI6I8PouPyCpBYkgx2seyx3pDyNW39htO6tQa/lLgz4HgCgXIikMR
eahAEpoKoSgf7iu7Or8G5/tZVz82nvNmXW5HWFuocdFD1+nK5Y9HJVQFQPnmCWGt
Mvc3k6/f0J0/nOiT3AHIBHk+M7xk/m2vH8wD4DbnIoxM7vdsT1/ABT037623znsA
t68I7urk6Kbhxks3OPmHvSzumM1lKIywu2zii/Cs7dgp0udjgIBkDkgAdUuwzFn1
LVpUbCm7wM522+E85RN4+YEBghHqdU/DC3ii3jQuQ+iwNKO8KcdVgCrjsmGilwK2
emsdz+fP9n995Z/w+wDo800oNW1NZjr8PbMc7rIPWgErL5I9vUV0c1OBfG9Adqg2
VpTEXCf67o+Xl+0Zsl9MtGJpQTZFpzV7CGgqWr0wFRBz7669jWk9+NSNUfC80w9A
GO5+92Qb5/0VA/OWiRk8nN5mbFZqxxZ4p5kckNvvzNSzJYD7WMomvT+IIb/d6M9n
7UpkYuCEsNOo4ZacEPCeQLtb5BI7Kw28MsrTTgn4+rKrYbHLONBnS+tfFmRDtkml
5AECTeCvw0Gw6scsKDuo7p8NNI+XsxE3f2nALQQTCFWRAiYoXORrKo0jbLcWle/T
R/nx68GA8bHpO3WJmBgvlDIcX10MtzKrdktOItQx4JAU800JCnWkv7+YJ6DxTNIm
pTbvXhSeAKGMRr9itb3gdrS4fxzt4efDi1TgTbi3CEovPBrB+Vw2Pucx9I4CIdzj
QG2BGJowuSlu87VpsMXolb7F/5YTc7NaFQr71H6PK3i8DhAowuxl4Q5jkh70fmWS
cPTv7/PnlHxsuvsGa0hB6jxs3NKZL5qpnZtRXCT2Dx9nWsPdexVywUWgn6rRD//s
gwmCysUGzEqJ1N1pc2c2CrTUqRS5SWl//fKBgcptMIktLP5WIMd9erSC26F2IY3f
ub0DcImtG8b+fPVPQZ293mIiDPXsMWQE0pG0OYlpNfX9Bw7KfH6C1cf/Dx3K2o+s
B20QoaOk75SvllylLfawvWihwHFlJYCWEUu6ekuM8scJN24RMcWBwbuSnpR09HEQ
OmchcSRKbFzlWl6h78jx6JD40VOJ++HhbJn4DRby2w+4tXhz+fsneps26XjTUDh+
t8cngn4qc1Klt4zwheeFeTBJSp9UNU3wJV8aRI3y99N04+3/PfPQY/tkhFu1AoiV
yhk53aqpSsprIW0mGGZ61FUAuUv4IVwZp6kUyOTYzqc+y7gwYDP0wDPxn+3hTqHx
PQRJVYOquV+nAvu3X+5SdAQKGfXXNZC/jctbEgu+bWZdN5EnHdhp2EJaFtc6RiIl
fKwk++f3FvhVXHB4YS1yC0GRbNF1OuU8GKHvlPrb88qL9gTiKvutaNNcasGhJv+7
WKvOHpbTWxTUyN7dbDlqtCDG+P4yHa/KCeN6tNprkSazt7CQpxrTGusF9sqISikH
FKYuoB/Sx/usKKr6MXESCmU+2jsoQlL4ye1fu1JrUgxMCrYoc6v8hj0yuTyUEGuG
DeOGB6MQdwSRA9l311WMjP8sksO2YOByFu6OdWYU2zIZ5KsQtXRGPUSxEyJoAB4p
7tajdhOQZr4bUUqr+i+LdgdMwuG6uxc3j4ecPPpkrdDcnE1Qfx9pgys85ocIoH70
frZr6+lxbcdKuNgRR/D3+IbOYOZuCklShLHfG28W2pAwHpRWXmYhAOhuFKc1KfVj
QZbd5MChH3nKS74QR6F6Mks/g2zH0jGwBnkRIJtf9SNp+90BEarhSFXZt0u/xUMi
2ZlUBx1fg5eCrjzqY732NAMI+zUkAtSyRO6lUdx0n4j9hiaOVaW4klijTskw+U3f
Z/o1Fgj1wUDR3VDFGepqq0XlFmEtbPcuyiN2asWMDjjPAMyS2R/i/+E6YBRPSx29
wqPHauyyHA8z43NLnzFpMIuYfT++x+EEnm9RCbmSXNXgDgNBYDQgF62CMeVxVd1S
+AWQC1bEeFVuaWijKaIOrt+317D5owWRSlHY6doDqMGgg/m/4rqdr1LWuQMFGYCC
Awg5zp+fklTC7yXZjF2LWMXlDKxDiBCR2C1aWHThnEr6990nwLeD0PdRTHn1iYaw
WP33Cu4hmvP+f7E3fNe/UIl1jr/6qxt+FbGWm7JA9pzOjESltpdL0a0RPBb+iuwE
oZFbmWGhW6x9ogeNd9Xae+HrZts5Fz/fcYLf+xewVjCEoRS8B3iinabjjPyka+E1
upCsaLMgXGGFSEA4DKApmLaVSn8+x8FxEujcHD8lCheFJP5OwuHaGuIIERcl/PM9
jjjrigoQJVhhK3EsEw+KIhKOlJ7UQ5oIUvqGB5xA5LPUR2Hd1eXRwwekDC/3bZft
7nBSYhabfFprriSfUP4SFlDElGnrq877KygzffSu4q0+uI9y8eaC65jciHwRdVSZ
y6v81iLNYHzK38ozxrzU+BAZ8iLQlLzTjW3tBDb83v8FPEnKQ0sQ83lny21bMODD
E/7SI/mc/4DBINehbNE3fAJE1M4gxbJCGOO3FTc97qRFYR5gnU7HSD59Phngy9FL
d08l3Rn3VjmNS0cD9Qp0Tup9T430AIDU19s4abg63czCP0q9g6zyia4aYCx4kryM
43gr/GQ7z9XX/JAgG7My+w65EgedmQlEehYQgBfR8qANp7XTvyfWNURi5+ERCGTz
1k92Z5Xp9WcARBYNh2J9hmN1Wirq0neWMzX7fqeH7F0u0MH6/kh9m0Vnlw5Hs7Am
NrwJIedr8NMaZX2KOSf8thkOrD2Mx16jJI1TO8bQEinDN62tKp1qstUZCgr0rhuI
1cU0FXinSjLbH+kvyWIzt2hA+qKYmc47LRsGJc64wcbaNuZK4dynhBpRXgX5LciK
HaLsfDSaFTuG9b7zEyKlYJu/apGQ4hhtCN0/hH0fsgbUauFAVNO5u7FzcXghcn56
R0KyTNMNGVaFM4SqI/2qDK9nkaGuTAKr+GwCo6iGEelOnHFcjW7IRfgSwSDsuz1Z
0f7CFk+3q87GTteuhY9Pl2UKA+aaVLUeysWsgdwLepTJ1fyM1o6z+XGfUSrvNJEx
6On+5PqpTbFz2g4XhevySIKA/A8QEtKmqk0LohAA9QHPC75G3nwSMTdhzvY2gukv
DzlXZlI1Bi3Yr3/dapX87CykrcqgDn6LCD0f5jlBnyqnobIz4n5Mr3MT+xJQ8xnh
vjgI1w+6EvkZdhPFpYBXNi9nvxKTIgHnZJUgu3xU/38jcPgXxuhE1vwZQ4eTyjbT
6O/KFFPu2MH6i23jgtcCIpRXJVc8XUYvNA261uTVx9pV5M0OWCH8TdvzlkDEXRRm
26IZpuhKxtDRgJ9Hq1mDG9VqBtakHbJq3WryD4coCVIDONDFWdjZQRM3h8u8/TWf
Z2ba+8URccMtmrwdxtY3b2YC261mgpYV6/tEA3ZTvGOormptOvlefRPWy9kSbSkg
MRuPUg9fjEbA9mh+SdE7OizJ2zX/AcKOjD/WPluxEX1tE83HSw0eke1sRlId+CwU
tlsgdX3fkb5QmISia/el4VRQKrR5fFS2YPyuxQyMOot++CgZ6D4bdNIDUUs6ROEs
yfnB6WBit8mM3+oMBFlGP0eSKc2whoHpD1IzV/jUK1ZRNNS6wkaNmZRlLZPf9k+G
KNaUUlvDF54xKBjpYSJMmRpjQhOnoOf7XszzvgRlz5hodPj972QsFU1fbdOmHp0/
DlNj3wMQY1gJRQvTZZLbehHugicyX9xe0QouXIjAcVYEVIPkjquLv5rI+vSGjlVl
uOkvMeXoRRugaT3uNpLkIWBYvfQk+3faIDEf/o1gLLaqEnyjzjzBJdTXdgYpO+fk
qX4aWZA3fL9M5SyYbHh8TInA9uLKAclwYOBKfNNIgkuYydRwWUWc4p+xJdIsj77z
4CsTnCdChkIiqiU7w5AWN7aurMLRmi4uz6FcsInu6rWBcjcNDbA/8Q+N7VX6UoXo
TBlxZFHrP/PgHRRFWtEJ+0melpSyuTmNl5/fMK82D936jTu8weWaeguqgqTgB8SQ
kBEmH8HSefrDpRLxE4+RPOk0erBVAY+Ww3knFV3kyKzJp+smA3js26oALZNwC9VY
0YGe35Nu9Vi13HSDGtdMuyOTfLxSaTj5ur3qncxrv+KTWfA1m39gezJY+Uxyo1vs
/XmXQULxtTPyhDXfppxotWzAJ/sAHmnFHoLIhqMVpJM92toL1g9y/AUczIGb920z
kwX1Ta0NUdGt/OOoYAIp+rIKdn30mF3YeeFOFi1MIEallgJy9uu1klyDbtMDJOKw
b2R5HmIpzwVT2auVwpz7JRBLp9Cw5YOcTvyAzbj5HJriAKlbfGsxaUqx80PK3nxN
KYZVey45TMCEcr2seFL/uBc2vIhKZPn+NUBe/GCrkQb/2x7nZTULiDApWEjPHqHe
CJmtERtBeBi6kR6NSXyBJiQZtP70qAiqQx3w2n3vFcGLr4ttzT4xtV7WfDlQZbfK
P1nCfsKjerrysnRga3VTp7trx/+jnn47uM7bZVhE5nUxuRA52zIeVknYq1DZ1Dyn
j0HD/7wxGFv5O3ESOFFUsmMa7jIHwNF66G7DmnWUmt5DTg/JQ+9DLbGxxCkPDUeE
LcQz9WkpIXXiYwKqZLfkWFNOnOsBlBtntjytOmkYABT7eiWiQGrgCboAIkglCDkr
dlNgPPgbXIpxFQHcPDzsFUPxa6eiaJJzYMsadEnNYgB279FzLOjaXPAuOrKzP9ry
TlcoMsWN4rGUhD7vZW60UT79+2X0m38+8dBBe5Lrlu7oorSSx+8zleQQWVzKlxVw
vKMv1/KjbSDeQ4tv74g2VcjSkKRByENODv0T7StDHtHCH7+kaTTDCIWgBpGGghn4
VzUZG1yuvL+LE8OXPadDJZ3+qhARyqhZRt/Q105siBsigKB2aflyfzKntdCCkJkI
POkFRxp/ct/IH3sKIHtms1QGewtyhGtZCgk0gBJoaUG1yIinYDYiBsiWpSP8VCFi
t/LB9YZJ1RgNjTtqvdBMUCEghaA5TnJzUimK0/GqUwHQHfAbsr3UWb8Po+V+Bxpg
DWv/DxiSm7Ok2+0PGBuCnSQsGsj1Fr2G3/Yv9MjogPLJQ5l5wD7xkUQY7VVmNoCF
619yfbsrc/PmojCcUnPpvhr2eJTBsjlM/hxU3ZUjQKgdukJuGYDB9j4LM7eTSXRD
EmzJds9Baov7FYLlN7Ma7MOV2B+dFzUZGNPc4ExHHE2nszi4WgYsw+uvWLNou6F8
KCO16KKD102Olpj8mNoC6Z2LsUpIBiYTVX8NjUf84TkWXFhKJK4RXrWeAVFVu2MT
Ne97UCR0/g+woq+t2wbwbl+LGMiwE4o7uNOtcl2R/WHOODHa09Qi6JpPCBfkhzcl
3Go/gyrFVquKLVoAaWZf9pQJH/Kot7pMX8oO7VkmFeteiyY1b4EKtJtqHARriKxm
AILzquGiTdLWSeY9Lqv5NhnxUSZgGxv6Mtl5IZK7BKB9WCSRKenVHb5ELt4q8xVk
icBAZJbRA401F+/urQwooEJaFMz/n+7ZamA1KQ650lTFPHgJeW3WnKeGD5dlsO5b
/7f/Y4iUh03tcahiOEX1S+p8rLuAmwVt3IL7IK8G5+MmYM+gSNBkU9/QCg17bpLM
YsIDIltgUpCbrN5+sLJA1dD5dLsG73YTQOqeoXUZuM2/Oc7cIICB8Jc2qyzoLp0f
s/JAp72phj/Ntb+gal5ONywOPvMV8cXFJNGThhLYX6tMWtHXPujRgeMg3ltD+daz
kA9sia6qgjsiTDzxaVuzh2w9VZP7TaIpjTZ/8C8uYQ+hci/b/JyLkTm/kkqgvw7v
pXdiJmG5EUt5FkZBpOO885xOnGlUahMQO7o248EnYqqa42mK9O5oYHislJ4Nsk4x
Vxoy9IgcvNQFhIj5znSNjsizHLnF7vqOHhIzZ7vVjHyxJ+RIQ8VjjVnakLe0HCNd
roQb/zp6ltUF7PTH8ZlS8Y3GY5ZRBFnrxsic4y8rH1QOGpoEVYN++KCMVpEbIrmx
w5QBmumKJ5S3yX8AiK3xIGJCjBLozRVUa58IewVJSq0tawFem7nva+uq7iza1eLx
VWObSlQD9m1/SIgV0oNoCsAL970NEoTNJduYamJ32W62VqNY5JhuucGtTPRzJcqV
/GiXh3C9e+Q9SOmyyKrYvma+YsmNQmk2xL5SgVX8t/G45nxELiYBzaePXyW3s+Zj
1UHkWvYq+gATUoKgGUOCeGPrH7jQyS9wmwyg/k3zH1JynQqroUIAh/mmyJfk4A4G
r+41baBf9VXKzgFSgqIMLzQxbUuE6mQt1TvkwIYsa0hsSApxrtCTTMHaHdnRn1wx
rjwZx8Lcx2zKn53WCpgLLxe6O/y2YSJPElIeOY2SeOAdVB8+u5XAtK2P85ludZnm
PXRxjApVjwWmTSN3ibAZMm8QI8alUWv/sUSIZrlizd/rt0+okSghoVUUl16Ilb04
Va0fH5u4CdPRplfYAihB/CH5aGeZFzrRKWoD/o1N0MFmyt9rJ7QBA4OVzH6HGO4D
k1KMeFEjFloMJX3iwhYUo+QSoWyFXCzFZ5WQVGAGLBB/R2aqg0O8gv7VQZ3xW0Y5
N+tNc0vVHK1JvW6/Hst18vcKHDHEK9m+rjOjAKbXqDg/9FSDgmiBc1nXStqpMbzo
a/JvRU8RlVjYmXxogaNyiexFUqu/n4wzplNAbH578J5PqZVa0t8heAupWh96fwC1
tFTxHmeGMiOESUfGXsFN7HFLBG3TuYqxSNl1l6Yv6rbBfiLrF1TL/wwSWHUKrux+
/7i64thMWcBtrioldmjMDM7KfzmxrJ3QwxM5yJZOz8Ee3kz6g5ubV1fzeGHfADB0
MRtKYwc0V/wjJmJOeCKgGhgOD6PNDTorq90YykKMNzOqtBDOVoacvUXT9Sv5xEsG
axSK18SrB25nLFqlZXzkzULIS4p9o6R6klU8QPOSBk/qhCXV4nifXFtdO5Ncz+Us
L6V8Sh4idbe+m1jDPmh/reuBNKE0i+xaPN5lmSp5qE1zJw7TPbiZMGtjnKV35mhq
3JSNEkx9799DT/NyhYA17bo7beajGV+zxArrONZ0P3eh+b2vQR8XzApvBRUaXSdU
bvk9ME7iV9SemfjQsC2gqS9X9UKAjwr4LCwXDqRfFESPapjYcXSwfLf5Vrk4fjgG
cmb8JPrIZ2gF/UX4zOZS8lp8xBGoE0FslN5b3KOOJI23qn5qczYl2ovX4P11+Yx2
hq2Hai8E45FZgGedENwEbI54ZpS2cg5b0BcRtRgFyN63OhFS5Y0eQiS8G7SP19cj
mE4lZKk2IPtmpTsPO/C6/ND9hF6YoDM5wJ/hD9OSlTzgzQWSBHSJpeCl0w8QLfOv
LOrj7hm5syeHMvBgVpSeSZmM6+IZg6M2E6YlVn6Y3pyEdiKN3y36EwRtrqpXRG3r
KIgZgFWSuRXwQJgR5XLX8jOt8gUzdkaMLMcgzMOxG8oEHqfXPAOVCG/Wg9mjP84v
Ym4SVhEBxIEYISLcPhp2B4AbWzjgBVGd1zAJnH7r9gvBN6ZkkN2vQyXEx233UXSU
e88fJ71Ly5Eg+FjpRFZDp0NDJGVB0tGt6lDQZKgKg8XLK/6QokqJOr9ppO06ieug
xf2ob3BcQvGh+iawgru0xvDGydXaBq3/gIrmdrV9iN5gGlJm/6ED1GaufgvTPUSH
qSEBdhaapkKM+LgqyRtC1L8tk2BVed6V54XrYdBUim9T8AeLhaMSCLN99dgOY4Bz
ibtNWKEMbr3NDzAxDFedSsr3quj2XHh3mrG1QeW/G5SyoEDyLeaNg6CPgttX4K6Q
+1/2qHyTFph/pP60WAb38n8BHA2SN+N+yqD1p1BE9vMXJFZ7JxoW52EyTaj5gO4i
ouvs3Q2Onu+O9PFQ27+QFPqWdjQazIBP/kTymSwU5h/yvBJ27MlIS2+/YKecC+Yi
H2yHvCIEVXsr6LbU2FL/zr1YhSnZeV6ruSnWQGjShnSAPmz0r2UYf3vHgyvrUn2m
xUkFEoKzypwXHr53jm2aiZxP11cRW3B1BjtESb10BUeRGNuv/acdhCB4AUXqmBDI
ra+dEBrV86qVUf40+rgcj9bz1sKphB1lFHMxMv7ZSIC4icaOf1iEUIwvkpmrIps6
Ox7MNy9cegOZuWIu7c84E07oBToTcuWNbihdPTljrwYxAcPGmLeEAdXHKHyfXL1D
qBBZZE6jGY4TAVE4ZUwCUJ8sqW4KRzs5fhhsEtmKsCEzK/4ldNeXI587Z+4BgM5v
bsHM5FKLZVUFmPtLxSSa8bvu1ANTHoROk5wFzaFokQbuwL+yWn8AWnxyoBxDnSZX
MKlg/OD0Wkjo4bRzlWaJT4asLGfR7Ib8nx4semCXObhPn+bULnR8+Ze5SJfD99yz
aVOz9obO7/1aS9wjwqaVHnW7tYBhYJiV5Go8Ad3j8/ZEPbg9Ld1UCZ6dUxoGFaiu
lv9rpw12ON9/SmoGnhgRLFThnpnd2TTYrnCIGlSVD+aOI6wg/x72nJJ+Zm+DIIdf
3j3Zz/LA5cdXFD/8bKZsNl03CjOrzS//kx09Pzd0YW7zbC7ft5sjFY4k96gyKNy3
/uzK1p8HrIpfZhvuXm3JnqnlOXXQbIyZNw+3DxrXQW8+aKwBHb33Asb3Q4RH40dg
MNXVetVqI6fL6Nb1p7cotOXhNipVTCYEeaqoCEMhUVHOcPykZSGKbH4rmoQO+mlU
MqTqBlcKLuh4TX1O4CB62K1vQ2VI3hFU5zb0NFfesLTj/PztfZcQERpPlqqqvbDp
HhO/eRLdj39yMsr/3C+owMoNRYt0JgBZnUUA9wevVeXwVkQbjJiex4eXQzZK9fCU
aop6WmBB8hmtA4ItONS53GLxnH5LvjoqhxneuPT/sZONNDS+6gBeLp2ySt3udtXC
eavIN2v3uVUXhMmpbzy+Y5F4WaQs1sXzWYWPTSRXK+4W/fgo8lw4gR58FdpBpuNp
TrVQtMJObW0Hlz/O9z+Crx9IVlou19crIzOXRPLXJg1zPXBU06k+G/aVq393Wa/7
GG1Ug50Q3SSWmdfM9iCeMZPwdfD/YvQwpGegbKIJENFwcEfarJUnKV7OfYIAnjiJ
lQM1kAwpHVQYuZ9E1Q+RR+qDf8j5ewXbHEpjK7T17J8+GH5ZUe31i/sCMhJfmin7
WJzFYjL4AlR/5z9A2ZAokRN8n9whRL+stAPQX+gLdLLPKdeLx+RChA74exGtV/me
SgAr4POFvPOcD2L3jNsQCbbacjV5eOGkNr5753c246p8enZaZWJKlKJsnxdf++Ee
MAwY8DUmz72O8ureo2Aa8yCpv7Gi4nsZ6EVwTmp+cNoWYGDPK8qsz/F5nJxwMILf
mlX4gccLICeVYk7H/O1+3e/20UiLn0MMAjKZMqehPJ2RYM3g1yjfZPJWE0vwAm1E
+eqUpUSBu3SzcPTKF5t1qeWXY6FvGBKSaynggJo2wPgrw3tZfk8BBLGw3qQGHf/Q
ZvkzhGzAXRBsAWJYdh1I1N6a2SrCz/aHpFdKAxtdiHTSEW2xtisPhepzQHzucFr/
3VOuKbXF9CZnAw65FAeAyMtZnK+6zP3+Q9Npt7KI0KDUIh33OEGMgpaV6prs+mll
La2RxVfe9i0O52ACO99YLmvY3FRhYRWPlqHuMW5X8dIZDZjUP91uaTh0MoU5kcAq
Z/X+0DFahoPbVwf+2HX0LnCjP3xRhf2Hifr+Tx7CMr/b4CEe/gtZIiMRwRAPgvdQ
jRDhxPzp0xxva4117gHgtmk6HpYt7w25xh+asdJY5Gv9fM50pmBRjk/5K6pDsjQ9
J56DELlPZMTky12vnlXD56jzubsvHXCOvPRZRmrYh3kTa/PGmfHBqr8I0L6aTwNf
N8ERNYpNW2NMGuDIwoiNUxIC8mpgxbtSELV/Ru3z0Z7gT0VXyBr8Nk3XLSbXW+4U
ybDVdTjdc9ar57jXQVjOLJondP9T0vFAhJpHAE6eTUOjD9fEI3Rgt3YaL+Ofk7Sv
GSlSXkZ7aTwTk9o0ZnIkjjVgqCvYKsWbmZtaDCIXMrSISVYZo/MlxJdVgf6deifO
GRdrR/RBy8qbVVJkI5l5UZ+J+Kp3IWRklAPJv5Uu3TaKlpUWsnPR4W/7SqvhL30Y
itJ4I3Rn2ow80rNfVMlHZVRY+f24FUYOOoGZLmUlRWfIiNoqdgCSQfjuBUSMqLCq
TU7FhNUogjM+rB9t9yAglepIfp8XtzmJKVas1ozDnePgsIzAemyusOJl5lOA2GMa
70cPQvJYHabUagXidA4cCaq3I+y/WzHURR+HJ/9V3YfEUCrjoHrOTPAzsX6lHPYM
RcqnJyDtN2WuQQlhDAMGNqF3YnU8MUAmLHRmTSMslCltjykl2AW1s43pIcf79geg
GojmQ5upNxjgJjbm3skHdFlpl5s6cudRtr/CWGvbZlAuJuo/hD1Dc4N0gjQKJw48
dQcWkkNNVP5sMJIbM6g1KqW7kpgl9tAW5n0iKxmndRTdGyKmpX+xFauNb7XffjP/
MtuS/of3uOP6FUSPRrPieSJMDYoxVtyU+jBJnZ6Vgi0zl/lpRsUmm1yJEtyC/VDA
EdiczEL82G/RLHmWEYEn41KLip1JZ2Ar9YZJVjqsuJ3z3Kln9fpVd6cbA+va88BM
bp4Efs4sIw05vrhPhYRXQATJhsYMyJ4jbkMJ12CKYNw4nMguRTJNhpMfJjNh+WAo
6ffbb+Pg0vfZOnhPvWePdJ3g7dGzpatuKM0uP7D8EZ9xujC8nHrnO9Hent7I1X3S
jeCOB/NIFOwvbwrtRijYx7RpUCcsFU1zQmIL455BncZ+IO/QF5n350rcZhTaJShl
fJ/PmMpfG7z5pZTnBLsOQtkmfymkiW0jzHP/bOMTHcKfDLakdneiBc69D7VR6rDw
n0uS6OVnTwiJoVOEVNJYP+2U6/CYQjqvz3sItSTJn2X7Bdmnh7/gwYxuNuHnQwyA
bGGdAsZ2nnyclWzbuh3wRvnlMAJ7TO772WXo7Zl4s9S40nhYh7wHDZCA2twe+n7T
6JLCWV8lIjyrxv3pJ6t7cousI8Mtf9J7o9AQV4ujSwlT5XwqktbsnHZtYZlDSpwj
U0ICDOoyOa23XYMMwbQowDrnpW13aDG1e3AcglgPxjCO9kzsVgZan++prnmd3YNQ
eQKZ6B7FCcCnznbIFJsU/YHDgBNGQxKygNVvOrbYUcxNjU4HuDqaldP7omepJy84
+sAO+eQbughiwQdb9DpYVTPTyxpHCvbAw1rBTV4Egi1dsSBiYib4yjm6NN2T8qid
iQAmXm4gUtFvh/7lXx0HWiGaZ1d38vchpQC/wqCVUapgo8NbzCeVf6r9jFZ5+IXy
X6QhK1fkLx3zPK/xr5Y/fEUcNljpqGvrWsk/b35Ce1glzcy/3oyjussBTIhO7zIO
wlP2TwFodrq22wb+8WJSSYM96bKGnSvF36rNEAABSUOaY6y3eb6yTtg/D8nUwsnq
530vp32SLZQ+TEpFaxl0IBjMKcbi8vasqcq5IXAgvNYPWaxyc9KuexhNYP+R/Wdq
J62q8+hVJqlgk/8m4F3DlqdSznutNppjA4iw4nqwKJsmU8fAtnfrubCNhlu/TYaQ
7po5J4tnwTxnU4Nx/a/UDRW1MP+Cp1o/Jbnou9X7w8HQ+q2clPr0UB5+l2Wk0iov
m2rBXh8wAw7+dHxtp5oEKaVLgt4qS6cGnAQYbKCRc4t0+1Ky2yrqU2btz3Yg6k6R
XYn4S3hnH77LLsnd017+zysl+kK/BGKXb845F1m0/GWsQsbCS7X1rsdOEHjFD+0K
OjJZsHhjTSA7QqYsAaARBydY4LZzjK6/nHojXG8HgwYGG8Khre9URinZZH0OquEd
Xy0AHZxwhxfD53/2EG5ruc9aiznafOLOWNlSubBHGhr+eSTPLY8xUo4MW/JE7+U7
AqOmB+0N8fNpjA1DU0jHl8zvfaqxaSBsHVKOfrWCGio0HxZ+cGKXINo4vbP5pGYU
41Fd71lky3+Qh65AqHlwNsilKimup9//rcF9VYZaAnG07g5/QbElVAA9bvpCuqFA
oybtCRUXI/SWESLEI+P8clfodp4bxw0h8kpIPvBYmeUm0f6yrgDFjzc1ZoaFfGLA
967zITg44Z9F9Nu/CXb3lmNXr4C0qAsKCK+dAMiwwbKShcVFaJhgBvTxdHXBuWkR
XhQkJS61Ktsn2+0h6uZhAkiXMOvLWgASYcPdsLbpcXRwmcq/djVxq6CV8sFq9L5h
q+sqB6RroLBFymtqgscfI9c3TFIr9yoaU3Oxxwn617UR3VLIk0daT4pfJf2aG5sT
H5WlC/eJHQ231YEroA/W9lCZtUDwJH13rA6lP5FA2r/UAThFCQZvjrl/NAUuBzKL
CCH300lAcSGYuc3OHSo7Brj6K0dw3kZiHeMrncO4KRk/1ukiRrfA9gm9bGYVI7Xg
72a+qgpJGi126D3W2s/O3CZZQK2tNa3ZS0j5SJ/YX8sCNJ5qh3a2Mzt81r5iIWK4
KxTLtEl1MszrZiRtqSGvjh/FLXr7a9+tC4qVZNs+uM8/1Ciz2zRedf5pGC2Vq0As
FLpeyPAg814Ins5aCdODqF++ghMB5Bt29hPY/6Gihandf45Vn2R2BYakNn0xZ5bB
TyjhisExtas3MeFDrEEgafe6Y+YS3AHYYsi7xaX1ZpP+sfqerHsHghB8ncengxIi
TUvPhyVMb3wRvLvJXLaQL8aIPNTnTj6bJnzcf3+XEgUhOASzIo9SrWZKAuBcnQY9
eHPcZGiZ8XOQ10jxWuvhxBcZ2Ob7Dks+vABB+meIDR3+x61VtPEOe9XAoF4IMGdz
/AwkrWtuwCl5Dx1zKRnDLBBO+AdY7ReyyHMhzs3c3RtsyJiRMADPozUaN3EAsA80
wbRGVdC18uY85ARUKFHZzInhKR86IKBnwaqHEuUVpPEYaSizqxxh4vmhHtF2JVed
lQiVagUPglSHasDmTq098FIhAsT9Bhcu9c0kwi6LmfCWEz3nYaTsvI4GR+hrlA6R
lja3/2LotH/31byVaDFfTt238ZjuZ0FlfOk5Xyyoojvhac7Tvn9feph7uR7Qx3az
9xgcClwXoAamZ9hWFj54/MawD3st7I+1ewYb3PTLI/f7lRZxKJHt4KScCaW+ht2r
X2c0tO2zqwEBZSqovn8C8gVW3CwDE3vEAq0RigWzk2pFy9jdxIXkkQc4TfwHmVGv
hZTd/DE5CQUjse9maRR9WllhVdExqG6fwiklw9L4JitjdEM8NY17xXjFonuEtUzF
6cHxz0Y3pMhIjO4lLl/qyyINJjkf35onD5BbCoaWsXIqiUyrdtVBYz1vA/o7UsBL
wB0itKASpC3Hh2KrS51S6efjkg8tPK62mQCi8vwevOKadMJaY1W5myyxI7sQjicG
ClCpfrRzas4bDLKZxd4Avqh3tn30Sb/xOpLcso7BTbc+3WfjpIa/ifBrcn/oT8gc
pPi5bAU8kFvpgw8tC+AyhvJXoqNbXqUh39pp3Ig5rMd33hSuiqXFspxJsXi+v3ks
iISD1QmNT5LeRFE3/3kQwZ2uG9ugF42DDV5CFLh4PEiiRCg7nD/1pLwcf9Yhr95x
wrdku2RG8u15jx1SlgnZh78C8Us2YHaVTIEjKtwFQqvQLRToYKdvbWfDGKhSKGoX
hKoNuQeayJGT824nzK+BLmTVffbzOJOmVaAwxgJpwRupTnQW4keqxus5bVZBfmgW
3+ZMbMghm9Kr/k04A5+qbHkvl3YCpPgPCPnlmE7HWAWrUiSqqej06dhRKvLmZZHl
XLBhz/M08EwKFctewSelY+9zR+6VOPZRNtLuIhTetAfwtFPND1CDIEet0P87sL7E
DlDiVLFBGM0uCdYeBdWoc47s570FAh9kaWMJkp3pA1MBJEVaIGbaeWRLIrKdkG0p
lsRZmY6x/V3JN4IxQrk31MjZU7qB5tt3i+RDZf6mz9cCSYaSg/dAS65Wr61cHBxi
jTQ8nNi23p4xZ2n2QMu818PwIU71b7h4edsiYIj5RPCcH1b/8M8N1fnaUZ9JdfXI
p/l4yo0077qt4JShk9fhQsl+fVI19HXwBnCku9LPP0MrabX+5gsT137wZYvaV+YF
Mc6XeWVOT9dADUHH29SvveVjR7RzjuD0C1M6pHL9SsY4tP2+CFELVeClekHOpmR4
V56pazxoN0jPru1EiP0m9FNmYJjAXKKqcufr/gFYb0xlG71+a54xZkzJ/IS/2G3c
DjcPoE8/C5N4UnURm5FM8lol6O2MRY7KAv0mLKBQrSnrSY+uk1P4v8e4dwozzNzq
ORWMMJDTddCkGdz5OpZBjZqLF9KYzRa7+NIgHUfOtBeH2DoexajVP/hRVhhMTwYj
YR1tcUo7SY8KK2cXW7w5eYgxUxcvk8k8rRT05FIrfXxDCDmZvhORd97eF9B/Vg7t
dSqXAOsjQw6hOpyyZuSYOf+izLLPZTVgF0yeK3VKbFexn8eQ/BAsUuZ2CINQCcro
lk94KxepQj8sEWOE5ZLoqZ2S1KhtZX4DPPE2bRVRNHcDcmAgjR0ajXg/zz5Wi8ch
GYJrC6sQKTLPnlXInqjiD/Bcm2JZpm6c9UFBf15n9F+2exTg4GBqWTb4mSywcIVS
VIjT1vhxVtmaRhG9YJcBSwQvNeYMTqdSYo5bACFxj8IUzlXXWr/nvKyGdNutxYpl
4tbiSN6RMyAM1+F5Y+IyAYjKoLkTKJxu/QRgWVJPxC7S4OH86dZTvv/8asdvK+y2
KNokUdH+AikzgcUY57NSB0UVBra2PmK4KsOb2dcHQYiFjMttEo2IzTAw0fOFzCG5
Vt894ipbR/coAYhxGYFxGqb1k2Rp4fy3/QB241LT7Oin/sx5Ldw6noTmL8S9kEbS
hUn5hug/WIuXmDLO4pz1aV5gzceLTVRMbRRGCcsDLjVC/7sA1JNvaeiPmETvG8hh
DQW/hYLmQUululvu2/IsI8QQMzPptPG/GV1J/0f+ElrYE+G/JzwL8aNcBWCf/FyM
DDTt3/rw4Qi7Q9OYHdqH3aG7vjqmQ3gavNsTBBe74psi/M74e+kG8ml5kNxdQU2D
0U+aWVfGuvtiguQ4RrmdOs6KZX149MczUKWlfRpGaGPdrSLhb4Ib9jsip4KRZyX3
QskC2xRCfpw6l1Q8ngebaewd0UeJUQ4WRX4I0YtftbW0ZobGVWwwGZx1p7pxcc8g
wZckkNfmKORzIdc92mb6gJD6wp6yspkl+WJG63dAmUa/ErZrGVSmlwwHrbIYoTc8
AiaEZ1erQxNrIe6OD1+lx2Y1namst3mGjIvvGeV9xbyeUDZ6Wy/x5WlAIQd847ns
JmtEPnvGL4PeiIesnBTnyR6KhNi+wSd3roUWsyAIbQDKgBVhTrZqrflK55sKQYcm
/5uMn48bBtqDzwb4xqdpYqouOAmYh9LblmOGBHTNy78OfAOLUM1giH1rg24e+Efg
+I4mTiCzsgIh8Qm/wIXGpaL57Pbn+ofa716n1ijiTfRChAuRkf5h+5z56/0CN9am
+Qt53iTa5OtmtPg9kl1XVrp5QBLFaKyp7i9w5531CopwaiGPncHb4rb2Ki/XJ2St
Fpo5cTbuynsKnEiUme6xM3wWYiTcHrdwL6o+049vwQ/j1a2UNHqW814e/6FW/y3Y
wMOLIpD3MbNQAcA7uZ2lYPnIhxFQAq/xrxJwZSlVPUVwgae3mzdG5KIbdidQy+tO
m7bTXr0wQhWBerstQ4SDLuOrq3vN0EV4uMtQpvBVfgghs6vTZPgGFV7Keu46bVKg
A5cShESUyeg0SExvu1UiYfw7q2Te12uvui0CUtqecZgauagq8pXgczUC2qoTeuOU
dmSDFzVRnt5QJitU7zSC4ROo+yRuJDMo1DqkGp1xisH/GxfzfiLQ8Dbs1jsKGC/C
5T77XMFY3SXni6dvAgEwMTN6e/jbgNGHMpwPwTGOF685ffECSh3G9vxO9k+v+nLw
G/QLaS1525mXTjAHPN56SQ5rP747nWxcGmljMw4UTYaTR0RJITA2Oh3NbBko9WO9
uYur/WD0UizOyCYG6dLLyf+qmiLFRtEz1i/tGkEddo72qF2DiMjDBvQSBBj8OIdJ
MAVmedo7FUvTsqwZLKNC+g9Hnvqs0L5Xx4eERmKddogViq0pvBfBFIDCAyxPxMOG
jjCDazT/vp088e6+wtiv2at7pT62Syks0egH+lfhYF2U9yEDVhGS7l04MxeFbs+q
HcAHkbN39fbnHEZRPkCOdOGd+rFNvr1ruOBUfUntzKyqgGKuk0u3ShGOIaYxYZn2
bSicFBxBrQuBa5MQay5lbUgtp5LjRVzQFSrAjOs/sa5A5kLZHWBX7znXo7kRdOyL
FaDPHtiNGYwWCYW8DHjFJkpiPHpyxzRGJ3Ww0uOu99eN8x/pkjp4v5o2Y0hYF6Qw
2FARk+K4Uf0LToBTJ8O0MCiuybWCyEBtcinjI6+5uiKdUD4d5DlXjK+g0ELWTRCW
HZgF+cW4ryycgBFIVZ+ASCdYdHZSxPmLQ5FZ/dN7IF+N9vE56IboHZiIa5hMpYub
aj1uC/PiIoDyDTY65kdG5tcooTT0cdHAjxEJojVBFzNo7HHMHE5kZeu1+QHlsnSG
zTvql5oN7p8o/7Z+jBiXmAgMEvUzusO74asH3Nqp+yNNt/xv+tGcvOKuIij0imEr
r6+bTcVklunZBWusnD7L4p5R8eKM2ofhGcXqQk095fVHrbTqPzoR8+FhFoC3Fn2B
FdbNvJz2pKTmt225tZVw6GU7lHNr7twgD4s8e6EPiDb/Ql6NjL83DQEV3kX/2VJF
2WdgzVwq1zurmJKTvpGwMBx7KnYKylvGGZjguD8ynti+/zFif2aA3JUsGQn10J/B
0G2AtW4oIUB+x2OBjGaatT+6Wn8v0/zqmuI5EXp6hgcDuxxPdWNENaBm5NMCHnuu
4m2duaCISSOm/fFg5samO5+KAVJRBui3RpSJi6+k96NaAYh5GfNF32O2s5zDW0Sn
V3sKskqymA6GrlktqKecK30MgVxeLrnU9JMJeaL5BICfg4VOT9nI/3lZWxQGMpgp
j82W/bwl6JKLCMtmDIt9pQEZXQVgkSKAaBuNRD6/wLHxtcmAInzLm8+zwsaGb4qw
qvI4VBIo2ySqZSMj/GQh7xYeLRblsJa8WRurBTBUw0w+Qda5dN1D/KLVWJDBIVkv
bv6e0OXOnZHuZMoBa3mul18wWzRGOopo/lnauDVg8hUBuiwBRVOZaNRneJZPUvYS
DDA1TALriWxGpmIeLN4FwGnLk0/IpU49SHybdsYeSILRbGY1RJFNCrwc4l2db247
elZMwtRL2wnMANtXoqLPlj4qLq3kMJd9CVnM6IW/Pm74vLU3bWY736k9y+QrsJ9T
vLnnQ56xMryAE4wPArsniQMXeJY//RA5FmC21NZX40tDDM5jncVyHSg00amc210H
qkBEoxrklgHwQVXl5FSVtzi3gDrXMOSJQHjkrZTxWWV1CSLr3RITfXaqaGPz57MI
56R1QSQEUmjQRnalADDWSj3akAzNWklR3uIdIAUQYGazcbes7s4rhxWSdJn/JKQl
ktvlO8X/9/mXMco/LGajU1UfbdJZvBD1Bo/Zf+FYEVFLPGyUy+H51rjbaowVyDnZ
cX+n97JTTTUdyLg05NDnCB5FXEdUdCNHCjOyk8cQM2kue8yj8zGsMKFpOb9EWITR
bmXS1qE6NggQcQlUmM2YWM2q2Xo4gP3TM9m1wFnb0DbXrKxwGZBPFodfZXt0NCCc
VnKGwvu+QdS069mpgrtBJn/MhKax0lIgUfcxFr2cxExeptkv+CJPaYEWnZ7VmX6l
9fCbyZUGomiGkhH0p4Jr40U0uSAcGMEUWSrLAVw210zeeg4+e9ovvf1M5fk88e0Z
pYhkOX+l/8phXygsUklT2wW3eybT5KjVNcry/wTvDhFkv23mDbRc91haJVZpVSPE
Q3ZPOPZZ7qOyFfZAGl4+T/W4rf4HmTNpX3ALwm6SdR7gBNMS10wN80o1jsEVaW3w
nZje16IBjiBbaTQ8aKGnJlg4bQP/bOKlIE++1qC6E73plWq7ae1znKDgErwv4GIy
etBISWVt7phmjY5E6RGD6uA/NBOmcGRLsMBc9RBOpzHoGMdB+lVIuAMwvCqz4bot
C2OVD6a47X5NYSzos1i+/EJ7j/o2g+luNjEYZjT51uY3eE0eJ7r/HkDG6gbyGsxy
5zwuvN9H1Okgnug842E0wgADs0vctzQyumZFjZT5L3gG1GONTv1jvFA9WTo2tpcg
sHVdjFI2eiGs3M91EeJjLV7y/D6Haf+sTUT3icn68vO02f7sVB4z2I6IwNaxDOcU
QNutZq2WXe8WRH00Jvill1RG4vtETRImC/30626Sfh69V4Eor/55rz06kyuygDXg
5wyM4zu5SDoAPrAWFnftNiOH56AZSiTh+6zHZEhmGBEzN8tubPAj8pJXpjiD+/tX
9Hzb+UrwL3JM78Zmg+WAw5bTv5GhqrzC/qMEnMEgWNxPsMgjiDwTviSTalB0FZHG
gkMw5HpMZFA6gYhhEnkg43fyQPoCoTkFLpDe1mDuYOjM6jWXvFswtFCTmBxjWfuY
+ysVtRmYdFNUUq7yEvK9Xjv2J2PHoPAoLJqTs979woK5c+aTtI2BL6pwBhGa1U7X
Y5xFitv/Qh1niVdH2Byv6aSlIhWWUu5IAHbJHZnJPToxQzpma77w49RKf/0ekYLn
nt0b0+NobcG72Wd4jPEaQxWH59KbivjCCKbPc9Yftaw0Ap96+nSqUs/3BqeBeN78
i5J+8oTVmLt0il82oMnqO/q4fMt7S775jMi3P9JAbqcgx6DkxkLfR/c3VFpW7v3b
JcZqwuxflypEHW9QgyiMufC3tIxVdvGllG6dHwEEwdCg3MQxs/xypxNM9ls8TewK
Teh5WefiPiEmoplwUDSz9ILImHLBKSeTj8ba1nGQTu8bZ2Wc7ekyCRJusnLgQ4Ll
Ji943QP0PwCwZueCIXEUzSLbq9EML/AKgtrwJTT6Jl6mN011cjP2F06ZUgqEnV4s
EofQEFjcEjtNtCa4N8koHvB1R+gRUiGMs1RKeqpnw/53HjZtlnowtgcteNmwt0f4
bxaEpuEgBxTbqQtq7kRJRUPv1dfQcGNyTNYLdfY2iPT6GHxrg8ByazDIiUpHAD6T
YY1j9bqQ9nLR+VxVWjnmtQ/WSPsiEejtXLyGMa/d8bDIoSdmLLYszkXFxdZ8/Dl5
9YNb8h8JhxGC4q8O8ofNoze6q77LZKc40+ZpWtdhR1JBDnSlGPZF/TMYM8eNyd+c
6fhg9x/Dz5KR4XLJNjdu4QBSIfJNHXde7T/AKUVwXwXqe263X/EkYWpyke4NmYB7
gy9ts43OGgcWVJqAsSJ9i7STmZBblLYsnzzwW4qhkJji12bjkcmAVKK5bidAWF+5
UwQeFdGfPw5IudLOIup7geUoFbKfnDJwx1qA727qEPaqjVeJzXHiW97JKOzOMN56
1IZH1nyUHyyBG/rTuRQHOSzvU2KfWVzznEEYwbdJ3CJgC6xd+ldPufn0J+cN1wEO
AFS4B37KJ9qKTelRYdTQ6u9zDNziOLVvUc1K0O0Mvs0GaptvSrSpaKAaKQ7bwrzn
5ihNMQQasQ5vARxYiSX/2RzgCvez9fU7+m5yB54t+8RO6lZhSoWVwVTI0iqltj2w
hTy1PmybgPCO1jLRN6u1WWB0Q/JYLDXRHoPzX4nERdH3ABbQkBszRvU7rsyg6ae/
6O0ok7hEdYOsm4P5D3sZPhppVlqkkfo6gcw7fBa/U8OMElh5bpwUO4wEmMgctyco
3aPhfsYfQdmF3tiC/LSEvIc5PgsYnG808DJHKYbdTSf9ZEQ51n3XFDYW4ZjoVzHF
rYE/dkXafDnGeszuYmFRrwP1S42HzC8omDAHR9/SZjHOHpgbz1/U0cZ39EZ0pZQg
PqxuiZHAQtt3fy0eetMwtPenMm8Rn+uf+4rr8fDGrdPvIDx9dgq3xOUCpdCv4Zev
w4893BQSvU64NWwojhx1w83F4ryha+S6nt4bG2yHAhIzOFRMHHhkWWaPlishyoWh
4S6r4PwPx0ry6RwIfeWYke85NVCVSNxV2iz6vfqNboUTWcVoBuv3HswPSxBb87H6
6w3wZtVeW1cHgWtgByuRj+dG6oMHpeWOCdXAphoMKfypbXP10pJZnqLxuhQ/Wp99
Hsz95lXuwSEfDmSCjjHdauYQSmphGOOjJcVRpOvyE+zdSqMa/1UXPOAuF/22mvID
PczbxBoOFHGL9xcwOvzxEq47BwEQNDcIjrY/Pi8tHhnB8Xu5XgbQIrE524SCmJEu
jm1GshwvJpOd3wXh0GbqYYYchAvHklI2vksTW77mIRrukeGfLSnwMCi9NRuKa35a
lowwUmZrF/j0d6t5Mfx6p8ig9A1JhQkqjVY6rRAtfMG9SCFJTO1aLNA671AGqWuL
MUtLXLr/f1PUlJAgX8BkQvhUuHb5r4cWf9KwjFiL7W/UBE6/QNz9jABvGznNiRAh
vpUKBRmM60brOQiP5ltVsM6R0AwQNjMl2FyHhD/UY9BEshfbGjcrLgXlydAXUaky
zKlrdMbD2ZbRN48aRvPMP28yrBNZ/SVGRRyETzajI2OxqjYMOSOiAlQm+RIC9pam
53J9vnpqNrQchvFh8OZ28RpIB20sHk1CyEXgSk8ZUpqf27lMx3a/QTYVrO759e/j
s/CAiJQ/DiYSuc3goH9tcNtserG04EG++RT6oQksXGVsmV6thGoKEM9CDhVXI0ZW
dDI+IYPoaKyDosLs1laE0/cxouX143J5H35PuDIRm/abdeY9YXcOefAF9L001A9e
MU7BuEopKLyCYFaDX0HiG7+hKRcv5gW3AavjVAOUAYQaxiD2NlVcJOFeuAbvbxrJ
3TimcKriVHPp/dl4WKCRLa/H67mI5haJzdkPW5d24h4gJ1KGGXRrALvx6+MZF94B
zEmc2qylJNJf0Sesq0wjp0rRuAxOlo7sDNlI0UKCEuDZVCemty5HsynGeglzPEXj
yluFg79kMhdFIrcAiOOVtqLBJ0IcVTdDPHfhJUwKMV6bULd2DJSNl25BEAVIDGnW
zrTjqM7OjHSwWMuVAivXok+faq6JAUs395DojLuljOcOJjCZXyxHq6LMYWW0HyAN
xSEWaul/doQxyYky8GAimtEzIgkboKnUBwOirtUOd89qoYzTu+4fiS7pfY9p9vTi
yWfkUIcQTVcpBECxiLZ1qLLVrkVniMcLV1k4Zv9jyvcymxWm5PcZUoNi2/Ydb6k6
3XWn4woRxfLDMX1yTAG3Dn9+avNjF2XqngExuZPDRL407Wa3EbEsdw2U/b4K7IzJ
pPOhS059nhMEbUA27OXJfg2kg4p3nCnBj6EuRpFSmiy9qe7DGJVIcDt458+CwnxT
FiHwXfgvrC3+fnu8FF08WEQ7BK+rTvZnc0CCj+SHp+RWS5erpYXe/vjmLi2KbgH+
Wvj+WW9Z+QAltYJacUpqfLtf9wZD19pYbdwIAifnbVXFxRFkAf0l4N+v3ZWGuHuc
LmH1dyZv8oITbtCtJiqATjmrZ0VAgc+/wxCBjqav3yj5lhykjDfMom774YR5Ybo0
+RhDgxb7FNG8n2QBt0u4CshGi+gE2DwwyKZQRQg9v4HdQbpDdlRxDhbLrmCdu+4P
GfLdMC59qE6sDUv0txjaZgJfUsAZ0h/3GiJ9S0r8NfNKdv/tNctwYyYDHRjRjIGA
eejFqWfdT/evnjzoXMcxtxADOgbDvVW+FpLckrrQaf6rcHgpWswee4zsTBTnr7Bp
hFXzaZjXzR5xzDyHnZH6XgLF6A7Mu+BdX9uu0CUogFW+XROIbEstXfqYvgaZaOoR
7yVUKlnr5x0CniSi4vUzBXOOBRYE/yQ08icvUMZ5DP/LEq+y19JhnBw2xmRXsDCg
fHnA/WTgmv7Bjw4mY2/EI3nsOPHpDsvLtLzlbfsIsijlmcQMzkSQX7aG6bkOpKFJ
qs6xE8jwa33TaZNpaBSIncRlkmsOaDu6cNjY97TxoL9mZzYGUR6y7AC0D0uo99yX
TyhjlgDU6z7gb15ASrJB20I2EdZc5f4jBIFQqI7Ah8cNJ8dMdQFMFpcadF1mza0y
yRW8RtSYbFOomke3FsTnsCwySP3avLm6xfWuVpd0z099n8YIkO8BZGMDwC9LcnAP
LXXes8Pn3fdu1RYzCbB1/2y/SGRJ26K6ZO6Oyk5JCuMgu4/FcV0e8xlXi4lAj13P
mmOuPJSAGT10HlefjZriJV9ZuOZW0p4jGPjW2fsDsm9PyugA1p2m25yuLM5cKO/y
K7FF7010bRzb/KwB8qxCNu//9Zr6nVfsGAV9Ga01oy7NfsA3D+En3YkacALnTJj9
zQUEAxtCXXS/DyxxjqYujdi8oa3e1jUZJ3TPgovg2TofCpTEbzbgbFHF3RVEiciC
ZqQSGvI1p096cA/zuLn+fjKkNIbjfAh1dxkzF+8TK9gKgTnmQ1g+SOiSbYoJzrsv
vSzmMqEPztcoLh4te2ubmc47noyAyufP+uKRnsUnuyI+q2vHvQuVdTPkFFANyB9B
tytUZ6RbcqwritF1ZnoXBeFwNz1vS31b85i+T8G3v8RhK/I3UBE2zAjfYt1VyEyP
1XMdeenAKAIvUd/10GGSXt8Sl9Yt7uVUF51YxqXsCigy5ps6yDmRr0rLNM5UU+Ue
vB3CfIJaBYv04hmEAk8983VcGsnKEg7CNDX8+PGDa3Vj/R1wKSaNhOwirmUd/kmW
lO3PndfKl21te9YKcuR90VoCUz04ZR8pk0n5EGU3jxg0heORr1aBAB5RN3//mhaL
y/1ay4XF5aF8FPnLdBxINX1P/WTqeAXl2JQMiJdu5sFt4fTqEeft1PtsOny0DV4M
nkdSHiHmJRnvSjVMh4kh6pzW9XyRKW+F6PL1EwYI0yXgRGHD6U2AmWAWLAyqbgRA
GV1zLPiq3bEhG8U3/dnZYtZTU6+0SYzwgOUYcQbpTYriFO+KoBQLH3bQEvtJzN9t
hDArFeg1Cyb9dfuG5aVleECJq1Jmn5VhovQBP3XaRnDxaPIE8mL2LjwlOFiVZrF7
R8UuG1LuEYy5uq8ixqqpcYm++Yc1HFywv0OiZ/T4EYFO0rZkV90+wr/sHSvYfRMw
sBVaS218loUvQMHr20FDaPA72YTbF2BackPOWLZaLnv5buFpt11DRLPGjB5X9aCq
J0zVpiIC1Rn+tYW+qOLPCW2daY0QA4oOLEspE6LVumDfj83gCwGHgCzc0e/KBaq9
7H3V0BJTXp3293Zz4rNB1gxU55gSn77JKdbHSk6mircWl3/6KJcuUvLSUzsbGNqA
KLxv4OdHk4TMSHvwgGSdF+AzGWJqYGSHpSgerlMtvqvi0B0tLkb1keQWkCz6vz+G
yu4eJJ9q98e4UNVP1RAvrXK94iF4+XR33e0sWqLNT1uDPZdEEabjV4ydNNf0hR8d
hR7MJkXxAuGub7MGcmLMDCjNsBbGhBg0sCuYoOhivY4QEeJOjX6BSwl9HwLz5KYH
c4SeODTGQACcjAXELHrx8PwQZf/N7KSNFx2csZxTyHVFYi0FsjS+D7+LdEXLGftT
W8oxRb1F8CSvsxnwdpsk9XH6vU6DHYGHNSn/EEIZoRJzQ7AsVP/gyG+AZlhPcwbX
nycYIJQB0lV4cHPN8IVA5sEN4RDHJecFOOFHRZmphgrSjObpebwyBok26u91Hpsk
6AAT+a56T3Y3bWTh25rnP4f8032koL0G6Df6dWUofO2Z1qY/VDwchI22Kf/l3WR8
CvpNPPSZ4gWh+dm4i5EKNPv4qh5PezZxObMJgLTcu6MaomKOutKy0DPrvpY71IDl
zf51BLcJVi6jO8WkHQQvebUWHX3y8ndoOKYwCsqXbb37mEHGMc/sbLBgY2afc+c6
I3sRmz6oT2f1j/BP6oKlgo2653n/HBDFPHMPa5XXrh3Lb9ME7KYpzcHfg83KXuEM
fv1IE6Av0uKkg/aO/lSrxyDWW0A8zbzup8DubPgnrqaTlLE1EvcqkUlm0xBGBxjX
58QKSl/L+DfXArV/Fmn/LBKx4mjOehztSP8stxCTTgxOg3NPKXciyQUCSp4segoo
vZYiyqjFLbMRhg3so4rkI1uciflOd0lMSvR5bxae1jlAFzX5IYGz78dOv4rXbdq+
hnSsUQJ+397h32Kl0c6WYSy/IRC91rGcP2PMVlyZBevH9CXhHrS9C2sRKl1KKqCb
C1+uj9wX5j86nsfxysgGq4EbSZX+l723Nu4Ctb124Hj1YZl3uUTU8V7+kGmorbRn
nNlrt+m/O/o1g8jLF/wP4VQyQOSZa1bo5Bv1hqMtGBhpslsS8O/jO5N6B7EfFZQI
bIjD2Qvm2skofs2uhUqkPkWaWbtXnmBaWp0EK8sv8G16g2rjKibDLUHPHb+TprNm
C0vEKh/+iOdpTDUTyVu6Fky0Tt7zUR2mQhs2NZZRUAok3JINZokEcSiuL9yjjJux
WHePe8ODQuA2M+mNb4a2s5vwtZ4OW4fu6vj1j42OQP6ol8mBNDgk1LUUoBh5a/C3
sRYqRsIVNYa/0TmgxsNj3oxmDOttyEIj2Ldv7Ry9ke1jNmWzdwgAEq8J8Z1Dl9AF
YRdaBoZ2et/8PwBFOmBLBUWG3ctpsi/cbV5hZw/5dVTB4MaqPByb7w0hC0wD9sat
9TIJYEBNtqp+uCBVKoQ5fTq82GPCXBWYDSbtbi3kZTBWEhJrjf3LwYgEwHMMFmVw
0Q1MnGT95Viy4Qj5QjnuWPYom86lk1VEfrhqSaiusQBpdmEMAg5GVCm7WYvCImqj
djvmzcmnTRFZCkzAjbsgU1Nu8yLBUrJmqLa4ynxyNDfvWczxyIfux5hvOfaspEbt
SyNbzZCiD+yRrK0RadIuxx8Qqm5rTYLGhWQxIO2242GQQ/i+iVM21al5Pwuql0vR
BWnQYZKoYqDqhoTFUBdpDDX/CJqEk/eo8xAOR4U2KGu7EQZKLWgzWxYMF+qh8PHk
XjRLdz5WH7rDnQVKQTjwWZTQlRB9tceiy0jPX91qqrrIDGaM6mAE2allqSfSvvvw
odnLM+Tbn+7FZK4UafQyht9uETFkOPaRvW1eGOmgouajn46oawUYf9GuISKMECPe
5D1/2V2GbLnNTQhRdDXTc89367HDTHi7pOGkzym5lkXq9bSmg3YEWdIxqm/c71a/
qOnfzmDv770qeLMaxU9L7LKzStIGYb33ONloRmswW1YA8naBxbBSUUQeeeyORJ6K
5N1CridZqcro+ULTISsVXluM3mEk+Nh2Gk30gJ56bxE5vkYseCTXpuMPdjvxu1Qw
bpul1NIOvuuBZSBCK+l/pkGBELFn/tkdFcCNOduqVcZ2kbOw+upN/EJOr/VbnllR
5YBvV+upnm7NqJwzLaL2K9BnId5oHbZDQcHAhYesmUh9fSntS8CISfi0ovmSlJgh
UVFnlA3H0jl8R9Sbm5MjJMOQK9UnKBXVZ8gdnzOJ9posKsykllWOt6568WHf2rV1
gEYVtEfcPcsQNGUIvrrkttoLt3v52cwIRJxIv/bvJZrdNP9kQYP6LCmg/WU6SPLd
578lCr2z6W6uU43ozdFfRBISNYi3FEWc6g/OPMyM+z8W/eg0i/lAJOVNDpFRLDxB
6FYLaQ/wjVhoR8cW0DYRyXXenoyeBUW+pyGmQ9peJHnymDizJI9yVJHA0LE9yofH
ZH/j8CBhT7KVZZJgvqHQB74XglbUxfGj9Uu469BH8JI4qI9DSPh/izGiTMM+SWw6
W5rAleOU90COMDKtrICw1HX8WJ9MdkkBdWgZB3v+wbWiefyC3t85GM9eggycFCYZ
rVJNTZ7AG3QN2+lTiUmBL6RS8fFKSbZxQXfqZtUc3Hq0hfsxdpUA8POBarGN5LwL
Adb1jdDDNOkljFMMdCmGTE4TT6loYagQ9qZ7yIyLm5jNeKk/QcH/2B6Q6tQDGdpi
apH+qYrk09A/bgxGAEyLcj9Cy03ctO9RgzMhJXTDQVQVPeDPSHpsM45YxjaaNsWU
DlWkW12h2Ws6dvi8xKTV7jbThpvxTCLNMPcaN+Uq7+qXao6q94+KAcddTrr4MaD2
N/wzPqZ1x5iqj/SqCMpotGTZ4kGiwk2xgwMtGMCepoBQ4/WgokOcvNs4oRoWZKi6
YS+rCWdsVYUbWCQ0ye8rDbliFJG2lJ2H4aR8D7duqDn7Sq0MPpAtOfb8bzOdGICz
xGzIdfMLLzDuhZ/NHfdykYDjSrmZjf1AZX91+ARHraKCep+PzwG3R2JoemPw62Fj
Ar//ySsd+8GdK8J6wY7a1eeo+P4tesT4S40FtO32ZHVTptoJi/A/AaZPMjvjcJdG
9kqhbyGvY5dzUl39oRQ/iRUfLqBuEEXTurMF1aNTi8of3Us+vvjZ6TFnOfG37FKt
eELK0nZqEP5WsDunEBbFI4ZkTtFf0jTDZc8qyGELku/Iq3XW4gE7IY522Rxl/CDy
u9ZJOsLurJJSH87QAzT0KK3hJTCbtJGmET1sxOVBNd1d/27M/nIPo6O0VZYGDKzY
H2a+ev64z8CpG9kWMY8aStGWySJS0SITjhW7snKM8y9EG5SIN79PS8HIzAttGTo0
24uWlUAq9RlrSM3Ch83O9FKqrJdZa0n1dp54LYdp0vbks0otHXMNf4s386K5CyaS
IRKI+UEoIm9bL/vuE5yNxr7MdewbTNHL66TU7KKqAM0UprGcFDiTNulPZLmpAvJS
HT4n1DrD3asmKTepay9eQbWdvnmoCfY0kzxnJ2KfDckhxGXs9dh6KjJj8ocbf/Vy
hBW+Nbkq+zeScV1RuCZe3XaA3gd1F1R1HhMaUKqPKnvtUHCOuSxaQzF90BomKmO9
8rDftRAX/sHl7JbUKGH1J/t9ddyqHQ54mEDCixIvSUvXjUukm2UmPaDW4FklGVlJ
Wz2I8Uj7N0Ub6vVTy5rOl5N/Yc9jZAjo/ztRTHNxfWYGOLJHsR7zu4S2AHihZd2i
RNz/VJWZ6Ug2qLxSrdPIPN7PUJdwKtrNoLWivdKC3+bPpeQ0LcfHkq+UUZUHTS96
YB9KEZjU2jas99yexhyUjS2u6CCLIQbZOGCUzFryPKZJ9bzbdAQKCXEAhH5iCCD/
VmGQ65d1CahjZVztCZ/TTs4nTq3PWJiqejtQXxy2oMhSHrENKLoFDuZawbEsla/n
fLRFLUFP/01jVt8MdhCrrd0AjWKcWBxYUAeWpSoZTXjukzXNyIBO76BAE4zFFVpD
6h4MbMfZ3Z97XH9QBPeILXJNbypWl9tylNpvPEF0MrQrcS/KAZ4ZVwQz5FbSJPos
vlg0CtEEVxK/klsCgI4NnIy7mK1hSyq9mkWP+oX+1+IOB8W6ynDUfRqqS1t0TXCY
rLU/88y3Hp84/qklsPoA6UGOXIx2GS3meNf6pOnpBdTRJvYa/8pt4upQxBYzRInt
Lx1eOJyZYk7EXKILZ2n+JOYMPLhgGrxR2N00MY4mpruskmnn7Y+G+zMl0u8CZ/1i
JlMKyVQ1rNS7roekyFV5tZoiNlaERM+/dFgspwy2NDxZir1DC++TZFEHTjvJvEfK
9cxQsx7br+oIrllb7avZvCiAi//AZ2JRVllY0fePGcZMP1h/eFbgIpXVpm1rbQzp
T5+0AqeXBWFXww+1mDyz74U2/ri6bM2AHlNkF+nsHoryzMRj2QVrEIs/jq68OWYR
KdgxRE3OOVUJxN3/4117Uk1YIikAg10WmTakUeohYzoLhxG90ZWnAS0PknXwrSWI
h9/yuPoAXojmOCLgSgW2kgJxTAxqdm8k3EMsOT/puBIgBx/otmpLiCBaC2+tteDW
qj11JKA+27qRnOGWdP+FF1nqFnGxmQDSn3H8C8l7zoPgoO7VjFtK8gCvp6AvGcab
qiuDZslbQeKVYJYNxK724C96Ti0bye6z07x3sY9Na5hNBAfGDBEiPff/ctlUNp0+
mvLG2KgG1JCOGrHlHcOqOFwLZfQ7hIiLYGgelsaO2Tepue4ShvLb2+/btmbARxz7
CG1p0KbHvRJAuLIlm5ZU2A+y9TD6ScevdDB1jMAMRjvym1wWgCiXxshmYX7iPeRc
dld8xzsQvJMf6MUqfZikfIwZQdhcfy5YK4WNZzYA1MrgKs+5lMxlkzaJLkp+YH1C
dWw01Ktdqqnn8XNQwEuoYTtm4iLhpqtj0w7rrYpSUGSaJTqrcYfCxs2HzranUJhh
ZP+yKWoHIrKKf232zMDsJq1rnP2o9C3gvC43BwEwO8gaI+JAN1ZoGYtWN4qmvY7+
5NFB+nnYmtJadrl5z2frr+hJUAwCr7N/rXqSKT6lz82dmNZ1QvrVfRRWvs4Z4ZoT
C2If16THB9w6UzuqY/MbCLvMpVsp86UNl0oS9kBFoJEwZG/l+BelIcqfJjHznhAG
X5OXq7+2+ysmspDgKAxkea8HEguGfAf+SYcWwJzW51j4zSEPz+Wh4oLt9wkNEmWm
GfdFHlbspXXbluS4dmtyNa6x0VP6KlzhETcAmL5NQL1FWnxjd4m5qt3SCBl75E2q
61gbjte5QGInomJ5PxbhZKDBk1mvrtinOW+SwxmRgTVNHrGeA6C8i9D0J29GM0+d
FW8X83nSBHtHmM8TfDbm7Jhv4pEsVqwenO/zwfbvaMFfjWJNkU7dHhxgd+fXatIL
wFzvCwuZZS8qVKWth1EV8dZcbY0r/ZfBFKVxLLIpd78vM+I+LPqq7cDVGw/n5ezO
kxIFapG2LlM/RnexkyIKm5VwPnj7LvlQF9N2L7c77qMsT+FnstP5gOBpMj/qL7vR
ICnhgUYwDdcqIxsJDVKBvYhOBzjJmRfbN1t6uY2Bcu6895hl40561XIg+BwhvAo0
X2MB0g+ewHU6MUpn/8le4VaGS0hxhmwNyPs9AIMDtjlIZaCBAN6rr+Hro0biwyYO
WE9x4VGmgZoDZaElseri4EAifk26cZInFrjiEMVlXAaArLo+caHB7UvxGD/2WuLV
1fUEwQBZT3d7m7JwCk4qgl0joEiZqMOZ9U+pyTpTBP+FK1XuxN3mKpU4Ph7lUTVj
t86+1xh7xzTRd6jGxP9nEh7ssD48ox7SyhYdcnbONvg49WhEwrcKEDKEKwa5gnT4
aGLSq9XQbGjYz5VS49WGGuwdhK0xSb6RXzOoECohnHbEOEkz+mJ9owjPtwN8IgcB
fFucM1gwOxKUu1xsKAnbEXVSamJ/z6mvlPVudUWKZc8IItulAUYp/fN9WgheOx6x
K+bcS6xmLRf6MspGbvIoh0PF6P1a3yUDCCJ8qOx5fGfR7XI1ztl/tURpGaA689DQ
S4sUMgACMpOL1vSuZlX7uEwidZU7nTC/xpmGr0KkR7ND5/4eQAdGvcOLi33XxEFp
V4dx2pou4+b8ZHtlZVFv8zY/OcDVnPYtl0Y/1k3uypcCFZEeEgLS4Xte1jigOtgZ
FyAAjDab32ErzCjSVrEn8+FFMrR1BDiDyZpAoLIRixTp12nzjBI4yp1aVAhjSu/i
TQlXnRHichPTxdBqYzYLZgkBQNOZDnn73YB4jmnTW/cP/Uz3f89BfQFs6/CfBGnh
jUqNLYdW3cX0r2Q9INNByISanKtV9UHgi3XBX8zZREocHCdGfvtYjp/Get2HbE/d
F7O0FrDY1zewpdz6dkBy0zAXEyi4jLHxq3sArMwNpMicOP3oSN/QqCoTIggxM0LV
Zw+lTR3zQGu8pg+vRgWBuwgvgn6g4BpCbAYMcciCCVCusKDnndgLbcInAcwzO7gV
XdXshbLj+uKgZ1KDWHAnf0sar5EBeBs/wubJ4+0mSkp0Y3+iG1Mi11wfLl3E9rGS
iAls5lnfPX5mh+cMlII9NUU1eIOCdprQ5A/tRg/9H5mRRMH14U5s5ne6PJ0/imRj
flAsx4G2UmsYLPloams7nuWtUc95OmqLK62EsH+fhpE1xXIirLEZ/hDtkE+PnJ++
uIHoEcFgRRpsBJcDsl92ROeyplqZ440zB5qiCmOo7neeYDu2Vqd12pr2xKXeoj0W
dCZ7aJ2KCKxCiGlgsWZcguWuvxQgL6focqJq3gaOIVEmOLo6+gGRocS4TXKzk6Br
tHTUmNZhaCPptraGERHGISgcBdN28QvKNdWn3/lxOetJi2djv5+9Id+yqeo32t4o
c0THHoTXAtG5N9q595S8xhv652lzSp0eEeojzrxwijVN4xhfmbbiiZ6P62U+EgVH
MYwBHJwXRxasuNJ4ZnHJkDKKgjpHj7LawIjprsXC0FUZaZdbPX4AqThRaZuHMzyl
BN7b5GGoMeUf952oqjBTg/fNJM8PP9EGGbMWIVpiitPvQ6kam+0BLolx2oSfw1ot
wu8wv4Q0UdpnAqhzTNbk4xyQt7HZTm3ci6Bj4Bq/WxQUB8RlmGpnEvySfI2u5hr9
ZlZiwLFJ8OniZQnRlBU8j4+yOONyoH+B7jN45oILmbNdBPAL8xyT86tCXVSWjRrx
RInnXaaVg7DTUDafdv2aVnXc4UGsdSP5wEOhk0A4ODEKjzT4U3h9ZQfYEKaWqqhA
wUjyAYbggMTHYjpPhhwLRJ0HKTfkDViDK0bfle65wnBE9AJgpfAVgFBAAIDtoOg+
3ka12hZMmLn+NBrJgxUDWj/rzIt9K6VpiuaU0Mn6qYIgZmLtlCzWfTILre6TN7+8
5dr1ciPid54NBKV/PLXHZGugbUXORkvSyK+PkD+UV9ZDCV637KHQnkc+refJEyfh
YIvPV5HRB4EqnzadVBhaYDSYjgcAUslaKjQQXx3hh9/Z0jtTs7YUwzzPjr160gCu
R8Hgvu4ihrD5OW71jycmvd5PYmWlkHsbCRhClp+taP0rlarqObQ2UUTOVGy/StxT
kzJZ55tk4r5VxfaE3MLjowLnphbu7t3731F+FoLHdz72Y/LYq/2O2imUcY4UKJMh
ukAEF2zpvOp8UP0j9PQd69wOyUjYleQeG9XRxB2dzjP8YHz6gbwBrVerOkWGf47X
QSZMO4NYHSydQZHHEE+wkhtA3xqC1gQZUeD/tOn+L/7A7IWtMMTi4E5CtEBVti9Y
557tFt6rN5h5glQb8/lLTYeaG3OFxzolepEKnEoURdnAIGkVWVw2B2YM/znR4McT
OrS8OFeUYXSMCYQdyN3QX5eZulyWDLtkDypJlzZh2JgNhnHSVQ87X8G0PkswdoCN
Rg8vOAMKwwBjI2KNkyNO+sEAbBhKMVZnvEx5k/dlxlfthgzREY3otTfp1BeKWuL8
fqpxsCIdv81AY113qprt21QF9XfrAKl0dpyP3orNsoEjgtiMmP6rGOkqq4wERK52
MhEXzglzaqkr99YOXdPjcks13FdkuM0DimgdX4wARiSpH3+gWL+hHuw5b9Ilu2e4
CrUrps7rFTyVn3aMWe8EyuYn2R+o1FEaGxl8ddy5K8havgI+rEL9mQD1vauKYUOT
4Ul7wsrEWIOY3f5ebnMoKdrd4sznsT3Ank4UoFRNvCSPofk9TQmkA/QFi7rjEasY
QzJF6dzS5smZ6rNtStbBGMRFc8P3xDpP1nmV0QkPtrQr4SacvYl4DTG8btiyRTxG
CMzTFaZAf+Z6NtI9Rv/FFwFcXdd3n9b5kdwE+5hxYEeyVND38tcuurJMf5N26xVR
qAnZOgwyCEVYNHjV2V4L4E96ta27XoTToTuKTOFRrgJ8fGxr5ClzQ9uy5IgK9bKr
i9gQRKyHIerLwVST3er1ibU7kVhKOkS6VcFB8QtFGe5LcRJovQ6YKBk/si9Ilu5t
yOs14Et344OcvPSl5EzKHGPzvE9mJsMxZbmff3Z4M8r8mQ1Xf8Jj5GPfg4nhHj6o
NZzM7Nlp5fO99+lASn+MFcl7AaoaRMxfiDoMuMr7IginnMLwHs6l3lwLrlyPT6MK
kzi/ZYa2F3MCK1gr+kv4GEjhwMdFQw4hjR3xNQjvx0Jd7K1YndUia6rGaV04A1QI
dTSkcB/qgjazyq4hOaqXKmxz8HsV1EfrfyHxuso9EEElJ+RNUIbOoKJeQN431TWh
KelEbQcbCfmr/Ecicj6h+u8G1whkvxlHZyh0sOoKyISFAKtouy4bpVsR8yG4Aq7n
lKPiFpkqcVQPnuSHOJQR7Jn7T9IzFET6XY541/1aqc0D568cL1tYaIfJsYB0sbBs
IsnxEmqUxXv6o3lNiuI2Bb2KVWO56KGMfsEWek1uv6EroYiWHIlCLO4Ufg43jm3B
CVcQSsPsukm7tiFN0jDkg+XZIZ2g6oT9cOPYOtSj+wo94otDfkWA6/Oi7fPwedRp
Hbw1YO7twzI2EGwdvHzx3EGVih55MfX6wi5EJJ4VNDUnY6gsbdKUCY0KOTqNCNNS
sXPED+WJwfbw/DqxRzMV32ou6Wz+mYbBrn7DNVzctAJABd5iIoHvtZmRAGTbN6F7
O2cBHZ2oQgj5nxDcai6esR00dCIdJsG0T/SZgzfWjt+NtGUzM9JS5YYlwREePksv
y3WBi+HvrMlYk0gWG+SsuJfT6MU8W1ZDuAHLQY1ts0BxLMtuvASSTTJbroavTyyD
4saofO/z+xzo7p5008L6Rh5pfsD0/Vw2MgEkBm/HBdNpTznrqykJMqs6D/QMadhY
7/lr0ILKAzUL4xXFsWS0dqNkDA0hArj8U63ZJ0KRxmzw5+lsH1H7Wm1JN39On6Jc
RijP8EDt57foPm7DGnZQ7Zm7mI5QdQHRWfCqBOz7g7UUku9wT8eGjuDtxlm7eT2r
7svOT8+pIy7MawJ119poeLglilIxGyA+urFn/cE6FnXIQnW/zA3kaGMiLG7RmAXT
nCQUkw2kI8FHkdkMynLB8cAOhPGdSHn0vrZw7WmcllPc9PYmMskIBrPGHDFzSRvd
lVkM2n4Mbspi3CBmSMiPIiWqA8YalVqKGajLIXlBSB1mXbHqOZEJ8RAEVWRsGibA
58racjBaYslBySUOAZSUdAiC4pL0viH9dD3pckymRecHWXzq8MYqc1V5YPGrPd0o
beVp3+jroWqNPLeXW732qulcTqQPIcVLtuGzTTnzvwXt+o7ceNnqzOQyvlYDCTB8
xh/M4X30Lb63OBqzZ0/+YS9ZQDSPKWJ7aZuObEXd537bD98qckSlQVKNwFDj5y9d
kkeO+z84DleYZBBsFVQP/uYDJp9Ltt4Xmh0nwZoTcepeqFPw7jFxnMBWAf2NPwF7
34gTDxg7s0Q07Kz45Tab3gA/T4ZANG7bHazDrzS3hew44Z5WCfpmWA/Rw6WINKc2
Wb0OgJQx4buZOrsPRLtsPbSQSRGxVURo4HxJmGcMWfqiBr/fjJElVqOtvHr2GsUO
jNAEEQ964hc7kfAoZM60tn0xp+fcd46h0ctJS5DGwQULsLbTVAhTSk/AnsVfp+zJ
sqjpq3n4IlDU/Qpq/Aap4ADfO2Iulcz//97LFemDpBM8PjuJ9l63XRs6taHGzizt
dZUXIgo06x3hE6UbpSp5GMbSuzvcF7zWNRnWW7OGco46Ot5HXS9CeyfG49uzJOxT
q0FDAsSUG+GF9D9oKKH7WC4zYVhpCuwR384FtiQ+xrRjz/GOAIReqlUhPAtYW2Pb
Xfvl5XkihnhSb7VIj0ibZyfMYg89nz+loKDPJ6SLA1c8HzSHZXeaNczJoXLpwM5g
BQAuQvFqK5rtuHZf/TAoG+BaLWYfmWnJnU2uB7lCOgjDrp7HTLYYUeWuf1+tByQY
iBZMyawv/U80Q3+qx1enVl189V/wEtH1e/8ZJ0X2bbxk0p6+T/06tFujH1At8SMI
Y/OwMcYhXZFm3V2idNt/Rdf3wRhKU0kv2ugFVp3V0huvRv5i2PeD6UGqDZGSlUjh
T8MhiM+DQJGt2+zxTXpslyPsm2s+e1E913fPrjinBInhksSrOQrzQ7qUZwL/i6b7
xfpCanZ7g2dynZ8zXQ1maqsA7HnKUkqlqT+BKTHfeUWZZodG9+ZN3eRo4/vsxbxv
3DrBBWcD+g4p7dKAaW5nVGFO1XCaLaWql73F8rEgH74n2QnhkYx7zYUnLZlV8m3Q
qdQXsUS9FpNSX4K33wP+aiwXdqB0IzPmqFhmu5ZHmFku4HNmPdtAFvkK4MF81nP6
yaPdjqx64QCFJjgxHX0HVstf1TAfvYicWokCmdDXxpjdOktLQhnkIpdfRiIGxyMH
SrNQxhxsYgbtFpW86NCutess4V5a4Zu8ueKkoQAo9j5t+Gd/ekip1aYy4L6YEPoc
AzcNStrV0vUeCNwNUNlrw9NvFbiz2//qJrqHN1+efifMMXCw+E62uDDhyJwZuN0N
HTM2Qpkf37s2WK/AvIkmGysUSB3JFObYvJQDhF6wc5usx2BFn4n2J2lpiHKIe58M
SypVmU97DEID0JteXeV/N61k7xUIuvNLjaHs89LLwMXresyD2Do8LcQL/UjT6jy/
l3oWrP0XOkWuex5mBqIrM4vi6f9t0Rp0bYi5sugQ2E/pNNl0IZzgyuI8jqJurZoo
aNMQngdlzCi3jJa8+zAUtqoIQxC5KEU3sv0h+0zucnXT6YdNhgw2zGszLHl/i9GI
Q8ab/gP7IaAIofbyWOGT0TaZr2qm8ppq6/1uhKIM+1kkZJibFm/x5XOlHuB1PMrx
qc8ZhRW4uCHq/t3yGqZgqEvDccV0kC0OUQdgVfX+RtVn8R4jje16HOeFulQzaiQo
2Wmu08KhtQKqRB1kFyLs/bqtJUm3SGvTVNh1xm4dln6kEiCiueoNNz4K4FSZ8eHs
q9C5MgzR3olW0QffcpIKGQZ/ZwQ/Y7RoLkswjqx94Bte8AY27Dzuw9V8PUdssPwQ
iDgBb8EsqKnHja3ISG8bvxZDkQ7Dc75JfhNu6fY20D1NmzoS4sFgOkSAQ0Sml5u1
QGv3Vsrx1XcgvABSwI/Q5Kb0tpgSmWnrF6X+z8hG6UY27hskIMSPGTCOnsDy8G2D
RpP5wIR/wHjN26zijHX83R42aJoGl12vjHsdV8MdHY/ZskXS4qkgTQABnHpPmol5
FOvt6Y1pBnqO7SRJvw8O2YhXfV4YGnwKuYN4JjXL571oZvfDnH0XyDi/eJFA/fDC
rxBnlTa3Zy/ilBVFbBA3CKS4QDB+vOYdmAPsRJJQK9scdA9d2ovRwOXQRGyjCkAX
4spCQ7//VoLYfjseqPbcVn7IAGIROWMgQLzNSPDHrbkKcs35LLsE22wZJUJRoS8U
//4onUkt6XGYE0299BP7VZUHq9hukpdCrdSh/+xEuPYaK5rHwpD+c2r38TaLn8xO
EC2NR6fhfiNnDbPYZ3rnFXwGxm3Kf5xb4NQlurvAxXWWa58SJIyj5lj6YM6TPmV9
KnKNadFAnfwTEvpQYxNZFb0QshcRkwKemq9wB3vCUQMGgtawq+ylSyeLPeR4ck+k
k7LD/wcrFvwVEPu/2Ie5U3JbDD/FuzjKRxxrw++ECY4OllkKy/rfmD5TIvZ1veuL
Un1unmbta1Z9k/NfUbbT04cOzHK6+l9r4hr06o3uI7t6Fg3a/wb2LsWtGQLywGzN
IUU2gaohko0gLoucvHAs8qJW2WKf4qttfa9/17K4XGqNCxaqmMIvtOjTWrPFzfr5
Nb7vvo341ZDkSGgLkBeR1MfwEG+3lByRuouwKFm07WqWuI8XeIxGfPEgIZvUFFgv
n7OqhZcXsdt+ahRonq1BwnelyHApil5bAqOaH/PFErOrI9dcVyHxDoCpcr95E59n
idvforVNZo0LkkyH6X1TbYfpdExLyv+m7FRBCoNNfnl/g/aSCWSUo78bhKUUkT/C
dDAzSFTxQruCQ7sIeirKYr5qnNX9lhWG1GYVe3wbragNI6JEHLBpO95iwk3yWzvM
8GkVi4SigDNXTYMqr2iy8nGr1d/8eTVxED5XyFJprRAQNLcEVzdWCMI6nCOyUQD3
po+nq5GsSdCqIjQnpzek4zKv1xVWhhA7gTX6fRLZFYTlCH/Xt4wec7Hd2TPx4kwM
zDTs0Y0Y8c5O57Fh2oz9TCuzTw+SvUxQY2e6OdLWW2W6Eg9r0y0cV4x9ufCa+uHM
F3XF346HSNzXGveL5zltY/Dv82190W633JIoklLS/Yvl1n0NdCm4nXArro3aPbZn
KjlMfCoOpY9QqoF4ODDVI0GydFX/uMbTV2bQuxDtxGLXlvdYDl79uysy4OOWXy3J
Mdi20QLm2KESF2p/GiINFoQq6QmtXw+epRXbZ9QnyVlfWG9eLL3MSYad3T5xF3sP
4nVFlXkRZTWC/iIs3feIK/TJFC/m+i9mEeANLoXFCRPdBdko6qkqQbPwsPueWvBi
vGsVsHPLqBgJJLIrvB0G3MGfKYEWDpb1MXU3mHhPwe0HQyrupuxo7LUDPSVp/w6u
Z96N8VmzYifhrn5dbjP6wAzqcZkAdy95X31yFXHv3nTtwhpYXR/8gQgstlw5Sh2Y
lRwrWr/loS8NoVqSvGXVA551y9YInyV0ZbYRU7IIUq1LcqD0IguqZ+3Hwo0mMKTn
I9hG7IuDHlEjEsj/kv+2Ms2x6UUosskx6RMHF2mvq2bb/eq9jfABFuZBiPzyhwwK
Vxh0ZeuMo6q966F76KXEDTizOlcBe1vP59RQL1SC1pVd6AsfvoBDklHoN61CywQB
6pBixHV1r9j3sHqu4RLxWKZE5m2wO52nkbUTEh0lDrJQ4iiPcerp4zBqk4E27260
tcrSBiHWXiuJK24WbucEp8i2MxwBYNaQNRs9XynXS3sSLspUoUkQHSv92TKD4jy4
cs8Vp1XP6d+r0JsMURRbU3R60UNPhXRr84TUkM/IlEdjPRlbaJw+AKy4mA9ASFJY
n3Db3oWI5bZQgPzSdpCC7AKNpvSCNuZZJOH9TYm1VRTvZLJKu6uphaGc+18HjYhO
BC3cNbaDTPVLKsFSWiKBhB6WgHuWEYNIW+uwMraII8W9Aj9aJZxscomk7poQPfQl
4OL76+GQE2xbukZqmKXj//F7MACgSNet4JfdVo9PVufim9m59y9UYh535jczDb1G
Bo3F9ziCEWwzhf3CKlDmugPGEDsDE7vXIei12WFXXV3/7yWH1yrx+gewjNbvHKGA
MptyVWPhCnr3SclmfOFN/V8+ERLBy7QqG67L2oQdwmntgfZlZF0V1BtgsXnFUeWG
M6SHG8VjyrqOYMamtqiDK7eVNveT8R92/seLMebzBLjn9xVDUnf91h4DEeoXPz6g
ynxgf3oCygNywhua7wSbrgNgi+HRjbdb8DfeicOyIObzFivmJl5AbTd8pMcC1h1D
9HKJft3sKrnkla9iHGQCvGSqgh14SEux1SzvpHEdXdV9Dhxq7XlOVo8jeSQ3EGuV
OrFrwY9yMb1oX5OGEFd4kkCPNHdpycEF+K+RXvJzkGl1xgGYxmTlZIEjkC/L0GCR
OJ9rmSVvCeE1fp0R/cFFJCx9BA6vB5T1ZF8tzgl63PKCtdTQVEFTzAx/IKZY4YCd
spLegiNy1USniYv9CZVZmxq6Tt7Ali8QfY0kXvcStmSWjC/btO4+0hzWDsQ3x5Qm
Do4HqYMv7Vhvl3Cn4NHl5sUEljLhxz0wDuvjUiezWm7OoW4+rrVmz2IB1hnQ5bja
wRLl2hEKoAohqh5Yi1zIsWEQjpeK2zqGqddY6Vx56EGU1QBcRUcur9VeU27ArlD0
BPF7HGTusl0MJN8b7us7TLStQXGNLjJyPnqcK6UyThc00ap0yj51H8mUYilR99c8
2tiw/SGFxFlSeZPs8Me4Ks6h8hvkD3djd4Tnh9xnW5aXKTLInD24opv0fCtcU2hw
TPKd6VTZPz3k7LPPRSBxdtGFXxPrEmS4GqUrrbZq5Qf5YieJ0d5hcIkgdOVg9sFo
gxOpuTkXHGkGCN/kbKlvbn1m9gKrHyioREt5nVpx3iOs4Ez1QhHsINhTXorRc0c5
N83c0j++e4x+GURcgUASefcNCvHhLMgjcaccPlxH70jU++ieu4/5cTNl6351Gj+x
f0FoDs7kXAZtpakaJ2YK//XzXpZvr0zjupgRWdslhvC4iYnL3O7zHlXRDUzzPY80
Lu9bjO1F2tnHf4wlQH8yLSgDMiYG8Nqm/m19BP8QjMWxAZxtBfpcxvmDTB2cdOPF
PzzQcTkHDKBToCBiuAGfpo2wuBDrGkz4XmvCeMKj18pB3J9KJTh5n/VozqZ0/hVM
cnr7AqafnYbYpIqkv/8SQfXPyHki4iR+9zlFAGVc88F9ZeN0SZzagJsGiLJIVbUa
BwnCLMeH+Mm0zWQVPTFYUlDiuEqjh7C+SmAYsgg5WaMrfwXCKfoSDuxxMko/uQDC
35EUAYNPDup1EqokLKV+Nts/RP3uTGDG/tlk/3gUv5/bvWjhwrCqKz8h6B7gAIkj
SBpkXNRQrVCZaFHF40+BvpHpypM+B4vO3m60JLdmrZF2tp+p+y27g9hne5KVyecP
AaLkC3m+qGJZvtD5Mgto401mULgVBFANM1H2HQRc7OofEsbdsQtSr969RpFyDv0C
y1s2e/f+H7V+9ryBXW0m2AnR6iqpgw8FZXBeRf0ntxaGeM3527QqgWpFba91lK7i
tsIJixfRqjSA0piUTNi27JJqMYyHPE5spOtEkpk7NK6sP0u7YBIn90elJ5SQBzLC
meFbeX1lcGOqr8XcYGgojFIknPC5nGZ69G0stxvF9LOUd/iUwRUs9vdoy5AYiDcx
0O2wgNXkpecMeencRyVHikgFd3GldouT5KZ70L7SN+xNd6onsqOayft8LkOYMWUC
HBs+zgsz6ebF6M88krZWfsR9zukm1FAG6cO/+2rSJlOj6juIBMyUU+3XCbDfndiP
z4nwrziXq5FJEdyWlLRro84PhcIRzb9z9umSghqGXF8pimbBVXsBRwYv82C/3oGY
GtLetPAKrLZ8dMIECBiU6FER9GuUl+Mrw5o+qGmIEYg0VNl4/Wv9bKS5l7DjqSse
ocFKE7nMf+RFrrsnwZ8KQxqK0xKV/rp9288bISdhuRBSxoQRSibrvqPQ2Ki2QPw1
qmzpHMbP68ls0zvbu1zbo+XFHNrBcgafPk+XjpTRRvRF1e16k6vZqLO7KBGAgA9O
fXJpY+2/5CRd6QrqfaATDFRdmD0h2Pfbs1hmxyTGfyhpE0UcmKlwh8U46oQ/ulOf
wxfmfWFKXZDHaoePcdpfoF6wZvsHEm8+Ulj/NfxOuVgOKDAYaG2Y419tVMDL1CVV
TNhOQvJYvWJCWBUkoucRUAuhoOWizRciS3NK96It5WlhHkuZ8wEaCRP7s8zZYGaa
pwGBGkIfDDnOafqYp2tzcaf7kMsJkXqRXDfMI+P8mLcMLIw6Nc5ijr7oSBM913TN
Pdh3AaTQwkH741LRcssR2GEv3WlYIhbPqrw6e1McZ7grCH5ugadG8+xX6wM6IZXC
H2QFjcjDD6orAKnvh9AZXPZD5ApKFMPpfO/7TFSCm0vw75vZ7g36xgUdRiSuG9ke
X3P23npo+Ap8Mg5xNcqSF3lz6yb1CVm7bhbpuiqKINRFY5NJfgkIFm3mJTgkqMWC
9E5+hIcMHHR5iMOgbKk4BKpY8YpbFQYZACIfHdzNUe+VTHjauSekXiFYVPPHyFUW
Jy4NAN+MoukEPC64MkwfUJK6BItGkdbS5lCTWXM89ofFTMMiSv4phxTIqtGhHnxw
f++HSRzaGjJFy6iXQ/WrT5Krp172SsHtqBFHzO6r185OzmiVMSNIUQbGrvPSbDg8
x/ULJVAItpefi9NAPGFxbj+WuuZB4dcRMPPr+MN++3/BaZmZa8GFU6s6f1Thptjn
3iLfsfp98KG51TKB/vAvIb8vioAe2eq+VbZFYAFLIClywtwY40vg5MEoEhy5p5WD
lxm0sDHpQ5d1xeHRndmjvJzgchmoh5PfUSOYxKO6fxNv07hYvWHQ8KPR1RXPw/7i
ab1medKP5P7llhu0UTS2u3+6ml3Vbx/CM6O0XYAm9qMOIOm6edYFUY3C2O32SbyC
YZg6aNdHa1QPPQ77Ut9Wb0vN0cUV1ATxBe+jjRv2EtBaOYJqBA5X70aiBqiHT+Of
H+DjY+96qt6NN2cv2yvzR4fAvemF5LKezbX1hCIGiL+rcG2ekvCGT9puERABRuc+
BhsVniCi5yN93oPB0ZkfXsjnI6Gf0hzEV+To7gLWFeyDNAmFSzZnERfKzgN3S9pt
EmxfcY8R4qSW7Y+pJY88QtS/U7Maf3DzJIW0Ih56Be/0utoaIV7MAMEeYdsQlDIP
F9I2RxOVrYbdI0uBThlZpHHRtzLdEs1/6FWDjDoaUxtKSf0FlpCePkoc8DirTmwG
sbknRmdSC/8zg0PbB0Ru6B2GzYsBMZUm5A3fZXtyD/2dYJ2JtXsrtiC5Ye/RRDrf
qbL9qFSU30Y8MXInDltOIBRAdUyLufF7bdrJ0FK+WGQjSThGtZA96SZLiRfVc0wV
2MvR08zqtzsbwUb8fSTnKKvj2iYN11RiNQ52eKW66d8sHpCBlmHPuGYIi9FAlLC7
Tc2TlqBOGdjS07WLeRRSSLCSbPnTbgGSk+Vne/taIJWzqCo203cAMEU1SGt+COVO
LORIwMEQXFPaKD003mFltj4wlKijNAVEg4CNE3r7GdKYtmGzzqI31ICyGwvTLV/l
7xsQjU3SXR5vBad6PxYMZmDj17/lW+8UVeSBorvRP1JC9TfPOERPY97yiFaIiwNQ
lQVkAP1pi7lFXDTi06L3msQx5/SGQxB5pibxsKtuwACOzuk3Ikiv5VPelNyfeGUU
zya4O/nmXKJoCsS3hSlT8Ehw5jcm+M7oRh1Sbj7E/Y2W3NMiniT1ciXphWbSXL6c
LFbmvGiKqQNzk4Tn+8BD4ueuUzBdj3gFBxUkZqaA69sleqUjjQjnIAreGPRR7+uP
vajR2J2MoKznDvsRcKgH7dSfIunsyqISOcRz0WWk0kJwERW6ed4egWkWR/t8Hizj
9t8IoEm753+lDPTurZHI57R8KFXozYnAHhLkJW9SujeUhNqvIUUUrJZs35hEB2bN
YZksI050otsD5+NKhAcZIJ5GNK6hoKjuAoz6Ey6T9E5v8ljCXF93LgXNrU29Kisx
tGeffb6MZUE9y2gXhLhGAQ89g+bWBiIOUCjEkQzw+/FKWN+BhaLW6OOpJ8hIGQ51
KJiih5UCCfoZ079v6GP39dAZqFo+JpMP2Sw0Jz0nHcpGIVKSW7qRIwlIFDWfMXKb
LlyyZVJOjC07jSG3FCimUAoFNXrYv+AnpWlaJTlQojx5N1akwcLn0GHNW61wzlhr
Xxxe46u8LHwLk4gVf9Did8DRILnWmHejw4XwRDCgzy8t0y7cCJTk3n73KzrBhaBy
Ztd0OBbkpFznp4xavzCTF/BBoO9pb9dnCk/PyitrjkcLD6TszLET78YM2hHvm8cp
bCl7RxOFoxjYybeq1oXc/nQC14GOpwnZElebXW7YJja0C6YtLlBiXa5EhPvRYOKO
M4tfea8OerLDpOjPAPR2DTOxg/VzVUHwr7zpSx9g1TecK6Uwz9VG2IqcthiQSynr
2GQS6ABT+xdIjTyXGsvIeUPmQFP7E6umz1e2sZ2529vJjHVP/u75J+g7XkrJSAM8
bv4seFqCbbQGMZ9svg/Wgs4nRfOYpJ+Bpuqw+j9a3E2etiUlmujU1Yb7vOFGQBHS
3rge2m/6vMGYM2oJoyrl7YBDG0LnkvEi0gixD0+XB+pU84SLBmf5P0wN9dgBOvor
/dVfELoRAqqgg8CbVzWR3JrAkDpa9sn9LDPRy3UZhbAINMwDshcqhiqmzDxHm0sZ
j8vgeL/H1P7P9mjWWk9OKt6nmobGS1Hke3G74dfsDSdryslTHIHxqJ32wR6C7YtD
2dwdLPZzprSjb5Q95espDDy4lJPesDmdQ4FsKR0e/WdcCt3ViDwKxyl5qxRQC5TH
dgFWlNg9p/tKg7KT7X73+K3TTMPMq0136XUnBAzeG+5fZ747WqhU5Pw6cywXdoQV
UxqBau06KDIW9qhwZu0MKeweO9C51REPO9uMqqd/jNtRi3luOtM87yRfMbI2WmQ7
d1ixug5ye5YxE78rtrP3CjU7s8oeduDPvl28vTdU+7MB319Sct/wn1lmR1/kAsMf
pi94dOffni02+2jmYi1mHb97Ork1xHFXyCQxUkPPpj/Ly/s3nwOiBHQ+1W3yTt6t
RTlg2jHN+eSgTYbentNhTSBUAqvAF+HTOBmd3PHtVdmYcRkOG85SJJ2X8PHyybZQ
D9iV1xywZBkSQld/pyFBefp6h9PkXwtB0+bPbjqwZD+Y/a8zzsBTezJfAfYSLDIT
rfdtwqq4YzaAM7fJlCRHG2JIBzw6J/LnABzwOnav+v5OmoFICO98yq18FknzNeWH
YGkdJRWuib4DI/PouIbFsw8x5H9DBMpRO5ESQbU1Xq8XMMlcmw+XCofkRkAwn4ME
YKAR8YzloDz5hXt29rqPjZqrLMNyMNlT0ilLSJq70hPXBNBFih6Ch90E5Nahlo5Q
9PwZsukg666p+UoxUpLZQqhL2YibEJnyp+lp4DQ2WsGwmilRmughnqtMmG8fhy+J
BsM/XK6YnsJDs0xVBMf4NnfLOIsAfihP0+4Y0BGmzkLPacWGW3govSGKGIT9IZIP
sMUURBpX+GFwbd6IW4DvoauO5eOSNubGqcE+KuWjahOIaEFPREKZtgVr/Fs6ThyU
7zR9KQHwozSUp9dx6mUkJjY3/BxFB0agP6yAmC9AyOK6J7QB80tw/lNw0v5570Y4
uwrc1TOXabrJ1dt4CdiM1/91Mcrds5JGr+Y3j0/TdJjrxJwpvwLyfrsuE6zLXW/2
/at2XC5mhm8qNzyAPI0CoSowwOHj19Klwun0lRRxLsrNJm9CyqcNCicLhsg1IPs3
MvsPQmymyKrY9anYxvoBl8q2e5UZjwUy0KvRvdFz8W4twHuM8OjeFNkUagvS1zgb
jvBo+yNZg4Cyk735NiTE9nOXsE9JfAtw7fVnd1tlHmw53h1iox7dBqSIBY4tEPtQ
ImZc1JV16Zs8Xw92/UAcC09R/xKgx9eImZDJXFzSbn5sUpj6hGG0tUqNZ3l0c8UP
n2GtrGQVo6d3kTjPL3sbNn4+z77MSiF4MpTbYy1V+TBsVfcBdup0uZF/JY8x9kEd
bY4WJCweJq6vxfVbgOu0XoiYx4owpqrTuye78TcXlk6Og+iAvKGIB13bJF/Qe8Gl
ZBcrBL/2qVMpGPCeObg/hRI94uJW5WO6quOuNo05zSM0eX9ylYc/Iqam6YAxPfJC
NELZjVYj6TR66zfLPYYY5djtd+lfZR9GZ1iW9mRQgakjZ92rtK9ySDR6g/oHGgHS
Ni5f5mjeSXkrC3mBh5xvZG/a4AyxK8qBA5UW1u/ALNsCQQn/poEDnPelk1i5EIA+
3oXVi7cG+IED4Wgp4oModwSG94lL6I9Q6gRHL1wIND9BBO3VZg5X/lgi63ivVG8H
Eevyi9m0/AoCLuvdLR8obQIbP+gzSoOJ+M/w0tE1JKDspZKhBcPP2oCKtpMu4GaV
bm1u7zUv78XrNTP0GBHq8nqzDvJ3VGFKNjD0TzoyQ/CL/XSp9wR8MP/cXUSPvwHc
Gs4NV97lu53Uk5J/VAEQDn2qIFGyiKR3mNbWxK3zF08VrfHpEdVTAQ2IHALvB0oI
POF0VYbCmIUFHHNQS1Hr/Q6sHoHFEbDRwleHPCSTDjUgtdzAFlVegTZUuI1PuLeV
cw81zvl4dWphjPhUdoiwa7+U45OO7JyldDtUE+lj9p22L6+wVDw+2eAJnSvXMzgM
z1YXi03FzdbBespvrFJWp56qMtErn5B7E3AnhGtIE+5HgsrNq79qa/cX1si7qZa2
gbO8ZU0F+ePhR4se/VnIi7eze/qvKGPW73q8gPSK+KfSw9/SdHhTZS2csLwiiX6z
e52gyzEjxAKBeBhprycdVgMWLQPnkq/2HFjUlKfcIoh8qN0zV0DHYwsRIAdq3tVB
/AQi+sCYBz/+gr7FxurG+LlIWj1RK/g+tIFokCyQEfvrd102XMIGAi+NcaAbmMor
zDAuOCulsSjPifm6jXdAifeJv/7bmfYDl8KyirUgyWgM63nRL9P+mQ6LJsvNsPlD
8cdwUyJ+DAW4gFAKUNc6ezxpkGaqDHsywIL0k6enVijw8S+oJAnICn+FvnFFyarl
bVOp3kdFEPkP2NLvW5AkSD/vuXv3ZO9Ucomzvne8oweW0VCwe27lFvKSNEFBHHib
AnlnbRkd6zJrqshfHVLIKcUYLhgnW0OgSlghavK18BlWWGNz3gWYR+l0YxB6gk9G
u4BFOWL00sm7SuxLi+Q82Ns/7TXcDSkMyrQU12yRJXRL8POc6XBoW3Xznh+HJ1aD
pDkr59bpDiAjTx00wPiSjLL6Mqlre1On5vuomht6/U7S7lNBROlT7MoB0y2Fvy4e
MCdmGT7IM3Ewkv+fD0L15UB7yT+zuac8xDCtdC2/b5vKF9T9EVB4NSBuY47eFvvI
PcteZ7/B3WRlhteF29cp5YfVihusjbccSWWowmagNGJNKc0MLNzztceicFfWN+lB
+of3la1qR//BEFv7bKU+3tkCelVhBPVlw4XMxtlr1F70PqmlxDYoVfi3JPMcjGvZ
13OryRvE7pXD2rPNo/kqcW01bjRHgkMEsE+yuXx317eSdHhKUdGLQ6Z7YNjbEChM
xtV9kIxCNTYyP5yIJnBO9Z33lomGevxDCZAoUwFDZgLUfysW+m5vrE4tn0raUMy8
3Liqaaw2PDc35MzUnG17+eVVQaREXl0I9PQxPP5ngoapLJmvQecU65p2PMbAf+8x
FBziVOjoJz1qwcStetjnmTvasK9Lsjkn45lAINl6D/VOlBkcWkIdPN+PPuiUAdFi
RyVzG+W3qq0axlgstfAraDb3l72eE8QiGYI+6r3K3hBoRuV2qTv+Lomj4o7Nr4bQ
EKPUVexpihPI3PhnB0Nhn68lo8XxcUq0x/oRirABqaJ8V+//6WHRyGnCjEp9z8Ew
4es/1p/L89we9JfBYR02135Sf9dNY///x/5WQAHAPQ1Su/rWeJwLwN5hR9dxoDJ3
HAWAevq71ZX8hHKmflUY6kY/I9NQy2Idxw2xKPpw079QjvLn2edpUtJJZOc2kzpB
cAQJvtpWOdvDK7oLYUOxklkKVabn06I1vP92oX/Nfpkr0/Xhw3fmkfPMi8jPTmtd
XrgxIW5aY3MVaaunqo8DmNr26S1YIBYCSwr/D9yIF720Mzvd2/xUvcgGzG/lxVhP
gzNuBYzowoonnGuZ256Lbumc92C4v1ue67TD0OO2p58VX1a4e82zc2ZxuuzZmnOC
+8Y8tpjY9GRziaWItnCvczhNZ4RGpDEHL/2miImCsmqikmftqC7ZoK/abuITK7GZ
Ooa6wiFEEBByXsPO6mNmKeDwu7bb4knqHvmJT4lia+fIQ2gaVqCIfZOdwxMQJy/l
9tWWL+Glr+HYyZ0du3hHDGq06NvNvI4K0XYpaNgYG/u/Bmy3c6xHZYz2joLDlWpx
pO+wJsaOPb2WBkLsPSGHItbIko+XU3pbJyK5iVZpaBE9mrTZ3bF1WaLCUOnWh2E1
fVJ96fPn5bzCU23wuqS/WbsnkHwhBLOJwj2SPEmiHQaQoL77QqScIRYPKGQZyeti
gFZ3jUDJX9nsYznb/azWlKUSd1LSDyhhkzs9YfxGuXrWG9Hk85/kOKkwiPZiPTN3
casIoKGJjtWP0JrA2/i7VIk1WzGKZ94oaUSCiHFuG7bw42uNmGuUFU2uSo5MJSQN
0qFFPjbEmdx3Ne06mkQA77+PbKQVWN+oA8CTHeewGwjLCkPYDag3MJ9WF8OuXeRp
LQa8x5HB2Fov/EwXg8ysI7wdP+a+DAPez+Clw6KG6aEJfewgwADx2GL1fPzzkmq+
Bci+CZwxIgh9MiAMFyakjtqwx3BXfHgLcStDvhqmIc2RRDVgzE6j0VKBa6sRqnxg
Vu4GlWvBbvKc/GtRksFzqJRYd9pzRbu/sJIiAZGWtjRJy2Rju0a9/R9clm7enS99
t/pjfXr9qphxMXOEaD02K0HkWGbwRM0TKL9YUU8Sbk7+YYHX9yoLg25R9JOO5i57
z5bKAAjjHXgGd/xk0moVQiB+QcfmwqBs6DopsjZHMXEjvBfUPSmLoCsvgS23AIp5
ykzD7DQ+VBDSLeTYGVA6BMcngaA+K2HKncQOhSbZSRG5bAwlxyoAMw7Bl7zi/iJK
aD6zBpoPa9rKqtVuxYLA3DDukBcsT1B5+q5a07bW8L6F/MA3JboDLYpIkIafEzFk
R4SBpx1eLvgD0cUZIn+XMk6AhCgK9JduYLwp/XjQS3F0BRFgPcJcoPZ2CdUa79rK
r+wGYR028uCkBYb+mijZVMq+JPJnV1qEjrYjI4aGlI43fKkwP4n7VHWrbGpsUc7w
ufGsWlU1HSDMv2erKVRb+L0Zwka/gozaaForBKLcJ1esCR9ExwphAFsNgCj5uSY0
1cxxyNvIbgowqn13y5mNvudZj1ogCsRLC4ydoPJySLiizDdyoKGHSrofbuLzOi20
roVCPDos8ADjS52uhCIfzsPNeIEysDFG9Vy6WZDP6hbO6e+LihfehYdeUfcZriqC
/mcG88bbLcBcEZV1zJ9lRYLWFXVCt3AwZfH14sPgxydGLjDLg9I9Kg1P0dqApAMS
qWBBotIpkG53SLTu4hj1etPFoko5+tq3BzyjzClEAJ4uR2O11dehrbwtHlXYn7Eq
lr4rvoBbulcpCLpFelJH+FwPbtoy/olRCor8mK7ECp/CdC+ILENegFpAi6d2GI8v
x+x1szZSQ2397rEgWyzSDb2HQyGu7kxSKoAC0KScmM2eF/KnONVYdF8Mk86aLNyl
6SAYtSOG/z1d5k7jDhCRrNbqN3cFabfct9OeW3yycLG8Yo/pb6occfptPy51qGmx
Q0Xk1+52pAuwL2hbws7fki/COgChueoN7PVJ/QvlJqCJR2dhsUhUcz7Mp69EL9Fz
dRAVHaV64nr+nRTOqitn3rESpKKvpwgy3A/QalF6e2DJ/e/HltdZcrA+8RYtVtdE
YCVpLBNCB8F3y3K8u2Ib6+l//dUPhcMnGgVWm666eN8SDw69+YeBpL3S4Ov5Cfle
22vjn/eebSlY3WptT6ZV/WCCzXXSeZKqBN6diXYtMrWGoNmssQkUxc3oCyRYfOHT
s609EDaK3oZaiJ64QZIqXeZSwWP9/4aMKz8DpTLLK6aN25RYsm6+Wgv7J0RJ5l6M
mozRrQq4DhUps0R+Puof68cXA+8eo0ZTD64y6aBkobXlaxJP9bbL2s0lN3PJilLW
SBZZ1SKAJsofoHlvXEgepi+xuVbBARACP4zoSKKE/J1VHjqiWo/k86DjZQbr9R4r
aPvzc08v8X1WXHl8IrlR4mycXQAXiXx+CRKjGuP615WHfEL78Vc4rT9xcXEsn59u
SRDmTipsg11mxJLIRAW1HZP5MHK3IBYy7jX2ax3GwytwZewtIbdl4HtKPeNvazo6
Kj2Wk5xEYIV2HpXrt/UUfft5Qgtldj1oEDBD7Ktb28dUCMVMoPb0FASQjMSsl1uk
LP5h4mw/3phb/4r7e4aP1qAmQZQBrbfOAH1NnxoZycmVgWEKvoIjWTlLSJgzc7Iv
fcjI4h3XDI85iuvPGc17KZaXaXcMXuk5k7ZaT4I0lTUU/M1X6hADcOKSxPgfnfwt
iLxutnOdS+lv6H77OktJA/HmF+ROKiW6H5mSs6qrVLS8ghhsxLIKYOVk+F91eDT2
SYwv8Gr7wbK2B5+/f9ZeV9CTh0SEhkk0yWbuf3HbZRhbaUuVwdgcHxE5USYqZ/8a
acRM64lWyBfR/5hnLKRKM6OH5LgyrnIO/cX7FN6KDyLJmIYADkwQAEt3PafnYJA3
2ysUp39RIbRf4CCtaPgzSaI2tlXt1h1t7eq/h1QwkDOFmSekxzyKo8uxDQUe/UIj
n/lF0tsjCrN8EYdIenrKyHvfP36xcI+I82632iihfipB8o0hUuOIRueSZk2LFP4Z
DOoLxB4K/XaK8jhE8PTU2PlzbtkKFmxe1M3fQ1VhUjmpgNzaKv/MITTWLFQIxRLK
IoH04oiyiaVtiiHbEZzM/OKo6+tryiCCZkRPClSXfV/0zuMiOzsLqnzcYqHYduxb
rPbPvQLWYhAstXJLD6VSi+YBKhNnACFs7xNwiLlI9b+/s+xC4duKAX+tYxDO+z+F
Z8SJ2ccU5OeSzT0xyKMP7FtETuY0N3FKdp2u+QLCZwarWT6hkTzL8mT21bZzJziT
lDhDotMzZyhigsgkrYcETaUN108MUcu9V4TLb8bJfynFFkQNHruGnlNvhvxJVy2U
0VMUMpoulGdxyPcbRN4PMSwE2m2+BKuZ1HrH+bmGLufzn9l1WNU0h/10cfbwzqM2
AI0WFpcb6g8HAqGhbyj7xVg13OQGRPWMwSZRE+LQkZiM6SHOo/CORmQEq4mtykSW
6rdz1U4IUa5Sbboi3qz22gGBIdX0p+ipnypUabZBptCpS2P0i6VLcKvLrjnS1w5g
AnLiIJaQsr5pEyWKfIzwWA4uwc91Ua18yegHimKiePcR2RQy3/cnfqWtswcyiQjT
fpsUEz4bi7GlYtG+HlDy5fKSuyD2iaXZMD8xjDZS3pGwqO3/ERM/sPuty9WhqUaJ
nHskDreQAQSgOKLOVSKNV2xayY4Eoixw9brh6v/g/ztAEo3A9bK1s4kj3ug8Yzu3
S44+pNVmesrvtxYmuMV12CVwZ9SytsGIoZpFRGV1wpa9OnmuKrbkQJCgmFK+X3I5
r28C6HIzaofuZthoXSS8XuWFhAj4V0RfcnqFOIXoftEwzXAzRx26dmWD8LVMcClw
CxZWA+tsJy+PbVtQtq98TK2oEVjC+OOJaQio//FK7Es1jWWVNezvRDaSILF1oT9x
F/ybFu5rGxEaehs9eJAlfEjhJrQgX0dx4FvNjSdT303BKqDeVwCOfP9Qqulj7qY8
4XAUsSv7lgOJKYyeBEPoyok9Qe81YtuuaEmUkwjEcp9bsD3y5U3cNnmV6COKGTrG
7T7wzm7+kvZQC0Ob5RAcCwguKPNOu7uY/Iyx58zOz5vTtbsXqGk2Fc1kdxdFNZ23
5uFBm9PaCue1MZlfD8WAopAn04gkNxaukFAObGRfIpRjzA2/7F9IJvgkqNubsS2R
Xn0YCrgVdJGdpWXOg06bK+a4wIzIRPwZ9JygS/AdLCJiM0IyPmC+jqE507l0UYsY
jolGu7pmLNpIhawyt6ZvukD6zVUrDtZWy3erKlq5OqOidGO+/pT1BqAk0iSHtg7P
qhzzSqAR5Zp7Ndz91iy1dClEZTreleCeJ7lVyfrrjJ13Jrg9CHGs2lgAUk7lP5dg
Zocfb7erHLbPha/XAI469YvXx2NZ6LWjgQ5acVHXqEkTpKX0H7IfhG9YBF+tnLsq
U0R6uTIevLPtUqkGUD98TvmmvElmSIyAx7R/aUpnA1cs3Tny+LM7WEkmEtPeEUqe
X10bdiSfdgC9Na2c3/Q5evjdTLzTJWzdiG3uoEj13NdfC5F9qLJ7Q0aqx39YIeJr
zuqOKfaQmuW/UpOsJISAzb/CXAckTeKydvOo47qcBCB/VOOOT4hFyJiet8KRP7DQ
qqyZjczmNA6ouZ0/xfmCNtxBhSTMN7tBu7yZN8cKLjCiPeM1L9KfpTj20kiXJHdb
pJXGpLlkfpg4U6XUEq2Ic26h4gjO8euXsaq3d0Xs0AqR89biA6NWMTSWXFQ8Oddr
3Abs4/cvpWHoN80ONKI4o/1TccF+1fkt76rB/QLYR01fy3a2QLFYHZiMsu3XPngi
UelDQ4karUI97Tehc4lCfBSQJMtNNa8j9zgqPrsbyioqwYaD7mCTrA+mSH6PKKp7
LvwbDnfvwsnRdCKDRLM590HOURYM7tVEzILVNtuKRrD3uxlF0HEDSbExTTFaiyb2
ve2LTcmN37SLbNzvbBdq2xJi0On6lbIV4oW7kq/DTCsxtD29idceW12v8FUhrKpX
HVzNH7M8npbbBygLje8beMc2xEjK0bzAUvbuiSk7DndOeQWeuFedESIxWfj/KT9h
XR5vKW18PJeC0x7kAA8c7qUtNfQaknmjYJi8zAJ9RSp03jLSnmRUwzQ6m4SADH68
JAzb0lMIFWzBf/fhyauAlVXV/4yj2keZaC1zbjka3KrIqp8pndD1WAVbuap6z5Op
JjN8hHJc/FGCq5bePjswNF8VZD0363Z9Ydu/L1lxnnDQ00NhQ1iyFK4HSaj5Vb58
fKa4cnlSw4aAbn3y5ZBeJ4WheAN1z4y30rRwOfPzDQDM4ejBDk/2qLt7Yk/FwSeB
TzuUDTuY+hRW4QSVJGhmgvERk15ZT4jqefwm6ix/UlJSc7aEx15GX9jwyVZmDjsU
K63fXNd56gFkKFJdIEUgLciIoLH5RNtqQ0rb/TArh1UOKXE6YGTEuVYIAeQjWkw8
irIgMtXVFAE+iLEz+p43JE1MN1vkjqtw4mQMyK+wuadOBzow1oBZXmJ9cYvCv+5s
PNSPxSC5d6oyGv5K2tQ+cLdFZT9U5WDKpyNFYuJNjvBowphf0DGRD5KHlZkKNRsV
Bpk4swPMIkQYV94QEY/jQ+LJd1d3ELp4LG9XvQ2czWKOalZlF/TcMnnQ79fGKSM1
LXoIuViWUiDrGLggxDacBsXDo12oR5Z0qjgY/inyB+OXogUaULz5MjVr9W1qhnq0
U5Gh6UkU5OPar+Iu/7msxaIiSZyy8sHpYw777RrCDHukY4ruqydkXrPRGaFWpW47
vds+40GGXtPMZKfkz/uF9xlKHuzT4IzG4MHskgg6UhUsxbAZUGDllalmArHRnVve
xUmzP0/EUDg6nYVXI4HNeMN7slFTXZswmKUoriM67/zep0Q7paj04kqH8ccXVnJl
TG+BbB6oy2S40+IpIjkp29xCdzcuubsEW/3Nf1Q3JA9r5EAwvrX+lD6lcUaY1oE7
bEIVwAdMJK5+Vpj1aOE7mhPsyMtz/sPs2aX3q2PQ3/Cqrzzfw6VahST2F/ueR6HF
Cuem8p0DJSU1fa8sHrbhQXFjrhVZeOUURxGN+w+oR+lHnQa5uHSqZYfM1L3jm6th
vo3nPZ8e0wCRsDdZ9JC4NxhuZsQkXgs1X20EF6d091PIQBEwOsuOodtJgjX/gTSc
PmIa0FxeDglqGO0aaOSvPRYWWdfI93J8GAksvDpffASnwPZpSmNryZN26lOQYWMX
ey09JaKrwkMlGVxEMDxn4DK9jvUsxzBB15ah2TOigkTAWa/Wot18+ivBcgj0hAio
oQNBF5CBk/4+K+AYIqHYuAjaczHQ7qHbw68IOBHKfNw2X9Y1bvHCj65vULnDPzdU
2DTKIvzGCSM1lCP0biECfiTNks6EexMMIOziikBbH2ShX0UmwvGsg/TEa+WdHXYx
OGavApgk2LfErwbg8bqf8bE14DT7LkKGBX3M7pZIC7DENb3hf2AV2PXXSHMzPZcA
qCQj/7SkcxQgsLDSjMEn+5rMOEeo4xXrU/bGt1uDNm+a08L0B+IZKFtd1h3/95an
vQQoio/uVRBfiUuZcujUlOn45p71PoRelkGn8tGv9EwL/Lmg4LgJDWsG8lbREI4d
wVMhTpkZmWtPxeAvzHwe+RWUxnpXz45QBWDxij5Wt9S10BXiZnbAc2/MzKI6od6z
Z+eG3tm2kXdEMRYTSRkQq45cvsUz9CcqMPixNg1sIjn6bN7CktBj3PpUtY+aX5Zq
vSGipuVIpRyQT8pqp0vrrYM+/BNAb3s5/1OchyGsRIoY/mJXx9mkWyseozzjQFSd
WBN1mZSIENcIjlFjGDmS/VT7c5ua4m9jo5nz7p/CFc9yuAI4c/zQlXj0anJWMYBK
yttbgCNSg7aDLyxnKd9kIqJhx6ioqOEakbbjouEF+Nix8soYC1aMy53+So60+LdL
+2xcy8FDiO3s3SJ8eg0lT44lcudwYDQ9x7HHt06ycpfxwmA14RLiQNdplwLX9zLV
u6xFduJsSJSZviklYFs0Ds8Oluz5tuWHLN4/uGtGAj8PI+nj0xqbeuP/OOgsQap8
xQ8WbWWOvfKIG8Lrs4+tTK4EtC9aQ/za1ZiES8MkdCOPFD4s8gCFkpemf1GmrTv5
yttk/zUG7RrEskXS4EUskzB5PNJCpbBKY2IGbNwSiVMUvxUta6k9fU2Z16ICjKml
wCUbTJn/OzWK4BZHMxst+EJMpOx3WWtQWZ/PnBN98696IdBqnzNyJbbht70y0Jlt
CSMVE7Pi19nV63C+Rnb7WyD/ge0i6VxEbkdm8vg0rYkk67cHdV1HX6PX005ZUnXS
3lwvRkRNyPInnJX+iKbNZVXKemqgyCaf91v2BcwEuAD5uClCkCdyugu1rtk1DjYB
IhP70AqAjkjPvbUlL1qllGletta9/wHWq3Ddde96sPk9ixKQWX2fnAKWizgcno86
TTgEN9cuEhUMgCKjla4/lGJcz4po4YnPghlTe15QLUM3dAS+fib4SkzLubbszXxR
0cwaPdBoLCC74ufoPjE55axV3fuJXR1jd1EdrPHf89/E6QJXZZmDKpCI5W68WvTy
LG1jYj5cl3j1rMCJWhTDJVhA1ImCB/HcdVJtQVaWPDxTGAtLvJyV/86NyMfV3zkV
+OGGdWVb0pMIJW/xo8aL8v/SYK41/jFjzNmeqj6aFN9FAftabJKef582uE6Pf4pN
PwvfRneXS017OwoJaSlD+WXU9u/oIFGSHvA8qr5D3qX+GNoao2u1I4DSi3IDZIZc
3f1eG2tT7d0fJwNHOTPMrNDWfoSvpk3WAmQi+9cbwBt0Rx+b0GSu50Q2eGX3MFDR
OgWNuCJfl/ATplmTuzNcxX1bpdQzQuYrIZReKAxnMemKYxIEbD0eKbQpzGnyVgdA
2Ci7P+JzHG8w1DTBLOpnYWcTb2lJhHTOOjmjJUNxhoMGwoWXE/nmpuggXDhlemxH
BatuDKG/pnkCZcjKT/rwF98NpXkjIxQjn/9+p9oi6zxLReONrTqj2oRKpvk9k0A3
Ry+SK9Zlg+z1gdVtJY3sQ7Fk6TtSGRN2Cs2NbgHpholudYeJRIzC47asTMT620TV
lDsy8maidqaRqVHRDR/gxLVTTqOVMBYLW+OXr4/Q1zyrwP3SRcVxGp3o6vR1ki9V
8iFLuXkGIupXm7719c29m0oPyiliv/vOLKT+OFl51kKLr2HhrGAqhlt72TM5Yu5J
4YIdxodbiMM3KRDravdcbj1jBlL1rDzFLXhh9AJH84OmYV9mm38mBXk8t/kzLFzE
fMCBEOJPor0+o8VKXpIpU6IHBbX7xcqsUw+3goj8+v7KWM+eR5vWYebKSQ3oZtBn
u8uj4WT3uq3MxdJKfmZZNaXmyIBcki/PHCh7zydXCqFCMLrlLENUHCf1grSbF68y
bVqzV87hIO2weE/WJAKLE0aA0bVkjM0uQyyim19ly3G3+ECJeYgYMnR5Mxwjbtz+
AqjLELITyRXPHwxCjNB+/AborSJcZWhA6BEbUwhVVrZR7MA15LMC+kUznXPOEhp4
qYiZrxoKHctk/kAkhAlF2Kjmuw/wRW5jZVGaunnGNXvsubpvTNEzhB6eunTi/aYg
S3lzBtPv5gbmV3Dt+YPdRX0+mP5IlmlaIIQ9imtKqU+FctUrZv/zeHyui5Gp0KqQ
v8U2NAQGugk4D7tRkURkkshVdvFNYd0jKrK0qX8tEX1rjm2jPddWBh3CnQOSNOf9
PhvOw6Mn1qSDTNWPuXhRRVCxJPdrY/S5YACnknJo3rJzj/dHGh0Ipomyob9KMGB/
lsLuvbYytG7fNOZkTcOM9VJLajAB9j1ovNvIVuDysnpR1QAme6NImGS9P8qON482
P9CgHF3zgyVpS8qwhZnf1tmHijAhvfUbH99AxpGcZFR3/Kt/chcdtOPycygNH72Y
QZkqSPfQfoa4inaM3cKH4CD8CPAj7ZiRZO2zEK1/bkBBW1AwPnp0nYovzUDpno+5
SqR8OQY069KgFPTbu6zrN2Biw326eHpD8qhLGsZEuhTUdzO7eieJaLVJzFvNQUCB
McbbcKDQnW7xJQez0nncqWtTX6E84eQ7tWWAEDQU8kh0ZouLH92MJRRZsjLGVPCl
F11zKyNSiuAPh/2H07/nz9ucsU6nuLC7h5OT2Nr6RzzlBSKiM3nUJjG4IyKFJiju
Aa+QaQ6BlRa5AscLsjpwQsK0fKfWqqi5FN6f8WgmbGG7HDR56KYLGwi0bD0FkzG/
8cjWDHww5oZ0Tx0UnNums/5xfBmTecfogXGwNy0pHmioYuEIWm0gFNaXu07Cv8ba
+sPsFTKLAtG33fsR9QuUMm9VVwPlmvVD/HZM6TQQNu8NNXkifAtjyS2yZyBIbmRO
wczkokhQR2dchir8bYhIReLSmB0c0kC/bIKfFyGi/7B4AjvYnFEoKJW6MU0vhv5A
YeXJFyLLrIrmCca1bOd9Pf1HTLbeKgSXLNpk1oegGS9qyAmW/bbP0mpTxXJLIJu7
ItU+NjOXnj00qBRIT2+S/E1Ze2apS4Xrs5xhVwfLS/seX5QuykIqvprFe26PPtcq
RFCem6d/Ec9pLqwl7SNPUiOIyQRTREr20OlkmwejeDq7in8xqyUvnHARJib8R9tf
PNTYIoR6CgxyhTyJyYV9rkdu1wbcWUuK8K17Z2kZCqVT4xaWMGiQnr9e8kWIUWuZ
KB5RUIjdrcorm/fDJc7cJ/Hle/Wby40Ic1iSdS94j4PMNbjzG2TmdxNfvipZuE0E
tHAey200j11sxC7NqVmzcIrzwTPNrAxJKt+HIH5HPbkxfxwrfdkBYFLwVBnqiBHz
Eq8IxR60pxc/V2Bk67dv9KOBziD6gGwcOHQViAnDWA1uD7gt+pufxI72SO6991pR
ik9d8WZv6q6hsVKz44pTlsqeeL1pjYDK6bov1qhArFXbJ798vpFaQ41C6nNAHaEb
K2MpxhwoPq+MBJA7e+BRKcf0yLBHA3O09I/6SNha5BivTbMprqd1IPXhwL81380p
tSNwRLlTL4CDBOfb5WDQFO8xTactk4+JDRvbCE49J8xQzByxE8/tMKr27Xpz25yF
6qFH6+66dfELSdijL/QTbVqTUbgDvmFxIcZS3PE2/BKAvwdFxpqsnbNahlTXBeK1
c64kepNt5ha/YALF2BZvzfrWWZHNL53dN5yITueTcTHjfQ9foZxPyTldJWxRq7zC
+P/WWU/C8eVwWe0XwqQKz6mGY/ZlSdfSdP4p1WdFnApLsBj87bnegB32mLctHNYO
Zw8IbfZ2YTMpXbq8H1/tyBjsDMRDu2lpeDmwgGpHiYEdVNzvNqaOWM+QcoHwykPN
JdoKkC1QbpdTHcMuM4bUog36oeDnH/YorT2z+HE5M7tpmIPgc+LBpr38oNZwBJit
BJe1KkW8hbo+Ox+DaMbLGI7wzsvIF1zIiqqCB4gCa2dVMF58CwS6tu1gUKZS75yS
BaIS286TJIeslCdaSErwvi37h7vZIjAqB7oHgCgECAH6fDzX+Z7p2i7dP6y+UBXz
LWlJl6zE3F6TqbC8/eVXNni3qPwtCL1p2uxgx1IqROeF8ahI77DT83Adm2KnP8BW
JuaH2PPsiSJDUav8KUz1s1mOnoZd1uZMgOVWMko8Yt44WY40sE+7+PlLMPEsjXeZ
ngQt/Z74R6R42TOB2Le2fEUTYfBk13SAotlPp7TuApLliiZZ7Q6hOhCIxMNvOfnz
ilTtPcVdLAdxQ7oUuqb0nvE5YnSfhv1fWPeai9A/xd3WnyQJPcPiM4XLOZ3osz1J
bzTpGR0+KLHNoHkS/EuhsGQ/IDfG1qSBWBoHou6VqtDkxIf46XRGokpZ3zdBj6pe
GJplsZOad7YWh/CU1ZlBiOnImhQOHTKy32gBSV87tVTykSkYDOEoVaYbDL/CScvX
Lh622ILbOc+azfIokz1NcC9TEYFVvu4l2qa5D/u6UiWxtmGLVMCJI2EGQfbXzRKL
em3qtP7rDElta75sBlKqbrmbuLFaWdTcYazxOt4Bs2BkybUUg+PEWQKehtfJ1fHB
nTUr8vGSqKeoLDwmlNAA/XyXODIciTlr8Xefu9LrbXXdQjd7ChBBCjA088glNKMK
6R7LTzKMDA5abmDXhVL1xs9NN/zvpv8068pwWk+8dw7NEx1Z+OabEvUuog75Hyfa
pTj8hBff+O7zt3+zbgMx8r9lkkf91CAzDHFrxthuZ9c7mGC0atk4IyMofXHPLy6g
2MP62PIhmrOoJBixGjrNCPftl4w7Id4jmCFPvnnJXVqLQBlda3nNxErz8CbmbX/o
sY8k5wEbRm1zy4cjXzBtE4jhmlgp06ENDDw1LYQC9VhTMq2hvucoBwwrpsDeL+bs
Csz2O7pjV2Xxwath+d4jd1m/P/XyjDptRD0B3AeJTPOT/OHIaBnZOmiIkpfuqudN
TLhUdiD7KR2o6yM+mUzB0SSgXx/RNCQFrwrLbtH3AXQdxEgsrNf6DGBrIL/M00/x
Hl2jogF3OcbP3VNhzH5x7SPa8A6iwJKHq6SNow6YVQkeKD/jPeHuUedZuroPWjuq
h+ZTuKA415XzRXw/08MgCeCc8CXNCTJ6RtO6/JnGKaDMcz0ar8kfsB4k8ovfhxCN
c4NXJEBRTEK98DqAO3PjVCVMaSyLjAoiXVthYzq2c+KzCCR4+io1zU94z/6cam9L
McwqSy0Me4D+RpjXcGDfNfTNEgv0Rw7n2Sq+VnDzmnbjNzga6WOhS0d1c+9VfvPr
XD9/+/PbdsnEmSuBp9GCCPIfNbQUmV80QYMq/+ShEu1uV0E/TXRaL/c0SkE/n+sq
eDpquK9QGOaQsDkcTlFrAnJVpg6SeTeGEb/ea5JMEFlpjMDqYdwuNGmGvP3DW9dX
i8MktqWX9SULc9i0ceU7KBe5Y49NLv/JjqPHJ4x21sCeLTsHKGEKE+Rsfr5jSd1S
xCpu5h84nu0jt1gXT0j0pIPn7lknFzsbm5zisFQLy162cAVSM9Ah6x2r5BQwIw8c
4Ni9Y9MN+7zoDpxX2tswN810t+Gxn1WJBujzR6IKhS34PgDTfoblEa8+MTXTARRS
5Ig4lP/LyifKib3Bf3L7BJ+uggawCH8KQUGT17bm0q4ImwRforCrENT8WDHewp/v
IyxQe3Fx1o3ei7F6v14gdWexLmvxKCbE4weZSAuyfGSv6BsL/xd0tjz4qeXltUvE
jsK1RJeg8H4rLIThoXvBckqvRF7HsEZ0B+mR7DncGthJR/YP6XsNm57A7dHumkoY
aBuqsxT5BLmVYWpFoqimjDGHGQAV28FXvrk8VVpCxWwwTwF0gix7xeOJzwrOpvt0
CGx/E/6gdB4swOfsdA4+K/6doTI7tRomKiZSrpeYFGGPbo0Z/+/o4PiCPzHlmgBH
Wn7q2gAuB3nVmwVL6mKKMsSNBpYYcjowk+0rA4zVNRRBuP2AhMVv8e9r68MmcfA2
5mAMTiUSeRzrdpcbqQPztachmuQiPWTVvgl4xwRZCN5XMADAQ0CPjP7U6ryuPqeO
k8CTcr7jqpER9IzQ5oWt6goa2/4ynEgODuwUtPnxEEhhy3dxQ/h0nwv6ByBlS3RU
oL4IlXqzcJ/KIcZXY2uo0FH9ResqDrB0FWWHduzOQwb7NdmUtMp0BKraVlMzoGeU
OMMrrh6fNphr0gUpHg9G5ywiR/vrEunXbMpBIiR6cDejdkSSJwCI/Kokt7Zjsp28
yUwvIv2xwcPbFWkBGlR1ieZPkzEjDoIhoBk9YYOWrO1vZpCMhGucF52it23sJxKI
8nt/5EKG8p2S9VbCDHCA0fV4F1RP3xvfbw1y8Js1gjBLvkVigx+ti7E22VibRcJg
7Vhb79uYaBnpKpl3pmmU7ZnF5iRcWb6YyE62a6ZUhAHriyh7VoxiTUaser3n1GUz
bLStAG5U6HwKN7Cxx/N/pZ0k4qvwOJmkeBJ3efwFfxDjbydHdAiiyYlCfJyLda3i
yjH0PfGbQc4lu/uopMBLdd4NMh9BhUYpx1o/VVicyeXn9UxMLAYZE/llB1zZ5ErP
VSNYxCTQJTJQi14Gn6hOi3lJ3Qzzb11llh1YHr5smqceuj4tD4Bsg0C83lYTvWVq
l4RIVJx0ZFtS1w5av7yo6qTbd0YNJNpPufJNZsGa7+AauK3MvA9K/IH5fl03yD+M
D0mWuwtD/0KDvtKahw52Ax98b/JV2NGBoz6wVl+IYYqZTWCygcNVBXbnH5ide3MW
bx2pBUKqRyF9WyUrb+g9ZWxrrJeMzJNtUFCSH3tFgeXnd3h0bWqvIole0eFR5bRS
IcG/Joklk/bF8YvEnE777tO1FX4GV9YB8FHlvmnn1kMpp3cCsdR4JRlqRoiEklH3
PL2tnnw8FGhEcou+hF5AcAOP4rSW7v9YS+bDugtsVybgbg34PD2zmDg8gNRpXiLU
DMk5/pyEnkaUUvRyAyG0pqasGltQaBq582gjC3PJukJZAFbmkhD3K8hq4UWjlhDD
rlJUPAdlu/yJOwTq1ZVZZygD2d5jWPoB3NGrIUQ176v8DfLkUSvr/RAtb0yzFr4G
J5FdBoyAGshNW4qkkuUs5KT8uwTMSMTJJ5p687vVR0eFPVD1pgO/BsS1TK4PFwli
Xcu5QBiSTE8VkD5MSbxkZzofuQAUPPzZuufrYrX9Ch1x5JDcWij48vrjujJFm4cb
F+eRpvLQ64wsnUAGXaJimjMLoqJdA0LY0YsshFONeT5+dZE6PysEcHhdv6Z4uGI+
tk5ICu9R05vwsVxO+5zaML8SwVn4pYdPliJulMyUn2VFC6AL3EOasApqMkfDCRKS
2GpnHVeWhkZxfRatGGbxia2kws8kvri/LP7T2duLLIC0lsara2JKvlZeT4C15j+0
TMF7ZxyCdLOOfjLL4OAKeTYWZQ0me2fCxaFeNYHvGlHe702ks0qsIrWdYTZOJv8p
rXZk5h2w+pO8Uky8ovP++LgFT/1X4UTGmo5EymI+8x6hrx/AXdasyVvMvUkPKAad
XHifvciJE/zzZtBIAXF8bjyWIuvOknJsVa84nUOmmEulFFZVE6MmrtSYCklEJsxu
ygVYZ8vPtHvUsEfU4okhTw5HSGgDJhG2QHfhlExYk6TbZJCNxqZudOMUc+T+9Qh7
Xr8kTHCz+GHWeVw235CwwTQDGCgaBa0Lbl2yArjis+aJCMztBQE/j+PW26aQ+Yxn
/shmOVPAn5Tx5Z4tkDMMIFSgx/WQK8tvYL5S8lT/xb0e4sknb2zD38+VxWf7L/Ia
Ln6QBaJw865c6Qt3gBs8PXkuMlomg8zR2bNxJ3Y1GwWMMJhTSx2ZUBqGDMcEjCCZ
DhIKtX28JwXQqRFXdAzIq2sFzzAaRpnZib63kZclQkkftJg7y8X1ix9sA8AxVGLa
LFbkFKWybWi2lzSEbyiEhake2md40fD5oDBPJcMtitsvi+/xRME0RHIDeGH2u+To
gaMled4NoA6JZqo/DivKzDZXVVnuwXX6IW9DdL4IAObxPsQzTr2C16+UF/RNRqeW
2njynYZ43PNrJNP0fYtdOrSv+khrbXCJCqqGjE0LZMeSKbfN05Kr4ooc45MsugM9
aEXpB9b69f5Bnf/hvFrS2PsAiaLVZZPCkJg64MPSpBCKyFJTNlYELFLs2IAzmyTf
vPm2iI4M0iTnLnjsp+KH6nyhuJm1jGZI0cbX6/xJKcwoapcjZOOCMm1boihAAGUz
w+ZLY6cwK5RMaewXrb9UfdXSqIQrzsyaYOpEX59E+HK4n4Y4K9UPgCKWRwOKGXaT
EDfAq+uuictoQXYvvurfkxVjaLKmAckfw4im0MwM/MlnZy1jVJDsIEJkLjkh8mKP
768w799vqG77oCwZD4GavtjonW5CvWXNjHi196iTv/JZMi+d/H6zZ+1HqeS6KpaK
O0AQBxqNJ5nGoqQxOBKTpcpsIfhHoUCsoq6y/cIvOaZt25gctwldNZlCaKSA552Q
4i6Ny5xLdxzEap4cQZn9DvnfDlFjB8068jHKkMu3EOW7+GU1CNRJP54tEiecA+AM
+V8pys1s0bYzdiqjVYTJlYUePgtFoUgHsBRWnKCMtcCkrgDNXAGfCo8VMKg1s0CX
FUt6mWRLOaEz1Z6L5TxZG0bMBIrfo9R4lzf/xmcUo0ZDnrNDk64fr7LslMm39eHm
2K24U7fUXEFSEC4hzozW2kdM+Op5Wr1PEMi62GVkL/ndwf2bVTVzGAPwqycV5VEP
W1Q7oIl11oXnBZ9WMJ8ani2n+dZs15hY2OcMu7kj+sPlwTAmZdXpDXRoeK5ULTR1
WPrdCPXMpfDfqOdwFpbLW8JiXg4NEmXxS9Nqz8PLR48kgYkpDj3onKyMh+4CJ7xf
6vfZnhe42dkW8sozqggkEaZJFbtId+Batgl58jJxnn5EUkvvv5enOT6392qe/ayy
Vu1KyUy2wJtTOmpKKVqQIQE8+f12jyZK/Mu6ZYzeQe4AYOfb11qgiQ0TrTG87L4l
t1sSJLVJ4lko6yPktoiwC2/Mg+coxNahLY7+9biZqOCFqxE1kDCDzPMK4JAz2i7H
rgzic/895X5AwgSkdBAwwl/M3TYPY9ck5nPO4cTFbLAo1c+rvl7hWLua5mPLmiBF
3jm2M6ecrurdsMtjFV9hs3iWgHFf89+Tf+HLBy1dICsyBjbfrtkL0gmfOs3reiPX
SYkucG1yAKWwktb/U3Xer3JWiz2cbj7WrSFL+2KqUQ1NqN85hjUQDA2KPN7ZrdLN
pareUHhOZIlT7+lqo2tx1Rudyf0BGgHGFTR+SGCRemynSGt5E8li39FSJAwZJR4A
MarS/w81blwPhawKZ3/jDBHKQ6WV17UfvlRJbNmvLm5D5Q4AhquJIb64rsNDY7AX
BjqQgzOJ004VwpbfVjvbs7TCmuCqEXncqe3tWh97FtB160BPa6ejxsfI10RSU50o
yWmIh1/EwrjrnSA/hAfkKQQgP0Ksi2EESIwyhjZp9yZEebD73M5dOxEaO/KlDph+
jYyfMjjdapw+PEtNKApwTuRrkLouOjXNp2bsI/I5td8HsERZ5BlreGK2EnBj8HRC
vdOqQzHKSCLn7+hW7xGtDNQ7yFNmdCuuG36CFM5ST5EX3Bwo7/8Ub+P+NbXpF3nq
kAghVzqGLIMbuvz4Zlmvj8ImD4Zfye3XSDjYtSlMbMc3fWIrVPTQzP3bz+pEsip9
qm5ziYfWEnxJQSJt/rG/rsLdzhlOtt4yfOSUd6zjjFVo9EOuLCtahF4Lfzx47PvO
6wa6Xx7Lp/Refgm+5hXQ1Bw0GRfTB04+w74MxHp8DnHhax46ppW736dbNrDKGBxy
JorXLS9V4+FQ/7xKZSDRcqolwtAPo3fSHo9k9fMohYKXkD5m0KVFVe1w8VVaULWV
2wkz3RgJnv/QxuQelA+X9mm0uMy0VALJKwO+wfJ3BPALwd/Abm1nOHONVeezZDHT
9YCG1rMp3oFNuc4pgrtTb+Wo9gV2goaC4Ye32A7TzjdmEUTMyOfcl/Cf7Yt/ozj1
JLJFQFiEaIEdhQAZnM1uXOQRPRom1xiGWWjy8o+pCpARHQjfGo5c2+NkP7vokW0H
8OUa3exPqbYKbk4EmMMLQkbZ2t5Z4GBznS3tUu83JmboY1J7Vo2NtYzrsgUHs80S
NRswts3bkxZSbGha7+XkSmCIl2CBTo2C1xSdfGTs9yCeQeUCjTUjfkyxOq8V18b0
wVY8rmH4lEjCnlthNBi4XilfmA4q8uq+tOpTlgOs1dTwiDfdjlzfYitDhHlmu8qC
0Ohsqq2okZn2D7B8W4J1YHa5/ihEOTKTiHwUchbwP4ue9AVg26qGlxcaE3AumepB
hl8cdFJ72BiS6qzExKklFv907Mza1sXG09GNazIUUMb0DG+y73J2KuS1DrTAq14n
fro50VB454mxMenYooTbhkruTv/h4lPJVl72ymjDk3/ghgmhiOCQ+qcwMdE8FQd+
UD+7GSr9QBs/dg+4twF6tD3EMI5p95oMcacE6qC46KFv4BX86joreTNx8rgvwElE
6nKE3z/awjOwNl4JlPBvSENDjyug8SwS4rJ6o7YhKiVuqp0L8Qoko2AK5DXmFLv7
Sww5hAFGde8jqZnNRAGA+sa2qS/1QM9UzJy5cEPddw9zmxEopmOAuhsTGtdSMuV+
ZfMUZSCzJtuPKwjCSPz8fyEQulKqwKyZipZkJT8TnTZAygWIzkEnKr8kTX45AHCt
308uchl1BuKvMdmzYTsQX9cZZcGHSppRsyDeRrXvOelGXRjYXizVpQhQeXPHw3y0
x9HMNrKpr6CjCHiDmebLFQlD4O4XMIq4l+B4PZguAwNMAR+HKXB6Nqmez01OsC0a
xM/pHSiUKYWPf4iLuZAkBP2I50NwJxyn0pvQlVvDt/EmXgHECnqEgMKvG7Fnyssf
LoiRu1t+XqxacmzlcSzZrYf93gkylKxt+/0ZbjwI5j5Wd+iAn2Hai2QJY7W5IUMV
0IncCQz2UpW9av0V2S8zXOvilUfXXPJKmn2XDpxNVCzZ2NFbUU5TIISVD5rEwiVU
wazqOzueQ/6A29XOhTwp3z7fu2Am7KkcUyvBKT8l/uUXQUqeEjogjvna1Lvw8ZX1
Kpzw98KtWJ+MuxJB9wMgBtxNeFWK9BqLc6tb0qiItXveEY2KoNJDxT2M4lC17Iu8
nSQkQE6sNWxftRMycEctrEkqvyhW2RdJ1LaEcwiSNHY0XHqf5AkUowb0lqeCqKOj
wueo7dZVxcLJPVPDLRBku5fTIrY1TQHo/BnqwrMqlcPKbz0msyg9tYjWb8fJA+pa
2MAi5GVVwQVjHuh6JOl5Ub5KFw+R2NJLPyEF2oeVvZSpwF4kuAlg7SNhIldRorn5
W2E3dp6pt5I5ICNnD2E7tJWfAH2ZEVEftnIYkBS990jtQgWoGfFaUiC4+wzZWNe/
gvZWvcVQ1foD02FkNd1EaWagzrCUKn3qzn3yxqqQ/Od9mXZVIvhDda0nNLOmCtDK
wOwl1lySmzX73Qbcf1YSVfJQK4RdhaPP+mWh/VL7ANb5LAwfk1kwyhBAbxFFcZ5X
wnwE4EYON8ZDnnzYi7zT4Lxj9tVd1YfbAQN4MTWJNV3w1EhVZpIf6Km20Qg0ETqB
eyCcKeLJ54rgQRt/lIzoKi3bSMDJOhXvyeMo4gEOBzViZI2IGtAeGjKdvmXIdxmd
kDheU1B5DDMeazlWtJw26ErYzgY+KNnf3ozk00aUsHgVjsvrbmn/YTsBGFgkgwT3
Bg9VLs7c0+zJ1tvzaqrqwJjGwtmsbC0FMb3r6XeVNcTubYr5T9/dtshNxhzOQ2Aa
+w6GlhK+T65VTGLqyGTUH7+0QD3WtgfTd/TjzQTyyNFwa4DMIJImyVdlsneeeq1j
Nd37Sras4J4XTRQpLZCr5xaSrN19s/uymmSPRjiU2tQApxZEuxzjU0/KVbDbOmFG
shc6c5RxvbqTq335a8TUUgN6AuDu5XC7sS4bQblTtQEu2tHemeXuTDMTogc1jLc0
UCzgqIjqFx1UKclxYBoLrM1+QeuHhQ4ZH4LP0zwj4gSwwObApSIoBbSOs1VERFjq
nDV6OObDuoXRAhMMokKpmaZiJGwSkAP3iKprYrLGyuoUVQVGgpaVJc3Gh0R+KFNM
2UQZXszagf9ftYHNwzZ+gI/puOKzZ8rLSRcl60SAHj+qmYM+tOfrIEFK68PNg6rM
bt+1ppOG95vU7ffcUeNGxKe1tdETYmIX3FcPxVTlxwTE86vGOkLd8ZQIHlTmXlqf
9c+WovhvWaCR6j/JObw8DttLfXx+KCre1zPYgcDZg+GhuaHnhV4QfpHN+6WphRlA
kXEttllClKJOrDrImX1GpQoK/JQ5tiqTaf+mIOCFEl00cGzGEVtmcYsjR2eIzyiN
LC3S67DgbufNkLsz0goO4im0wa4cX1rVTxwQRgCEzNhTeAGSUXhjDfnrTeyQGe0z
n59uvnnpaJ0riiS+N5lIxzdOchRDVsE31nCoxEzjCAwFvLy+VgJww18Lt3Zf0zot
jehDpYlRL2xAVbuQhIqiAbA836lL1yafMm47T1B5ZMMOEv9VwS3nr81HZiZjh0JW
osF+2VoZPktXI/zb0r68c3tJCuYNiys9EbqxwnLe3CIOMPaJPrkXohFG4MKDgq1r
HFBPUwPffN2YkIxdJpHYLw2ww/s1v+V4HQ7k9el0XAbH/IwPFmiCnmvt4pKb7jvz
tOUSXdbrD78xae0agFTmNlg9Mqw9pEl/6nHvj6DiAFOSFbyNwpAvX5byJQLYPEu1
H6JvQa+Jjibs9WwCIjCUTZE7BJ9QNHwOVGrnrabVf4kwGhajqMulA7Xe+5divKQ4
0huNzvn5p21UFRjf2aCMXV4k1Al1mK6ov4Ei9zdWRXyrwB8cDlZbjhJufg1QgrnD
KHvdU8Xc08xdqdepd/UvCjPSXCYALR0TFvzdIN6Sv+9LTqCIgs15qNKAz1ysJFk+
8/EPokkmA90H6WiYLnHG+9QSXS91TXDVFxZe39RqOT8MegoibtE5zfZTxxcyDEn4
NvSJLsmaEaUvkG8FoM5flk5i+PnYaQXvMT+PrDyBjaGnVsoa7610KDxkPXbWyMPP
8Kgr6RTnzuwK9xQqCvX26VDHsDcAAuUlqZzdm8I1f2HUpoaPu9RxL+KEDNZ5VaUA
/MVH2DM2UMNX5CoAvTVOcQYdICcv3p6yOQiJGfUwiRHsoI+Q79bPa23xzE2vTkLg
A56w9cfEFxYxRtPklPgvR5KPkYXM1kdcC+OVTePKF+4qQWhEM19Mtq4qRSrTf5Em
D95mcu1DjsMzW+DTb0dpUX8XpOG+q4xtH0fadH5TVdPJKzjlF/FjXk1VUFQYmTYX
fIks0Z399gMoumq4vgBbS4kBKSQf3A5j51HBBErRtyc4ezuOzbGnuFc7J4rXBz+F
4mr84MCSyXR+QVg/tlrZeh//npeXVjSd6woUSSOvuJpiUkN+LfsnZIVN9lfHTQpg
E6e9edaVJKL0SZvKlvdjEMeXegaBr8kO/h/V7CQ8IfuOlLTPmjRAkX2wPOGQELz0
HWFndMMTANaMEf5D1mVAUhGcITNghy8gXI5OBU9635civlWdeMPZqki+wy33yrN7
GoJ03ic2RV4WtkY/LDr15xJHuam3VSAntheL+67vNIRhgR47665erQe9zDHO0xPc
O+vRTaZpVww/8iseLiHKWNhpuA22NWz/hIljj93ha8hY9hru6cWpxl082a+XEt7B
7Z6E1TV6Dtkb0C23m1/9sOtN/vftCQTT4l1oyUmOGswmHkCddK1egySsNjAWiM7C
7soXof1aTA/iGkr04G1b0x7dcUpAoQEQJHVvFxyRg64/GTFRYnHKc8MXjZI3sEFr
ur5gPVcG3dvIrPhv1pYr3Z0BrR6t1cOxbmoEcVn8sONBy+PJ3JEXmIKqlw7+dFSO
wQwNGz1YjBIuyAR9gz3rAe8YJSi2N5Xaz8QK4kP/pZ8MLtv+0sj+UE36uk+1kc5+
MWoPJdEzqnFfE6XVhNlN0dZHj2trl8AfbXJ71xM7bRr7d4arQhZ44Si3PYIXColc
lG7DN9S9zbm4pI0o2/7C98PAlGgFz5WfBPR5HMCZIHWNoQmakhH8tknDyNF5wJFX
+j0MNZWle7N8OX7JcnPMGDGCmZsjQTnkxE9brDU4Qf8QtiRtt4jvKvRqHF1rWNbh
oAeQI4UWEQDz93IV9j/XNZpb3lBqnD3fl11L45Yof9rHnrzAt57Gfzju2YjWSs9E
E3qEC0N153/17ZdCdAhrFZ65JAy1JIKGj/K4dMEYKxfe/Tn6AYXA/VM4ED1MC7Ey
h1Idv/HwGap8wh3K+NYJNaqbbu8ha9KD0/OHUhTD9RsgoKamueoC1YYMxWuovbN6
Hk6/jI4or7URxDrKgClljG+RlMLm3vpXSz1yOSufkjk9eqFY9gIxdXXrx4t5kOax
z7EShzwzLvQaYL++Y6p07/6g+KTC+Schmj39lwlZtcvDVfOZQL7qFARpErZXNpsd
gJpECa9J4xIO0r5FXuZc5d3a3MsxyU93StnHeugfzXRt1vGnNWVJ5QcR+kWJdJeG
Fna/2ejr8fKHE+Oci4IjuIeszVWov8RB1zqrRBZtr855YZZlOCIST4yS76kXT6BY
IXGRhXlO/02zN+Ym2cduYZGH94Efe5A5fm+s/b5Lz0rJDqKMM5ST9IqbFZSRsXXW
gG35chjYdnEEkpxjg9NavXIPp76wdHm+byCQgpiC2e9lSte83incezkyw8qz8ZWL
n1D+UIZa+1L0/DpkV9vWMzLKVfoMGK89mIXzrEEugR0U4wjp3i7Eypfso+F/p0p2
kT/QVBpkW1WMeqwBeiFDqxJXLHSn4Cy+9WlpfFY1St35go98UYW0Yy0ol6bZItMN
fN3LUCXy3XBQHiEBpCCptgTtgsPCk+RZaTbKpToGr6UebHzPF2/aml70FKZWNB1C
aO51p99Y7ykRa8YuF1dpmH/IRMLHv/mV0lsUAbBovjWDKO2zhGSeYL7gSDj9MD9V
az9SOSl2LKQOHg53ArnvmBezZLmmtVhpaR0Zo7e5v4c4OapdlD8tlKsVY+Cw7dN3
t2f7jBiIdrAlX7fz8sIpRIZJKKR4yPoB7tXikjLx5/NVa4C7ZC9g7Awr0iEhwRII
/a4p0SckzgQejdUYn1bbb2vtCKcXKW7CNgROfJdj+HYHBBH72kf1Ru+P5j+SrYDn
d3Zn4c9/taXsZxG1cuRR2im5nunTp7AW73JRdKHfqaIfoiwyTvDew1DfTZOxw/V4
CPoLLs7ol+Poic8lDB99+PaclXQNU3gg9WQ1HXO05gLLPuX4OCGth58hukmxOr8c
NeaTVd+GHmc5WMYZ+Jt7O4Jqk+CuFIqpi/94GdsSEwZOjIrl1UWPi/zXaQfRDXYL
x/IZKxDu5k6ZBfQJKN+wj+M26GVoXpJiJtAWjcMNneCVYFA01zYotr0U+/0oOoLD
u9fexvNvZFiOHvBGmWHibSu0x8AM32djFqeo7g2AzjMvJncHJMyavLlJe5EGZ7ZD
0f22f1EpDgEKFxFDa0VxlJTzzvh55YnOiFUkMcIXTlPHFmsak15o8iqLTKOf+gpV
AfC5EbJyMpceDofLRch6oQ//c0cLhAGnwelmoiszbQwoWsISguW5TH5K/RBtJ2/h
CrzcIHcBm+o2a7XOmRe5WZs4Wk9JzW6hJeNhtHORDfe1llBcMA5gXdsZPLJpLJM8
4YM7wpkGISr2G66C5o06ZXNMDaSzZDqJwiiazxX0tWtKPZEWzB5eu2MtXhjS+F2s
Tf02HSmNyp1bTPSRodQIGhEqQ8+XxtqG3SF4d4wshXBr13370iuBrltFyHp9Cmd8
hL7UE+vVqLU6i//A5CKladD3ypjl2zcxYPXKhQZnlKcfy5i5AlC+vVkp1W1J9kX7
obrzbHex/VS/ERAVBjvES7Uv9orrXupMlc2KboSE5wiCi8KUUDCRMkA3GBOJqVm7
yOS1hBYkzfSqiUsjfRb/MVDm4wvleyZ5I9aNjLjgXZUy6s+U604Xh/PFshUugc2Z
glQCAIdG64EDW7IYW3vdNK6+tfA4FS03Xbg7LnQIwqQ0GUo9crpbYVu7EAJioI1o
lpurHEAW9imAPpAY/q9ENHBSH7/cIIVf22hQbE2wm8QUyqYe6vPl4aEVd5sjw3gg
H5I1p4XMIuXsLPyuxlOShCvhTNrf3NrOaYAMkV7LM1tLMz4C9raRKmhzjwnb9IfS
UJDtxcsX0+CTOwM32iqnbb0geRo3+2GMJ1A1L9ge8TA14gbxNwOs+n0FkUU8xnkQ
VWZtkJ9AXNmz6umGpUJe1e7Tzv5pFJyybNVHbgc+a+l3qE0hX55Ygm9RCqcTF2+t
SBZdyVlOOwnE0N+potJFYaoFHvD70/9onhmZsIv0IaagpHlHZZxB53Be6PwKmwBg
n1z5DH6WWJ095xAcA3RZ7nyvgeQmlh3IarTP6DxRicDg+bAo2uHyHx8SSgiFWinD
qBCPzk16afoaezqMqIPUCHGBh1sJJtPQCPF8i6bV2ECQgIH1An8VLGwb3acMTGrQ
EJVgYb7vc0ZaDIkn9Z3mGyl3LDH6doBquDTAQcir6ZMuZntVEXOmgHtx4/OMu07K
BCYjTxOt4+rCxC/Rmwp+iCNidEm9TAZE4cEjJASFf/DS8fQq9BjsXGJte2CtrVeX
qpC5KOKsADzcSkWawHAdTJwzkRggp4CO4X+GobuBorq2JLzvhb8EnFVD3eNv4BHk
/rAFQCITuJjdw5krrUT3+hMBiTryOKupyQ7WQrj/DJush3nlfV5CxhnYDOGhKBPS
DstnWq6DnpSk+UEl3jZFeGBGsVW4+738eKGMnUrU0deL29ggkvJeAG9Fni69QG7d
MBHStepkfwp+vZqqWU7HDbMMZrhAo66Je2GfpXCDOoWnkjHAUISFXWQ9FKA0yPER
l/xgN7VZh3W4b8rZehRbqG3mYPDpx/uTyhSInBDXERg04d8jJ40wqjITiKHFd4xt
gqjWzuEscQmveMJ/jQm2axTF/iKn5apr1w2yx+GrowFWnO8LAAaZhNvHFQg0MI9c
J7yj7KK5axaT3ijwlVDW4yS/pIlCg+y+2qeWtsUzOjUWxIuS8//Go6UXjidarYzM
pqZoi/NlRf75NoI9FxhGP8K5qGz2S5wJKKhAmlTdElFLthj5im+Bddr6ognG6/Uq
Ocd0PqMBcXBQRmqxi5H3zc1pFUCXoeqL/zBC4uIlCyZdYM0lNL4jM/Jf1t9BLDAU
eGXv8ITkAEuimJsYr5WxBTDxZTO1ppaNlBq1b4XdNd4tHwPLNCpPyq9rPDDmdxK1
RCWWZZsAzA3w7jq3iJnAZolllEKVvId4KEz3VIHULByvAwGbUPz182R8QMN9rNQS
YADrbFnxoe5BTtMe9CK/C9NpFYFT7IvrVif7VWMGusPubdclRmwcp4GAlW/+KC5b
RA7tS9kP9ljVJ9sfaOup2Oao9onb5SMinmjth+0OiBC6jvl+Y8qTPZowhfGnZJU/
HQP2JS+wpXjy8WYmaPjMxgsO3abKkfKHAQfvHRPdySUJutGt4eiY6wh8Df2fJwZu
nZf33d+1mxxi6JgJadXQ4scAyMVRO8mSLykNO8dYASP6mc9p9q1l4E4sTION+3NG
7rAIKjUXQmoUOYrDqHN4zbgkY4hnDN4YiNZer+HW6X6lck8nZq+M46/GmvKjEIFy
8q9MJT0EO5a4s7OISHltjX1RMsspZmBJ9gv36/ea6nhtlBaJC5nwDZTX+a0zGNqh
n783t2D7VmbfIkbt0S8yUizW2c8RAbhmy9LvTCisI79lgJ1E7zkTuBsPNAysAsSB
3uQ2mxuEses9cqG0VvG2i5RGH4YwllNZXfbUQWjVENwRe94yiHMrNRavegtNdgid
IoomPfJt/NvV9bp4yC/lVBMKr4t/HaZescyyy2cHwy/tsNh8GMFCAouvouJ7wdi9
nwjwNOEjF3+vQXuv3j6ns3tXFwlHxPIHHxU46OhKIuqbLQXp7Sou+6ia0gcgJWPx
hXwJA+YnN0TS7BTPaNY5hBIEhxvMzjWx1mEolXuu9D0B/NtKlJpehoTKly/yqa6+
bwBOYdlU7QL7H6weja94CC0o38EzcIHU6votkT/MmsJTltZWZeJ9zUZdOrAFuviC
39RxvxmqgItdHgICpmL+a8DW45zQhr0MmDWM2rUs0j31+r4MT9dbc71VwhmeN0QW
2N2/s68BxwlMwld9xBbtoSanRBcAIF4YZoj1HpIMQhN59Z0O/zeJ0VDJFbNK2qCt
+sO59a9Tn67ulV1l+NkPYyPrXaPTfmwGZ3CkJueXYhXdB2YkNQ9XgX+cCDtH1QFi
mMFA7f13zTYlLvtAKymOTfQSrEV5jCe/FD7syqiw0JC2jSDbeillP3U6dBC4Ck0g
MyT1WbbCRIYOmA9EsVI2ckdjdgTv9lt4XVeXlNpRzUrj6wbuBuwKY7Mf2jz6zGHp
DAkw/ByZWipar7CxeaYR0EuAA0/cSQm2zLq/YWf/wltSKRCc95LJy1whzPI03/D3
fTB0tci68Je2qos13Clr3odvMwYteTwKlgA7HQiboDB/ucpEsKVbnen24FPlliMz
eKbiT29JasozaSNXgtx9h5w0GwsDhSBwsojzRJRw37hTtEugi84C4zuKnkdoyt77
YBSLKypnPRNakgTHf+S1tCALFRuPlkyJerkc13DNCdUVHgzser81o2Li5bhUTV/i
4F32BYxNSqesshVMQPCIi6tg4Skpl3OAZI806/Qk9t/nihZqKsS5nLfqXH/cJU87
vqpc7UCoGGC2RRVPU8TNVJyy+AqIHMXIJUjA/mdelnOe+RswFFIurd1AKRe/71wO
TS0qBckpxqDuUkWFBxGvS6tTcgWuYFZRKRPsxoqNGNfInILwTHEHaSamXPFVkg1y
2eqryi6D1Nw08qAVya+h2wMptpIQ904M+UeQLZJxhLyOAC9shVSfoT42QFXCkKqX
mGoix5asUvzE7hVAK4pBD/W7ATi1Hfb7+/83Vc1rgtRzsg+Hp0c4jMyDKA2d6gTp
8eLF2achLEgcbSles2sY2yHJucfZ4zx8wzQjuVTUkXKfmY8S22sFiF9ZWoQ5J+FW
rS+EcnixiT6aKzpd89FqlPF5hkGEKlj2vlkL40SiD2GUggj1QonMfGaNXQMwVAyG
JezLTt17O8TPjVd/W1/g0w1hae7R6xFQW4Oa3RV8iTjOPcGI18/ZKtFQ9zRjn1Su
wlG7KbI19xOZ2IFDogfaCNbwi6rNLPWdBpDOeU8UkDaN4tb9+cQLz5glHmgfgJZr
8MA6jkJk4Uocpus+red5rmp82lb95rxZ2q4GWBoVimejvkQ3VqhqUeluiztgbMug
Hy8dbrhLS8x6xU7yp5WwLwkPYEzDxf7DI2g+NaMsvGP5+rjf0qUvVcf1KwpXQGuw
hQgfL/MGIvKWvm6jAQxQEjy7CJ8A2OpeGnaicRkIcNQJOxzRwSDLmS5Kf9Nii8Im
nM411cdnMNip7xa0scrS86CXh1aYsBrmSRvcDA56YjiPxiSCpefFyhqL1LI0F8ny
h9r7edYnjjynFtTCvt3YdntGoSetm404JXPFbOPiPpytckSzZx92Vmv85+vn54uQ
cb5cjDnMfBngwoXjkGRUkMUC/Iy2thAk4ZqSRy39T2KvgnG5kQFiVwR/xRp7XdFS
x708+tCTpYrOM/7ew0GOBFKE6aF2L05JQeB95tDz+E8BhrwiWVfh/rSGcr0j08p7
hiD84iyntKM5hwO3za9i5LA0eFyDuGMtkJOEVZUJ8UvEmbnJ9FA0Jd8BkSQzSNXO
cLBpsJWd5firyGKH8dsukKR0O5K+ODaUc7L/SLuP6gwdXkO6n7LeBfODMxMdh9b/
H7YOK0jcBiNDZHNNLZHvi/KLr/mb11yDEfJ3V1N3Eqpj4eLYNPl/uf/XM1Zr9hcD
NXhni0QJ0wx2LLpL57ih6DtbMWhlBJFijGgOmkU0o2t2LNeVQOG+ryzpXJYbuFoK
X6vBlxve9SSEGEiN2h4OxmtkH5qmw6YMB3ITxgyb6bxzMK3LpBZldHS5WP1oagpc
q5iDwNTQW8oDVe6moSvjYqZRtwqeTwdn1eWXJwpyga3Ya/ISF7wBpPUeGZvz31lt
W/K/8XL+z0Afg6yVeCZAP1iH1P0oBG/P9ITcTLjXymdbSzd8TjEKc2u6aV15pamR
y+u/Pv7ouz3HMvSAcD1zyoPD85a9Q7qLLbwlbs/7zGkbMy+IJ/AoGB1DKqwAtnxe
q7VxN60dCoIpVBngcGFCq51h0yJ096JdYvNXCo/Vb9nf82jQplby2FBgagwRe73M
J/vGeSd1cBthtHU2mV5QI8f1wbJfdwnlPeCNcH9IP5ba3t+k0+tATjYqd10XDar1
mS3RedhLuaBQN/jexqLmvuAtz0U83bB7+lQRyc+dGUKapwoyZrsYWI5w/twQps+g
SzbxI/KtOUG3G41Nzu1i/tHmLRAECmDYhlReCzsnAXP+IJlmgYSZHGGHWnVO5ceH
p5XxKnrLxLigr3+nXPavXxJxt5Zl1Poqka6ygoTiTG3je1UTiMtTClunTJJNwAQz
iJ5Jfa9ef2KJWm+R5DOBUoSviCxAYaU/gG0kaM6FLQOELG6KxwizlOshFdVDVyUQ
1ggaZtIQOuSDJD/657tq4mAYRMmKWIsss29tqS1vWT/43ccx1BRw2ut3z4/s6PQg
IoexCa8HMyBVbMBYAEAFZ2/9ZpA/61bQ4KzoN8KbafXByL5liuN4NuPA24/R/se1
s2/ORj5sy6KiVqI6jgW8+wpwEYlHvzsMZAzR5Hnuhe7l9MKre3EVQL2PSUtaJBZD
ADfbmDvIZjxoU6arwvwYW53uNONC+krPUinQY2pjGkxD1rjCUvflMRcntBNpgM0O
3D1QOUoC4jzIZYR60lGbpY0nQeeCyBuHpVD2jotyxuGwY7hZiztij2od8207ixIW
7GYW/xc4xZMBy7r1X7by+Z4VKl3Yz00FRAS402iELBtlTVVFKeBHNdRoiMhNpan0
BxwSvs4q6Na/nRb5jHnDqwAkIXHkG2eCUbIvUIVT+k7OQX4IpSW2n5IJuufWLA3p
COBTsBgkirK1yQlY68Z+bcjet5Z/5yF1PTHVh1M6pxeGxr1fImKGNnjtiJWvr7H8
ASC6H0hBkPCxZzcU/DsLVbN+QExukOPExl0AyHpBRzcyahJbUlwRW641zFe1oX+g
0u3fUiLi0YJ0kpQKx6ypySvgzr9e5sNpNy/VLJF0D4gXw6zYuAZGI16ghMaBrhp8
NQCPeaIaf5IUGzdMMvWGNfNLjGIr8hSP49QfvswSyol3cg4J17C+3NXKZEAhICWy
in+78zOxJ3xMPm88WbZB3ErXlmjDEBDsECCka/8eESbVmUjUqnhrA1VUAgalGaX1
nlNZioqpoDU7+kZbyQzU563DwZgX8UrrcaISZ/kv99ik/NWcXOKk+CsR0Jpqow2n
6/4+pF+6W9ucXaDMzB6qhgPEXWpxsbOsIUOzN49zXkMaMvHzNFvMlv1Yn/VbCSoV
b9kkT/TGco8tdqgfC6iqRX9mDmIjL3vbG8Mr3n6L0yUipA7RsmRkVgKOxOJSdWYh
SaKrzYqtK3eXVAXJgyH2kiOgahdGlVvJSzWVdYA0kzMuSrRp91CVNLSI/OLu4zjA
5HmiyUhlZrTly5cauBYwWIUfCm0LDXEi5v2Ur55TFDjv6JWxMf+iUTDVZQvPYUDy
QeWIhebfO+305eBxOV/U9ejGenMu1VJBTxchQBRDBZVbkCjPi0U8gqyCp7gM00YF
mEvVqqCbjgbqcZoCM4zEMjSLHEmDNnsXflS/MybFNMUdLV5pfFJkaCpmC+/uT7r9
g0lHDvTPkdhpKY+4vjYEE8/A7DO5KDiZv/HiU6HydZv20s6z1RuZEmw3Wlr1+TcU
B3FeBZO4ZEQ9HcNjrGqLKVlLAeXtHWGrHCfyK7UQEjFAyd2Oei6lDVxBQbvDRV0g
TwVfKZiNCFo7R4rQAV5XQs+LM/hefc9SLmneacGEn9/MCWMHBU8fdSzOkdNLMXui
xThJsV0h91a528rt/Nswj7JgjBQHVDrRW6lvHEg08ADVIae9v5Z20+TXq00+mj6D
Nd6D6550nXZ1xNcUoRl8ZH1oCOqtFxRRlTjsr6I3Nrm4kWyILxKmSUZBUOSQgKs2
Pa9ilyZzTqvTG4BkESvZJDAlbc6F2K+YDjnUxrDYmUSU6uUspTgvPEP6H9kt9mVz
N509P69wlERni0beuwuQp3TGbFpfDy5CFNJvimhAaFXkqjW/K2b4Slnoo1HBQwgJ
7BjeQfYjeYvRbpgVf17/FS503PF441WgyLM3US0EFfvNRr/zDKM/bW+ern6ckFd3
jPZ090/23azhbup+mHJElXIjiTMlUCtP/vzgzQtghg47YueEyIRXAZYN/LKYsEUC
uCnGyVI5hKvReCdb0JdAdRPXI5Wn/H7B8k+MO1WEjOW9yqmeBtcpNsLy9q4Ft35g
5dV0evTbl5nRX8aHiiLe5Isjan3WAgPaQ8jc+8X//30Gb3wfroQlEfF18qp+dat6
mQuZAaiRHgNA2KnwgN4VAKbUxFfEb9WuJMSkH2KExQqux7SliKq0o94lv/R8ftlp
2njTR7seKFsC98RQL2BdgXWqFPkxEYmFlWaMwOLmZJmhEJ2qh6fDR91JB8Eh8ifd
gQ6hTtetMg1I1F3JmQjzr3JTpg2upAELU59w2RRfOhIg3r2x5keVbVZgRwfIHLDy
k1FA1LQ/G4avXoLDJ8lbfxBuFksAoSOj70Kf0Ck5EZ8SHOxFRMQKyOrB5oOet9VA
JFu+Oq/4bjoWkRNAP4tfOobqytp2GJMQ+DJs7DXz9wwwwhiirBgLyiJ0RIrXKYWk
r4jRnT6So9kreyXZsvLmL+FuaxqptQgZ0S1A/n1BVzLPU25LG5r2kRpo3G6CjURi
x3gYbKPgX6YgnBg1DYjF13IrwDduH4n6kF6mu1zlp//Rj9kThj5+3YpRXbDuPh5F
xNeqzA92ep3xegJsizCMr4kbga4nAXp4yXtnyKxgDoX6UsfzHdYy4rCdhpzJKihX
fLYSbyE10hl2G1Iz9/+g7zWuoG638L2v4dQZfOH6XVrTNdIOYjDeZYhPJX3Wph2W
1gKQN3L6I1+24/LX7SvrjlhGuPYnA38EzbYYVSV/84Sc7uzx+AHEcfddahuKzVbr
nb1byY2cd7E2HoAmar1wapeW0gEJ7Ln+m5+byJ4voFQTT2sUgmTxoQctpT3FMx0l
GrEJGAiEOo28WllLWkGoeGHCKkM5l+qAZXwYuInkB7P3lvBVYsvqBd5n241gi+uG
ikACUfHJA2B5FypJDCCBUnoCbtVZRriMexqDUy3Cf9KGV7p06n1K7pCr6rY01QXX
WcnDF4rthAa+bPJvn0uw276Y/LzeqSJn7NfK40RjxW/lKoZJb5j+MBEyPtlavYBy
p68PBga6cOafHk+kOyenwOq5qR0jQv4ZF914AUCra4xlyrOOLzVjqo6rK9nfqyZE
wahPn5bxl5qKgp8tjVmu+1yKRjtMxIDXqR8NtudPVkPyZFC+gWS+lHNaOcknfJBu
FeJC3tIByHu8B1N+Nw2OW5/d1koZVE7D4xO+pMC98RsSlpCmuMj7NRZnAVtwGRSI
FRRR8UrmEqSWrMrEznGhQP3kZDsODVOQX11li7Jjy8DUQXm+CFO1u2xagZKVNK4Q
WPo7Xczq0HNzPYL3Zprop+4AQp0cqRQRK69qesjMW9Z9SPk4vjdTvBmz7jvFVhlo
GPK3ozjtf2BjkJnqUSIxcdoXTzwhrWuBdw1g6qs789Pp9PMy80kiWc0S53sc1Txx
ij2+BlCXqMAr5jWmIpqTGNjgjjoVQfuOZnPaaYY4E6w/BfekMMLT+iZXzEU8XOku
jTG5+wpb/AOfDk+JZDpARxdgMfqfxRZrht+kASMQndkjWDxYHKlm1udyjhUTIccY
PmigM0iO7qXGOP9Iw2VTle2X6t+boNkZ5KZRwrR/7h3FNk5i86hohhrm5xo4Mks3
XjkBnMmrEtxOMSiDvKyLeWBBJF9u+GxWVXB+zc4r2uRUwQv8whYPp31Z8Q/keZC+
yJvH+PWWYwGj4LEQtIkA5qhY46CjCjN4/sp4hjqWoASchaNjbSkkZfiBmI5atBDA
4kXzFwYnffDTEJX+Q65RskCnJ3jI54vOUpG97WjQDxnDfUXsmoPy9UsSzziZboFR
8o+3J4yYdDHozNLbdGTBpuqZAeHaXSrbMa4wuF7mfQG2VE2UQ6i1i0u1YibhP719
fYuRx+LiYFx5adC3T5z1zIIV/okJB6DhUn7zgAR6UtfKosl63h5G2wckpRtEUI6T
lzw5ZIgr/9QN136CW61Tr9WISexRXJB4hN1Dgn+AAKQTIxqeUc25TfWMlBnGOfkZ
6XSV95SwCY3FnnGgptdkf75zeomLJTO6GTbkKf554rwbyXt1Tf9pmno+AUpjSg4t
rP1C6mb5JuLwzZuvvwlws7HbNll61ZON0HWmAch2dtfjNRnj2UCnHgL9mNpGw9/B
D1cl5wUfozOhTMoeWzTCT+iXgWz0e5ER+uF1eiGOk9TZdHnB48rxqskcTvwrVbJE
DQaKicyktEmlJVdBHL6WvqG5tvdK15VrwCtc1oCmF2bVbY9E7rZCkBLxuQ2NXlYi
EDkwOlmx0tGVEhArvabjHphN88QBhgvoRiFIzrs832mhlFssctN8pYGMSSuOFa3y
uYmDtiaqHcWLnvFfU/hkyGfo7BNZQdZ7HyibsMtMjAhJktvmr5thVH/b0ZBpqcTs
xC4hJ+zz/kwtGbGbLpq1yP603BQ8Vj38HWKYKi+1mhtSCEzI82T4CKDgyGO1Z2JG
b7Kn0DgOpwwQitaxPHZl/OddWbtSvZX2BGtSTLgKSIfv4mxxra1U+pxmuKzP24dz
wS9z/gOvUzcr46N831DBPyJl24ChWQqrHYQPIGfd8fVr4pPljBwfN+B2JcY+eYoH
wL+mMtPq6yOVngDhVPRzy6HDgXt0nuuP0+Svb7/AqeCwI2NvA6Ritj+/z5GZ/IlC
Hr4qfXQu63AoVQtJD62rQhlDxIS0nCc5rFU6vLdLc8namADGpn+pQYusJPJumDTc
t8Vsa4qUFX8zAKfEDO/of08B8n1zVk8aQCUVgDCmwVHfmwcmVDOb/6piPGn8BPrF
ZCLKMFilnmm0pS38AiCEfmLzh6ACUhG5X1OQ9U6Fhms8Ucwco8tRcxgZBx1X0ixi
FlNs2pkP/AkY5tO2xrHpr/yAV+MaWESRHWwtMmh3PPK3pVTdCmSv9JUWJ4fXVOFB
pYF7e82dXgET6E0sA0TcOJJ0L3v7ztJ6uFI5wgSt723dpNE+wIE+JfYRI6vgV8vj
px2xHWcszSyRlF9ueJIRchw82CAzK9iVuVuNqo+1b0Bb+1n51IbwMUgHdiXDbbti
PBpitLLTWlWUW/mdozivneoXzruvXDkHP5kLYuHDd2mXnJJnxBj7Rz38Xylk3JsF
ICFVJUDQhvF8lgey5XoxRHPOvTHYa2Pwv3tjScXxnR8jTp2eaGETaG1QDoV2YIdF
Urv03+toZhgKGBZcmGa0WieM/j222kenMy+mFDmg8Vew8rxIuCgSTKiWUOzEEn1f
DxVkhGCGwa5UwVEUG0Z4G74YeMFk+AAiF7GAOLL9gU1XeueBUH+QbZcAGZZB2H6F
AjSf5P8QqxwDwfX7wbYaDR1edl22OKLIF4Sh+Y7xvDDN1xOELX9hatUmuIylCvqR
x6YEITEnRUPog/jmsaSQcEJ/csU2eaNYe1smUlnukr7v3a7Go+uGur45FYVNs4yV
Gp+g3sZfW66BtPYYDxcqVIDjxGrguQx4caA7N1VqeGfWaFscofUm3c+R/IkI28KU
KwyQm5umAMGpiPEDnNC9wY+tP5kYxjxThHeHfLJtPu8NHZFmYzUdrRHLB6E9vwPi
sEHhUnd8Pz/YSkAbGtkx11L7ClYmtbb2p9wd72QTq+ZeT1KCXCTEAfc6bsOQtEze
QsoR/Eo6u0L7v/kQJCKRw7BHkEoa6RMsradqpqQsdoBIfMdN9xCN+8yRXowueUJC
ouibGGYKr0TahRa9/hNwpfWdH4YE+4SNguMJHKV5Yfm1meriJtcDVT5I91n5LplC
Z2N6/o8rvHvf5BMFL9d5nBRel1Cqif91eNyrd+5+mPG7hatfNc2b9iNge9PuRkXk
yoZAmGsqEkhzo4t+qZ+QZJRp8j9uhw98zZYW3CIONocf57Fuxcz7ksCpbNEQAtNG
pO6D9hqEKieasokAtd762zYslI7h2eiWRMkK09PE/sBRZwUQ0oOTTYfIuhfNFgGf
NBkvUThrrR1ZKVvLyTdVq60QMKyz7BlTRDqaqWoANDiw/AmiKUQp6uIFfP35Wj1/
n2+BdM4g+W4xKvK0WWeUoDTtoCCuGSP2YTMHFkD5+MqqM959cLod4KwFfdNWX37e
HC9wxyyDG1kKrNu85o96u33VleCjPE0K1H6Kj8Jt/kSd3u3GOej3lFIA2g280b6x
+7q6TivV8A6blOR5RZBgCl3mQIxfRB6Mka9xPLjaLYIRS3POuLi4U54NYoMPYlSB
KAq+6kfvZqEic5Tr43+QNCWuFDS3wPkif7eHuxmfw9T1NADfBrNdTvBC88a+nD6r
IiL6wgUrKWc61ERmLR7t+878KDHkGnpJD3gnUBqVBhVEFGuibMg4aU/tKy4H6kqx
S8+30wwB1+iRlbKKmuyaD7diuPgSo3O7sVDvTJVl5xf7DeMyuNaq953GQ9wiQg11
fWnNNyUy/TFx6XTKTdgOlqv5A1l0WS+9qCbtBMr9J9AzNCrQPkJTfyZAtjRWFSwN
bhyZ5GJ/Olfa7t+YO0GcDls+ayMGiDBPk7B1IMsrFeHrSahn3L2zzyAuqgEuJCQC
kHAkGyrl7P99gSiDmUocPKwvmHy2J3c9CwABmZC8DWpYeb/EeuCVgI8Vb4uCEfPK
F+hdRgQGQDHkbd0EoY5dYFA4S1QUfDrKjfO2Bp++7s05UxReKOxGcG1MZBmsYMbv
dDldgy3pnOjVEbtAE7nhmPnQ1zfuvMMMJdQQ6unnuHJ+RTQUOfih6+ylhPAuxNc8
OkzqjTKvP1czsGrXnZ72cKoNHfHrg9KYlcXlOXOsYEKkRK5jl9DypUho46EmzrC7
Qy4lzyr74Vya5wxCAt7NpBHxlaMH0EoW6b0vez+EiSZDe2wIKdAzWptofg+aXLpn
vYZnWWFoGUUovQeVk5nnj432LpDw+Qb8uKf3qqs6rOmMUgnhjmmWmqCiptDCHQ6N
+Jv6ZP/SEuP60LPXl6bkGLk5JlOnx5wX6PuD4qxQ+2F5lX05o1dAa8gLqpV9sf6g
uvWwWCV2STokqsd6BoB83m/+VIkM5wFbs7fGISNqC9bfoAkpJcqeapUaUxo3ctO7
63lo3hJe546DxUEWPZgsojVc6BT77nr8PILVrYT670nKwWLBEQuXRxqiBRTMB+A8
3cloidJ9k91DNLRKeoI3SghHTjBk4vOlEswuNFnwb/LSqCY7nqotF7uFvGGRJv7P
FnvUoVTPDL4klC/nRX9dzI5e21RLNiFXMqiNKKzT8rsTPSgrMH0hQ7tIml7DgFRd
8rTUTNk1Fok1YLWvgoUES5I0LDSIEYV/UFrSDE1sX0PdWtUVFtnyp9TGGJN0ac4S
dAY5IZPQNpVL60lCay2Ih6cNLDQs9+evvjUdDJTCzgba0sAyEeUwHN/Oyf+QcVXv
Gd2wScIVLpn+X/ntq3xbcI401VBNLvSfnkE5jmP+lfNZTxoPxZU78Ui19jUHCcwu
Xxes1FS83qtbYsdOZTlDIvb89W5I1XPlgjZOfUmAWW+TqssldP5XRzFzoDBk5Opl
NU9QzkILZ3Rn/uZ3qcaPmqJi+UVTeVbepYVComYQCNPrf/H9qvGt4Tmc2vUvxEq7
VQXhsDE5MexFM4Bw9H4CqUfu8TXEdmpHqMSO+b10kBEh9fCZvpP+aySYB2RwthHX
HGWZ7C7vmv7pxqtdfLqud3meKjSPwhQ41ZLvmpM0savZVOFz3J/42YwIXzDZyB05
8tqO9fr5kq62Q2bh6/9gwSnUx+UfT2xOeQeLAqq+DVSXfyIwownJv9tm8ygZaD6l
DDXc0ugBLgtDjuCVwZMpP93hhZEN5nW6I+N62SAMIR+YzaP6pPAx0xjGNH+L+F/m
71JpjaTRi/vwNT6X/cF19La8sp6ubz8qfSWeqi5rAfasSAMU2evvDnYYvywBmZ3m
M07ehWsVMa1JwGmk8CYqODXe64y8ZqYPxiWkGZKQz0Mvo9zpTSNKhfqVqIkmcBOE
VzDn5GhqyeOtGmQH162p2klIyXjmxwdIDvdqkDOLmWD3eRZbgIJeEKuXt31yz2jL
oTxzl3ZrNJlIMLVt5lM1vJbatNbLmQxPRhVX/X/ESbcGMtGSxmiddhc6B24X/zck
DR9Ttr0/jPRDzyac4Ra2WjRW8yXqkVKkt0K6C9ynNJWe3Pwq4yEX9AqKJFPMWd+j
ey/3A1y7X9wKT867Gpygc8GYYJmm7Ku4PFfQxrV0X7u+XRSKPg/nwZSwEuFr2vyX
H+mUlP+KXCVccdtyFpoFUTYOhR7fRBSRA6W3qjkdTI89n9zMCSsAsMnFvQzi1Cd9
XDKILPUur/5C5mm+sF7Q6iMNQ8j0GZ+djJeJ0WQRg5DHiMmqCTE9TVYoHmrvdXF6
7qbIUaQUOhI1nlhtLiuAA41IAgHjMYGwtomUTZqf4ZCWQowmfgIj9Op4DWZebuQx
z2NmpjjOvQXRfdj7JMf3r8+y0XNICW09mX4TTdHcm7k3VnjT19hwGlMrjhN9R6QU
3p9X8VomAxd50ownuLqH9unRytujZPTZi0I2rssCVnUUX6Fv/I/BXWAPHtxQQx0Q
omWQKaz1sjfOxIfxuEEpZ/ulWjc5RgifwP2Rp9huhFglMRGZrQWux+cu6pmdielI
SzJokZq136vP3biUd6QyDTQBuNvjKqu/XDUPhOcS7jmh+egw71yJulNh0P1HOW6z
n7By3nLcJ3gkQ5xz4OjM9lvHqN9EoyyplQa6fopF1Lzs0rxIix6dU4YqhWJb9Mtr
bPZjs9844a2aUqK5f0FGSgA8+KoNXQpGxCLlWi2l+neOoxYdNHXjHPN7LbXVN/LQ
UJOCHY0RPjKCXQEva3f5s2gvg1Zgk6F2LQL6ijVWqeX18O3ysJcIuI2Exa1ztJMc
MXBYXS5sTMMc13tNEN20S+v13JhQDol4z5FG0S4reduCdyn/8IYOSyTfMm2Iwo37
4aFG7l4daFXV1OXQ9diX3EagIKnv2yT9ELW96HNjvtIDZBfwHXGmT+S21/+hkrvR
VqexgHNCwZdkkbTipeOo2fBV5fNF2/fMtFRmH7FVJKUemGNsKVjM0GZpPXEKxOLk
aJ4DJDfj/M8aELoS6xfyiwFpjoVvCnoO6bM2X+D+FF5ferO7dV7j78B+hekHkU8z
aDsP1jy2zU8lXLjG4UWFVOB8XVGPKkjOLPdCmIBn2qbyo5dMZMIqqFNAq2LiLJuo
Tr8QeellmZO0BRvpFkNTRRksgUw5zaarM4uG7Qdb+Bzox+zB4l72BCQm2cnqYY8v
Lw46b6muXR34TNOHNv9XIVTCO0PDAH6tRWoJ9mJ+j3qhIM6jJ2SKnyNwZex1vs8e
Tqv0d3KqBEHFZsvcAMN5fyCNIELjO2Fa/VClgwkd2tHbU4uSAqkUv/hUHqzj5dOo
HU6hYEQ/8l/y0rPptxuZfSm6GhAUEpxxexUP3qM9ymb74BBDcYxpNUzRyMAvSfef
ATcHz154djuKtn4hTzy4PV/nkZUKwePNdVY3ihlNugDkv4Qiidkc348ybHn124MC
QLZho4DEXk9zSbHdZVzW2sHJribD+yCrLTJi66bLUNCtB1ipQUgtpG6PqwI5mFy4
+ydZywOjz+i51U4mjx5eWFzmjcx4RYreeVOQsX84wYQFN4PwQKZbyhFznEHarZ26
OzO/JZEV4aYzvZm9jE+gJ0WC82SwX+ajQVX+s7KwPMQxsQJGtL+RT7WgD9bzQdiz
9zN90iGF7h4p1yV2RHX3CtaPQk2ZfTdTA6kiRJM/mOa2wAqIrDAH+N47p2akB7v3
mng6SGfe2CwnL1hw3tiYzjw1wldKIpJ+Pmy7SwiRXWM+1CCawIvUKPmHXoi95A+a
lOSvcvJSPYuj/oluguo9nTT/xBxGt+XkQD15C+oGAYfSfSyHULjISn6QsXquadPV
JfZEJSJ7UAdzDNIJl0RAP6c6pN9Ti9COyZR8rscGPNAqDOjZtBQAZDiBiI80XgQB
jgr4awASKLfyVXMIPM2HxlsqzF36cfz3BW4dYTYhAeHsYuAJZQftveUm4HOXoDWr
EMzPcraW3HWSSVXfY3T2Ym6vSwzQHz+3tx9A8wkJXjA4MU7U7ILJEtHiwVbO1vGy
CqW2gXXXKh2xFBhDkj4F7pIjf2QEWYbkHnmHHikwR+FYMKcpUQGeQ1RPUwByOseq
IiKnPgg4i3EOxp7cTi/wX4cH4y37zjW42GYP6mVBIJWcf/4FdAxzdhGqrRm2xmia
fWqqKXOXR5oLwU6LJ2XLTYbN5GPaaGFU4W57dp3JNUC04qVXRFVxwEEq2y5zrTXE
lB/erod3iQl5aEMeNNWHApqM+iwSHx8APwGgOWCG1DC3LL4cGyuXwa+lRtn2+hh2
gDqwTmaMc+uYo45EhqZltMSg11+HFpodi6zCc3BgN9a07vihWtFH9gdJRtE3mXTl
9NiJrlonZm0xccNaHv6od0CqmLQZ09Z5sBIIU2kuwG/p2sZoEEOX+c3dLpvp3k3E
Y5jN0d9rSVLfYnh03GKf9t92YNtL4xb+SzvqS1I5ISycYVtEzza1faQ2ITTq5/Dk
5UAEggwvD+d0phBiIEZs9Mop3Z0NV1WVaITTvu//JNL1x0rRSOc5ay5/HisTnwbj
CGcva0vkXz6XPVzGqhZZC+PK1yyUg7YEGxpXS1haXSPZ1HgUjZgJC0c46I4FmCgc
De8qsl47fBRmU6E0WGL3kguNwQ0u/FgRxqyTRqv8zj5gncUAc+DcfUIyWYvzMUIl
8hYCapdjeJVyAwkyEvAvhvdJbqKP4GC3G2Zj3XemP1Vl1BTQwsRmZc/ptbEKc+iU
fOZLCypTtzpRSy4PzKWcIHugQdkoF+Ojt2rSodpOYXuJ8OpU2d0ncwrNsWhIRxQq
25kNp/oM1iEBuTecjwZ06SLX3Nr+xDKdSUHlyPat3BQztPmOJBLR6e+mtNAob0Uw
SDgTo1h6x+ieY1iunZS+Pt06FTAlUuY4eN7rIcSuHEDSgNf2dQ2bXK9Uh7pjDF1M
pHtpHQEl5rCKX2w/8jrEJuBvyPE2mDbVupb4mERR02gJCYvVN/fp0s2I8AQmA4Rn
6eL8n3XHQ8DG8ChhrdSm/sJAMAMWewsrrzxSMlJvjXR7rgX9spj0dC/MEz8h91Gg
4vBUwe6NQCxSbXT5BWdKGOqkAEx8TXP3lHx1U7gVGNlsCxfubBdSfqKClrjSuA1S
hxm59TiE8N+NWSj1EyqoTibARkeUyBkal0n/NruIBsRpxYgpDaa1JcYprJ9p2AdK
JvHRoSVBOJ05IQ12blbe8+BPe3/msnx6+RLYUHEIjRjRD28+fRsaoO4YsF4WIeU5
0DZIgT5/Y3xLbNqG2qFKEryxYvdXe+zNIvcQi/3csNCSkS1TN2njqxYmh6OpBx9t
0s+H8cPx6Y/8CJVRr6i9lZpJ5QTS6zPgcvBNo/iW1U8owSxS4+JLi5McV22E22WF
8EWuPzNFDJHSlTfLy4NRJzkF50Z7TQ3Ivs0H4OuFJc4Q7SKypxO8aEZs2QvdtqK9
g9C0DgPig1E1Yxc0Y9yzvsI4TrOCWNmz31zUUV1jIrig/MVzwkkUjVHcjbQ4f0I1
UuL3i0S0cYvXxL4aYVv5lcKrqYIKeAW7hNZtpJOuR+B8z+tvax3xjr7VbTk3J8Nr
WvE+fzvpCHGciJVW+yhLTVlUD8ujeJyMz5ixvMOJ3cyepXyS6s8XFcGGlkWRnmMi
V72irVclXFdAMcxbKesW4jI8ZGyi0+AzONLnO/SHOqBGZDOtAEgNQMFqE0LJa4Zd
LwCfyo5PfJ31IsTaFDiJDjW6Tq7L1S/9GDio03C6PuNAetXrqgbYhS8l8ZNwDN8u
4VOH4x+S74E0OlLmnTdiGWodzDAin9ziByBEL5ke/f3u0exGidMqPkcHB2Po4vO7
KNMglfzP9qnIiwNPbefgO9NtEpR4eFVN/JCqct25AdK80AxxHD1UbWV6132lklUx
BFufGM9NCVAnwjLGEtjvKUqczWJbxI0YGw+R0HdQpgpiNaotLVIheuTMiW/GOvcM
PB1Y3vsm8VJWbXMk4lXLdJZ2j7v9e5rW4z1GgLbkEOJbUyysdGxN36E/1pNGOWv1
hnKNJjRoVEpACR86E39imsXlwMgkLBzRfhpKuhOJ77BzsjTEU5xddrdgBetwrdVa
7aPWKRfoeIMEtvC/mf123DsYYXIYDb4KEnPPHEMqt866ZHaosyonKlYraAdRHCQ2
Grwz5f78BOnLRflGE69vD37czxu1p9HN8dsLnoQZEfBvjJTGwzIuX9UyO5S7o0SG
EjnevihE2OcLkEYrdxx+eSCHjT+/NE7oAvKCD+wkTBTrCKSKxy8MHDGr7fGwiaCt
ehmRIAQoZTMdehZzpbyxE/rhPhkUIyjzEdnkwM9xkw08JAncboA8TsZO++Lya4J5
ljAK1OpIX+VOoSPAb3V+riH+jP2n5EUL1K4nq3zWPaM/dXpurgP3ePGKJMvO7bLP
wtvGlx1yRgV53nBGpE0ikaeUcl8GaUXrUWLERIEw3DUwkzjjUkUgPAqGMC/oWcPQ
fr/LQh6CtW0mnnOFkSE7dg4iV3QZzttmfZDlTdFPXXJ47U1pyhWxSgmDb0euSKXz
/5V/uVn0azDxtkh8W4vQyjiuTkdYhf6rY44jiT/UQFs3UG2lVK0lndN3D2iXhbg4
3MyawhmwC0smakan1ejCsv6NEH6nEaE4zPIqzfBcHsIjBxaXC4ATBMc1PNep0OU6
sOvqAKOuO4V7VzRR9Zj390vg5ntXZWXHmpA6dyarsaY5COt0Dn/Tk9TXua41N3OP
bJUfLVjqv+9J4VcRFnL8rrbYspVUj2qEFIC+Rq2oiiegACRpKVNPzj0Ci4PC0w9U
K6w8uhlaC3CUFaAnYCcrSv1xQcaVH3jfL6Nyw0MbTP/iYzeT9uNcklwrLzuGz/Yp
LumTWexryUEAHIE0DnRHzsd51uoepWLc+CM+6CBqaVcKnsRvGW4VajsjX9v1hoT4
VjiQn+lTAWqakYMqSk6kjEmH8t5MQ6bfg+cSH4XvVtP5P+uLEJe+98UHBf9m6n3e
hGC6iQPQAZmt0gB6oFpjMQhQLVSF4cY8oyxvHxayAa9oW62CnnGQjHnvF6MobZLx
9nT1aoosbf/b+AH86EZjRIRCdD1n1HKLlBWjXP4FJE5/VM01NXSV43kPIFbbq3TJ
olV7AXVwsZkS5Aj/cdUgafIgYvys8EQeCXmvfxzRRnQzBlo70XOYH5OWOMt2Hgvd
qHZtpOQhBBzRXSXhoLPsYV/snnkq3V7AHjSH9UAKW2n5qJaX0WFdf4OsZvV5SRfH
iMNvRJPP3EfUm1gvtEOQDMdciKKz9HozW1q6ujdOeeo21aFC09qyH1fW6LXlGkW/
7ggytKShZyFpDpQkVmz4FcYlznSO9duDddDEXVR9sI3DQOZDIq8INdRLAJtOCChB
MMo04Arh5MppR+XOVZ7xjUnSTw6u9n1KZKNoG/JUbG7a0E+F5Zwm9qtf7PYBnoI1
rc+4qQ44fUCyJ3oT6jt6hF8DBHyynsMxiq3jQ5o2ntg97SlU1HTHoNj5NowkGG+m
yMZu1EEbe8KFRpzr7DmwNiqFEZlwLjP3AOuKMvgvTgKzdxhuvlLRMy/wQC5HRdXc
tHJjTcehDYbGB78NgirRkCQOYs6S875sTRHc32zJcmqyTFPz4Qqg6Dao+Zs2K5+e
8GBg2sXCO5hPAicKvwEU64zE00of6OXhr8+igBg7TPAIMJFn5QJHarRRLlLtB/Wc
Mc4X6yi0nkDiBQEhxjwgilW3UAsQvrhwPJ02ap8cu946QgaOn527QED01RVIrQuy
Pf4n6l9uRa5qBRCD6Ftgs4fnrDMVFaS1zKztxoGc2tPlCeNQEkK6cHXxJqV/URSU
G0WZrvoGz3FET1J15lZ6l+3kgC+xqcnVES8Aje0kV5bnjfiAZzHgUEdUjMWmVb62
Kp5RBlTYsirAH8Fp1ACDRFcFD/yE761td92VqhmwUC+nDsgZqKhbKvJD4iUqDKeY
3O76+g/0ZHZPttMS1T6kaRaBnYjyrQE4TtvsSeRIUhH57ozrHilO0Qyg1nIRMmQz
55XBf4oCRSMAzxgoeKoK4hc8p/Fngb3LzvCn0bTQTacrvHLribBfs1tkZ1BapXub
zD+4DTKk89/nFAtH7v56oVWnWUafndDIoJBeX2YC0CjO5Pn8waKV7thzLMZRxbjF
6OHPorl/h2YwAhW8B0wkcSVaSxzpHGXRKYt/t+rw1cqVOOUCcq7PUFYSbMl+v1iD
mRzMKxto7DyfqVm0noJgjnnYDCD8sc7fo2dInCsw26xJPxazwoaAGmwjcegxce6s
+3rEXCFeoo2bA76u7FcDf9f4Bu8duDdpTBZD8Mk23mhflXmY0vYG7IjVM6DhlGY9
5NkbHaa+/q65eV0SdN+VOotYEbgC2Di6rsF+6gaietftKRzn3Pe9KZytZeRQrIMt
cjaCWV1w5G5QPFit7+fRL50QrDtIh6qo39xGadR5Xg8n9vnFxnBoIPD68sXUV0Di
6Ux/zL2xi3NkD/jaUDx0SZcJibM9n+Wlrfks6DCT4lsyK+Sprsty+lB0FLTa8D3A
gly557N7s24BIsBYoRhiAEeVU6w5zTSzXLDoFszYz1qACMMk2sj1Jn5cbyFt3g2f
rfbzOujsv+8IkGH8OmfoQhe8y4txa7jkjlEpyZ1WzfxNrmpfmKVN7e78l1rRzA84
e1WMfmevAIJdJWSmtLtSrQ6axu3MgQBNdcHAeZ2/M+B6iTEdVpj7u367uPLHTaPf
k6lXKGMdGcL1Qf84F9F/Vojysu55JBbRqlkwO5LRUS98zDyaZ//r40/C6Mg0N1VJ
ZtioMwcxdNkftOXagi9zjNLUfQh6s9qfnXZsw0E7QsE1dZlL+u0Jqi7dNRisPVF2
fvEXRSTLHJWG374Gdt8TEC1LD1LKpRIxIhtJ3TOF8kmywvX8T+zZgjrF37Tb7EbK
1mTFS91DynXLVOL1oi1Pq4yImf9k6ShpcGlfhAhNmov8L725zAPIfzP1iAI1iFW1
vrQyJcw90OZeL9kaiSslZbVk6yAqx0qFcIvMDCtnjaJ0ndPSgq1G3hUIeU7Mpzim
n+n3m9ZtA3cv3YYWiODgdIVC7mbqWzRAqzlCwUVnea//cg7mYCVbweNpvxTYUFnn
CQuxAj6ZZF1hElen8LjUNPG4MR+tX3U7LHMF9sdAwY/pNtvZaAA4XvYqARdB9ulY
U4diKxRxqXB/vRVk6fV4oB9RLm63957YUO3GTMFEL8kf0aTAIPipO1E16XSFO/VM
AEPKvQxyRKs6CLftLB81t6ltTzY6JYLLQugASjGKgaI6bNyBh4aYDR4bb1D01snV
VIMgzQOM6Lp4u/9X1J5doBQhsTou1y0TIdKfRhkfzKiKTgbyeDbkdP14CDM4roAG
pbLxJMZS6bpuBinDdepj9KlxerwwiKKfMAPmkNs9kqqb7Mk4MJj9qOu6gWv02HE0
YKoA5aRpvxHhPXsdCDAP+odR2R59YB6osbYMw8yFY9vfj8Ux6ppn9egFNocb/mzz
eV8KFUxhD4EU5JbthkOiV7SdqWcneOFDSgvj4RDf+iiaViP0hDyL7qx9pbBnVfjI
YE4xc+u03s14CfZisz0Cv4ISTs/XSN/EK7I6494WpChkSf3jVvK2DEHm89T5E+L1
3nrXYp7xyNMoPkoUvwB42o6bnvQcmj16jUTLVz5CiSFNKg8vTdORtcWdngcyfneN
LzkCG4vsK+3vThJ0VRz21Y4VyDpavFksKwhgy46UpCPaA237awgP1P6PCIMIBQ5U
upNzg6eJf2skB0NCihPBvcAD2hdo7ib07xXdaE2SR4Xx3qnJi20Y2pQzGNiMsaT6
od4xZLdXO98nYwCyceFXWsYS+cffq3MW6pTOgqyTPOIMJdKWTnSOowR/FmCxL/+x
FB5r9jqJ6dWAaq2UZ+bcrlAjXpXDlW5yX0CfE8WeM7OkImbCJf43vtrkEqpot7cN
gQWywdTSf/pOQYPfXKoazN9JxEqtibmtjURO070ESOXHCkfI2q5CwoIOhdbAf6xr
QPltnhIM38z4E4dnRGtfbbvns1nqey2unThtnw3ZRZTY6VoBr7B/OFeCJd9kjWrv
i/ZUF0IkcH17NT/t3JajPI6EjzRgarrqauBc95QOGNP64rHrm7UcCJ/cly2gsxjQ
VSdPDon2u6NFuvNMnFWFLhY0ZddqNpxF+oCp5CxBw3RPzal2Y3TyR5jtkl7pTpzC
Pe3s6nwkCRJVE4+plTf1xn5HJ4E8BOY+508bi7iMb+AS6kJy+sGh5hn3in6Xxfpi
uTiI5fGGJ07DsgILQHbvdpQU4vvRrYfl8IbSrpodoY8DOM+yrMkg2D+rkOWpti1g
jHctdULt96Wo0IzFnPXbY8MzHZvbjoZoyKTx3JK9Qmn9ZbTzcoAiDy5sMnf76Erp
nGIMayYUTrHi/r7CyM23Rfqnbmuz2mN+7cvLsAOOmeLwVZqOll/ujhbu2V0F4O5b
D61Q3SXmEv9ST1NbbiY3LDaciGpPmRYuWVLcVr7iNjL33olxvJtaKmfNEXusJ+Oo
2lwk1P85xv08o/JhB1ddmomQYvT54o1AhGf+Gkm5LPVQD1HWJ8EAhySg2yE4fNmp
uswU2uUQ+wG6OJ+cHHM+POSK2H6AB7IkZOvySSO6ZXt8ziRcceC0nn3P4tnf16Gp
+ybOgY9LUK20W/YZtIZgqfpIPLvvb40rgIlC59Hj3k+PMRFmhSWb/3LTcMyRC0AB
ZwhYRvAELzNYHvVGIZB5QzTlWagWFPgaaDhkkI8yCHx39BQZK4gTTKSotrKoByxn
tDgGsuPruQDmcRQWyPBKEFwKJwCMQtXe3XP/F60XO/5mq2L/cEbIKH3ekbJFmPTN
2weL3sQZ3OCVyfpHOtXksCu59U9rEmY0atdAklASI5ySXWsxRDrg3x4v/tUO/6A6
Z30e/MWg75jXdprj4NRXB9b3bPkxkbZYjG6C4OstF1ydE+vSEtZoweqlJgT5Gc+V
+L/oDzqAK/7Nyr3mnb2er5aLWIebD9XFZWrFgGftvAaCrSuTrlf/dLQeKDgjYDd+
NpmE74tYNRVVZLarAXbhxy/saL6xcpVmtHL8avPU4/AfoA97+/TiDcKXkwawdY+c
cZ+7ObzoVssKIz3+FyQ4r/RsqMtH3OuUkeCqDtiT3ZINMToZzowVgT0J+veNEkjJ
fjBTDpXnkiEPsTkN53nI1dFeJ35M3y5P484DBGuYVV0N9csluoGNWMmJ4fZleM0I
/L+8KsgNXCuU2MRbVlfuQcVayWqk6/ywDYCnoLXZvmHE4BMnczx/rUjcO5XWNw0i
h3a+4t3ztwbx12WQJqyGOD2ts1pbD1xqWKpfPVtl54ZJabtvaVXrzsN7rpkEQJCs
4Dn5OsqOhVg2BG1S0Qlde35EMdKKmiBblAncccx1zUi2nyKDW36j34ek/CWRM+jG
ekW4h6dG/1oWqxFF/+7VXuRRkVqeuhvRr2Od5yNV1VNDEJ2OgD6hVrL+rhZp+OPc
nkXIB3AjE9iexh6F64fqOu2tW13EaBBx9urKGkeRdAImw36oo0lF+bVcXwjXIK3e
L175oiTpvwTUZSLUbW3onREpqw6VgxyzYw7AdzAbsf+LriHaRC618Hqk3kUUeo7l
bLkyxV56FQ9PUCbtqcyXQr4PYUUQqva10bCswdWyvDXbdHZHLv7/W+Njo+cEgfLp
uCDWcPYX2++Xg6bG07XKWrM41RLbRLbFRRR7oFEURmkwDhB+ukVUoVKATIdceTrx
0I4R3uL+/OXOjeTBUhFVPlQHcszP5nqHsogUlyIuxjZWg54QljtYiaZKBPjezErA
mqvTlNlp5VId6NBFicy2o8tFJPkKeAWJ8jMXNnQoZTgEEd8YypAdF04WFAPUWAcK
0SLA7K4QrYsi/KbOT7VzN3GZMdda8PSo0JE6Nf6eVU7zcGPf3ZyBNasurq/hwZsT
7Tti649g5zNWzcOCCpZKr2PKM7BQSzne4gZzpslaVrRcFbmlClnprlmAxmUv+5il
k3233uTmc1f6gjT049MI4LRgfkINr7PjMZQVyywNO6U9XZs3lr5YZRk75FOV5Jgi
+fQZgvfaJ+Rs3diYYWCwh/WcSjmcj76pdL81w5RsUB0uQp4vAQr5K3+YEIVSJER5
i9PSQdyOw0vRF8jEXz9aJUB8DV/XH3SAPs3V2bvnI6kXCsWrAKDcCy9mBcRzMIhX
CT5jxHIFGB5yetL3GH6mE2tlZyGOzfTvGiMXLDEl3Fgl2Zzk4vO8ELcztfIH95Ky
NpYXVJSsbX55GJXO1QKZGdl6u4Tl8dOmWYi731/7EU2oQmVhzVDwyDqht8yNHkYz
YRhF7uhga23cQugdz0XqDreKeykv+3uDmMwKhNRBC9eF8RbQYSHKW87HDEDgbZW5
BjlR6gVYr/F9i7Q6QS1PSH2VPpq/eSjK6FIeCMfA292Y3m5C7YWh3+L/VBMPhrUf
SQ0/wLuS2MxUWTXoHc67vFZ7KqyYnmCalOsrieuGGLY+rRb6B8aDFEls58lDSriq
hcg6yUpSBTqSDkygjcFmUtQ36PPwAEHY05o5U/bMGzeCfz32dg/05P1ZDzOEkuk6
dvzatl37Uyww3aD6rO1NgQKzagEPrdAy3QBGyoE6c13Sp5Y0xa/tUr3ST4nMpkDA
xZ9Jzg9U/AhhUFzThIgOstPcDsAh4S72AJZzxdpaulVzn859/OeVqiWXC3wLUmnN
+E7HGVIDkgxo9pusyZ1WqZUJDVz09CQPpx9MtCbd29GgqGpNBYV3cDwUdhxQWJDE
tpiFvUXEfOQKE5BgEF21ZrJoZJZ9pBA5VOvLlU4OUYBrhP2v4H5TE4AxZQ8bYN+3
qIkJ/mmITiTWivgKN/OfOvHiWLDddY70Zsyst9hgWOtryM0AGSq4i6DkYxrGVYUC
VVz78elmk+EhngYs3BBm1lcuCLgrJN7mzTm5x9wpaQzPBotpjZbud9k9ff2wAHSs
5kpqzBxVxP2Yg7nyarB5n4r/2MCsfGFCFCdl+lZ72bA6at1OQMaSb8PG0p9jJ6bx
oYMHBPhvkXBbXfJJcFLxGF3ZOjzgznW/CwkfoSx6Mwxq4HI/YwwPW9ouAOD2Bvht
Xue6lhJTa9AXozrrb2sp73JpfvGKVF+Tnl9/SzzZoEJ6QZ+Y6f7iLVhEXWzuoB51
ZxNEaP0K1thgJdS3SLMI6aUsqsJzc78CuhP6jBhhjfzeJHzfe9KNw5Fq9GvB98FW
gAYm0kEZ7KnKXMa+ddijBiS9xaK/6+1MmaYaeQk+W37vvg9Kby8I4duUM99UHzuQ
I2z1whJc27Fd6sLIN03id8r8a4d9mgEjekIpZvAPTKBvRBMeqGw4bWw92alJL3+p
OF/6d1kq1MLy4ZGKs48b//klq1YWH/hMs99AQPQ41pnmpq4Np8rBbZ9O8hCfYWOB
ggvNQMOZw7LeiOfdiOgP5x7fygqTy9JWG5G5TnAtxSVVZTMPgJZJ06qWc2RBYm9m
UU8Pic/bqggOAzYnwTqhO4pzPziOOO5pgKwOIwPdwI4tgq81dYiwBZzjZuor9ALA
7QokMZGmUIg9zN6JJ9c0pZyEBjLSqQxZAo+o5enWBiwWeUDjEDIHQN/WohnX66ti
Y16jnf4nRa/iaUMNOeXi5Pl/x6KJC2msanlAp1mF/u8ME3jn/9Dsj7RqRQDe840Z
8iokcBz6DGX2cbJZxMDXk7fkPfKzteCxW2jvjdAXPK9CKEtSgSUx3LisypSYtIbA
z2F4tIHEBIImEX5pYi6X7NnwabKli4GlkYlrfTfFuL9wanf/9TyYOb70rtMs43EU
8DxourNqOoMYePxc5mLuHAGSTRdz565wMzRGql6nvbR9FDoY6hNHsultFRKMQlYg
m8u2O/VC0ufRPiUK3SKS7LLsb3GHrKoAvZPlmGTZWs0d084NsZ6aXn5xRIcDL7CC
hiMFX5OxbwU73rCIlBt9UGbghHBqkPAJcL1iOv4RczjpeeA364lzQ/YkXch7vcx3
yGWzmHbw57tjJMWjhP/nLOt3RHRolWxA9dUkj+yfg/gzl4Mim1+tv2WDcOb0M/0K
7x/WlOtYHALqyDEByU658Ht6I/ZGz2n/f6DNiAa/NtFQ46fiYGY+XDdcjJaTYZDm
gughuSgf8MOsRpbC8kVCtacFe7QEFBncjQZhcjABg/HGd7kpaq5/LO5+tMhPyjTl
EW0zcIBGFrvJw7YYDNVb35b6r8RMUMsZ7OzJJQRZVZWWym/7rivPoOFILfVjK2LW
yfzk+wTBBqlYhyFndiWUAeP8Cr8qIY0WmKsidYlSu7CEAqrntFwIJ6Vvi6fHlet4
QjuS1JNpBf8BHzATokzD/z9S83yQNQss511HT/f0ZcZf5DIWss7fIY2g+il9hBrt
ji+qlaWBc4omrZwaxHy7nElmHO8ze6arWOE4IMAxw2XBV9qz1IrgcdtCocUcnLG4
1trW33PP73Y8gifjgqCxlEH8tR16aSCmRzZjHDWWuMQoONgXkeZWMv4fAx8vMMcE
77t0KhRnSYSDTD8WyFfj8qeWi+O1X7N1Qpt7j4Q/M8pq/2glmO1aNEWqRvS5gD1S
sEypgE6L1nworf8jrm1wPjwP7HTBTJ2Eu23zB157L4T+5W5IWVk/XUQIO+zQj3hR
hfSHQcYcLvLmo4G8QxfTEaAmKSx/R0JyzsSPhcQ2CWwG6D9RQgB0ixkQsn29ontT
Is2OVltZBoVi0eBtHoPrqjJw+tpJeiVQawbG35X6Lb+uvsga3IVHoc84vxjHVuRm
HcWeT8GgF4NbIhB3SF7rZKtI347rHL/YEpmupMg6UP3anQPmA5xTKPkTDc7nYYRK
fd6QcgJs4ZrA4O2XaPPFTyWil6dSnVm0lDCORoN9O4BTkSQMSfmJEzpmg4cU8nc+
5lgttupB9Z9j9LtusTK46x1bxBk8gDbuhRxLER7hKdzQqg8uOBZVDxDzEoPGGT5x
m9AayI2TB+utLeHxoQE2dZhoBjr/CFf+D5uq0d2mJgmDiR5z/iGDxj23G779lqen
vxk9r3tggwNahmmmJoRdJEtlpUrsyYEAo50hf+rMWRvsW/ABRRZbxejklYN0YC9+
gN6muJD2tkLK3LQ57DZb0jTnCGEgbpxOr4zFWqwFzW/R1n2/FyOu4qL/uVOni4ig
KFh52QbFI0iH2nCat/fA6tzwASvrXgzrHXaq/nzcOGZhrakQZADOKj9+DeCy/c09
RGULvjw3/mrBQwSInMjiqFMxSV9KYTtyGePw75kbgA2nC+w/NfTiR1RtwyL2a4wv
BC1EVxBYmD1m5skoVdrrLosNCZ8KeOgtEDHKlXrJbXccfm0KBN4W2Ll07sFABeSk
SvFSMbFBU8/6op3qKqpBJxkDFF7eQKW5kKINMkjHU/ytGXeulQQvR1bOCzjDm4OV
ydbavUl0XOf9kzrVLSEqbNcECCUjZOJlnqjqALHvdnk8nP8XaOCZ3lxRd7XQqqBU
IarhEJMtRm25K81wJDJ8pw834lroHgAe9ZKPbpMeoSX5CNlImhEHFAn59vMjBOpq
RGJbfNYvCxrluAVc36w9J3WA3E2dirRFwqTUBBoJfBKvZvVLzxmAQfeHPly1GANG
B4f+FwUwys8ufR8arEsrw0mM6sUt7JFzi+eBCojwHF/AvWQyDMEofRE/C7ip0sfP
iBhmzHj4XnnvvOyrxoZbIrxT22AtGvGc4/nvUVd1ckDHIermaoSDBmsk5Vlrdz1q
irIvACbRcc8bjCohoyPms884pOBB4DVFMOmIUOtPrDc/8uju0cKCiDF3B9Wn8Okd
aH4w+7BouOwtAFx7GEavGMYl4PtM91JxAF8wKr78pTrKPDqPP4tE8gcvz/X8nxti
OiQCg6ja0j0FvWZCdZdpYM0P4URpu5QcUlsYbBR1pEVhGfJGf/uF1GiWuhwV9PE0
qqIkzMmm07qZwGOJUu8BGqA2l2lFN7OjAKfBv5u6XWEs4on1JmpQZqhB7bAB29YC
sCHRC0/PMLbnewqslk1Z5WcHRyVTA2fnimigpuamQeiNqO2arr2JhE0jBIl67Env
iJ2iy5jdrw4GQdDx98pXt8UqZXJjsq4icOngU1Xw/0t9uul+TJS/T69cztmI4EJX
d/zK+zL4etIpU3Nu9af1wK+BVJMXzmImRdTQF0TDpIwGpMf1/KRpY3jdBgmrtxex
Y+gM6yuPgJm/67HGcggICiFYONeg5ozimNSGR7T9wDxAVzauHt3lMdAYPaWx0Ao6
0qfaPW4KI2a6VU7+/+wQMcqnvWohhh3ffaHs0yDymkOOutRcEKvXtGQXrPKjd94x
rgDuM4S8LmTSl29klPyCzDwGUz5Gf0JngjSHJMMczyBJqZ5Rvk7/E+nXGV34BywT
yiZMAC9IY7z9OTSkVuEv1am5uoU18rlp1UdN+1k4idPgOBCToKLZ/9Vmk/CWiqHo
eQdaTppKZgEElrJrQZSGqCV0XFU7RzYNKNVChs2k1hAbZrxTXG29BJG6qe898QPC
+Cjr0z3rkvdlhcpXHArPOKK1zRLNsY7XIxzf5eYMBMd7DpKzsB3dDjg2R5t9UpTS
xbdGZFDA8LCdjiJhRESSSyIPzKnwmUCacNvRmYnTS23Xt5nkP0YmftY90MaIXWXW
3tEUnKNB3Fxm9yCl7J9lj4/ks760dTr+pB7vSwHyPcKWU/sbV9TX7Eg7JZIGppnj
WyHnDURFwfI+mOYZZtsCBPnBpMBVeEVimVI5TEeTUdT1L8DGhf8HUCJ2y8Zp6Zch
yd0oXFQTyVSAUv9szvIeUzaIjtm3CFE3rAkLnLvh4+Isebkv7tKTPCTqzbKkyHdW
BQ/6/eL91Tg9JbNY1jCxfq01/PlQ/y+T1x686AOBOrdy0z+qBXU0VMNClmXifvfa
AeYV4VOIf/LeP5Wo+/DQdwvpBzYpPgg95PZ2PYlWPstR+gaLMQT7kDMvbEvOqmBP
1NRFnJBb75JFWwdfv/E4dtODytdh5fFbcCr5yN6DVfNi1NlgAbMpT8w1mIZT6bKH
0zG32pq6crwjkioGenrthFb4Zkk3hfaBMqtzwE0RRFAVE9iWoE6sGdU1nzazqvgd
qdSoKrJKin6PEBdg04uj49beENGx7iSZVcve7+emlzH4BHbdLxg7+2rAzqDMqtD8
jT3isSh9zG+hEVrnhg1oq4g7b8mGt3RjcpxVsaDRMb2qMIQAm+S+EXdpB3IsMkw9
2hssMikD06wbaKKzdOLHHS/6g3Mf/RQEmyeIw0Fm/RxzYQD1EVoXIyeAoHOFTIlV
5xVmmRYgUxuDwamyYVgUVZxSi4/mz29ncK7W4uiG03lzF5vM6sz7p9qndviMqqm7
7fsmnqdFaWEPSMTsyHe8jOFi8zrzR6eAWK+UEMIcYzrJvELKNsCmRPIzNqRuDWIz
010VYKU29Dpam7HFEFTDbtB3Ws3sW/IYUj3L50Q43/QQgiffKrBwN7usFmp0ruQH
88mRnq2/o5tkw/CGpif/X2+O3HR/UTV9SymhpbrJzzUTrT8djSJC1nR7MCAHIgxk
hxmAiB45k9geno/3EnZ5tde3Gsdez8SxNyh4d/F22PLDQFnOxb7Mdq/5ZMDW3k8f
R3tqsPuXG1BJhBM53CurBGZ7qq3806/nBZWBxl1x9+qV6TOYMKEvqiCZcRSv9noD
fmta+wTMq3tnld5GC3ktLEDPpZnF3ivnsMByvY1xgjFiapTu7WnWrwiv2PEwYfBf
ejKsR8o1KE01j7WfPt7RydrdFPKkSCOqkDqXlBbMqiRVIIPehdyVbHdyZ/vtoS5N
ygS7qs2pS0P1T5YM4uQ8b+wyOE4kozBtkjsJrJYkdlJTZfU/0IY/hNBKFZpg5DIv
J2yEdZmuR/450Cb3opXKfwUjvC6ZyKWxc7C3W9mi+EKrYxE0tylOu4KnvU1M5MMG
g3zOd29cA3WYv/XXyNXKrUzQolp1yZMMEevEijIpDD/iWXtKCrzsnOWYrw0ziUQn
kmcYBbGrwJnLmOu1X2L2+21KicWRw4BGh0lckuZ7X1rNaMavWzQO1rid9f1v5igl
3e5aKFt+YihuFA2SSt56IBdeAXgtchgLpSMV+NS2aKbpQJMY+BlozMPSGi5MN4fB
Ezk1YPOC4jwSkA8i8GroRgtnN3IHXLmvKbX5WUpbzbokHgiRYfzOffI8zv2T/r+4
J+WynkAMszrWLNDqOOzpDGUcnvIuvx2dSXYXg88Z2/jtc9XQ84+zUqE7Kgb8RxRb
yVnn6JdUErDUFQ/YyvY0Y/MamwKqeE3na0HGZBrcMXNCn45gz9txwQ6wAhERMpMg
5awTP0u9tDHINu/GJqX4VCGyBVUfF39yXWCFeS/2HihKAtzm5xXtYaDTvaB559wf
zskQBALG+RGg5lM1w1okWva7w5WdDnlgjQQDN1YsxQmF3mJ2Lmw5Gt1wMfwXwn/P
ZskILvcMf4KmOwBjVzHaG5HcqfX5ciCft3XGEyVZaS7dG9aXTtoHJzg8fzLJosXc
iaKwJkgPe8PeLkfJFQArNt5ouZPGMygDN4BNg6SVaBFTlnJ1krREI5sGf2aLwA7V
lkXMK49wOin0I19H9tK17jWX3meEsIKFGnQvkfJ3nnJoirtvWh8dpgoJnTW0n9Xy
tZtWwM/3FUe08Wm8O15F9w4XHDpsXVohzHr83ETTw0/jpBb238lB7yDDi+62ofay
cEKT3GE09iiwzuMWMU2N+thCJezMYRndbo+Wp6WzKV317npsnm5g77GyxDhOkX3i
xSyjyXavlpqT+1mPofCaKTVWRGT5LBdKyyD0kLN8FetB5g9bbTOZC86cmcI1sajD
/BBpxOVAhijzbIDSniTcwPg5byRDPvioKM8J0n4W/UqRw+CXY1Cjrbr4JcGAFSiC
p4iZjbBCBGdNeFJclg4ZmkVHfDrzbdYmn1DlpvZaijOfVS+Flit0SlfoDkoFX0JD
KsyJMtKrkKmzD3y28lQSKIEKNE8lEPKk5SiwxM8cZg2HysUR6okxEbLy48bHMeuT
8v0k6/ijjwXBe1mHspA5MlvK88/uvjehjDKudkYMoTSfe/uoZ7HtPe07WCQNzp/Q
F1FOyIk2493bNJFxgGJRTraYsPmtsYjGijph9rNvJi5UGXFG9MB8EE+JjiK9dzbF
AigcoAXRFDMPgAE7syGcZ6J8Fq6svN7PsxaanGF5TdtY9PLf3tyxCqObrd66XlXf
NW0J6/C0PguHfmnPOUFQX/Avt/vN1Ds0nmMSOO0bhplfGKWNUpakrbZakZSi9thv
AyyC4iYUs3/5NmSKM/Eb/NMUh7Wh6VJeKxqJ97gm2VqPRCpN94HcS3jU4v61dlc+
3D68QPEAftbhHU5a9OACPHACeQAQg6H8tI/NSihab88GdqRMHT8ZyZI4Co5w4Diz
ruNtcf3auPT5r7nycjBKx51dkUJeaHWIu+WJSeQAo5btl9atz+l8ECRhV0qoemYc
9Fho/pNMvPCVcQkYJVca7G1o6Bfo3qcCJQjWzHqnlpvyo4UAnmc9oguVQx7YOB+S
KxsWhspTrWXuoF3udeIkI18fGmslp16I4OH169/AwGC/Ps1sVF9aXc2Ky2pkPdWE
f89Kn5HcJCzYnci2NsaduTz/ZoYL0TqrEGFesrtR+VnHpL6UDcJNqzVT9oiNtwTu
mET0XYRZVQhzh1RPD5nK/K9Gw52NK7ENVfbOWih5/PEeAcU8vaKkz2UuLu9XEe5D
J3tZ2roOe1BPw/O4O/nepWy14IlKggjs2lSvICBEyGjWwDJb2TO5CCEj+uJAu0Gc
8Sg4Fe69MnQjwsIfyHzujcv4LpSJhJMQ2d0rLsDtdE/N0YlwSoKTJ5P8z5JIV5h+
yGAP0PAW6lsVfbedXexI+SOjryCvfGS8L4rczV2uoyts+IWGjG92FCBRQ/JPm6IG
MsGWwpNJ5jhiWITxzOtbe7j2VaKiYOCjW2MMxSVqdyAhk+TsuRC/qL/r10Ix4tCe
ItFYIB2zymqwQPMlzulPrGuoC5Yc78B8q8PHsIJu+1qoUFJzWCYDNBb15JQBibKV
gO+KsLxV1u+7Zskx+sTLDPBOifeoN96iIXMZVLv8PTa0GfHGvUVQqrZF0n9gPUjb
XlSlkJMe1y/3oAZg8BCY0nz82tbyCVjZ6nTmQ2QF571/145szekg6VIpfIOqcEFC
scGJgcj0Gkrl+LRuKeYUDgn0GbcCb9ZXjGeMLNFGa+sbbnxWbCyiROlpv9KXb1xP
TSr4Eyb2uijK4zckYE9ZGDgmAYP2VMUKEUNgmd9OzRMitc0gQMGEnQ2WqJHZTUBo
HsKbK59j+doDv9NlBlD19XxGkuVfVwTcN4kTIKoU8CdBCMj0EkqinoWyJ/Pn88jP
FNnG772H6lZ1BLiQqluo6/iglcqgINYEbegVKfI/wPfETMbIGjTkCzj4ZqfRLf9V
2x0KY79nOPLMOSuCtddEUJJLNxWO7BAIdJ6rxFUe9cazTfoScvMnvdi645xvUb8z
hQaiVaFz6tVt+Ss0AAEOUF3PliB6trvPeuGchz/dabFfg4oS6ujgdA8chZNL+yJr
igX7ep2sWPLbIT7v72ldOQuHKfwxeet2maslzY8LGPiS4Ex8mwvFz4/e56UPtnnT
aPa/LhN1OYofesG9iUkCHRyfzG5PUUqF+zyuWM+CpdpUMNK13W9kVPFSBg1MLFOM
Ir9kLE7lJC0ZIX8/CiXt0WcqrGyuRANyu9Luu0Qzd8XPYSaUVHP3FbWnm8np7ZHP
UQvNwib3WaXrCIQEJs+27/zkM9BAXrgIzMHkGM238vUlpsOHGtAtXTdFEPgHGqhn
j0kawL9P9wEZI4lBCgqctcVk6o6laNaQw8WwlpFmujn4MHS4OPsL7Vl2gaw55UpQ
vawNslTvF6Et/kAttWoPAhK1zpC0Hr/VFmAIZz/lC4wGbFimoKLL52eVS2C7ImQ1
LgYM/TLpOdkNLDpvR0NjC797n7/YeUZIIXaQZhQvC++spp2kBaIIq20aP/XvBD57
TRvpzOvNolrQAJWkJyf8yQUWvgAkaW3UhLx7qBne/cxRTxj30hXUw3bY1LV5EsTH
rCnPAw5AH5gsoXY22tNVFR5xAd8S9YDjKfZw0CYH2vWgz+jrBJVcVEdSnVmU50MH
dwDVxKP3e+ijRqx2OBG1G6PL3UzZp5+wrViM5/+pHmc4E8Xmu6F0oJxWyYK8ETUV
q0i8K368GvUR79kpPNUQ8tyInw60B4iEhqteuYaHnt0Pi9vACcFS80Heqo8b8h45
6RjlAn+komlQvdiZq6Dna4FMHOIdMqbg6Wy5qcmy8/hJ6iHpfwSQ/LmlQqP9ORvS
MpkDtesGJBuE4UyT3ezZFblr/tFar4OCCJ+2O2fE7FF/oVlAVFosebF0qrcZk0Ri
Ou0SmJxDVDYrmOTiHtZciRlKG7TMkUelBj82JuaAw0lXGlZXkVskG45VjNCwb6QN
h2IooJ07uhDXfsG56J0YDQmRnoTQc9VArXB+37DVeLUTRAwAy2XvidvdbtBhvNuA
xh6IbcBItk+NHfmPyI67BFzL9nAPrvEPylx2P+pq1d3LnV61Mm6viCCVIQ3MXpFK
NBbaIu+Dio6imuY5YRqaWo5Wb5O6dCsOiByYsZVqIV5X64qYZPmqNDpQezjaucSz
RHPgOj6YSfq6dwgkqrEZkTJbCx10b88swWrUuXBEiAllpWBYE0VqkDINlqJNUC5b
QHQrhKGQwbPQI5cZvpvkVPBQ4/FSZyddLM6DWB9O2EdWnaO8rdyw2fO8azmf5ImS
e2N4KFTPJ/SUT0nfrvdCiYGKnvI2gYbffJ6OUKiPORNEf6EzWF96YLotf+tWWMq2
Sg1vSK4HR0Twxq4JaJ3Gkwqcq4eAAbXxFnPl6wc+w162t4Hs5QKvBbfExAJD7PAh
N0rq88rZaoCUK49F0ZB2XS27/C0lEF2eweZl8k7UarLVnAcoJLnaNtLmqWE2F2Ss
phXd/MNvcX/LoQdDev53LU38MH6P7UdroUPK4hN1pl/AlxH/HaZY27q3f+PuD2/K
AyKzSMWENzkGcCA1CXQakJhHNmXCrldOfPqyDKGuFGKJKnsvecYkzlUH9pFTJ00C
LUraIOPxtwH5c9IYE/fxV7XQ1hoJVMDkKlf3zsQFGx2GLkL1cm0/eDq3YIUp0Mb4
Xqymvdss97Q+Nq53G9VRTWzfc2E/0OTlOlBbXzqBPE/IqNeD+aQOx8H1MHNEMM9C
KWAtV8CQJB1ywOT0q+Nsa9pXSSy66/LxjosJgdbMXrFazcTBqrmSDt8/TSeFK1Zd
EV0lXahK7wEcYw5bg8KfXTUOtMRJDS/OiqrpSzCuX/aSmQxDl0YB4hqn6N7SXejM
1ZUvJLlnPVScwaQqnvl8Vx0dAYhsBoYpkUIEG8mPDyt8WImE65A4NGyp+VzwrxCg
Q4cB2JzSnpHSBvusNRqFuGkKDt9DbbNuyHtKjUueD9Ni6MdjPzX7CiQMMrvGOeYv
O2uyEjevYJlwLn8TVhpZ8r+8wB3WBx8/1onjpG6E24tbX+NLVwSsvULCfcNU5Asd
SmeTAuOIS/PZ3QzE5H4EUSl+cQ+tYc/tvFT3kY5fZFGpv7dZAPfLEiKisUjqApsZ
vX334H2tJXNBEF0oyi/hdJj86E1lxCe2rlaqj3Vp+We8pQYavsWVhACpe0o5fiqk
tE1oQ8wdfNdsPEakTQcxrYcK90yVyyewthWSLMo5JyNJNio3JwYge+DCfoceb0jR
4Yz3kunCqPGRK23+hhlx3IYIbK6YD8VD+gDMB29/QCTU0dxMWT7teYBnsxogzcdP
UjCkuchn0hs5X/sohY2XYjVoDVPfGbpXWp1pPK9NL38yJct6JoZdvc5z9qc5wItz
dmIUw7Z8WUw4v8eaN7BBv0vNqeQ3EUYO4CAwTz+g/NCKS41hULZ4usiLGjDtZvjw
Bpf3PJtpRklsbMfTxQIVimJsHjVbJC65Y1eRRU0F/1rIVWwvxCciM+1rvM0B15em
Xjc1ONj7BAHvBEt5IqkuiY5TE5lvSuAD6tQZfBvdFN/EJ+Y0sYStWJq/TqPvA5iP
YaOntTAM4+jkAYR7IhABwT7DbIl2rz2fI9sEVB9KRX6HWNxFJTn7LL+VrTSd+9hv
aimxnsDmL1YBeEQdKMNzt/HMz1hgS5/w586T55nD2Gx9s/BOk81+Hyf5PXzeqWJC
TWmJQ4UGgY6sqEsPEBOcjqbn+yPvxcCemQOSVvOI+0A4Foe2jTtSpLOvLh8fSxoJ
pNosJvNZLWyQkiiRpkAb4p4R59+TAfOPlKsSdveARhnFwXolO2kDlHEt6WAFPqRR
i8IDgIJPu3lnyaZ+MkUSbY7TuhzeHzUkrGYPH7asgDKuCwUYx1yWLpLOjIjHjQT0
/2tK2F8G3WdT2FQubD8SwdNo7KA809i85aVBOj3N7x9eW1yZcFFF8pVDFAOwCn1I
xdjnY1uVZq0/EHQ+Nr37WrRoGIifyOyNVJMIAAJJbfh7WJXLr+/QUEJrFLhQmTw8
JMpiO/sKwlLuiv/9PNPWZTlwh7ZX6W5saiFPgKJKgd7Yid7lwxweVgsB5KnHRNbi
QvRKPN5GyI1onWzLLQDqQHMxJv94/LhL302Q9FRg044WBpTnHJfwXCkMwqTKFtV/
hfpukvGbkLYiqChvj4wLxsgE4UHIqlc/3GmK+h6ZUWmsAJUO6sqi3ysCfdbdBaCS
Cy6IY2faH4A1Tf6XVbRpbv8AHX9Zyv4eZl/PutQv9jjzmGe5ZlplzJwQ5DnWexcA
8l/82BcTsayyftpLbKE17emc2WEkQX9K3SPyVhmQi+TzeMWQhEOxRZ6+i+2K9Ti2
6FV3bbJBdl9xlt4QFaLJf8wMlrka0BHTwUeb54Q07FV2QUkQD200DvwmiZXWxftd
gHyEYuhmzyZb7CkeodrZTkvKOZWEF/KRCIl3TY7FxY9AigTzuG+rTeeMWqHAvNzL
UfxcsWFEvHy/C8G5ZsQ433iQVwGDsYSMgVlkvxXC3/mDkjjO/fpZ1uJ5Ov074NJW
ooTCNdTWd/g0fLvH+sA/lBcoFj9/lL/EGO8iL/6DlWIhQPQrCNuNkvlFMOOZ/GL1
b7hlkAUwB38czm3LNTou828dNPEX8M79gm7Ati5Mq1xgH/E4yJ5j5Z7PEiywIgll
chdrdxV5JCL21SJ21SzoBaNcyiRFAxfnkeuHT+nfs/rGU6fum73R0waYeeClyoc1
koOz9Za1/PigiF5Ee3O+2npKaXGPztpDlC0pPzjXF7n28QkZ7cRjac8kSFZlkmYP
YwL5oT/4L7iR071//WQB/J+dZnO9m7SskezF9qssaMsm9A1biXtzYQoIg/KqBX2v
E3Lc7j4/PNIZX5T1et7JnPS2LX+uWYspfWKFcWqhKcu3uw2yUQrEMudO8zxTdSGX
n6JV91V9RJL22NbncwpcJQXyvGspcTMSVm27FHw21sDyg8lp5t+mTeaoGlcMXsA4
QaYmUauAwWPBCpHh7jNoJ4SU9uRB24/gw4yACyz7S3YSChX3qx7ekpAE0i43xR0q
J92fdi5MEa2KSYZNXdKwgmAJ+TuEalUnaejIJEIGTMWb0UbObXBkbgpc0YofWnVu
69gO2Xy7egtRyt2Rp8qKRyigNjkT1rICY5/+z0/c5o/yT1tA3xP0daESk2fwiNv7
rdmrJswRjoFHzqFJrJzkDuwzg3A328CVVXE4R/oW58Fr4xoFWdwV7XePxkwHkn/O
+TyLiWdFWWxg13aN31vhxJTgH09fE0vhXKzIb/nzjJg5riFhWTA4TXSyn3+m3n4T
GY8nJEChETnZ2w9mD2OqegLVO4TS9S/5rJabrK1GSWPkngvaE2fa1J8f//9vp1pm
gnFxxnZ9M5kICnQmN/hnP0tVpF9HhFAy7iEF60OZReKSGDsLMNL0wlNS35fdN2TO
8b/13oeyyw8Caun3ag9FyhmTdZjh+gMLZzVHhG4ApFQbUWeXxhBLmGOlNQlL/DjX
UqmbY3l1JyNxc0vSA9xveVLkKRiX5JCWMHJbvftaXG/aZ3XvHjmG7YPKtOJTO027
tId9tVF+B1m0loR7D7oaAy7ijpTnLUKMnqY1VFCKmSq4nGYwxMwRvurAjvt2Y9o2
uXRhjyr+NEu0GmQ5GThvNiF4c1P+4e6ikLcyMQaLegLVUfG+7NjTRv7cAA1usw2D
7O2koQ5zKhWA7dv+/aexjPldyAdC+Q30kvHtgj48hJfSt3vWudXWZLicQshc0Pm9
U+kLaD54kZKfE1OaU3Dv6EbPw0FLwUmXruUnNBQgoYFrb2Pzk+7WjV1tQb2MXJDP
XTiQVV0hzbhz8jMcMM8gtpb1uD5WzFUxLJ89sCtQdfG7UCuN78hMpg44L9MHJmsT
XWCyLdr7Img+Idn4eVIfr+2YrdOJ3qgGtd/IejA10faGO2yPMA64N/+y4bHc7qcU
4tO6B8AV/O0BbUjg93CQ3xJ7gmBtUR6tN/t9SbdQBVd2DiaqbV7uwrXfeoA+6VCM
Jv5Allklp3ZZA1PTDqQKwkxjh/eKqFBjihIVp7FerjWqaVE2tUumpjTg3McteyJ7
1Q/sjtRzbLLUnB7P6xyV6i04tATRwdXwXcocdOSfWxm8EuUzbQB0z1SfEIPz6uR3
yXrsWyjZXkSGqbdn0oLBkyOCNfYLY/bKBN7XVRrd4suev3m2mttHMEFiMLiJxBhC
tsXpCXD9qAzFL+MvMstu45drSV4/Lf9V14vTaAOi0+oMRLb10wtKc5f0W55v5VWY
w9YiGP9Xzkrr5l8NDXn4jhkzibLYURBSlo2DQfEEbl5rxIhYzOR8adX++ib4VSvp
9W0s7C+9mD5baz7+PDbmYDiF2SBK15GBEQ8818yeTeoFOoAUpyEOODaWEHG79YTA
LG5QnHtQtBpXUir0W6NnZYnMVPtvkcPm1naeuWtmxRLBAMB5lBFkd/tUKUkpOqWN
dcCqODOVEDURwZlUelO/sHeRxLC605JcIvpuQUEsKenQXdpcHwdCXwdZsJ6PYT+d
JsMql8Vk3dmhGsavOpkqhmgFpQFnKyg6lXdundewko9woMD1AsMxt9MoFimb2hsO
+9MQSKW4TOMc8r4bRf05SsfdX7AfoHTsv4/IdVW1uCextywG5k7BAgSDSfI81DeF
wJCh05KMyttsSmuh31D/dvExkvz6mvUw4BVaIgF9wOnMurzmXjNSeg0+XSlJLOxU
+HGs48pgdMRpSTUheh0lfwuIS8lCNbf/JlZma1+cig3rjDJTgNFBGY6X2S4Kg1is
F4umLHt1k3bWzolZt9HCFP4TlkH/zxpwI3nfib0efsWZQj9KQU6JFt0u0gV5UF0m
+Mx4qzgO8RLLjjnwsGDTlWqb/RIkJcHeQpUwMtxJZEO+HMoD1DMthrHLdk8YvKWD
C6jP0Y4mArDHP5qdzVM1AjQxEGQlmyfwKpREj5sTx0eSWiYJBBeI77czCAK3TaXq
0Duj0DibW75kLUOd+FrWAAn4zpCNN8RiC+HfbgeldtqSB7TAKHh+27mkE8/jP0Pr
N0tt+w0X77htAfAWAzg6h2zBvrxW0HgWQGzwImf5nGvWGQz36bhNrdGzh3sUg40g
QC9GHkmNRnIvTwPWGpvwjeTGXahlnigxbhE2vmskceC8mTUP+DDFqRexXLdsK75K
pQ7KOcgo4Xe+UgTWD8BA+Pe+zT0DULbTv+uZrOQXy5zpXizi1iycuZsZjq6unjfL
9mVT+NZZat06Ua0ZWf5Q3Oo9nGFi1AxmTvQGM2Xj1aRdc2mejhWhoh/hMe24OPKJ
yVUg4e8vQixEhKwHU5GkiGJy9Wi2sMSfxekKM6jQHRcb5QKPgqzTxLg2+mBRY0ui
IefonkS62kt2RadwwbQp21cwvHD1UuUKDN8XJtNvE2iPDaxQ9d8iPAL1DAzTO1os
SX0CYHgsDou+iVA85jsf8vopLRWdRY2pJNpd9QQHoUMufcK/1VdknW7wXDHV1Q4U
RstHLKWfThGfwrw3bw9QETfIIn5x2ylQR4NTEuPK5dMuvAxFGI8CrmC1YUMAfWHz
X5hgtxXilnYjXngAaixvpLhIYJtDcUNwX6LQZGZbe1DOaO51ffSmENUiMgQyg16u
+e66f/YjfT4dnxwrWrBJ52IfZrZarB6Ri4TKNPg4TjE4TGpIAes5fcMRLuX+CtzI
iN90fH4mSkObyPAMYVeQxBYjZG4y6mfh/+AIR0d7TTGrS79yicJnXSkXJ1m9cuJo
1W+UmoUOCdFLN8KmR2UDR+/j1IjTzv36Vw3pxdEQGxxWiBqn1DB4c/bLCkMcdYax
dVPOfiC4uu+nLvx/6AIV3Nz4lH3NcJVDBp2aBWtFp1b5WTqAaS61CV9OQC+XmYyY
0V61pAvexvaJkWyLgcdZchYftN4S7rkh8sshcwwSueaohjXjml8e7nfc3nEBowjh
bU5112ym8sJ2tKEWhnn3cU1l8PkavnNY95lZ7TEewaEr5VwEfYJbWB1bNciDq979
SAuRXoFPKdUHYaW4K3mtAwluT1/1xe0nqjYoXU9BzYgLS3fzU0DpGpez5X4QNPwu
jqoFxzlLyn29Q2qQWoz/qdp0sf9xo6f8u3kkuHuw8196kD5WXlbUkONmCuwMV1le
OZVHDoYevrI6awOg5sdRiYfMqpDl6kfUoYIv6+92NBxrnzjOxRcv1ZfkMujiTB0O
mFdQ70Qt/YWr6DEAEBDlKCmxRK0Aq+SDOspTIlQg3LmjqGeMudb5vXTHNP9hy0+R
auuXdRU7WspZUURWKGuhKkG4LOuvyvU/TweoHKyUpdkw5FpEXh230UmnsKpFq11w
g9j8IZgj1XNuHaaxII7kXBdwPR0qyKxvwOuomQAAlfA4JEF0xYfFSbFUlOFqjsZ9
/xODwyuQasHq6NAcUi4TNDYZj95TQpf0E0KaLXlQE0kzPcg190cqvq3TkyXNVyqV
7YCey5CK5rKdf+ByqtZLCjkdJT6CoyUGd7Bie8diJ5A/2P/hmRGzyUMI7ej8Vwow
TK6OOI8BW0i75TXDTJhDluj888AMGCd/lQaFNhpBb1EYFgbVzObLPcDTlGxJC8PW
0fcarL6MhFgwt2VJt8h68+cXFf96o0JQ1fN4MelPi5lJC0eQ3vwabNo4bYm4s4GF
DxDDJRa3Wo2VsLwfYBRJupiwC4PIBvOxpbgCiMNlx3KsanQ4KwV9/0FYJsFLl7J5
Et6YaFipGM41JzZi0As/3m1znqkLBgV1TQHWD5AGB5D/HQmuRPCCmRPtb9FVxeQF
D4FqoecvkD4K5dZ4Wok/mh5syRWZ2v8s9fU1Xyi8yf5TZSZmtAZGZKYVD3CAaIDy
DYqBi4/9J+gOxecuGoUJDuZGCkJ3DdeG98Pg57M0ZgR4eRnWHLWXEYnp1IiBml8n
ckmtUf9GWH/FUnp9DpI3tC9H/kqqE/dhOYZvHsxBhFQOXtNIzTPmvgid6VgsNafR
iIn+c2+G+7X+3mVBikVS6CX0G1KrJPSttWtUrBNzAGoe5iaGF6WdnxQCv7eFpHp0
3nUOc4lttxaoUZh0J08TWhxju+1LtVda9hDLcxWv5+f7Jao/Ewl/iWKmK0IJ2oqT
nyWRiYOyopKjiwwRTWRxs2943qcGWuBkV/67yWj9LbnZl/gk4mfUuOEC6NJf8aEW
BZHYwsOSZmgQH3PZotTvIBmahxTjwyZf45AXVPQF313WvFcnbQ1YemH5uAvp27wz
5YQYPLFPOuqJsGGKloMNzxmJmOvpR6zpYsUcTumISm3mFgP5PU87gEkgLdU43sCH
6nmfj91HsdubTyUcrTgIffYvNkgOYLcfcHfCkLc9dgwyjSolXq9EdFjE03EtmuUp
AqzBf5h2cYN27KPCbyAuR2ssdpj/Zhbi8DCPtvigrbvpgWbuBALrLZ581TZKAlLA
jYjxVlTPgiT5If9ym8xLG+hwSGyhGOIS3wEleKsyVx8suDvDz0EcrK02u2+WTDDB
eHZSCvCq74Zve06JrkIrKC3FHDEIJ70DLFjmG2L0iQhyT4kNzjnzJbg2WKA3eTUB
dOdeQN0ARJApbv0pnQnhTGdKmwzBNDfI8gGC95xBHmE+oGAzW5cspEovWI0r5ftq
aU5kkzsv8IpHgviJPbJaWenlS49peXGg/h0eqddywMU6n8Ukt7k8znoF7Ok8gudj
ZrglwH4YxYljun2UZIVXOJZNGdkRMSkMyIR1MBsyetCa5E5NDsFL9wj94iYv9dbK
iGKsntm0bzJ+xCVFrwkxiM5bSRpiFMXD9pmdC6HW2SKwfKh1ClcmCYB3U5MAMZOh
RSe/8UPyZu27bNEDttJiphKfINycTDKtnk9o12VHdpNrLKl3syo2EabhW9K3NgBe
lrSxIkO0Kaz4dAN5pXWTe74iQIB6OLuyHKBgqJIeArQzzJxwSc+bl4tMOpfgiMZu
5i1SP+7ly7eaYkjatPbSvheP812GaWE6+COL0eJ9E8Y6iqtQVL3lLwbqJHyO7XVw
ObwLyaoML8JyuN2cc2+pvivuXwZc6n1/nqDPnNDi/ra6TcPmHufy/W2mAqrE/8tI
FkGxOjMYZEL+rFhlkmLdOEv/p9rFErvYsJVcJfcKlbmecrWvrrwzNvfgQFSSZW/e
M7Wy/ebjbjvz8/PzNYVtmOY8d9k++D1b/O7b3zUYSgWnD/Hh/8ix5pnG3lkiSUZ9
BGwLDRaPCdIuwUn3vMQ0zUX/IE6lhU0C2+wK7BAsECaA+vYDHJDhuybFNrnfuBJJ
Y4SBJ7XrOrOcuPxC2in7S8+btZXoX/TWKqLaaRRTBHbc1IKjjgiDKf6NBhtRtpan
Xknr4tLzmh7qnV7ZA+T022b5NVoRZbyCt7w0JixyRx9CyzJs+yHP1QgQiQ+VN7pt
yis9JuRIm9VBsLGie8fXqSx4zdpBXFWOBvviMAgYONSGbbiAgl3D2LWARmOdBFKv
j50F8mbaHqGytN5TeDOLPa4n2YmwCERdwV+dYRB6If6FcSIEZKTwPmI8RMtC/R/6
waLN5BnbjAJLdGfgOT8O8bZdA7aob5RkwNN2I2qo4RKngDeX8wMBg9RPLryz0epd
orDdZQhx/NZJVQuF+VYH0/8Y92bLuxVkelM6SeZmbzlu/ySJ6sTJZEJ27paGGBFO
fH/96XD5ZYnRw9jN5Zh/VcgaYxY5M7f4Uw6ut3LEMGm0StCKYkAXgn9cuoxQQAu3
ZHRIsRRAqkBG0QJ8K1CPgqaBWS6YToq++wbjuOcy1WxdqUxeEuNMR8EByFIMS/G5
a1gNiKVMpLqSbtBD1Ukt+/d+r+NiX9deC90TQtopHOfnf9tf2ultiZASrXm1lbDy
VEAe663dD6FKDseZPLf/lu3MJTRcvDVvFYzO4II+rTex1vNNkTdbRuNbGZbnt5ax
quCe/pkeT4MflGMpe8SVWYoTs19xMuqpjJziNr78j/GNMzbeeyUgenfVRUYnXDAz
nujS7XsNeWD2QW06mAMHgNKODQO1ThaWHa4z5eqYUnYIlWSKXMEAZS9r9FN+VSPE
+/dVZ2Lk2t9pnXZMyxOe/SNE5KNowpcGmOp+PXCBz5RiN8M343K5uTf3N6+Fg6vc
mx0QwUdIUOJFk+/JVKsCsvPELu3p/766RoifsF9biQcm1mLc+F2O2H9jqSC0zdhp
q/P39OdYZZ/lZIMrFN1GUskUBsvx6akESQjHIAwYt2de7lci+APKeteA6tTTpzc5
ZOnkc0q9K103IlnsmEbVw7yMH5+RmPA1ihuu9KhNkWnWgnMA/8mKEp5rJcxXNaqW
ipb84y34u4yz/TOwUAEihIH9dgak70LmcSYvhq2w/A3oCUpJ2K1xij3Wlp9pfA1z
mJEKfSHpI+7Rd4xpVZMegUWDYrN9v06t25185S0hhaZ+9bV5AXCtDHSk9jv6baQB
O8Q4RGW048lmuGVE4fU5pyR/dnV6imw2a77fRbNyofDBIddpJ4CbR8uh6RjpTnxx
znQTCdx9idSp7s7cdrdj++nV5Y0Bzfqsifk6jIfwnxR/PozxcD08RVvnlGLIYMT4
GZdkryo6jHGljQ9IMXs8K2iHgKltudF4ffpKnmaptzy27fdqmurQm9qvNZ/JPQLx
8RwpE5o1kgJuqk273mFhhhn4vBG2kQLHycqGbDnaiAkO7UAp1EUzeTynTX4tDCDz
8L9wp8r2sqjThvscU9gvKIp8GG5YyTwloWgKB3/JgS3Z3rjbj/xcNKzKm2dFIB+L
NA0PEfgMvYCq+7W3lpOlZg9CVgUdr5ApjKpVesEyAp9GIAEtGd1X1DegVoETskrq
ql3F9K0rUoMxcvVeELanzcV/5bXB+z2V7F1el+fa+7vrslQY98YbTZdwyxTf1u3N
a05EuI7vWy2IYIJ923MsaYBBAjDlofw6srBBvQp9TIF+GM11o0kC5eLVvaMWZdeg
dYglU8cD5TDYvqkcFK3wOmlq/EVqqdVHQ33IHM8oCuPGOixy1BtCownZxc4i3Ljc
J5RW5Vd1FI4FWYDZPKyLHqlAvrFGVLAvQh7OaiKE0PcNJrFNuM1k0P/vXK+oAmcY
XYgwt/GENdU9C6Jq7WyNzCkZ0/GWuTz9bNNQ89b0YBCkB5Vq1ETQxaITGcIznZtS
8tRShDy6AHnmxcbf7eVecorVbOyR/s+s4lySBQuAp68IBAmY67MLm8Qim/z1GzVw
DfUWqeGgp7KLbPgSSyiwGkW4RyT740C242wn+iZ2mwJ724AslmOcLPd2Zr5rOGMA
MwzUrUalQrGRwdGjMSwABFL7oJTb6NQ+EitVSxDrD5GEp78YVAKwIvBlnTmB7t8N
8fYe3cfhQqnCLvVOyOrJLjbaIY00WX9s1HKWg1z9MNQTyONIby3x4f5tI8aDL4VJ
jtYf2wNTavhtJsUukTAFS9dXuaRG6BLwzHBYnk9Y5ON72+kZdoMIXNGjF2T+GnEq
9tm0EPkJIuzxwTv3uGlzK/7RyZyizI0vRhQxZxjMuNT6XQ6ZD2TtYjPT+DvXGJHb
yNQFXfDg+w/XTouvmoFnf3P0xyk9y87ov7Y1BAaeK+ZspjD4tupHcR61JJjfG8G+
4HM2B2pY6JmrkuUPqjZKBMd4gPuIHN3djdUyIMELEP++59/rHbncxGDP68iEIHof
IxHtTLP2c1sNr/Iu14x/8MIIEXnl16zqwB6RfnzWB5BVIznk9SnatBkIywgQG4Ez
6YUrw+DqdJqrCHQzCMFmy6XMD6paX/ywPTcLAMD+sa3Ez2HXBoHVCfBd9snGbPp9
QEh7g3ALul1fj61Xxdfh7uy6b9wPlIjOloRacwfbNNLLRGAzsmWcXwcZNp+ftlwj
o0xZ9D8dhwFDg/Xc5CsRtj43XKFJE5NeUOjc8faJzuS/Taf9QWbwT0uwtAHjnAY+
bz4elzAhlfAQ5j2pkGupQiikmB4r3eY9mAlzfFkOyr3EKqGgrh+DthWCvtd38KsJ
ARPzLwGJfbaCTfoejHErN3AWS08anMG63NfentOpp2R+opqvZxoTF0cVhxtQb3B2
5AMlyCQ6yWVQGB07Jt74Yofx1Wzk+0tF8VUoue47gfRsyHSb85BUbhTMKRcbB168
uULChXR3DpcJj8RK4HGnfEZ+o1DhEoRTh3b/shxSFfJldLo9lE76Ql06zIrqdt/4
tHkgiQ/u78PwjGZLN2v0IUscPNXK8wLsmsLHkgZ7l1gB/mFnp6pEXbSeKe5sctus
BcD1j6RpSiclQiMGXGju8V1fJH6yh2K42vOKGbfgTva4bqNb9QrkioE+iIjssG8w
r9oTINwAnlCzvUyq9FvjDMEia5mYr/X3dVZN6fA3ydOsBWZZl5XMceS55iyklPec
1/vJjEUG0dQg4HdYtxvRr5lveXY2mJwR5AcOdzATEumEQiouTEA3is9SY5L9GFuO
IoRjJhksb64rwnrKfM/OFKkVF7I6hp+MicAyqOJkcqZPr68B/QITL/jaCJzLdixb
fScZ1i3ovZhje3k7D7mAPWfA1AtYMLfwGUyRcDQcKcvQXhGb+tfTEfH/K7IWStME
L9VRlX6gFNigYZYgfGOfP42163JWvLgTPkolMBx5QcyFiMXSoMaa3LqKzRy8vjJ2
QymAcnke4x2saq0m7DhmiU80nvPaGG7oe6KW3W3rO4Hdj9dOK/JyzJiJcuWYLcep
S0OAiAI/cpN1QbCSfCOMsMd2+aNQ19raY8rxsnJy2e9BgBtLBuMxYOMAQ5bxi19K
jLFGI3BqEW2OJsZ+ueXZ21AujVSfDqeNEOVOG+wUGTt8ryCKX0cHfoyt80J7avoN
DYmvLDFofuvhU+Zq3uPVmvIO2tfnib8s3QrgANQdC4EeZqjU5nRy8ySZF8Hyao1W
mZIOM3HleBUZmwo44eQifwWwbBbzvSw1tomUOjyOPueXvqMyUyLs1wGBhA1yi35q
pbMxeWBwSzOkYe125Vi7DgTsYW7L4JKro5kqrrrOToAb8RFjjgS76XZxO8WzcpY5
QT01iFKo9s8v3yZTh1OYBE/qABgaEx//FFviaJ86vA6xKpYesqcwBued1R91UUpR
1FcR5DheQXpjiflqPuqHMESTbItS72hCsVk0B2uKgSVJ+VjgMidl1OsqisRg9al+
b1mxDWb2GA3ruIf/OFuiGIO65PMS+RKdatp0F3MD8xbiHpe7sHyfXZCan/3IoTDN
KIs4SfnmDNrd+UCC6FplvDRL9VJAsimBnrpPSCYqAAR940IZAAfG7on3EZ7Psjow
uR3/6xPf9VylqUwWO7r8LU8BikweqIsPtvWXgPjyH1WRlEcv7mDOO0LwidPuvQ6S
J5oGle0eLbI3GPPW6eSz2kFbktNXP95nEQ4Vbgsom4fBZxS4HZR5OzickD5Pbauj
fTeUYy2bOwRM91ho+eQM2fmrcTqeWr3AFD7NQUpF+LAjp6E0drTGGOSEaiCv1sR0
IgCK3qV2ImuVOba7rMBmv+VOV+yfObT34HU6idZcb0tGcaVRBbrkMoSRHE48jqWW
lCQQE0pWpQHkLduN7rUzUReF/nEqRd9rgelPqAvm7NDpSZ1oLLeYZ0ovs3GJrikb
VxEGXh9Zj+suu98eR4p8FvjbPAwU8k8/kJ0xUegaEq0KNpsR20V2VzKwqxg2IQod
eO8Ai+H1dweuo4lkUjAyC3npuz2uCVLtFazSGZOa/0XbiS81hWgsFwzczOQ+Y2Cn
0hLUQOd+eblHjn3BGI09PRJeLdWOJIZl/M1piFAXHjTMrTVkwelr+bd5n4Ix8YJF
xDK+rhohJMiWp4JxV2kZbBY9csePf87Buyx9mkppx8LvjqxcwxLLUcZbMRuO2woW
L/WIcGjDbGNyFqAQbbZPydOHzsCU3ep2vQT1gBWzFtCbUegIcH0xP4FRYMZXaZmK
eyG5WToHXWY0t1momMVTzUdBWzQnYUm+PK9svOE3F2C3DdAcwCc6J4sOlgQTe9Mj
rpManFCHNuXzcUB30QMiS/S4QhUcR59yqMq4JqGnQ/SzcPB4aO0meKbh3KZuPfWe
/oWfO1urQdIJuAlOv8oZUPfnwqyp+H0DYh//mS6GdGE93u/FSAxSJZJQ7MZ/POqR
w7R5BKfspPmn8OT0r/QD4cK17BKvza+32SI0OgHIfiAiqV6U/UDLc9wFTBSBmlxM
KT+zng/y/SDr4LgR4ntZ47KBQQCHrJg3jF42JkCE7U2hBEMr46f95yLhZ9hApkVL
j3KGBOnQCwbZ/j6KEM02zBwY84FhhgGV72uUt8PgTbgFRxhUAukzNxke1JPW+oSE
yZCY6HoTvtIGmE11vEye8hgUyX0dGeSbyE9yDYWwnIiJiC6RGZIiVTigPp8ZoT8J
d83UrkUcOrNoDMb+O1c6KnTXTelu6seVCPzQE7TbdrOwTxItXrZoht8/83hMoGRi
/OwccD6atW+9rgbZrjTwJQaCu1sm/9fOrtsy19iau4NkdPU10KWChWep2mqln7tI
wfdV1cxfONo0TQ3U6ZAjVEqlVdU0ZphpK9+McG91r9hl0CoCKBUhMWsju9MtxbNE
xFeNRCCQXfm7WVfE2pbptOaqqrz7o32CknxgZ/boUi+FbAb3eJ5KquW6Gscpk7tB
BES/njlXrVv/CQgbR5PhZ6fJnUfjTmizDXNdn5j0llxya0T8pIMa3eHu5v2vrxM5
JEosYRx72OuWYk+m5mNaR2ReS/KtnDHTtqD77aZwyzVZttyxwRZQUwCc8c9+g3P+
uBSrGXWGKUaLc/WvKtytvLyrAxPa17AQbwUwBIb7Cg0xa5cXFzJVqEL8xjtDpKmf
n/L0am+h+8Gfd+h1C+M7TOb7JLjWNy5BFgTv2ZZYBMVruIBp3b5pfvBbF4bN8qvF
5+7xrrvezp6u+WL2qqr5ID8SAcV3s/xPgPbXOQFTZjh/dTJJbk1WYmvReA0ew+/D
2LFNEaZmznkaC167MP9SdMyXZfm8zOVd8moj4386vdVOVKeVRA62mxzxWlLwFIRM
D18I50fI+7AcIItNpYS3b9TlLtdXERRebhUHxstT+dmGHGn1Gv7gQ4pqKh91SZPf
gcL4Bvr/RaNWhIvDLNrFuPRrmfVWGFAL534zhLUz5tpiHFDRUSwI8GgH7MDtiqvt
IbeClNKuKHeSdmVffuHMUVTeVWwgWMmxC2PtUXe4RaQSHOp41rqGl9j6655QqU8C
CIvQMlAx5M6E5PNJY4J6Wt7GtgLd0MuW1ehgbUBboHfCCKudXdKU06UcgYBz/8jN
hki5qB2LpdGz4MZJzMbJHwM3zj+6+QzmdWWc2UbDwYt/GIwjTofh7u56kUP1exMr
tf52Nx62gUyyZtTbdrju6RvNyd7aMlyJZf5JNXUFoZ5h/8eaCdpsKBPBwf6EQGuF
gJz0Z18EuKpMtamgUwBROO2fWLHV3aH4KBXCZ534kkrDOJpmaXJvtuLRiDzsLUSL
UYLQAtDy9xrr6Yl3glpsDvrK2kTR4txKQg42/YvLgW5FglZj60ui/pUG/2+TAhN/
pCi6k/mS65UOMq9jSG65fXqtq4xA4vO8bKYsZqbdflayNFVXx6H8Wyl9oy6tZq5d
Y4eK8UnMGmmYPOGwLNSEeQiKeDfJqqBLzeScUwBNrZ7y+19dhluUNg1eSxDQb/Wb
da0J7Rpm78pY7mJUR+pQUBEfAWkj9+I5Z9M0kvOujWTs4VHD2hxkpMkCM1DTStLE
ZDwUVkdRroib7+oPE3OFkpSLRN1xG3k710K1qd7OzidmQ/WTL7ie6SocaVRW06gE
FHGuEy942o5GuyPcBxOwJBYdiB+f3izAiPLBiCKRJMUTtDiz94+WVJNq80mrNpFv
vET1waSZEsy6uc34l6OIkoTbByjCfkw4LuaPz3I5DLdKPtHwyEzAvCjqY8e90Jen
BNG4eT5k+eeGRTXVJDwmWKZscbc2u+jjwtijfkS9tNyQMBbrMxnzyYRtKGYiy97w
uvywUu1sHP/PEx9oiqtzkBTbuxFuKJi/2nPnD2VWLuOsC089oGLPFZiHaO15Nzvf
KJ/VJJgBVc7+s9biG/tcfeASCCO5kbpIXs8qN1m7EN79R2F5XpWT03CnlK4plpgf
xWP7ntrs1IQ4wsvFq70tKe58oohIxzqUbmPveQpIkLJel0KdNn50CkG2Bh82q29q
HsXxI0ociTnLkVTdRz6QmHbgUao/SeJsVMz6fn+cTTNB/kRV/Z5Tr14qR3gDbjEV
nSCKsVZGUuJ5Jf9OtSsLGUrBfIBN6EGfENadelKnCz5B6Fa1w1cDDSfEa3ryLGaf
7PgpiLZA4R4h9BzqqiLDHfPkZz15Ddtnxg0C0w9cY5y4cTTo15rxGcdCAWs5oa6a
iJ+C2WEy4geRVeD8GejroCP1fAeVz8fPOmfqeWqr2VLIZENX35jOWa3K9TK7unYY
VWaLmChYcQZai8phUtTG+Hi5nypsITRVtfGSCMZHWWpo4ynyc2rL6yOQfWtKWsyR
Nay/CbCX9w0jqmufCdNJVoioDOUr0JGFIkfOvoxxvpUKx/weenYAurjWVnqCCEGL
Js/KtnpqKoPrOMiAhEAxTdu6nLp5C9NSBMkXv980ps7woeYJs4biUk1mBZ3zdkPo
aIgNHiT7+68oqge2IVPmCbzLCRcaSFXgNQ/3w/xQbnWpzeRazcsYRy59PNYlhk/Z
5jWxkzEG9mZeAWvhnDwjSvzn/axVyK9iMCwYuduumpY7f1pnc7d4u5JasF156Ih/
wmlrKh4entt3ecy0bApJvBcjjypIvuNXDR0Xnx1ws7jlH8k+PNOY7gXVDFFluWo2
D9pdAorWEL8dmHE7CvRvfzZVJIfot2Ae9BI+OC2hPIonbP0rYukDt8Gd6dtDlpQ/
3GWB7MfTE9bQPRBj8PXTE+Gf5VEVt3F1GTiSb4eruzw5knZkfzsqJRnLL3H3farB
qNrt6sSHcAFLFdNzQnSOzFP8A2qvBr8YunItcrA+vrlTyB2ZfUEArgwq5S8XK59p
Xu8B98sXZFLKPQyF5oSvJurlFN0ak1K+JBXr3eOk0Uu5mc9w12KzI5r4pKdNKNUL
pEYNNGM9D/sguj352agF2HHPHrvB0AvVf8lxxGAUbHL+uWbM0TewSo6V5R//MXXG
0/LMGAO6ehPS8YwDXtglJXENDYeLwFsQXY9+W8nTsz1Iwli14QbDfDlD3P5MCaWT
GVlsjE8cuegzmcivz9S0GieAWuF1WUr03hx8LD+qy30/wkmWSvaJLl0LY8Af4el+
I4lgSoTkUVH47tQoDFVeQTooQY/xuRDYWGDa5xX8ahXECJl5pSr2PjIdADNK/dUY
H9NS+3RzwjkrWXBd+CL6gBOOXQbqzLt0Bkuvw0atwyNCJW7EJXiyxrZdaAWZP/8U
ufcuD678EieSGBA6RjRYwQ5lTpy7Z9QBqCNjbZTFmYq2i9k9Q5GF4j7rm4Mj4/Sy
CkXJzszNk8Y0W6uKxbpTFabIZnPvR2npVOAN6an+UmWZ9rUK9TV/ezpzRD+Z9qwK
7cR4i0EvDyiSBkUVHiq/sc9mjZwOofwZoisnlna/tjNcYdafFduZtytawMTL6S+j
vvIABNGhfDjjN8wEyIwiwnzU2zq15izoComlxUGvBgYIT4E7C1KZPWAoLTAw9ZKH
ihg+LqH/LfMxOpffoI+lnSY/7Z+a+/ukqgUurwlsqcX8tzwX2VUXUaS87iR+nGsk
NWiQQnaLQcEBCIKsV2ggdcrAz3nWvL4/ajYpWFHsBl4jXxWjG7KDjsCtriA9SVP8
Ox/8AlEcOQjs+/SHFAfMmM4W7t5nFcNGOizxLmrnzH9jjuWOzKnx0U6aAale/Lr9
oweHWQBJ0evjgYzC6iovPhC0kT7SkA3mkgJ8G5ipdVbxf873/Z+c3DumNH/aw3cx
z5jcg36u2GUx1KjAzZacIVBVMVEKLKpCm8hUFMQZYNMyCQ11rFx1/4I1XjgYHfBt
uz6GD1pdJ0cBeV7qcEjy/7ctnkREH+D0a1cb92C7gMmyaDw4MFeUlqckboGMWQCX
IxN8kACe2b2R49t6v/ZPEZ57JGh+QY5cy3jxwplEKvZJqs8G2lBjxsy1jxmNOTBM
VWYEHsff1BlkEDJcHgapGP6Mr7eHxsG4dNcgczB61Rmz7ldFB5t5jzTs/KgPnf8I
pkncW8Y3gaLnky5ovmAnbnPbvLhvTJjZXGqEIqs7N5+W2u9TV4zxMmUI7rljoD2+
SoxQ1JCmyXqqWLTd3BCxVcjdi08VUkUbGKZIDR1Wm2nVwnO3s94R5q5xjgfZL+AS
i+lBPAMrYR9mSNHwD2yGGAxy7ditmtF9Ah5Rd1DU0fQ61219BgUFzTM1Gbs2xJ5D
Np/w0SJE0jp8FlFueSH2WNbpKahgXnewCglz2Zjc27itzNlkZGCTOnGL4iPenkJ0
ogsOJd0Cmcy4SY5lGaaaCS2IHI0oustTAmG+mP1CxmgbZwGsJf3sWWGKL2P/sRS8
Q/T5ghQKhEBzNKtTNdEqRNrmdhuqm0zjBt3vBE2fJvX4hPj96k5fi0N0exca6W7+
XWZgAGimiWeN+Mpig7IJkBY84YRE8n7eVscKJVVXGNfKmieqPIdRx6IaxWcmSrXg
UpWcx2j/kCkrmiM5jSxqPxwcWTwljeWCuLhsYkmEa0SxkwEGnawUH/06AqKesWgk
7Ca8+AryrrzLqN2shH06qOfPkwF2KsH90H3xV1TD08On9Zt026xGfoSQva9zeg3L
dW/F1EJn9bNPljlMlxi+w6pwzkuplrhvNYODncowqdY0ObxQPlHWz/AQqAwHHDUy
mg4+wzhlHyCVRMa327xaPQnwZyYwdW9lUNvUhrgHkyfJzswkF8znJvwbJMB9bfLN
Bkot/mI533KCU5iFngVoMFtfrsAIB6YxadqukeVJddHXg3HpVBxkoQ18N/wvHvOU
Qv9FB7CRjfFhXKrCdNFDFa7OkKNhfgL3WVOkbKPKv6gdDcMd1BWwFO7sbqVI4hG6
4Dp/BF+eeJpPKYYR8R2xUtGaPtOy8VUHA/+O2H7/U1HP4y7nbZmuErYd3eCVbIXl
RahpKirBkp99LbCYHDjrDYGCIuXs3vYi94UTLKI4bVcWjAunF4C0zbuqNlDlzq3S
woHsKrjhbjlJp3txpHikB2ocpwnWlPPTu6rgo8reWHzQ2jsRdXnILJU4lrwzoNQc
UlTNY6XcPRbF10GipyOBakjUzxdyvR2TENsLZ6OM5JmkyZLh0UybDt1IqFPIdQMK
1d/mLABqclqVH45H6d/m4BIdNNWiqr2FwPz5OCR0TlpJSzWU8pSA29itkoroiJub
bVCM6g10ifSyWtiq+G72lxJvwBD2jxmh6zra9uUG+bI1LSzSeFqBON+T9XjYM/6J
bk2q8p3IqKnpoKdsqJwBQ0dyO4CVshc0JjlWrjDFhpL8MEIG5JrOcJ5jSRQHtUB/
35znn8QuEx8y6BY7n5BR/oygUGjDuezzuiqK8l/Is0Pfsu+zb2q8UkaHizANudq3
6nZn3CyF7owmmALJcba25DhtBK8ZlOL2u/oMMdTOAKAjGc+5mXVnEauKvBFduOgz
BS+ah3iszditEAnly91VA5YB7OZhT5lX2CEH0PoAM0gyxe3ccmBxrMG/d18z6cxa
OKZcOkLqezjxPYOeFqtlFFfAsBppv4SWwgngUA5qOgQ8igpb4vhDpixRXNHPMktq
v0JPtYipDmSXzcrzikc1+Qs+GqgifVRDBgQPzccUjL+PtVLipjV8jxFRCwEfAkkv
k94gA7HkwZHK4VC6JtCEW9n21wVt4m5uAVzU2AQ9rcVT9eZSCrTDsxotjFtI7KDm
KhfG6uTEq+kMRhalyvFpVzpFdO7LZlYpoJZIgpDqs79JTf0VSZIooYZVLYteDpgO
bQOxOql6g4KoGoqgsvjOIg3NRhtlypbEKNj0LSwuzevyywMS8kFrmTFurZz/zBbR
/OLC+I0K3t3bKeBj+t0PfCkKthcjewf/SW77/2mPUdddF8VBZsFqCbVGBw4tpjNR
W8b2RtasDLCZ6iVem2i7r7AiFrTEbHLSfICDbfPubHlmk2KjBWNDNJfpA8OhnjRf
pScHT0LUOxfzRmHUofOc8gtvDxm432Yf2ffQ25N9A84Kokb8VmEEsBsIEZliJvKq
fijZJItawNoY6aIZBO6evE2i4zO4IYqA7v7+wSOxOePvxqbQxiGS6PsNXsC5TswL
BrxgaBhhcbTJeSgLgsA5ZYXN1FvHjXapR4rCr5ez1/pQRCarvrAnXwA1TcNw3jy0
qyYBUWuGK4CEZ4zyHoJ8XAl67qG4fgcUNdSbmkLYHmX9Kz7T/g6yBTOGdzsDhRoO
FAEX+dsA9x0WLmFciG4n5KKHzRKVdQj0NIbmLrgQMTEgKasPcN5gG+ky+yQHG33W
PPWmiDVnYdlHpJCqtPGbO9xsbfFxa3ZM/ojJiTH/xzR9a94gPfpsHWD7sQO9j7fj
ob1yljSL0gC23qNIhAE/iiLkSmwhQQbLoNvtpwyzVP2EwZ8py99FoDSWn1xPS/0/
Sv0ji1Om4mhtEPzYjGDdWBYitNxNalaXEc0ZqeTaw1Qtim0P4FQ8ZalogvNYh8Vw
SlkOBlm1OX8a649YiiBjkYlgXoEMrw3i/nFqXx5yEkaU9cqyaFEVISO+5j2nqmTT
JvuAlLj8EGA4yzYs2FPWLBlhw1++8dZx9eoF/x+gHK3V5+hOq+Z5MaErmnDA8avZ
eRlT8ZTkQML7xxbPtA0dj6eExfL8A5bLc97lLqz4H8eE54MvVuF860gTrUdpD+4n
OG3Z0mU7R7Lii9mKcs7nqo6/nTDjQlWyWLL5J4TjLKbcyjROOk8aSDc3bhNt3/Fk
6CQzZG++Lb7SXh7l9velb9chMVvOqkfjnFhlt95s0QKQbzyZnJnfxMjkve/cIt6I
iV8FV80FKI6FluIwvBtN1zBIP4px0rCNx5IavHdBA+ui1497Vb6L5zQPAP9cjfIt
DU0Fnd1P+5CpbGQhFJUHuepIy9UvMFS13ZBQZqe/fXcQKXvasVIWxwJdMQNe7jPu
AQkopEH6wXXwQgUyBAV7qJ3jtDsPNFkC4uoTMpf/jitfaLQLEPP1g7YpqiUHOjHK
7FhMml8ddT+Sxn15JRvqLQiOFSCdUP4TFeIyl2AuCTsKuuRrlVPCyu1kJfiQyb/C
xhPTjNuDrOhyxPAPK4RnGqUwntSM3qP8s/WL5mIu1g0upZWoGPKMasS7AZzafByq
1cMUS5bXoRvnLXRMKtrpdWvIv2CPlHozDnbovPcedKdtjsHkrKAe89l4DkFTss/S
ZBo49eE/T14SrvcQDvMywvD7PLmcJs6xkJpXIi917xJ7oEG6PjAn0c+CJUD+LS8B
th1yYNNPWM9ucRsnCkUqnXdD24+bkwGLBmOI0cD2iVeBbS8EnZqy2k+NtDDGBxL0
cmFQDIOEEg4glhJMy0yy51F9npehQ6nsJhPiou48EyT7dP4K0xzkK9ZZ7LDp6Q8W
NTMO5YiURdtV6oDSwzl5zY9EkSVfRcquwWdP0wu4XCf0nbt2HH47UteKb7U2UQ87
y5/cIEP6Rjrc304kWm6SVUSya0q9RJf02GoSxitnXZeHNSppBxsLbZlV2JkBxHVP
C/l2IU9PPu90CQ1/hAknRBZkeJBliXrxu7ObZ8KVrCguqAWlpPe7mcCSNG0vRvE5
1+MG4L+671HbyyNx94YR3JbodxkD3/z4rNS+F5USHeMiUNaNJ63IyqtqPH/qLNC3
rwqE6bQLdNxRMbFQp+2KwKsOZE2+CE61sIOUvLEMnTVTnw3QmpYI/q10eMSZNxo5
hDvAXJt0VGNXODWrrJv9bv5hLP5omHypwlPac607jXmciXLbI+vaM1uHs3D+WlPs
+eINTUPiNvli6eWykLQc0LAM2N0+10WpYrGoWJ4wLUDbjKK0Btxvt2LOATRCjaZs
Su2PPI+D+AvtIrFnE/ArLcbhkRiyZ3ascBHu82v5vcsxYCf7eIMz/HIRwz+BRnpT
ao29wqpA4wSj/v9bsYsmcgyOpU5XsPkO2YfX7LmjTw6TO6Ly+xtLtUfAQRDxSL8A
WKQ0xP58e+WLtspluElG5IbwgEeI1hcz6MWawH7BkBUrimiPUSC17Ci0XVu93C6F
aj8naHLLPAf6yFVETQTMq64C3BOC0dc87O88fz8g8y36O0rqaNsHNKaRXW1jh6L5
rZ+WrOhf6YLm385l77oERek//0a0H652DOBYL+cbhrFo8GOR8U0p54jBfCuNRrwr
69qQE+0RCEX+ZBysskMqi4YWPIcDlv9mJC6CfShnbqyPqotC5WHhFVs8zbEE66N0
fKoKqUj1LGmJQpzRV679sWXp8+f76D0ZZhs1H3kYV0b/A8ephxUSh/HTjXH/2iv+
RqvcNoaJb93rrdfHNpcaZhte++YgQE3JRIQgw4uv+kS5eOvVPuMmwJtxl8nIYPtr
uQUujDNrftJCk6b1UrbZ3SGjzvuyTwtfUTQMLpGdeSNzHPzCNFCmeEryDziRYn/f
lD0DHT/OOnUNYX9gRrDXwRExptSU2lQRQa8AKnRBxifj10M0w0QfCvhrBbX7ncO7
Fyip+p9pg9GhlCpjuf7E+ltL24np+FQ0NWWW/BOsB9N+KOvrIojbClEs2sX22sSG
tZd+/kjpU+WkCdWc/C8rv0G0GygdUtWln34cHPOX0UU+k7JmhaCBwaouEPA9F4uM
2zuulgKtdPLFoE6/eUPSaJPiwyicphKntoawRHlSRkob2gPHwObdGyKtcfX4RK5k
SRT3qxdjvnmNojaKRiuIpSdgHDkzV0c0ruwR5btWsIq6z3834IIjt7ulA8/NeVCB
AK+Oac7foXeMAmSTPkL2f4/2PIfDsCN0fXIx2+WlUaei3I5HStUXCmF409zColBp
snW2F2Tf4e1D86Ur+Cmi2JvY/ubsgbsR6xBj+V1tZjoyKQk5q2Loifqa6Q0DWqKW
/hUuZA8KwHgZS0iDpFFxJUe0PiHg2vzwc+S29pvYNXVSWhXei64K49MaD/QS/wYZ
PYTc/qn6ePfu3AgLVijM4Mmb5cU5Tsa5V0wnpIV+xNoT9CnKQSeFwc3GXxDN/ZFi
/mFj0mbpIRjNPMBFYCXXusJ7DGa5UYYp/sq96oAwJfSiC/tl5IGAUDL74i0KTfcw
0cQxbsx9k/XzlPiSA0rzuy/F9Nj7f8Jyiv0EAM8gFYMVSbHJ5aQDW0uMgWVu6wPf
xRjqsXXg95wTkQjnApZ2DUCXV4QKQwlH2ygmhikpUsaN6kM/7jy3faVCsZ4BedZ+
i607edBK7wHWu65wZXGZXnDixRy8Cpht9rhkPvNnVzf/WVhWGSbugtsAf3BNEzdh
aCDvBkdiImM9hfbm1TjCg3M2hvWh5nLRp7E5CNwVsYsgAfxS6uflA9SEtYlomPok
eKtJNi/Uhka43wdQGFUrzJToM2s2RocWfBVF03IYN7ngN/+d6dY2KRSrDzita4N4
fXpNqAyNAD9IGra7iZdQkIVLBriGnVoDSy37oQxs0EwSZ32bpCPg39WnmX+di/SV
LbvcufsTyPhye0cV8hCwuehjOR6YNA+HGI0MKcjRSYmm6JXcQQxSMYm+un0yTcwk
pqkhD0BRamhPK5vyzsD2fb3RS11PLUFknpYPcmxiTMUVXOtTgp7LF7SmcnP2HFND
R8ppX0BImUpWTgYUAfDnK2yFXmTsmETtAh6vZqjk3FHl5/xouc19YZT5e/RnTQaB
Hyz7BxiKKQOena7CoFOspDwL3Jr7zqlZzY/GbyW09DEC19rVXPPSXpgB8dc5LZ2G
KQABbEn5JLdSJfiAPyEwvp1dZIT6I3pKYyNEKzv7cVsUKdOcOtTnwi22E90CIwt4
WvVz5qB5f2EvcZA5r8qJHxylX6xCUPESu3rLGlsIuV8whZ9KYAnUZEx6kThwR4KK
2y4tppP+HoSQUzTnv7zPFets0p9SaQ7w/S7azrSsn2ah4BMxFIbt+v2VPmKY43pg
3IBrUAUMTpeymsBT3QzDhfDMIvlADrqKODl8hpqSMQVxB0bry68uifYHhlA421Xc
7073EtEPtjalx5Tk/2tLscdtfF2hRYy07Nys1YKrVYV5IgXz09a8c2Rh7zpMBErW
aZNyqnrt7L3Jt6o5yvGQiHd6CXYoLBT5Zd6DGV02xoTfSWjm9P7IxjHx50oWUdDz
7+9S3hSr4Aa4bsbXMHLeyctAevOj2MZDGJy3//aD+w7Oe8FU5nVCA5wmVvmIBsSm
TgAy8wf/3fo1qyEbitGUtkE+Qy/u8IOXOqzRAgguFsJ1454mKl1kIPEM9w7t23ea
V1tIXmdUYokzrdYUxpVGeiZgEH7nDcTXwUeU93DIe+F/EwEljk1RQqFA/tHg+tHw
lXHNaofGz6HrtnG6tZ4M0Zi6AKE0R/6kOwmq2zbmC3HrVWIAnMY28jEML2kYV2OK
PONUTypQ4qF3a06hPeu4GIpKi6+SsaRSTpqHU77EMg/xpV8A9NDASgVQ2jYHo4Wf
Ouaw980Gpfga6d2Yywsg3AdP+2iK5naJhIdtT2FUNitnrYKxGQbIbCpl+1cqMFCr
TuLkDeyK0OGy07byWTI70YtAqRjCTbrLErogqZHP+RlxS6awF3dboCG1to62Nu2o
cgYULrIJvkpFzWSTzT4iuCz0O713YhIhxdAp5IszHpe9NaRVQX5DAG+ccPqbStMi
+XDos988lHVjtg91Ffc3ziWPD9yfhLAmRknlLVoKMx5qDxvgdNvRRU7tO0esl5ah
MnUo8emT78Jemmo6LksCyoVzCCSOeJW0ckwjEVcYvIyXuWM1LvUHaZv8eDyJH7oJ
K7YY1xNIKlADPE1fpemNOuRRrdy3v5FHZhNPR1NUts3zoKt51vIaPhJ2jsvSS/Do
NAJgP3X69xS1uJT4HaYY9MzbSxjqXJJj4XaZ17XJV9C6Jko5BAtX9PtAm21S2Ku+
MMaM6ppRaoLA/X/2N/A0WxT1TnUCwLztjXbth8omQhsBbt929WwCA2txRW3hxNyO
zxP04Fxpv4EeA06kImgAUinGWd9xveHV6MHmbCTBmNEe9EQdUMxA6vsCVFvMsEvJ
iZmjjgHiNzsNCcxlCYX+xLX4cmHjmRN32LKlik2nkOVEZIRYCcPZ6LbC0h0ZMV97
OqwMHYAa7yN/yKjOaUul4hfdaFX4S2rb5ERGtZdFZieR44p/3c75PpOebXox7FZ5
GixNfvYCba1upQdjgjtfGZQIwsHk899B9tO4CGEXdFswAADTfPP+qXEUvRjkzq4B
PqnQEZzUdXUUprbib3HR42L892HZGRZ1VZsgNFs8xAqyKDxn8ymN7LSPvnRaESG8
17niBd6iTqWwKAlJSTEXFAHnH28hUO0Jc1dTIA03HI7ET8oA7qw6re7m6UYUDj70
/E8QKjHNO8II+S2o3X+5eCw5Pgn2tiLM6BOUeGmglw4iXGG4DY90jnLT8g3W0/QX
Us4f5ymdZz9hnIuf2WN+QO+zq070IjEDamKXGj7duL2SgUmjDQERlhFV240oNoe3
1qeastvDgy01aD/80152jbOvNriDwWPHp9UpCxoXArK+8hqd0XcqY1jiPHstPWOQ
lnPkQY+MBJEh7p6AmarB7BFRC88iyU8qmrS+42baIM47a6l51J6vB0uUPaBT1qT8
IuAwFME3J6uiqiKpjvYipLraZE55HZgQrDJAXutwykaHWsSRa8C3e3KN9eb/xYoU
OgH92dpo17fetCxH6tYOv/E8VxycGYuJkuCalpehAx4G7hLNpSCnLgxIPjFZ23DI
qni9qd9t3iyVHzjVIQkX9w4k9o/Tl3yPLoMrxwLS7XlPxD6NntJLd5Q0HP/Ke0IK
2p8aXZPdUhLwjfpMISM3nz/t+Yds84UMX61+rAzthNaEZ85CaLkq8jh5rOJ1w/rd
uFCnsG+lXheHz6vbInVgjuI/TiZ8N7i8ioPxhYxwHaUJBOBEKt6sjvW+L0WZ6IZI
kwP07b3y/L0kivj4q0crGTL+afsKDMoEdEZqHZOABCpQS3yWcISKk56cEon+PF26
gVMpm5EU8s7ffkmnnzBvbzomHHF3uRkDUYz9Ez+Mntd6DJ6XXtziM64+LwToqmAP
CS1z0bL62qKNktTQlZdY40HnCc9t3m6yAyK8MwqEe3iRlMPEwlS+IhiImY636H+E
w59fF9moEo8rbiEcorGZet/A/YzXJ6agcgtVF7NFfGf6Ziv5FSRFa2vo8tuehrC+
g5JlqRxSzCW+2xnRtklHHWvndMlPMZv0nFVgK/iWw72lIvcXQfmCdcWjuyrYOPxM
WZZbAEKgZ2sFGRZV4RB3clGHOaJO0N00Dl798WszrJD6AWlAwy6Umq7XNesyfnQX
VqbL309XjPCUhcOHvTO8osBfd3FP8H8zMPvhZKZRylCb1K8GyOScEjOLJyZmBbnk
ZrZaSYcoBGm7DtuKZZ9GikyzoT/Bltsxmxc+ZLa5Da3sJfwaKZER/7dD997jzd2u
a34BYHmcVt+CoNWgg8f2T0CSZ0tkAWerPF1mO03IgQpWTjwaRXySma8Rh+nku1Ng
Qgftimz0X3yob6CrKxiGqnBTgAO4goIYa3ODQ7ZUNkR82tt9PJ7lwTbO9257CZ++
2ii5HOvvomGFyBZa/+swoGkzx+IKwYCdeI25keivLpjDkddQ1WnaRV4MgndC8LBA
W51ZJQOFc/PB5m1a4aVQqdZDq+lhQro1bZIwNIqRYwfGjzOuC8OPvBtkpu+eDVtR
On/7AXCZ/mf8lBm+JecyGkWj8ytqAbXR67N2oCLOzm09GZ4xFma7UPsHQA6kVcDr
DD3kTILlOxrUeX20koI/iAi3q4/C5R0+CXC7R11RqZtXPfz1t9LZlLYnPaK9EyUX
aD5DOhP/y+AdwyrJE5pWynxfaqEQgvEh90Bc8ekM31o9iG9dj5G0wW0hD1J/qPs7
LvONqN6fAQ0rJZmbj2qZM1dAOBHcfLsQealALi+kWebHJc6a0Cd61WKMF3pjF9rI
JUUErf4Nh9oALtkCRHYSNPu+O7rugmSWhtNYmoUzfoe/hmO8firs65tuvsSTBaST
7iRSh1cCOAWeJUPm9oGUOsM0B0uH+cfGsc4wcQpNnuYOaBs+n7ygACOhUdd5LKmW
K85KNNqJL5tWpayZxqaNe6Ujr80Kgb4zBiJCnWxxTRdqITHEhRnyFkETcRULhfAA
ftNErL2yzvS8UDJDnpcGT7+S0Oso8k8KzRwVOmuKn5HQnpXzsyF8RCpE4kCa4uN7
2nWQECX5qyGm6skiWaluB7RMWyKCOfBRtk3fLWZrwbz5Q+K+/ZZnudSmfi4yHKL9
+psvWNrfS43pbvo1U8vty80VKboZAj4ndf0ILwRrV9D4ixF42UX7UkjUsdrqM1oN
RPD28ZNLQTL4Ab3dq2JIPhRgBAPAGRO+IHUe4+tyImCZQ1Lxvdb4LV9K9jTLzNwi
sI92eYsPDTE6kEJ63MvG8TccVNwuYqIMfem/Gh+yjXi8fAT7y9ffuRCy+IOjbUBT
YH20GAx+rlSkwqanDdx+zzBh06iWiI7AFYcC2RSECrrtCCdjULZhGh834vgvgRfp
NUjSqbKH1sFgIcSZ3NWjpAflgXOFGJdisZvctOqSgFDJ2Le8ftotC/uEKhDAAi2R
kZsDrtloFy1OumCJ/GpbxykiOeNMpnIlAQLSYDKGFMDIFIOezObYDfo262afPzRu
/fO7c0j1budLAIa4IqeOHhbitcAQ2O6S3BGOBLQ4MBSbey1xlvRgR+itqi5C7UCP
5GpNMGRjlnoptRHmYTFvhArH3Vv8MiiC73/+NlpfzKFV5jOHThJYqCkM/NsELjxi
7kBxzEahGY07HZrsOf3q0NUirw1ovd2e5JuKOD4DaJ8xVfhS8HJ3SRu2fMw4OLRf
aHlrR/dcKTUx+1+6hosowrTtGeV6n7q0WgfkDCE5ny8vp7Hdnr6PZSWpVm3RTSW6
2G0q7JlAjfco6krQsjWLu4/sHZYdBn73YS29ERZya+sxx4XpbdlyNlDNarK3bwxP
ppNczkkNUbl47oMU5A63DwsvqGjYnEi3utdiXysYhDdn9CQUgilf6SzaRePgbBnr
nNwzgW+bibskjARcFq1EP0q7e9igcExSPPKOJYB6JljKE5o9sqaTbK4rsEn523lE
fzAT0gtcTppJo43+jip758NPT+P9YEeHbxkGPRD8gdBhwrTWpzoIK24TMyb54hst
46LKF+hpp7IXW67XW/xPz1dxHCkgf+nmK2buFXgIqxrCIC64VscF2yZdppAbNzly
z1d5DClWaJfqNf1r6SRL68ISJryssY5ESRmstAE0m/Z/4BynIFT4yjum+V1qTNJI
NsW3GFs7Tp/IS6qtxj0RNbImWfTO+0tzhMWZqN0CAp06PbZrkgm44dVqfKC6zorr
szBcVZc1zE4XQElCBRuxxR3mIXoEo7XU/YjEFF5OPPwpik3f2UOvOW3apxlctz4P
HhAOTXJYkySVMZQW64WYjkgDOAXA/qcb9v2jIIsdj2UXNK2KQVrxL5hgjdKKROM+
iWTamSZ4FROMd0Uxr4knQD+M5UlBV9n3H8873FomdBQCizOmeUwqaJZZVylcpMij
RB6Qi64oqJI6zQgntdNgCJyf6Z6DlMc5VWc5XaOdS88T3srD5vKgT/4J3wlofS6e
PiAKRPIiMgpd6GIHuzNei8rHmRCCi521GI0yqd9ZN4Dhk3UB0gI5WGfT1+yJNqbY
GQwTlpn+T8COmlvbyV5MMe+8wkony64k3Efqo0olotoz+oCWo9B+6NFzieUPwxWO
dq8NFHtJCpb33lsYr/BAoKjCINKCtZXODv8MTTRYBSMPrdjX+jkoSTxt/vJqG3a2
kyutnbUD4IfiHGpN7CZyPvhxAc0XSpg6x+z2HmL0kNOAIY7+1e+JlqIw3BBenToT
pt1TEoqbbGJ8fY63802OgXNoRkzvHo26fUoAsw5xHwtAZaiCUU/u/ieIDL7YdUJS
U+z0rBY2gE+S7XH1SlTaFRFf2unc1pJS+U07Mz2CT4O0vK27KiA5Xux7266e0iAY
uuQFHv3Ml6DygR+tAaoWZwp3yjIF8VnTRf9BD2WD9bmqRDUyV0AF2veA+IIG+OWM
bNyMN0Bgjqbc0+xvZWh02ZNNkdcE+8+2HvmQ7fBQoE87BLsMJS+tW/Ux7XaWIjVt
qLz+Cc8JhqCxRjS4qmEQmJWWNlS0R8gSVMTvmE5coRQco063gecAJgtvDm2JXnn5
OGoGX+DtX9d7liOnJLGRJsAgLkeVYghpk25XzX7cV+JLFWqYvyBk5AjMrYIhgjah
Gk70yRx35DHqMd4Ci9s3954SR+8IsK8Wlq+T0qgAx66wwYrwmLxVYGXqOKm8EODX
wFORHobG59E0Q9FPeBXFHJY0LqtlsRx8F1z+sGEcPbarG/M+t7kH3yeSpGqQlKg0
wD35Vh7F85Do7PkNfCNH4F8OTL60PtTroslSW2b/TT8DAseWc1mUMqM8E72Ir9z1
PBpJdiQHpotA2GhYwpQbAOH4iGZUS0dMoIGGjV3mcgOSOoSU7CJoZ0Lk5ioNUXKL
0dp9rBX7ch+wzexa6imWPEYv3nYsNDx0rlIYqzYhTxeE4elVmDcr55sUBufqHr/z
VRO35cl2madSTitSGt7HUxdJYMFvMg3mCYaw/0PVeICtNBSV9sIITVXVWhtj/W0D
LRWvyISqLUn4MvXuZUYx3MTdNmhZWI94ZjeszaaSb9aih04o4tp3+eawPF73xI6w
uo+PmGa8AXhHwuPHoLMZ3FMHi1XEOAxMEKxl81cfarWA6TmQyG424D7NHWNnP9y8
kFc+YRkTGAV9xmDLlZL1v79D7R2cdSkR1HJIcyMmNz5UFCjT8ZjkaAo8DxDJ0FFv
lxGHHQ6aENrcpL5BwfxrE5KD4O4pCjWuTH4bnncSo0soy8xvDGZAKQRRU8kA15Jz
pKVH598/ozFDD6WDuBOxLMlrky+87WbzNAEu9sKkV5vI4V0mIha/xF0U+AUvAoot
LebADNFqMPyoH+iu99UJSQsvDxQcmetfgNRcyFn3k1FhsFzrzTD7iPsEaNPkgQ25
+1janH/WHTIPfs3tD/IwE+WiIbkC2iS6kYmEqEm0TLjKJ6fZ0exAC69QQMCtUQGD
AufIjtbtTpZVf2Y8/4+6pen/BGoku3i9tVQhmXoB3+r1a/JAv10TUmIaweBLIhzY
WJCtncfVGJj14+hLpdhemfbpp5i/BMcC/3Ue1xcU0OgS/3wDLJNUgwmA6sKl9Nz9
bElIM6Eg3TBKCKQ3wTCGfHYOqvx6bhnkhIlZ8uieSVNfdazyJZmAAZiDp8cIvfT+
zFpJrt6sV13RHnp1mZr5b+8JUCwsAysJ6tuGdRTpE3sszKSaJTl3oWdxTP3uMvbU
Z4z8k83ZY6EfWDoseQfNMCjamXKiJ5SuXucBk08n7bQysBibiUWoNjz7aJcJI1sE
otIOxRMfkUOaUpdxkUHZpzm2xqyl6iCcr+iig3Soi12oTh6DC2GuQ2o60RubM8Jx
U3mErlIwFsYGdEKUGubDnWAnjhICqjZG9P0nQ/GM2DG7gNQn8mCyc7wVH+xRR+s1
ZonL4s6qq4z23kONxEIn22w66IOwciYrS85ZKSqpwsnhdJy1UEF6FrDmEq18RS3w
4AramHtU7StAvdkNj48n2kNRtURzzvZq89jlOTtXeFZHLEN7u1OpMilUAZdah9HF
Pz91yE08lThM8BwGz3+yBbcErhQzekebjT3XKDBgE2GEvKsnLeg5/eqf8yqDVzwp
PmHoHd7n8qbRC9ZBjsRno7c6Z1Zsesr/dwvZqcZp/RpYko7N8Yex7ndQKiSZgO/d
jbd7Wv+9y+cO53S33m1qv4B6yDBm4r+gXd7mEeqRDadAZI2r4ydaQPtQfCluxLbN
NrZv7sKFfbX6cjWrK/pCvBguZkJE/VfjBWr3Dz8LUV71ikOYoSg6JA8HK50xY5Uy
wp+iM6mLG1VS14LO2lEv9iQH+m1EP/tIb+dP1lQliMjZmGvi8oLMQGAAAzJF9+/S
4dP54STicLjTIJPincEEJFSFqcZDvPar5G0vvONwojGF9EiWZdh9f+8ZsM2YYzZS
4Nr5xuWpj9TtlOwlvDM0PXC2WFd8aHxtB8wplvrrPt8nLM+Ry2jOCS3viEX/N/Ru
+6hyreXFzwQvRsMtRx/8eOudGTc+zb+bw8Y1EzobJvGB2cSHtcxHZjqnYtltO6DV
kxQ3BWDENeASL1vg6C8yLCTIZD7IW7IX9Z6xkhTP0EHX3wUZucPoRCls5v6+t8t0
zcRLPS456r4J0qbq/62VK2/2gIBJwOWDoFa8MBhbrw8koY8vJj6o4JCQIOjGKIzF
sX3qnXApgoBVMdHgW/87ittg2SQo//l/s1B8JviXT4ipORDCYbI+5tbl2ZcgXlV8
C5i/yJ03hTUerad/dwaQHCISMx65uBH6tOAZ9VmGUqXx4gzkaOiIYwzsDihIGs6R
l0OqrVcxkQyxB4jCej4tSXhpsmqaAByysqBmN5Q5V1l0KgfhV8pxf64JMI1zbuIj
tX0sTTzmJmH01kWrXj+mxw9rkaA4C9Xzh7Ot0pnUmNufYEnPjLxqcFr8QIqsGlOi
Owh7sTuyjhYloItxQTfhEaJGBIUx77ptKiVOlBN/G9TdLArB2/pl5K93p5PEj7/0
bvrNJoHR//joJTAGHWOYbguJsE9+EZROfVtdDWBL76P3fQEHqfqAhl8CyD8cgnIL
ChTYqTLyrWRRXjY08kNRFy/37sxl3Ue8ZcM2W/bIc5dxeHrERcFOUeK7gJXC8Uvy
FPj/9mQd98V5MJnhVCQaMoYBi5YRgSPxqdHK3gXRSdGzFCcbzdVDrt3NI+egDIx+
jqt8kDzPyUYbf3MmksxSqh1VCTt1w9dQOhTIhRemYBa1BuntSu/zhg7Q/zCmYDng
PVgadB4Yg+WO9o0sT8K20DdMq7r+C1C0tkWo5+mym3E6zP7gIK/OyugOk4nHtbXQ
3zxGDMJ6C2Jm6HJ2V9WlxpyQNNQYDktq50Na1BwTuJjIHVfmXdaMXSWuXrhInWOA
iMGoysBakdwUT8XSwvW/5C+gpCwK4Xp+Uv9jcOclkr8J9G19YgQFB8ZIpXUoQQNz
f/lUIcR+WAwsyJ0aMBQ6QnnsrcEoK2QAwUlhBygnUqPUEaTBEGR8LJv88IwCVykJ
uKCHJtbAptihlsZZzDV08KzHHBuFlVNfTBQjmkwJZWfx8twtYSaH1UDWoZpauFmC
Mnn6Ytj0lJZtEL9eGuzmnZBllruvP5g7GWY9ZF52W5uPbQt4D7cBS1wlx9ZSHEeo
BCevEXNNqcvYNNvRa+rh1bjXpmTUct4hV8+wXy+wsc5LD0RuEPoYsUg30Ybypv5f
X27xHytOSnlURcpV703Cc6YPzb3w0qsRZec2Huyq3uJHN6OR/Z3mMdvBGdlOGLm2
3wHDAciOh/4xZbMuunLxpMYfDT6MHNR1Xdo942svQ2sRAZ7fLFqIZMGRrjwi8hpr
KG9VT4rbBdZF+jfYj9DfHfMpdmmQS4WXAwtuIbDGfeuUBaLRNpntzu/USy8lOxZx
i6pdq/ZGKMcCjEQbM6cAVEnxgb3HMpFEpuGxQSYUWozJWOn6BAIHw0NEYNbw+OEc
5lgEB9skps2i/nidAEB0LizUucDxxXkkN8VmzvaQdykM5W5O3HfSfI3iJ6oY3l3e
+0SQ6GjF/mvjRJ7Xt6lySejVKFJQn1Q+3LDpsvc7vReyHlbdDKka//Lv+dl3JRhl
LkqyRwFMOOVxqQmiXN9PU99COqklE225KNPCx8GoXykoyW1Pdq+/bQE6X2r/vVgD
RXXE+4vjSMDrsDPn1DEaTNeR47+d2RVkEoEZvpZJbpGs6XgoR4jjsrWJqd+gkb+l
/QgRECz5wPHjz1N9rV/JDTaRBeC2dR2fqEkBPaVf8Q5/Zp/SjBsC5XCyHxJdsTeq
TnrAOOZtfzAn4srlHgq8oH2rlXTqMRaExbXDbkQfFiZdttDaqeLIN9O3Bl8ADFOg
nfF0QR2s2pQ3zzUuH0K5TxPdy/ZDOCaA0FJN9cImpfWIG3teDeMqi1wtpQl4j2Ky
pS1eY9vUgIahgjlsGosUIndBFtwtWhgqqLAb4Wt7NAMjTWNwmJjr5KwyoJ+AswvF
o1vRjgAYVI37NVVIVBlLhfO3gn+55IVAbvFl19vBHmA+BvhxK3EVagLwhp5Th9Ko
D6ReCAY0Y/W7Y3pHq1izBLhhAN/2TYKDO7KEZN0Ef4GcysspBv3Pl4arpQ/KEASa
JqnUkhldxd38zZ9w5ruO9wfCUPuG80GH3ee8Thzlo99CTHDhYmzW1Ae6mIAxx4cl
nrNK4Qjkw+q3Zw/VIQCg9ygVYx1pD2bEfiYxPSIody63mLtZMvjC/oQpNzhftutv
bniH5NQupi2sYyKk1QFqcG2c5peb8HWKVl2gmkWRAwpH9sk+xRTt3lFElv8vr2dm
KafYl0+MsLmKiscXwWZXjhE3TRT5bTANPYmoEokgOJItRhptjtLKj0Vs6Mh5JaQ5
EZn1hYeZu1Sln2lIjsfWdnzEZbCwsaJXtm+LAUZuAVEGgUUoB/se2VaZ1n5njjwY
v2FpjlsUzIzvS1248d8p67v2KmlaWIzwYH48PBDDBxASbBYnYFGykG7w/C8R71Se
wUY1faioK+WbBaEJJpirfoBKUU8SToAV4R7QcUclZ2sqK/4K4l/t90bf2HrS0Uv6
sVDmEQE2rXiqLxJopt9ncvmUQ4GKCTmBPJFPlMgvGErsf1l9hqH+Nosfu/zykg+e
IENbesVFi6ZNzjyRjlkQfPiTy+ct3gemR/4pl/boSDbjPrJ8Jj0e4dZlbAxdYTO6
f7k5OMYQuR4iNEk0ex9xdnPKzvPK3AGqIudn0xg/YyhPSY6TLok+uXMwWE/LAEF5
tjhtEWIWW63yV4dKaj14KCDmwTMr/4qcz+3hCsoNCi65uhk/fQVTgKyjZgLGE/Uz
MEuAfYGraX1yz4gPd0WENRJ6VEESKAUD2HtbqVw8yF1hqCrAC02w0bV9ZeiO3piX
xXVNCXgE30xmaVDmBmQ6T5w+yjbQHJAgY48kMZSvGS2r6R+09nZJEuuT/r7OvgSD
xNZ9o7eu4dsXxgkyJq6lxGBKHGcrFDpK1F5zMbwKykz6eqlE3KrxwIg+THX/OuFU
g0FhscsWJ05bckoBqvndwimcVxfpmCdTs+FXfhH2L+ctc9Zt/Zfdvk6czJEiHRtV
RVL532TnSTO6Atmum5XR4Thp80qFUN/a8cvQ3Cjn+sa+vlNTo9eXQ23dTYtz5WtE
njgDBb1QmM1NUGY1Rh+kNGh1bcgrdb03zm3pysoBcRuSkiffYNOhYslZQq4re9je
Nj7BYujqjvZKjdUvLDe/x7Zh9CDsEuFZ8smel12JN0NLxblVr3hQcys563ZGrfuu
djKTN0hZ6Fzwojr/gXqM3I13HUdkfLNlbM4ulHxTfzCxxzW2k0YgNU0mg0R0xDt5
ulw+VGPZOkEp7fXIVnLEj0t9Mc0DZwbAVM4ftv3GerCLuf7iVHCwBXSxb9WsiPmU
rTDcOch9PsmUbkdLXa/ARuSM4LnUzDRlu3alXMpGPgJLxbTEcgxKcj8wbU2r6XrH
X0dJqYL9IvTpUABsdoUYZBLbvh4E3AlUursYRvYq3ZrRg/aFcRs0TTrsGNh78+/4
Lm4swh52n+/e9FHr7g0RyGcePxCSlEHMzeXZb0hVe9vtRbAySVNoh15njereFBcH
y4/vi1onpYRNEqcGuvbNO2XYF60AtkDe2215Vv7FI0pwn1uX9Evt10VlkZAd/xmy
RNut/l4am8W7+Bdm0fqSldxgvtU3hREfdcY9u112zuN7pv8xYlTVYhSiCxXn5z7y
yrQl+AlVOALsCQDWEgJhzO0frSg8psow+RnEcmxY0YNzw6I2++8gaO5KH9/mvKES
3xp8qRcjcIiyb1Ye4i0Zaun3GVfIBBSQG0pqXv+WEKfc/7PU8iPiZ+3v/M9xMpRK
2h1vBtSYJfZNaNTlIvJrkCbk/9pkCMZOnbvyADL0ewz8puolcdQp1C4JAxwT370v
t4BfsJ3eVYNP4QF+vE3J12jJREmvVL5uTRUO6Vrcobf/my+KJa7XHYGuApKXAlRW
xdmIOlmsyoz3FmibB7NuoseXd6/1ijirhDCmrkWgHTDvA6SHbLJJJgZGyElOO9st
mg4An+FnQDcXgLl44xWRfH+nS49OV/5OGj5jhoTRTEm1mQQ0KpuiIJ6dTurMO9ci
OUtA4SVSKLaKR+MKhWIfDSDH04lI6jL52nkfDNN8oC0IPJGCZtoNEPBGFHXwky5X
MZAr4rJ47BYHgfE3T8ZtuK1Kih/q0ZMRbO9Qgx9giPWTuINPDR4gxibX52RORgzM
zsdLuSVa99K6ZIdEHDaX5lEib2rAAKcAyJiGowGbeL3/YO1v19n4iGPbxQj03Cm8
wqQlzCXlEHQmvNQ8oqUDYxqoakOKgwQdG8VXbu1LkPEDHdKXRbIDk/L097O7sL5J
G6yymUrZ4yP7I53dhTp1XcL2jTpi0OlpZpj457nMVVNuttzJ5TUlJui63baxYjw/
PPhbg4OnqC+EuhUlz7J+Hx1Kq/YA8oifabnZRTUwLhm53kOwEkccfHBoprBObz/G
/nVCX6yYqmbJytUI7uX8q+sboATncgjNx7VWw/t9nrZJLrH8sRcxC2PPWJj7zYNm
T6SXUmby+AcZoRrxrpOW0v9IKtJxKT+JzaCs8LV1nXp5w1hvrbqdLYUQcDXmhpQ7
tk2PA3AU+hTN5CtkupB9M9ZbbRTLtodpP2BuEbaOZVOCLalFJwxgqrdiFpfmQOLv
I1Mpa8VIJ6Wwd7eVZvBa74u/0WuNNwCK5dNwm1o44CXv9kHGMuZDzY5Feqca7Sgb
ODbZYc2CTKdM+g60ZS0zkY7+A6GBQNSWesE/vr+8y6DbO9kTIjhc4MafMal+kF/6
68vF+FTrE7S/d3gBcRWiJATdbT5csDLqIBXH11WO9Gl7dGrsQymDENgJC3wxn5uH
cKrASRg6VLr1jLuC/TBS0vfgrobWz9ElLkgYsF+jSdexO4RIe7EvSpFk5iZ9IQI2
ixB0pOJ7LKRHa8gZRQ0QYIWbN2CcfB+OFdluhb6KU5R7NriGile8IGcLi8FdFFug
rrDnfEPQaJUVfeaILusXZhv2ioZs5LslC6ZoJ2+fbrWW6Lb49Z9tQm0RaGWwbcsh
L6tZlI5rJNnRFn+YHYqJQ3yGaLhdPT5v/z9rLApiumG/KsAzkvDDdwlb5WFv0Qhq
VbC+CxNuv0DUzCpfFK5DCqtJvcTuzoTwwUL76z8tAUbt1gxh/n6H3cX7IqhGsSbU
tscNl4sp3qbm/4R2RUdOfHHZepf4RJVkkJfzvd7xpHd+4fwI9KjOPNZCzmP8XPSj
Uc5m457EDmmO1Y7hGFJqQuLvUoZTXfilm5nlI04M4F6VsZzBs54kGXnzJIptSJf0
zqYIXE+6TTY37vGu//V4p/e2jG0tBa3DaTNaWiKxNvhVXSke8ScdOUQqZsWbSNIJ
HA0G+mXYT3AtLEewwQ7pE89FQIRDPgeF36WAoAeqYr7ceKpUV2f7i/ciZ/sEQ+1/
uPht+TjUzsfAusuKcEUX0dunks9hZjnn8IXm9AQhr74PSfdECv5tkZE17x55N0Qo
jAU6opGPpSJ+j4NAMqXPb9qOSM2j2KYB983ZsxBDQ2MwNUdJMPOHtbqNVBwDkXHJ
exzrAhLjBiVtDCcJkY0nwCjVnISCTpiiw8YAiN0Ak3e0y1JJoWZQPutWT4GqQinr
Wpw40LTh51ozzaZEwlkr0wjMEExUSmyRTE5gwCc//cGzOnr1DH0xjrwhowRUk9Ls
4rnXSgtg7R9pjoSnln7OwyFai/B+fJM1dxrahaIK2wM1oaHWMGb0NcVOs/0NIFlC
e+R7VbugoaIxQmjYAkmcKk/NF0WHnuHVuhj4KLc1EQmBlpa558ydOyH7rOBkaUfU
XL/JHeDOwhFh1WjGAqDC3Z1riRwQe9cEOJv2kFm0tUyI3fPDnIigLWSaUd+beVha
sSsc1UVzdhQndJsKZrt2S+VlimylRtbjonh7eIjF8T6OgdKkpghZY339/FKGPUSd
HD3S9qLNvG8IqDsHtYX9u5AZloUu86AOele4EacHWMlrFlxa084QQGAat1vI1SIZ
FUsX6fVHjhVIfwcdNdQwHfW/Iz+yXyYIxNdNCmleiRDHQaIr3PohewjAeZJeUK0Y
AS3xwilGVcIVw9+/yqHq4iXxwFn59Iif2eJUQaiBxjGWJ+4ETcPPb5vl5e1FdvEv
Lt011w7tkROJiq6vvvp+3QIFakkZMQrh+kCOuvIKI5cLZRbGP1han/iGbI3NFYit
Cl5wVZOTOUy5gDYmI+4UMcxMiVvv+XvhEs58d1e8a0Hmlj9XX/JOAHEyeAwSdcyc
vRxYZQsQ8ufv/iq8KMfzhjrokZnO1pD+l69RZqIzRd+4LJfp2LfYcpuoFej+f6Dw
OkYBXUy11aKOvS1xJH7iN58Aus83TISth40mk4k5Xy3V+y2HoPGp5/OEiBwmYZpX
AHQ3OYGL75D4nMhiJrvHAHjcvdNchvX36nifXxg50nIRSzE0dTJ74Qoq7qBf0gLS
O8ysgV2qAq0RMxVoDH8FGB87lBq01ne9Oxm8BNd9v/tOmNEy7CR9RizrBUytf16O
mMygtpodZ98SFP7sR/x+N6vG8Sug6ehs0twvzX+hB/yVE1Mvp1Kcgejc/dlqoIBx
VjOY7hY/CMxwZOKI0ZmiJsCfEq7bXPCBAessnejqJq8s75PPLyA9WW3SvuVNU0kc
LZYK9j604XlMQLwHJRwVXI+k5z512SlWIS/oAdXc6rEvE8EgU2dJ+VYHOyRVV/5Z
xB5ArV5/H7HqXFBrhw/1WFVRpvi7UdI12Q2vAULanc7eVrIsCdVPXH60I/eQflmO
V8d7yP+ZJnxZXGG+0RxrxulPl/aZcfgJV+6nCaO0k4Oo5cm8/gs3HgDBkSK6ovPE
JwH+OH4RxD8d7zDyXTJ6+1n8iamg2JbtVlW48zY2j65TMH/RA69tXrrqfNIWWNKv
YMLxvTyjRid840FLeZ1Zew1uwMvmD3PFhvL6suiLkAUzLGmJdWZ0dNwbP4KyELNr
UMBvB2I6YzTrw5PnD278DoDEF4GBa5fvNOVnX8ANPkOhzyptE1UhNSRyFf2FhCZT
CRkdzsioHuSyjEPT8TKK4Bai5zoTwMlcTsZh3EBnkK+9XJvOqGTgUqmxYyoET/xs
OU8v65Q2k80c8y4LNdJGLjZXgbs9oFspO6hXO4oUAuZdx7Lp4lAAsaI2wUxP0Xn1
7oCu13U/OCtejxZKGDrSikwmVRL4tJ34k8smkMd8ZHjBtqTTpVnkM7hrEGJgaETV
i2cQOTvOYwpYUWSReLsBAAGKYRv4pk/5TASjiLeXmNl2/uY18WGiObT1BTKGN8Fr
UvxFDDG53dKJRuHjoBAb/rZq21DR9iLBaTaV9Ds+BEioZd7WWXh6NbcBK3CjdGOM
PX1qFO/WgoBnXPKOzDQlb49fzD0GCEP4ff4NfJP7Dv7TD6imr85Ao6IW0Eu1lhQW
N4x558hHuE2VkyLHge5il16e3pZg8cmtoS7BAGxJSbYDEcFtBbrfHOEw89bkM6jC
nEoIdqt20+RMfccHhdGCq1m+dGBCkWHRIl94wsY94/ayu4LldjxtFC/JLW3s/81a
rafi2Fl4m1rIaaSZFDbWgwQw2Lr8SDsfUChTPkakjC52gaZpSbM2R2ulfNRhQlC0
yfxGq6fx00B11IrcsRmtvmO7vAyhSnIupDRoD4JZeyBh7vRQOdAmemaqIcoV3hLj
CDRUa7qaEALe1PFJXjOAdlHtw2ALUgoKL5Kix1jKS6BpNKcMPR4RGMRg18geGXKr
7lKmoigaD63XAT4GoKTVAiK0dH/YKpSVCpAHvdFn0UgDNbT+gmFg8AOXYtYE6NPa
EcBXX4ftrp1kcI3EkFME5BnBEGedxi6HNMfSmLfRz33S03+Li8dj8JHhdLg+9E0J
HXZ4DJaO8EjTRmhZn47RwoQqhnLfSc6IgtI0tWHpxpa0FVi31di/ZdS2qw82FxvJ
2PKrURhuwKD4Edn0htVHxvZ/L3fop8ZWvy6fm1F0fp+77tVZRk4TzOHFPnZ+u0oi
ILB+rqV9Z41ZZnQJlLtT+7Nh7MFP2JM164LcpiCS2fC/SmOA14E29L36iG+QgYGI
gbDwww09mUsa/4ysEn2z3j6l10CliZQJc3s2lC3yOwIppbO1nPFGGIOHuxl+Lkkz
4mc4LRf8KaDFO8weiuyjjDmHK1Of9Kp1MXJQy5GFZvLtc9FzCplIbxbBwMZQgFl9
iG+PcAWiBoOWaMCJEZkXwIbDZxajmt6HiQzyp9eqkaNLqNfpwo0Qj8aqMWMFGigS
GLoA3WG5Kq5nddxCNyCTq5x6KLfiERCTpRgeOfIGnQSsTHEdga9GWvzFVfUI5EVA
t9D0vKYNuqmkZcBayMqRju0RXgYGRjkMhfCV+z3wteItRH1KbpkRP5VQazjak9uM
JfkkF5iFa4k69hdRJgPDnptVbWWfeWGgsOmfXrYyTJJj97pfV6pXDBTRBP+zpJ2T
2VZeaBeeAJfUTa/GP5HtDXbBH8w/jWzugC6DoGc7XzCITQbo+Cpm6JbJ3F5S7lAW
2S2/t+Ge0q+5mikuE8uxkoJ0Xjd6NrzbsM3FVCMPTxpoZ769qH9N87BsIJfoFOI8
xtmeLYGSAtbaJfHabXHP5MTMaZCHSveeoHIMQeH4/pZMOFmGVMA2bEKQt03RQpdv
DGZ2Rqu7/Q1F4g9G3imsqq0s5jgM/YwKJPpLZ2xjBDK+OVOPJZ7X0dzXkBT5wSEq
qpLFhRJUJriCr+UdnThoRnJTqbTs+xluP488a0de09pII+3ZX6JUSKeEuUX4gvgO
p+BY1ihApnsrNhyX8ZpU6IlRNt7+kn1NemLI5RFVv5ye2P+btRLbFtKzbulsWGk/
Ou6bbG93FWqDRosCfdbIZSkhzQytlbqDW9buhOxYcNVcO1GXDSL7U+KMEB8E17Rg
0YJWEsit8Zb/Y82kDbLgE124N+DXnsp8g4aSvFwGtOXeM+insWT8F1FDZ/1FAixb
2bpjoSsu2AM6TpqPxYlQGUfCoUBWvZpr8vm6ItMTuvjIyC1L3KCXy6IYi24uzgip
1dSJFKYaOogbNCMLoOPG/ED3mObdrU4uZHhQ+Legl7Qv46vFpqiF90rXmJPbpT2R
jJNz7LmgTf78jBJsmeJ+OJgLp0N1NvLt5ANGx0oZchUyt04OxJM0QjYwx8V4FaoB
Jqin2VYDtXgtHRDjnwk90zAcRItLZ9kV6IaYa1o/L0i+88uuRlWjrFbxGLaYxg23
X1reYw2Eni0csB2vztOPQaEnC5JmboAIi7OjA7T7z0gOYpyJ3+65cTbhW/u3TaRv
t81QzZSv497dFmILFPh2nr2IG8xMpnB/DxYxocUvvCeEyI66roa0NgNbEh8d1T96
i+3Fvuiju2TFQi9yiRQ6rm5CVYZ7ye/q4Nv8iCBwyry9YJAnQvqbQkUG/wwAwG5w
s+eJrONr5IqIGvbd/oIQgcu+wTHjoPUZYMNx7DhU4TAFBhfWBQIjp0ACUjQtk0ab
h+/+QsBUppKf6C4R4aRxjLB1INNMIgGMTmPhzRbeyceJIQWFjrk1m7dOu4XBCkMw
HSz28SDKKpyyK/S0KMagUxxolX64oxQ1vxzJlVbsNmlG2blK+ms4j2zWBapaQ/cq
IvsDQVJxO6Cj1m92rBrSJJ0dTHJCS3y5GMnm+fOW1i/Em1+IaLzerblTZNqm1/t/
jxBZt5HvqkS3nKNEOP6G6vvJPXxfV3l6AKGZYOBs16BZQu5ijGb/8Sdvoaw2bUY6
M2EGgxauIUsbAWNshHLe9Psq3J/TIog/evPKhZYYkfDq2o/OV/6IA3NPPFToKLsG
qmnC//QHqz8QplKJhKsEQ47p4qld083WJh9JMk3TxCOOx1xYFRlJU1OIyiKw9sYX
+BQkY4GbE9ntUb+OPAhN2TzGfY+sHfCOZ+8u8DLl9nueJpIKkkW+2PLA9sjDu5vV
6h0kbrrQOHnXUagZzC94ZIYk5FcAb79zFi9G2JFWtQWQVse+C3l511rHr7litEYO
LybIw5vycoS8nryp8voIGjJh4yHl0J8SkbAkC7IvjcDwFuYwlz2eITz5ERHKs2N4
/hO6ETwGSfXs566ZGzlVxyx4i6dp90vLBB+tYBf6YQ7wyarYs8ZCpG1iOnbMmYo3
axulmogIUWuk0m3e9ULf92MnEtII49WhYiLuTFCfYw+hY++2wmA8xdOnOeyy5dWQ
z3oJK+Hr3zd5MPasgf8WXXWBFifqiqPPpGcaiXaAhtp4IrwV3ERW+RxAbMItKTaa
gwZf9N/LqoH2aTXjpWg8sBHQQISrm51hR2VzNO9t/krtgW8NcPItqajb2v0wmNHj
L66ZpZQmjMipunVeYNmDiNJTLQYLlcUD6NIOhAM2AXTm5JcGDijkyQYvl83uo7gP
AdH9WWGAL9rSgT+wS8h6F9+kVMkA9M9KbOsj7I8Y2MVkhvfnDOmfo76BL9fms+N1
yOEzaeR+8JhCAlzljge2oee4D3QkjylbxqmmPhUNxemTI3PpV5H1kCeb5dREWzcy
IhIYfZ+m4eNiAKmyc3zYamJ+pZ2MQ2mHXBDpNbr1vJVgPIyObvOE6HyQXBsd2HId
1QfOgQ/it2buq8Myrtzk8BXrF6+Qa+f0FeBT7bodIPRiWg9r+fvRmz7HVrfKwMfJ
t5P4s3TRaFZjS88hnOh1Eqkm2DMd6knS0MsfIqzG94Wn2BdrNp7drOkdjKrJ8zpi
IiXvq/fW1wVaAMS2hCrg8FI7IzF+IxrsvUdUSNlY0t0kjZmX3WBYlpGyBIJh88Ic
H8mNQAMjA2O9NYSOAKo0jDN0P4aVc5X5qF5qJC/RwGwt4yL7e1mCbda5L+5RvdBw
AnWFGfQbmKRREvJ0ympTrwcgkrOOSkj/8PxYwJZW9aSmGLa/+h7sHtNHcqLvrdfF
Gu5d2S4oidplhxFl4UmYKIn1dTpKaUiDmPeDkIB8U+uZngfx7jvOfKmVsfFMivJo
m3BWvBE87nwO8wcKyDZ6COzesmhjfGw0sMs/cMprr3psOru7ZeraNnDOcKAahT3F
+3Ov/qj+A6M+ypV5iS6ZnIhFDzz8LQ7SdSleq7fpWSmX/4zsCf9UlYhTGLVByuzA
rvPNSmUdlT6X3xZdlCwkhmVdlIv37zdmS8MDkCsRimUOgA3wkCKa1952K8bkar4w
i0KI1vhQ/M54b06BczOZ4rJFfOTogIh/ZjatRgGKBdjB362hNX0tjPB97Ie+B4ca
w77wluZCLd7axASvELBHeH6H5v0xv9U1Btmx0U3I/0EzVBJA3yRGQN8udBB2oY3O
l/P23erXzK2bD9ducm3yFbLHOevsFoahOaoXaZuRO2/O4zd6XZse55yZeEucWY3y
WdSEvMCJcZtbyDlAjIOaIPVnzJp17qTYEYfY0C4GLRZplkJIWLAFOFIwOg1NQ7c8
qFNhYduSAtGTIODWvHH2f4ZMKV6FYGiHLyX5QLo1j5K8soaZYiO7ykdSRUBF+X3b
aYunMojTCUx0/P7DizaA1pvOVz4MV6JJe5gi0kV7sz55Mk45RasNISriHxp2/Dx1
IIsYaiA8wLhGyr1RXMz98DN650wqYhRUvdTLbtFT275lsun0QnoCPo0oIBb/GJNd
t65unGU6/DJxnFBaPSybGV1VMY2J+VT9Vto+8ms/XJXWtPODhe6fIXJZYKz6vlHx
i7CoYTTx2f9PWwqNGs8bS3mFFGYhvdBNoT5p67X6BGCrFengS6KD4o3Bd7fkxtkw
PcIh362jibfsNgEl4b6Oqb/2pkjfdiNjeQtlsoVloTPydTY8xsb0ht8TZBTMmeg/
55e64AtwgTkaiKvmeTcXM+4wNc6eGY2LZ5UVz/CzOR3h6ceWDzJzlTtXnBib2R0U
gSdyv3wzy6ThizzSbrzw1tJ8pFEhoYpUX7cM9cEMymBgcSFd5o3I9B0LPlRzRZx0
9gRxIrXhHyZWQ5S3EttowuDX+rQZHI7ahRk+VJAjm54iXQ1aVTcsdVAfRspi9E0X
nNp+RoaMHb1CxKKVFbfP4RDPQu5jonZxbCHDiGqWqhfP4/P+pZdA/zjzJ7iR/V9a
B/5qMDNpi1Lucfj2IPgqlHYoR4wjF0p/iAgxniLq49OUdo0479iClRNQt/RUIrXP
IriN6VeoDr+iYk01h7wfqdmBSUPBnwQ388rNNMmEsoOxmbyKeQWC3n3v4RWbR5BC
ugWmPqsvbAEsAb2hofMAXeSKf4jywZJutv/tE1t2BNrMJCCW9xS2uB5aH1rY6DX4
ZNLNi6Oy4GQdIdXpcoGfvSH14Om1w4tFsum/g+cBaBK6UEvk6kSWnEQGSipw3sSE
cWLc0Xf4IWe+3ELFxN7YX/kUfHoFDzpwCE2uFcGLyOnUsUaJzfhC1kNYldGE1pEv
CV/Nks51GriOld9Gi0EI4UkXu4W6d+ZHZbKTBmJkD4y2VVJVkgX35n8v/OZN7DR5
6o3BGejTJrC117ANheIPsadSxPi7YTvJyk0tKt9SfRFrT0sIBeTV0BBAFitoowFH
4EsSBTV0mWbFIbvpZ6zVbSxrjUWI6NstX7Ey9MLPgEn6Ok2wfGMEcAombCngPsPL
9fhciQ/rmcPzdGWfp9l0+yGvTDom+/J7wsyrb/ETeBjT7OaPAvGnVY3z11sr8zZK
4qVh58ziGjisDeSo8LUtDwnPcwcabfTznd3fgOYmDFRGwMLO8AiXWKkB5FGwRM6W
TC/GeWZDlwcaVc8AP0S25wVxBt4mhQbrTBvM2UdD2rXbIzTT0uzNVYMeFrbqtunZ
n24i7g47fsar5McpDTZtYRjEejY1DeoGxjf7O8XVEANLKMspHxX+7F6vDm55rbOX
WvXHB46gyBa/4i/t8wZt97HD4zK+zze6k4pmtwHQpPIGcCqeWGtPqOUgiZZqgt6H
oXN+dQcv5ScfzH91XDF8C7O8CTiMF5mONrZXwn1aCVMuCWBUd243Oo51uUnjCsTb
4HrsfqMXgFkHGZDdcH1kLVHyo0JH30/H78h02c2QiaPYVYsRs27o/DQWxZG1YOeB
NRXcYnH8UBjuqjVnncXsyp5SDd000gc8gebLLqxTodbfJ5aSz7zDolyePUCmQlLT
ErGLHxlkvYL+MMiI5cj9rtQEronLKWdP/Qhwlc94+Z4+cp0+pQV/leCDcQ5DslRm
cEFyrFqzlegbNKsXUeWwPHWyp/qQV4r+2/YTHkwzvEI7u+lkiI/7MYfocrFn30pL
XvFRLzJPPknsNLhM2q5SbKIa/EeeOFOofEkeVs4t5TOtr+C9yCNGIPLjCbJ7xnui
r7WR21mjBStlNaBBNJk9XF3WrH6KdjPvhfF9dLXjXF9kecKBK8Nitagf1GlRT/iG
Hn9NUfL9+zaATEp/Dlyt262C2FBHCcey9W2HwffpgliF/LqMuQTSFgwB1/0o7PIt
3t1pbaiwczVLCU1Z1V6i61FDc03ULVfsuDbPdfA95abjl5oGLTpjA+OiW/IUtgNF
LDyX+3gJV1da0oB1GEfymCHQaCfO/jIR5sOgIC7Y4bk27c4KFvls/FjJX8YhaPfv
4lXGtcWbkA8oEFngjainok20UhdNzRrdb2yILhGtVvjg86MIxnl+ZsHo0wUfuxqr
IuoKUeu70KYPW+81hAMiG8LCX21k5htr8Hpg82Mz8rbB6qek9R5JQre+m9McuDLx
+/Lqev+EMdo4xLbHf3glcrBJhiauo5IIx/u8H3P++4+iJ7e/E1tC1rhWzYuXjI+2
jjCUfExtwInU87yJufvlFFaKsArbg8g3RNv3/NR2vF9HGEVVAry/UBokKeGMJDjA
k5O+y/fgUy/kdWoz2WfK/u0cCj/fhs7UEP8l4LN4IUga51BHU8tydiI9v5YRCj5B
RNWnfTee8J+S8QwoNvKgClEFIbG42SFsopCUwPkHwHT5ay6nnB0CArMPO+JQ4YRH
S7mXhLxqCeQV5yxevX6lwff3qX0lvqJ4eiFXb3F/93v20RM56GMPo3gZ1S2uVUui
XVfRqEMpIwUkkMK7hS95aaQAH5ushCtCV/OknS2Dx4ROJphzE3app+m671zJsxea
ey6cIGxvCw5GtFpXBJ19xCVn9quybQU2k5ZMbI7VEm8+eeo8wdUf+HeIn62f0pmZ
ZEASVCfgRAiDBC4O3czLLvGgjPYJRmtnVTAXDVHoiutkOCVifo01lzAqW2bbnOM3
2/Af66/CoJoJd1pN7vfptzX4ugVO/bEm+I/f3sFG8BmKfcfJuiaKc+SiFxpkrtav
zjymxpvTX3XVkr4IrDyuaLz3ozwmx0Av0XaHRfspo5xhTTK+0dFbzUrARewdHAgn
W1hVVvwbX1LgslDcakOE4uoSuXyXP9916Zs22Vawm3sIWu/jQAsQcJu0KthcdySj
qXPLO652lgUYCHkIsm+5MIMSMGPjS1vcqRw4GtdreVoCj7yxw/XizwurkNbRO2WE
u1oZNgo7l9Jqx8vRBCrhn2TvpKIpNlY+LNgAUn3QVOv9YEq1Iffg/bUwli4nNNTd
ZbZVUqMWHiSHBI5LRBmiyqRNNtGgjnC6YG/byMXDPpR1J6t81FlbpBxl96a2UzuG
5DZFVaiJ7H4U2xRfluhWOC1vQhVq6bsJM49MzFbOh4qu+sVKiirt6AdQ0I9WkVj8
1KjABBYszsrK3BA3MHpZSNGbFQmcqNq42ZlzN2fzvX1VtHrc2gIGmvWozezggh0f
D3EYGDNrRcYKQ28T+Op1rqowi/kmnaGCx4+J2z4SrB8LeP1hRnvUTTR/toJByAkL
iGdo29uPxWs/k1TbR0fCtavSggBbmTf9ypopJrUMPQuLmjzNs/R+oBkyrSu8YYjv
ajjHZzT4l7ByH8kFQz/9e+3ixF0YCOzQRjVH5PtJnRhz//aXe0JgQVWyAl65dlee
duQsO1xxhbS086qMBCC2jJA0NWBpgHbu58++8rPhRynKOvdTrKHB3JtrvoFjLljz
sZxacYnKRceUv/qzJZGsZoIW2MMBSuezXgb03ajv22gBqPrQ56r0yaxDw0lrl9nE
C61er65jfk/jC/Ju3KG110e/AVOpHGDXRTcJQOMX1u1xumbt+Wk0OlM/gaH2NgUw
JpZ+a3CoZZkxEznJhlMXmqn56XjpkOB060ePI5yTWp/4HwI5al6M6V2EMWpOunzr
W0aJbf9O4oXTlGH52qiLvmSUf9iCTE/+l6hlWqjZM8SCylUIsuwlYC39rTlNwOjo
eZGiV4np7BCuWzTJDwblnIU2gjmtbUJiYbtMcCherc7tHpSlWU+M4PB/ywA9n1mg
pri9BcmHd1yIYVKipoCGO1R8iiPmgxPoLhdK6sKW7OCa0aGKYtYkvxRfBI2T5q9l
jrk/fShUNUKavOQUCV6OTon9IHuv8nRONXzyE42B9GTwlkCJ4A9BS6n+PpGLMqhB
mWTS1+8GasWvpCuc9pwx3/IQa6nuUxlcbjBn9aXB+dB+B4PKmPi1EMHehlu2by3Q
WdalZs4IrMeddlpjVTLXJ+ZUQJqE9PJ69rWU/7GCW5TD7i9ibp3DoD5PVYgZdHYZ
82ULUdbUpHVv2MoTozZYhgTjA0gw4kDPf6/GeRdD7jOsPhoZqxYTXda6YFLiouf8
ThPxI1k0kqrj6KyI0hyfdocr1bfWQdFpzJFxy9bOm//qqTfq7j5PxPoRdI03Judo
PerTPxvPxpJK1Oi0wXq/w7n/aDi5kwG0hCdbf8tG6zKQVOTAFyjtt1ruYlQ4tU5T
5cp3Pcyqgn+VsfNQnBHNv0C32OkiWk9BzK2fvWMrtyV4cRloCG5MDhdmGEpJ5jrq
USw7U8WrnR+QVAIDmK6GnfjPlTksIwBnkzkhrjEfTwoiVxSJ9EB/ZgCWKLpRVTVH
Rc2vC37IHJjnQM5q0dsQ/eLtD6ZaU6oMYMi2B212CKiiNxeziC/6uMtImy5qS4+m
Qh66HHq8r3dhRSnYrS6edmTiCIdDUhY67600I+HeVyUiMi0YqbCUulpN169/IRNY
TdEubibNgxA5FObKV+rMNedRe4m2CiGUTkbbNnDLPBeSjmqJPY+Z8k7Vl14Nqh4O
Eqkwnz4GdXxW0Tfg4+VO7JaWbZ9t4+FL+KLGdKpohW0wAssTmujcZXSRKYBQNpWo
Te6DlG1OZ3DHWW5BIndlzlGBrEq9ZG8L8CRo6etZHg/hop8QOGaHMAejgN/HXPuL
7RnHU7XfcAGVRXYvndvpdYaybfmj6AuEb+GLopbfS6XjypBdax3RgxI7rK6g+syf
Xcxc1kjKZx4Zzn+fRjjPL37Il1vYYF693mRy9f5CMpzv9IQ76ZWUwBr/xdNE1w2H
T+Ol/9Y+c9u40QfZzDQv1F5Gg7p3umeAG11SVd2Wv4Q3sBnk8Xqv+jRWYQD/bneO
0Ne7NB8NuLX5UQgcOKCa+5MFAPZSAQ/AFE/Ppy+YQeUr8Xh6Ri42jjZ7LrE8Zc5Q
iChVMn6+Mhbe/jlHAYLi51KI0K1CcRQne7pbB6zbDh4tkroUzrMHE0t9pXoEacAN
tJuzaspZkr0zNibrnJhdT7icdePj3reGIXnR7n6jNRgcVpAi2mhaMXU3E+q5y7XF
qLVergxbEoSTBarlKUDbpQCwtMTmzKnWvQ/f1uFWLomevmT9SzRlY2ryVxL5xe3t
rNriBt2lO6ABVQCsPGhVrNiZA05lbDmpv1T+2XOU6oZUXBmb45myzNJH4zCzbIWC
ijL6aAMZDrXORQzQC2XOz6DIAPIhTNt4Pfpqk2IN5JNEGbg9+aHqffANTfNDwDg2
gHy5FWlINzR0gvfJX50uV8AQuY7vcJdz/EP+E9mLwMVrHKvl/Gjp3kRJPqDAGp01
tMD+XXXYar5Mj3/LbU7B5uEwupidX8tUuvaXGboeo/eH47G0/0NuEhI5/8ldfWTa
pzTU1/C9S+NTW7JulETsdtYg6XdSYpY8TlsADnsofL5QcITY7977NYFvu8JztICd
9KvmzWV61ZpoN/vqdFg2OoCmD6T5xKLEl6j7pPCnNransZ4NvuUBio1J6xCWUtYN
LgCxpGlzf+jMOtwfQ2+siEmAXyiFwGXXHDB37sDoxtjo5oyJJ752FcVf8/mEhQhF
D9AFjWbDYGY9FF97gBAfR1+oKaXxliKDZRXrM9OeTEKRjWDOzY3C+v+ddQrWj46d
qixHtWwgM2C+Cmt4YswdLUfpgiEJh7fZ/qLjEeqvjIOo6WKcRwqFUz64iVsbCBIq
Mbo4k5h2yd1DZhU0jv05MIZP1RAymtwOkcPgbNpnO0SzRXJuB03HfaLGIUoUbfVA
8Wd2pRfnHzrfe++ROT6GWKLg0eVurzcntNxjW10WsduuT0iJwUwANCIdc9ustTvE
p+sDfCQOpZYaNxYv76yUxld6bh29tzSMr9+1ld53XE/0UXu6OgGQ5YIcEvuuFAC7
5xstaoqIRqhSMbzyvX4PUpm0rpPAGrrk3zrpSQlwEW/jGGqCJ2cxr4Ca+7z5LIHF
xl6TTFwIFwCkmiytXTJaOe7f68oPJSwnVuthEfVrpbjNKr+Li6lwbJ+yEJHWxe/7
AXABU7fxh1UtJi1jrV+Qft1XZryH/mK/aBc5aQzSTVTRuKS/Ts3UHCfo6xQudpF/
wNwyPrkwe9VmX18dQDVYaI0aFg6OZfc4SMeUCHErwDX1Bq9lypP8aI+DMlBtmD3a
+b2M3mT3xDQ4uNpuTSmzHyQlq+mxO+ILXjQOV2l6If4CPg2wchK2oyeyh9nGlA28
NmMGSAviU4Tl5MTsOTkvK8+okroHyC/I1yRHIv0VSKhRz7LAIi2w7QIV1lFdHpE9
g6gbxWci5079Df//JAcHD3/Mwl9pdB2nV4tLMTn+T8q9jyEuHKii0FaRoihwpXhq
87dAB5OiVoqSXNmkprcXQuKons9k+DxRlyaLIV49ybNGuyg8UX39Eqpv5Kr+X3w2
wnZzatjFGJVDybsB+TiSeFgQTyR7WdXG1hk/Q5nk9ZRfOQuM0LJdbhr0r1ApPfwz
7S3ShpRm657jQCwPaMISKtbwOEKDKJugMXL3YrZDRaOEusWsjFWUSAgWB6J/dVAw
wRt5eVgop99a2RzzkZ9gjeDvDgR+WmgN4g0nPRuMod1KaYud/HCQzoQzJvGZvjrf
c0uh+56C6bI0x32Em97LVuhhmdcGmfHvfojgNgrJWcTcY1OWi7SCKx4ehlfBAAxJ
rwcU46ByCFPCa82DA8hvh0lEHT6sx/4zmP5kN5nKLw9zAjDQJsTBYK8HmNLR3GRV
mpRIWmveA1QhTECVHBxbbLGSioEYNRRpsTvzMuLopUTWdhWSYPfPMTozO0nLi1BG
uwM1h7q7/WLes9pCzDXZ+S6fPVxnKvjXJq9YsXDHITqjQYT7UP2ImlW+yL23I4Sg
dftMthSCtIeptfkiUFvv34fTRZgTFgLKoD6pnIERL3okdCWpW5RVoOCrHfrd75s0
7Dn1e7D7TKCyNlsxR4U5KkDliMmf77UrEfVQ6K1JR4ty69QRlDuatsBflpDU5DOx
HAixRT9CtqeE8wIpQCz/spTdZ/MTD40xScXYlw39gYxHmkzdbuC8csK1dGOYFD2k
UynMk+/hmuaJ0BgkLUjzdiA6P7GQFwNk3W0XYMNNPkxifuthglN4A4nrtUMcJ414
MA/HBNSYb366V5YIJogzQI0xvcZjAMloXIgLl2eST2b3tkVNw7Pw7k/sH3QoLeDY
ykGVpnhnj+AUxz9It2Zl2NsQq7ve35qVVltqfYPgPuvRYt89GKcT1zvi9h9I3WSh
DGHCt1KssRyrI0PNaqEQXp+7Ie7ZLYLJpRPKxcK12no3I0CO2+HJ55bIih0uEbI9
HK0jIKu1/bb/R3nQU5iHOY88bViPsjgS3OKEdJzoTiKwQB/96Pc6XBYJpgM1NsJo
fq/2IyZALcXoZrCu24wx4v3TDhgAtW2KGE+dwgkCZTnj5GNcCTnNqEDgQBAOzcZ9
ZG2o+n8/a2ZNpn036RqjbCGl2644o/VDFuaoIQC3YXGz03PfEHtKPeItQufIaxom
5NBeOB9y5IgM07iAroUjgQIrXFhRTjTXdnPLMuh9LQDVdSTWnMVqbMCFA+/M1gyC
qeaj9w8w/UeUNOHOpSEXvYA6XYi09PCRxEAdtqK3XuS+DpSplUkM2hDGU0EaX/fd
m+2rAxbrlJyy6HAaP2U03AYgAa7PWE0eSyN02rSpsf6XYpY6dnd+mg8Chrz2ulE8
FBntKiXQ3UqCwIqIIKucZKIeRnJ75C86iw3T7Bi+VLf58gy2k4Ef4fcCDB4ox13+
rxCJbu3hTunFmlHnWrmrKUVxlXvvvdEwW6XxG0cyDYlfj6gjINvfJVmXixkGWUyt
AZSD+owdgjSaT63s263q8A0NWQoNFG/DhkXvqwD1KdqhJykmh8txLrQm1P2lNU8+
0VoM9UxlTkUH0Y5RBPROF2mkY2eIBxWo4n7es2BD8ZkJ+mxVR8495PQqoorQhryK
Md8oI/Dh6yLAqn78GX/r5kDzntxP+ueE/HYdUegLvF80162pG4l/eyFgJ9PuEt1O
TCNdf0chNPgEL01oaeY7wnxVXruwera24C7MxyUyLqj5JBb0jZiAMmWv8dF5ryDv
K6/Sy2SFN43utXsMgDxpcuo8nK4aVK/+H3kv1yyj0wSmSL8FJv5NKCw+E21dS6E/
KI5UlO4ntSj58Xk5kMmk+60oqsW9Ay2aliEVcop4zu2u2MKynH6YZr/sN0CYnKCb
DPpUzxlhEkxmonJPJGaxz5DTEKZ1WwUDtEMiMGcEbye7/Lo53GJ12Ib3ZONS5jNm
mzjs1hwCiDG8XrcEeSQMaEIHryN+tGD8FRqM+IEMzr2ozOEI4BDE1X7crn9M2E2F
7JPT66LmVB6i58ExITN2psfm6bdx2m+E35ZfDarzubGRrm62tQhP8hdueiyvT3cr
fCzsRAVd9zPGo9I0Wk86J3Jl8K4ForgkTh9jJsv9wQhRMAV/4e7kGRdDkeagmPdy
r5wx0oWQtfGhwRx20j9Rh0tDcUzu4yZzSZ1riqtbpytkbxUWmGtZ5HSv3rMOMI5P
V3VD1Vj2PZo42cCpjTXj2txsuxZt9GimbzR5cTroUiCx1HigJfUO0dIiBcs6dI+C
zjMKnmACYqGGBFTgvgJLaa/4ET2ZsZdE8KemTAtbVtB62+l2n7YP2Ezv4daHcnjB
aWCwtzbnqT56QI0+4rWkyp1CKU43B/VgxOYOU9e1g5ssqLnzUartQX8xWGkSuPuE
kCETtPMRf/LAsFbA93c8h2+zktb9DLB1jyieem3XAgD9t/znW4H41OXRxaBEkU4+
SHRDyp1HIuQMQ0BwyXYFH8jI8SYbeAgCdXbjTPUiVylO6H2LE12HxmLeX3SZcTkU
YpiUBxl+UC2jbTp5bcqxNAiJduWS+ZRKBuAMaFazxEX6BMLuiANOwZokmE4ZZ/xF
rz+OkGWV9CBymzSOrvzgsIKYakBKyGuG3ztovsHSiT7r54lX7PWUi9XWqqL63as/
0ctKCgAHaqPFRbMpzrHSIp+7B6XB1rhFXrkG8NrL18ICqr3F6J3pdfOHTVhtatCX
u4ZrAYU36jsfZR5CGfm2MguLoyizCfY8DOvPXcc5f94dcdj/Z+489VYOU9mBjZcD
JQd2KmeuepUhdINi50LTWkXt/GyjwnfcOsPOutImrVi/XaGWtB2SoiYhbBVrgpst
I5GlppFOHt7tQKoeKAArMZ6Wu4VOSexcPr8pKoqF/CjsHUGY6TRj4MXaBObcOjS2
Nlut8+JvFV5JboJ1XYmtihJHEA7Mwjh96eDMCwm41BubLipoxylpWxewgGAzffsE
XHTK3hMFxlxf9jF36VDnc0fpODJEiiZxggj31qAlrLi0TRhcVvXk0TrSqIXl64CB
DbVL52i3Yqo1YX7ismQF5THlsnbDdD+3pSCuB0bQABWJ42Nr4xjYoIKeqepRo0gZ
SoJmfl3A86LB6JDEx06K4JgSNPEjbsaAwHxClHW0wMsymh18DXamJQSzap5rSzFU
dNdecJH5BCaWPYgARTBXKwj+8g0Nb6qs7aRNkjht9Zrp9dB2QQjSZcvPN8MVjs7m
qAXf39WlU5geHWKboeP6Qm0zsuxoIcVTnHutiXngRf0rC4fsdrMjDfMxlu3pCiOv
YlCy0tl/TYMLJ+pXSvsYoM2FbpgOElELVBfpBO82fPi89qMfDFSAACvRTIOIn2on
eF0cpvK2tevtRykXssBCFEN7N2yda3ar3TIZ8fgZ/+w4wKF3ecKB1B5o068VRrMQ
b/lC/Bvn2451YXIdqCN0iO1VRr/tWajfzfR2lgN+0EVAUOEyQ/F6kUnwiSl2hIUF
uY9oYcU/S6Fa41feos8FE4f+DspA/Ry6xxJvAG1AkVp7zYkaPTRRzL3e96T4C23j
iEhwmgyflnSWjFfXnJXqDydHab2rCG8nccQydhwFJgdmGMkn2LLoAAZh83E8mkWE
l66gGKOuTjOn6zvHeUUWBpRLxwN8H6MJ8wi0bcvL6StVXg5HSf8lQcn4JFfhjSJK
OlEHpGzX0u+tUNcEvnzTsXE9bpVeNFndLsnB83jTTBj5aQqfWqQ9+DNeDWeHsOt3
6WozuKnJ+aDv/IKwyyZ7Yd8GstIl3iSmuvhQBY0YjdriF6Mc0wWuvYgzYA3CW9Kt
Em9lDsLBjK3b+SVpEXKU3fmzv+3TL7d7MaAwEj8Jf1p5Sk5U5LsW8L7OS5NdZVZg
ygg4dr9i3cyWlzGD1JRKisenn0BKwBmmbxMXuze1LytFbzj7gEzsFBmdjLavWnQ1
5/3La4COsubQAccxwOFDdIcNPqmZ/wl2g0qh0SBbEGHpjIsrUlFG72XlNkhBRXIG
8XUMBRxBT6TrahSeANhhVW/mMy/E/9uZDryRKMOHNzo+oqQ1oOcQlX2g/TFYGdLI
EcXL5JwK04/744YswVIV4xHf3PnF5jGSyvnIcisI7j+Aznku+L7Z/o0p1XAwE8Op
tfR39yUba0VLV6XkDCakNk+0+d+gAH3S8ZdJVoNvnHk3XZWVWGzRyQswiG54baGG
I6W+yTeM7Mvtgw3Hj2q7788tWBghT7/tNZs8DufjOkEcVZAVWHDsexh+ISmAXgvl
8BB5P3zYhOVoX/1Z8ibwth7KSHkaJYP1XtXE30tnLZsvO6AI1GSB97zRfOqEKf0P
7WuqSVhUuW+Qc2DBht9tl6l2VEt0Xts+LCDIsUDaXLb7oxDb4sYvSVgIxk62YB/Q
S0Y9wgxJsrxiv5i5JuqGoohUxUgfnfnLe0Eh9C7HOKihUrz9Gi0Ki1/PDOqAtcdY
wkWYYChmq4sa3lTRnUbZ1V2uuJ00N1uDMI3nwcmo47B93i6BPEKvaJRnOoKSY1sm
gvtGUMwuvwzeszG8LCpBo02ecFAyKD/T0aH71wMs5rH7VAy0DDNxezWO8YRsQDgO
6w76sFP0R6cvV7Zh6SDy9G4omtMmVu0spcTSe6hEvmrfny4AOrqVArEQjDc0m/Wf
gI+asbzpuaUGSh/Y6eXBKK/DK/UuULmhIObNsAaA+0NnXRhNClhyVwr5KGhR2WkR
Ou2LnZPnuH4EiLODyqtaeQsQvc6b9eJlACGvDeHKzVMzvT9GDEYMxp/NY7zD8TFb
qC8/FzO0f2mXWFPli4wjAtzGGAstPO0Jt3GqlYAKScjboytBQT52RZRPhO80w4eK
Za19laEupI1NhSmhhpuh8LhySfWNPj9pJyzDMVjHXK2JM6k4lgUd5c0Dax/Aeq3O
JC3bENLXh4P8US8kRTh8ioX0hETff1XFRfES+2fSoQ1Uq+9GTqW0S5aLN8QTB7Lu
nkhk3mOkgQob56oqXItgU+0nG3MaqQWKztVaID3iE/ZJwMhu6LCZjZbST0QgFkc1
KXiGAJutcjahxNhj5cBrJuhR1uZmUXSeicrrYp5vEaF4/WPBwq8HOs223XVsdgs1
1Gox9NRaMgt4SaR/zHq9SteWHgDQkW/+ogffoAEqHerQm8eS3SgrV04Fm2aWFldo
Rwg/WEptRzoNkGg40Dh5RJ3NGMY3HTnuOqth2oEbzNh5HnQ6zLxMAODk/Pe05ARM
wCAOHkO/QwBHtVBzZq9dC7knEqAXQNjC2AoKLy+W6uq89dfRfyzh3Mz3XprZZCid
x4dWSlC/UyxmI4VeZjilOO6XP0kIbcJ4UIS6JPwKoFSYWpCP6uoQE/sTVdFXkNVV
+VWdTpMkGN7Z6DDynjh1BSzR6Zy2sMTvcurP8kpdPxoWXtawraoeeA4ikolHAf3S
WmciTKaA9ZV8P+6+0qDPyOPO0TDXWW396I7tnrRn37LzzcIg+n5ZGZ7QuYYJ0e9I
tYUQQMUlXh6O8Uw+7nxW4kZQoBJ8l6rXT9KSjAiU2Rp5z8GVGapjdHr9VpNv6L+u
BpzAyKtECg4uCK01GCVRoWihmxiYYnE9nLZLmy5eUZ1Dqhu8EzDnawxPJ9TOQymX
50xpU5KUw3mCz0gBnVUxf0w882IEiiSmNX8vek92XvX+MsCAeiTHbH6jh0yPmvC6
ZdYwk9qo/NGrIibRtKgbhX8vdW/tS8+0IiC3k+1c/DfDLlY57B4PtFVHgA/1Dv7B
Q039lHM5J3rzCDcYyuieS/prcC5yX5MrLtEiVWv6woTqpr0bXt3AE8ma10wQiryi
8IGHjBmDFKEAN47JGC6Z01T/e1QPpscdx9YFbTREqkPxqpCyLBA7zAJZ1LgMCreU
uoKG7lnzdrlEhN3T0IriL/6sIER8JUA51Lz3IA0hHZe42us0sdKWvBMGcH3d3c1p
xQCa/YOlPOR7355Ps1ucmz+htpKSn3G9d9Q/Egswt+y9/8V9NjXZjjjo7SFkLC8e
zUm+dxEH+z8BSGkxEziYehI9y4VoS51M4Fd+nvPzAqS4MreHyw8efu/asrdEN1A/
QsTK1pIT/GSXlF3MpvJAuvL7QkHX9Dc0KbSt7qDZyAFp2eTKIRGIhAkLk0Baiul8
gvaUHrOO1ge4FIOTuQG7sxcXszTaUemrvTuaRqBMwdGq2e79kXLfHvfRNMAEas52
V4uoDVy/A7/yyo6p3pMNl4H9vRW7t59E+2yWW09qgSygCY7l5L6l+2ru8Y1IroP/
SqIrtOYuVWnYRDDcKVf/K71nfHlncYwTPhDh6PVENRP/Ssii2eWjDAfU8f2c6uHc
FCISSnl+qCIbJ7o+tsPkKkqQC6+ckkp1I2LiG8AnpnkP/Q1x8TelwXSjT9XdWaqD
tI0PaBKloZAI5tW7w09A592x7zO6qLtVBi6vqrgDfV9DqLuzEUdwskbsmdrn8fnV
dLoZDeVHLo6YZVY3l6dAml8M3urcY7i0jwJnQVpW3rwfVL2JX9OH5B/fH/Bycz61
xvh09SVkwFxaGFOiliyDTa1B+crJNExx07FJ6JrpIqx0JAaFfFFEZkfD16vWElTl
7Mc9cM9Y58yfF8nnSu1nTi2cf0I2btO+VAxz8JWQBOnF709sBzla7FDYu289Bh6F
EN3151loB6cF2qp0EsZmd0i+0RYDYzVKuuGH0ZmZ7jycEcKabT/lYc58hMY2JMeb
AhRBBH5uRCC0RZ76U9dhWaWRo45oUPdc83z5EmAlXkhuATXwFOnMmbi78vYQil2t
OL06mRmGbZVxVyrqicZmxwT/iI3Q0o30R0vQZpLkoUCBjvhmKyDNwyDFa5lD6f7y
x+60tJnvq96yZLIEGi3P8xZkpF94WR3u9pY7FV/kidFHcpAQkxMWIU6kYrFj21kA
kSGqHWXH012Tz9bDGAm3LxKqdcDrLooI6wlaSGCXdbeI/073Cc/J4wYIjU6vLcp/
LExJcf1qbmFe9RQ0Du6V3yucFipiIlp1THZY78o/4FbWrlrOJ/ZN8uIeV47mXIXS
LkbGtFBE3pYaiVPpg3tteF6uIv4uwswib/Siqxtp7F7JGdbGyq+qG2HX4gtGX8k4
ozz45aIh5v0N3KqofTWj91qMaGx4fXH8z7Zd0E8m+LC2YX3rwVjsA00n3p7kGlk1
Y3ADgL75aU+sw7lHdc+OHf1ArGTe0Bu4cSWuvo+dhjAR1j+r9bHMOC2dque1wsCf
Y1EGe23SZOqM6tRb/IrjATusuTOMhq57Xyvb34zBW7SNs1C6Fw3K6dfZu6pTCKoW
TX1KN9PGW9YLEXJ9+4tBmhyiuZM0ZROiP4KIkSfaxg10rcodNMbuAUqc259KIXsd
KEVhMOkDF8FwlAk4j28wotMINrTrHOhq/LqpkDsSY+7le/FgsSOyupNoYnEs+2eE
Nv2RkIIPHLpG1RijxfncK89IaVSNx7l715dxRgDo/RPimW69743gcoE2u0JoT6XE
h9w4wF6yqTTL5Dfi7Fz9Ac1Q0hlT5haAXjCb0U6ShsPKD4gYIaL+umASNDZMgG61
4hdskWXkOD6y6UZwS136samsyQ5A1UgPAaNJO10JDeBK5jdsiBV+85pQ93uVXtA2
DfuqJ2ePxZlB1QAFWXbsxPtZ9Mq81AZU/zzeQJ3OTX86l4mpTr1kvk3y23eFNamU
j4jaPFzhyJSpCW4WyOlWuZ3TUAUha6vuMr/EAvEsss68EnArP6IC4j5n2Aatq9Yn
f9IqxK8Xg1gFFOR8nWiparwPM+KcGpoVR6p0BqKQGLUugZu+wZSMLKkOuCs2HDwq
8qQgJyop9g4PO5KkJCSpoO09aFTqA/58h4runDxlHy883eQmqqV4hY5w6VGDlX/U
oh10FFVjBUAprqRjj5kH1B4V7QQBhxozKwr6ht34shlED03c1PIwo8Dhj8Ov0Zre
OlTG7XGmMUHOfLv0KZlTD1EXXRgMMr3X59BwLIyHebA0txc78lX2nWK92nIHMLYE
2u83xYuB9GHzRDRhFUiV9OoL1j0xXkKDD0I8auvDIOZa8IdrXGN39m1Rt704cJch
/9LJdEwBVGGOMhzpT/TBrORk+pG+YeL3EYs9pRasd32gKTGRKGKjkvVN3+TfvCf9
dQGB+gr4orc0ZRySrQdC/kp108vvh2XHpZcBXoYn16AJonAfYTXtG3eASLUcv32q
7YshF7JPaKSaJNNyIAuXKH/vSx3MdS8MOocUDV8uEm5tVT1SRcJQDJHTiSmTT+f5
QEz6gj+V7QLbe5GPqnxH4BXs362G7rovUONs7OhAQBnGjvuEvz9sSWPdh8UQeyh1
3wxtV98BmZlM1ky1n1o64Uesj0ilLB5IYVzzK69BGeHbVNfn3CbAizZyoOx39pbl
XTI82BNRxqxUybKNYQCf4VRzL8BFqGTUWpmBOI64q8vhBed9HdXJJxSqkQrbEqme
6IfxraaBTCBFMbAjLlDTaYmv1C031K5WbNlEWxrL67kg2tqPocblxlmy6N8k+EvK
w2jt7sXPwz3t179wta+Nt/hfF326qa2mq1KpnKPY4OGTpOeT2aHr/+DeJu8yb/JQ
Y6mUqyqJ3OgQwMLroPkreiFiN5tEgsAFk/3rVP2rofYT3FD5uBovqt21bMbWf6Lb
xA09Bf0FaamUZ6AZ1ZQTxZGxq+Gq4cKuihmKfGPrTaTm5bL/A/69OvCQilzLtUnf
FYvVMCI425UXSKQ1hU9RopEGvCwdPcmfpRhvqlXWa8xnkj+8m8mnDl+epxCue42m
GZvD4G9pW3ho0tuIcswEl+UbbvOUbiwuU6V0nrR4VgtNMcqLIPIW88euHIrjdmW2
pEJZ7Z+2Pl0ZwjMVyCQxTdCa9349YNWSAWorLP50c5GmwD7NkaS0njsGUygiAxIW
ZoKv7+d8DXSFkoz3pRjfUpNgGX68L9Ohtb5XlxAVwstxtUhObflDehtu4OF0gD+j
LuddRmRqHRPZ83/tr+3/LFIoVSWLAY1GnkXoHNulcCJsi67yVEtzm8FrQWl5GH5G
VKzn/UhCmqLpy632Op3soMWQT80UQoRxAbGoNwrznMwfljU5ScJElgxGjh8Bp74p
NhTjRaQ4A5rG6qIdyKPBzLQH234O4rWu5+uz41OYyPMvsndHnMYppeX/j0C+BypI
VY1z3ztFoI93ttDdg7knU/WNtQhWT387mVTxHxhzBRztecE7Vc2JcEdSu+JxCuSC
J7vKkoJvEP6QBF/J9i3bBgqyrJAjrZdJXtd8SqG/Hbr11Y+VmtMgBY6mFvCEw+HB
gGkGyKR1uWDD9YUKlKTczQPo4Yf3GrSg4+vhIr2EkZg4GX3P67R6muZUQ/pP/dFv
V9p5bSegKq3KMkaaSpaL4tqEQ3gz2VfXd9+M3ZAiI0sDUq2ufFwQzCCZDq6ObfOR
tc770TA6EsMhe5xnmiqv5ejjm/iHv3m7uiV5sHMHYuIvxV3mrRS9ApRyBBZN5Zb3
jDfGJr98f4JhvkHP3R8W91t5YocYl+a0cf6bIJl+dlmoeK+69kppNwCLJr85YomY
/B5kQkKl6owMrojFIjkOMOGDPLzEwAuuhYQgihmCXnMSKguLWoF/vQxGAMorsAoL
a0rfWAmFg/sM9VBh84uhNwxhV+ELtpDP0tZGBidB/okDgltyC3te3iiUqVsyM0B0
diLlWOdXaanAkcFh73ROFd7aUqpRpCmvKFPSP5dsK7f5AnHRc+qM5i8UB+vYXi+r
KDfISj69n3NXKa5RHkUALB/wVNp4HUZudJb+io3WpzdP6fBzCYOJn9s4ma1/Vw6A
On6VlxXQvPJ/IGG0DY9RyWL5eYBF/aL1s/l8y3/TSxv/CLUQECKHiET+HCnvL9I6
/etJwa71DspyNFHNt9jpNlc9cS594f7koh28xwR9GziUAHf/L1QhoIQ1tILVhjl9
eq7C0G5R6/j6lrhKfc/8vouf87oawjVtgSFki8q34XS3luwIx4MFQVN4jKWBuNfk
XTWEc0PoQldqu+6ULKO/Ul2ujdMYaq0njRZFE2V9TMuVr72t4QKH/EhG3TeM1jvB
izZKhfchjsVkaqWzJWvbZ4Fgi6rGvGvwTsnF6d7PmSCN5Ukq8s43aNCaoxESPOZg
5KwkaQRjvsPwSxccaDgXqtl78/tfMIIo2sWhJODBSMWzUrQGMj7KwywiwRaXosVc
6zr4ZVVm1MLcgzn2jVNnIXsftZd1deqonotyyR7mnEwgEq2KVLDmv3T4ZCsRWgLs
eL+ikxPm2OraxCWSeJdZjT28wzltV/rTESBFiB0CtyMF+hnlWN8gCE2MvdqZW8f6
A1B1k/cLdhZghBh9KwXau3VQSIy0CQi3b5Si7m+uq/pqvtZLNyitRaAPkgsNrnWv
HbRow/2BKTr8c/AsPDtWs9CFdr313gboskd9Tsgwrj72vom0aDfKZ9m+ymtzY73a
6D28rPio9T7aO6Qw2K21XT+ViekY9N3YbyhbKxbm7mCu8nubbr6USGEF9sTvb511
BVsFYWXRH2URCLAwwtD9oNyHOQ2SgiVozf8yup3jgwfztLPNN6SNtXqIsAui+ZYw
RNuxgn68knr5BHzSaQgpcuYRvuOg1oypfW81evHqopQ/joX4vr5OeFZDz/cUy2W5
IFninjDhUvM3xgNsr5ond7x+Ct+n1+/00J4PDJ2LxxzFFWNCJxaGpjquqqLS81wL
YR6nQUTbVrWVvwuX3m48mbnqcx0AfwjIHEpOL+fuC+Ga4WBLj1BncTm7g3wB/UiM
FR2RPiPQa7bj9m6kNKxRnrcH7XjFh3+vplBmED31uvcrDBsDMyHZ+jFo94frpjMo
aufe2mzg9ViUrmeTRltvqH2XDFoOYt+JaYUgpuFowqTeLAQOkqHnIKxQh9wftbBq
Inh5C5Y5ePLr635taBZA/cXhMz7MAiklzAqLmfShRE0Wgv2izjtQa/M+x1bsSAny
dWRMCJ7bhl90vrO3sHbp+7X/uLjR88xNOK8h5BOZm5M5EHHeqYY5ohkR1ipkRxqD
CEnDnwkykumZs+0UZDfyLQzsnfJMCeb/XqCX022TCkNPyVL7LZ9YFc6ABx8kdT0x
5md0fwI/+idWAIfHnVa0p9A0Kd4cGycoN1VbcD0gVdNp4G7/XUklEQk5DzyacaAV
D8LRlntUJC2Je2mV8O7bfRGeLQ/XxMV7+WSMW4rG8FzCUFhcMHMwcOApcU/j7mfq
DfUz2H9ETyhdoQhhjsoRW7nEKtHNgVcS9+O8w7d7Ghei64cnZGcHibaPoKLT4IMV
Cbz4CNOwy3ZjpG0wMvjM04mnWoPu6dfXWo45Uo5X28ddw36vE4hGRDpft+jw8ad1
YijGhyIwd1rbLQ8k4jctZ4G3tqPo0hUoFK++BJUSHoGNsOP9Hwv1tmUASQ8oiujF
JMBYWxRgSNuiHOm8mw8zj2z5FtlPja4S53qph0LNiCQPJK7xjcTPNTwhCckT7V5j
x769h6rWQMStfCnplF2utyipoVX7pB2gn4kyle4ByHILJ6v3U8ASRTFqEC1oBAsS
6ik4ipJyTTOQMNnJBU4Kuzrb4HHDiE/Y3AsFIjeHr9+y5BVrqJWMGW8cfOFK+qsL
69/yHfwPVPaG8Jj8+spTis/OR08p/8cNDenH2HEh3Dy8XtLhMXCsokdR7FHO/GL/
V9KD3NT4FpRyyXA3UNzO29oI1+VuX/otSm14+Cvy0781meWOgsrZ+g6HEUkRU7RC
q2UvScUTs/2cHL9GDp1ZriM7HBG5233KSa0TfEL2Lwg7Gn0owTiYqFMmNf9pklMW
Egoo2pm2DdsCr08m/g3h5QfEsn30Oosu1DY/PZuKBLDYFN+D7h8AVSR16I3IEKeP
9W2AD2K8y3VVCdpOM2DMCR74gPea18cWnOUs+SS88xCB93Du1GvnEevQvfwjH2wN
Ey4FVJUP8Hl94OZ5qRgSsAogCq7ke4x9xDVSk8ep4T0NF8u82EePm7lLapg2Yp5s
EaFTLaRInuzq1d88fRuBD1cGF/1yu4lftjSNsHM0O3JelDhOJzHZEDR+B0NtnXig
WZZZaIi4nr4JVvwlIBQzZaraGib3H0+/Z4RI5YPRi0P8y2/jmqb43342fK1dt85c
/qrqFZ+Mdfn9XpJUpwjmyxUrEUeqcXHX96p/3dzwl24IgjQJKGiU4px9jkK4ht+n
MqLs6SdAfx8x/gXZOAWygN3O/0XugKsVGzoODGZRW4C0bWGYcaL1ISm57/mYA0zW
+1gEzUPXS4Wn5awhramH67UAHMcRHuIvaM8IWlAqYCQH3MySklnpB7RZyfJlOm+D
5Dfci5WDVx3UhxcQjtTDWSlD2ezgk7Ip+9NnX/s7geuXUb9p1mAr8OzGkE1EFbFR
hFmY9cUNiY8I2LsIcATJN0qKTpe1LI0pbCY9037EgKdsvtHXAzUfcE4Y/z0P22kp
i0Vhe0SnF3Rj3S9ftJ6Hj/n5/rYoP8B6wL9e/HPd47+dgu3X0MHhJotZpRKlDgKb
Z5DLtgI7mnRf4ewxqlr8rHM1oU7WIxMhd6LGdtTpt9OPZRqZ1eitBXWV8CaYSwaa
Xdwen1xPEtKXc+o/xPmcrhiL9MVpccXHZQQ3W46nV0NbwGf4owDXuRUIcC3CUdiz
UPzoiZEwoG8YNhpPY699RBJctdr11BN0hEN89iABVz+rkl9ClJraqUogMYLE9lV2
b3GAaOSzFr7gIGZ51p0TCotEw/Zsm3U6eQdmd0WSKkLHpJmvruewk3OYdppCXyvu
CGKk9P8TmgBxlzvC36zzVzutCE5uzAnMSyRY7oXinJqAcjfJ7UMccv6ta7Rcpz03
K0SNgfBu4eq/KUDJsJUfthcMpICiGru+1fcaLd3Di4WpZD+/WNh/b3E8h3HsrEQ3
TREKWMle0bRbWNi3IqrrN1LUOl3ctMfRiqW9Sx8xFO94soba5PnZ2+oIOKjYIgK5
JrZlVI6ifRfV/ZEExBiU88FpEqbv+Ab/z9U3CiYX88nULzTxFCPPyUJlTSA1axgN
wk8u53bStTI1Pct9VA8j+hk5kiYcQsnwwrbyvp00IwXxHMGnbRNk7S5wztg4maDD
v4Xgm3PdyYwnwTQgPNBaZhi9gF0keYuBvqyYrXYITjdJ+6hWT8J6a2HrbGmwgfMr
MHO55L4ACs+pk+WhCgGt6wPc/JQhkqQpmdmevyrj61S9SDiebGbcYMOB648QshXQ
kc1GkExiUh8Q6cjc51Dd2tbp9L09xxCzkCwSZ/FBojwbC2KbsruCSxUKCbwYFm9v
4j7kPTOOBauUCq/I0IGtoJHoyAfkQXMUJTw731AinqWrwbkHwQ4pBMgsYCDHu6kt
aXTw/3KtcnMW3Y3LnORVhw6P3AnFwjNipRpeep/3UlDR5zqiFcge072Wgx0DmYy5
nT6LK+XdFGIG9ZXVTsXgVYVcKuWVIlEg79VfbqkOtJQ7rlcMnQw8pHd2HRwUEGf+
6u18nNlZkXhBIosniTyBG+3Jq8kmwgFGHktMh+kHq4Sbo0NISstWK4Vvosq8rBiX
MFGOgF0IJXlk+xKxNNanQ4Sw5hb+jD/thqNqd+mExYpa4jG7rZptx7L+9vXMr9Xz
wtzZdiS3GJklgYQeMyHGytg5ciREXDiFRk7QspJR0GOFY89JNDFVXDUeDbZnh8qb
Fmn5T71eN9e/oaJjnTrdRbGw8/ZcIRbPRiQbxBKzsSlAHuQMWC58rr/i6UF/T9K7
P/KkE2ytC0KK1K+4O1E20YWxmwXNroN5gPymxh31haV8aKmywRqQUgqwerAU1KnS
oxQ1lU06wufIA6CdoQ1vA66zd2OjpS9XZHKd43cP5esJGRSAz6kbpW6RaE2yrgTO
FdJaR+wzrcAkOiTAcxgJLrq3ebUarsuaN82CuO0Mj7HonC7lGkuPBQiJ7I8+WUn3
NRBorDqyYDn+9Yb9h/w51ni4W4XaRFCYHyTwSYCw6mCBkOzNuJdgHO8fIDAiMWHJ
+YezDCXeYXcWx3gwDpWio00zMm6I6qJTIfRjX14V5KtGt+ghJUWoBbbidnK3zCRa
eZQSJqQ1JPueSKKWnB2pw7FVKdBWxRNOh2X24H4fhPhX8fAOgf2fjJ+8Tdb3RfYU
MdUVCBS+c3H+Qz3GVBWPfmTwwMT+eNV2BPyPinSxFJkTpj/5xjwsai+KDybhrqr6
RfJBjIlMSEfN7nEOJSTUVVMhfzDlvYlalKLC+KSmBCwRXOoMnFP9yEZrJbMk+XCE
bp7tkYT0Ya7qI7Sf5Fh1D6vN0nozwSmfzquk/CeE/roulq+sE61aYDXCcRGTqUNc
WmtCVc6Ylu+ao4CCySy0kKnVYL5cx0prQFOx+4e+KYjiHxxdrNRn1li8psNwPqfR
UBoSJg4Pf6lLrpgBLW7OebYxcfqKBfA27GVwIa/C12y0eD8dtbapPepKxtAHt33V
v8IXSOCd2ebB+c8zJyLxiSrNsS25fQvyUQm0MAOrjhXbxuh79h8JdoRhLvruu8MD
VB6Y9l9P+K4iiVpn6pKLPglxfd5z2MJsUiR2OTHujSUQIuBjpCi1w+rkVWk8rh57
eyVoUJ/9FSOynxtQ11+pIjtl3Cf+0UNVEW8nbKldIAvZcyIe6hz610DWNWX1Vt/A
hiMw0Zn15SiUZe7onnmcyLV+gX80ejYqgqYtdUK8ubcVLo3oGA4cs/b4uriiXavx
bp2Jjsv0J4hVJt/AGPjoKl2mxfwPksWP0WamHXg3yP6PS6/Z5ieq/wp7Y59zeuvS
eJnHYvdRrcLBzY8KtuCrt2VQ4eyCJiIzbAQN0fh1Gzy0wmhxBBC3LCKQrrip9FLT
elXcL3MVwBPk3T/A16N51Uthg9tOVXqyQIKbci4SB8aqDpQPqW76WbmuwkWITLVM
xbed6h0YSEDMWisEldMAo+F6pYAOP6PVditt3srpdM96nP0Pl/O7YoFs+tdOzchD
buTq++5bVwEHLptgbnefxPd+brWTQkJZw5b5Yr8JyTe/0gJyHmKml7W6mq9Ep102
OIrxwJ2xEcujW0iYa5lZ301jKrWzlXL6EyzMHDGmXHpiWentx+pPEBsLjwIiKXuX
DB8s7L+sjlwPi9xp/bh7fHNX2MLRiKeG8yvuriH6BAysgti3Uct/l1F6XDIJ4fc/
EB+cpPUNexrjwllrEzhZOM4iWJazxYUcokwwhB0CSGdPly9lXW3kP0QFvey7eG5Z
cU/Enev4mZg/Yvezq7s/m/tIOnsiu0hqFv/HETpaCr9Qo2Uwr4qZafmuKn88XsEJ
O6Z1sv/spb7m6wYuNrK57ng0jkfqsymLrrjU44brGRXxUDo01QBxieAvVhUYbsvy
Y83Cyps/SzcBgMpuoXdPiDxjcH807CnL62BDnebeq2bYqIf0MSbZk+tXc2dknPZt
Qpr21qhVsX8DKjDwxapVy8vfZ9brjFJ6LVxfP8EqhqFQn1wmuAuJzL8nJn0A2Am6
L6iT/mcN4+f9Qfv5U5ORmKxKQMfJ0XWOh36+7bvykbH7dPwk86380FPLFLac1ZUy
HRmjob0GLU4nEutYte1ynYx93jPmXQr3PDMviExa496lU6mP0kOmZn5trPd9o4IL
leiyEqqprctvSklaLI3ElhfdyTdrwUad0hBk3zz9gw2VuqeDt0aJTCVom+4Sba0V
aL2Y23g5bT/O+O/nRB2Rlgb2cAJcHArih4/anFIM2e8ygMd/bpDpmeYcjazBp1J9
0XidGmXdkSe8txMXuSAf6+bib04q6gn0bEaVX5316SqDU5nQ7WvylyT/oI73QhLI
IuF1voc9yzvUGQiqlz21u61r/ZRt55HiTgyb+Q5e3QvSwSFf5kV+ungzA8ordoBb
dNmecxd1bCjeZ1l6V32A9aGgEgJX5u3WpfovTWHmQmHDqkszxSg4PzoI/LMXrWOn
QhTjM1uH6c3Qo8rQgek5MgaWAt2X9fQTgMWQOSFVqh7rIVR9HP5p90JQiCBDiOIi
JdcLMOqMkzin+c6BBKguIxMBvLnhCpdAE/jSduFnBy5znLchanjrEQt28Ws9GujS
76kPFUjQv/kbss8/1fMV8MeWlRddcptzGUWMdlpI8o6HLyE5evdTJ9eSHmuGeypS
NIajYx6U+hJgxLtLqZwBeB0iWx4BmXjz/K8WgrSEjjn5z7UF5/aKY6Mio+gjrWc9
aBQN03Zg1jpsRyDpDjSaqFNbM8k69Ryj4reKxbcV5HxdxDzkoSAQx5y40/W/Z4Ya
AI98su4m2zaEAZ713yJ1QwGdhvqtoDin0wVpHFajwKGW6hxPSr0MrQoffKVN2yCc
qNkHNxJCh2v589N0LuDYMuxg89vVUu821CTVF4u17fHjHW4RltIIE4nEkMxz8GqK
4IiCAnfP55vLdsVQfZbuMJNNcS0rWN6Bqe2krY1GfvHi4rykHBt13MczPpTAWhXT
IS3z3wFPECoU2OftnpktGuFMPDD/bM9mnBe0PUrkjPsfrXbN8FeDsAzu/1L/DakC
qN3FOyj+nE5PxhsWGMWAx505SmkDuhAB/g6Zz0r2areYxr8fo52PPxFCWxoHqwk1
F9K2DzeF0dSAfLkE06vUeIKXcFokxbD+p5urQkfIwRSC6G0huvDVIhViPxdYFUJ2
bzgt3ZsLkxJ5gvXlRhB51/42LUfpVNIv3q04Ob4JV4BcZnl73y0HDBUvYzZIt+zT
hU1zTVQhWvemn0yqL6rfHAbs4oOmakNG5QHkiMg8R3JBQH3BfLnQEluXMM/Ujz7a
0IngATSk7nTlSOORv1ZbaVqggXYJg6ucsk/3hCdu3fTxVBwIKeKE5Iq2sW8edNNr
OzXFKx0iHCg9M75eIfxYDfAznWugX64Da0LgMO2YrxM/DR281fKI5zBMPRvSXrpC
6eytIkw++0mGOhPhH88izcIGwbCF69tS9919Adr7mfvC6OR5Jfl2E2BrG24/ll4X
NGc7HW6Ac1dY4VT+SAem2HG7UdoROaCCBK96OFKCe9PTLgwLMqbM+xUl3pAKoH4z
UfQsDBnNW+Xe8URvpX8PkshHrw7chu4kf8Wt0ggB9VgqkKj+8dyWuv+UbPIrKCcx
uWOFazqceLxa04sWM2/QQuA5ZPseVS3saegXBEQHGsi2MCYbw4dwcTMuheWFo9Xd
67XUYulxJ7xR3V+CZG/wOLQkykETPhoT/LQ9ym2Fkuu2SOD4kFHmxROPHvZBTqEj
RWKQe4ohA0OkBuC8XlA2WaHMaHaYSVJpwFuiO/l92oXem3ej3O2dlnLahXKkLtLh
9+ZK+G55gM95PDvKPZzWqkl3b0/qCSwz8iE/gVg8FG81RWLGidcGytSEMSU7tJUX
kgtoiqFOP65TR2CqGjsieIADsm5d8lD+mRtTVNbCeFrcUeu+RJ69U6l+sSBqDt8U
NdPD2sMiXAYQi76buj0/jTUuJ1eg//IBWh1F5FHo/HMR50vOKsRH/ixBDNeon03l
VfUSkWR+3DE8A8Y/SUvEBBFzHIFODxmfQYirNBHb3W0P0tYIRUcM+IoMypGyrbw3
g0mnd7XRUpUpbMNHCkcgGPIpmGsloBClI4xHUyI5U4+HTGYv9KrIMYAkkTYlcTCl
xy8cDnM3ZYnyxx8jTug9Q1z7UmdX14jwzSqtz3a2HbNgVNbdCTtZq4tyLZktDeu7
Ip+KN/XB4GDAG3spxeGSGsMAklHI4Ls6gj6Lb80y4irRM9RZ6OGwjt5DTJaAqSXy
jswF6B44+u25Rtx+JyVTCuB3q4wvx4twRVPSS++Cl+TgM+J+kPv06sJuAiJqxTh0
Y8N+lJ9+LTeE3prAYNbsE7xY+EkJT/9nmytOYSLj/iG10XSxVriTgJo+yDUiL+wc
0VevIjBsnBFiXLZcfvtVa7K89UVNu4hXAq1oU+ie2NKZU0wjvOWVXLsRLKj76AA3
dcedxZ8iTm/ZgGH0mC8MpgoSzkuzT7yLsQEQZQRlnQWbdXdz+85dSGE80ihtLJNl
wCF5Mdr1H2CUqbFsbI4S1rbPWoa81OhMfh0bUemfjgd0QCNN/rlCk2BClSlYQN0m
nwT1gFdX04IWGRa4jseLlkYzzLcoNv7i6cTPHgwcF2x8HxDeB3fvzik5oMKpubJh
mhZzWjMgW3m4HJordl8Xn903Lq91KC7eXfCoLe1nTt0rMTCU4oERxfVa8sNG7FP1
GCMWPTs+Mxgdc1Yz0ESNsGirpneD8d4nYymVL3tcJKtJnL1ajVZrpcTjWsf5P2R8
MQbvpUc5b0G+ir+sepLSZeC8K9OqrKZs4wImuWY/9F3savVB5wxDpGDa4rp6i1Ia
U+TQ3974nXdk2k3JidPmpx8xsaflweylMnMFVUctjURPBOM2GRWDjr0c7FyWqsGk
W934s8clJ+xxHBLj4cvl17wpmhzkYpE0we01+oK3JzdGsbefw8UcOjTq6paGO5Y1
Hx3Xw3698UPxFkZWn3vCbwbzwxf4Rs7hG9lCVwtJdAC3aAJM94ZPSy0vlZqjlWHo
NmKPy73nT1A6I8yCzkyShiz0gDTkQVYmaiNgERI0aodwPwHTkSKlcpPOwy11PB0F
uNAgvH29fDlBW69xVOOJ5/wvJa4+gpx/7dszhwRPetxRdrFw/KzoNerLrQLHYKEk
FTUid+pTxJoyRnJN2vw7XfzsYR85ykOfPKK/Ksk+7n7iSNC1rYozPgtOmn1dySE5
55CSOLZQR0i7KuhvqCAj+IMPckmnQzQss2YP1nCzNvu36+i0ooD0HQDGYjHOG7bw
1m6ALdnCKMwTyimEHKFeMuy2zPSmZdFfGhAHEFpiEfSV2bOw4lse9Bx4vBETFTcU
23PC90Idsusky708B47zKn9JIruaaSg9PF2gbCaw7lh3jKX/k5kpeq3XerUn3T9k
yb1k3eJB6pzvrXZEy3DYHl1w6AKV8tzmJWmdga8zSqBQfkxQwaZN7/Umx6w5Hckm
JSCTuht1aUDeL/MB3Y9k0lxz8ICZ9AluIVIUezGBsj5LQPZPa9OwsmhNnYtgsS0l
rUrvOO5MTmvDyNh1K3D9TbIPF8SL8Jt1cclHA+c9jaFUrzLKzdVZ8NBlunLwp42c
VXCm6wC8HHO/7U8FgKvdMl+7oLbdNN+ptm/SCwtFq9Zu5HsKXxmwXF4w1BUwI2X9
MIckDaN8rYNYbY8vnfRZg1DBYeMb1ySgOB7/U832PYA4NcJTaLrs5U4ItNKc36le
4I+f1JzxLcDAmDFy4TCYzDoyOVQ/pNTicLUtEOMM4h6ZD8TPalgCgSpMhcNwmGfB
2/Y1eYPrKqC+s60Jk4Rc0V2IfsuTXfyMxUQsUPQRddj9u7o6CcV1EX0LoSu7bYKq
WvCqrQGaWx8/lB9saryTPFttRpBLKX8bbqSUDV5GnstX+iFOg4Uf/O3s1Te4pSSx
vLYSoYQPGYl6k5woaG15E8PdlxsvEU0vIUjhZQ5am4tUaCQyBYP2exgpnaQZd+xH
LiaPpGhR9SBCa/FGwffqiatt3ClLemFzO9sMiIfs2XBhXRBpVuwbUqMOjR80ntF+
dUR5nrQ0F/2NAauAXAkSnSDLkrV5PtcWl7It1RQwvrzccImSmrQ1Lub6ukRfYhe/
is9hAQ0IK3Ji0sFE78idMgzgclfskoKfjxaZZpSHzJcej+Kg7eZw4blfYEd1rU7b
fjnH0CHpZ+ibiF6Fe7cxvGGJRQX9dbqZfypaOmwfhKrJgIosOM2BW9REriA1o05d
rTmtbWiGAUn8jqtXDodtGYK10SOB6n8XILqKj/a/CAHuT6YCPr3AL19NIrpaGKwb
yiK+4yAOlMIJ/oxpkfuzwm2/u4LhTEitHnw/NZFC+U0C0sdsxnAHCTc+l5A8vmaw
pRo0NYzG3bVwSB2xNXaW8F84LyufmrjvkBGtbJcfHXNwX69BYP9pQoByrNESvfy+
hsR5Z57Nyzqe6zCPgMsxL2mGTL855aA9vruYWCCpsX4mWwvC8MvUWuqWNigaR3Cs
EAVNXEcZeazvgAXkG68/eTXpqZLGl7Ec3OKftHsPjVlhXa2Z21G5kpD6n38quhla
X//0FA0cxroI3JrrY2xI4SECUj8tjRKxhD8kZeK3qBZl6hHezX08uoHx9iI5YEh5
xu5IdcpcCQ8BbMm8LQnJpF1rzCclVoAspl8tBU+IVkBcX8Mbw07mmX0+9l/ZhhoQ
P5WRjInOOIvPKlM0xW83I3+Tu4uTV5cPjJL9vdxSjEArAEb3QKmFaZOrvCsvb/1v
aM7dmxOcfIr13jbROUcAtr7KeF6PzVPxSUhYlhGWJ3J3Xwsnyt84+qd8EhM3wMW5
A2PTymT65+0TOiZylkbCOVWrBg3nxAzry40LGVBBtUYUWfLGe6fhrn4Sc2yw9zoD
5KaTjoOgqauwYgTH5rhLUl7MuE10RNjnoRb7sndzMK99tJIdS/iGTIK0BQj89gkB
LvuSeHEXE3iy0Sv4J/KvCOnJKktg8/PuPoGfLRO1wiNK2saNsrZKZy1ox/cd6otf
UWRJZKpXzvh+5NJIr9tUMUJRLOECYM1exuvIcPMtznr1t2CkCXd/Bm7Ym+azDRL1
EFnVVU3796PH7lETk13PMYzBPhHUz9e7YSdaLLuBMroKLtfLmlr+bEbsfoTTMWda
1bmMrt/sA9azm1NTLfyEtVxhjjibhwLEe11FOhj6ziZtQ7VCQzB8brpJdxXqHJnh
E0lgEaR/MPYHhN3TKxNJpMGj3IUdknBJ6GQv4s7pczhHjO1OUTWdAiMS0zW2CAqU
/jNApLBctcpcdFb/jCXaV9dZ2B9h+RCqnvcN7FB+z8Xyqmkc+c74TRtjqGIvXc5A
1eH0Dg9IT7aYorYzd5Cz1hdoEKmliiSOXLx5dUafR8R1NZC7XFtcTU+EKRk+K+ke
RMi5VGUQNGoip1Zd2dP9iIJUih5KUP8UgFpM7WvfLSUfY/B9hYWBPQ70qzYobd2S
7JvJ4dyMIfAEHwUNPTDKsAIQoWe0VKCjV7z9ppxeIPf7xB8NlMSqJmGrofM+bVW4
5KbHEuj8TW4CmIZyZ2LrQZ3JK4ujpXYfKWFt4FM8KQZVr5kqAqNVwPdhZrLI/6SX
8/oWxVVIm0pGZnFyrnlZkZBLJO8DrvN2NtMzbgZXAge17BxdWQPIVS1aWTQmE/qr
h7p4qisWig+juP4Zlq59iywOUDVcek1tAXmknlNDpo4PPAEjdHcZL9Yusew/IvEw
txvZXaUAUIkL06oVipiSIbWRbo6w50OXaGzUNq0rn3mn7VJgFSmdajucFlIuMOH1
FojVp4+HGw1SPIU+MduF3GHs3qjrDBvZvbvOuviCCN/G87Qznspj2YgdyJTuNTLm
9zfLEWatV3JRBHRRB4H6u31lKG1ELf7Xup6ylmVz6GzPE1D55RG2a3I4NgeNwByn
vEkbk4OLy8rbilGIFUp/dUNcSQHUYsubwbEBuHPkUdtoMHEGvKbga2C9Cvwq0tq7
JVJFSg37mfWxf2HHwpNzIzn7SRWTivZShGUGVAcceQVQ48WqImrapvoHF41cwRUk
9rVtm5L27CP1zowodIAB2BRjuy3LPp2WXUGlokGaxS4gy7h2F9reX2EYdmLdrHVL
i6rVibx3Bko0AHryERKfRBtBDoled2EjF20KTVd6wSSUhxc0f7E9UkiVGsTjhgCP
uGGPJFoUS5/X0mq6P8yxqRLMsA1XR8MmyKLVDIzDLUvZRrSHJ3hUJ4Gy/sWJEkyL
gF88iRvbUlT7+epVJg75imGPwdv5S0YkuXANq1h5TXhH54X8DCas7CDDhnsAN1Jj
ADM2F3KRN6E07daAMdTDISu0szHqX4romFE5aG6yeBpvq/vT2yx5CNWHFDfmeGey
rfp5MHz8GXBCXOKx230/7S3pRJbRdasCTrg0VYiE8ZpGkO44PzYu8wIUZbzDl1cf
S90dbS0i4q1OB1Oj+17ZhfHJ/9ncutnLGgFUMvtJ0CSGODqMuoRDwCFn/b4B1Izt
XrUlOvTuTnhK9uVUlNHIuhlVgpq0T5Fwx6/3SvT+LbdqdKOXf7U5M8TZ9LNWlj20
tS4nG+S0MQTKq1wiNOhSa+HGOT/ltJ8PjPAVE7vX1nvpCJjzMpD5p9shKcN3jRmk
Uzkul0ns1o2vywKkdjqb6BcbcNqB9IosiIDyLTGyR3qWlr9TO5ehE7+guac3CaOM
S5ghBia2/nTi0EHP6j3VF7r380AJ5dF2ar0NY4D4uRpgg+lUztveu/tLjsfErLfQ
jhhGP4mGv7Z06lCzlZdZKhEGaphUp4rbe+naCrCallihyjB1nVbGDovcYXjtGc0O
HnIyABxKKZTLcz0ASL2V5obhAhqyjfitHHAI1VF2Medi2noJtlBYbN+XaQhMsyZC
zbkIeSczm9UZ8oIPxGM1kJbZA7o+pJupTL412R/QDyzkNrARXzsbqEw+5lArMtPr
uut2pT3lw0yZA+WSzxBgpKXrgS9iQZ/cobk54hF/nUZZT8xLpnJq7D6M4Bu08hqx
7dbj72nzSPvUmV1s7cP9LQ8zxZ+YzI3LTaAES5288k+2VesSRh2Cz3l229IFAwG1
wsEbiVdHrNeV+hXETmJ7hmRXfaf33DuLvNB31PC1kUEhGH/+FxUUNI3bV88qE3S0
R2+ATFGgY2dO5xjKY4RovHOo9qn3GHuCXkC8UXwjw+M8/XubvTvslA9JT+L3Xr5X
GEa5qinnFvTuZQIIURAiYb0kPAQ7oTyeurJ2x3CzanUL35gGD4lpixKUnAARBp9g
bJesBabFhzuFT6ukqJ++ByptucEBeYSUWJqr1KNmXKjf5H8qYcOeS1pqOErG7XYu
z7WNleeg3SZQq+xWBFhekP+ywPU2D8kk7yyV4Xx/A9cbF3swgVDPoFCxMf66GCl6
jz4HvXce8MUyXsALbC3ngT3yA3efPR8Vsky31AJHRHnx0DSCNf5KtOHVPsbmGtPx
UUCbDa3mfZDGefW+y3GJzPaeVuAgw1nr2XBpcqsNAgLRc4d0N2VLMMwriUhSEN+f
GZzGlrQvuKxwQKpQGi39IEPQkGFrJzkdqtjfyT8WhjHvCZ3y/4Mudx4wpTBC1Thl
6T/7ahy1ec6OD8EQ0MkRr8aw11hsGSEYbAPG54TtQgi94t8HIVq8m7Na/udo+kT2
QRIGxScFWPWBktgf5pNFI4uQWcG3N+LXYy9No1BVAWrc5ySZP0RKUJDV0ilIq+E9
4pJjVX5pxjrzlAfC86GEbFcM5OIiik9cqAAjhoxF46Y+Fr7zTKSfecDpmXldh3gW
7L61O3vl2OHS9j4kOwdczu6U4HCdfoPd88MRq0ZHjqWhPxVWArAugPt6rpLdM6Gh
acX7LPqPBhmoySzidiJbrjDniPY8D71nHkj1P4ZAzRiQNih/2APGnGd8B6UK3eJo
lkAejRttbueLXh3+nk8PKTCWWAg38y54KXcIEgMcS8GTO97hXLRgvqMxijUuOX9i
5HJXNPfDSTxJMTTo8MYXhjPYhegC1/uzhfSgNs+uQG6v3qQYSQYRDQUt79mXiXaQ
nQT5BSfs+wsiK2sfQh1S+WyjapVx5EC647VFjqPh5j2zgzm5zJnHIG3bQkzrOyrT
GGGO47y3ZBABXhEY16qFLERrjmWcNDLz8q0BOgpSTwlCSHVavRL3MH0odcx89BwA
FPQt9J74L4pvYu+QzdhAMRISdaeVoY+/Vt+KB6D6TMYzxo0/AURwSFq+nqWw8bCA
yK1z1wdoaz7IWt1/C+4zJx3e49UC2M5l00Jq66fou3qxjZDnckdERvO8W3D0Gh9E
GKkX/AV6kGKBcLOx0q794fKa7AGHi7u/NfPfBx+dogfbVzJ4S74PRH9jxqw5CTzg
bUVRbXIizD9WmIb626/fjBqPHnFyQq/0uESw4C2gfYVzGhi9WIaDqjsp4LNmcxNL
TOLyLE3DttMk1h/cfHyjh9gtW9MMU8dq2AGXUtJdDACu4sq5/u2fezDPhMCnxzSg
qqq9JwbZniG797FhMVsvrXhmKRxktaai5d9jvkIeW2fwpVuPcBID5CgYQxfK3Oo+
3O49+Yarbh4z68f63IC6YM0gbrSRT0JMo512kLA6KCMSMLgD7z8Q2gS60KqpGMEM
Wp2BTNLJcFqRw676cCmRH+JulG+n/TfXJLf8MhwUZVv1Cqf2FXSPI4SiZc17SwKJ
u6/dbevU79rDXGXu0LYPMyep2r6j32ZKGGk1SJcfyJGKTN7t/uQIJnx6AGAjNbn+
MoSnjXNKg4x24czHa1h3ltoc5Eo3uZaJH9lhVJ71NR4bsMBZfJJoWw/a9zjIKfdQ
cAKzlxKLezZ6X6rX15AXopcDWTLYzNe53ietg/0eAUfrgE9ga3ig+HRGE7tnkJOl
2l7Br3aWjY6SW1YjENRl7r5lYJNP+IBwgnMVm/AyMPLQaEv6R5Neq9Od114sIvSf
MbVv/J7IVWQ2bUna6mZSxI3ZtcqP4VJULfM/WJD7GHcwhE0S/8qOANN0a2Pif21I
pxfVbVTEZtZTcm9My7XENPaye3CWqIEsjJjWZwXG+MHyKxDuhSTmSX3sVHXAvpMY
sG2OMckpnrwZa/xPXGIb0qCDJBPSK21lh1qQiTlILLYvzZJGSU5QHFV66KqCpJgv
MCFt8zZJgS7hvsULxDBMeDP1Zr+hjAY8xycbABalkT22nvibW2e+bBsBKvr0zqDt
W8lHRpDXHpNBJKmpbSScaQEdkd1AovcpEZoOJg2RPYAwFdHPOqmqyThuucV6DRwd
PwWfaiZMXtQFgeBNDwiY3m+44WIsjSbbe6IdG8J/6ZautglqSHGb/K9zF8fGPdfE
VF4BdfQO5uS27Mau6m3dLXh467vPiKfXVxJ1XVXUPV0vhTURkT0T0t3ZaodAPCgt
XYeMs3/AHdoAE6BJx57avuRynEPQiLwbuFgFJvfgCJIv0OxLYSV+veK5OEe2rr2N
Of4EjJ5UqW8hyUUJhZEZ9X2rp4RLfF2+wHJ/XRJFa24rTwBPWXGysqMsZudAWTBd
C0fwCCGL9Ds+Zqs4GqL76E9lC53r5PWaIZ3ZkzQ0ih4rfianvDKs+pUojXit2S3c
8FsrI5aHRvfic71KgawZ3RW6GZx/o5Fp2Juu3z7H0nEzVnTo+NvW4sRfi/9ysFOx
aGVz0MfZq8hrCV7P8r9IHA4iD6xPPz7mCjdeQ+HULKz1BTnsGz6g6cTFVGuB36mf
AconS7wqv4cGvKUtCtA8bpO9PqoXs8jsyAbdmEftUTyUR48C7i3vJqFSfPdBpzpl
B6fE7SibNWnS5yGScA4Q2vrNJo8QK9G0AnY+r+bO/8XiTXYx3Zc8kptVzV8ALg56
BR8nGq8f7EHBLZrg0Zh/ekcOFM4/f1hWhE8OFmuOzNUE84+hB8wERVbJ4gYCYYob
WMXpLaq1lL7vEl6IAx0MW5ksApXYwGJVutGeRdKbpoNLSd2S7NDnBaCMjOHuIGMY
+60SQ4z1uvZzaFyKL/F4M3jXNKZJO8PcNwcv4dD5W5PNxKTn1klr0MFho7NrBznB
N4nbbE0ZIZX12Jnn96/gf4SK1LOCvVAJb550y/yOXp/GxKgxBVR33WRKgmBgiC4K
vEUbb8KAG0IclmdAd3aZsLuvfOPrS4PBZXpCqGkf22P0hQ6u+ZanZx+9Qvf6NADr
UanSEROkwuaqOCFwxG4zeiW5whzGvMsVFxyhvQ0r535FXG86SZToEgMJjWbZZ4LF
jZTbhcHef4quJu80P8tRe+y56stcKvJreW7zZX3DOIec2h0f1PIVzS+KHmO5JSbo
ScZr5PsaWzFRlTEhKaPK4uLZF7Li3fD5tUTTocLhoJiIy96vMbf5v5NfCJn0/KGm
tHJCWjgFsiM0Lazgkjg24bZTwGTmniMuhLjklrEN+8Q5llsiW5deBu2PLBElnq3l
ZjzrCtUag7qn7V4B/KGr+F/0AIX07Ut6Rc+o6iMXGNP5oEGna1NfDZ7TrLEcUwtE
7pSxcaGF9UTeF4r0UdBk/LsUJ9qRFHW2SIKhiWLfoKnPFQJhrx5pO5GoR8c+Jdft
0ruIPAJBrHU/Aoz5fhEkcJylYnPS26347gwUsIp0TenjKsoH6GopPGXyxZeTqzoV
QgxMtxmbUO2gMzIM+ZxgbMDm8YPqGOPm2lpMbZJwFTErOKOqcxPSKvYnhvndEegM
oP/a3ZSMFcXrK9WjsmaaupnshTIqsU7wvNKN6pnj/+1ilSI7QtmDvXEWlXayslDG
uQ7VS/LZToNR5v2jqvQBw5JPvTfMyeNzaXylEKo8rG+sLxr+8S7M51C1SkHn+cGh
CpBGEh/Rs04O5YfzF9EFicPcOpaSkRsBg2XDVQMeD3xBxM4G1VeJGQ3jCd9eBnwL
RckrqFd70K+shjIRZ5E7wRsFv1sYC2ufowXWV4wUFUeDDBnERl016Og68F4jUXc1
5WMJc/pZENWmN+Ab+0/iewrI41zkU7IGZvx+QsafkRJ4dZ4IlMLPcQxZ5naA9yfP
NK9d8ZdLVenVzBCKSfTuj6fWeC1HFV5quVvzOUG9mUI/HKvWJsaPD5fHynROQAH1
SypWCD9GsLmAWK40uepTmHqEov0lQmtqucpHcPXPuoZYs+Aow3j53UvDKfOoaZ8i
xr30PpNONf2UM8s2dz21JS1JlXb89uxzPBqAvW8wpiZcnje8NPHj30hZ4aEWQaIs
UAsdc1sX8gNWTAQ/NRgIUZprIHWDuz+dODrAe7Wio8H2SGecaTR5TXAh0lFdDuPj
zQeVjDSvlgu2uwripz3S1y0HGWdj6YC9AaoQZrwdzz72rjk5SpLRBrZowGFNdtZ/
D9+gAcECs/qNjIVu1e9C4Zph1fNUgaJ7876wtiSSKJ4a83Nz5MMUzW/R88bJ66Lt
HAZjKPlEbJUzhLA1gkS53ft0xwVjQntaeRdjn4SqhZHK/AEQiDY3qIHYvQS0DQ8/
fJhYOHIqsj20C2hlZkBYKTSqFnVtMQXC7MV5fjKRMyJ3jWwTZ1ya+JlZNRqoWdAe
8FxJY8MXQVx21G9D8HNIbmq3QpfUkDaBlLQGGWeEW4aPgPJKCb3l5jGitJ+zyGfr
RQFYULcgiqwho66sA6p/SfXglwgPrOY4Zqo/P8b88ULz2op71boY4dkbVCM6GUJB
iLqfnNEgcw38IZoxN/T/PawC6jXfTGFsCXerx5N7uS2m68fGVm+nF7wQEpofStB+
XZGmc39xcVVeZJmHWnVYinnUtdOV3UZ8rPEz/c/e2fMB3JhlTOmL2gP11Uk5GgNI
sDkjxlNIF4YUtqmmNamJ6S3cEKi1BG7xNPVjS2/n7RBIQ7PGuQQoVAISRGmNxaNd
23Jg8mThkOvEpnYuohkH9UJEy9CNKODKmRZmN95BOMA4nBcmXyYwZCdqbo0o2+0K
hZM22fB7DFMyQWEdVmScD3WEDQPMwZ+LHbh3GSt1ccmBzoLy/rjvwVUd+rLaXyek
5YiifGQFigMemUFzzP0E87YgmAXpGo65B20HI4Znp8fzYq7AkrtjQ5Xe0s1oXxyc
leNHdgP7TTHOxnEoyWNlCAKw0a300O4VUr284lSm/+0Yb0sQNa8DH6cEjKqNocdU
yGd4BLVlWDNmA13P+2JzmESeyimD9gCKVGWS25dPC1uva3MzTazSY+O9Lc5Ww1Je
X/XRyD2wWf1QXiXkZUXZzE8RRa2c2XoOYIHzEjY/5vaxnHZmrYxT1J5cBNTmiO0g
mBXvvzmzwJvj80HHfKQ6KlpylkZi+Fbsg9iF5G8bw6SGnDySy0BPcHSrdF3EpPxJ
RsvPG7K0Ziy8a8RbDqzy85McQVaQYSFsOAM4Vrhn4XeW0lOkSyfRHQCotvbu+UHI
aPW+XNTZ831gl+xBda7Ooev7pBdFm/bfk5f0tDVgpsnARrghtcZVgWtMczG1OT9P
2KgBgzzqiIUsnJelWj7dxTIzPRnAmf9ITlSVDAtiVE1/Vn3WRrNw3HP62IgwDUTt
ueQM1mujHVkBJ58QTq8+jwYCc+RVqX5MKbid2pn8VeaupgutCFufTrO7XZ22/aQh
UgwKVCi0i0YoJfJwvsdq4zGvve1A+lM21anaaE5qPV1tQ55y+ZibETeUa684MYAq
WMFMqMoTuFGIfav1kXAt3MUpg0TdTS+QfS+9jxWyrFpE+fM1+vESoQXAwuzAv09l
IerxI2lfMDglYVDaUc1u0r6xNsYHW0LqiVZCSux2jQ8AwN8OlRrTQcq0lUGGX7ZI
2dlilHDUe8/x3Ud8yQNUngR0tRDNJDXNVRMAUYq9X4xezWTTekFMgBBSIaG8dUb7
I7J+jQVx3Oe219iAV1dIcayDChoSAIR15fyk8bGqwalov6eBrhft8eD+v0fFj/L0
k+YiBzzBPLt8qIlmNWiCP+hSdzRVFSFPt6RuK5v0lKOyjOgJTxR63zJpFgkl1f9x
H0ze8sWvCySaYI1+0RFbTeHpPeZtnyAMa935gY6f5k2pyopJHWCRBjM2JerFgcnI
hRvCs3XVX81AFXwEJ1q1UFBKORLmZI1yTRfixbYaiXfv0oR47i2BYEkn1krLisaD
8rWMbi7yQl/ZVXD67Sc63DiIVw+5ri9SUXaFqoePOw7oLsoWk5xO7upnIXupVcG4
UX0kpzX30K93VrQcCYP8Ew+v6qsaXw0cD77VTVK44EUO4WnUl93tYo57etlsLIyE
LhSnYUcu5Y2WPbC/K1gW98h9aDe0iAhg2x5AHzRuBe1cJm4QnNjbdUSQZ8QMh0gA
Lv0rx8z47byZws3j6TAuohtkLEdGiaDSE2154y0ohC+Lu2OgRt57uS68QF9XqqIN
qFij9lUsbPFWF88IVNkUcwATcucGmM1MdIUyDS+XbdXnGtlTFYLWRvXqL3G5ssHn
DdwmdHqQSyaKJWt0ahmeZRWabwLkojXxzLpp+jSPDOF+VfzaP14KFbWlpUbGIBDw
ffAB/HkZ5Mv17XLojXD4K6VbDId16Ko61iCBT24rRDFAmr5Vm+ZEN/Ca2dEy2IbW
X4/LoN1fwJWqvMKxE8xdSNNI5scANiEgQXH0cTUPsrGnELPUyvLWbklhbK7m9bur
WVOxcOwYQcf5P+esTH/zPCRgTxNdOnjF3vjuA/PLPaDx2e6sISBK/P+tIVNMImp3
7q37WA0qaK7QOLJ8FPOb/DbZUOiUTHP5BK0mCk5l+LbBQC3LsLQ+vNuS4XQnVLto
fthDfpn4YkFyGs2AGMb2VrcHcUh+XH7u6FW8iCHEmA2nCjCtJ1IsZCytikYpBrJV
F9ecZa1LuzZX1Esr1ynqbRmls6QvICGlKs22Uu626S/ufSlayB8QKd15mjGKVm1b
trV+HoL/IQsBAcrfiXSrH+BBOfPrjtE9eYD6cg9P5RZpNvqLXJrDwp34uB02Dtak
LLxZjX1vx04iM7YXb8NGbor1bOI0jy6T//ravS2Kb8sVxfv6lqubRm2oLp34xMBL
B1NAfK6HDdM45ocpcQlbYh1EjMdcTjMFYOkus8ZEXhUfPehWmMOLLfYZubbqYpMh
l+8rn7PFdvHyf1BKHHGQYUTKd1QyoSUkuWbLc+C5RqezQ9mW/8JQ8Kk7cXMCHge1
lf5+E2QTyd06eT/PPgbk9Et6hxE/SyYQ3vMwM0L7HIhxD1lJC7quQHcJ3vadI9GV
i2tJTa0J67kbV5K97sQJTN/yRUN/UD9zAZrVTZnyFdrHhxPEQGbat+zG8Zg6VNtR
ilf3GdmkeYcPY0Y6TcwHePdAwuNTxY3V31iHiz1ugyGl4sVBY4UZbke59vHK20oU
oKoU7RBwNedVO71rTokmfIWYtRTMsOGVPjgvtcyOCLbnrG1eju/V55KHwajeAbOZ
D49ESRQBrW/JWKYKqmUdcYqx6w5KQ0LCg1EWpgguBKHUYhVz18IjG4gaoT5Re6in
9rAKuoHKc5YYSBpHEDqqK4EVQ3hNZA5wL4ycv71nM0ul1e9rxyCmj2u4Sb1541xU
9BwGzB5q4g+GEOPoQUnj5pPW5s5FAhuM44M/8lcLk6P6gq/6zrA0PEPqEfwasYGD
flsS6T9zKpvjesADL8M+o7x0+vlve5fXr5anyBqJ14jBBzSr9agjPa6/mlhebSBM
kHtZ+YiKIB539jb/G2VTnuK0PiMtv74TqAdbB1NVXN2zfH8ee65mrwI07Egaonwy
qlWjnfZJy5z49yvmsvmcsM4b5OOMhwCiZzfzc/VYts09XOPFW6R3/8hmrph7iTUI
CetXJX2tgqAM44jI8P5nEz3kDwWvQzxQxANGp0qLFLiW9H0JQX1OpgXEMGz4JM3r
jU961zqRrshp1AHOvKjTN8nFJ6U6sWVvj+fi8DY23l2KQ/UHreicCXlCiwyZC12e
BZHZ1KbMgBP9gLgMnF+vRm2k+Z96cCKXHP1/3f00tV/Il/1+xnZbsT91W6u0RRHU
osENlgHZTeWHUJ9bYt0EeMhX/qzNAN+QqQfRkhMC6gAvTkNKGOzAeYlxqNG37oZs
GqenuiLsA0+2B5lcwBZyqDnJ7YqjT5JbhlAR38SkXxeZfQnKOqtQ0x1s0L/AdF8I
y66MpLryNgwtR0AuFUnR7dDKiy04LMFs/9jxHjnQ054bDNFiupafkjzZ/KalspKA
vd81RbkI4149NTVW6n1+xNwhUXab0T9wR5byvb1JRxT3j8ZnjwkCkHHJYtf3cr0P
o8QP3ifgtRU4IjihmBEHeBfzuoOi5YvvI1fOVAtIQSYpyiMyygHSRovDUUekWjP3
wPFvk9yADorSaDfXF8rsRFvijvcSvhWghOAGEFRk0tXZzls75vgGXgdpd1Ikltfn
Nr39kUl/py8/HdBhSdAd4VbelNHSJyNtjqFxhfH/rp3O9i4VNuqnch7dhfqeZfMW
VsIiHHnIlN+8nIGeicLJ3VfV2xk3HQsN5mre6zSLxrytJOp4/eeqeEcI/pctwbQB
Uki/Bhoo63UtumAvfULUcIzY4ns3v6tIaAqxK5vy34KLpNuXwX0jykcWzVArDYAU
0GxtOTUy4edjZZa4yDwgcW1eDEBxTJGFYWSohhgxU+bQIhWAM+YD97jLRfL+ljTs
S5cVObnzD0tPZw29D77BJNvh8CyJa/aIs3wZPSf9XxwDe/t9s3jtCWm82begpahS
YC2MnIwsO1OELFUKqwtuz+MFibDubhnoa265SBO0oENazaAMntVEWnVIOLclHM8S
tRoBauSoOONiQC2cFAyzv0jrzpaT4K5b7AWLJpLTUDms2sAWfWmTFty4aRV5Dz44
TfEww2pp9bPcRWvKLQ6rVy1NLyhLpv27QRDe/5VkGIPY/buPq7wZb1GpNCxNEpB7
5I8nD+sA2CvyVf8VPHLMXCjB1aOPSv7r/WP65oDcu/IucxDjzTl26VbEms4Gyfro
OCcyr4i7LYZthE++ozte/McSedQ5whF0ktbqr81Qc4dkUSKtKRR4Y7ShhRaIzkce
Q65r71cnWcCkix91e3u9tBp3QCrTU6BXqlGHlyKOWBEM12wQuin6x6VniDg3jbZ+
qp9D0I7sbfMMO59YBgRt4KjTi4JLYS+eBOIWQjfsKbSpU+1c9wb/CDPjL96pX+jU
BkDWLQpgbuXYS+hb7MTPmAN3i8JqjWCapOXcTTD0zRFt+/8a1amoTS0xXibmPgc5
JkRQyesyJ0Q0HkoTmtEZTkEbIWkHKIFe7u0QLqUtCA1RFMqqLJvgT3HWavcKWVrS
44Sga2bnNtt/4EtFgGO4G8LD2SZzZuY3z7bzvGGck00zKyCQxhQ4hXjQGtqyOUuL
ExfU/CFNiSdJwm4S8NrheVlbTUpjM+9aCuKI5+Ng73MQqOFWyJI9BvnQivULxwbn
bAgMc+GatY4yoMfG2YisOcZ110a42TECCO/NxPZf5oiShWpf4FhJIKi76N7nxUAZ
27Uuxs/ioSKxot7BPyVRe2NvLzxnZ9pA9sGjh+X3Crs6VyS39xYrrswRjV0J5BHV
bkxrMBazGGLZ6ocVR/7pJNTc4s2VmhXxR31OeELvjhWvLIp91RHTML5VxHYSz0T+
xfNJq2QHiD9cCPK5lmctsq6cQENpJoAo36KwuhBgSnvFdD7UpNFwwyYnVCKMju0B
Zvy1Bl8RvYCXkMd/nqIsViBTv5jpSxBzcm++6q2bOVVOMJvUMdL/ZueN7ktqlcHN
Mkw9GnrQzVP0HK7fhQwaYc4cBK73VKTkjR65WZoZcOxJI04qgXj+4e5sFxwqUJQs
ytMSaczux2+vyGr8ENVEZ3dkNk/+Acu6HOQJb2IOlgeLzNti4PfeuQSHTiXj129M
w9VhibJbcj89k5KnZ4ti8gRD3QXxgC4PCYB6uPzEMsHiQ4DDLYCRm9doBihRwV1g
QYO1BHcVwNK7fYH9O2cPkkco80usBOw1FWxXkqc8/JdwX0cH3Pe7qynwLLtMj8Jl
1yB+MjfUW6thm4WQnw2dG8zWbdrUW/LLZTZ8S+d2EDBahi+yy0zS9dUBDRExrW9V
u+21CruUCfnKhiQcsuoNcfjjBmI/zJNdZKGb4/GVjeGwbTmmttELBaGcGPBA67ga
iveq20uV6Eu9xjv5YkRNNII8SBjCkNnKHd2AXGkJ2kBJJfAor77XykWxs44tQX0a
kyfZeX85IV8w9LCgt/+58mI0WqHtgzXNox6Xo6PGS28OVyb/sCLGmozTOT9tVk8G
yYdBXxS1An+k8et6SKRxVi4av9VfHDDe7G34QUbeyvFv2fB4DkXm8T5xQ/LWymBL
El5RBMw9cxWjGvgpM4u1loX8/hDE+ulo/uMNunxCSueToZveLFmMPa2hWrsSB1JX
44cBfYa7dyejgUU7BeMB4PBFONaJc6Xe7cvsqCkDvt242gol2p17lfSY9LyCZqJj
AtF5RzKzOvPculg3tHK3LfsPA4pO+daperPuAT3dMl8Eg350DLKzsW+yNJoE29EP
sYaAWhpOsxj2CtADGxITmY59wOBWpW2RYehAb3QR0UR/nWdDXQE1Ie0Ir2UoAafB
b3mHN/H7sDW+5oPMDPBn93mD2//MrKu2ECHyy7PAEYnm9QE5uZNbhLG5YmrHcrNj
qNqNHTwUoSRbwCV+rvhQ5+IkzHiF+3Ue8mk0c3opPuGNxRSBjTVS3iFjR53nRhBz
FzxQUSJkqEhj+vQzpwetYeJ1go05DH5ueayYs5qFAaEpWyC5dB6BsR+5lS9r1Gng
Wlxo++2ArfRdu1OmoFqnt/suIpW3ySm7ApxYKNIEYg49mwwREcuo+m+ElsXItYL/
JT/X0rpa35Wf0kVdZHb464AtxwuixVcPrz8zWkADaRFbRot0JD92oB7Zn6BchL9K
gEF59hmi3YranqObtV+aAzreXILvtcjIIGNToj723YeDpY1hvxjhp6ybt7t05PB3
usw0WOzI6J+ilwls5QLC9qjDgMKe81dW5NoED/q8lDlc1Gp0pPXHXHuvlFgs0TpJ
sPR3kNM8g20xLP6MVjlkHTFigSOSi436xttdFEL/Y7rfNFX1lEwrHvUx5FbHGJXz
CLdYVtkDEtmfHzJSnrNFEWuxM7g4QWTq4+JbeA1tV+mgBD3cr6bRg9pG5nvWBZ9h
UaYGs2AsqoS0H+gtDw7ZKeq7I72WCESCMcBa68IOAPgv380Jrqm5Y1cOhUGnq50L
8VBVZRTZoyyZ0SOVu5sA3vpVTUYp+hmrSStN/0Vxh5xxBfOidcwCqUyAbcFSWbfb
LN0F14CGMJga0qhASKbjLGpV4mCGKxW4ssBERS8fLv6k/8bTse3ZbufQb2F5HpLq
2UfC94RwyllJYRUH1NUugMr5rCfNwqtA5aokHHDZ2xPBP0Lr9K1DfVtUviTR2IPV
xRfI3oRMmmmByZRZvg1LGgmU60g7rhdvPQrXLA3nSlMQMm01PwOBTnPf1bPQMP1s
bD21EK0oeIIfGd1AKiUrUC9wcXVbWylyL6OPRWuFAzPdvNej5gsgYJYEUhnHf2/L
9939HrU5w66TPbIPHQq5Bf9Efa695I31jsIoXsRWdJRCSwwP1PIXcXjbxXsOnYWw
2K+yeoj4TV++oKK83yvYtp8dEKTMSd9gYlIYNek8FDnZMRciO/q2UPVJCK7tmcR6
pjGv0zwDxTyR0tQVefL8pgKEb6BfFPHs3Z7a5/YdHfUH+WQK1lj7NEtbjdNrGN/5
QbT0W2T+nMIL0LOqS/Udr21R6UNTeV3pBqk4jXRI0vfBanqHrc4tbFj4+PbFzEWf
g5/aLfOo2L7lmQ0mh/BSz6MFLQ6nFSutRBYXMzn2zs6gADdjI2JFHdC36G8n44Wq
Sd/005xqWG0AsC2aK/064rg59xI6ce5jOh33NomM/hU77KsWYNaGvi2wr1QIClAb
HmQ+d7l2eFcoHOvwEF0bTTn1EY+0L8i6wGEBg59G2AkH8zUWH9PLly7IlzCUWCZI
za2fcM6JrX/R6fvRqEGO9MibLBBpj43hh7vMDpCZ/BLp3/AlHEQj4NTtFeFACdkM
rofCfPvF1TCxXwcyq1SOVQeaXA5WatJDhfXxPdM464uoVT2rn0z3TWfj4IpbSRLT
sVQKdtWppwQ/Ct1OytHUrcCxX9bsT5scxL1/NVyK88j08y5mkAICmFJRQaPEH38X
B5/n6uYuEj9bi7Kp7lyhVadtAOHiHkoGH/I3Jcgu2o8CaYbIK3EhwOLVQgvUc53w
OdJpIg1GbB84j/Bv1Z8B9koLRNRhfwCHNycrFgCaAzS0AL8ihTDclySq2f+Qnkdr
GIKAPOhmmr56dn/V2LdHdSR/eASMN1bqye+hZZhCaDSwBA9fw5xJIyBNb/GGvRI3
2lrU3li3b+qqtzr39j51EtIcd8kVffEOXnwNAMtvDejoH13ZE0p7rM63DnRxLmfO
BOmZT7xF2XokWdkq6XqR1Vo5h6ockDLSaMsrxW21mrXdGvAJE7TDJDMuhr8+EMxL
xKRaZ8c4+/iq9a8OSIbKeLvSQYU1UiDl3s+Xg9jXj6lXzQqQTwrqg354DVouHTR8
i0aIT0NJTHmiiS8OreMP0Cg8KzwfNtvVpggPI9kfpJfffirPND7nivnGuyrUx41B
fc/KD52O08ln4PifK+RU/ypQzVGH3ncROk9+h8vjvIrvV8G7WtFu3+sbrqXeEp6N
kC/IIMgJLAh11mgjuCaElzwkhI9RP5DjwmKo1aU7iLSWVtu5VCq9/3W5GU1+40Vo
p7angjQ8KeNM7WzotFfTc0Jkfr4BFchRdRBxf8oqhRIusLBv4142wYZpCN75wvUH
bLHNe+qQk1U1nhtsl25GwaszrsmYKGMNaEy4Z8avTrEB9mD+MCR+N3w+L4mQUAH6
wxp0rb0UDwFZ4XeuDtE3naCmWfpP2azOiqPGTILD7BtDYUqc1EDfJKRUN3XP+cfe
0ZyCmN1cmzU7UlS0u1o6wEn2Ax3BwHkYYV52vWZg6VYNwzhgO1MZjXaVGx5kDkmA
4H+5PF3rrz5h79v3R5fqy+rronKIF48dCIe46ZPMmHWFShGlN2FY9N9ZM3n5VW+e
FZUx1JJ2qW1S7XHrC57EIFxzxVM9l3ys5m7iZ297tjA7pCL6SfgbR0IvLYVRqY2T
M8VFTvt47SMAQO1qkigomPrQmxcAWNF7lf/Dpvbi+3dxY9DU1sWy8Z2Ydeni8K5q
kFAf4GX6W/x++UpVRCPUl3Sk89zPH4vdiMwQOx0mFhRwmqVywmAOuCQaERoHr/Tu
uSEseN4/LTRkspjULgAGW/3bwa+5F5pDv5bK/uZEyzMy16JuzAxZsHXUZ7VIgKup
uLTc+xpeLKGIBFBnKqNyEue7kVd/ELhB7lZ8C/zXyPU2MOkrKW3F/aKV5oItNJeS
9/NXUZ6rrZUlM8CSgLnsLjYsPdlek7HgzxpO2/2fIb+wEO/rpyH3zABx8qmb+Lyz
5+zquIN7uJ8yiyocEpIv9/0t3xoY/cUJmRb6W9FSJGf5XPUYo7gv/UKQSw4sg/tW
cgiZuRfLVgZ137e6U0TGoWtre7u5HoAyrpEJXN+VtAQsOx24kqjXsRrvdp2GTVt6
lfmiTm4RpQsfsucbmIH2aRmLLqSyHAIiJL+2jBMPWeKrT2+Y3UUvxsk3Vxe4lx+7
VwwHZhXX1jmMKG6N+JL5au1Qb9hRsumXYtSzZczg6Qi9Qsc/y3m122o2mxufX8GN
0pyPAWY2UwlZ2F+jti4c2CkTyAVQO707t8/FhZzyDh+AxqbFJBRhxoywzdNqBfWo
iuaGeJadpBt4m1BLPnmY2mI2ESO08E2Wqmj+xiOIcNcfQppCLmIX5R+idBD+rrGk
BTQ6ppFxH5WswsABotAcsXMTCvPtd+prsNhCXCU6Heniymk0mtohBIsWVAVj6qi/
rD/5OyxK4q7el62/dOz8Jas7e9QRYpGK27nv9Ntnuch18xwOBpKrn9zK+xkbhwkd
UtN3aF5pi1QR+lx619QvcRw7xagDcFvxbBOJyTL1csdzyyEjFtmAfD1z1BQShYym
ySfLhZd82vSnCU+5pYV3uoR5l3s5BjQKydR6kASu1iU2Sr9ppbWH/xSn2nfciauc
MsEkeMfx66SgO1Nm95IRvMnj6S89vXoWgkCNtjGb1ODnsKFsS5JBONTgCnMzhX5m
tQ7cl67OflhFySH6drHo18EX4OCLVyRPHJL2Es/W8aD8Va49+W5APEiruWdmM48M
kq+cduzp3Ln/JTWSXSfKUIpoOJTfHNX9Fk5Clk+/ve2dErfz3Twkg0468AwCLOGx
b1KZsPxGhAGh+ARK08A+Sz5rwmGXTYZDv/1HuRvIjpm7gNKoimcv9qi9faMXREyt
hDcBunD4l2HtqE0wPfV13XTCBeAvA4/aB+90fHz3XmslWqYKQ5jx3pNNNqK0MKPs
Eca0urCBIFqXG6PIFRnErXfMs2/2bknKMUvTHp0VfTM3v7FAJt/K2r36PlWjwtmS
8UQsXFC1Z+4tML1c94B5l495SqMxz8H7CKsqYQIHfbPbr0KPiSedZc1c3tP845om
cGHE0iVj6iF3OK7IzaBc/Ara38lzEWO3BR12JK9SRgVnUf0G8L89YGaQhAIeCAak
wyxfB3dfR8FD05qHUN+fyRgHOnCL99hwXmQUonENOpcNmdPfVGHYZXXKoTIpmRGX
VBEvhetAPZ3FqWTzp/fx8iTE9YjrSywglJJmWMyXYPHntfivCktzQ3sTcTSzPwL+
4aPStps3FUs/qQnaK2orbvJU4mwYLqqFPynDdyvfFdcT80N4pRdhWMaGafoD2yle
k3/6wySXqwPbR0LFCgo+QAMlUp+fo098qUgOFjcX1RX6ocAAXVcxqsFtZ0kAeTlc
Fu1g7PSB9fpLMk1hHQGBjKBHCQ4PyNu9v3lDlgE1KNKGF2wlf06i69O1a5DUXGQZ
qz99asU4zsSusH/xlvkIhBsAeXC77PBPwIdUkXJxT6AWeNiE2rx6aj7enbSfwLqi
7GJtK0uPhrFmO1caaRPMLEeEZV1Sk6zdUi+6Q56SLg+z/tiZWkEyM9/bSaNGyQoD
j/SnLbXUjmiw5JrY+eKBkZbxtcb6x+xE+pXv978GAQVbOVm1tuYv2KqTEsE6Fc25
Up6PKe9Gq35vEa0XTQ0zorpTCj3nOKmNpP4KvvqevePWmlQcHjwi5lOI8GgvL1bN
T6NgC4wJE2hD9lTLat9MO+d1C95K9SO81VWNpPvDl8uRBjuJh5FalH0iYVtFM9im
GWy/fduRE8hvXlpU9ca6KInavm+Lbk9qtAgYwwTMHRpRuMvD0zLPI0RxWKCcteCB
FMojO4c/QCHgMChiWLxir5zAUH7D39pMC8Nu7hDJBbE59Q1eMrrG/c+tvlabX9lJ
4GbxlRPTjcjn17Hg1vT8lfgqmVIGZi8hInGhcn0pEcs7ZZr6DT9UEH1i1Pw3+aGf
QS+/DSpJuIoWdXnDEThleAx2OG+BNBL5LJOEWd/QjP7QK4uOVU4OLYzg8dLg+gcl
Oo2fLMYH+W7hJ2XGAiJEOe+tCBJUYOA82WfMxw+YmiUy5FIP96UuLuKR88FfaJ5h
bd9eMp2B48+pv9mnbV9BgaZhX87d9m9Zm1TcvlMJ+Ww7AXudoG9LSp297P7uLPPa
HAGAS1dM4l+NzG0MUdYaTsvToYEKKj6ZwkE16iXkqu15RI4gY9PbgRTxnDqiYLiK
V4n4S5uOAwcbuRjiZ1O3UdWyjsteR3jD4U21TIzh4yyFL2AgcvQV20xce8FFGjNN
KPmzFph5qK5Xo8z+j+2hducgrIyl2VdrVgy5cR2DMAy0TUwrkS3yaCiKEW3DTeWS
DVHfy4YgeF6ICTHBXKqzApgm2fAZK21hOQg3TLVtSpwu/ku3C4Pa9p899HgmmYr9
YTRNEMIw/WHKv0nwLs/9LIDkEkoibDcReA8gjvQJ5w/SBkjpS/cPbM5Y9Za9rXvp
3O8B7oFBLSvGOtRqLP4U2G2G7lxxJNMJ5r1oSorNdjhVBz9XqFi1isDB4+PT5guF
r7dNk9t5rYMFQuLTRXiKHtD6Jia8WxoqtPgteWwbFPO1kmG/tRzL2ylMFUFSTfLv
cxZc5TtANvHWvNBNT+ZuzUIcbrYdGUnhYjUcWrqpEEpJEkHejc88Uo8qDXps9mYk
DTmbM0bwwwydpOZhii+bYF3PWneBm8Ud9wpRGY38RJmwQqvaxrLGYhhqVCYTH8Be
valOEi0NMRrOSRWJe8mPreSEAtdMqha24Vk+aSuDftnxpjSEPl3eeSALbwVQeXUW
ab9pyLjQ36hiUyHHzTUroyFlgk1S67FW1UCPyTS3DrNePjyZdDglyVCRoVe7G/V6
G2g4rlsOx431/c+vGlbGmTfg6x+TgrwOFpk/Gcr2i6UlpIwHvGrTLPUG18pdP2qt
Y2L92CyYd1SoGlFtfE7fgzC4yJRnpyitCspc0sCE1ZOknJfc8YJye1oNIiaFjllA
rJF/vmu1/UVk5GJtk9Gg243eMAAyBs9qgRGj7lhDzC0d9z6JtJg+4OThIFnWL8dw
ect9ib4y7QgRHn43fnraCl3GAAr+2B0mt9rncYYvxciBbEko1WWFxqmbAPGXTwum
wcjKwd1nsSpghNdWnDIu8GfXpsSeqKhlD6/S6BB2keNV3XzMNST0gJAkdWnvVdqQ
6QR2qEpNSWExEQx2yb/E6BbfVp+/dQikG7tv1DDDIXmCzkHqIB0jopWYP8OcZyCt
w6NfJnHiKh72Ep3UAMEudBH9gjwV9YsGdYDvOs/zq4KBwloaXeMk3R5M6RYfwUXk
eYV5j+V2ocgtXwem28lRfN9VYoOU2t1nlFyGUxvLJpcNQFR6sqll3uq60lvvb2g9
UrMIyNPuVNDtWHilgDeoY8qiM+pIYi8bqxKq7xgcodii5SJS1OKb3Bb0wGDa+UQi
svFi55wZiMaG1ICznCYkjbq51sJ1VSeQO0ADOA1hyiSrLXFkz7gFECE3o4aSFvsK
zyDast8fCQswi3QzjcIN8YMtO9gRv2f8mdmg1iG73naa35DuT8DLVKU7/DNm3F19
wYmv16VvyJOfN+u/cDLIPd7hO48gCmgtC7aIToHRrhanH2x8M5MejtMRpJAaM0e1
ZSGUI3qH4VwNXQ+bOU4BrGVfRxb5btglcN3agsEBYCQT95UVx4d2okqKzMHfQqp0
uDJq175zbhA2rnuCd6dJlKvwjmoCQdf/T1LBcucT3G2ZvpmdLM4fTa0AKypXkv+j
nPTXBnxYia7XxjDlVh42/7pM2ilw1Xy1Xo4oYmlRJFGudmXs4AIg3Q6oY6vKT5Az
y4kwlkGRkAw+GhHlKpsXPQ0pfOvdbKYoiUqxk547OuhZOybFHVhQ/JgXSDZhRQaZ
k70yCwokN8pvAXyatv9mBdC++WoTG/K2po4dslafAmVwRBOYVu8MI1sgaDclRgVN
WxEX5GqZ9frDrI7vJvtLd99g0HKN9ViGznAEHJbmErd2lxRKPV38EEFkzMAJ2xL4
GtZAoQhbEnPIohizw1xyO7k9qqyJG3rPiRHvhzrT19sRHky7B0ShfRHD2vY5Htv+
r3c5jRxNan2tZvyqdbm0zhAtTzRyKgMAHIItZIhs4FsWqL6tX2vfpW/NQbtsB2o0
0TPTphfWo1p/JWxuzSF1f7cEdjgHS/ljQTxxZecYks2hlvo1n6r7ZORX3zqpIRdV
lwySUIDHe/BAAmMlWiVZvDioKLX6uVuPqDGd11dOOzyetj+Ue50BSOTuoqos2yTb
vB1dztKAmlokoL5QmlSMSCN0Jb7EJrMUbWIgat7QQ/G4JaIlm1yltZKx9Rc7APLv
M/Bfy7hLTV933JkA6aWu2YMdNf/zzG7ODpVJyxy+lnAwddzhnw7zpSp88lJZOnUv
If2hOolqKf8MtArpszASN+4Y4cqVsLxO9KbNpmL6etsVC2JahtCe2RtkKOhkIXaa
qiOumPQUsCFv89cRKffXBWWurtza3qapvpq3Ngp0FWJTcpKIPSrYUHoOM1MpAaik
/384T/0aOrE8jQFFxNRmgNVUqiW4CcKHcJkkcL+PsQINKqALbSiZdeT7paUTsCoI
pWhOBcNdIyCMv0xdtN9fTJEbBS1z1q5KBc5reLvL6OTWYHSbBjYtHysDAnPwE//b
uEF3DPYhq1xA6YByKcJflmEMRSMJ5G3JT82Kjfd0FKAGD0LPoicIPl9LX1iJs91Y
S7Ah+mn+Ycexg9vTudBwHvFwEc28yyLyk9DF1m3EqmC0j+URf215MIyRZg6sw3rD
vVjK/gQTtHVzwinzLhwPapxNVhvGHJEKUmxPsZ2lOEm6njPI9QWo0RdV6mZCMSK4
pLjBnVAw4kbWoZmryFSxfAa//b+1eLfPGxWwpg0UYqbtTuKlppmZR7aOUpMUPIPy
ZoQ+BQ70OPQ1RjJfYvawMvYR0FTFd8NjA9rgUm1A5N0/+L0YcQn1FLl2NBIkrJxa
yaxF/f4HfJbCJpHWh3VnIlpSYAfoJhI8NQwscKDDF+NUTkB/ABYRsD/vkqXBUsmL
YIN9aWa4PXUXGW1j7Vo6CV9c5Xr7y0KpftErf4xpgBPOfRdMBXM1dhLOxEND0BUe
i2FNq4N/UYCRlq0z+Prv78PWSEIZJhg/13h0OwBo/Pz3dYd0nv1NB0vZSUi16dsQ
T1YGGTKLbaznmDJqYbZM9KKVOGy6Ag/MXinieBtgi/7qOpv+W/r2NYJGtjp79qdv
MmSSOfGnrdyKe2z91WfN1Gv7e17ci8mCzKXVdNDBSyhNjIUqy/iFBTEmL7wVgY3M
edVSCkeEoc2uHUo0/yeHeeB3+ZaTETAT4KrLW3wZ+aweUV7lzZi8pN3xNzXTJp20
hS/HYttVwi8BqGDA/REX/nFid+aPTivb03E72x5ZPOPfBRDOSzN/V60MNcjZw6M4
de2p2DIE+SY6G2XijNmMaDkzch8p34xSIhKkg3PwkROdrrYsBPJjvVE6NPl8tAzF
1ZBRvIXGPscXLYynq74yD25HerYmHuHDzTbr0E4UkI31RNbQGPhsIJwrSsgqsbu4
eRNGT8BG9zqt0Y07pRcSacznpfDsW+v8PNHz2hLp5CaIVggw5vLqYzxhStRkf1Ra
RfPt/OysNP23FT2+HMNGP3UghLz9U2OzqJS+iXUvxTsSeq56OhIkkyN8u7SLJIgG
Nq795GOPaFRaVw+Om0SUToOeuYuvSnaijAR54m//ialLsqzdx2jXOT07Ne7pUQng
lXEeEGHiGo9U5oj621lkV6QyzTRbkK3OiJNQUOJrqafFVTcFJMeIAyMXqh+48D09
aJBIxKf0akMwMim10ZaNiMCEbbigh+LyXiOieQRVi+9z/Luu5Bxc3O+/9680IKMV
3qrrOHE3jb9GtlFm501izn+TLrG4Jr4twjNBBNMOdDmTD02xRL9LjZh2BoKdjOdx
XPwa3N2tlblxtkk3mLnyQ8EAKcsq7DVrsUNt2fED65jY387pS/xtG9cfqlGujlqZ
IId2+LCXBFgF7hOxYI5ZJnZAIxTDksR3VI+6/y+INYcFxpHpB9Mw+7epnhj7cRrR
9CQ9omZ1rfQ1GNpQg3eRKWPnkMIMSGDmUlD6vEmM06LEBhRAEao9rA0NB4VSJrYo
mnUn1ytpA3jlbUEzs0eCUEkKcmpA13b7xzMz1X5A0iYqcMRXSpC7HwlOAazydJ2D
zzsWT8RLdzqpdSsQduZLntthDe3cAShM4tKem9CGCDsfjplOjBrZiByzhtKIX71X
cW2AS/BrBgrFiwutBG4AsrRm6F6zosBJ47c5NzcHyscozCo/pNdEe2UDWRobN+rl
W3J555KwScbpJAsh+gcIP8x+L22omP2XcvruBNT0lymNYr7oVy55ncb8KAdKmJrX
WppC0N5WJ5LrffGSicDMVHg6kzvgrGEsNde0J9owB3RLVodg1F6L4SB8DrSXdKdT
LXC7ofmNhajzG2c33KqzJcH5uOvZBxYVczCrEXDdKDPTcCdfned188E9WfTWEmyE
CEF/CYGZbmYDy2j9Pzn4nL0kNOFs8/TPZVQq6bp1HpdYc+gFE6D4VTDI9KspeonB
SVU8V+/wVps6Jn63OVRhl6lMc/w8JWt8DLvtFj+smjCoAjby/42TuvYiBN4UFWpM
uq4kMQP1RgyL0b3mQ1eyPf31BE8CW8+m3RB5ypeob08mMrODi02FKTZawKZ+0rX4
sdtwPNjDb8vMEZ5e7T8fRt+SwnM5bUQ/Tzb6Dtg150T5v+vcY1rJyxsRJWsLKBe4
ExlTcf0jL3CBa1JkS1V8JUIukJ+896n8AmNIM6PNYnTPRUt0uJWnzimuRH4EH9oo
vqmdBMxnE7Y3pldYF18O+BPaJl3Ui+p2Ck0JQbVAM+o9f4cPm6HvtoNz+l0BzPj6
p9b1u6gnq+9WP5gaLiV616HuyDEyHPJXeq890aob3MrAw3z1Ix58OTIQ/cMUcJla
gNHI+/Xyp/TXEQgWP2Fk58sNNyD4C6B1kGIXuwwMkLL6QPm2sN/naMOZpSZuht0S
RT795pOlPQDe6RKJKo9KJFchNIiR5JtxuUPwb/Q3mx/EJxQZ129dtQGA/QQzQSa9
wCHJ2k+97EZT7/0mUb8zzfWU3LFVeEjweRztRRh7637FVSDH18nXWk6hzv4Bn8LC
aP89aKatBVDMk7vANWskaYjGRhYGJJ/1pBLDhziYoTU4or0T6o/J0RLZIUGLekgU
thUsu29r4OoZJlbExKNcMHEmD8g9sg2zIPDGxSzE4QUHmFK7vAqizWQi60InNgNi
67LhX/KlDodCZhBEQ0ckEPtdieY4BxJ4qjaUbcdX6/jLBtvMjj1QsA/UCSeIMrOW
KUjV/MIYtoMcDk8wZhVsqSfA84y8s1kt3IN53X7Z4AysdOJi0KOGX8GvGXEZPzTU
HFSoaL9uCXMR/+qJqr24xsUeizg9WVAWGtJyVwhpqolFuGyJde1a28RcqYK4GFMb
eJd0HgQclQDRlpRLDWwG2K5Gi2D6DRHjfn8DBJCX1IWHp3JalnK3mi6zS/YK3eYn
KkoLhdDV9kqSCPEGtIa5bUmxQMvp4PBgEPImVkV67IVT525VFUhBqU3VSBgzgXmY
PTC38nsw+Tdbj8Dg3wGGTGU7Ia2gxS6/+P6z8RGZQbRN6CB9U6Xom/VjDyzeJZoE
ZB9A64TV4hQq7uA8/+3qyss82L2RdQKIDlTmWgzBjQtuQz9weSDukMvnNBFVw7yB
ZJFanIBNTFnZANe6Sy8wmo8Br+qBu6qI3KyuXYgcyy/TdIfFJ2oCkZZPL7JWLTgH
7a2+0dY6gTleDIRO9xt1S6eap9/tUkWxNL79cm0tyh6odCqQrqBk2Bi8/HOVDK1L
kKBSYjHQzayvVHJ8VAipe9Fcz1Llb5ppRih0uvYzuwkgwH6Jefl8rs9suViYo6DK
tiKwEQ8OYTuMPMH3QvgVVgfDNRNSnyxUw+xVV0RtansX12NmBzjb4+R69ed8JcVO
Ycnp5tSBTB4b5V6uSUFJgsDwJG+uhUUzrNMzTCivzdhEvpl/w418x+Q21/gOFDHP
awnJxEqEFP6fb42fofCj7gPjGJd/XfSc5BEdSK0PIE6ftllghql/B7fYx0h//vBn
fGVk1kGYJGn4+q6rPN3w4wSYKttkI0gXcAU6XbEL8qrwwyPkm+fPEpxP5uckGo5m
PUtwgfaBhSVGurN7ALHJKCSssDuGgQVmbq1l+EQ+18whKHgJE+yZX3MsXo8gbSzI
mASthFIkr5n+wefIFB76fP6ESi2puxUVfzmgn/CtS+aAVJunpd5etMqa7Co2v7OS
54m5hsQ1vXZ071GN4I/e6d/3I6s4/X/A6IrwvO8Yu0AE6B4S6kupFKSHsTz+V0tw
KTRs4j3OSeL0KMwvR+BQKYpQb67DAb9x6xKnJ+4UyT3y+r5xS3zxesNh7YNLnsLh
DTwgn7ftfCfP3EMEhGg+RSD09kH8nBahNR5/Iz5IbNWeHj9pWxxwSbqpY71JnLxI
B9CgDE45LwXKB8yzJ5ig0NBkzBXF7jGTHO9q03asJDue/V6G/P8PF//fTbgWwO1t
FC6PxRXadmnSpA+WI+xqAtiGU+8Bor5U7+k8hkhyn25k/aYL4wS8TIc7se3yJD+J
6zXCdC6hddpnsJ6QA5FzDertBW24uMqlREb+qEyPlId8eChfWCIxHr7y01fDb7rm
XIOXOxyx7/8Vr4/DWXQq1BXtlnwsXHJuNcck5KRG1Ylg6+6iMFBmSIPW+iLB4GY1
F9emaOdyqL3Z7mBvNwjqDuNHWK05CTUZyEJytH4yfLKREqmjdA5u24F7h3Uxor17
Ge5+K7wtwtljyTknsJjWFcuRmefpJ0+37sGolasXxozxKFOM1lYvt2tUToid2MsG
ex+kiKnbNXmXoC2U7+Z5J42afi4iV3GbBAFxnuaJYDP40Kt8dZ6sgNeEMtBXlSNb
6yu9jJHnDfnK2vlzJNdHtCVlP+stU2Tx39n7QTacHTON1+wuw0buB9el8k7pXN59
l9TFCyGc+EhAdVqjq8bQEZCMgOkjURsbvEvfPARNYHOeBE9jHxH0IUZ5EReUUI5k
3Uu3z46aVu+U+w9nT6HLvQ/5dq5sdV7r8+g1gKppJYsB9El91oQFbqJEhHs7xjbr
Ua3ATRBYxoXoZ4nkG3y2TbSfZ7Cl9F5Mv58PUuurfoJVpk9HFYYl4/HZMtNGeCBR
XgxWI04r1LDmR/rOzfzQXLcCXA2JH68VxrP+HXzS6G/QE8uXV3f6WtiT9JRzpDgw
UhEAWG+fl4TeWSbQ5WTr1vNrr9bWbEom0T9pZuM4LlWH4I2ShIV2VrEoQicLvyi0
V3fNYmAwnRmADdG8HqYkld8xgqrdOC294RC0kZpNXetuKCE+y1wM3Pg/ptbVfB4M
CDUfkjjPGZNqW0jHV1YOfq1F+lMiaGpfHvzxn7ErhkWZwystcU65Nvikbq+hex//
jLeE2hJGuOAsjVtERp/+5VkIlvPxKD0zqxtz8q+j0Qrmjfee+AErSL5+SIwf1yMv
OGct9hbsWuO9S3xjwsy/DWE6DoWZfe4PLCNJETa5A8ue4TiBUa6BlmN335Tpcoyj
5xIWgBsL9dunYQYGOneuPALTJGHGe/BOYoM7pTUCH65uykEdlAirM7XSvrAm3OFa
aMI7tBmneR0OZ09zasAv1QouGUrg8KBFaPwGQUeu85Rtd3vm8bTUHHTc2bcEpzXn
QvxmzwcfeLvI1DLHNwGKUkWs9hZideRdO4kQ1UDtNH0E35JCgTtD+/+GnPX94liN
0sLxk3vNsSiWJwENuBfv0aPpLy7eSVAVGLZ0f5XG4F9osnB9esqDrqofivXJqAK5
y48sxLPIAMG/r9BmUlRynypWqen4tWgvQLOah/Htc9FOO/dDJF2ln0/C6iWOZTps
BGeULvMDcxBjFTHyRPIu7I9wcR5RXQcUTNgc+Kt9aTwE8JNvlPmGJeu1+w672eQY
3Zb7Ion23FtWkSQKTdY2J6zSZ9EUmzM6FYlMyBrIMfXMfAHUZYpYPdCHsIgbLBnH
hxOnbv79Ms6tlLDCPtX0E9WRWY++z4V+OnjxRkdnuDYVjC4RzlgVF5qT2eEfCo3Y
jy6Szg+28J5VZ4oHcL0CstQ3qqy63JWZAg+sqUixQ91LveFqh8o4263M+lBTcojq
cqvMjto8HRBbdh0FMDCfAAwyD/DgQXcS/2G94r7HRZXRIYlWAmUcw5G0JFX9ZFee
UuocRgYVvnQsKJFsZ/54ceQ9o9GXf54YeBho+0BOZM/cGBA2IRsXmDY7mqKjJ5Pl
0gg8tnSkGXa36E2+eWebPL7T9MJ5EWh5doo8gk9MkrWV9k5t+1WmDqIucZoNTCoI
Av9BFyi7pbFukgiWKTRefRQqgokV5YaRpUZ8E22JzeHPeivJaHBns8Bz2VLw1p1Z
1YF7MzEPtF27Cp5qPAv14XpjOt1SCoNJme/gJTYdjjeyf/v9lTNpvQ+BByQGtJyO
XWPug/yqMyuhVUgPG3zM8JCYJ+oZeAlDG5TNgGHBQWkGkgjYF9PQztLvGYTCMe7s
yTM7gK2Zqq0ndfCUnqjgu13glcnJLsU4ExJpS9YaV6n1wTMXFQybyVlz/B61+JHJ
ReS/IqTHGeD83UlyvjzkK7RaLzSHh44zmbgAKdOO9KDpECnqqUx2mqeeU6okXY04
f9ZlS7wA1/hYEmclG2Ju584zpl5suPD1M/uz57Ni8zCSe+SNJsrnr/xqO+D19g9w
A02Pa/02OYMM2ICqbvYL/A4v0dR2gnfP/fYFwQ2H3T27a1fXDAC76JrpqvpSNX2d
aVExQWVBadf6yTaZLmTPgL1SWKVt1QC+O3WUS5o4lO0CnUgHn7PSoFc1oZLQyEbp
lkK00SRreSLOzxymg1fZLEotWQcwiy7s27PXxlUyokNMw6yvpseViPg7GPIaLmEb
1Zkz66c1RMU92WXvlfmqYZkhmICH7GTfCe1uIUCa9cMDVQQ7q4g8+WrbokPVN48J
xYd/Re/gMDGbUzZ68YklAtMV6gnG6J7FeFP4OS+nZNdIdJTiGoeqAjezDTBCY+g5
JZQOQzZ7hBxnRSCHl2fKFyHIsWPta5GrolEoEWTturfzxkhulLGvlVnnn3QiFMIV
SnndohtMzZ0VB5v7i88ZfgulC07qhwh/9wJUsZK7Zq+tH20lNkejMB4wsQ7Ez0Fn
IIJ2zem30c5BWvIepfOUaWeDxaEs7YhDOYU10wha8ayQs/b4jw7N6YHKi0/SCZ9Q
qUaNLS2fU7JiOYADtZ1c4MghpeptCjiOTp5yNr7gnsBzV/IgSSPQoWBLjkbxHd+r
xmy09bLoguIqlU1rWp5iS6SOribfdUxEU4xcoaMkbL59GzfIN35UhTls0Ehc+odd
G7NFQLOAUkdiZzE/NnyLJvK7sdHYXrYTgMj+5AaOgpzhiq+yzWNWWbnIRdILxxju
JtY7pztWhB0bXufRJZlK5AQZhrq1mX1llQLowWa2N4KEWOkOPQQmQSPicoguBSG7
bP0YrTyXrpjxFY6fT59G08r81gmzHBGQGt5d4KJTMy/ZuQlFkQ28YJ4lassdVaHf
ai/BMw+ptuTGwHfDMNO4xlDIAlP8/QaDqm4Wen78GuWhfarw710vGyQFp3Y29HOO
O5Aq0e/MbPOgiSVrBVSziKfcE3hcxKfvO7AuGga0QS264vIK7iT1lPZs4lxFhaMv
2xuxmjGGGk8xBUl++QP5ELltRETL6CqczyvzvAWFbgLGjyYIxxSsHYTEQeNxQmPe
Ikle1TjhHIjxCa3+PxOQ+Hm2/bmXV09OyJrLWLgP0XhsPJjzF4MzajW/dFKYspzP
Q1Mf+FbH/YkDXVuc6wWCnM3j5kFE6hJGbuCoz+IaCoWRKabYkh26A9s3bPqcer6s
idui5kwmmaUSUWOnla4N2LNCGRGrUEMABIxwpAaFpdl7Jl5jXm6MsDh0ZbOapM15
66QcJY5duPXbOLKx85HKAGV7v6uX9bLlNffRgABSV7dOBIa6MX9gOSVgIA0pN/oH
2rbOcoOTwkqiU7Cf9QIbBxCD/t3rbVUpQ4PHCpoDmfCntdTcOJXi8fJnldPiseCa
+ony3+x4BST+ltzHDReVy3bLNLOP3gufKxxiQ3TOpULZZuVZzEJaQNS2FBM9T61l
xlWe10LWLAH8xP5bnuRjPjNvG+WOK5VbU79aRNEqhIG7mRZ2YXBDnODjcXS5mFgM
3F9g3Z6yE+XAu6kvZts5w50yRLvzBZJvcnFhHOSru7Xc8jcwnGu9JKeudCGiF0o2
GB2qPmSGKiW0tVV1fVqHjp00GoktQXmT1/AtwX774TD5WykbFfYWBH1EROQOmBxI
kiuz6/HkWnlkLOKK5nPnWpA65rgFlOmZrfLDPx2BdNQmB3wyofX5E7Q8f4c4I3YP
z9dH3SddEzISpCLZzFHykP0Au3+k50Goq8/xd2bJnz6Uw6BFTg39gpB4rojewyAB
OGJAy53meLN5kYD5B5CKSpLGqNDDamlaxpxuUjqqzfMaggfAvFnmv8oln7MfzqVN
7qzzrdZsDTQNNCRv8mvcF19tyEJahzyWuEWZdIr/gSsP36z6slMNo759rut8F/e/
WzGr1mR+VAcSQUUb4kGB3NP2Iz9SU4nRsLT8Lm3mggOIbafW8UZV/jb4sq2wFRK0
H2xbcu5pmJFzHLBOX2vJNh0w5ZCDzx1XVG5hSW4OdACOUf4jB0qCm2Jcvl7KNQC1
wOSjjtx7nLm/O252HLm5R1cQWtW8pZP4nxBFtYUE2Ssx7gdAGCFPVz2FOOTRDOTk
R2IxFDNpKg2ENTiDmHSm2B6rhlFvRkQEo8nkc9xOapG7Xw7Qr0ijxBdhtfH6pp9f
059zNslzFP38bSbWuefnQm8Tg4LkwgehV243VEgkvZ+7bjBi3l23zQ9BNhmR5g/w
ljBc3tilVpmqZBf4vRaafZUXmb6Yw3B8Jl1U6/6ae5UM3xmdxcd5AkGM/v/+yZAz
Sc6nabw3cVq/qz8TK3poUtBBV7xIZcJpYiugjV3PX+zKfTYwOsZ20rCZgrSWbz6p
gFIAEmzjMnLNe8T3B8Uvd/JJw0de7VE1IoPoX6iCD7YSqxyAQwS85dUWWCSvDFL6
Fsib6ZvNkPH0lsLXzpR6AxupR+G0vVDipD0UU1V/4VQbasZwlZ3P9RlO3XaotOjh
xRweCEvG5GzRol+43vV94HZlWvPDdn6lecWqf+d8wd5EVPbnFjSFxbHmS8NdZT48
3QlB+P7vO4073x/fdnZPfgSlgR+ztuAXhsU8mF64EZQPSIrOfw3ScJqI6GtIj780
DHdpz3LYQXvaLeq4XGS3uxtfx+2v4V+WTBOvFo2pXHpPbxVUzY0o54BLQtIOONkL
/nU8aZsgLQWHRaI7IPYInKdSYNohAmIZtKDm5ybpQL06jZV+0DLSnPxUdF1U+EDP
pnXtQWyqcQEx4Fk0V80MDMcJOhn2LMnb6mczu64na1PjgEa2cnTp/UIwOesdqvs2
WAgI/ld2xUrPP1KbSU3iT3lljyedxurmcyFT/wPbPEzg59ckZWu9/q0nwghdjlir
PSBavXMF93alNvCdXQiVHnTB17n3L12OOAzJqfus9IfALzQPknIiiaSDCzjte1io
n/cbp5OOsEhTZdIB0rnHsoMios1h+U8mL611ulpqiOp43hxHwAKFlZlc3yDHigHT
dM3sfjvMTgJXIdJLtinWYmSjEY7wPuf663ReevqhiHfFTRwgREwu65jtplQL7cdw
gWHBePy89CoxN6YdrOBiMj/EMMAzFBb6T6MNxCy9iH4RL6sp05viME/H01PBZswM
WVCCAxvmZow1RP3oOv7wFmc6lJgbEFRmV7ys0zsGkXcQSJc9+To8ZH7mpIZ2uU88
rCykKYJTSWNBVO8TlWhnY7qTW5ZHjotvfY37LaPxFBxQi836Uy6h4mwP9Srkg3kZ
49WkKXkfV7xv/czaNnJ8skjCp1SWUvZYjE6seQ75mK5wIOz2iW3OufCF+w6Ui6tK
qGTQ1tFiY66Tt9fnoOwRC8TxitaNyzlA3luRfk87GtXaF4xEbpHxllZLep4qLEpE
Jx3foNVEYEZNH0L2Vr4fT6CSdwVmsdV7MFYxXUwXdNqe/fl6MVvppvoekgfhan4m
nJZCDTRF/FQ0QC8XURHgxfXUFY2XtIJUbsYgRz0GVTz72a6MxNhDXJjkpaQqTE07
8VNQ+MC1Dn3ZublVROYgVJnnU8G1cYAq2nV8x7hIObXXGMISgUazlBZr/miLl2so
uS9OnJqAaek4REVeKnkpHdRu3NpHvN6gfmk2LN6AcrPBCmbvHAVoElSuMvpP2Qlu
Ghp/PWBJqSdime6sRn5RCv80YlHn7qZ7YPCBvt/oMCiv5lXIBkA84LpC4bSMsF4c
IWh2kbLi5Rn7AkRh/rkOtpLYKKKww+r5+hVtzSl1VJpTUnU2H+IpWuaOH96DNWdw
UcxWpfmUTHQ3D/5Lqrq3CAEqmWy7epJlTq9WQ+tT20VXfaGy0rEc4kAYVnl2OxCq
7XQ/QRhF4U8Z2UnFw4XaRSjvPWd5zP52v9jP6XeuiiRhAbAUFNkhiSluQSaUV/Y6
7lRYgKHS870XYnooKbPV0D4nTGoNZAGPNkDOs8xtIqS6mfSSl9cKq9EjxBr05rz7
Wn9sUzN3La1KtV7yoYx2RebRNg3PxTzepg07CnJ+rUKMw069R72m34Xm29cyg/UT
1ZxBZjm+y3mpNkLP+nh6dOvQTuxr3M4cwsQpygR3Jj6l4eLJ8+GiLQnzt8Yy/1tX
UtN8IBE89+qygoFaUYtPTiSEeFbz5uP4LIOFAwCR9YOb8bZASGYBqe3Qq1w4w4pU
WJfl8eJX0ru/RY0QRXyJEKlsDDMKdJAMDggoiC6ZbV/UTbK1vlLzZYkDOCF27V+8
lGb7qpXbN5fyj4ako5DzV5gyXoX8QHe3b4all3ZIu/0OZvWQT0zVfjm2HItL8Zv2
YhoNcwJgk52KUVGu07/msCdzikNVbBQJopopM/NDRvFEGxBNe8na3riMhThfm45r
QuR1hh9JqyJ4g36HHuYuovunuOUaNJy6v3gKZBmKK3qzemAl4I70I4PsSWGfRoTH
2jhdgZFcf1vJpDJ977UBgA66DkgS5eFmdk9BymRMjtj7jU4ArPGDVOcVhrHpXw2k
YUgI5S/bMopFkwhZMKOmOsDYS/EIL4FoIAAeIT9e4yhdqlja9IDEVWvu2bAEb/wY
i1TJG98FOdu8OI3JYMXSnkrLbQFfK5tmUSINIVZh2EB125HTLvDAT2tRbJ5CbGhD
6HiCCLonuVnL+8yL5YXGvBAkCqmCUJOBMboyibC/jpOKTsz8NC7clqWRY8c9Ffos
/t0wdfr707GbRGnUcj3JEeVK5erVqoOJfQHpU7s1lYrW6jPb6B25TE8fQsGRHQQr
odnnr9Vfv/7hQMsH8W5xfcsH1BhtY9wlZJlVa9FTL1+aUAHeC4ZwWT5ZoIi1Qbgv
MhyfkaWIi/YDtElsYu1ndzzaU69+OcQs6U/matBPc/4guOmk4G8IRs+3lNyZ/C3V
BhH4HzEtxvJ+5Y5YCXLtRrPJcobj2gWv8g37B32VU/HcE37ZWef0t3p8/4Bi5Jcz
Q/JfdxFZaavTRAy0WkU/LqmY5RKNUqpugz5gPloQgcJJfMpW4/0pyglRWZVejIVz
mbsFOKCty4Fp3NlEOPoeVNiK1yVRtFCGnhvP746HMOXlvDTyqmUhGYdyX6ngGdLN
UBkgd0XgSgBz0E3OHtWMIRjsbOFDQwcY2gqoTNpF81ozQmaqYLnoLFL2IwlflJqW
e5Cs4PyY5B4DN55YDvWhSxAC853XY/cGFTBM5ShotKjYaSoGpZcAU22u88UfsN39
Zr7WDBtQfBMoRgIfYQfRq7wS7AP3+LueQ1nComGt1UpzCRb0BkdQANIt3Laq0aPo
kr/erMZBqHctG2G5WDBOL6b9spOcsy9QCB0fKmWEdgx2FMARNd20TE4qhKv2vozJ
BzfsFaH6YcIduugqGpkTb8F/OFoQTjdPwGgPdSmu7P45miDt8jTcvmWEsvqsm33c
ediZW7jo1A1FK7C+sBWoOjQfiSygIZvNLyNJkUHAgGld/cycL/Gxvn/Jr9qqH/4v
DC4zwdl81kOdlIOO5Hs0B3wkZjZEFft3+fODHGxFNpBKk+h454csBmR0vjT6oOGk
w/8nEfTnT8sGb4rJy+h7z075b7MSQfwKtYGi8OxpWkafSq1RQwnZqAbUl8QIvisH
emVfieBsBlhfuP+e/k5lsaLWLjQQ6V0vcCVjhQOtZrMGwAMMmymF7CW+6XlenTl/
ARmJJIqnE0RDdpWPwgx0sd4WXxtfE4gzFYpskx1mGh8RGsBIsLaaj4bwn8dn6qLj
5AgJs3BBt7meof8UR0EceS5K87ngzU9A2lInaXDohfUPP3xEv7+0LW5FGSDeXig4
+C+Jg8On53nkXmvDIPQ1wS6sjKzB9IiuaXVYIp7mSrYov5TWopZFoREILtshJBSI
7+6+Q3KDe9m8RKhV8oYPOF7pJghHCRBXBIP71BpVo9MkN6t5UGDHJ8n07kBI7+33
Z96shV2LlM1rGKKKLCei7NjkHZiEfMscOlnBJnxr5y4vLmCLU4QZOmIYa61GWaQZ
f6nK18waMzu9qSH8bCcCgxTaq4R8ESWFIBvd+o9gNCPwSvZG1j4GXcnHTs6C9ZAK
FgpgOFUWQ7wM4F98WlAY71/NH/XXWi+TdCwV0yqw6tY0BaNXqrSa6NpzaK8bu2Om
LTOUmyrbHA9+H+fCLQ4z3kCBAru2IRRDhrB0WEFJ3sl0CmmyzkCKvThwFv6hzJhH
PhZWKxSSgjKRS1S9elQauuwVsk+xB4Xk1AL8nv3wVb0BQfVvyjl7WAUsGGHVMiQF
1gD26QKyCKiICaiGRAbFEUnBBvVnLBwuVkSWGaUaD8cowiAVVWjm+oaw9yxacQIJ
IJdQSZjJ5R9QMGUinMRSlI5N3pd6bOxN7ztwd4cLlXScEo+U4Mfrd4s90l917fF2
EI85QMo0gcGTjA7Qe9CwOxJEoSpC4OBDQHl20NiAmruplUAILXFqc5n6bnhAXl3o
biFrtr71vvIF65ZW3sqF8c8XeZS2EPrIgC/IRdQfv+c9TvldeCy3xRuibae+EKlo
tFChHp6OAEIKeXBkfVJl90r/1aghdtNa5NueT1lEFU0h8gNApsZcwoUbjbQLSSKr
3It4lcPlzVGWUBHnPx2EHHcbQgmCz95PLEEHpTvpEtbkJ4JMMyn71MrAzC5VLpBw
J2A2/Uu6B3rzF2J/2PEX6doexzrpxXuYGTo3GyyJuPlGR5cfOheIhytLUBqDPoO1
v6p98/Wq8K/b8mGXh+6bOEwN3SvGQhw3oeWPI3BqRFeL3EG1PxLZYpDbSXLO1/ib
TXazmbA5ynDpK6yG9fSEQ34lCZ7jh9doe7SkeFdxMCGBrWYl9L+kMi5yAm/NJHbE
CvhDF/nALwungTZMIs0iwPQ4L5Mo+qdhe+ABNKOOd6yVMYbBnPouc8wdvbIfJ9dm
orKLvFU0nTOAX97pJk31Z9iw1lAz2gH9lJ1lLz71k0XolRByKqmgPbOTb0Gcfi6R
9FfVNNUcN2ifZzSGP6sd9io3qdjbdqMOZppgOZkeizH4g7OpyMHkVxduaEY5YNId
qcMq01vYF3Zbf9s1diMKWuAGQWsf5DZHO5Vc2k0F1KnEWWmk9K8UjtfHkPBe9ayI
AfYbHFYgUxwBWNq7tuzjsNz5veMHIZiBidsHrhvGOnvi3sz0HmTrEKdYssNh+vUC
toqWN/QYgU57Tk/8+3e49iBB52/346hyK5MJRR4Kyx2d/6Hz0iRhILEh5eHNT66U
5rtQ+BR4EBxvj9755Jeo5aY41iyX6HVQdPx37GQzd2XwznD/hEJq0Py1ZkUdo8ul
6I2xjYamrt0ZvOjLknJo4PJk9plBDuDCHM/+JyLHlYlA66XdVLf51Mjr9RX8faX1
KvZG775h3Iodxs0d321D8L6g1Qk5deC3+9Q5k4ji3lkkOEZsJm8YHQkW5y3euUpS
Eyh8AJfHc1Gvj6/8k5ThbYHMeFlyd0OQ0tlGrt+6QUgDFB/Nf79kajkR8TEhRfSh
4T2Hi+PB12p070gdY9KT34/Pz/I8ikuWDI/3aeNCHsl+c2mKBa9EbOS1xH388uFL
NQUEeg9oxHWO3fdfEB0G9lS7ce6+NfPgVlwA44P5Fl0f2fA675Ew+jv1drspuBZt
vdip6GyxzH7p2O3doV51v3mbVJV0UiaLYIRw9hpYzPPIdxgzoixYY3dLp62sAfOl
47+s6g1d3YrIE+TPmtNQQuaPbz1jlhkmPxvuvrLvJUB/d5WVzYiIz8xzQWYxKf1b
mAJv8UuD8WezLCOBND+57rDn9WJT/hfHokuJwTEI1XXg8MVJEY+mybqjnaK3y0pe
FvF2a4ESfxPh2pEO4980PbMt+X+uzaCST9QKrkrUBSsaQwoqJQWZ5k0kTDThhCxf
J17CZn/6houCoG6pueXd1JgjbLju+xPQEm/EyF8kf+PgssTV60oIHeuBxvmDd4qh
WNYvk74D5+F9IjrRsRorCgUVIkabUupjQCEGrtcHHBy2NPlzEcP+fLansPBh2+gH
I4YGiP2c9Jxp1Ug0qZG2smUQ2pkpSHrFCHsvYUuhCjuKwvPijIr0Y3tHjWL/Lxzn
iMGZ7T/WxsY3DFgLKNPQ1G0AqOowywxNnKBWAPxirbi/j89oMDaChOxGIiU1BH7b
dw7aj6c5PlPsrjfLHj4CGGZFdq661Hprm1WIrQ0V5t3ydhPIx6b6/C3LXckgw00g
sFNWee4gl/Vo+7xLXcyaYNT9FeX7itvT01qh4R5fTKyDrd8mcCor5318on0RDDtD
/DdJhmo07p64hWAmZdq1Y1bbRXbtpu/fIT14r2dHfPCBAXrbkiJtdDtIjtMtaFz+
J0ZV9zu39Hr9iF7hE2F96W748QK8wC8S7ao/PnbJLNpju9DE1WHSghrcNLzNefQn
Yqv4BDR+9Tu1Tj2zFuJVU6WYOj2XxkVzcdave9AsuyVowBvOqK4g2X3gw4rHilOA
nLF8wH7b5ppiJaqwhYUO8mVQUhaNKntM5Rydrv7cOVaV1x8vUW6XiUGpyPig5138
ImL45mr94++LquBLH/65Dkc/wXbMy4oNFfVVZSqbYqdvhcN9egoKIxK4c6pqduTR
Nmk9VDTEif2v9Am0RB2nIKyWpo+o7tKNTf66wXZ0/nUc5te2PhkGt/g4Lc4RS/Eb
4WqTgJgI2ppbIa99E4J2003TNNdqWNkkWGmkChBby/C9B4GVGOmrcpWcIeNUt4FE
AYQMbF774aTjrjoZuU6F9+EIGPZh6j1P9RqmWrsp/hRAL9Jpfqo8cXHerV+XOL3o
mg3ab0Gc6bhFZbz8R0rGyoLow713s65Ah+wxd0C117p4LQQLA7KsoNjLihfxVV8g
OqIZ87gnssC1ifn0jTwqCXDyCRGmljugMpwD9Tp/HTDoj+gL9K93teojeeYRjiQi
+xIXuXDjYVw4MDtMGKYCn4tfBlgEQzO8Ad4SI9EmDX/B1kvZpM7FOWR3FwagDYXc
QUmr6qugsKPTjtz7IqPmbsTU32gwRjXDo52tkHj87kPXL78aFolLi/Q44AmqXMJJ
xjIiFZTOL1yH5hWCIObw1nxgp508OmWexrkRweEq949lx8WBccvhUUDNNdkx6j1v
hMK3ooXCXBGaFZl13+wHCZlyqC2wKaTBleoD38sf+CrX/dmilcemf7WvSqiA404D
u1qPQBmD9/mxHEyFFQeYGaWCzm8brT7AgzPNPPiGj4A7iIWdK6HRtDF8BWseTTH/
gQ0+5TlcrKnhqVSL9+uEaQQpGVt34sVzy/63ICs5OMJVD3yPO90EAvrOCeYFERUF
caPEn0MKle/geXUpMfFBUNFHCZLJU1r516ILsW2D9pB5kq6ixA/ffyXlidZiXJnI
jhbY3d/b8XKcZ9MKqyYEIO97rUtUHfqsW0xd2ndQBs3Uz7AmnwCnyJW6doeHSrMm
+nP6+a00HU1SibbzNJoJEtbFLzssVnW5rvq41bp7+S0aafhLrHHMn9DVAB2hX2Ch
GQfpCwjZCAP2GlgYGTP4AABfHDvwjWFK0tBFgGMGFe4PS17xyGmkkNS2h4hZ0E8k
oOt8EH4DbvtX+yk71/I+Cx9bsT/bJRSNHcTDvuWs3Z/KYI3zzt7O9/vRp+DaHbc3
a/K2Qvqb8Sf3F5j9l5+bBSFRnWjWGvRYIAljOoeru7q9VYZUQIpvZivM8NQ3EmCB
xG0p1gSkXOJ8cjLKiNnWU/LY5GQeKxRxRscveOdy9X5CbUtpkTZITW0WZ1TcqXp4
ewn37KhI+rkkjpB3AONR9AVfyeF1YIMo0YoItPKlZ96G5Y5e6wBTx/qg9AaugIka
GBE82lyCfscNuBijaEdMFHogBv7lqAj+RMVWwGbmWBeJcIrif9ivnbwaqXt2BtSL
gCieqKoVWVr96PG8pPc5FCmHy3VyDhpVZiUEOBVYzINx/r69j4bZgi/LN05Fsg6u
ceDQA5HI58fHmJez62TxK9HdoLJguap2V3Oam2q0IdOm79obb8HME/SQLMVaWH62
juIdRfYs2WChORWuKmt2vEtuCiERYewerVjvpOILTgVK6hPZjYv2islJTtVOj1Aq
ZvaizJ0Z/RFhbVGvW8MhY5d677OK5HUms5I5oyRfvMu3vHpGhTGZ52+bcex49B9P
FrfriaqqFAcnd5D81sAsp4v3JJBY+2ANZMITji9JyNmDa2mxmf96Wdbwc21231L4
9S2DNsEqEPQ+vD9tpDUrXxyl+LOanuMsrxQcLPC1yyiwTcGH/pmkfmsEnUdLHjyr
5GU0MpofpR/p1qDRDzPiHMbA/WHA4Pif+MBeBq7k8yTPds37oKCiG1YFrCxU5po1
tq2Jmkaemq7m3DJrUmfQCIgX24extYIX6Odp3Bz9Byz9UGFbuq3cSl5zGHUwRKRp
RLkOrmHRvVstxav3S89kZJK31pYkRGyOqyLd6kcNi9++t/FJiYh6WqmEitaGHNbQ
pH5287+8DP1RiQZe6yAje6/XYGN1EA40yKds1Ws+LK/1GE1IE/1ed2CV9fcmda13
A8WSfFc39fKQiSzpIfnnQzhudxAO8jYr8gF5jY0K3W9tEBAjiSEOkfblzEBMJG5E
cB2bd/Is/IeqjD6vJX0S03ovbMQDevrQDNssVMU+mBt8d7id3H9SUHo9q+JTyi12
xPDgSWFMC+l2Q+erokOMY1DHNzy00MqN48J+4UyoKGrOmenv6Wojrg0fczNl1Gwg
YmCXaGXnB+TnalIJD4TmRtC2t9dL/czy8CBMYG3Joq/NvpJD+a5Xjds3+M/JqiOZ
lem9SuJ77cVRtauFqSlaUPVJi0YWFcFr5a0dRBn4RRPSuwZruWpq+1TFj1kxNNCL
tHvAC11iHtKOc39P9VLrd9vlRriYkG4tr+jqwFxs5UzAUgudMp8d7tAs7xhjVSr+
cacBhtTpLCYLGSMR45YNIW2/coXQvaJ3gPeRrtYAtU2hRFoNY9rkqwtu7umfhbQE
QdxIOEklYQxACkMPCVcB9GT9MzuwZhhuDBuCh/piDDJkS66/V/xGz4Pj6+3ll4mk
XmeC+rvzh7ydyQf4S2C3RuG3fJbwzDTQHY/y1T4TRbfqanuxA1VyPLX+cqOqY3qV
FYtnCUyqyGCr/3Vr4KCKrV0yjFlRR60bN/jUHrLGtjIhMxdQtI+U3wSovXsqm72M
lX2uy2v/6fnKdgIxsZEp/1Twv+cptS0lU5vMMHnOcAIkuRYEP211lfUogfE+8Rsj
FIE8NKmuqQQvD33AONdfBSG9O91HFoWqf8KAwo3S01S92ZyO/hFiddyX1S+l2LxF
/uAiFjRRBOa5vXW8Pnu/4RoDlRerokrE+YjN97VMRu9G52Wy8jq4T+i7UVPdYWq7
Vl49sInqWZjJxmbmNuGhZYC4tMkFZF4skX4VEwRTqcL4lG97LzCEhL10r3suoUY3
DHJEpO5vk61gtxfdwZ7e+TeamluOl6UQK4ls3F6KnQmN93a7s1PYu9or6J3Vhacv
e5ZAlxQ4/fMjQfUsGkeFvYUuPlCDg/eUN3mQ9PozSyVja/+h1/C3dLlu7vOzIc1I
zY0l5Qyvlw5KTE6DOsDPGtF52NtvcLEevoQveY4uMvt3w/AJ2LLIgkZgFuVsPrDD
v+MgYwvicwGAshXma1yE7GLjaw6bR37sLoU/HRkJtOQmDu+M4tOx11az87QHzt2G
dj1gpGDdHuusbPDFOani2vp8dZa2h1jX0jo7/s+tYE86+IXHw0HIeI0zh/ATw3zP
vHr+HmYUVTT8Cb+jBQqAkdLZQlhOJffxFGf+D4Hfy3q1vSuKxWFtx3TIJmVTBNwd
szyJLjbWIe6i+r8OYAB8rGL2GIqnmBzKl0aWMYSIWBPlOvR00F4AZQk6Po84Ia2r
Xr0mTQzM/d/7+bvL6whH1PufN8Ssqgl3lW7+scpsDgjnURXsEYaAI8XaPkZ+Ifrp
n43UqzAv2ia5CA7EDAMvQEYfVvANq+eTvJhUAMH1DdVNh426Z2FDUEWtcw8dfIaP
KC/qkkcGeeHjAf/jvyFOuiVdc1AEjdG+IMF/tzR9KtkKH8OJutaz+WG53hHHoTyL
v88rNPQXgMamCgfrmCgLTa3yZbOvlnIIAntNa/ti8jatdUt7INyBzD03xL5IcriM
cRIzS9c1dcg1SjrHvYs9auZjf1FhKh9u0LWVMqTvlukkaObNWp9Q7CMTb/2sbbor
dO3Qo3aI5tEaF6ydjV/HaK5KC2DyJo3rM7JvOwr7WGQzMx6tNQvTiKKBifyAYZ6S
0JbjWUC4WXjHWW87yQKMYOeAuaEYkjesSzI41LNRt87FPmi5qgPxZBILRSwAX3FU
AYkVslgt0zmAhDlAdYrjs/53Hh/psgUfCmwHdMGwQcnxx2/wF9sqHv5MGXryoX7b
0ccGGSJiBJb4LR5/O+gcNTwUhZfbKnpk7xRosxoQbEElI8lz4AjRgOSvZl8F7/8s
sDZe09Qw4HslJExr6sSRcJ0oyEY5BXXyuexIegszJx9N3Bd4zZ3XqL4ygGMHjWPO
uviiZQOdnm4fTfKKePc5Ns2ORsd6AY/Z7aPT5z3+0PggjYTsO2YlCD49x/+OLcuU
a9J8kegTMF0/feUsmOqNXyrXioJZJ33cuASPobF7DHJ6ofazMs3PWKo6Lmowdt4Y
WxTf5GMsHXi71h64dM9469VtTHeXbEBFBxD6VTU/3bl1RaH2nL7gDwD+l/RV/X/u
Oie2/v9MxcVyq9nUtGsOLeRiIF4n7ZGWrSTxUoD7sPKxN61TK/mi+dEyroxTrDR5
rdWz+UmXNDomE3pZUu+54wopbioEDvHjCtX3ehxe+0BH+YcPTMi0YZLuok7xhrgy
BBCbgihh2xL5UZE4kASHaNVzexwRvF8ZH/pfHglBcuE9MhQ1WwinynJDQ8MUrJiu
vk7zUxfseAhtXaZGrlPYpifW6Da1uteeT/px45Fi3qlKlXht4isdroVvrKQvmSlg
pand7Eo03I7br8SQ7BdRtlkpxQqjUVUgpR0FOqUxfFhDTjHRTay84sRpcMxLHEFi
lttBZf6ARSQthFts94Cfc5Ij2Tj6U+hQkEGvsBpRVfXfGmuNbYLzfILZtz0hWmQq
fdnN+C6scNmScbZ+sP0OlNUExBAHYPtGhbLAHNtEIS/OT4rlJin7Bxm8Z0ouoX1y
JZCFGEMAtwS+kI+EypcOUxO8EsAEi9LREnrlrBV0n6EiSRGbjNGSZKS1Jb0lpor2
tw8hxqZ+2TPOgaJtgxLoH1dZHqkSGJDxey9TRY4JTqjtjQTghBCfPyZg0usPObGI
AbnB+VW74txgypz2H53hYC7hCzuwADdmCHF4C2JZlSlvq1yrUDBnIKnmIaBLz09q
5jR26HuO1IAWRrdQplANA6Y0v6aTWFNkjaYOt2xUA1f4eiYi1fiDpx2qtWXvMgIa
yKUSC5CxDuiy1i1Vwa8zDF1yobQtbXK1t5cGglRc119nIV+X49GUtRh83s0gI0Mb
NPJVV2W4dWt6CWf2pGG2RX0Bfm8JATYdoAsS69wskTbAHuLt+EhIFjGIWoQYfsZ3
LUfGBwcEh11Vti/Zm1/dsqmhHWpEyPfFjzvkcoavxydvtMgRTRUZLK66gXXywa/9
Y0IzN2anpfaeDw0Hdg/DMX8+sqJie9/1Sdu344lfq+oe91v4QdKurwJhznDAutPS
AH4oPr0jQCLoo+TG5Vp1jJknQMw59VF7Rk0l329LkEAF/TqG++oyTEf6rR+kRcnD
9Zuw4CXK4uQM95/3RQmx73Pmqshw/VH4xOaAfCug8KR56UpNZ87C90jZXzn9rGyZ
MvcWjNOnHc85KQfWvYomv13lB7BIQcyThmouU+0Te182lIwlG+puYwtHCWIcrHMD
1yWrShpC0xuRq23Q3+OBZ1Dz7G9i6PR2hiAfBiptbjcJcnugpbUQDcTViY2J3MKo
mcH0cVAcoxlikuWAbV7uOTPlgjniggcXAY+ieI2X8/tGCsL4rxgBcwGOk1b09uCV
5uiuXHCTp3F6Um3TOCd33fvMW9oEE8+QQXqLn27ZJHU6Bg+nyRaOLDrzz3sOMO+d
Kgmihp6YHRSo9ImkvvDX0LKy23iM+F0pGNGsV6az1eqOzBUvy4WTqycc7kXKSU/K
Eanfyn6Gut8Rh6W+IHttXKZa8auab9RayXkFlnirYvIkfYxzZaq3nQMBuitwz2hl
itD0k33kxezkYGiLKKC4j6AujBt+IglaAqk8p8ThsKJyuKTzd1bm2co50B2zzkvG
ePNYl72xHkFCrSex5sxcoHrSnMw8wORfxD/im2RablhJd2o+o1Nnsd4W5BNVeYwn
Fq5NW10E3DtBU4bUHI8S+ETxgAjH1wSVUgJqE5ax41SMRnW9KQwfruLN8NZG9LHY
jCabHzdJyVOC1AQdB0dFvuAYz+xgJsFu5PT4mJQRoUvLRWp7JECEdUFgHSowUZKQ
KQCDhwm/xwYnct55d63Y+nWLXVSNv5Oi+HQ8AmaBuj4FAULE9bVUc8VrXlof2zQu
EAAWQRGX6UA3E12v2d3cEeoRZjXMEXa5CuSlL1D5mriY9nYb48Hh5rJgqmx6H+CS
hvZ44wgKyfpqJyR/FUDkLHeGaFrjCXzmpKO79huw+vqLOwGp6KBk6M5kqPkqt5Ix
ahUsAZFgzHsKFbvW78YSMdQiGpn4WK4IwGM1ysqbM0VhFnI8tPIJjfusq2ykA5WB
9rOuG72vNYThzb3gRpLsjQkvLz4C0ThYH9K4he+r/fcofXvPWuCUtJiRwppy5zIC
HO+OJL0af2/pNxUMsZTan36jMnc3bJCMzNboVuD5aD+me5LTgPY3Q8d9FH4wXX/p
9eU8h506hJsnZE8XEyvcCXS67j9VuIiP8myo13Dmwkk4ZCpovPRUeOkTA8/NUIs2
mdf6kJFPRa+76/jAd4nsjSpb5vvbkPJ0i3bGcixLAFmees0JmFBT+zaLwuSyfuiL
6nJ6G4ILdLp2HKFaVRG0I8OO3ygf/WFQZGq7YcvYYelb7LbHuyjqk2I7QLyZjwKd
efVft1y/QMXrqJJ2moEs109ra2cpnXxXmd1FVHJgM0HzT55HMSou99+a6PF3CBsT
qgEL/Fg9E1T+/6Hj+iRG3g0MreD3I6Nfv9/8y/hVyxdUOXxPo1+gtnGtDcsRz6nh
fJiG0rzGOuKjZIPIBmG0EOxQAcTFoZJTT8x5eRXdX0K4HSwhBUw0cOU5zlNb4upe
I87q1vPdlxT3NtNDMvERpEWtfpiPFBwWcZLwQZ/Y2sO26769wANX0sUwTgrl+vh3
quMHbSW5l8hV7KAjnD30LUDiFl9UDfSjvMvTNvWQdY+CtwayR1jCl9nBcQx+/Wn2
PMCivadRNpEj7PBgIx5rJQ8HZ+/Gr1i+NL3h07y6nZCezMlzFdmFjW1MU7OlcQm/
9WP52prtNQrBcyxZbe+r+yFL1Bf4AqZbvrJQO48NKuZUircWadytSH10byLfjT5w
fCVuYg8nrBipoyDIcWm+KX9a7vohYoPRwW6fQZmrAqmQwKbBBWMX6+tblAuj/q/3
N/jBhDtrYub9kkJQ8fby/e0PoI75mmVStcvrCHDcbl1d4lhsdCi2BIEI6vf2jyqu
eHpXz7fecqgNtHP0zcN87MA9Tuw3mvrKjY1x+mEwbtCnpLuB0jKLSKEZWUo+hiEL
oK1R43sSlmKIPfX2Ri3jGLxoYN15mf2DU070JFMbB8RelCOFltzJFzWCqvtsebke
hsvPWi3ARMRrjG4Igp6YUACg/DFjIbINhEg8R9WbglDMUzOGailbiHpB4Y9iujJM
crsf/PNSr9M+5kwonYI5r40VZo9W4wscZIjHy40qsHSnPzkKtK1d8aMUGoGmnM+E
Dxt+xQsGq4HY4YH70RgvYjiK500ozAnD0zhhvD+tTrVU5PJCXgxm1wBwsEm6c1n4
IrZh9w3FYOpoHhNbvkYHxwh7X3PqECZzRRv3NJMkTbFZ52WwS6BfZZslHHv8YYUA
7r2jlr8xP6oystJBHTH6g7YNXEbHdjc40U+/870dNEKAsO10KRlBDK8jd4XyIz3/
rNzol1TC0nFF9Y4caieIIfY/M9l1ddAWIOMIy31M8Gsqo0y42Cb756jHASAm0hw5
74GdB3IE2vtd67L72eYYL6R3dteNTTAl6oNqzg5kCy7J7FBbCwg61jnooxlOXy9U
pdiWRdIiv6QcnbXfel+TjuF2rgxPbHay1OGwqKoQUeY6NiGtOy5yLQ3YWwfi+tlN
zp73SG/DgUDQMjPVA/+WJP6v3oJd/ZQIupa+Non/ItXLuvgwnvTWjEfbxG+7LrAm
jRV0frp8DMjM08fHgTzCQO7zE2P9mpjM7iA8APUoX+I/OhXOLt5VFSQdyKNXFj8V
rO9ACUbnYI6RPuDkN0fq0ClgFsjManLjVs1DO958EGNcEZRoUbWSBmJ2GbA33efg
0Qi9afoMdC8cGROZFMtBRtdMQgLW73id+O4kKsIaBglpxxGGLDhG6VRaqs+kkF3z
0IRZRB3kSnuF3/6pISFOM0nyv/qa3r+mV56Lczuu9UFXrNov1+dE+2KwpnwUfxee
oFrGYeHKlwlueREQtKVe2G8oWcdtf/3Z9D9gLq2YYkRvrs6GCg2nDEo/zSdZflk0
qDwxHXMsEl47nqUowat/+QIw3X5LxDAu4lzVlY21gMj8OOjY606sZ5eMsIFNEn16
hx1lPrFe6FuDAwoWa6jdZ0BiLCgWtUHEiPA9zOVyOSKD96+K2wwEZb+MGQ849Dlm
knyiMAqzSQ9hF/J+eOoojGexrJg3lp2patzW3qYWByKQPh1Ou/JeFv6swfGnCfmA
VReWTTNTON7xWHRMnSktqQPcsde04GxSergTxT6XxayKQ59mOHQIoXKzz8Io1Ucl
wCP9VkqoPIXr/XQwCs69aWBwhvrzA2C2O5UmMhBQuqWGXJfjQPP24gXkSuBLvF3W
qTvU7D1ZyeWLi+C92qJN6D58GYwLYGDahqB+NoaW3209mBqGux+oR2qmq/xsyVCT
0RbPJeYgO820TdAtVRYABI/co/bH3R+kPb8/6hNSJsf5PxQeaVXdLGWDORKW3Xat
GlHdglbVatTLe9smhIRBboQTP3m411q0bNYcvLOstnFcO1Nn4d2Zsrvn0w3iE03T
Yr1aLKNFpPVHEoimJXrh8hBe8v2rYD5Y7PWA4V8XlQgdZPjVf8TRl2sn+BC7+Szk
YSls6JD90DvsZud3rV7ggkP+xNy77U5jlRUlmobUwq2i6Q1XXEH+rnjCmFy7TbxT
xFs3BgHHor7Zlb2upYs5/yy74mNv9sOnY9SiWLihlj9uQ5eIlC+Ifs0eRczw9MPy
gBxSqt0px456n1DavZH4S/6eO3U+9FV/9VnbhlEpoQSjelkjf2TLOQxhLddPNu44
/hlKNHGLCUNwrU4ADPDX0yAeky9IjqyXlD+PWxUugSmsNPjdugp225g6GVXRi5Zi
jxUZ2wI9boQvzg4hV8t5i/yqVR/3k6RcE93tXgcHX8JuONmtbkd12qWpiuc5+Jko
9A9uUT+9LBtXzPE8MsrcWkz6KfOERwVv5BM+c2Fli6H6P7v3ewkThGH8eVZGtsQm
XKw5Wl96ltYjhtCwSnd+HknFQ1RW6IPNTTpTmp73cLMMoVyua6ooll4ojNmmlSld
Cnx/EJaSIaR9UqFWmiwUi1kQIohQUB2Q47qaMXHZmzjS8DklrNytskbmiOpZ0u4+
CzsJfGtUNZhT1SZExZQeAXQaGSk4Tl73D376utB8mggb43MUiodSR9WKpY1utYmA
uCytLa45spHfLLWEr46kDuLU2nLOVvZ1B3HWX1l0hcxSieK2PJ3yoJPtupA/gsOH
4zByaUqu7hvddwTcQ05U/9v8HXcoVWblLmya7AD/3fen1TsVteMwZCdlV+v8SZbp
6UWQOdrktbW7YK5yMLzfGfzaM1F3MRJ38mBboWhNtZv1HyFeCgt8X5MwBV0w3bd3
LnLxTq9x7fQFXzuBqGSZU7zGrvPmoXfT6gDunQbG4m3rwzhoeYy4Iuwyol1jfFyC
TPD1044SbiNI++o3Do/gWeBCbjgP6qrb6VulVn+i/thWg5LAGKpUEPpR3IwqUxGG
f9rrrqTIVNot/tpaQQzxhY+ddJcgcBD29z331po3RS1PjUS+7kOTZy49LvSADPEj
9zXBNC+sGWNKwyiimWpN8DUGbaCdxjZIEjAkj3X6vTPHftSDavFCTa5+JTuoPPkH
r64dD0HvzXyfX3S9gzeQWcBzseoXjun53x092acodoFpBT2ZSehZ5QSo7R3dp8bE
pFglbAeO5Z19i885U34PnnXOi0+HInS0upeEbhM/ZAxqf+ERhn/LMNb4nqnihsdE
ijjA7vh3EET72WqKqGLZljOUR6PiUTGuu8BLjJRLsHqk/K0VOo3cz8iIkx+KR1Ft
mo9KGEDj+nD5yOhUfx2E1Er0TDI7+LY9yuVdfC1Hfr8JWq2u8jp6QJmzY+Xpt3RB
XF5exzshgXcUd74iFJQAe718/0B5eHbZzIQg0+jR2HZthRSd9T7J3V7B+XSIrIVN
yoFZf2sNJB7DRewYN9u7qzSipeGOr3pXUTCOjhjf6RTzH6rKflrWx8Rlc9mgrqSY
qvrnB0N0WFVG9m9fuq6oOc9xgkcq0HKorXZ6VQgTS1PLkbzazSnhmV69rPM4Pl3f
8BYx5SI6BwMqvs1GNCAYpbFvn3GE7tMO88u6RuVeHp8kSpOetl3M5D98/TeTABJA
B03In2Nbu8L9+FVnTbL4XtmooXzjl0Ozk6hmkIDbVRmfV6aCWCm3HjcNtp4k56hg
8BuFnfGPDTLr4eVWi3Zrx2GgEieae1JvxpvwTOt2PjzmAjRLlQZult2BOufwPj0t
0B8CgbefP1OVfZsFaXfp3pgJR6EuVv0SoPhiWm6VwgswNAPsoGjAYgNBTQqzZQWt
5Fpl6n6wWcwXiljl+x/YLAUy0mx7R/QuB9nhcBpQmXcmmivHJL57CXaQOqMk99Ip
DeO4r2KwA09/igj2/m3EEyFl/hMKA0zMEAwLysziXRSxNDBZmut5ykrM5hDJZ7CQ
7nx/gGZRiHaG0nugG0/azTLpYPEp4LKGbETT3HOpGPpDU6wua17WrLDIEady8RJx
Cf0ycVZo7O7V4NruuxVm+WJORn3Mp9poe19iiI5vp0FfhvyEMRi9GosG43/cPSIi
HpS4crKCJEh3/HeMPt0BmPOQYDpo59fb1pFypxnbVYqP0F4zVnr6UTcyiwCbjied
Bu/AzZClsc1wNM3ej3fMYPdULGTHy4LM/iHzLPIczNOWksrWgRscsFUFxcAjeBCm
B7p9snm5DUkVQre5AHBsf6i44aCowa2dT9fz7Zakg7Wvz90pRp/lJuIqEyWDpSYH
7fhtY24dUrhLiAlkQdB2Qr22EB4f5XB8rokg6H59KVqC34npV5iQeXozWJX52zBj
9XCeYi3OiBAtDmWhuP9JfONJvlixRsQo2Z/tJ/391Xg5XW+c1xTNztz2CNp/AQOL
eoRdMApflmwsVth1gKKPkLOaH/aQZA09Z2cYp9Ft0yJVIg42mu62V6UlBwIvZG67
cTKASB8eX1kocCaPJf4s/EVbYB45etHLxcUqqCVN7sRvp7niD7S1iJLk6vuCdpTJ
aFccb37wEV70dGZwQ46MIlVinUEfOiFcUTA2J+aqF1IZzRd5UML1bjcaYRmylCu5
B2iN43wR75d9lPuf4zMUlwNz15xEprfMR5BV82LbijkWwZczLC/4L5PkpYDtdTtH
wI1Rk+f4Nf5NXlM+brpRbG/kuqRIoEXn5zcJCkIPwTAdx01ZVMvyt0Y9d86+JFCZ
JQzRh9wl8rKbjzekDQnvMl9JQX15HmKhhEahPUQDxA42jBjODDUt43rXH1uThVT+
wWtHu7l7RI3WkAirhB24n+Dw0GbZZUJAJBUwAguqAb1sr2VMUOjskUFPJXDytA8X
vNOToBD52Cmb9MuXYGN+Vqh3aiqV/+6Lmj6+XjqjKKkSTIuy7uc+4Yxh7vPgqP2u
mf5ZjiG8/S7sM7wmFVKKxY1WrzvTrjogCFMIAfRwcSX3qF+kY92j191TWvzsbBXk
2HblmdARQ9RynW8TPeKE/07xCMAymu+xYYZm+kYOnf63eJNf/AsV8zxS9voG1n7P
OevRVfOfRoGu77cT1aa/7oxncPlQ5A9MLr7wCspKytgniNc6chMsa6t+FR9rQbFd
dFuEP9flSCpsl10DJbmviWAPjQjJxWqAkqbjeghhDyjp76Al6pKQF6DNSeSLHK+w
FDOuPRfEDvz/U6Xrw2hCiADm8CBx/1Y6TUbKmz+4e1k+k/97Djs7/JmUem0s4f9s
eAVTeVTDI1FTpjuT1cqyXD6dchGuLi4p+n1Kf760xQxucaGm1Tks8JgJXtgAsGlu
uKnHXW2oEglhN0iR8Fvmyi3kpNwPnMsir5JGGNvFmgYvRooqsg3xDnyKKhYR6uAf
9J5rY5vWA/OzPUIqYm9ckaSZRMNqQyfMJO9F88cGkb+0IQY1DDWSVqRJwE899rPr
ZqvNJTrT3+usdd4TFOs4YnSx82c7BQDcUEeKjaQNVt9DqzBmcXhDD1dBrTWVK9hn
o6t0PZFX7nXCYeIlXUXHsRBH3NMHDmDiiN3IUFT1E02t/qFS8ebcnzyUC0u3RIla
yKMjVpVY7msk7517Teb9zZpzJEoP7MEoQHF63HHsR06+sVcDolpyIB43OKxmltFD
Wh5EUIGWZtLIzKjlihsT+xiyNfs3L3IibY/U09Z9f+BilDhHI5LEKT5h2PBLbN+6
0HGmZihvfBh5CGWEVgh/gD8Q3Nzd+wdPKRXM4ZPb5jZ0DwX7CSTBiMKzKCCJDWdu
F3iFfnfs3iMqZ0wUoBkph2pCzBAsMvHtsYwngBNcidJJflPw0M9D3IZJ0Ta/pKJH
rRbA1U3S8r7Jy035gBMxsihV46FgddvvFQzOs9moAlaHy6mdikQPkgm7EPFue2Zk
wrHFohN3o8v0fZR56rE6BNilEhJ7nM4SzmpBcRv6eAehc5/gjrk3H8k3jQrMFEvO
/j94XvcmtRCbyXTdrSBklXBDYt++HRcsi8JAoaQY/Lqnu5FKmckBV+LfhLVhj3gC
F0fPubpWZ/5H52gsRja6VJumLybUNVAth8ZOp/hmTixJufiWdHhNoFm5pvgFGJwy
+4CtpL8teRwwe1ecR+LMAOwsi6cR4TTSxhb6O88JaZgTZaPIAnSIX9waE9kS5t0J
tQ0CbbEKHAGOQheV82A9ONKGpqERICCxMfHt3OeR8PAdOMfI8DNlbqGwxKtqV9kP
ZmKR2a0FhHhpakphgwd1otKLQ7atXZ4O8gYg4xnRkiHj3e+MLYl50vODTRl2Ohpf
YJ0JDBZ9mygZgE/A7h+nRWogiVNycQSUT5k6ZCHQRQxBnBLoGqonHGZYI+p2MlY5
mv71CgK1mEg+IwpxC26IGX/OMqx/L7+K5ADJrJa8ZEII5dPkpluDtMY4IInY7kRj
O8lBRCZPy5RMQm2Uz2rP4hlEqSiSOyNwUnYPnQSfZu4ZaDSZM0+8yXsItMhgWrLe
ISmSoNxLyGdCu7vA07SMhcYt48NhDKYXeOxqJ9UPAIPMmDjP4Wb5CYp2vxgvLqlU
/D0QcK82nvtmF9O/A5D/7772NOAbiGYC/F93yblaUMsOsMSjYH1KaGvxfApYAkz8
ZqCXVAbahfShtvOWv37W7nZ/GSWLnTzX2kXrHfoa/JGHxlmOkOqje39CUTbD1rSk
Rz46Tj5Hz+IbD1Lmp7Q19ZtIU9f/La+PALUEwPrGcqNzhF716DsRW40R5cnk4m/6
cQO/EKB8dD4j9mEsLGwfL89qUSgtfEPV8r/+1pnZ5U2BiR0VeLO9w3Y4ZOwgA3gO
N5MbnrOfUJ3yZ4mB9RrHWEywHxN0AuytEdT3hTPSyeuzdNiAyOTgX+TNX/9BXoT1
m0Va+X81IgaaSkBZZS0bQVJx+jO/id+PupBDMmKHcznESa7fmhjY2qS1YVdGOrP1
kHh3TQET4FY4jD9cgxxMwAoYm9E2fpnoy9f6mwX/cRmdhRz9BA1pcIIQcN6MzoIW
FZBcLF0shie1HdJf0OaRdRG240UEyfmLWLtA/lWBsBoQFuwvblinc1J9ZMi5PFf7
+r1JHX5E2hk90yf1bj4El6bRiLkj+i26d8h+id1vyuIxx/0cZhLs8QWDoWnY8nx0
cucwqtyDtt3m1/pCqL/aJ2IRZe3zshVJVIJk/7cSBuwfueMwi9ZKNd2Uh6uHG/4w
jTBsVtRxBOYwTYp58v04DZCpdxfTKtf8oKST6eN268zq+KT59/k4OYVoknREJpYm
fkL4DXLZZUSIKC3MaM/5roRS6dVcHlFOnP9aRhUtu/eiYYBYDxdKYDWawgkc75mw
SycspeTafKk+6JSv2SLOLUf3FhtQEFkpCd2PCb99/Rr9OZr2PZJ2i+fLb2lE+v61
0/t/EFee4yLWEec5vP3krVlpKY4NbwnBVBY6e2Tn/gmOSlz3xaUFtuki+ygkenvt
JiT+W0D1sB0YVm2DbPetoKLtjKY2yQI0RN7eYA6nMao6SBm2rA066prliFcuhI8K
LEbxfTxsa4rWInBcJRUwepkTmXMTZNESyeXKWvwzIYIdFxJQ+X7VzJFXyHmGK1zw
ZhGhcwDda3Eh2sAX3MKjaVT0vFtAgUeQep/jMoNOtrOOo1QEkuH0/RpYyFXDxzwf
Y4NWZNQH9M/ChOrIqjXMtZoo9/xufIcTRsUJfWqaYLODRYMHaYw+KbPdcfy/gzXL
IYFrMxyeNVZt4JbgURrwAVllua6hRm1FiHXYCY8EHB5r69Lr2RsdOMKKZsGGXEXY
IVL7EQ/fRk9V4xbaY2bJaMIF0IaQI/kXaeBOTtUDLpEvMZc9gVcBmNk/vRZHroYL
DG9G9tLtNxQZXgXYhTbq3SCM99FFHONTVyRVvhyLPUoEDPEI/+97WdLKzmriaG+g
+0KP89mdrntHxbad53D686HD4+dqvMBFhYmkVloVegDzX2r7iFYfJa6lKxODK5iW
IlBetybIbo3+60lFtbhOLNeqBFk1msE9lmIj/vnQHoYKYLgxcShdBIa6KfF1QTIr
LxXAlq4iBbMmFqGpagXdNURMGkR2SYLtHvSOU9V8Nt8qsx5Qayy15TT/5oUEt2FP
y7yzPjNFB7tX2yliS3nWTuHt183gbRDWiffUk2e0iJM3iJzoARjj62ACazWevR6J
5SXZ1whVYhT7nMvoVxThpaQuQOUZxgkNF/zLPzd/KC1HqyMH7o7B37shqvrxwKGm
5gLQ5yV06BQVp3wV+OW72VXoW3fG/YdUAKBul7/IAdkfJoW65fiLC3umRyl2KoDl
rTly67zeaA0ZFbR8JqeP/VU8GcIMwyzFsDYZjKIQ31w5lGeX4EDr33Hf5dRN1LrN
lpG8eV6AAygsTXCpbWVYwC3yPwlR+rEeSSIjmluZJs0XRGqjdi/RIFfUgwaHXywb
r7OMWE1iR0vQ7j4ZVBCSHux+0iMJlb1lqocmH0Z9hJFG04AFTrXGbxlpS0wmEI13
xfyOnagiGp/NtDemxG6QSHbypS9PYFjQh5WHYn1H8pIZPox4T4jl7WrugzSPRQlw
xP2rQrXn3wf9H9vjXiHgrDdmg/rZlpD0B18y8GyH39zd8FyV2vm1W7zeQrSrjjqs
lscqkcgTRGYokU1qaYgkXsQMaGFfKB+VZZOHKclrsFWWwF8csj9gIR4GwL8jTgja
W7jbMVSjgvDA+90UH9ka0sMfKmVBXV2WBJMXNt6ZqMhjNrxKIoeNQ4t72OcSjmrw
aHTmvyzVH8d5h8tqoqS0Q1VlFzdTNPuNHBLWdOOKefritATzoPCgWb3Ro2nOfGaI
O+ZEQMzMSU+rh/QMrGCJG2IUQKr8mkwTkg++LzD5T0/9A4uAjAT6tUOtJy2QG57z
2dj22NIwHef4/XjVtYU2kXb2P4X7ZvlLxWv1HBt4rGMUfeX0aMrmdP8QGfmCce8r
jTFViJQNkzLT/mkxqw2T3rQZCCCOLDkY9aSB4R64GHiIlfTXInfNY93ucvLiWIV0
SfSu2iAA9QLDzNQM/fZaNI7IuEYKsoTn0XSw3WkfGr2U50m677AEzthfelDYYDvB
kcV/ilpIX6ZFTpTW/WQMY5EtdnN11F3NkzDTQgKT6JzAKQX56vOviKAdaySgRlN/
8TFUG4SfrnvCqcPeUSEBlEUuMI+OQ6dbYaCBWzAdkou4+VgX/SeuNmwizhMPLTkQ
0eiqvVZiha2TInzTE9RPB4nK5uYtcEhmfWIt81U6tbfnlHxdPG4Tup4cG2LNB2so
8ZNJUR1LTMHpNoJC3fGSIB2oyMGNF77qimAbGCQgOnyu8orBPBZK1bOttJkqaDj5
ZKBrSf1SResYq6GmBfjnb0+jx7G+h56/l6I5bP4kYRpRgTW7WxO3H0zZQT5ldvS7
SUrqVZyW9+CI7xCder51HnDYVjheyN/IesoFeSYjmVa63rY+7Qm6vXv4eWMjuVCQ
UAs/UeVpeZW4q+uroaEptsysaFQxgpvIZDOnS/UWhToBcAS7zw3x/PzSOse1uTsH
1zP9/cjLbWB/BgwM8sde+7qtAJ1tCSQWWzb5ezeX3pexcUKg0ZUe0kXbbF1th1BH
arvOTsHnUwuLbj8Cc5iiytiYOa8L1vJfjv2hvY0oDFv6C9H6ZIVZbQfaylayRl9x
gab0/znrtJfR3Bacd8Dz6KTsK0dZYoIblFyjmFtVrxXcmCIokl0lKRI9m+HxFsos
eTMzTkLZaCb0LE0bwOFDRhNa63TQjSGAjmep4diEr6LHpEoKFBYVCeCUn1XC+eAY
Bl7BEiOi/GFQlJ0AOcxa0tNWbpX4mfawIYZeJ14Y9C5R7uZ4/4yNdVWcHdGaFjMc
ofPjveR3NGq0zA7Idks5y+hqwUtjH/Dvysji7mhgV+icr59FIW3VMwKiEG0QeIJ+
KJvc8AWbQSTqUfQeYpo7CHN69VHSjwMbUMknU8Zc03B8/BZXtibvkVa7l0CMB1R4
UtXcrsi86MDACjldFQ5RmCmT3oGZL9SrQLkN8AmEWeGACNEjnqb2kR2JHPyxdExB
Nju4KwU+/vRv7W8Xs55ZZSQVS4VxJ1AW3WbZUqRlKVELblGq1XqoioyWesm5J7q0
GlmUL0E4Wgl9ORg/BAq61Fu3nTlFaTsiWECzNMh44kBND2D1AxF1ZsRO4gtlk5cE
Mu84WSgkZRAGJf9cmouJHR3FiFYj9FCejIphGzPUvXEPhZ6rQYasM/cM5DL0Kwqj
gvfoGWx4uTFX5kpoaFJk380z9JXsc3+VrCeq2OeUOIE4EKgDq+bREb9zdQwHLIoO
jGzpWcS+Iwiq8rFaM6rRPOoiOpdkS0qKvq3+vjebJ9Su0KmPOBkwe3Ra533fSjyv
h4UTzqWJ01Fy3e/sUI9ZM2wtwzRwrI+eNlYZJ0VHZoU7ZeRXiTCLymQ0KxVKxeQR
GgJempngDORwziKktEsuxxj9yd3unV+sJ1jVMZKCBYPwcyskYQQNBdTy6vfhXUCB
k9Ph6J6k8UWa4jOy88HYLKHJc4ygnAj6rRuOZ7EBXYXjl282enrNrifCTBkSjaeX
HATKm0nNE/fLT0c/E7aibQuyNGWj3g+Xe+927JCkuZLYJOTnGO7dQXesfePVPKOs
VxePd0qnKX8d2bkS5W1S2hmsrSxEu10LDNCPtt/jZTWPjdVGiDrvPGMqOMZRxHXR
AZscOBlbUQVywhQuIer6oQyLwAh4w5o9+rMYDWoGbhiRfLHAIr4Ce7L0PDgTlmFn
lg+ZA0yymFzkWWBjbhiorCtlh93EizBYhEv3/lGRQku2Cz90sSVDD+w4IVP7Q8/u
LT6StcDN1VJ9GFDy+CsByZXqJnLlaVI0Cmmco0O82FunPyoF/CGSg0ZfNgFpP8e/
wA0lJySdyOyIpwVf/QQB4OQD8RdPmGjb8m4ThiHzTxPXfSBhtFey5oWmRbzP8Ps3
zIxTiQR7hK0jf0Ljt7yq8NJoadp5tjkuJiAfiweNZhPY5IP+gyPs3kf/JhK0fDWj
DBZ92Ai3DeznaxpEAGxYmj52wJscdJ17F4T89p5BONEWKdUF62kUiZRjeCYRmH0u
MKcfaXSG7l9q/+KUb9Ayb8SYgpXfnCI72dLCKoxBjD+C+HayziMXHOZ8JIlZa9Oj
LegwF69xvTS6Xff2hxGtvwcXvuVYAhyoK7A9+qFwuZtAmw/dfbTYPZzHmD3MEX7v
UPGpPmns+t8y6K5PYA1cBtcbmPjsynfMJu8G0O/oZ3Qkh2i1y4f/Pk8oRcpA1bDS
ZapI1TQSUm+4aW9nP/qdq4kedpl1cx08wF8665ffKPwYQw6lPPzIbbAySBLaNkXQ
BN4aaj7HPxjpMEsDI8cqRxroR/aJcr2Hj1STM5qjXjx6vqpr+ln1wdbboomcT0DN
/nrjJLUJUsopefrVqixYGWFQjezInPeOguWbFY+RtwfP8nA5cbUGo8MfJ55NyWdS
amUoc603T0rk8yVaMl74msXXNcMIFcwnmQfPjD2Zr6hwFza3UNZDe0Ew4xtlyLo/
6u+EQc7u1Nh1f+N/72jP86rjcIAnUuBzpziUxJJiNc6bKctphja/E4W/UGJo7KRd
3bjOBVIWYiQWMaMNL1/4egKduGLgywlF2cgBXD3uJ+CvN8quo725qEWZ+Ww8jQjP
5hZYQ2rmef4oOk7DxkERc+qHp4YA+Z0oLJM5tHpsTIHR6CtQ6re36Aldh+EIFzrX
D0j1LjP5MStS02ZIJBTVQTYoyuJhuWuEYpMdkIgNkFy4gc2dRrwzCz69hliJHVwg
sMSQEI3rTQaxk1snVyzftLDOiAdmfkg4/C7+r/fBRUHZo55Out82PORIJhdkgq+/
d17VMoTvrpan6J2xsT3htJcaKTRSOGSI8B5YVvyc2lBbgyuW4BCGj1dmm3+S+xg9
aTurVvLQ7kVawX62S0hDqdbm1mTWzjzWBsoJNg+KN071Ld55XrTD0kxfqbfaYfdt
9k3otQupDTlg5xFn5XEUTSizfobjQahXrE1yO/jGv56Jp/D+RPTKm0JfvEXPsJLr
EUTIZVm4/xIE+Xs7OI043K4qvtd2011l9dmaXMqGCsuMEz3YMXrZrgS9Ei+MK80J
YPidogaMEVghZvWZrJXMnqFJRe1iLJ8t8jClfRovFhm3xxzqg9DaNrfatg6p/zJj
6mCv3KZsXurttVCPilrmP3OJFZSXLGGkSnYtWL5a+um5B3N9cZVt7/2eqi7lp8ZA
MY2nR4V5X/t3w2Fn17U0Pn+7Zx9ESbOGHljWenHJNRbflxj190h+/8TDMNkIZUS4
VZaiH9wfOQ5lg3RwMokNuHIOo6UZyyOt/RL2dW8CO+19gK0d86bq+uUWmVybrQZC
XC7MwRlnNmaEo7dVZrlQrgGg0xuFa8rNg3ZETXyZv3u6A5LoyyFlbceJV2zX35nP
Xm9Wp3H4fMRGvYN5Swcrs1bUeWWBgB4tPw7uQh2R7bmJtKyLpiTxL0tN4hFj0zX/
DNLrGSFHb1tZoCvUl+zFUfrZlodCgC67TzmviPpGn2M3/NsNn7KE+uJjpwBkuuvE
h1EZONHCD10qLV+r97CjCJLwr60Hwk8UL05unVqQalARLT3Srit4YmKPQN/I51wT
VVga+OaBuch2FqLvZLSZvOQDVoBg0KNQj+NacygJr+Mon7TFg/Ueglk0ySTe4xcs
Mg96DnOlhyPzMv5Oto7D5YhNIQFuHDExgZ8UuwhR8wC2tgySvuFM3QRdWHD+mMwZ
kUKr8Auyj/0v6dsBG2MsCxHYBQJkuYGPaHsmJXZan1jeerGNniSD9ZrdCqlbb1Tj
is14roWgPHjS+FZHA25D2dUdHRtYaf6kWDQBLwSNQV8CNZnOWNrbbLkIQvlPtY4+
w4Vcgqq7C29NXzv1/sIi1174joMul+RU0dGpRsbsSJb9lUpPAnR0sDf2ibL2/9iM
V+52jX2Vj/Pb5L+/mF421DPJwAji+sRSsd1OAnEhPAnEg4vyA7lK5GqYy0r+rO/Z
DFjLyfRnMT8LDb4901uaqHyzsihhAIMeoQ6pCYV3qIxKyfTA5sSubSqrQY1vc3C3
HFVOkLRvQIUg6E47qZVrUbWnoYcML+ZgWSC2Px6K9RjwodKXPfm5I5BIcqcMbKmY
SxKD0Cxc6YZ/VU7i7dhJ7grGyfGVDApRZMA3biq2eCJ/Xfs0zm21cRNtPrqGle04
ZiSoflNkVoE+veFtVwsMGdMceqDvbmbjjlzfMSnonfNJbfa1utb/zOFbKnFX4TcT
t7sYb23lKWlzBsrtkeV1VzBHonf168vIaZA3QRIggw7z/am9+nC6WHAKB0y7x3zR
pPfI/ycRzSFNzeWnV4YG9lBkfRSfhj1m5GUxFUh3OEUY9IThGwAMlGnQNwQgAklj
I8ba0SZaGUlHu+QflDyO6emvF+ZWi7dzqtDrALxkTIBgOSwZ4aS4jxOCQ16OYlQk
geqABcMQ354E1zjFAqhb703Xv/vzfbry8apJISyCHwMGRdbpoaD7SDFlq+ASn+gr
JOSlX+D1WSbXxGFlvePYMoyfng7kufKk0vRov+JSHmmbEymw7kVCh49jBicfzYP0
X9tjdxNwFrIk44L0NxEeyD5Kuem/FHm8cueDTD9hGV7LL3TDTc/2QD3g9hn3k47f
RCCBYYHruJMqwRERNGAXBSdQDVtlNht5dc3bgeuWI1ap7cL1lcuLMfvRtNws3apV
8JaoSeBPZ1j0aNmhRn+vPWoJmGIf812CAbzrnYq3KfUY/9im6Q86RJGaPsRybFz/
2qm5IPsTB6rBC3FijcouUo4BIZCDfmkR7YVMnN9LUXegZRRtO8TyVz2BUO91xnZt
jEYCl0FFXEgqwlTV98RxuO8kQyjvM2SyjGifp672HpiebC+VEtR0XVvbYYzLSf+p
wflBa9IQOEELIu/g94tXH816IQOooQqRf8Ijr0CIWt1SFcPhRP6v7WoQdBaUwmAQ
onUC0utWc7ubP6MaFHEGXPaJ9gNlnstLC9/TMMS+JTMNJcS3mdVa4eP17zFdSeQu
u/gpiyxnODFigOr247xvMBrlO0J+dZO7gbhjVGRTfD4F6eGPA/vXnIpNFR85KW9c
Crtybh9THteRNRp7rndlV2Av0qkduS2FiHb7KS+ajkTNk3xgzx/eAyHFA89hBf5N
Zc1WV0sPlcBumroylPxkkxtx99rEZ8b/oiHXEaEPvUkmuha8NoCC80Og2wtoEJWB
jIPOiSAhOOs8K+iX2bdmVkIKa0PKL5Ke76m0JwMieqPG5ooY6CuCgX168l3hWkzi
sLQYeYAMnWJkZRky3sKr1jha5Sad6NDTecDHuiTYgnmlmTqNtYS4027LHxCgb5/L
xtywMc6aC3hjO9id8H/sBrThpcaj1l0B0Vr1W19PE6r1ZSwUuOAUjLFXeqg0kSWz
/wwLAqCgT9quoKk+goKvQdArrd1TgMUVUm4g5KdeML9jGp6b+BeK2cMRut59BGDC
knU1uml5nTrwLgYP9iJ0e+egCwnzBnlCMPZ//Nhj4Wi9VbhJ3vNEU8RnVTc9Rw/X
NtKE06Pp2xPHnBthJZXUn2Bf9MsetxxmqVSKr5SwuM8Qgl4yN9jaQxkwqGE3InQt
7Gv/2N6M2gmgMZpFgKeIas71G5aiGjmpJ0ct166elr5Gih2a4B9qG71hoVbcs8Ao
eb0w6K+VYrUsdxFZ0064C3+BU1jg+cOSBA+TOzL4o+nL8gJsAQ8U/4L/rXrPXYgl
0nNQP793bSBj+byKTr2OC8XLoDFWhJRm2sLlZoKTzX5jeCxAuiig4oizIvTkejtl
zS101xMZXz7fsVBSVIdaugaGFMQsfGh0dqMbBYWJkVRUODndjmiMqVYJwV2cPL1Y
BbSif2zd/rRLLWHWznTLNvKI9xlqsaaQdvmN1RrK6NNb76UJRBOqEDIIWclke5lr
frBfPvds8LA+OyQMo3vWbPJiKKrVaQgULUc+gXdDXid67SfKlss7VUjf2ZetY1SQ
QR9Tple55p6WQtl9kUtl5IdceTp47STdFIlPFJvOy8ijoJAW7S6SpFcMjYtdxKOg
XvpFJaf3lZ59YKfBb+pS1NPTAznbVV/Rlf/IphOLshFs39QA2OYFUR/4EuMasmak
aKK9xxFP26LdLiQ4J3YO+FLhKfYXJuNwp5exKp7iKjmoZSzWpVWCcDfqvQZKnRU3
Vv/akR88DbTELqR5UFhgrlphS3NIynwvB1eRjqowPQLbs8N4K7YkxScu9NmdIKQB
fp2MNzqC+I9NOpU2xNBXdPXErA7shhlorVqkr2GEIal8TnT6OYOxurZGx24F+EMN
kpL89RGlqaqBmcBM8JoELUyxhI6Nmng7W58jnWBxXrTRNkreE9Xusoazkzc+odiI
zd7zEAOXoeatNfka41yl5+0nKAJkDv3QRqnFe9WoxE9+rYfDBMxGBYz6pUvWL8OZ
dhWbO0ms6NXrcgGujXqsbeb3XsZ+S28jQqkrhoPL9fZwe350xDY0Wkwvm+yoRcHh
Rz7GvrB1AR/mUAcQnaCCyb7nVuCPENYbaBTKPAGxfwZRCtBn8SEO8HDNVaQVZ69o
i9ql/UsFMMZEX2ZjMI5d1sfHjDGY03h/7L0824QzIWfR61GCbQ+Hb9iOBKhfvL4C
bWdEZ7V7IlN6MLsMilN7lZhMrMa0Maz5bxdUgfEwba2VHyX+Dzg93LAB0ES5xIez
NnhcQdr9sV7IWdcuMk0/wWwsfntdMy95tiDIq77ibJjcFdVN/bxs1PKToqxVtYgd
4kESpe2vPDnIappndSGeDi1r420dmN0vsN2YXXC4tDEGZohCh1YKUN+xFoy2cMq+
Oz936XMsy+Y2/IdLgmR5CEyHrxBFw3Dc5732R2TsVbUerPbqFm+VrDGDGckCvcoU
Pj33Dhm9DCskTbqDXZiLfSj5KS/TKO9SrwAq5XpjoDAxtTBv0/l6sSBOQNNmKqV9
ENA27x3xD5OSoSAdFOgfB1DBNPWuY7aTNU4PqGCegA0t0zC4BO2t2lacrdN81ciS
IMPBDPX/G2L74OUEUDvLx0OzwPYKMfjq7EWpdXYDkVnEQvdGtUJpaSQVPle43+8q
hoFaG6JzIRSnk+PfxQQf/QDtOOzEq3qnjCjrgSAZhp/oRF3pgDIbtKeamWK/PRIq
y3xjBDETbyBySwXt2PMftB0KPbra7eS6qZ7rjSLq100eS0FBTXgVBpmILpTNDkPV
zzPzlerZws+8CyakCVFdAJoPf8uorSDFQ5YILb/aMX6PQlXXTZjWx6NTQ78KcLzH
1u2pR55RtvbCLt7KfJ/xpoZT4XUT++3jCwHyHwuZ9slCo23xlxu0+lmQLM5L5I18
i2ni+WtGIOcwBQgpVjlynj3nFt27x3TXOjSJ7vGDVJ252BBRV4SZCrHaOy4MC0B/
LrPwkmZMZ4D6/JxGBAku8VCN6NBiLxJUJV9zRWM2Zr3xD7Y7atfF83TJNkFir+k6
UhjlY8U7eLehzRuEsObhIc8D/BuCK6hhn1w0A3DZDJUVKFJEa2LAscpzxZ8/hdXC
Lj+5tK5z4ND1TQXI1gAHuMcE8Z2mD6fGQLIZc0H1LBtzZFXuHzfoUknKnOcjOMZR
izch/VPJwWZ1PjYB6iRh8DebeGZBN1BiY5MqbE4CxKZqkdpaV26Tmuwt0LLWwp9h
damsV4x63Cc4OFdc/TDhQHN161LxFWZ0B3zysWSeLOVRN+wSm3U7te4dVp13M4E4
q3QO+zKu8ZZ4K/L3bxuzX8qzKb7Wi7jU1i6MKJN54wkTYk6qmmFS5aKmgJtgz5CK
h5IKTjnQJqfzAdFt3ppnYpq1JGdwAgE68B/RkiK2FbUDERdOUxL3p7420uNUyPUN
x0D8wwPSOkbIQnPN3OkZh+2RK54Jn5uVpqUEsSOJXkH1Pl1wICcjED7g0j+YQXWf
t7vpidIvnYNcfek3eZqQf6MhjuY3Rg9Mf8JV4pJCPX8Z2Jf6/Fn/0J/wj+3eB4V3
TW0/KsJ5TRMnhatZ0W5lm3IhyGxQIFEECsQb+8K+FxVqrZ4tUq12S+DQJDWdw8wD
WoTw6ZuCM5JbPKA6QDb5Ejv64BkC/o+1Onl4akLCYoYWsIqHudUYi1+FEOJ9Xc2D
pTMSHDOegdd/2eeJSZGSq6O/KWrxy1d5THPdcUp4PItZYl0QlI+J/Msj9Y+rl1K8
ydUH0tNnKEojExsejP/CEuPeWEQk4pSyqj84qn1ONKJb67+uMPKzdWMmVvoTknPW
mFG7yc62uw/7DqLTSJo7MRIIQAJNXnr3GKmJfRD1eI9BMaAbJXsJDkXZ8KV93ilD
iPo1g6nQL7PymveDes7NxkdozqQEDVzEHF+nuvlHKM+D0cBLACZh8RcKHsd5JyKM
hGUUA6vfQ26Gllz+fooJ3Y3BuJzxl5x/di+6mcoC9cdiCFH6nrahQiraFe/g0WXP
EEBoXQ/8/Vvlu350hU36fVpor4oWzX8Ty4IwkuBe34wi0SBwRMq+4P4seHLQlkIJ
onVg+HyeBTzIGT6Ex4ZudQmtGSDePhyjRb3QVIYYSGSTnxJO613g0hWLVmt0wOHC
5QzFDYb+gvmeflbrc1Y08W4mRbOl+/XIOCX4c69Q0yYJ+TC+5HmJ3PGNe1rf98xs
SnjkPnkKN3v9D2T1viY0TzXT6uHw8RqVgPVhAohzvytLE6KBBqea461AmLhd9+xw
u8sXueYgsX6Mwn1VBRgKRrS9FB7khiROb+apS3aQzvqeKYZsuo8bwVKW9VQv1wTd
EhEUq7R8eClEx2hOCjU5Fkrm3aAd4DJ1qmTiXyUIVNEGnXQeExjgzq8kgFBigBSR
Dfr54bdHuWtMW2hFeWI1veKyBkiDMgkBJOOYI7J+NlAPW21p5pHuDy0vaybhkGlm
9jmEk5oWfYHClvwFDp00xHLn85r5UAje4HTjet83tokddoWkBycfMxUt3m2F/gco
pmXOeEUiJGfeURF9DeH28OoQARbdmf/xa4Pc7Jv7niDs3g70Rs1/A+srzbAYQhUP
ij1HbSvj41CuXmeitWVuNY8c2D1oUseoh+hFdzXv2qw+lyQgSiSF/Yw8rGbuDvxR
LOjdVmnJJHS1/vT0UpTmfk7do+S10mJ/ED2whndkHYim0g69Nzrz/Tj+m8Rby2YA
Eoz7cVZdmvDm4hBbi/njbISJyKYOl3ukCtnZwACAEALXtyHtNM2rD6F0c55Swh+1
bytU4IvoqnQIAU59Lyy3A6ZXDok3X11oTCXJmgGQc0e7MobiWZiz56E2VBFGn7EN
eUpTAfLWSM5FDzyoftNUfb4FiwhyeYrS7dVhB4V2gfamlxUmK4J2zE08XA+bKtDf
0rKOo190Utw0W8Bb2dkSOG4nv7N4uCbDeJ98se3smBVHusVWlFbpeiYC7wAcfUIb
m2P9BoDqH7YmSMcmQ9xEPyj15uYkBbRrr9Q1dYbu/Cg1D0V5dZKKWtvqhmkjt4a6
W/UV5P04mXj29lUQP2PQSWKpIxs8EmfoQDdnu6tDZVCt+FjkJznZW5LIdqr9M6L6
r1xClwIv7lo5hemhtC34USpbO12ULOs5ts+ob8Fd6rN9JjJWyBU94No2DC65TErK
mB8E0NrqHLowSgixkyZDgBBzUromSE4ck09hd1n27/6VeoOaJFZs53SFj0xUSE/1
tKz/h0VWYNxwnUbmn/iAbK28xOy/prvyLrqUuZzBaoUOqyVM147dsAl+HQiarLoF
/nA+dhIopCnYOmpL/KjPHZ8kNVrkiXen9umCf82orZ4RkLc5AuJClFDzfFEg4hCX
9tZO4/vO1AR6eMJK6IWXJ27muQ+s+Pv2eX34gK/nStP6R8YXEUyVRSkc3wIREDF4
o1iv2MyOj+WV57UuzPeQfl47NBsgWw2vRUcZnt+J+PNDiecM/lccI5s3zqi66atT
NuLv4nVG29Ma27lNZer5FmvYxbH/5KlqpxgPPW06NWcb5Jsssc7g9d4K/7vmjwzZ
MK99TzVfO6S61wGYQCFTatfqgEIhhpKfvz7nUMzDSlVPXsB4aTbKcZTSLsQuz42T
SGEkWLEC4g/E3a6lai/riajRt/Bsyjyavm+c6pSeu5O4HnXhT5QEGCHIWEaogYYW
Cxoid2qKw+XHP50Z10bQXB1EPuuH4fkNwQeh/IK3PBZ9mHy+svOpVkp9AH0lE+4+
Qs5x7v5fDyfOKBcfXKPeneDkgVObZ5qVeh9MMomTGmVS+CpO0OXMVjs88zTVbbsy
1u62uEoPji8Ngh7OwhmBUJe9aOmS+zu//ykF2k/GJwxcv2fhFN45PaXQDiDz813q
+CnMAmrGZOi2IdFhsxxa3w0ChBcIEH7EKBdLXxpbBkks1cqduzwpycD1COOcesah
41ZBPqte1r07rEO7ezIQW22gwZELNuCQulDFsMrFLpyexs2DP6b3DmdrYPSOYCEa
T3IwHyFbsqwzN8Xa2H37GazYN/8HROVZp13lphpq5rqokRGzm84rAcLihkeaBVrv
RowaEDghW6qzKeQxFXpJgnJrmq/jOwxQSUbiU8Jjuze6rRUPI/HRmyQnBKJkwlCb
XM2fmTviryQ0oPbjdfd+qlsQZMWlI1CjcJ0Ea9RHlZHYKwHqeNrUvuNBYYklhiaK
jMCfDZCuiwrbTzBbsj8bZUwp0YuIWwlLNU1Ov07nlxi/mpeK4yMHuO39IFZRxKhY
hLk+MojPkbMWvSuhgCJU/3vv8uUTkdBhYQselC2ds3ogdoolFq3p0biOGfmVKiSu
PdveM5h29C6FANavLKlOCJE/7Y5988WiSZLJrd3aays8Ykccg52U7D3GdCC36uQO
XqQL6tRSZ3kHzjz2L3UyY38Wo4ZZqFXrkyR2vFFi001bxQdWiJPU31mDViKOil7K
tk+JB57VaPW05D1Y11VKvLN5dcqEkiwVUZjlcteHBLDnWlBkAmiVFxeLKC5jNRD6
eBWNyYL8D+3i5dHuaMi8VtY2p6fJH2yQGLjc7INwkqwoC+AsikoauatQNdbbTWV/
HNKiAVM4CuErXXa+bJ0eL9KWHz+93dUSbqn/3t0VwRDKLAhjfGu2LNCALLrbDfA0
2j5MHwulWaruEjU0TN4eVjkD8NPtfFlA8JXC7tNTncXwPFWoftqqF91hayCLphqX
pZ5JHrZGdPeIjoH7/kBO+ElblBUKFP34vj223QU/pKnmEDKjHizS62U83r0/R8y1
BCdLHsV7LMEeINu1xUrPfayLeTG4go8VJqlUswmdCTY0RGsizmLk4hB3D4at1O9q
h86fTeTaz5EOwg4lM4B9x4yk8zZ72+QFrf+AtYtN0uvvEn1KUZniuRhPs/VkRUKk
Y2N1ib5mRI2Yp+VisRyJquRZjMqVulccwInfHKP5N6DaqLClUv5GAqkRzp/aXUsW
fJ+7kVA/MHTJ/c9+QcXuZg4nCr42r5K5JnKtrd3gC7dznYQwGlCYa1/mkPFT0U9w
8XpdBEXRzbNIum9Cw5U0ADSn+8KfRf8ELHUfTSN7w2bmZoHWm3iW89BAn8QiKtf2
UV1FFOrmtw+ARvWR7seMJqpqNkNE1ka8jfPGtGiimHAY44HYh4UF2zKwJ7q5iIFN
QDqC4SYHaaFCV0yXjCMMmE8EYS4Cjyb2PIc4tu0KCZLorPFdvgolF0L2VUFQFtRQ
1N55p5Edr06x92oFvivkItuGuPcCZb+E/ODj0HFJK/+fyYyvYpSF7ZPcXqcYBFe2
z0hUck44ySwVtIz6dpdu/UdHOqihdoheNvKFH6hFoVnLbywarHpfdNdHyCdvELWy
3m20VxBbuLI1TVVe1xsk38LPB9Cmb+a4xlHPSOXpCS10oMHUGhxcu9MakJ8a4cqi
bGhgwi+eiCohF+N+hMh5BY2fNil7cGjdCYsdRqT2YmBY+pSZboqsY31BBIdm6Fs+
LJji4fHiX2SYu3+8BVbEV7zm/inr34lrfz/v/c+IuzYx1JXglUDPOX6QwIU6eQTw
lW3UhvgPqEHfkcD5Sr4+FM/N2CKYT4XD75n58mXtC1uHltcmhKT4ZZdqvKQWrTtM
ciTLqc9B9oepOcbd8jDnNTDzcPM85KYhoVp1qBjYICCffmDckgaUWyI47PoBiPrj
6gaFlVtMhX9wOsS01uAh5Ov7mnTT472KTYDD6sfwkICw2EpsKZ96NLecWGWq0Epu
Chs+6xxRmB0i63UgOuyrjL/PwiN+mDVsrorK8taI+gVjIyaLVwTabqrtFnMd1JQ/
kX9dsansukUe/DaP9M1RSDLFNAngxTsf+HNLK46uPMNKGgv4LFPOwLGxvDxfFTMu
hrE7hEr220evXTWU7AsB6gaiI+EQqpauOaXtHRmR6jAH8+NSsl8JplyZOJ3K5z83
hnuorwTv2tp9TI4HMj5iKpXD718NZFruu0QyD593PULXBa/j/0zstklqu2Tsw/uB
GVKryX77WJI4l25okhd8E+uGmJxmoYFuxDc5NQpRWSM1TbfLhOG+eXIDwiBYJeoK
Gr2ZIjTdkyDaCvwBQtL4Z9LPtKS8WgcMoOD63TM5H00RSMe2Ud4lfm1ZJ504I6Ib
frtzDOHd4T3ZFH7oGooMjrk5XcmSOK6ahzw8OLpkDZbkr0m88xz5BXGakpWVdtXM
1WZOcEp/oxVCGObh+ID4pWv3vdYZKfNr+JFiZC41c71CHGx+Qj0Q6IfcV/GIVI/c
nNEePpdYoKl8J0UfpW2LRBLsZMezwG1NLGbiXzFomu3Gjcd0WQYi4QF+mKxecKxC
ouSbkD+r/M//cHV6DZXUj23uBV/j9jOZkEfF3kH2/BfLkXmK1SC+lerKwEIOaRTW
BFohRH83KnMlHa5VMn5/fluu1ga7luCwJxlronWgKhvOAogOX5766B9uMTzzxvQO
bw30mnUKWWNk3/AWlqSfizFuVAW/FlPDiZ4zfCp9WaWtQOxcFkD5r3yw9F9dofuD
Zn2wKIQlGVmM0druGgJlVHcLUqe8TL02e3hCyq5elU5i04XZTUdXgTPlUv0DTgbJ
gJtM/FDijLGBR22Kl7opkiSInNmgmVRxTaHri/Y4HF8nHw0ytMXCgmm21fYjAFju
7mQ2fSjTkEitYZhbOpgjH6dXXBE/emF3GxZ3SLIjLTUJ7wykl6Ijlva7tIfUEUcT
TvR4kOq3+t1vamRiP/cCB5p6doBJ/qLB9jHACfQS+vAwCIBc/NefDMmjKGkIAlFg
2Tw7wYu9YSmejJRIMZbay7UGR7pSlxaInOnEelmMCHjPzaRVAFCKhEN02x4rp/AX
VrylH3yVm+z4QAn32NXgIXncr4p1NFlefKhwnCG6quv+8sAiS2gneRgKRSoeZe/1
2R/cGjDH0P9ZuFAjP4K0YoakgG5vB6VcrqYww8SfaIx8Zu3HdGcosResigf/3eB2
WvtfqB/mhKdMu/Prq0/J8bJQCc/KkAFx9gntpXyfGwbO/AEPW2Mg6l/fpFyTmdz6
+1g7bJiHx2XA+o0BCMkhVIXpN+1UuHXSSInTUR1anfUgVgGIoXNtVJhW6JKK/Vci
x7vtfb2dhuzSxYZ67d5Y6m+51GfaJ88QtHcFAm+lRTs+3uDwfGiZdG4U7bCNQNmF
jbomcvnXX416Jw1D90ufNW3avZmYwW4cEUhuQZvjkKCGfjCGr9XfemL2ImWiwU1C
MCoigIu6m9WZ8eEP+eZ/wl1T5Up1aNggsafUj/72452Ej7+v8Y5lYQ3HuE2vFOEd
ODzZnAEpz3DZUhvJ2QBsjuUJcZLnBu1ECZc0HUG8RCqlu4pCi6wV2prsTz1ZpIVm
zqtztdrpO59zheJYcswm3P+MkeQYTjd+bx31sfJDf1cuTUcuCJ3cXtRJcnUT17Wc
OzO5wlaBjVX0OuEBv8wUOdz3SqLvZxFhG72qdRj4fsGf6En6fyQlkzXxuGZnqRMm
oIVVnBT/nhY2RZCypgbuZTTDBEm0FUF7OVgtea4IaCBpSviFQyJpJeUL1l/J/1iN
ezqqHBa4XtoYkY19A5qbWWVpqyA9NztPXl/Xz00ngGAP/4aoXLpV2rg2WV/8c68s
xuxfaWE9D+qFKohCt7SqbcQuEC6M0YOk5c0AUpDOOOH9xwg713c9CgENBwxMTKvo
d99X8GzeS6GJDd6Fr9K2UBdjCMB5yXPUtMCU7xepDbFld9CHOqzpSs+tSVYwKb/L
n05c4EdW2/vmtGhFkpd6uwrshvJfY0zfcbd2HbUi4TmCBsxOxGWvcEC3qg1p9hYs
T+t5Hg6LwaJtRc1ftqTxmdReGZyMcvX7v10NpsbsXMJhN1KKmsqEQ6HmusmzIQdP
FgBIUblgnaM25U1ZW0X4TTpHI0PED+CEID1nZo6TOi4SqjemkPz3aNVEvjnizaXL
dzoh/K1gFkOJu8EF9RPaHXF6U1WxhLo32fy6gmS/kuiMb1ip2C0ca419FLT+8CCp
OPDACRYg0jd/930kje2sg525akb4c0Lm1vfLbSO+bTttqbOPqHGtrG+OgSpLpKsE
VL1A1LHPFUEMHr7uuZ3Ub0TuEDvphzDoUKsxxuSXXXv0tBtI4kcg144fihVFRM5l
W0bXZD5k1y877jonYPIHD3QGcgpNTSP0CA6/rIG22j3yM3kayQ0f2FjygsxOaygH
hxi+NTIKgX58tk7+n9m4EXcTCLfkGcv3EHexCOHGpNV6+9ulF/aGJr3CmpVf8xbu
0zZJ3KTlm8thEFMV/dLeLKXdnVR9PkXA3pWl/O3W/S4FS92s+MzCrdPQk8Gu+T6m
1KY/1fZoIHz6WU2UJgAUgfGCE0HxwldVv2AgBaW6K0x/YFY5DnDOFqTl4gnKZV4c
7IXGr90zfBOP1uFXHAtVdZe3C7YPkk4CKGXlss7D4CTHeA7dAeeBIrHPqVZhux61
8kRM6CAsMhSikkC3a+re0vffln2Eqg4Z1PEwIZ7398sgdJINfolGQuoszSavqHDy
PeJN7jUnf5ymSRonDZjuaEncQpYYdzRDvsn0ccACAQtozqU/eSltY1+pWjz9cWR3
OQPnWxFyGcJNKtFC/IYTmThlWgTb8EnlyU3qc1MjPOX2jlHNP/65PpoyIDHSWNvx
rb0z7cChNBJYVhyS7+SofFxFj5M4i31jvWxeRQMlDbKrWh2xX2PPP8bBTDFDDXDL
vAgSK0ce3mnG8rScYEr6lAlVcG6TwHNUTwHdJh8NH718o8j62fbzb4EDUsNOmPgZ
Exc2gu4SWjloiFUt1P6/w0EUeF1OsL7peEgtwGQXO6rL0jfQRydJLO40PWuImDKc
WUUhOJAOAcwjxLEqN0QITYCt1eoNgEFT5zOZg07C9+7k4nYy4PMiHN3EBZXfZJ4D
3NzC1sxDwJO9P167R5JkqUwt/jeHLhT7XEVz7Tl88CPyPK1rymFfkygYW/8iuKUL
YruMpuOQvQzd36/vY43j+kKt/1//GhMciCWiXCsb33cNDsdu824em0Su+WxzwzoC
H7dG4RwHjqolLy+mL/F+yb5noxO1+3E12uIIobUyEQ7yZMVOkUu6deIgwP4Weu46
8RglgPyDKdbCB2zxMiDJLrxyjGPVa0cUoht5VSeR0/WFPQ22PPgbzcdpU+dREYcv
2WbchjXh6VajL8waxXGnbVELlBko48h1XZKIJa1TmrfLMGMgmzauzJYTkptfQuIR
JTWlWM4+sqsix4pI0rWviNzNNmUGQYxZl72wF5SpRa0+C3iz9+pvgrS99XORIZwM
7jRQulohHn1HjSoidMYeYffw8TXZpMtQ2NOwZo8+u5N/6WKPQ8FiwHc3ZYbWEo2/
iHRXF2QF4w7GoxgS7gLfIyB928lRvpdBHrAHQcjvOGz/vcs4+9L/hwR6M9OuC/7p
iaJJtb7g49e+oNiGMcOt9qNFlpNZobd2o8QNHeQ8bttUntZTVdtf2Wr5qaX4qp+A
mwwxre9dt6vqt0os1LOa/dkdrCT5uTLoLmVeOHA6Xnn2Th5td+q0HwbjsCdxp1UW
Bx2Y7IwSYJW+NfBNZaZGJ0WkAcysxY0tX3Hg8mh2aJyjl4/lM/+t3VN/UnHTf/Rf
iN1OeRkyYGbrbIQWHtvmK2KZRBA54duu2yfscDqWf01GNeW/juqUUKzntHHv9DCf
IEfEVQPHY2NZzQqr/L2o7NykpRVECDDRJGH+N+xPVGXIGeUYzuyB1X+U2Y6to5Kg
+Yp/cE9s3P4G0cRcKe+ifyqXZrhJw7pFdzqndvpch2t52wrwnyPjCH9RMcOuexQZ
oA0NUtvzX3oMrRdmuGs/XNPwHmTz4OWCU2L1GQadTZUyFpoqJpGdM/HmdTlMUR8s
eWfTkYCJJYIKcMcQfH+gUUUZWXIf12vhjcatYDYFq4vXFXPB/OorHZRw8HDrYu5H
HprkrouWHDd03s+XW/e6pd55IuGc0T3CrW4eu3SL2oSTgUYl0ifQw/g5MTQhjVMu
vSfL7Y7p1YQn8GydPK3Kett+9nmhLO+7OD/rY1LjgXevWqyd8SHSK1mKG0XvE//8
s0j9zh3HbNO+HvyL0sOXXjZGPShVXY1frg53+yDkCxBKjtE5FdPFLOYkwNnMM5ym
GISMdSOKxGZjQm5Dz8/VXrId5+WdDsxxSVdvS0PlnmNArX/9Da1fKfk/w8G8FkUQ
s4UU6xJqKsd3j26hQ1Mmi1ryQD+8M3vEupDhh1wAQ5Xc957nD8eNJHsG5BCCuqdT
Gb+RIunBRRl2LclEV1IuG2SmjrI3SDfyInehKlbAmUeKaTxETohM0E59XSeESI7k
z1MOKao3abAj1UO7DL+3axO4pbjQc9b58zjh7A6r/ok+uAX9esI3WU6Hvq1ksMqs
NdOs4UAsinBh1jgqD4rWGoTzvHn3QhUj+XWlPQo3S+V6J/cWbUpJAVt/Vi2FXZHa
9ql+RmM17KIorujj07J37Tai2ZzoMGsRTWOL1c70j7N6Rb+Auh0ldn4IAm0Xb5QK
PiJWPn6yUXr9LQm3ztpSe0Zo3fU/U1+gaDjc2giRVAk5Pxx5QOYoQfb2lY6LKGg1
Lfl53llG96cimWrT8B7/e69Ba0bb0P05s9MLx1zvEKuQstWYIHWtf50LMfm85qSv
OT+Ax2SRMPzo3JTNUwQX458BVwj08YG0SPOyLH+TCIT4x2l4+Kj5XU3DGAfp00e2
S2nDT3B5iV/xeaooNkV+nvIUAXjYfIkEor9IefS1cuVpBRJn2rQ11M1xDuT/aWfh
ftvbK4qYAHQXm/qOuEWuogCyeMy+XIP6jQTQ+TgorpZ/jNriBUMiFVgVY/prBZfM
tZiXujTg8tVvDvppk+8LguCMF3zVNSZnY25ToruQP3DCzLJLIrJWzA73ehxDs5jp
hoRdWSPzhLxMsFt4cBrwlGfU3lriFLi+ZLoxsAFIWPwWlEIgRlDM8CmgopzzzVG4
JXOW9E7UyZtL6OZ4w9ec+gxd3lAvdg5IdwTIQMsJ8KasM3njOjRn2Et40jk/Pt6y
ekzrSPZVT2R562VwXCzyOyWWV8TdkIZxQi0nYzbQy1fMDO7P1FX8kutLRDkrwlIz
ZZG4aAWrW2nlY/5NDU4mXC5YX+/sqR2qsTMZIu3BwhpolyAlGzE01l70aMjEkaZY
3KXh4HyEJs+WSOhGW4Do6ZJl9ubUtJPlDAeH5w6neAV6HffPpxRfXA5MWhZnKqwZ
6hAnu8dbJp7vmpQeI2NYnXhn1a9MKI/xMq+cYuyx+AmhR8MncbNI+Jthh4k5Ejyh
UqHDEh+HZ4BfrwwlLTFkw8u1hEG85McjTTFPQuD1O3+PpEWZ5RahAl5xyYQirtHy
cy3c+Co7KO0AB2YD5M7FKVALY6pSBgzUuKM14w8otX/wjKU/2BsiUyG5vKhaoPw4
dI9WfDRLXzZJzI92eQkEIDNnooC2zwIq1FVoycGjEz+vtOU4SdKkLVdt0NXAG+uL
G/mN5LZ60rASNMpCfwGrndibZA6g4g09CHb6gp0V5XrzKeaC9fIZkRmh9B7YnWCz
9nV5PM/dz0G8D2AWwp1pmXIQZTFwUKZ3/1zpDUISkDnuqBxY2nreaAEQaH5Tw2dK
mHwD2Dyh41jnj4dr9lDvpmHU+45KuDc4wrXxKdv/cfodO4Rh/Zs2Dj+BOKFiMryw
adlYcOHmRs8+n1BhTMkuP1EL4Txk0pot28FDMLDedI1ZZi2CjLSQPdlGCnnkBOjJ
Nokt7jeuvimHyt6ytH05rxmJZtaa/PSFxZapvXFTpdRcrIH92k6EfrqL1C07VDhy
/w7P+6JxIoSmyxDM4wHW0V8vZmrytSYisqAjEWHi/nb+o8VgDQ/u94wAAiz1V+3b
Q7CdXYIM+ncNiqowZNhnGCfwgukY2t1wIf7cLL63GJUP2tmiX9ykRm5CP3VsYUom
2ZeuI2/IPMHlK4g7nQV4ZI4+sbumOpdlxwwhinMmNljRN71Pw4Zd0peHqu02y9lH
NeJTWoAZCvVHfD7Cz1rICOCggy1jIY+JEhpPrYR8t5YIf6LThrYY3jUteJ6vAc/+
B9Y/VrtfmEMWUS8qG9OcpMNTugzXbKF5+OthXSOqxib4sksAaRTc2wDGQWTD07dw
lauhAtYJnvJqAUFdYfXnyb2ytWk7jv5Gr6icmew2GOUnHWaboAuQVwqkJr/iP+VQ
WfpvgkNEmq28eIBshQSH07/dh1PkQxCWOzPFXF7bV3vxnG5gMNvTHSmcpSvHTyH1
kPlhwZ6ezFtC62IBEIBTMnZqGDn28MU9hrZ62RUad2oQ1n0Np1+Y01DUHGtMQfJA
zw//AaMooK096m5JoM20fTX00bogaWaMUMv/a5o73WmmlNlsuF0qzSi+Zv3IxWqE
CzfFG0QAaxQxZqDE23wqe0nIxZN6pfX3+aewTlRwyl2REEkySH0b2nZ/Tc44Qfvb
Nv0QR7g7sl0A4Zr3ZHGZSkN223o02CqGf1TW79WFNGQuULGA9LwclExDTULsn/NI
Q69ZcF6WsZfhVhCW/ie52/SmjRjNeshRLtqKMgJfRO9RBqpA3mhH4cVMtXP09zYk
1XEfc9GFnPQ4XL9SdCgpUNaW6oaG/Gtm8S8l57yVgpQINh92vOMgyMov5/Jkmtr/
Qft4JXOLbUONQsvplemA0GRdRUco6tWMN/12GHxqY5nFCxc/pi6PiB4ZdehBKHRC
RUITw6gF5Mqb9g5kq6nNgmS2CqQI5wIvejQwO1zMdJedD8MOK75b2IF5koo/lnZw
s8sXWN3tjTMInt4OWedhsusFIJGSpRQrLcEGHeyCLm0KeFF5+6f4mosyGU4DCHJe
4pf7vEoeHfv5r7ObhgJv5Yd/umlMSUjaGHjJwgNgyQ3fSEGGF0S3+iIRwMy+XF1F
IXUkjGhTt5hDg0yLmKikYrRU7Q0xYuc4CUm0vqnzlooEnVQH174vkNIt6Q0CwgkN
2NgL0LP9oRN7Rx8lLZYlAWjFxKPFCCcKKw2XRvdoURRcwkGyoH4SFS1J4Cf4otvB
UWvkYoQ/KYWCnUqBT/qmTXomxC5uNHL2FF5I4lHP/5Oe8RzcG1RbAyE0O5LLS9dg
Xth5r09qTJVta392eyKrU0XUKVN9JZQHqhNLx/t2VM3NnG0I+4hcKqWH2drwzMh2
RDCDRcVjNKxyzFqo6RofxdkXXTPAcfKVvv9kV31YyQxlevPexMqDHKpxcPJjUbAE
rE7EVsHWkzYQJ58KUodvaFq8jj30xOOrcPzdHqe9A6hAU1s9fZAFtaGEtIFlaN2h
5DBqaUbnNX9pD8bJZZcKoc6OZk7LX6bsRNbCYkrBuWFvA98TubpMunT6WnprR2xn
3R1otVonHvJaFxHak6M7hRWJDgRjebSNsiZRTVGPhu26ZgqfnH0hn2f8MvSHPgHj
4ezef+qoZt242eyT3J7kk0hp0T+eEI2lt9lnYXOSMY2B/kyCFxFZXdDKcVlfeSBz
2hDCFbU+LkTmFRBS1tc17GfXXFAYb+GbXHMf6N9yvumoYwXePbcB8ZokGwVY+f8J
q/GG+mJtyPef1z6MapPegEoHHTYMOiITHKWSqk6VsAJcg1bq/c/+jkkInRTGkdFU
fitnVUXnStIKs5XRcEQ0L+UTG0lME5A0olfPGiewoK2uEmGDaoIh+3lVqpIQVroN
dnS5w93fAaUPAO01+DAAZI3yc1o1UOlFc35bGX0/y5g0bah2t6mGrAluMXPFMjxp
u36WAlAHSpW7tynUpjt10llaPnzHFlL0lkVAFt0nvumBRdgQZ4ECG86/Oc4uUzxc
g59jJOx3dfZOMFbJFxiMvBLqzr7BALiCqclP2pFWROOAJeIzNfgPFjnObWi7fsF8
YAWwYHbsVDXF/Qas0oGodGqf42LRrousKv8mE2aRqQL70ECSx/CDijRzOneZgW4R
x18S9mFPOvMc+/+gnNFEm1CH33R+WiRi3dL6aQ7Syma9hQaSyTg6SwKZhv2LG9m+
n2b9CNCPTb4kCbz5LRp1DjWXX5wV47rv1YYuhoE70JQdNeBhVPKW4LUhpvpYfabn
Q3GSK0CsQJeykZNxU1Gw04LRLp5aazlCvXHhj7+zh8qfi/ukncgIg7VLG7O419IA
dLe5E34s1gIWBYp8nJX99ajomjTj3/8Lh7bks1XIcWLiDFzDpY9qn0vAppT/9sVf
fVnBTLUfgz0atmwGLeXca+vBn/CrYvXQ6mfUjBK+wUXKQzkQwcOROCmVQjD31i1p
wpe6Q4VLzV9ZR3q1fb1UZKtqQPL5cZu8Ysi/oVzwq5i7f0dzC4U9DGrXWMS8eogb
MnpsugWGHYNf4ddoTCPpWbPWhh97SssEyYsumktC0yERuIiYdsYwzJR6If/bs3KG
19dXBXlXvomxuwwmKmdkKZuxkSuc9BGSMlvoFqC+c8IWJe+Vo2bBiMO+EZjvumTZ
QpTB0FiYf5EqM3Twj0i2sRZPCT2mrw+NLg8CpWcZLbtOwInXIKvHfopuo8GqSPiM
+yKOltkaUJBDC0YCSMWgfenOYIt4t3/RKIsjNmOgOO+wXE2NfzB9Oh+ayxTUjxYn
sEolPt/hnYleJYnch6V5l+rcuqjkPFLRmLF/rP9+Jbq8oHMye5RVbwvW0bOmKGIW
eEo0qLjlOdL6YEHvaQB/M/mNUFxU66638E8xe5hqcl4qw68p1Kk0/Ibz5i/wupgD
0NRQt37jZ64GO1+hQKxdVd6QYi4EQ16ro61TKKLEc9fF69uREIVBoqnfW28yNsHw
xaewgCx86s9cRfd9tMdTdhEe0BpzWtHazrBfJOHrq9CCHPchKSQGr1Kw8OsTmw2S
af2eUva6vypcgKhpjsxVdApja8hkCM/3nAJfES8lyfOe8uSTjT3qc+YVsgV+5W/X
Mn/RRLnrcuhH5PonpTCxO76yLDAK0YTIr+IwuzWI4w+jXIRqGFV6E6tXii2dzvPC
RzfZYQRjRFFQsisyDP/UjIslZG9BPdBDiKi//YfYM+wi+MHidExjKCV3TqyBKPlC
ryjGBtLPwrTuwbHYygx5h+9iea/mj7XBD5zjLsZC2vPqeFGdguG9c+Ih5wqVM1uj
mr6bnbgIEcYSld2bfJKk/1xPQHAMx8wi4Mrs5qUvVS5aRU2xttuR8VMp08udO2n6
gIqNRnVyMku/F2SLYnBc9nyRYT7gE89bPPHJkv9AuJQgEYPkg2bG+hbl2nGCKdnD
XCfxROu6nJyPPhu5xyntyyjzzqNGr5pw/9hBdBiQOW83P0aQna/Q684z+KHjZWuS
QtaqJd5uWxqd8tul3cAXjZjoz5ImOySlT9zUoRZhwDE/fLi/jmh/Xkq2XBtuNKMi
MlpM6z5QWabTEJvP8xfl0ikpytDGU9L95Suydxq6nv3EdXvXuP05I1oaC/YzTbje
j7MCl2xrIkeIAp0Krl+BAKtfJLX1m+Ip1bc46ubUgHjSCKFsZl5BtRLA8TYrTdqy
Y9Lg9cNQeg0K5upGPUfF4/fKW9Wi2RwKA3/bUvvArlw+uCO4NO6E+A+Gyp0dnpPe
zvLBx8FK64liZ6bqMmCT0061La6YjRiCv67QAyx3n7vF3IRmFoO43GhcISyC4W4A
EWcpC304eIhVJzXWMB/oE/uCfhyw1UkyBP9v2i5DvrVYiCU8m7el2rYC3LkuWlxY
bWF/r4MyRCoGCNE30eEcFieE/jQNj2Iggp0bSHzJbJfiVP0JnJR4yvOHJgVNj8h3
KuHpII+lSsUzAM7jElcMxTn1EqfPcYxXzxK7UsjNUX7N66Fh8+gg13L5gPiIKIHB
m4x/nnHbAWkJRuY0cGwtHDdgJjg8oBF+a/hqji9nB0mmWNZ5L0Phqctdrrn3UNzS
BZnHsh5yiq971hr/Clr7Kb4+PFvdinelpkqFJzR8Byi+aaGzlrsQyA7v8emqIn3R
VCLFgjhvadog2EIgj7QlOwrWa9jDwvJT54yE0RImZYW0jL8J9et7A4ClFXBusM5e
rXmXvwUMrIa/l7orv+m/YDcQyxm9lQxRsPYmIe5nnh5zeR2ndmXQza7aQstLbHgp
M6ms29IMpLu9gZqV3XIAH7sui6fWeCxICbsI17jDA8o3v66fzbNOwGBhl6UxDlk7
qExcp3nfqNjCNlWoZVdINYxQqsKi2ejqLiACog0zNbzuP1m4jC5PN2bfYbFwfStE
VY1JnI+x03+LDSSABIHcMsztYgehC97q1DfHcYG1l/gs/CFbfY6oM9eKD/HncOa0
EhZzneCaG/CwM9rH7KwLH/ow4sudvKctsYnrk+e8X+Im917OuCYMmoA4lvOo7TzO
V20MGRJw1CYcXeSS5i7D6hvkTdFskK/SphnmLHcYTg43CTgihbHg9fJKntt+GENy
ax6vsiPxkA2cBURYjTlD2sBYLSNPcaV7Bb1yaym8SY+Ego5CnPeXJBU4y64BpfzU
IvaSguQHDyl3DvoZnexPJcUvN200mAKf7c5ON/KJpQ0B82qCEahLVIeuy/6LCTcF
p2WL0MXKbruKg5Pb/z5fk73SSmCB+Tp/c3JKP6UcGnMUbn+2iCUN0wt2drIq073I
ZHucSdGnqYiGTCPO8fKct7wCeFWAdfMtxVFklV2Tr9pe3zp4vfq8xN1HmdHNUlVU
zlcxQiJ9f0YkrkFMI8pw8TxNx1Xq2TfimWGybpBA2XjImPpBEZ2VjDNrwiGZWPcJ
WllI50lXzFktRyMoIrjDS+Hl5ysSjXS752M4PbgA9oVoW3bcEuFnnoTcSBi8wk3Y
CymrClTlVMLUiJDG42IE5b72d7V+w0U2/yGODSGLvNfkTeWDDfs5I9lZpX8CEGsn
/5cH3uzRKltWEdwL7FnktBRzHDngk/21nbWX9l/wxWl8Z+KAZbTCFoYQYJKY8de5
DO/Kv5VSo87pW0sW9Ztnmg6L96xYRA5XVtCgri+ZeSgBoDm96AVSDevkQTEkXH/C
z4KeIRlRLdtuLgYzHf+rxgC//0pLUprUIdR/1RQUas8rmPllHOz/anpyC6ELim0A
QDSK3eBaWwmhVh7yJRQprr9nfWKPw9j/Js5yA43TLTSnYdTntTh/u8JK+ZfNPvEH
Ej9HSSU8eWWXu8hVbX/oH6Cj4qi7AgeXR7ZMnVhnLV5txxZi5PW1YhL+blMtoLAR
Ba0U5cLpfiHPGb3Prlw/k8pU5Jfacms4OlObnSCGuj1l3By2zKeVw8IfHiPNhbze
37FpRPlrUsrBuc9imnR7Yg4/y+UVBeEXkSBeTvjkRraXv6by1GammtJXu907uVsQ
B9NoUNvkMlXB3m4JS6OEQ8E/MuWHh7DwzdbjzNc6F0Py86fwPOuLBkDB5tbSdGkH
unJQ7yM1jXaW2kcD8EqkOSmsFyy38xwZKiS8l6/Ctvc+h+AU54+BvnAwmzrR5Fvu
L+3UV08kqoUX8yplC66Il7LmhwL0JczvLC+BA0Tpmf7//mtCQVnyajk88bJlwPrG
xMRpHhLn2mz7a5H8lYZI9Qy4w2bcRRfbDX5EcrPCsdQ4TOgdzELcvKqMd/vGLMCr
QJlKR2+Btg3zxFJfPfdlVDEB1dzWJFD0Yg+JEUTRgzNYg8IFBW0fF9QamVR+mk8A
rqqsAXGM3yxf5TOUpbjVbHN1gcxYO5TsCUfNq3kgmBVu0Q3bzOXKCpbjLCktj4Wc
ZD3vO8kEZ/oPq+uvjpQ8PhlT5fetb+JiYnvVRw/Zq80+R2O2FZm/BWWdZDKr1w1H
xyY4JbVcjzbNmmeq2zZOA5mfFNehwHKrIioOVXeeo1Kh9Qx8/HPrxlqMi7ke2bQW
0mCxVO7D3C+HQQAgOZIpcVpnkV9KlMddT6f+cPidJ7JKn9VnURg8wxgpe94CLOz+
orFK2WyuWKed7vOTnMv+hTHI2hIr9Pd7qCsdwZIndC1afnxTLbgjJaUjHo6y2rBH
df2uHPPXSUt/Qh9Ob447XZaBrVq8ZmS1COul0y+OdW1z4DaMbI9izet3Cf4YnIT5
3RFmHpPaAacv9Fi6XnmarZ4tL3w6j3M5GHGzvMNJHsXv6BSCk0fzX0kF9pLViLmn
uMSGCqEK3cLnrOh6PUZZ67S8py6yH7MTpyOYfEoQiNhHGR8/5ABsSZDwzzGutNMV
KyNjLFcRDRln4Z9F5zO2ItX0PY1voOMSCr8dGd3EHVmMpd/fiIjFKgJLjzbMJLDb
C/vNANo4leXE6sq2WGnMFc+lTbe+euz6vYGnubfwChdc4kDaHlZ80i/Edn7FYVNo
gNkcrWvxlppOqgVaSOT3p4g4+nTOLdek5frkrakvZmt8a0EZ8QlJNppQ7mBeZi7Q
OELX/o4a9XHbSTzOGzx/9podm/45cz+Fo51Ti6KIgvwIOcDijScwwX5LxvojVvTm
KBnd6jSLEcF9qzTr175kIAG8+MOeprKT5qdxam7Rd6mznBZ+fBSptg+LfjmjR9Yv
JlZsMXIkpiXG0PZ/eVmrGTkcoaolgpxbI1QbqatpEF5oqi9uDMyWkUGzAwh5fGkf
7Ecaphon810l3WRRWs5yTF0uTskydkjBuWUR0m0fRrMRT2rU3lKhTFpSHHjI6yeh
tcpHkcr/aIiJODxeKqsX1846qs2jQjh2VHaMCcvzZbC+4TLM/m2rbi1sERTgcgva
gQcUueXHf2mc/9mtTsn3vRYomtc8fYyFJEG2Dc5Ql5F5HgREKh4dcFXsWsz3q3sf
7fc2F8m6w31jJi9c6VO5s6j9Q7M8POw0EybSqO4jt+OxWC/Ph1FmdXIoCViegDXC
xKjNaDvb52vgqZ/c+hWyuzTWyGN9v5RzB42RCKDeSL+5YBq9IGnLbhB0uC+wVzFM
jJLy7R+1rGBMRZvYBUEsVo+temIlCj7wPKU5LZNQKqXp6WXFmB7GBAEQTOVsxg+f
Fxm6HWONiYqN6ppNoG3BlkmT4802dgiCvpN+9XhpBv8S40IOv3zf7O/c7VAlXoRT
lRUsp6D2JTmMkFckA0rHhpHb0XGdtud9+0/EBSTa6FVX7r8zFK01bImM2CGoYupN
/k/v7FBI7xlut9lQHPczrvb9AXhe779vZ9oinuhBJuaQuPyZ5MvvArowNSQCLUl+
ZRV8aVQ5dNa4FHlsrDxQcMG+R0S6ED18VQtxjQ4Zm3kw3GO73hSths0bQJP8Hu7a
rXImGo87AbRnTaSOFXtGBKCz5ZCV65VslF8C+erXZ5Puv7OsN2V4rqkxWYYTeqQr
tQ6b2ndugYHDyUDUyzhoYRSLnOuw9FmkbAS6mRqDXu8BKadwsu2230u5AD1la+JD
NMi2L5nLZe2oNdOzxkxadk0RgEKSjChcx18PSSsls9ijTSd3nkZ/wj0eNC37jK7r
2DKevVhSby+5LLCbUKcM5O8loSXzXxORElC4XOY7tGpjben+HbBMJz0GDCMeNRhz
A/7ITnPdbJ++vkxochQckXhEWXWdvJcJkwM4ueIraQhrNjslfdpSsUFhUtmogd8K
yKy+F3RleEZ5LMnR1ea2oZgvIQ+JZgv962qK3UvsWs2Yt0kEvXxYgoSepwDFGEFy
8Lc+0BCqjtTUpGjj2J+NTjC94gNMRB0ahlB8Dh0gX51unAT7HzSiLJQoI6AyzAMw
nnNzR4WfyHTSkPIgswTX+hDBnXjJLVHfEk397mzH6yz1Q4mVbe7NsZKKNWUIsos6
uQAF5rU8LxpUS85IX6TPk0hRd6d8Q2qYSYUn1mnxGK3tfOyJ9YA/NBA4ckk5gXqe
9HK7Mk/4Rc+XcjJs1IY2LTw5490k1CBzd9mRbzxNZwbOxNIjkEDjDTqWjjPfOe3I
MiT1qbcyNt7qLHISlCpr+0uYfpTxqWLpeK+baaXJVBnMKUsyNqaZX8cZXmG9mHdU
LbXO1pXlqo2K7NQBdo5GRAuUbSXnGMFLGSM6Un+vQXzQqyPLozMpwwh1NPyS6ea5
9k/UqZYrjRDtvVDNDulPVz72rflNCeJG3Un2IP9WhgvwpZ/WGtjvJp121gSayleC
KyEfQSc2Cmrc4FhB44g8pfCdAwzNdo9Xb+esWQdD6myE0mppTXRZcX1hqVPjbGIo
XhDczPjurRot/rXBV6smX7r5l52dLbFDuXuFfwfYSoIq7i5/HqYhDv++2dI+q2SX
bfBeeiJkmuXIHhZLdIV/kHbZArk29nXt7CxWbmFjQqxVcqpmewZKHbpzo9Tb5Hge
Pvsl4RZltceB3cniThBlqEz1nv5h+Vy1m7M+U5Y8DcKnqTd3Je6gVN9J76nAzSug
h7d0ehVGG2igWXzcHGa/VwdsnqQsBBtB+oLCnTaQuFNOU/tUSgDJTmpInOJKKcY1
zROW1m++TOSz3G322PKoiTQWR3hRJStgZvGUEnpg2O+PXePqjFC6DHszmccPn2Hy
faNtN82xPypC/tfqNN3FXM0pdcaqLNWhiZX+jo4NtxBGL5NmYfP0sW+snoqFZ+sv
rEXxohbLj9PR+KvtBv0hVnlM5xiImTAcq2QZ7rEZaU3Ml/hfkAe4YE7xdP8rLb/A
FpqsQYAwnZAHxTBeFmQs23AUHohRmtR5/MmpDH9kjx2kjL//CdSUkeSZRHQ+d5Q4
5oKXJ2xf65KIDGBpLvggE4tZQzNCR5WUJTLcNjRRodAPDj2YJBZ2i3GV8fOsXtDo
GAm4tVKkrBWbQkQFv7JTQ5+VlV4HEvsPMxNU8t/MA7+2QOPkzI+8d4KYRTbzcvhH
zmhrnmygNqwEq37UGsY4QPleQ16iRqAkKBvUJsCqm9qULHGgmgXrxK2bTU5yGzkL
3m7gWpXgGr14h3usHpAD0NO0kXo6SBbZUFGAx8BrxKP3tlBCai9qAmajIiBoh7yG
UXd56ep/CP6hMZMTHcb9XFzeFIWf1xFl6hwRdcvvXSazugdiwsVoWregtD7Mb+dc
pdlwiMLcqlFtXTjtiCvixmRFXHljJrBVk70bgeHJpbcfK/RsMqXj/wMWhswF5pw6
5mEcB4aLzJXAa+6CEOIWojl34/TUxHFk0Yo/nBdI1dIj6oHPg3bWBTrrnFCSBWRK
Q5kLKn9kketLUXLQgx6AUJImV4qKHfUZBW/cdR/tLzBaS4h3ihx8viY4SD55RB8P
Js8wAmlPJG5DDoUZ1q4cqgKee0TcmSSCFSz0LSdbnzlkDmQOoLhxpaxre1rU9cKs
vNfuZHUfb7eWMPZF9XqrIlze1n49E8dmANxbmAIbG6AcrO8U8j1zpV0qFwmhQvxC
80ujrXcTRKqPEldvFho17knwqU1kit/uVwYNwKyO6uCXNILdfvn1bFhWlI6fSz8X
Gzvwt+zydqJXmwHNMc6F19KpJ1TiJjUNTykW9lClb3SqWlYy4Z98t82bFGOu8n5T
OFeUTyPCFy9vMjN6/z6uG9M81q3Ht95yE+halar7jP49Mu+SidR7ohWhEHfTHKLI
Xzi4X81mkTjuSOBhux3e8/afNdUDXGkfxtlvl/onwHxO50zKVbuceb/HAJjG3uwu
lMqv25QS7ZwIZ2PmaEW3xX0xVLxHtYyrPbWeHlItlS7jaZCtLyNG0L/W9Rj/f51+
pr39i5WYRIw+3FPI98nOaD9k2mafWuWfJpLFscLQrUYc15XXsmzhr+b4LSiGCahn
WdSEBfgoynupr3MeP6LhPDKHxrU8EMSaXzWN8v2xoEuQW8EHAvnFX2rxkg1LCeeL
bk/Ok5kHf15GzySnIO/6OVf8gyh6Qps0bzgEMzlf6v9piOVzTVQXyPIpo5hs1Bmn
dTUuj1xj7wS8byYg/xP8R+C4MzmWNY2rm+kNQvZnH2d/25O7S3/p+kGRL4DlKvLR
cVJ0AdF8MRwrtUhc7drsj9IYlT9SfryZOeZi6K/Qplh5KvFVIdHVW2W5eHfgS1b6
DIzx3dHzXVKeUXLdcorh0/JAGdd+5hvevWobWGgIc1Ee3xTN1crSCEfUpOktpHkZ
HLdtdh/r4CqnZaaEivN/x2sUn0VmpCkOL1zrqOkWnDMQnGkLeAPnkM4Oxia8T0ec
8RZRjfXBQ8RT+Jtqk2JRJS2C/oZIPaYuZVgkQguark2CQPLV6DyDBnfxVixoqMp7
0C19Ki694oG5eKfagaYVNhGTqWg06uswRgm6zCqtq+tErxiZxotnx/L+c3vKTkes
QgtQCHXI/eM1QSuZ8QtOtfZCira9IqGiarjTWuMKk5bfK2PUY4ZjCkGkIqeDQeMi
A4pKBTMm458JChYTYTm5rCRRmsP+UFI5dtG4fDbzj1UhiiFB23vppGA9oR42IWxE
0R+d2bknuUg768wcBbFx828jOou1FCfHI+6gH6aTGuoZq6lFsKannQrkebSApXdu
6dxQkT0zRcgSY4BH+BaqV9yxW0MiXfDBY0mPgY8hV/yID6yBdcc1GIieE5ATfd0a
1hG5G8oOCb9sxsPCOiyWne12o6xmKU4z8uy5GKVdYrYX90Uci7fXKllcD8nq8dRU
G6TjD5US2pPR/K6svqgRPNb2CFM/S0KnsR0kG585KkMhj4d2kX+f/xFqm0gRygBY
h1dvUSurhlk1ukLKCsWTa4dYpRvqg7eC5pPteJe7jDAjmGEvaH6ULZqrB4iOb1el
P+3kB7yB3Rp4RBHqKKUZq15ojEmsB++urI7TWggYQ40StCNUnbhBbXX6RvMFDHas
wZfNfWjmW1SNeOA5eQLBoe228RhOVeZWw73O5Rfd+jpEQa4ZfET+EEn0n7EJKv3L
aqQ+fxuiCfhXRDdBp3pJJCVr874y5fRFwxNF0YnQAUknuVgPXQ1DUnu7g6LJgzO0
L+nS5smo2UmlBzs1LdZxzINvb2z3V/ddRnC8S/QZ/22OI8dFL9UHaQ5mzzTliYyW
GorqWgaZLiTXn1XK6Qt9zVXBet0sVqaqUz6dQvFz7pvf0UIYvzyefi1Ka7jQ0mJZ
Ewn3pmfNDEK+Tq7Z1As2b9nGR/C2IOA+36FEtlxACmqs1cHuSQ4e1fSt95gC4hag
L3EvibBDSHEWiAxEdTZhEqrHZTV+THs2VakJ8NW9gR/fT/PIfuUYlm6OlOSrkv2n
FVXjhyj/Al5s9EKKG9wXuxOPikVgrMSuuSrwrdwlXn7s6X0TxpaslVf3whRp0c6j
5gwSZank0L5TPu/6fsuE6KbLDmW0NGHMUpHpgktRC/3C1husaSojIJaJ+YzzizUQ
JSECv6zfN847FQ29bSt4OL6Nt3kZRYjoyORBr8ZsG2R3RVoRNvvPmIfi1Bii7wK8
0HH/uruMxDgbpROg6QypsouPOAzbigg+xWbF9rCt7NUicIsptswOre6DjnIysfL1
Vdx+HfTGJyCMRuGR/3Bi0WtNQxT8Tp6vFGkiFasV9M4rKfiMo5OknN30e7Dd1m+8
Y1pxNuRB3UP4zUq1D8gNyDxn5szxvpX1SrEYObve+iEQB09+C83xe60ZRhc/8jhZ
VEZqMhEfwTPW3z0RE1UjEUKvuvTzhHNhl3JTyCR18WnGCFMk7XiFjt2BBCjaaHdj
dB1RsvQPwjpclYYuM9jqwn0YWH+X/Z4DaqhaoFRo3Ix2KCQ8jJTZDOwPsGeeCi3w
PceLW15hKxIpUlrIAyHM8e9FsEDGzD86Jy7t5mkNDlp8j4QScERp16lgGmRq9XTG
ZW/tsitact4W+39E4sCYAmqVo0VJKq/mkDUGbVZoAUUzuKuhEVAl/Q0yrMlzp6OC
r8mY6cBwqxei9XzPmP1hNDN0C16y7xo5YXroQwqgJW68VvI9Br/Ug9k7et8nSo/W
LeIoNQgtFwQ1/+93s/DDJQSZOliJMKN2yFcBKervLB40u+JXmmBJifkvo/eXN1b8
/jrCrpE4VnYZQrFwH/ZAJEgl/Tf0e0Lsrc500DpbJ3bLN2PXfTWw2KtYoFYuGZRJ
bYEzkdDWVXqZAdi+NTRdT7uRFGF2icveSUsZhXWfXQPV+zVOKgyHyw7FzPABmzRK
egoMx0AHOyKhqZ09dFE9uoJEz05LqFiwy1Jn3oNH6ovjqYBqSfR9SmTgTUAoa+5U
q8eliGDTMU5NDcDR8QS+vrVb92hV73KGSZFkji5+3MIBhDYG7uQnjmX5q72SyqJz
KHISu4W0klhkogj2AYqOlWKo2JJjFQA57vZuGjUBI+5NJIK4r8oHARkOaUl+Fzgr
2faa/4R3olBloAMq48faezWrx5vFf/ctOeu/W3hj83UsJ8zptwF4ncN5oaCUjSRC
zean7qockX3heWO9KJ4SPwJaKNMnxt7CThpVmaxsDp8ewLi6A2sXle2dbcVWxJKb
+7yK98KfxQFIG/klIhSASVfbG7/87AFpb10g7NflipYx0AkfC9MY1K3QzgaHYYP4
0AVIKa/z+sb5sYdjNyzqDiTsF9hizm3DUUOQYdIm9iSOlVoZhk5s8yDy31Snu2s9
91fRAcd5PKEOYL8LvTFMHlpbf8oLAVXFP7b9TE06eHHdJRRucEUYt+j/C6u404YW
f6cVLWUtS4vIRnVYcrncTe1ydSEKRVIGpFpDVKxApvIOhV5FCI69hJ2rH2kfqAN/
n9WfvqwlqgZCz/SYv/n+6zMLSsVfO2z9zUbxp8iYpLnEVN6vyX9vK/BAzBc9P5sx
wvWcyoD7+tUAgj/u6JezGI2YLm7G5NdYwE7uRjKJ4VKDmNXcEMvX4eJe5/2OG7+e
wB7kObcFIewUOGhS5pFv5BojMEWHCVGXsh4BcQcboRmBaKD/VmmNGH3KANLnwF0/
OsjRuITMabRmhhRcLCuzxYbdx1pj0mf1Y4olhUAzb7EJoO5f4d4KpQps+T/Lv/++
uVWEcHLv1Mxn8OLHX3hy74rxwof1A1ST1QCPRXjLRKXaJTjknqd2AVxcii0Lw65J
IbNepkNndrH8hNXKe9ned9LkS6t8oCAfGlAS0VJPf1Btc9CIAlHNGoMWWC0NwT1A
xxkd5Co/OLiLwyqgTJM78YjIEiK/IrcTHsKP5BdzngFe28zLQAUugiEIs7xiYdQC
ttBfbJCkHe/yV/htFuG/1FoyXRlFFV9trZb/gLcX/lYKD+DDcM1mNMMWwEeYt84s
XvXdrFjh8uEbiORq0oiLMAcqZnU/PHPYj3exI47zC36sutxNkCu+JNNo0OyPZsXK
lpLqyMWGSdzN3WQFE2jvJ81yQUCEmqNTQnj7TQCFswrbdcbzr2pFkE7lS1uEWa4z
eQkId5Gm713jDKDQbM0BM9fHHPdeRzPDyEzchCUFBh0iO4qHfwsXZz7U3RbSW27S
7X8dy5hwCe/VwbPxvVxTqhE9CsJqD7oam9qdP7FMEw2VqL5Jk/tRWV9ZPiWdUs3+
UO3+VeNk7tZPKhekvpN19tt3kWItpL7Ae8vTUi6EiLBUF88bwcVDvxBbbjFY5LuX
z8jcKevAiQsJGKZ13pyqYh7BAWo+TAqZY9W2p4EQTjss++MMeCw7atanR7gzPLc6
XF6iI5bWRi1ysxOl9gSpN4Bwvy+aFxGgxqurb4MZTgv+j31jxYan7V7q3RVHlaK1
8TGbodhZ/6WYgIeZC/BIuW119vS3MlwVViTiVThSLLAlwUGbmTPhLV8jklP6t3Qc
7pRVVxG7CNaq4p2VKOyyKbZ4jc4rSIknfN6qwOpJjbwo5vbJ1zKIZuGh4Qs/mFVi
JgqvTfi2CS8btSOwF7FXy63Ezy7jqXbDHKff3PnhNHbJGQ2wY9Kq3mtOgyTbZn6O
VJC8eH0Rl9ew78f3roBWFI4MrCU4CQQQ52h1M+IgiB53BCVP7DA6Zzg5/Yrbo1hp
/DdK/FVhJALm0vHF55iWM4wK01+U3jnCIhH7ofuAeNLtKjCT4Z+CbQ3NodvYVs0s
VSBN1sJl8fzejqp8wNzkD+X0JS04CgAOsmm2dwTBYgkWPTp0Do6fG/TAdN8aBpB3
Ems1jmW17TeWB1/6ePywhLVA2C26VHPlvcVBc/yY4PbHfyyLK5Y5yknT9YoWawez
qFG/PBmULvEGtytvO8P9AP0aeM6+YRFjcXSKJkN7xQIwvQ2i7jRSNQy5hezlzkAg
AfNc8pE2YNfMeeK2HhRa72HVa4/9uBByZ9j29uQQ6NWUbjbJHrFEMkMj/OzHS+LM
EgIhIFJAIQhVbB83aU7NOsfFJIQ+uOnYosUfW9BUuor9REV4VfNO8IuMjNeE4hso
I/ml0OMx1m2ymaDh8zY6kjvzs13NptSkzUwBQoRyWN+yIr1ewB6NAVAI3hItKmNY
37TfzqnS9ZvHZoTKN06VZcsZ26vrK+Amjy8meRNhMr7kdgqb8bir+OJDbpwJiFU1
7ODEFiZd93v76xG7U/6LYgJMKxbNUg7nTAQ4Wnr/tXQHr+rQjR7bSJP7GAFHVvqb
xCXQuQ0USca+lYDIVZxoo1+tw3vOgiHt6IdqXi4juWLyyGDbTiS/uEkrOdaz2dd8
L/4i5tnTYW5CeiN4NgbwgGDsZ06rk4Mk9sgBPg4OC/z98/fwZg6yipUmSFtj/txh
g+6CGpoZNJ8RWSTb5gE+jrL4ZA5mXZvDWKMDFVdfG2ECNV+6zNMO8kDv+ISmc7km
lDlhcJJ7omlabrvb2mUNSyG65/QBlqtUGAZYtjay4K6B5gLYyrVwrbT1XHjWblAc
nIeQqC7G9GXMEhdKXG+JlftjlJLdtGEOxb9vdtfND+LzNptlaos9FKOsGbPygiJv
i+kD9lSC6u4CddJl5NQP3LVJU5GxumXFBEuHATB3x0o14KqXV9QmBoh9t6E1KX4g
9Jxlv1MXT2qcgJZFfsWf1cpVxG7kTyRfN4ldB2dP4wFCi/vUFbDJIWWeZoCOwMka
Qxj7Bwq44uGBDfwHfKB/YT6I6AMoJiO4p59WuHs5BZyMNvLhBLYzbuyEDiv37U8g
voQzzayRVRoKFMUGuenSMIyLafpA9QSg1sadLyorkJEDMEqTBcj2adIIyhOMprOn
J6TnOtUwSEQVr8q3fLKaZY5lhhT8k/HdpHMgULsuGPrC28ZcsJXS6i/+y3iasaZH
9+j0BIdtqe5vmOkFYSYQrM5Xf0RfFtRpVot3EZbsw2GRK948azNP2FyFf6O/FLz5
9+3ZcBxGrEH2TMYxE2Nhx7iggg+Eb7gz/Wqj27F8/UZgJOJyCsB+MX+MLctZJS6T
lwywCAXck5HKTWudMpz5PnfJZG7/Lj2OnoHIlIkxxk2fnp3j27+z6VuksXVlSZS9
NbcNMqZ7Eo3ST5ymJBRXyoJX4SX+teuD3ruylB5bYI4D4eSYWHJ12ggVebhd5Ewi
JKlEwP1dXqgCpjwtf1Xs9rEcieVaA0qurfXLbhMW9SfggWAoaZR4oc6K1iM4Qegi
XORRr1IIZxsE3z+69QxuzAdqG+H9GV3e3K+58uILRFIwr343ootzwCMPnDA5/xwa
1VNLz9ErqjBgEjCGtgpIH0+Xore07vY+fryi8LiUxJJmMGOK6XQVre12br5atLWn
Mih1JImIZPt6wNMUlCkJK3VUZbeU664DRxmuOd8i7XtQPtnnTVeTIusNwny28Kv3
7KzlqewylKq6mWzXZUsJibEHWx81dPxtHUEhNqr5yc+sMuPVtNOaQrn+tV/t9Kw+
cOwKL/9nyHtD5GoxuH/G4n9GSsehFfU4exkLGftL91Yl1ZGjsrW2eB5pvBEVmxbr
r8LuAtBI2Mb17lPo0J7eO/mOXfTE8EwbzKg/zoVsi7JC2FkwSfWJxHP9igvewZsQ
IGso6JzUt5xaSZm0xr7m6sjzi29aPCXk0rBZUEoDFumRZC8PyQQWTE+mS81gKcH9
4ou4CIvkooOGCsVuyV0nJL6xjOUzhZbMsFWtUZ2FOrpyX9oSr+SWKkB7QWlrp/HS
QAz1atijo+aRmxMHso84IeP4X8NOQcDNU1juX6LPtSksV/ayQAtFWILLB1WYXqZb
J1SJQUTK0vrAKFKi0dsexIVUIsjRLJrUTu0/CXy8t44Rh616Pq4er1Om0b01i/1b
Rpmjh6Th6Zz8cWM70VWclUg1cW7lL51SpDF9hgbFSLy21H6VJLOXxxZ5uQ3ih7Ca
PYIT3889Yi29o0+x3A4kRLtGQylj9AnZzEECSAG1OS4opVebNsFV4jl4K4m7npQq
gQu1IqPK5jK2StSjWAutgCHLc7/AhF8ltC3cYxmgEoAvzPZi5i9gd0eivalJOs2l
UUZVULSTbjZARa2gn8AM4fG+wHac6qiOH3api3QuBw9r3KJPLGimdE8qGl1gwpoO
9kIBAnc2Nu/noEnaQP1nAzAo2l5f2uQxITrnjniFlk60SrDPfsH3PyIlhmPcxmw9
QKk2Vn1ZhcFg6l2GFrA+Y2FknOsXxQExitRz3fx9TqsqTM06bh+DlKn5Mo32UF5L
M3yxZTN3uxhgB2LK2npeWxlJlwvEvbPiog7IURiuXr9G1KoJ60jA7AHxey5kPaa9
2NyfXlETO3c7bHjGzbI4AGdBTvZYlW3fEi+Hi+36SxyiVhDW2q+LlrYR5azEI+zb
g/YObdekfHWkkR5Wt1GKQZbA6CUB5hNkMeC4V7rF02NeBM3MFY1hbU+HxcyYjmju
UcwSgNzeftsrOFkswnZmYkutfETVyR3hs/NtNBIW4DAcI4NmBs3hieAoTcjTDLEO
QWPoAj5gpAQjaweWCUreti9Y4w7jbXV0X4InibxmFRHKp8RmkALO2s1j7TDja0eA
GQJGz/Y4z8o9XphYDlwLd/uaxFD+nGvGRFHxl3JIWbMhYJZbiTEvjZB2UeCQXr8q
Z4hxKGQ6hMxYnh23hvh9q8vCJep91CtTwX5dxiBkcCyzBShz/EJ4+SDWnO0hTZRW
ivSwAka2B9nigAg2B/7DX0m30T9+VQ6TdPz7tApsqGSGyR87+tP+gBBVkbANv3EW
b6FeIzQOMytUqwk5YQw1PDWLvWEbUwQX4bitmgs9lskCTMVFeSDYm6UACHyzk05N
RRE1s25Iab88C1Y7JWsccTjFCFPQTRuJfsd4N7uZAPz22X4aETgugdlLa0nYTfv2
W+EEt0Dcyh55zN7hBbggMgFTlY6FdFuWbsd9vIML7spD2mv0Jbg2EmQy6qJRgYEF
XANP9dkI3dltU8on8F+asd/KmbTuZBlNR6xbhYCVeL3Lpi69Ov/Pp/3ZX3RcGRox
HUH/qRFesk3WVVNvQ0Qy1+YhyBJPWIqt5PxbsTm89PC7l3p1JjcNzUOYF52B9OA8
3YJ0aFAjIfvfPa3cf4eLOlMjUHNSl91dYVn68owFNXODtn/rsIj4scEvHnhTCn4y
gfX1aH3q1Dv5c1EeNkW+ancGCMJPDgmQoPSm3NcrG5e/0Nl3RwsATY4Uvqq1Uomf
3j7AYJZBagXkZ+66dNitd8q1gD/054mbX9rQDDWZmdzeq6clH0sQsX8Fm0E6IkS/
UScCdUVJFR8knuuC29dFLa/yASSEYNLG48G6N4gfmaj/EKyqJpwOod8mztLsWcoZ
Pg1nUTDXbjg9JVXVFCrYM1ywooCR5QJqn7mj96XQk+H7XzDVoud7hEgAHf01Dq4Y
OnHGxCBu96ugeyey+Yoyax0rQ5/vQHWoYMdo4PiF1FJWqueXjAv98pTBr7xzRFe4
fuXQT1du+ETSw7jBanPZ/vH76D/YEAG5YsP2nNhDdb4Nnr6wTfx+nyivhvQczRSm
eKuHOcgvFpxRqfM/5O7kcFpFBdAXywUsqBFJYOfBZqX4ph4MHeYbUXFcQ7uVOKGq
j2fbEEz2/YdI+daGB8XEt4H0Kd+SiRhCr15CeOiTARZcs6mF7mGHWMtQcZwJRGLn
DVu8t4GSWhk5guWr3EjCPSRnVyyyRfQ/e3xlsRyXlRo7EW3eSAwQOEELmZRJr6Bl
wW3iRc0ie7NTWq0BLw9pY3v4e4CDQHEpyWo4S79i06hG+bNvYOqraS7bDI3TciM6
VGbnc0Cm1ktxOSzhijO21cyr78hndPaO7kQmh/X7cF1VVflHnWc9Pbbb3lH2N4JR
Db19U/ty5RJ5q/Q9+ZJcQNeIDEcToV4AQ3g4rttpFTTAgUBZmUp90pBXzRKGfFC5
UlgGcyYWHb3oNgbATvDZM4YHseA9WMnMSWMM9GDDbDKjdhknyM5aDYgh6pgMayvx
nTSaqKFM/t5TZirfCw1Z2gXrdRv8/RLTdXS5IqMmtH3x2vXHPfrS8lOfN2ECA8IO
xHo+nZjJjfcJJmrPQ5CP6Z0XxTv52QF+vA5668d1rrtdVv7BAmoiPtIQIIAYiseH
fuaCvBlVxj7/5ShlRyRaUXbJwNvKXuBRTGIXlxe3bGdlcKyhsCImt3R+KX8wGb+z
H8V3nvV4jaPmcYe7nXDbBS76jQyoLKxAmgUNBKHNYnHri0jGaUxbFCSRg9c7Zt7X
jwoJG6JykZP3v2jXScT7UnD7q6s5438mOGHNxEKID9EVQupIoAWQjBoxPpubzOE/
37bLkCJzsIhx82dvKIfQjJtzA/sItHJCXw+i8nSqkf0qTWq3jb7Pr1VxFtA3X+oK
i1fi4yReO75RfnpkSnxu0aU+cTNzjZEbfYKXd7tAok+zxY8RUm5nlasvKqjnpyKf
ISCUnMukx6Y4GL9DU630hc1RPlux0pl4QGHJOJEvyC09tpdgpZ1Ge1dc0ymTlHlA
nQBtrKTovbesXQe2nrhr+xGZ+C+mA+iREk+SOJpj3O4Q8WyFuoTS64toxUKGBKgG
YcEF9rhTLNTkvAjXEAUNuc2fTzH/zVo7THO9gmnZVlTuC7E7m95vky6amo1UDlMn
fZqYX3WTPw2AkMFpq2kvBT2IDMZpYDLUXKx+bfahD1wywSM3vd18KTHEbxFqplNR
NC7PzLmA25U2uok3oS+FwT115oNZ7UXAjVTO8IFRTzI1u6PIwnCjw+aWfS6bGVVB
pRzQlY/zsqCdLRWZzkHABgpPhGpZyAWJN94wex2iD5vZ84P6KPp4xQV22QoFpIso
jzwizwfMcOUlJoJaNwPwqoj+V8AgSRmzSBuHngwXFhG7Xese+2DkHdp6IxZLG/8C
d3G1xWJ6WRpbg7TQh3ArDgbsPxzO+7YgONSLc4cv6aQfSyn9Eb8biSy8fm0+5cdl
baANTl0UeFGmjThuidPljvWrReYvMATWi/jgKl7URb6qwaF9fKVD4ncedLlXjdCT
v/iXRrMopFGncxW0r6rdJ0u9PdaMTbAzZZ9VbLiXAUBGmJUY6zU0LM8ZPi7QqAOF
o1djPqSn2wPJNIe/sYc8sEjAXaNCrmVwwAZBlIbA9g2Vxw7Apwu/X/zavXAZ9D0z
rJvZ/swqhextyPDW2pOE9gYjiWAsF34P6CdkQ41d6PxZxD3V7YSgvagT4z34zMWU
ZXnzBWfDPpB86zQi2MAqUbuUl+0WbtQk53aD71zWz9t0QRv7SiKQHGeprSYgIYeb
ToWsN22SEEZyluMLyKCSQW63ERCkV42rXRd8hpj0//cYXT3DauiQTTZyN1iZXQ68
jwR/cai8hR0ki72wzhqVUQ0NBb9fezFgSlYa7uvbnej9oDDibZOgDT0r+EQSZq0+
JkUihficIaLaSfFkNNtRXcxhpHk4At6TtOe6VYxxdONq6BisRNyNpVceGeW8r68T
7kjOwnVmqA6Aj9TcJkMrwhVUdzQFijDMR/FegD9eKcZBk9uy1UJSGgyoN03zfLSY
PjK4Y/98bDszpMeusAdFUW+w5milgCOB7WvClRmc5KTH+p0lGaUCNDmU3uegZS0R
ckwT26rSJNrQWDhN9YlSA1Gges+ZK3nAlUZv7fjmj4KRsIbUZuI+R9TNAqphKQM6
HMsKp+SO1ztBVRI4P5WFGk+JIx4B9mbfhwUzT4x/MeHMvOtRXCaXyoLIwA24Nvi9
X6mcU7kWpqF0H7LkvkCyzjtG1x2J3tryaVOF0BudWiDHOoExrDJrFid1IbQGaFBj
DDzZAyLaPp5/26RfogBEzaqT+jtRa8PP2nvpDkdEdahyvcdiryu2dmhdd3pa4NRr
apYlq4ioqPWs2sQAwlfELmmWWoRI/Pq0SM8vIp6siqGGN284JfiqT5xRZWhukVfp
HSX1P9oCT6yMeY/HXiZEe2lUhB8J4okQfwKUANmXpwlYS8gr9cPaoVEi6DFjmXjp
ZV8omk0ol5f02ElS4eTMOubQLUb12vPGNktmQsCS/jIW68UQy08L7vZwA2+Vgsa+
CwSUK7OibkI98fpNy/LTUnuJNwV28fw53vn83Tjdqq2CCnHPIl18A6ARGxlv6hYT
/xyqh6y544ZnkR9ja02iWMQ8PbSQjW3fVcqtdstCNaixxqz6ZUycuiB7huzgHEVG
g1INKCpNiSA82Xrbs2QyQTeTTKQlwUZKSWMAZ/P+FD4pKYzcIrYdjEDuFqXKjQib
NaqEy22iK/YAvIFgZdXnv1ui4Ei4to53ofO22my9VukROVITtMQ6Wxp5v/ykb4HB
mV3eRJT0MxGkaJ3bwi50hd9IakG/zCYeZGJv9sgtWCNoiRpjKDSFUeOsCEZQimHs
GS18M62quhEaetIO9X0aR0ABo17OdSFrdlbOMSo1yG13sN1wKJupCXExQYBIYUgN
iwOPRMNxK23eRcjcD2Y+1RSDPTpENeLcbGLGP9BTCHhdF3qa14bL9W9Rk+/LxhGD
LGfsDRmjwJDex45mXo/KP0SXgwdesVhYiwSnWf/ts9UgoyknqpW8d6rY4aZDEXK2
QF+Rz+uDyAEbrB1YVMacjL16Y6TPP1U0I4EGEhQpxIW/MjZcCxansd3YwxT+Wld0
cYYFXT4+CfjS2WoSb2KiX82gGJoEDQL6jL4GQfU7e31fNmY4QeJG7pLgmqGQ297k
8YXQLfs4tRS+WojykGghDo7RkXqN7JMWpjmW6wAPCLnjDAazB6iSrr0QDmEMs/Bb
3ZL1LqvKPv3dbeFHNlDANzcVglELKmsdN54it6nbAcQW4gTvmqNRN/ugBIjJqRUb
vNuiP5dhKVQxdKOPVEGNs3M2uQQivHKr5glhbrgZVmSgVpAj2BwJHzKplEgcRG4t
okwheee/+/3C8rRedVYevAlcAG6wIgXk1PVDKo4d4hCtN2VYEQxMNSLff5Ih0gp1
r8QcfZQnRdhakVLXMnTVbljOMhuAa0i54VwPtmLFXDqE+YdznqAfr9JWSwQzm+OW
cAV5IoHX0Xm7KfO1zIiBlxshCrEY3Gcfl36T+e3Nqx63L8uJPlFoThKA1Zg22zqB
kmgsaYqKTURcVo6L2nNadkf4IZysU6qdwl9e5QGi3nEv297dnz8KOqMoxwzrmT6l
VP83ytNSMCFSFQew0sZEtwi7maY53X2r/mmwNs27BDx5FU5Mrnp6yF4unul7xycE
vBH8Ur79QLrBi5jtaiiyinmE5vQvk8/ZfL4/SgmZOgyu2h9V+XWOik1eNVyipSZt
NTtUJ/pieSu+0f23B7VJUGAdTSg8yIbUE3gNtzqCvB9MKroWfgLLwborxDjz/KbS
amp4VhPO4C4ZEGhf4cwfK3ujC5EwtujGG4GdAGqnPPAeaZmzcaLyEMOM2uHu7qOS
O9YltSw0vvkTIsEC7wSu/Vi+Bd8bnVKu6P4AuZJSJeHJNgLvcM8rv6B4P6/+QZtD
1eWmoYS0mKOC7QwmfMFq9Umf4AOIs4oSbYp+Ug38N4zoSMtjnoPmYuyU0rHRojyA
VwPEn+XJ7wygJNI/EYXMb/jxz+m7q/sn76JWuNvBgqc1QbsUecB+NTi0rf+JZ2GQ
YuWskjTYQYpL97SL3gBzFYT8V+HEaJKtFFEFJgf6VpsB78+W0ZrB6fyXZURGr2Fq
0YxZiOt9fbXsWySloeYhhb+2lytcT+zckj9Amba7WALFft1q2l4pM5XLpI4wrioN
INRqxXsMFrFAVF2nKSTEPsMbN+wbRhTcsoNyFx+l16nafwSywQ4xZaLTRExggTrx
lfNdUuyfILhAxpcnKrv+vfUkVsfi1lKl15VZfOzG1rEt05t2IkpnmNYG2VZn2ASI
Crg0Q56yVn2QuwlAVsEye6MMaF2vG+2rnhlorMF7Ra4YJ/nTlcaO91s3Q8Uh4Kg0
swKq+1PwwF1/YbJmZdPXOvgFv7MTZXB5mFAYCrS4oaIU5CGRoqI+Y4ypOtO0pnjE
ViNL5NKEc3XvAFHttQ+tYpqGvAZhSm4Sx8SXRVcI34qx6HXIdRpWqEL9uSTmXqMN
cjBZkg4dsEFzpsWoEc6ef8JkBAxo0QJwk7JlFGeT7au1stQD7krYR4AP5D1Tkd/5
eJsNYPRs18TY1tO9EYxPliC1kKQJ3/tPK1AofjiE1wSwTb1onNuQ6WQ7i5+d7QaW
jI+ay8udaDJpASCORmrhlAmM61ghwJhHNty4mcOtjf69jWNmNdisZkYGqEnQEx8x
kGnE65guVQIcI1jIsL5Vj2KZQ01IKPfOkdb++cXhvUREOeoXRuIaE6TElh/MA0Sg
t2AUm9M/KQtogdw37GMXH0W6jM/8TPN0xgPo2ghF/QMqq7p7ssRP8VW4cSCL+L7x
+f3gCbB6pXBrkfjE5tANKC+WRTLOFymErlWU+9Q+LVWfxugnSSz0hagdtsMRSnDO
GQtRBCPp4Eh0/Khtc/q4bZSPYHsz1Qp13C1iKKJFJYphSW6PFn8LunE3u06uphbj
gW5euG0N4z9qB82mObGxacQKezcPnP5zCdwhn6OhbP0uEAj3EM31VHEye4zeOHBK
5sUccKQ4X3GEv6wSvw3nHGXMdwNQT1g226VegDhjzfmG6saIrxAh4pDqenFTDbqM
/Yb+MYV64Hv+m/n1H4zVBrLlOuPERkkb8RQeGWtCoLlROHERa29st10UdUU1sxbs
1I3nI08xJygdMFZbqcHYhAikvt121aY4Nku2PphUs4BFIpw8N0HJxfCY54n0nTeL
25zH1ZmUG+hIhocO4CCC35KsQMy0Kakx6OB9I/QC//uV6KXMlcGW3RApVQvFb4Kc
gMF7dTVGsfizeXtvNuot2Xjmddnn3jEH+5eRPJzW8H4wT7ERvizgE3s8SuOGqgZW
ScIKI0uMCnb01I5GHJc/CMAIotWwMB/3jIcEuTp8kmHhGFE1Y95JdJgw375ylzeM
DTZisPQaa6jGgIRE8w37gxYsNktNjQQggTYUEROoWlhNSguS8MaibKs1CYD98Jta
ty+ifGU1GZltEtcJ/CC5dldz9tqOllTDg07Lv3F9iT5yUhF3dQD0rPBiToFNTDek
hqECZl+HpUKuNZKf3QcqI+Yi0VacSjHFJUN3qmmzmiUDnIWleIx0YjW05BlzUFbe
5hZ75l7b05EfXuPvsC0uUnQwH8S9Pr9S7xlpkgKpmvsDuF9aLFafM9tndMmpNsaP
k0/jwvERiFGvBf2bhdgWVEXD4MmF0e3AWac1s0XDGWOsbbfoCj6N0rhCCUjifOZQ
lY5LZKzq/U2ClXdP3JJp7FwOmr4BT5BqpaxSgGbUR6CeTXiyHkCpnZZjcICSQC0a
KRp2+/0fn+JtrkYMPNfsPjsIF5kLSuPUx5Jq6uPRGunHaRxXsmYTyuYH46bh7vqs
uFmg+5gbHLBuQWIeuQVEJwJLqg/YJJkOS5f3YCtNm37IBkRXXzaOQs0AVaFqbjQb
+dRFMWhBDSImb9FiiMzHnU0IDRrgKzEE12GvfFx+vjNMeEQn9mNJ4a9T4M0Cn4Ad
K68c/UhzuNJV1WucibHg0I9TVVTbfok4Ne0sr0sl26hL2wCg3Gnv5OzH2RT8AhON
RK1hrhjQ+dly5E9rHdqvEZp0oqAlg0pIUkx7H5YH6l+NoNsF4nRxKpSY8mertu1E
V/gU1Gt5C9cFdlsGFp/Xr2+yOfRaoHk/Cf7mKTnHpQGJ9xn8erLD5mLTMKB0GU+J
GnYi6fPzngFSPgmtosfvWGchwULtDrXeKhtM3kyJWs1Dl44jMA9csYpTpJXjohts
RH46sl6Jg8YDpeTW74kNYzX1B0bL9Hz1Be62H6fQWPNHvy5JjAO6YuZrWlZzNt1m
qcSCPtSWCtzsk53lRu0CJBkyKUjoQNLD/32e4aoBAvumvnOzSsfee+2O3qAPqEbs
98G5UiOQ8aqnx0mPBtARSGydJeFEZO1N0/A4C7mPJvfPDyNVC9vaX56lfEyWDzHx
P4Ho/R+dSOz++SxerZZBS1Lvvkjr1X9xEo6M1vehram/WP3Wrf2vqD4oLuMTGzAz
aZNGBpHgOPQ7H8dVu+3tuGp6taCwodsyBh91dLsQPpDMCPRWyhsN7yzrgjHjcUre
SM51Z3DO3Utia6jzTxs2eokQ2TmG2zZ/cw4dEsUAKbpsH7FtlgBtx7v91CyrJL24
QqQVCeKIRYbBT5R1+k2TAbG4/Is2L0uYu0HkhvPGo7TjSniIUDQXHKyYxoC4Kl4z
o2UldLDiqPqpk8AwulUFbXdMmEPyzAGuHNGfCjvpKnuq6nQ6l2Fr9fhBd77rfK7H
HPqJ2+lA1oo+n5tM2MBqNwkTompJjKyDZDFWjCMenupX42LrK01jwuQasn0AYN3S
A7nvjSd9MQGzjFsygpdJGTmQp1tCDHja6Njot2q/O5tNPCKpISpR9yNjEmtNPjIj
p4t2QJmJZC7jOtZMVZKw0A33n4LTeAytbCGuLPFA2Ayo1f3RKF3y7+wQjcohj/qZ
i78PAm5tgXsiboJM/4+cqpMcapV7kNNX1C2CNz4kYSX4Qs88kZZvVPt1/2BwmmSb
sBNqDO86JmUk3oqJIYsGk00ljHyZQLvjXTY6FV4JuTnM9DvYwXLfWNzQjgXhnNZ3
2UB3j2Sza8Fk0fvYvrdtHDnIpjkDEHBder9F8ftlSXyhkl2VEGpeis42KXx59tJa
fQDROg4mfZNhSekn+wnavOEb7h3ygPZjDfAbQKf6CvLUBqu9jWWOyYJJAiGb/Q7e
KYqLkBRuKx9miIeU0oThYvaJZ4K1hGsNc8BxwazFLaVZpV4wMpj37+JDyTqwqeXZ
7EbNp/l3GbH3a3g4zjZTmVjuBAxnSEn929FRhnVsMI+xNkuWc2P5zPZr0Ke+Zkv4
b1f4mKSmFe/UMvdo1XsrlPKOt36QLP8tk3JCFVyIWY9rzPfMRJTeWavelqv/1CL0
HFSDJJ7Ium+XchZa4Ibfo+A+ySTCCEkszmrW9zuXv+vSLkQM6gqKOfZNhSUEMwzG
w7GhnZuJe4ah78JVKr58RHxL/s3ynNi6XGOe/MdF4iQRlnvKzph7N5Gr0Q8Y7gc1
YOo8ZvrpFZSgPFi6v2hUxv5HuNWhIK65f7GqdLnsSayhphS+RqhJhhZyRtHsU+Hi
eYdQkK2z1y51/Cd9um7XbnnoDa2jm1vs2hGNikktH0EppBxYcF31PtqFjXT/HgZx
blMfuk64WdQO691sQbfg3UoVvi8sxRmYyTvi+qxyxovkyNXYKYKzd7Q0h/bSjHju
zUzvtrFaaiJhOvl7D4fJPRw7DMJedRoLwutbvR17mzEK+GObf1x2QpfqW+9xWxaN
S0ZwcOwuTLiga4eOq6fg2CIzOmVZZg8DUAbQaHTf+qIVkzOIdMNELw6Ec5VbOklH
NvLl9t8V+MyVkufF1CO4WkzMp0bD9/AWvVUBrDbqGl+8uHwIk9HiSaeKhw5yhVB8
Q24qzPOL3OPMooAJY7lbhOapVJY4yWDShyIdaENg9rr6q62p7LC8sIys08CWzGNH
6yapH5FJlpzphkZKDumgTyrOJDDEndwhKnnkf+abQZjux09uBaTjozVaHqm1/xRV
8iEt2A7c4s+po9jnKc06GJpYNwn1KIjfT+WTnQ9984BS3vjET0TjgS0cawXrWJ5L
e3hUd1cX8Vcffp5OlCrclZfJlQpS5lO+yH9vJo20wK97RPQlFj3M37cIJyU9dcp2
bBeBQ5fDpdKYHSRYSvMcX/kDIFCDfI+6fBpUFqlyjPr21I6hk97HaSpTtqyv1bUU
bV/u5aSj76i/hvWnNhP/L1P7hBS0Td1D+QhJyEk4p8lTx8gt5OAEj2aruz4eyMWZ
+irK6SMGIVmc+89Od7q4B43oqmhyRzxPGVA5iYH3IiRz6dHBCeMpxS7S5vLqEYjh
Iz2mipMrRtArSg5WpTxjRLDsghK1jzimuFWsCQTBEJPOFkcHRccMnaoC9Coyuqz6
+DvsnDuaKgqNCITGnjBhxWsP38Tb+MEOtvckV/yMi2LyHFRgNIZqp5utUG0r5wjZ
POIYeMn6t9FO9uVuWjfuFdLD7TL2ahk4ZRSzUTyC4nFSpurX+2HY4tj2w8sNTTpM
9+t5aDlS1fwBIxccaExZbcbBPhqxvmA6u3UHKqDGqx5t0AbHpOOX4IeGbsw6ryi8
O4nom2ufg0YOAl+jm8A1/tWRVI0OEddrn5UbsbDQgsKzR3B0+kaRXxAZCK55ow0J
t7iE1UwKnNRPn7KP/1tzW+/9DIH/35Iy18gwmOX7it5rK+V/2shBL6/0Wx7lzSVm
RjjdJisYpmKHq2ADdiLMcT/XoqPl26gqtG2yf95vrbS9XP+HVt42qlpkRN1TUJ06
6PdoebWVGcBNfHALqkDdL3990eN1qkOvjHKTBbd7XVygBjxlPrnmT3DxanMqt1s3
M+IzFD6vHlRqkXFW0yaHL7y9fpeHSwPwPd+HieAiEUwyZ5hlZ17OuwSXe0ZpMiIz
VKSu7KsFn/Lixmbsrz0rm3YqW9NLohsO6tL/IWogF4YJIExkd+m7rOKd76npra0V
y3RVUzfPLVS+K95tlZYc+tsNT0veqyePtNKnHbfoMpdsFm9UmYWTjp7zk6QwXHBb
3QOxxDdhqb74u8csTO2GZSe+Bod/L+9ochNyQ/B8WCOpL/1ofy9/5+aFweLu6vEY
a9mqrA6/cWqprPykPBvWh7tFo3h3iZk4MMHCqQRX8syUN9C0tuROSqbP2vp8q3kB
x2dA0Id/eWcvgWb69KFjExMc0BjtWpmZvKJ/7AvIw1H1Z2zZJhx7VGyeNARvfuXe
Cd8LRdu77caj995xHK97o4U8zzVJnYlnmPayYLxRhZ0zybr8uOg6M8owt3cD0z6q
j89pPlGt69TiVifY+upgzdS5JMwSCDEhqpVO403o2IMoyXM7e0jc889jTWOiQnjV
DVvsOLPar0Grt2uN6Weat3h+WhPNvYY/2qz7InbUioRKDNmV2bvuafgmygh1kNlw
sArKrFC7Ezhox1yD73S5Ek168ZhkumQdbaJgB2k8edlHxpOYlZsjAfs7XfrNU6uD
bHl2pf/CT4tF+tTJ5q9eb6eBAolX7bZlOVBKBeSEQnZ2BqoMH8N3WTse6pBqJoKJ
ZOcbL/G7appNwyeVEy/gk93Yre+ee0v3WyNrl+0XapT0rVJ0IBkyDJkbTg2lWvQE
zG0wWoNSH/y5iYCOsokR2dFbkT5rrvGSVevC0FS/4KLez6tpsTztMTPyO/+B2/bc
AZMUhuAEaflGehAh1teQtj0nZqhrIO/onzH6X67gOuN+brg0LO/y5jYMYFk2EMp1
MFdQ8ZCGPwvYJzDV/+KRaJVw0wlEdWqVIufkH6dm+fkSl8K0E1n6JM7ctdlNMzfj
jbcpKySuZSLMOfyMXhD60TXR2edY3Gy2A3y782mj8pClvZHCEpvyND79kXOBpIEM
miAHMJ1oUDhgKsGv+Ha2MUkekM61BFKEAfJOREookrX/Y/lKXPaRAHEt50L4Qlbs
8MP0lqapY4eu9KQgsjRCQziXUYuxXT8jd2up8lCI7N6q8Ia1rv+0Rm7ep75DgePK
sbnorWhbnZW4zRugmpFSVJjip2FAIY6x/Lo35QB8TS4YraL/Q8DHD94dUnnsiYyT
hB2cJdUF0XofTmCSSx1BEdU0ZvSfCXHnrOiRbvhCEhNsT2ubeXOlUmg9RjRt3jOJ
ygMDAJf9Ng6Ogk5D/2Qj/yVKv0y/feL4AzIao3Ls49RuFQq7FyDroMRTYJJyOJ0+
XD7O2Pl6o+hkfehnb0+HnxxM7c9lPytd7BLRz0BfrVTKDd3nmixcoDf8sZVwIn1m
c2lMiR0Dsec8iiUkafeBd7yzEGIgCATpy1aJebqVt1ScNByIiNf+iQcIkeE9g46R
ejmJcwYvjI6lSJn/BtHWmlAwuPEmrQ0/5EiPmwDZh0tumxgBKIlxtV2CkgnMBiJE
R1WyC+C4vE2fu7t3so5zokt3pGSnWJ3Ti2gwJ3P+AlCx6ZfjbTBgVzRR6joUkRiZ
zKfAEWueFwI+1cUK01w+DeomLUWxH2zEumXpB6T1g3Nh6GwNvIaEP7wPZb9hcUG1
FIeSOFSjF++SEgWRLNnnqPzxRMs4Z737jBB9BHDMApGwD//Zk0Z8NbmjX0trP4XB
96wawVWkxiJzvz253T6qujRL9NlBbDMCfRw7S2ifrK4tAvXTo/U4A/8wQlfYGeso
nEfcUh4rJlf3d/ItCyyv0MrW6I+7nOvJPEeTRVKcFKjvj8XIxYVnyyD2FJ38g7CR
3wARuBmHr/x7N9dIBG+RATe1lrZqbS2mdqmgzGI4Vm8UbQsXV9tTI7jUuSkzKhxF
b/hU04Y2Jb3U50z1u5kVW4Y+oKMcm+kGDE1m2TC2B/C612k1V2BLQyy3POryWuh7
SMXcHlNaLySQ6VTr/mh0EUtzDqCmCqIACo2T6U8Skl2AwXECB0AuB23KS6sA4PGR
mlwFaOyK+YSPUno9ntZc+eSxE7fJxIwLcg89iqYi4qfTcrDGyw6UGUr8pFU92nE9
slns4SWh3Comkdzun5ezVD1T28O4KhJ+4J9VuFUk17O9iDVZ3bsQe0ZIAYON01rQ
9V1WZ6BOldKpv1QKd7P0PIM1VuA6m/vdpHeEZJnkFrCTH+0ArsI9RuwahTd//f+h
w1OxcZyQMx54KsrGbp2e4XeDzLwC4s/UvYh0eAvpn+VjBX5/Hgp+oE6QYiDPWnzn
4SrZ/IAFvHFHdObcP8iop65c668J30A4ljzxkXV5LSjjo34FZ1M7+4nkut0aMNaI
IXOCLtNyNaO04MHMhFvCnVhwB5K9eYhIcypkalipBOifC23JWQ1hrao0Zf5IftUX
IJblPPScbEGMF05Ux1XMhni+1cAtwXz68zM6UZjvCvl+wo8oOcpi8Q+DA5+A8o+h
bT/cV1J10+ParBAgKlEfBXBWQKGGswYgXOCDIYaJaFFHO+SDn3jiKRCbh4SYKmrz
nnTxqNF6J9b+owBEauYgLeBFFB6a3v+euQbjPHSXXHr4kuLSBFAHiK9RCzyfOE5Y
RsHjjA5uLDy2mFMBFK6rxxAMa6kxWSX7H2PwGLQgYKtf/u1b3cZhcncBcUSMBR2Q
sh1IK6N6eR1NGebk855f+DSE0XKLIg2lNAvcfGwRYKLM/8OnAGNktM+FaLhnSM1f
jrS6tszqq4RN5NjqbyG6lpV3lskVRQDRxvk2Po+ufwSizE7irEyw1BRFUOKq1y2d
hb+QPNesgL7uqN3YTpnfR9Q7yZthEJAxooj+R3jUppOWRS2dSZAaTemQafJlQmnT
MUyQcNAeBIPrsmctC1S82ryZWgz0OfZqQgvRBW91u/HpToXxt+ZhiVnT13xVmnU2
9ledP9j7h/vm7wJ9qVj6a8Cd3JgRgyzoPFoP0Ps2D3pUGWwUgQi3I2gQ/P/TJvHM
FaGnqISs53fQO9zu78VLlGlMkqycw4uX1wrevAfHvmMzviMddeOLoUq1RQZNfYYA
/KJepBsuz2f/vFguE/m05iZYS8rTO6yHTqjy+kHUqRGW8zOyYfZ8eT+CKJKEi7a1
A1uplGJqIa027vv7RvSMdWOguizxwwQVGrmQ8iWsPRd/id5CIvafInOHHTr1EyxP
3PWpmSua09S1ye/edQpTkPl0RYUNUsxRFaEL0VT1/m6PQ9uip9rORnsC6EA9IYkE
t9PmoUMfqrXxOb51iP2pWBKPFm1M4kTZUb06EmV3TN+SGDvciDYGtla5+AuHaYy+
TzCPGX6c3jIivRbZ230+RMXaNeX6khyhahqjvGn/e1EJwp87ki0ZHlvHJGshFXvc
H5cVDZjcgIldtWlWB6dFQaXcCO3tba23u3OD7Ct7jHuS2FayT52PjW+pTP33e861
NtbtEXJmtA6dnNzLghPo94B4jsQycNqx6e1/4yhVWIV/8MUD2qE66cVEWpipXzPQ
3l2+MLfO7DCUs/nhSERmv1Jz+8/MiFKMbLrOLNO8PB9aDRhb3sflGcSIOOybWlfb
8sEZ+ESwV+cAFo8hNHoMtijVGehXVAAXTE7AKzoaH7mxbBYJqfZndgQN0MHcv2cF
uItKV2kFlOKWjTymxUObuDjQmev3EQYyiqup9cghKfB5wdsVGIsh0Z5BO3BYmAOA
2JfjGq/xJg/NmWt8PFFElR2shfoVML4KIvUhY0U7ye2jHsJ7x4BItGmChYoMY8Ja
Zckh29AJ//SNQlXUFX/+WiKzlquAYOl0gncLwKN9EW6NRFwYzbupoqDZELiuR5iH
oGldAH2HGvHshAil2CyFW3633tLlkxE65lhPYXzdKBD3LqwYw8XjqjsNPfR0Uyxe
T9E4R2QbUktgS31fWM9ZvQWHUQ7M+wSG78Xsu8Fjg9yRvoBxKLwZYJfnrTLAIrMe
cuukLbS9yc3XET+bKCS7ofTBzUB4fDQ/RSY0atv8vmleZiZ3nWu4f5iKpTEEyiRd
Pgl4n+9LUkgWs7265DJz5PYQkWZ/Dr1Vft9rXeCjTxe6kNdKy0fmDFOCXpcwR2/V
kidHqt8iYgotcPbknu1XIkFOS6j4vnn4dTLrZ+rdfcZfvIZTjRV9AcFXRK5LfChw
57nSE22fRg8/ycmhNOI+lUoeWWvVY1fpgyXhDpZWWGi6e8sBt4JPSkX87R3hTn8C
61JjQFyJ4I08mQCxzFNxCYcgtOLQWTvQR58SUyEf9Ru4Go2mzbUPo+zxP4gZ9ahp
/pPPR8ZCv/hgCGEvEGEp97PCnBH2ymccVtIBZdaaWickQkLagLybnVh0EJoUFW+G
1iqH1ChOt9IQEEgS3hkbOGP0KZUQQYkm5/NxXdMnTIk+HYDQpr41uREgKsF+RNMA
Ya/ogBv1Dn7to77J/fhFlGAiVj4zF1QYWtAF8tc1jY2mKx66+d4hwka+bewpqfwJ
dgd1ALjC7xLnTe2FukX0jX8y2D64OT6TiXGsQV4c2hO58fVpSXxMfiDQGzp2f6h4
3+QsOWD9PQrzJjXR0tF/8ZxLE4ukNdeIy6LproxVndu3gmiYr7vOvpvV5k5rHZ+R
+cy48JLaUEiz2ObQ3NzOWdCoLVhmOBGfKjY+3l205anNi7PNTLQkyTFI0D56nZtK
DWLeMqignSXQcvc0u++F6guKqqlav0cXyFfXuI8/QPhtvr6Df1gS6yP/BXi56Dd7
bJu/XvWuJi7OWIMgTrnJVB0txk71Xcc3ZA7O9r9r7T+JFumiGv1iOHAQSWfpaDp7
60GpCfJZyTW+W1HtOJVtl26p8n+HljMm2/bTWU4OG/DwD10eqdkooXyr+id4UqM2
ihiLiWbr17jrv9hv7AfkkqcnZT10QuhBqKyOzMXhZZDfz0rePJETWBQ59gnMgEY1
o2AexnzPWXwbyagrNBLH03ko0uqfXV07IffSLZSHklpfsHpL9yRqtMZQ9vndkOZ0
pS0ak+fep4lFAbt5iEYydT40bBpfFdo7D+fZLQsPL1RaB9ptaAgWBb+0Ir8T+4Z7
L4VPRx9QvzyE/pspmoaz5bFKmeKMP6JkiCK/1I7SXcyrTUtcbMNeAnj19pur5n9S
LMq26FnE7nykxU/DFLDCXnIoxLkin2/duqtM7+9rpEyrGwbJsCdNBDyT0Q11zhd5
RHu1KFefGkDBc4NlLOa1gxVPTdrlmjiBQAMLnOdNvSW2qjR1M8XwP9/mCGacg9dH
KRz4xFVDD4F25BuPABPwPeSnwtSj4eJNAXjJMrNFjeFinyZMeap9AnAHbZc1JISR
0PQU1UcwgAU0Bo59WcXzuP+GmBs3q9jQnhd4j01ZLMYKPxRZRy25iyi5vW22vmYB
lTM4SmnXFTNlLdtbJ03IoRUKRYb/8uQSPsZO+7/V7sQOkiaJZDAfFfp+WYUd6LQF
JbfWBWfAcpOStCmhQzAOShdnUJW6PL+TJ+1C1uv+pSxhlZ0jOuT2DjMigSd4fGto
MVu6clb6w19rUQZwAhSfeMWV0ftyavj+wry4Wo3ifn+vdWKfr2c/Ix6IlD9fMcjL
i057P9XRtK1bcgeRzZPbV9YUpj3tUAEjT4bYtqULDr60/5zVpAVRz62AS8iTqGL7
gER2JWGShcXBuH1r9MpzKp8QW4+1toKAwFwllxV8GN4vskz76DswkbCQZgLcLM6v
FyGseiHvDnBIE0yECvHQGuPhNN4tMUYeG3MdNF0kHYm2ZAQgPfMWX709Y6rfeIW+
kULOqfIIwiwbIqlq/yIlaZsDEyp2WQOiEKFgzRz3BBfKP91j941jAae2U/8gXFcc
MTaChNaLmw0HwqBj9e47SEE5iA14L0oNSxmC+9mvnyRQqBQCZ/o09nxzImHKb80z
qJC0sheh9tASRDrlQDyWfyzGy+77QYu99XVP5LwLkX3DeKTxQNxYLcciztJEEicB
xztwngjB1lED3paIMLnXOlUQtjnDo+B/mUiW92DMEd6SYsej752Xj4Ryagfjon38
BCCvCMvJ6ZMR1Kydzpi+UmMf5ugVkQg4O/mUPWmh2ixSMk8jmWGPkObADbVkLmjR
mDMWzyKmCmPRbx5IN1RaMeeKnWTT8j1gHSBHdRKCMOZUc48eYwdQX7coq1sZX/lG
c/i6yAHKsq/xnP52DdIRovuVSkgKXAWv6Acn2DX7EBpbd6u5XVa0E3YkZ7Uv+rg/
3BKNgEYAw8xnwu/8PanoFZ5AbTGbQ+a6Qs827D+JytdRpMWeskd+moINxCCImsQL
/g0uNhlwwyPM5hQHjt5TGpROc2Q8IJMdSN/Kg8uN3TOnPWyoINljGPVTrAczFm9s
7y7dV4HsO9hxhMCDEgNjA5KQwBcNgIR0iRdLpYPIIke/NtglEa3OMCwSJZzsmWnc
cODFeEf5tSEawn58P9sT/Z9g5qtkulmFgglyp3r4OIs9yCfJi3eDE/YNrZg+RT1+
uZicfHaIsxMmb22DkUzO30HMNU0fvKG0Cin+fx/c+kAmRqlU2W479ETrQer+2ZvQ
ahl+eVDTTuQDpAHPCpd9r+eYPXntc9fjTtxCCcIAW3e045bPVUmYvsF9oWRGF58b
NBgUWttG77SGuwtDEPWvvQgB+KBEHXWVKI0Nty8apb1MVBkhbT5g6/sLgV7eph/l
qSsPzXHPAjjIDeYSwbOb5/BoT8g9sZ1KuUSI9CN/YZ8E1bCmYqULJiPj2wKu7fQj
FDq0JqXnJkFo5G12m6EyeF10AMLb8HyC9CFuixMxJ9/QWyGpEsMv+S4w4V2qwx2f
/POqGkVT05IzNPFvTyE1zyIeJEQCIzH/E1JZSaiCJaDMGJPjPY3FgYuMqxQaaA4j
dPUk6rxhDrgX0q6S3/7NYObAKPDR1tIYho4FWgr25p/qoKNg7+9TGLJAXdDY1jsv
YDaGp/4g+ixnQ3wfewe/iPRhJ5SP14x0kcEO8dpLtALHM6E5IRnqXCjwDoR34B9J
miKzoVDztZRCEVkHlxq4XY1GUmu7MekhFW0YYIbL2JVx+tS+t4gFk3prjAza5+D0
aLo67b7IBW3aPpiQXZEHJj8gBSZ1lABjDrNUp2RwkncK894V2ZECd0dsE7D41/ku
fuCv/FdcHqyqALjdytCXo4Y19M0Z0rbuAx4FbLwEiUxvoLmNKOHyYKP3IqR56eeU
ZGaR/ifN1SYaAtJpNgXwLFg5SOQAVb+4BJ4VWAPKcqnbAhBmuBNJlx8C+J4g9G6J
II2hCj4N3xEcDqjuShcDDmb6sTEcanADKYBgUlAbdOSyfsVExV5QdpcfQ8yOixJb
A/W57vy0HhtkSsEE7ERVvMYJOQ31IVnyL3dTSxNbjbagS44Fgue9aYQQGPlWOz9x
RV5nNYjgM3t6yCZ5pDK+Jq7dwemMts2JA0aun2oKKw3FCDTuo4x3j7a+w6zvPxrl
9B+uudKFWZwYEL1Ol/m3IV/kSvyeFpfNWgVlPY3zZ7f1DYtn+qGOUa0tvHKvK8aJ
1jqYlUrvva7NUloWTpB6NzRi0MewdaqVtyLXE8kCIYUq407NugV0KRwMMhgcVW6y
u4J7agp+tnuWUxxpHvF+9YK2XBk+MvFGq9IHaWCIDaeG2iphmqpTZSls0CAumNg8
aZt4lYqK3HVIJx+8Xe09jCIVA7IEkN+yy33tDeg1RPF9KLY5Z7HARHh6zo7T8S3A
Go2/s22bOi/pUJjmfSEG2hGh+DfeAU8Bt5CU9tF81GYcEnBS8ftNqVldcjcNLjUA
X/xAdvNletZ2nahR+X+OhQ0xC0h7lLur2NyMybKsDWL0kIoLFp5P+fGS/tWX/CFV
RcCVsXXwCjSAOfEwGJwL+MYWfc+qzJRSep45CZ97HBjbLw4dtWllcuWIjWyfu9fQ
TeOf5uUeJyLlkMTm2oK2OtAvSThK2AcmaAFUZ0OJjk/Zy0nRDaKqflok0RfVs+bO
91pmgsLrywVkTpc409tjjm/F4WJeWFKImrXrNXLHA8Q6pvt/iy0Jsc+Vk68IWLp0
czUm/eLGinZ4DufZOmS7x1VAbe3npiOgLE4vo7sOuCiHr26qR41yBCFfYxPMX/8j
+3sQVG198WN+MLMKfRFL4n0K6Eio8CO56wXy0KikpEM0SQHBdzKvkNDk7ffTfvxi
RtE5jTWE3r8t+N7qCA839uxDyUReoG1MF7NEoUCrFJDXaGFwhTMACSFLpKTiPguk
aQzfQhOu5lrlVuPAtJ1RgmVKenPvYzpuWOxhSI1m8YjMGvcIeR9xhTTe6IEINqiD
t/SMHugR9Scw4JFv4PDxxg0E49BAD5wdKZ1XgT5QJbmkh+i0qItAOHFiilYosQLr
nV0F+8wT/P7QxwhJR2w48tj0TxkNSz8gBbzxHvZq4dzZ3oqhWMNyX8XuGCC5Sx76
EFp4v9cDTVIb0EaZ6rsL7Mkp7KX0PgSQwrEBa3ASvXc9uLboVEZsfB/ncOFJk/Uv
3uWmqNFsF48xODL8p+7PZUc7aWph+3d9dxJ5czl+5hFNVONV30I2zSCqlnuijMTM
cM/qfYAEj/+8ehH2bQAdS+JHHGlOTLxR7rfWtYG5KKLS1rda8daFaa808BSa9nWQ
IS6QuLtg0O6mRsUbnhPUcRqdmX/7+2lrkbflLw94uG8YwIrld2Sc4LT4zpihV6o0
vxdS+UYi98vcfHnwQY2+2Jj7vkYwzs2+XVqCJ20+2lglBqWI53d+nfmdGDnE4Rnq
iohdsAfkKDniopgHcGxY5No7j6McPXJXXkz7AZ6n1LnAJlHsCMVK2gWFMeRjUG9s
r96FSfZMQ/f+0L0t0w5SmSu8kS8IHbWty0AffuFo6SuqlbElp9Euqu6cYBxCzi7C
L8QyIbOoxC0IoQEATrFI/19YlzCdusSn0pK/sixLkpL03AZeFGsgL5m7oVv/Fsbb
DzceaxeMnFpj6m21IFp1z1XnmmnXusa60a2V+pPgpVIFBctS4ut9ruySDBR+noF1
dxbkwjwLEv04jhS8vpP510y9S7Yur+B3Q3SRGTBse8yXvWTD0WI3qBxrYeMr48lS
+ueZbdWYr9Lcefq7RQUgccHAaDX2gIQza/3wLHHBnHoxgwwX6t1oO7YDA0v8freQ
Z69VCAcE6YtLd8HS8p4EqQHcFYIsTiad435qgrKjmVsdIxqgp5IXK2Pc9UeA0A3r
vQ6b/qN2xx3d7lb555YxXYXx73zN5U/uU8sanHOiD44MpLeaUnbZrlp5+oBBlEBw
6Pc1AT8T5gtUo+6wGmW+Hp9XxK64Zk5U92afyUmkyXxPrZBDtOYKeMsglx+Qhpyb
UCvfU/Nf65TkUZus5iaPjEPR9s4nyAFpG+iaUAQ8WV/HZh1ngQSttRvqmCrPqTOS
b1U4WVEl5h802UHzyGzPUCs5Z14QYEbp2JcfbzPiDUK6rnW6YyVo6cpAnNIKmzcY
HEni2Bi+s0tApLxIUdrtdmx3i8lkr5r90uuSKYGnij0G/CVHO9vlm5NmFAmSd4en
/CDfrYlQawP2IR2C0FAuuabkhW8cxJQlKvt/C0NPlC6P0rmDGaEVo1OSos0CpiCx
yasDcQ3D0dEjbAqtq9f6opSPCoPOGPF876cFWAy/1ILRu2XbP8B0bOAIQqoeebMA
kQeA/LqVzwZpcNjtTWdljO7ZLQSHXwoUwIFxZeYc26Wf1ELq6b5yIE3ZB5hy6eXA
gLKUEi9+mVU+VRKYKpnyebhqpkJ+Tk9ZzDd/SAgy80Ihqe7VRP9ZWCCEPNKNQLgI
oVeoLwWjgyvhSSeFXyo8oOpdJnIGJg91FxYABwEEAeAUHNtdvhWJqrtJKihjzg9g
ob3JhyP8wdB7Fkc3vc5EGi5lWmC+8o3voUL6a99gCB5sHgtHrjJWD1dqvicQqIlr
Ue147vNSd6mG3KX4Smeza0CY5v8YloXKDNgTOvmjULCJMYEuvQBakkynmJex2590
+4VO2CpQV6mwa1kG23ITWghPjotlPVBkaXqbhf5Ldec3VxT3q5ZeYggiu2AZcHjv
nL1vh4cijmac2Wip+qP/zU3pRLdPZ8nairs3AZw4NCUcwDusZ3nxxKMeyVqEjO7e
Bn+skNhnLk6GJNuEh0zsQw0Y4aOTsmW2djwVgxXECQg7jKWc8M9Bta8OzHvt1Ojt
VimkvFVbxX54osoTt2Pa9o/AUoL/xhI7t9sjcbpHYTdy/rD7aVTGKdROUB+ew3MW
fFj4Rx+ME9M/I1WHxMkMg06XulTceR/SUeOFUp5nfT40r9o4aT1zzdDkZq7/q1Ui
HtOyc1jDvmXI6b5hxWVPQwc2xcaOSelR1FzixW7lLJVNcirv0r24CpA3oVXA6RQp
RnWVhJhVu0thchyXraO7wC5GgDbKwLyv99/ZoK9YfzXk8y/XTrzkIZtKj/rHcnEJ
sFBCEPVVC8fSzIxWG8r87TtUdd8qeNyxGH1NFw37YzLtL6K+NrQKOCv9b8gC4qby
Ote65Bp5AHqI0KkqSP98/Y9iNjlmWBV5zkyeTn3NbkjKHlN9R5QbkOvrQStPaO/q
Yy0z5EA9FA/ZUQSqWMutPndOyiAGiNpSPq2Pd3yMyaC6/BOJJbT2KC5QbO08uMUG
x3mm8AwCI9YJhlNMOl1v34ZBaCSWBEu188h4tA83V+tixpeXtoDAq6pN5p/0yMZw
XDErkT0eSncsZHOl3vSgh55Tl7blYx8aRGuVZleRu1XPoH3n+iXCy7lpZ6BtZcsA
0/SNB/ANH4dQaO6PYJivLmFWb2kWCiNE+DyIAOBk3R8dk3cciakmYhvRQNaiFBsv
2dWgQECrVvelmWrk7ZjpByfcaiUsgyFapVbF97Vq4dATFiW78saMhmIJy8AIJ2Ka
/B12KRuK8/phOjqX27d73S/RfEsbiS1dUOr8/M/QO1kHaRowkUQUB35mxf6QFnUH
qWkCBUzU17L1+cQKgxCxYHWhA+A2IBPkvk6Fh7xmr2S1wXVNcfqsjZRvPQltudPY
lZRMjSzaf+25Rwj70U/R7CVO+bGiI8fTzxj8vFAymePE1D+j2x8/EO/CvPME/H/c
6aqeP814nslDJHJzvOA4RPcbJMTqEcVqqtZIwXwz603cJTgWHQRzldCIOd30pfka
idboBlFJ3cflzeUESsAkbtQNkl9KBKK1QS3b1vaL/ILE7QP+OjPmkA+bJZcWRTYn
5yU/b90OWomkSARU3MF5aJQwcq3xnYd+PzN4DkZRH4X0lYM0nIe+C6UCFaZlPXoW
/Gmefyrv5oQGKfQL+wBcvnTtZK+Np3NEqTvBzPM9ntCTJ3btdsexUZ0qoChQ4XLK
DCeAF+qvowtGK7znEop6SVC13f64jK0W9IIviPyrbA6wOMs4O+kWrawsaibf3l1u
/3c3TZiRNC7sBDqp5svGT1/KheqQqDPpVZP1P2ZbmE1Gmy37ljS1rROGAy/aq+0d
QueP1I0AyA5d+vx1GMGSlcDw+/CONenE+p35WNMlNCArkGcI0gqanClb1/P9buqx
OOnP41pF1k9+iUwrGvUaVF98fSFQI9b6AyYeYasp6TRN3QrwakTrlhMuZDDhzYjp
faXX1Z8EyiUzMbWqe1aIi5WdAC0ZdGE0wo/+FXZZ6qxd7JBQsL26ZoIt9dqqfMQs
pKSlN8zA+XwlmRoU2SjBDVIEoTFJoDpjDrehnuK719DbZVXtjPAFMg3/D76ZlurN
wvvOqiRFLp6uV3OzlyZWT/EtXzcVt3P5YTkgNRHySm+jDzMzyWFU+cBt0xQm43/w
hCaR4cr7TMDnZv1LEvQbACWpgAZynSsq2XwshatJFTlfRbs4BDVxsJoXACLWobEX
ACcGIXQNNvuPUek7TWB2CvzynBer98wIIkeZSlvciYeEHNSUm2B9bubjGEI2b2uj
D3puYPCec4m2i9GPkqADhVu9T7UlAeZYMwjVeLNwpcigGmqNJ/L0rj1c1EESVsAt
uL72ayRvaAA62q3sS/Jy5U065THNM+ML+P4I0NcbQghjnwW7RlDYb4ORJ0UqVW/Y
GuUDI6A1JEQX1qWTw9f7jqH9B7xSee+MuFufGYNSFxPbxh5n+VlV9IvkHDTYZpwW
GCheuyy+pZnvPENNmMEDxo4+Nmk00dv+8UvBmvZ7EbF8lyaExqgjTZBb9kJBvsuN
Q2wbUQn8f+VoivTvZ0v0x9O4Ya9anKECFBzqyffZUE5MmAYyD9volFj/AYukQCWa
eqZI2N4R/9vUfIJlTNo+SaZAe8e0+Eq3Y6LrnHUzSNHq4R2SSiUqIAR9p00WH0GN
dTr3Ul3CC2/05qg3of5S9yiSVAaYyvpvPNmbiTwGG4T0MkLbtpUsyYvPqPvdJXP0
x0vvOV8OTsGT8P3hhQX0lyKc6+piR87/ICi9aIJ/nnSpW6fDd/urHQu46SEuhOgK
z4JTNIN6HFBfMM1XJ3+veTNvYlhFGFJOT93phm7/8EJCIFc85xoUlDkk0nqhtWtV
Yi9O1Bib0s1ySKhILw2uApwyeYcj0yN/Obx96i+EDKrW9XbXlGk7mng/6xFQnJqU
zT39LiFRQNsbBL9C0yHv6FFdxWK4GIc+YBPzGSl989ARnFzuSOWN9VRZQLJu882w
EMLrWNw2eKTbH4+tyHvcRdguWnuJNDRZ0dg7aVNUvDegGQlDvZb7aqsJGbPqdD5y
EQqgXxc6+ecrTwFTgXTKzDjxvBQeWWC0OCKtC65P8VNXx5rSKcuPwyJNlN0/hH0C
fTQdH65P8f6U+0vH4s4ilTRVLPWWfmQA9y/CpYmurVgIP+FJXW5AbloABRbe8+ta
I4jXb35kdNX8bS0BM1DRPNIj+QwlbkH9Du7V4CwgnRvnOQJkPA2SDKgtk+db7EIM
k5Hot/tkEYXwnF0Kah+fMNhVFwW7posaLtDNaw7PzJ4br9CrVCzS1fbigwGVcSjx
qrGiP+qWk8qNAmGLxV1wyrEVsziDHwAzPlxsdp9XOs9KwsoiP1LFv8vUYIk/GY20
gvgiRPSt9XnXaZHK160jwpmvAUjRmnGmg4112Pq6g6o3X26lEOdr7S1Tb5ImTHIl
jZjKTFjbbrj1IKJEKDDvsgfVByIf/RdPfw5K0E1CEW91Bqiu0AA9JgyeVAh4Zq5J
Q0ERxIQZvbHuhtHkAJXhcr84ZHozmEFVhFESyXfuhD8Ja3yQBiywrSVhqIIdfcOg
P6pLCT+RaW89ODnFjlG+tQseqE/uQ2SbvTuAZEMIWWFcYI943MYhEgADticoA0Pe
WTd6cF8Zw4lZf9wWZoTnrV5GM6/5FaNz8SNH7xr4+y5oQnedhlRwzMPVtpPLEcUw
WAseH7qm8NJl/jYt9TDJErwP4oupZ13vjz6LL/sPEcGRkzZd9KD8F+qPa7aeKqMf
ndYDhfZPnvkQM1deZ8zczMV5r3Fru+mmLctywlg7+PwQANSCuAAOCtzcBXJLeUqL
Bms50jBS4tHxBUaKQNvuhjLwoWaDv6VoA7HcF92XCY61Sm0ivttmQxHdpfQbANgA
HlGm/L7HjbH/gnn6kXpY+3aM35YFdedqpMp/+Bdyq4CsuWcnlsDMOVuw/5aVOoJI
/t9QZdzs+tBa2xoU4Z2gHY+kVP2IROj80ovyec1eX4cJMjFT4Zv36y0CIyvY87dV
UaN43M1n5TFxf7rrQpkvA5ezk73FCkPB/XFrn0MfrojQGSJWTtM97tjtuzVIFkjm
CeJHjSGZZmcC2mtKQ88UOYUBy80rqXn/5F8Uay6fTK7jWZ++ETjt3Sz6/C+2W77+
ArHDu2SkA4dMQa5ow8+v5MojwsXVIMTesWvizsTUlW0J+uEJSKYoMgQhsQt/Gx0L
vgcyFhG9ImnAGxKZmJ27sYIKbxs9sK8s0VtPAesEyBPbPuDHoYthy+PPkpa5I/1T
25hPvT47/kB8AJNJhNByktPLqWWpbMBYKzxb5G8wvb7U5bcrQf19+U0PshY37l8A
ExoJSBSdvKF+onM0N0jFqzoelGwTx6eaUuJmGiYiHl5K6c/g6At4N8A1YfyVE9ZJ
yqMaFuMjPTGG1nBYTu1zmJWhJi5oUEjBcEc0BU8yRZTcIDXazL7NTHOsdMQ1Yvm/
WKkMvcjB0SKFwSoyjuzpAyF9UiacwGLez0py/whyuTr5z3ulsYxb4ETbTAzlihy7
zu6VhWJ4m5RhdG9QEVjaKoxIzSfy4Hx5zNgR/w2OiSbdIWUNp1ebzeOtFApQ8br1
RxjTtqhUPCCvMYQXbKgOHo0rQN0Dmh+JV1HbeumdSzO8KstlbqNW+15dN+B8SNs0
C7uAfglPW6RyctzF6A3X7EALpqyr5Oi2iHBYK1fL5hQg5GNVyNLco5J/dWVzTFeK
lo6NQ04SHsW6rGdacFyIfUgDm48WtqSFuakB2+tZwlK5ZgC+1+70SXSe5Unh7lm6
yiI+mtSRSezdcRlpnixdIzhQsFBfJj+ckWEpgiQZcbLyDoEVEHnvipQdvhrkUI5N
iRqE+ysoRHGh/9+y9Wn/T+Nk6ndPXoWQaKPNGymcFuT/vOa5f9IuKwJfaCfj+9jK
Vat5rjdF/DHUtx4tTZde5sIV7sjdjaHKo0V647QeBKh0jCB4p+fV8Udk1DbPrLW/
M4QPA7T5I8d/7TaSnL2g2e8JmONo1LyWmbZ4YDA9pZOcCHLWFAVkAGoO2qYh1KLP
BVw4ccbvR8srVSNpvO0WTfTxsdHs+H/0/4dxkwvUFwFfpHRFbkeZk/ggGr0iEqh/
NvuS8aNtZv///wnpN+dFasvvSbOHqrFtr/Nw5f72jFJOihOLKoF6mV0rk3LPApoG
b24fLglCUFIqB5a8YAZhT7mQJMHJRqszaLmfeA/3g56hhEEiyX5xMQjPijxNB96b
8LfgDzFXpv7y/WL+AcV+2+Uyrpek7pM6dvFBtpVQMcluUBdLEkz1Y8uC/YZkzHJP
UD6nsk7pq+BY3zzPOezoS6UdwYzr7chZyIg79c3mV7sQBZDr6gDkDmD4yk1aMe8g
wYT6uvY+LyWhkZ32+yfCxPlOT2GsUHrBMO8kvBM+EF4RdnGSltRSzHIntrblG+M9
As8+eu+BEnwXWjOAznbjlNTdvNkZZu0BB5uEshb+dD1WxYxogPeh0Ni3dXNeu98Y
bR9X1vVh7BGlBjlEKB1O6xfTAQLW7X/MoIcGNEma/+XcwzaBdkF6JG7oZyV+2nJz
Eyt6odEcm4jyteybWbXa3LY16LLamHlZzo6sGHk7Y6P+/urRpzh72VTD9rxSwsx/
22PNzzebM6OcKRQHe/O0279XgFmcwO5uxnbq7xUadWg2R/mE9jaHYHYe62/oneKh
a28jXXCWA2aZtXRkrLTg+eTgKkhpoRvDZHWKagGTE76fuyBvcLtnjDXIBJFx65uW
Hb1nmKNn4AKz0x/yIsjwVP5Slq4IfRNbBf+SjjOH3CDNOWRTYGr8EKQ1duGkXTpv
M8Xjn2TYYqayVhZbXveaMLDt3Y5b3HtP50/6PvbTWJ/QTTB5X9B21v4DjbdP0pkI
ym//26Eb42dZxgYxLlh1WKCG7JuuvJNtvc6WYW6mAzc2z8Hvg8clTE8TLjy6I56J
2R44IDa0an6CSmAq5x8o4TA8njku7C1ANhzt9o4xZyIMrRA4xV5a6gyfBOw5xuOv
ekB0YfeP20t+r9XJKY+TTxH+JZUa93QxNuRgv79yaSCtzrJJBJewBeQjKgGTV5D8
0iiI17ouKygCe8U8sn0Jvs9vwrerfTpswbA0e90jaueF0EjkWAdwsbxP/uOsBycZ
h/Y4Mu4+YNqOXG8r+OvRA8YMK28mIWWfMyVPJOnrrXYHrByko49T50HV/q7n8i/i
63STLNzTRJK0b6DY8ENL6ekQRCxP+ovCfiPmT8B0sVeRO2yz6RJAeb8me/cdVIfA
dt4QhItEib2y8h4JjTIS2ze1CsP6J6PQ960PtD5XmgelD8B45y3JFUmFeR03nRWe
2e3VAT8tQEWTFha2fOsdSMlA4SbVVwu5EuCvvrPy36vSpk8W5yE9mXbKz1gasl9g
joDeFn+ducoqmDwpo2j8cRcyExRUASPO06wljXwwkA/8TG9mq4ofczrjYzBFAJKI
DI6NpOAr3ZLCAlszJFV7KjBZ+y7WFfv66BidvZ688rNX1q8R6TrBxDGtpybytPTV
ClZbR58ix2Wo2FT9NgrIYADycRwO+JZFxm4iNSI+IERPDObTbBW0z/GwkuJvJ8Jj
CGMuozeQ3qOyx46gxZQhTIKU8VIEzIxJnHVIFWhrkoGbqG/obf5FPZg7M3ixVfuq
y8ZzuxzC9T0mjU/3Sm1DGhp9uaFTJh11EUoIShoQ/0DwulTIFvcoL9yTlLY6H5BE
nFLqHG5hOcSjZyPNXE5V+irpa/cy9wcI+5elfxmXEOuc4WzlCZSZoqI6zcL5AzkX
kX0X9a5dEZ9ufvWc8fI4ftr/+li+kKpTUMVsU/VycgCY95VnLkhnUSgWyd66aIby
MY+3as6V2z14Fu0yYb14KX5w2INkg+A0RyH+E9JxcWOAqHg+VdLceeT0khtvtPoN
gLMjrHXXWwMsnrAYVHFr24ne2ZbxnRdkuL9X6F69J/wgJLjM+AJIDpC3FoGrcQLB
T/LnXfwrJM6Na7ge3q6pvNhOhX5BO8YKc/dyiXNT317Irs/Ki1eH7NcWCTcrKjTa
Ai4YkJPVk9zPkq+g1NH/learOSigkxAmakanbj5a+E+cAnhqw+vyduteOqW+yywz
h1gpinbwhB4zHiep4Z/Pv6NTGQpdjQ5w9sxV1AXEeIb8auq6iU+pBXlJh3TqldhD
GzjpMuQJB1mg8BJv2hvD6m3uhkEjufXFCnldpdVej4C9h+9ROnmYTiEajDPW30a6
lsRms0YOIO2rT+Hkn22Et+nnMqI0cZiKWQr3VKBPWRhjPQANtrXVovrukluwbDmX
h06kqAcPYkWCa1z2LIk7zbcAiOuY+DICPkVOSQcRN1c0SpfTbWbPcFMMaQVWk1fe
Q6FHLvOxt4zQ/Q52dTtwVy92wfPggFrrvcx/0doUWmfBAL2T6GigsgO6fZsgIMeS
QeL1tiyyeDM8eNAS48IVaSzRX4efmH3xXKN/NFQqPFMB/9YysEc7v0kOE8aSWB6O
d370U/I+XFgMt1Bd7mkydFf8BWpuNMkrjsY0cHvyL6ikMUeBkILPipjfu+X8e460
6p64XDhQwTRSHSBlGtb+82fvGYczAHXEqg+HobKpx4W0NtDJsWEmqATSL+J1cV9o
vLHWKsBYLVGcAgLgTq4/FW+KAws+ok6NdfJtM2OI1iEataAcQEwKFvxb9lfK8Rx+
CGemBDhMvCOkzv1N0109dZNuH+l+wFhifDK7/G6q6cE/uTE8OPOWCMroL4B3frVJ
GuMtCqGMLfeDM44C2uKsIgZvuU6qtjpZltUDb/QZYwXIAn6ZOf8Q4KI/b6OXk1Lm
VwZLgWUqqSCJql2llIacb7j1/OR/tBQuN4VDnHPnlRisUdC8tfr9lqrtXRiuNJxv
bGETEj9jl90BV5Xd5kB4YlKsEF1CZjQkLHGF5wrPeuwoGQ/gaFKKEOl05mNjHaDh
UNe9j97BsoJvA0iShyKgzFM2QEwwJpA3MNOa+S828CGRfPJsoqkOo2+NnPSwestp
305aP0k33nUwVtVfMdv8b2jrtWDd2sfBAYKborz/pLTP2mhg7swoLq3Rf9uiH/VB
mWzEFNLKs8U9Ae/oR7vvR/ENoPBB42LZGeXQ5gXgR9VohUztCRaPHLX4qtk20E8W
nAwjBk8qY5dQgS0GIi9O0lJ/ejXaALEErHMO2MUUAnMC+ZAX8fexFLaAWeF3Razq
I/zHyId8fjkfL4GXkOm+s/fVRGImLrfP0phz43mzIB3PAD28I7QY8UhTNdRhesYK
oHBUISIsIveMYv7IaWbGkSlHRc3+6+6t3orOVUIug1jmshjevcb2A1Bsg6X7hd6r
05ellOSV8nmWrLDDxSgkv1JcNr9Jc2j8Cly6DOpAVpxT7CzT31UQKHufitFhHtXK
aG4SbdWWIsKE23fHSviaoZUY8nT/BNhy6orSEtVfTqesdfmov0B/33zmNmNyBCvc
U/qQy4tgPO29QaEh5nQEzB3o+k5Sdm+J/8R+sWuQ9BdISpFhsDKIlUh2QeAK+U4Q
V0K6n58oNNK/vSs+MXqgwYWprGuPSoDA+trFeDXjxKYLYO9/jHUQs2EaL0bF6Aih
2ezAgW9Blt8vekeMJxnCbG+pxDmK5LHWMjw1rGvvIYF9NNeyOGRexy12rRYKhtO4
V59RHs304VD+cPNm2AGmbPTPTpHNh64FYqCSZcQBmSw12SvcLmmCUoNKbG9fb4hy
xB7WCOxSkEu1pPKD8PE6ZTs0p3XDJJ/BPV0rtHvVjlQSXDdNeXa4tvQAhfpYNWxE
s2fhBb3R2sn9yWa1UJm17DpvKCoTGxPRcEwhDEjMDZDTv9lOsHQh7SmX1niYyVS/
KfTMtGFfjOE7ADRORKAoE5bAxx+TyXbZbZaMAB+aebidURsx4J2i+soyJlH61H1U
O1BCt2HRlDYorEz44vk7JZoS6zwpw7e+WYmWEdmWXZZW5/HPugX9IMoWIfFIC1mC
AUVH05z6zgxDXN8KrgZCJMHqGPYGXuSwWUru4gtJFdlEN/FA6De5alChm5OcDktS
le7Lu3IMcjhbnjEGbcVHDl1O5kIusw/2oXmTbzoAcF5RCzfYXq2erB8TOM6hXoiD
qytLD0/R3SSb7TxN+2y8I4zpy9Mt+HzcVLdqAzX5YW/nK46xzpBGnEbSN7rXT3hk
13pXQ2kSI3WeN+oFDfTrBYFnwa8CfNlG9s+I3aEf3B8zWSmTcT924jyskycbMD7d
blB5br1Zs1X0TqPUHRSLvz4OWGCjQfCdx4+zdHvmQ63oBpY9C+8yxAjOa5nyMhxF
fdVBqewfYrYidnSaGCNEP5gO0nua4bnQhWnh/hHnY7DeKP5/jQyZstv6SPX/RqFx
nfYUKuWUOzP/JOAF/feVyRarqkdljDDqfpJqsqPhmFSf2h2N3PAYR9qZmKEUSjVQ
BPdc1pVl9WIi7Y8mNxaTunmFNCxnmxRqTH2MzBBb7b5z6A/1jbYvXURmFgSNFc3b
ZL7wPdFyEibHW1+BaY+K5vNwYIdXs3c4heOJVIFOzksOrJk5B8ge6z7CKj0YRhRw
s/uL9DsOI2AZXYx01N3mgTXmyzCDcwNibVyGcC/OymQg0hyEn7pz/jIuYr/i4fPe
SGu0jyqNaTqPySkkwA6Q4IJussGsuI2tiamzyJB4Obj/k2/mkDmrn5WgxVb3c3wP
8PW7OS6nAvohtlBizAHjxGcLiRRPDdjxm6ZMUQuizmOjElYmfiu6x8CmksbYUeio
kvFx+WrfDdsQad2+9nzUWn/pREUbhx9dnuxMyBgUCy2Ukxp/D5r0OOeOmeilJuI/
9FZYwrOzzLHp6sgSdiMVvo23PLFLDLuqwCCqU2mTVCk5PSdlpjAJEKC7J8BBGlLr
E9IyIGDeWGgdl7b7+a/j8rB/4RkXtJrEX99WZibxLlmhfreABCzu5Pgkjvaoa2gc
UMW/IGUIH6f6OYBdS1F8VAdnyUexN+C8YwfFgK0JcxkNtUSFNL9fTf3vPpa+L9ty
zLqIGDiVSiXEtIP6yQN4FPF5IRu120N0ZsANJbFzv4dggQTTJaqRUDUk4psNwhRO
QYpqGqE67CNXPA65ZqhWAZVjVCSg3kMWuGXgI9rKRrf8JakzTzRflIwp9DoAxM1E
vNDySyAUQKtAmyy7hsL9SsRDjDwpOJdXWF1MDVfmqQV2AucKs5Yxf5LkKHQ8czjh
cEJ9AhqI84aKFFgru68LvwECYeobGMVy0U/TFiTEngPnPGHUSZ9YitAjQ9/josbf
IW7JrMUkdGHixEl3MECko7fpZ9GpybrKZ4N4NrvKzuE5+mSRbn5Wd7I9oekbzdry
VDTDpC5fn8AxVCMd1P3XDE0uRT5rrOSIWCvekNP35+4NWozMzXda1lddsG6KBIXu
FRL0nvhylsL9L4E0Xd5IL8IPfiY92Wx4vu5FEMpOMho81oD7VeJLHYiHyZM3P1iO
USp4L1Ah9j8Y3df67/zOkXobB3U1L536HmgC96HaoYdXHhhFyVdcyHU8zbwaPkBl
136adlZOc4amnRjy0e6SMVyTzttjucEOhTYgtGjNQVu5DVssC00EDm6Jl41PBDhl
dHpX7aHmtFDNtxlrYa09ua72XucLFrJQ9VqfibjwD3/s3GZmi4Z+w/vhgqZ5/FGf
kC0aJ1gppDcY8pgRnEQWPSTVdv8/VQENtfsfpbd77omzIjDhvzmBnIzjhrLx6Qm5
1wiLoskdnw3MkJglj6pjwtarLvBCSvSyQVorJ99VYYh81MPyYGSkWmLaNCjqU2gB
JSpz758VYybnojSt+AqKG0WuFvHR06LICs7MNvItSY3MfdPfno6OeCoAmNdW67KH
0/X8paq0h4FYmB36y990lPI5YKgIuTvtQevU8L7ynsfM5Aw6dBo94Ta2Yk94g6j+
37uL0m/ItGVdJIimxxuT8c27o3ORfdaJ9E4zxIALCj6XhBX1jJchLUzA/cuN4OQj
7bwc2po97H/RVO19o4DMuA20HCCNnzFuix7M9BXtI0XmRrb10cnPMdAlauLzqWT7
coCCPIwspMKziWfCQjUxrcUwAYWgnsxVFIyIJGzT6Vvm1uSsYA4/s62uHCEweXf6
XXU83ZSPUsM5v84gnhiJZ0KWs6SPTP8bVum4umHd33+biaQY+/2BrbGg9DpuZRNz
B2pgjrqALTYmTOSjbuUPkdjXk9Nl6wDTvw4i3wGgz0VuhY0e3pCdDz4s/bGtrC+M
pvVsMyYLOprYJQWKeOQFAz15eDxGJOLs7/IzAgo1Qo8FxoOiWQjgUhH6AN1lB9sM
YpenRxj+rOe7vnauRoAARfdhaQkzNA4W6C+HWjfZw1ouvTaKf+8m8hLJtWAHkcf9
klYhl/k7Onwj26XU5N5UBGPXdCAUrgx9RqOyb72EpZFYIMRnLBCWcFx7IjAUxGfA
jzqQ3uUm0cF/OOiIevOaRJwcNhfbI7VOBL9F7WOvLkdYipfzoKbgVULiNLmVf1nq
3p3JlaKq1Yse/DNkzNCJv+CGkmIu0kpCIUFyTCWmnvnTzKOQ1FOXCQXqsER7PeP0
wwyf2RFtOvhWIHpW/t5op5hFMCOwukSoQ5JHj78CuJqCmivq9P1QlRwaoBVDcefB
uh/I/sqpJGH7WZYkOlLM54Vh/51rKp5pndRX16FK3+18S/p0fiomF3XB2UZOfb0g
7sQK4tFli0qxmewb1y9yIwHNDJCg8zIKzWBbyNdmnd9nIAVctbapUmUVLRo4XLQf
wTSmToIXaTHmfVYI9QJNCoA+5eCkYGDHw7LH8IDW2QbTBf8jJXWAS7iFSahHoQ7/
c5p68hxo122183dx0QY+C7Wob7ZvkaAf1C+7aVDtYErY9yue2VfUh3Mi2jePDk5a
YdHXgUUcLdC+exV22zvBkV63woAgXVH1vpk/VdGr/8w95+qL/RIWGSv7CzqCmm5E
0khAM9ktjACi5ZTUlXS7hiJ809lk5TWplp2K0bCS0h8u6+Ma+cWrMeLHlHb9+FTf
AF/F7WyX8rioeCxQcsnKviJlnA2E2lhUieebs5pKS5oSjxgx21gUqTDI3GlQyHiV
WdmASXPXM/JHAuVEuJOu6SMexUGksbzHE16jeSce4NcR0dCS3QZ1oh8iVlz8I3YX
+93yxEPSIonM30bGGKcw+8y5PR1KMioAYX1iH9X8wlZZYeE6bx58WzAQohA509FP
wKK52bJUxr/YvRnzboR7Q42jgw0yNQOEq9I+3q7gvIIGrgliVXZYOWkj3cEfOwTr
Qav4CDHCmDTniVjYWJ7RbATnvMBZ/8a3ZY0jho+MWVyjwxTuRZeeXd5nbG53885m
NVWB2aj88/zUaAvqalqquDx9qWPssCsqWIHNLKBXdrsPQx2ejL8xUTqPGYAx/PPk
yLS3J/sRKMPmtdbZ+hJGKC+0gwGAtVrjEnhxEVw/z2QWY8nEA4K8q9bWgjJhDX+V
1BNh44sHJk/WldE+NKGslLIco7gpHObDGmhvOsHp/+Do28wzgv77cNLfGAKu3ipv
/fD3UWtqV3HEfrcPt6ZjQ+8XosShfVVzzD5NjqjQTGQihx2HhdK/pP9f+VbE5UBa
Sz24W8eqX/QK7j3gW291i6knZFRj/eaA1IZ0WFwmRv/Hj2zv5tCDZuedOrTECjD+
LL9DFRfUsDi/33TFNnNch4PAIfQXTSK0qChRo5h1+PAC3bsKsljHgYP5gqqSQcsQ
yT73iYbNW73qIN6qN82NffuC3kRbrb6ziELGR8NwYoBwDwJg60jgTNUQYIy1Rl7G
9kN9YuPMfRmTL8Vv4jdeD8h5Ax2kRATz9DNK1ubLO8yGtdKTM6prdfI5vMi1FeT/
1YUwNrDjlP+4m8NqUWfidQbkOeeKEbBgHVP042BWcDStu86vY+dD+p7Gk9VM2Nor
C6rBxTn3tpNj4CbuJuVDzHFm9UiMqu+EvgezrEGEiA4ANZnbING/OeV+rf+f5Yna
cRu89/DL74elJoY9MShqsvx9/mGvYL5gvx2+t59LBoGHzEna2U0SjHJIG5pbDvfn
YKI0Iti0TkPVQeh5zgXeOs1Q1z8l7w64oBtHf/ROzWHCTViihaW7UFgB9ClqylHg
tmxY1U8YxpJEDmtLLSzj0vlZu6j50Vk6Y2X6T3c+CjnwGLcnTzpkW0xRHhN7o4kj
1h4BAJL10YxKW9HH98NYXORX0h7ADm/MSlZRvX4kB3NkAsPOVmK5WRWFTZ+oRciH
Z+hl3TVJBplR+6j9vbVaF5oBdLMoORuPejvTe6H2ApJzjhjYRnGY481lIy1vbo6S
VxIWEM+BSXFydZ/aTxdoZHFDVkD5r+MjHqepPoypC6zIb9zrcyc13Eq9GT8CICl5
mrwQy+9vG90o09uetPONcwm3u5xX2J6AcMAn76r7vxQD7Wx+nL1eo7HTojROUvMD
BlhF5aJ07nvdcLPEkP4+1c/6E1TGB6I0/w7tUQtNw1kJhBZPwgJNInIvFFe1NTVO
vx9/sMVNTOFp4Htn53DzDMr0VslPGGZT/KeNoqcRX9AAg6M77VvhdT/9BXUKyUTU
/9aNS1jnwdAyhhtgjo1CwEesFWskY6whfKURUnHfLYqhuvQUCwdOpVAxhdHXI8wv
OGYFHQSzMWp2xoShf5trcZJbly288l1YCcTHYVdVnPOZTvH6+DY9H28C6fAF7PCJ
W3S96cQdi2hgskcJesP+Nd/tpeWqIeeQnvsRtPfjKsLLzMKi59RRODvJYBNOh5zx
s3tLPAdOb25zny2UCXVFUNXYrikCYRJrQdQaCVe8yWyioIA3ebOL+u1wjL2SMp+L
J55MG8ptpqqXoBZsjbJHbsEJjRwfs6xunaC7py/nx+LosSOtZKa1jU88TbHBgsXk
Wv0MI8bJ6AnM2d/EIP79IOJKONbumwc9FWEiLMoTF+4SZ1USQqI3cpPEJKrCvvn5
5pSC1ewtZ7yNwUCBPBF+87gu0yt4AIa3hL3O2Dhgtt6v1k+3vjabS8QISdc+QHdM
X3gawdviNqkP4NdJSWBS6il8frUQZ8mSMw9ALjhc4SmKasDEI7EgPwi3+muMfECD
g79TWmgqNL7TxiTtzePTOIVNXdX60xPsPWFgflWSuPOMzwoIwfMjBh7PWF0QwR+P
OBYBMnCTfnIEme9D30aSv2PR0G/w3muKpsDqUE5vPtgjIPBEJp+dUROTOloFe+w8
W4taf4Cfre4txZRgrvl2J2jNB7sR74hoV8hFR+eRkm97LQy3xLidOood/PCW5H0j
GuBRJUrGVlaLKtIUAz+5oOedYuv11OvJZIoILhobdSBe9vutLv7OwCWPqB4whFwu
A4HjcwuUjTHeFX4OiYPeWXidgU0UZKxf5QITE2fyFtEyxE4DLPwCC35fKSqDP0+i
eX5TPeCPOCA+DPTu4De6E1qKOEG7dBWyoWE82KKekzX1/kPZQgbRyurAL1tW8DVW
AU9W5heAet0c0WE4B7AqkYk9GUxHbIAMfuUNpbjPtz39H0UjjaqdvdtS116Pm38r
N3w65BcdTtUnepqOJLRwocDPITABu8VaN8SUB6LO4dy5h2dl2XJfE8opdTnLUZle
L1bndHibiGmb/vsrcjK/2L90qmnMv+yAgr7n+VsuY+amZwsz+8TdZjtUVZmo2vVB
PNp73EdbUpTlfpkVXXt4OFrjUQSAgsc8SQiIgq5PXc/8gdtc9mBXNyf6Q40inq2Q
brxPqey84+GmAxoy4P+xLkp+nvs7s5E8DD1th/7Pm/Qd1mnRup8sDvQiNmKxjKob
+lz4BwHziznQfmk4rxhP+jcCKCwqYzPcyZsU0iAK9OPxpUgtWgPccX1dhWpBy5Lm
N/gNn46ZcG+Lud9epOiuohhV/TRuOA6+nSrcUNsYYnZQl8Lnxul1Cn7N63OWVzZw
eAGH/RNBY4JbWqNxE1Dpc48zVY/Sa9vmr53+s18FqZ2N8hJclac0W7ZbzAfwLypK
y79MZobx7+KlK4wJ4kPE/iDvlEAs5o5+xDKkSqjJ1OgbQTvMSliKnerlB+58KWYP
3tMpAPOPxkx2qeP6Jychq55rLco5qzA7/wFvGlckv3xX6LvOWc0TRqUWFDRgdExu
TxdN7s7DkVEEMNkaboLJ2SmeTF+c4P93avOZbapwsJMHe63H9DBiKTc9XF7bsUi8
UqXnouhf5o+BCEQJYaGG8jeW2sYE2mryCzQ08wIiFu1EGV5lG3GTgv2cot7TLRvd
pfNtxCICGqnKLl8PR8H46Y17RgFCRQHsZwEnv7tLrkKVwvtzLA9OZSJgp6QiO0Ts
11HeqeDTRlpiz6t9jbx34wkeeQJOrVtr6a6zxHJXQZBHzXqjzU/AnJeenMhqRGmx
ybQ8CqctH5KzMW/1kMTE2G4+e5L8vKSk6IoFaVVtI7KVZ+yPG5g9V7Nyp2cfOEy0
NyZskrk/PEtxKoaO6VOvSHjiMcGAERXFq51dUiju0QjBcaaRxZWtWLdFe2qO09di
9CUlp9Mc6nZZlbjjfyXP5yI5igHG/HQcokv/HFQWGAJByNNhJOhS1RCeJLbd/yxD
Ua5xKc8cL6ZK3sb0vMV0bWZSK4xjjLFWm0s/nvmNx96UiYd32dxDAePVAw+QW1vl
eFC54A3cVOe493zl8DPO6cbHy+a1mEEp1SZU+mlVeGvY3SIxhOmtcl04deCDxrfW
0uPv10BAtC5W+WIIjRHYAlvR8nFwesknGehlwDmvThQX52miG+E9y80cFNGRkhyq
FPYuOqUmiqrju/IthyOM+OlLFdTWb1RU8CsY45XywrhNalDJ+w+IfDw1gZvyycuB
wctYOieyGoTU0ThSyMoajHMofI0vjkBP+nJBeuq20ALUvFJvBJLk+9ZCdVraeqj3
c/RUPTsiofNdGifdUrBuLov3jgpVD6emTqWpSVUy/xCkjJIttwYFNL1ZEufchttS
lMP41OUcQLwFJVw4MkSIT7tV/ysoKh1QWqFtzQ+1U5z643tQLaeuvXOPB4zCviUH
defr3ZEcW5vDaIkYkXw/KK/it/wVwJqLI4P+cqMmB781RzUfL0lUPJ6pB007uLMq
w6YnMFb6SQIoF2jVb12fYAFGMThLhICfxBTHNQ2+iaIPDmMEoiT6lzFURIR0SB3D
3YfPVlONdI9nHL0nhxXNaIrX6q0Y3kp/4llvvSAGYRF5A7elLfcBtnEngSCGeUbp
JmeDMUOQWV2uCVDgZzBcMxq/aVTeYEdjQJDrdq9ubNpn03dFlKIVpDnpjsFPzmD9
vxa9lkHZws1V/r3O5DsxJ5rikZSwhALRxA1HTpu/TjItQjABlouTNnO9S1Hysvm0
eT18LvJaarj27N84n1Y6A9UbnBIVssebHD1+2N3Z6oppr2u1JxozulTtTILhYzeZ
w0ndyHUVrqSGJmIDRCl0pmgGGFcuiAsXz63BnZrQddhQ7HQGyvE7H2vSAXnCHbZz
brjj9Jtf+W3nNug3Qm/wp4DMyCFH1ITKWwt7iKk//YmaVr8bXF9MPmrF84utStSb
Isiy+5nWG9KZx6wDrJVcY5z+l+edSCsRX3FMj5Eeprr+f9kvzYq9egahc0+cEQHm
7Mdp8gTukaXkf8gEa5IiACsLTTlJPlQMKNPTdDC37IhJ7qM60XR8tSEB18h97YjL
GShtGZQREEhLQO6F8YvpIB/ezUCVNX0FqIXC7/aWtGDvWq6fRNfBvKCoDJPbm2Re
rMlGDM8ywOaREkaY8Ek9EiYJO2iZbliE0tjd1UPet5gUw8qJmVlgCe+SXUAZJWDE
GUPnl7GJuWcbuwCWowbCFiLpRnyYPqQJttwkegkEadmoFPXxOBNxyznpP6l3Tsip
dU+bctj6fHuzqwjxGUdOxx0KPuu7WCIlsFJFQ/1X4oDwWKwECQEiqa/1GsWV5dFb
h2Wq3SIAytHRsBmpQUMNLyK8kId+rQ9uVGGhbheG2Cyck7QjNYYKDPo6/21vA0FG
HGbKQYukmUq7ScUjQxoW1C6icGfyN7qiV945q4Jm58Ktl04P8EMuct/WXXejUhft
DsAkc2iEvQNHjyTdcYUOrBbgtjGdHEeeLlZqSYcgpPPvpPmnp5u2aXJxNSi2diyy
T99JPmu+xAHBTwoDtsh5RumwEwbP4qeUP41VcYxmx65djZQJ0LrDBbuNqOudWNZy
+GFdQayqMeEcw5wL/8KP5Y8VGFIiuc0fJCJfViZbACPr/9rGwO1FZTdF4OC5wYs2
MBz/oRPgLidh2AC85veAg9ahlmvin0owPnQn8S18LGDtZyaZ1aleEIQzb74ag7V9
Gb3lDMxpTx1Ku+mCYTz2JWoMNT+iGddj5JqeVxN9Q0VGHpnkY6o+LnY0H2oVmGzm
snl9TQkmoNbzLtryQZ/njJhc07in/9OIGZf07Pj09/x1EifQFMi+BI5KWrh2JP+5
BRTA8EvYhoIAIDUl3Kq+mm4mZswfp5VjKOiFXzybkS7eCyy+7mE0cKByXDAG3ACA
xqfD/HqprRb5orrTPPSQoxAGotq9Klt1csJxOlySBPvBKEEVqcjlYfGmDslM1Pth
+U5G/BgTKaYWcgLnvtUu84oygI4xGaY68HzUrEuv1xwRBw6JkeZGhmvp1eLzjltm
XSpbUBLdegwsblcsUGksJSrqxZ0cE+edrwOvV7iu0eE1CA17Tmh/9KjtcdIJ4Fav
fmmlf1qFW2I8tM6K6jTm/YKim+p4qJpGNHpeFX0DRz10Nd4VJnVqPH6bt1RMsfxy
P0l4SzrOEkJfH5pTbGQijnO89/adly5IvRadk9d93l/z0gnYIS3ok+ihin4RaArd
tOjtPNnO4ggSewTNNw4uMnbmuDB3Ox7ofcjDV5SPu0vN44cvnhY02VJZqySl5ksf
5GzKZTHFI0lVDw36FRHp15x1B2qY8QQLQ2FJyX9wUWFoM0olHMBUMY1ju0LM9hal
XYtX0sZ1+HzIepsxEtv/8GAP8Y2FsPVTW6ajgTTSpLXnd5rh6fGanI0UA5WEdQuF
FXDMQyiBkv0aoJp0z8ngiO8ka3j9y4dgH/dD18lSGgZrlVa/Fl/NiarQqPYkjHwx
fRzm6yPEtGWy1HKDFN7EQHkERwgHGdLKJ9Vh4jBhwqX1nLoqlQhzk02J1/C6rnpf
fvchQu89e1Ojb1iUxdbo+Pesx7glhAYGI8HH4AzmlwHlAozq9pNXBGy4vQ1GVWaa
9gSS6jBw5m4uuJgLruhg8f/c8iilBiwcxlCP6a0d7rAWBJczaUpTLy4Iimknz4W6
afriR2W0vUP2oQTA7igh36KaS1CpP+W5x/kG07ClD+gzyGWp/vDK/3KDOhL3has8
K24UxNAdVvSF5TNrMTgpHKUG0du7G6qFc1PdLnicJWD0+kmzr6EKjdXih1xk2EYn
/g/CL7Gj3BgkT/3UJ7hk+iWyvcfsgVReJhtfSg5xIAMttBXEp8VLFCbiRsU10o8s
fzcSnlm117c8oNwNXAOMB6uAKtnT5ajzrFbrMgnldhEzc/liewva8zhHDAj4ELaF
XC7a0xbeuydfiUM1YCFhovcw7RaltFQjrU9lcVBHOPAIAX7SvrtsEaiRbdMl1R6t
ayaGVk/YesJd6p/38FGH4YJDjWTZS4tCmwZ+1qQvbNCXoyT1HZWwke4ETDBlR2ZB
wfen2EOM9sf8OnS98TFzVI/x1wxgPlICHtcWQY7ZAXlSaH1/xgkv8PuK8XixWz9E
BuYptkgbrfqu54fy67GjXPQyOsNYWORtJzet+cYHKUUtmUojmBISzD8OPZCInW6w
VF9jvBP1EaxYQSVo7YblJbfpqskyp+2t71JSyJTbeqMO3mWVTBLTAeVkXrX2MJC5
YVyRfYtbhQ2X4Uz0HVNecxgBealn/BVrma0FUlzk7odqeds29cyUfobhVbxnRDhb
JjDhIqqUzXp5bP66iAFSfW42Ksqgj+y/3aaFTIFTr3tfkCmpbPjh4IizJInBAHwZ
OGwmJab2QXRlLvF7NeE6UwIeBfjLvheeRtEhzOMlEvtYzXe1ae7Iz6UIleX63OEC
4uW7lmidQMbNw9vDlB3Wo3tNy/X3HdwKzFB0VilDZMDqwkyE94iG7FkF7Q9i4PBS
kK8Q//q9hDvK9j2lhe+w/oUcgBhIdrGqosjki4QZEYpQq5m/PHRbUboB2orDs9Yd
0WHUe3szNWprwotTkKJ1VtWEOIskkgjvemNoFGTBVa3yoS7eacdyA14xWk8aQQJU
Nez7NCJRR0FNNfUxmNtTCCbbSWRjQyU4KnDDN1GQqa6960s7uZXzWZAVCnMnHFJX
eRpJV3qLBOKXhJD/WC7HTjstm6dVhU0suGKnMar/NgT8H3vTgLFA5QMaNXbKAP02
txRjpPYs0uZ12K0Eq7Fc1hHoVJAuiE8JdfoB9d/7k2BDJP1mGbXPu2l2k+4PzQKs
ollLopxTX7csWmkB8Wq+bIVeEMRYYmJHZNTDSPRsgGLTX8OB5nHIrg1NvF5tYB8o
XWJLEwhWNh/VY44pD9LnUcJFg+SwYTeRYqBMyT8waWUFKXUmZlgkjgMqXNer7/KE
DMqFYPEEfrm2RYKCrtYl7rAuXWoLrSpBut2Ks2Ice/WX1603j+qiDZGnZQ7dCEYU
yVTvG/3ILtxbHekFf84llgBIoJaIcnEfYAK00BJZp1kMQrvMmgAdCXECr3UeGgdR
qSJYubhEH5/AdCuAR4MAntzYyytphZ1MVwMdaBHHjjznq78NTMzFa5SDwsV9MDW3
QXftJLTQHoUyuImDxiBrZ25IGXJAcANPZqdQIgarNNRzWFZcrRfJViHEVBMxikcq
c6//r33Hmr+bVH2KK+0CQb+VNPn9wg7ObNvPMCE2SdpfFuFDBRHFcQc6hsA3yrO9
IkWhbOyyGww7u6eNC6sV727l+FI/0iYDWQjp4n5zmWDxsTdvyAsvFY6ZvxoV6bMq
FL+M8ixiHYRRyc1VHd4zDZEfOcl0OD7uYgijMvriugr/P0Hk6Zz5OpzbgXGNc/uX
9OroOaBhiJjUFz+FDmBW+2qxrLJ6mR89Hfon5cfSPsigHxX0mFJ7PYXHN5dnyO/W
gHUJeZQWItHd+QNlmJI2PDzBaX0nXAIMCqcLmCD/HZhU0IuRYDsbEIApMK9lAyaS
4tp+PT8rwGkDyxG8x3YDE4mWr8qoOCwxNCyMv52ZMCcIFrrZtqGQpM6tupakDCxv
ArGjxl5DsSjbMakaABjFaISN3QRW1iOuPrzsCkg7pQHEtsGtV6GeX2VjsidpQANT
QgYojyT+YU9kOK1UQgi8Pl06zQFe26ESM9ce5Vsa6W1/npAorOdiUVuddh1uOMgk
8ElmTTc9Q/XoFvLN13zWNhvwUAzkpmuF5oBLc3ZZo1FnYmMDNwpYeWEPgGcQAFPS
mTrndntfBX/ug6deyyhRnG5xewA3+KbbZTYyuqK3OVwdQdDUBVIieG8ze5wHSLWr
5fWXh6ypzJi+U09XqsmWUXHFEloK14sTFiyBkSmgE0wtKPrgkEWzuULmZZTOQYmv
BxuIg++w3wIm6wab+SS4I/KPyscoFkD1OA2MWFprt15RnvCvOuYlRY6HAhc+celD
z+lRdQJR7ZEGfJXC75SdqkO4i6vvam3GFyJDQli3g2PKj/OAfnVw4Z/6KdcnmgnP
oGWNNrA1Fsq0WVbMOQ+FGRQFXpFPOpZ7+COxmtJDn/4PPq961N7lbV0OCQMvUL6E
CUfMcUkWgiD8bmrhS8OB6NS60ZIM7mxMlusD0Vnxf2o9PnAPpDZr0OC5FBc37clQ
8H0CnE7qcESNLD0GpP2wer8vxSVPpe4SeIoPIlCwruISR847Vrb6v5jf5/3ifKJ1
S6oaE53wMMTAGc2tckkO6MY0pkjia4+Wt+pKpOws3fPyhBetQlfq6lzCEELd2z3c
JQFhINrEWtrdBPFF4ES8AaRHjrjMlbwQ8xrR5TdRNJssB1pkZolnb9qKdj2/9uZx
3okES6YDkJqC21OiyS3XDnZgUwwGXEPyUjtQTeXXpT7wwiHo26ZWgRFHLQXFmKzE
fzBHdMsIJL/MD1+Zk8JjnpV20hGsHikdt1c5lWh+lmYzhYQkxYbwskmvLZAVfmy0
D4civyUIOpsOoahJ2JYYEUMBaho+PtJLLru/hLjyLsOvzAMfrYkPwqiBDMP5fEoa
zb985B2ZWkmvGs2gVUHAjEujmb/SQsHqWnPHlsm0EKvvU8E9yLrWr/aYZ8Z3Zl5C
QgUuhQUYCXw3ZHPn0Ky1AmMx4P3k7Zl0G6x/MwV82gQj1g7MwwD3r9oPXVqj2JSj
WZyy3o3WjrltEmTzWFnFYrSR7uOHdN7DWjCRDr9afQO4AVYtU7kMDRtkbpnq+Y5w
ISI7+HTdxQ2aiOmNWNr6iQv0lkxGy1/OgAUhCpbqANi9KFrjnPudHCucIF3p1oOx
5zk1XV0W8LaK106VacEthum84TGDeyAjgYYZfZesGRVoHFjf3hT1yRcRRP4ZOC1a
T07rO2N4ontFnDKt/280De2vKgkmtlEFTAhUTeuUGa2/Ta2WBb1K/dQyJOkWRFns
nUPuC41NtVknnPMxg7IGmYJLhWtvlw/1YPFSaXjs3n6Y6LI48xCyP9QgPdLWfWYO
JdUDd8ZBGRQUhNCeJmH/068eCeHCJ2kgSe1hhJU/oO56AFa9OVlEigy8RjAOVvyO
h+QeHT29Hl4xJwkUxfALdj52h7GHeN+Qm71HF8KkOMfqWfU236Du2pqM1fgYnOQO
ylTQ+3OAeZdING/Xfgt+gxl/hROOHdWOY+xpZMk4bbG/Gbl5SgcjtOILGsX6xTKR
2mSN8YyZyhFJTJofq9/MqP7JA+M9Kjfr7FsaXzPS40GwY1gpTfFSQYVEg/uoc3rC
hNOu6BYlt6edPku3IuY3KGHd6xjAUfR6KEoudUaPL6eqw8hYPS2A0/TVRE9UhU74
EFxgoxqcKUQPqcm20FpRojy4kL5k0Gg7tifp/NYXuiVAun5JIHpBdCIPQ/A9E7xH
iNol5p7lwXbDLH8ApbVusS29DifWxoeU0nqOexpbCL/wh8sfCPm+acm46X2Ix3op
CRzRg8piDdE7+bJ9Odeq6ricODlmix+c67xOof5ifjE4hED+UXIJiJ585emEb859
RV4zToVM32mcX25eg7jyo0d7OQgshoKzw0Ugs7pUcbYm1wGQAzaVj3mp/rRHkzXg
62QGVaZb9TpB/fcRqbDeigNRFkqgbI+ZWpBHCEY8ad1Fm/FoXUJaYned2vnWF3GZ
FN2aWuQCccZNZej1VsDeNl42Md2eF2N8c/JcmiQM3dAl/MTFafEfjWZDH4XIphEO
tbCa2cyH25JkzAqsmr4AcfwqMRy/E2caTCG7boH6KKV9/CHLFVr4pHMlJnmnA8zh
RKbKHyJrpJonCyD3Pi2nR1Iv9isXkOi99joOF4cCJMa9ANkDZGPyzV9fe7iyrTGw
N9dzXiy1eyXE5temVCQI05ha+aA6hMMe67lu7hl7aYb2eJbww1YEC1eSM//TSARo
4hkDF4aZREFsp5tSK25mio6n9QFmVSHVF9IGzCKlfHM3x82OHm16hjnpm4uttxc5
Fz9KDPbKhlZIib36AyXPubQPV8Q3zR+uIqoIQjGqlEDRLzTllHIq9j3bFtMxGTYr
OkOI+/zSmPDSpuplBftPgBVMRQD5TgGjuZXP7qdmYGLBQsk9KlxJX8gCpLdA6MUK
i/shNEQ3hOOs066GdUyxt9NOAU33ksme8x40ac+NdhU29BkixFaRxn6Fyv6W4DX4
6MygO6AifcdBtS9kMKL4sQhXQiW6454Ns4PIay27V03CwARE/BY0mngLJk0sqpia
vB/0WdnBnTq14qNhh/lZ7U3MONo9sRrV48YE6uaRh/ozDm2P8E4f/zzJxBhSiwW3
q1/T+swVds3Onv4j+KYfL6ferirH329bBAgQnGhBLJIMI3XHEn/YyUOyQ3xpd/Qr
MZl7D2TIINGtJF0Dq7VZXJ40/s85uWO9LVC7BWl6wG3xu2Jg5dLEsUsVTSrZlqKu
2YVZVpJf4/BbRFa+znW6ZmDdnEXgSgs70dsajZ7pom4Q2ZIA1ufFTRWOAtVBKhvH
/xwn9u/lKTt0s9VMMyB7uEA5ESmv1lAyYkhYiPHTwumXukyPMEI7e1EkUIHYYEWv
LuZnxRc4HrmY90wOMOcHuFzeNZiBlosbHDslZ9pT3Yzq9cWXqDO8SPPfWV8YIrrB
Ufj0XWvLrabiQdknLLh6Y/ujRsvGxjoNMegkcuY+z6W2w1J6aLzU9a6QbURx9O0m
PnMwQuIfaPZN73XcCw4SfFCPsvGmQKdbM2fUyIun6nvF7ssrL2IjjXL2HTPjuJCo
le1jDIi5RaiyDFAj3Aeqx9WzyMuyV/lYeu2Pqmdvp9WXrUVTB+N5lp26RuJ1thXt
ttTTL35uFrU20cIYDq5fOWpFDYR+ZOZ41Cx/bV0DifHJORtei6FOkJ8jFirJ2cnb
fexLoISVllUv9zFH/VU9VjKhiZ2nyFbibB5jGZ6YvmTtk8eJyrEOwWj3WkSK+KQq
mqlK2D1ZGqk/3VwawPfebP262zwXuwnSIA0+TBRVMYoWCrJDlcHmVNPjFxTAoEmC
rh8g1Rfh6SzgUVjszV+lOhqWc5BJ5fS4zQlSBIC9j62dQpy8gARh6Xft2OOa6fdU
amTuyIkJyOg03TgKFy9WMVWD2+YGGlXgOy28hbfP6Ogdo+A4ekV7X91fqkS7M9xc
k4UFSz2F0xBoD0tf7TSif3Gu1qDwgEIm+vAFqFYJUIHhGvqReDI6lWkMgZbKB7VA
1hwMClbpnDYrf0XNO40yzeAXlnBfbMiyAwmKGd61puN6La5ZMcqxRP1pkfjPRj/Y
2197vESE/rJ1ckRS38UbLdeX9MJsvlAifcK3o+NhVIzhVBe7YSUmDIs3wBzEHVrp
KOjN6Uw9doKZZCsXGfs74AKWHS9BaQzPO76w/CXXXfr9nw7oYEcEqUhFLfBKb9F5
mmxG3O5/PMTuS97oxjAcHGb77KXMMwTjbAYinbq47p5FkaDKPH+pf7eBEAj5EwK2
RTn6VNHzIbxh0HVHtVW0G5Zd61d7UHCp/kjB7XtSspRsYccQtQyICth3LHbXYg07
zK+XD52AdS/94myxjCrmVJ5lee62WOVqsfgXiT2G7V6Y5M15G73645zNdQPhRjjJ
ZoiBEmMF5uu+t2433FuJr2qrkTugbDnwSny6cuvcEEPw6S4uENA7ydA/Uw1nfU1I
qs5BdlB39bvSi8KBm9j7onFbQQijisGBeZFgHbvcF1xGGsI5ymegjw8wZP0Dnihv
eJ6ALVr3Vc+4F+TSNJEj7OS1/l6enO2bjppLbu8CP6y9XrF552PYPbnm3L/mWDS/
LJ+i1DUjPKSBCU/Yi8LyHqxgya/3t2ybjWTvaamRKyxFSal4mFJtF6tCoypIivRG
yMS1wfg17I0J2sq6mUVu4FRPWUA0mcueoKuWzeCo3jllsK6om4Ur+RgTvYpSt5E+
8PFPLwYmc9rH6gvsf60e0CEw98gCDFeRi8NzI0Pz0t822q8ZnATD1wz3dRt3FNUY
4TjJ3hqavzZOQhifMgubTBKibIkUqssfLLbEzXf/RMzZnPfsE5BVbw3AzjxjuGLM
xptCsDADTeols2vC4CEOzBDLPrPxQJWNJFmwkFcKsqBrx2o7+Xx5TD9xUJEOZVBi
CghQNsvrbpPWqJQUmgYt6omZFEafVUzYOzSAujbVNWd7q+uJKW1BQCtMJMsqE7Z4
CrgmOHayAvbTi4GGArzyKbviSxI7VBwtzO3qiXRNY+Jehzo28mGOdZ62lw6Zs8Qp
0vPjeJ7e8M1K/L/XmU3Hlse4CnWzEsZPz0mhf+KaZ+lNOQ7wX9Ov84VuH3Lzjj01
+B7/wm9e5Zg1EMT6jkJeeorTpUeiHQusLOCt5xlWAJxtDS6EFT6yyItalnF2mcAW
sJBOTRmd/GCX4pk2ryj5zX2jkDZ5Fq+VWJmJHlIVsZb/Tw7gypyKoeeMP+Lt5UEz
MV5Yb77WUs123LQMQf1QrScJUOzDccZbd8NrrDHHAmWNw7ppIiB3CAicB2HL95W0
GMVE/ayVh0MxFg9I/hcnkQn9xUdmQZl4e/01PdRIxhL6cw1TBZfn0TJ56IC/DTe4
111KN8OVNgFBzOVstKwMzsz2cjvhU99oIEKWEgSUmi+tcPs3H/st9QKB21uDzugO
N5UVQtRfRpdePjnBWze23jtuqHAuO76Twqw5XTYr6WGX+GqRFynFQoADei0dqY1V
UKPU80YXJn9hoG41bfdJHKjpNzvV5jiSMjR5ERtclfdaWQkgOZKxxqS1OdV0CZNM
mhPKWlk/sMZiPV0XIctfMtHbM5ag0sXLm8z55S2WZox2LoCH7wU5Wqz+z1LO6pIK
jFAxf9NSxVIRKOHnoLsmW1qOLjs3ze40bUm0GJZ9+4CGW5QxMDA3DZ+IUy9/8Qps
Bw2oyZn9BVOOpTPDS6+95kiiXxELtyYiPTv70e+48HAcCbJSf3ubmWtmx1TuZfou
bbSHJEJFoKQnky3TkDCiYOlqX9P1kRjJn9ma2yrJQPM/diz1J3kKC24NKy8BqaOR
UQO0Prm+cVa7ktaBhwBDH7yNvAcs2U+s9q4hTPwhGPafuF7x+jQp5j4H3MDvCRH2
uJ7LvbXir6fZuUtyxeohGvJqg5I5Q2crMA61IU6Rq/TiLQdx6wG4a+s4EM2EGrqS
PvZ8XiRwZJFiafNDe31yNHFhTEqEFOYBnN9OSo/4shjgYYq+m5kiBE2HqKTlYPqF
CQlYaSYL1vFwx+9N/sU0RgIUZQBPtgyTW+VkUEap748aZJFDnhh7750y1gHRZ+8z
0wZqvMpi3b2feBd8smehItf+qIKDEwznfUpfobGfU79xQemjGhYDbncx2sVyEkHb
woSTUCTTP/uV4Os/K/FbqQZ4hjDR3aGC6ppxlFDBmTkon9pBU6kNDODmjjnea5fy
VJlYbEScWxJodMEP3SnCbYQhD79k9+VY8CteZEQCeViWsp6on0N7YSF1rAO4PHFn
aEymUoxsWjCuHy8UTHyf0tEV/pKcJAgxPSMk/Y2GZ0XqoZipR3n48LvMZrN1arI/
z8Wzh7ycYP2RXdCinF3D+07+4jxDBn74dNO/TxPhx/hKI61MLULIq2MJTVyTGxxM
/UXFXabVsl7jpwWOHfGOonU17H+x/R54vVTDA9H2s+M4kVsRrHwidgmzswpJ8KG/
MKLCp4Wg9hNAvgSrjHTDrjhH45+pj3Nai7e1/ER3JTAdup2HNDzrI7SpBKlMWyqG
FHA7VYugSLjzAFsF6APqJGScEu+tLI/pvpoQGFPYthJXkLWTcmFhMDleXFzHtewx
KBnf8ewgdqaYCIr1OxFwFlVjc5nd7XeCCKkhlPf11xwTbHhFyd3rjFPDQ2199mM4
I2v7JX/kiobA9X8tJ+VOlG9GJROblTYRcqnhajcNm0Y5SYqY+0J+JnlaRpfHYXuw
Q3IWk9YlnJLxXq1+Xkd/Gfn+W1kmYdVm+I8cq59T5gb48PwxeMkbmj//WdLqu/20
O0IZ9nFtDdwDn+A999MdW6hHCTwCkV9vGKELydvQnHU4NQITSoPGY8qRypp11NNM
gGqDdf6irNuoyRZn0midJq86EQKnTF971V5X6EFb+7YYa7wt5f3yOzV30L2cjgTW
4LXjATnUFRcmB+/27loE++x7jp7IlJbMCzFsspFa85zQjcJO3SrxF8vEXjjJKfgP
DeW04NA30zioA2eA4PWdXIe0tuZEW+7htQV8MBmPUgDY+OVx76aBU16bfoPC9NLK
+6WYFae+ofc1L/8MTjDN0fQYRVVpw/9VLhv1tBrnp5py4c0BPE7c7zm8TF+2hJTt
98LrtaWjEHYgNQLkOH3jQfBL4mxe9iaMJLmySFmK2ds5YuONUmoQ6iQ3+S5F4VRE
AYVSzyFBGbRGUgAp2wG73Ted5GtfaFwjqP4ug4ekx30femsi1yFoa7aR07KajbZn
T98AJLIHlvnGPyNK4lkRgwD7kGJsdVLfdNxTaJOlwzveXaF74sWSMOdRf26teJlu
NF0vC5+hh8MM6BeDAy9f1thmE1mIwpclxSdu4N+RrNjfQcGgfZciinIa1Nr3kGnT
21CplSA1rzArAzHZF9HhvPCRvpKRb6FYJqcHkxiEbIqOuOIOuZ3hMUwCdHsfwN3T
b/DRwQLgY5iPSV8GMe670/EJC4wKxBF1IbEbjir93B3Ia84P8Gydxm25QPkfDGf1
ZTKEv5bZ2ggGSh3N+KNBJ8VnMrnHZHwIZVM7jIQ7WCVaGMfsIT+kOJ6bnjitTSw7
tpnNOIP5q0ah71ZSv9wYA6lgabXSTjcPNl/2LKXZJ61pgdEFA5BATMcDxNjXG6zi
VcG+ODA03+x69pauEm/+SDv8vM6jSahlzwpoGH6WVAvg9k3RJzbS2fUC4J9N1UCJ
XC216SRvSdc3/uLhOctXrNIWwuH9QzMjKFKj8MBx35wSg97mNmNWbiIeoY0UyMjL
6/NBsB4WZlLeK6LgyuZdyd2np6JAtlSd7hsD3vzIWHb2H45oKQqY61dEeVnYDwgX
/kZsYwZFYVWqo7AuQERxnVp8t8KSIDUkjdDTJBtTOYQe8rSJfX+3p5BUjC9LyKAV
VmV0WLRUqDOvfvBFeLfufnGDQo1nlwUW5LO9TaI+42U+No629lVeUMblEl7AJvMB
H/fJZsx5Eesn9nFlv8OJX7fFN1JLvt/HkSB7va0ZqIG4K0IF1gElXic/nS1G3DVu
3QL+yApRizGTDEq/a5z+V49dHtDIL91SKbnsqRafmJQWCZNhY9aie8cSdf62xJPJ
hZV8NL9U7LHU9QUu53/WeR6ycV75MRtAvtAswkCaeJVNVaiQJ8Ok4ODSYgRi51HK
l6ALE6HhkZvJPmw2bVuwjFX23TryqSw5mndnP+jToTochcUp10Hl/29RvJlYkCoJ
VO4TxxdZQAW5zhhqsfur//I3GMgEjwG0fW+LR2hxEig/6MIxFHB+A4/Zn6nEZ3N6
lxhjxJvHMMUh1SOSNCJ1D7fvCrif7AbcX7nI2jcKLtJZ1AKEXb/n5jBPas6Dw90K
T5R9UK6CyZv3Mu/PIDIarokJ99WWL42imoGFSvELYBBntj3M/+vWCxUf9d3PASiY
4SdqDnHBVi3CoxaNFKPuV4l6vFNnYUIf5G7BbXTx6AamJgMnQcsKjpU/J5SxVOaZ
7w2hW6ZpzwjtMZA6XKRsdpBJ13ZVYTD2HifmILhVtRjVcy6OzJssywzHcEwkohV6
YCYTjctIgsy0CECQaz/1eHTJdn5nNIdYEkIF+3cF+29pccpalzED5pd3vUms+qva
PJMCM1bo/mDfUGPvcTopImh5Utcw01WxNVNMNicGKxaa+sERsV5v643lwEL6VTMz
lKI9s2Hh5DNMmr0IVKJCnT3enY9b2Y/ueyxyu4R+CJxc8gU1cuxt6Sb+xpCDXCdD
aV4J7EqQ2yPELIsF/Rq65YHZcPq8P4BH16pkE98BIaEfGXR5jePI+Jz+tMn5OURu
bkEi9CWDpcGfC5mtNGvuvREurn+v6nDEh8jhBrc8GyIrlbgaw7+j6XtdR5NN/rPg
TjDXAEv3qw3k8GbeS5Cn5xPiR6Ycz/M19LjbKFiKA6s6noo/QeDbhC1lUFWo2kwQ
GE6G2AZaWEEZrTqRs4w4NDu7vgLLB4W9lEn/Ha6OQt/h3nPr27rU7IOAOdAxyki5
V9u9FF1ijbnT1zz6+ZPtG4bx6Qkw6cl8Mj/iI69E0qHK6+TkwHG86yPqZ/It4uKb
CDIDa7IEGWOqXfDODQ4ZGjxrqdY5FfQBbAJrpmAe8DoUC0K0eAp0gnxn2PvrODCn
h5kyqFVhbrC37U8nu+MEHp0mnCDhA4855kapJE+rOFRHv1QTR2qMCqsK07eNY3TT
iOmy0VOgMULthPrxHwjcupDrvpBj32Y2RUyqgbkQ3IGWsBzOQDunqG00v2SUYXxN
34F4T1sGRz4Vpb/eSZQHPl1Pp/cmpVXcEfBeb2VQYrGHgbn/QBInzJqUliY61IOK
rC9gzlPRHOag5r71X4+s0hlySCT9f2OW33R2fqGs9wy+f/S19AcjBwI2UET7BYdH
CZRzcsiWyugnFH0lpjKW7ytQ1onSKDKm6o0yZ1l07gJgfjL0pRM2q+Pn5Q3AYN9B
tpNJ/SzYwdUOAb4yI6GgJh3yJF/6ypma3gcLKZevQEh8/akuwgoyRSDWTKPkBnzb
o/9LD2VplAg1QFj+PGQTMVRhONkRi5XhpyqdOUSyj9pF6sJIJwBiWIzDsV+TIfsi
OPzqGvka41tpUREpO30u5QstNNw3MP5IQ4YQVZ4U4wH1oXqyeg5Bu+auQ56mXPNk
dvYoLC6s6xRt0aJkZNSVk5oiQh0mW7U6nY/6+cL/qOM6Xk4tLPbBMKnNU7vF/GW5
jlJE/7HEWyG75WyrRKxvT9nlHj4bMEI/K30fA+reswHtpwYk9WLDMfRiLjpqc8Li
vgCw2lqg8dvZ2EIk9Qk4baJn7oSYlY1lt8w9mq+OisyReRWy7b9IT6fso/5Pq3lc
sogDZ/iF58lsU7c3pOJO5ZhBKVqUJ9ncP7jWWMFjqmSh5mHSclrL3kINKrJso63L
WfxaWnr0cleHATlj9AOsmuu+sgUcokHOejmLjt2SbV422n4f1QCN4EedTo6z96h5
qcT41Y/t6aqrGlkFabMxbh0D84eFQkcyLgHmW+K7JTIwE7aJIEWvOpoV+T11tWib
lrlHnl3ILpGtosrKgmE8xM35gdAJ2hB7KGW4R8aAdg4k9HboUJKhzDR5bUC44x1U
CYF8ImAqNB42qx5eJAR5Bw/PPaV3GCvj57GdUhY4PVhda2dqrxQiMpMrkHKfIXBy
9RvxfshDnvIcf981Z98twlPndi9JM4EOZImh7vI1WO7Exl8PfEjEzBvjk1b0jSKj
f3pLswAsBQygoE2oK/Yhc+kAfbBr0rUT4d5+9LH5z9eC1mgp+WdKihnkwYoHlXvc
BO4/GzxEWKAqXOHU1r7dOXAump0LJpWNh5JxsJ1bQqrTOsDiGOkFVLD+fnrsbuOH
bKHI8mwFL691oHh9S4DpQHE84c8ryaP3ugpGJyHbxdrGKdRrP58y1xwyKQ7JEqrh
hI1nY7+9vVl2F7NIHF7H/idzEv6VtqLGhhmYxCurvawbBIzjegLxGdcZXgkBQMKq
MQJfZ81nx0fyJ8SwsLdkOpD/5UKe1On59TdMok6NfFG4rpmzhmjLYo7GMMZpTClA
drtLKNizE36wRtH9/Mj0NbNnbM1atG5cdOqH4LWxWWCN+g0/Vmcot38xIqRgWHMb
/1EXOo1inrQImJczeY7wOjxr2EapsxENi1Nep1mQtUWamlUmgv7Rc0b1w1Qx7LPu
O671XetZyUY4rTTgqhnzNKd8qWWnzPBL7GF2UIegXrvongDdjrwQQCaLyilxHsQR
8FwDBW7GjdhmGxO3WZ0H87LBTnWCpF53a88ApiNV7lve2y3UKNp94JZx3MqIUhhj
pvO5YTxD7cvE3QRfIZEwp6Za+M17KaqXZ8v2jMi7qRfT27C24jM4/qmGM/fd6ge3
ogioHX5aHXxYZduW3npuYD1P31solnQvIrFtI30Bf0meciVblnQXUMysxFG2PMVQ
c3q9XE/pqmkYQlSjhOAYvS1QDMeT2Fa+MxRVSysIhqw7D94oLD5Xgja5AyAwZA58
NQclq2m0vBYl+HjeJn2tj3p1ahVQp5v5e4eFrD1HaSZsC0RwzF377a/oyU60GnSS
PR83NeY09wRIKMqfDTjdBFtSeIg8j7ysHp1uJTOfJQH/+IuYHQNtYohgXfmsR62N
MC53nIsPEKvsDG384CXMsrkXjboi0db4BDUYvWuimZxOFC6TARvI34ZGwhghFt6t
HsKuiP/ruG+r+XPLi9r85ak9hAOWtXYCUDW3HUNPYgY2QpAqXFe/jZit5LrLtPYX
NYCKfP2K+mXGv77Bc2Pi1plUQqu4ksFydaZQhgYyQ+MEm0I2AxlVzTieOnNEA164
c+724WQwfTQ7t2rjyCWC8bOyr+5P5X8X+mAY78+vlw6n8ZgkfW8wAKPzmAEGFuan
ql8T8gHXAUFGSxZ7PgMLRffMoy3LPjcv84O6KwwLTEDWa/zj4UUZhUTlzVeXFx0A
QO+g4jeeISekC/3008+MbNe1eAqGoL2CyZP1CZSGBDHXL0VEEktd2pQ4cIM65pWf
pumnXOrtgm4VBro++9cS5kJ3fAKiDBPjs6HTZ0xA+OQMzL9K/r4MQB1SBbidov0H
XHzFp7OHHUQTK0NOiboL5dCYYPZ50x/Fw4qYxSx4XT9lj064hmz4T8cjEFHS78gB
Ly/WJTJrAErsAoBNnn2CFU8sZNebfoISuRdCVXa5VTwWX7tozuWLxO9gMK5NS6lG
e/AXyZnC0GEwYTiQWR8fDpII+PQbzljlEAwbJp5ppTfE2HsT3diuRKVEsyfh9lij
hEosxVvIH0+bfsGskc82NcucRO7EPBvuGd8vForssmaB8T0XHHeeo5vwDbcuy2RA
dP0mCiwJuCELpJwlp1il+Hzl0QsrjsIx9aJRS38e/Zow5+lnKG3Ox7WTzPiRPtJS
pl/e2Q6iJxGpXgLtFLUns48448CoDl1HjYaC9v33xMpDL+rsHjKjO+d+ptTaLYUo
oqEFipwTaNGTl+6ghYMsyACMWdN/Sauu0cHhAEj30IdWXTaGN9nuqjJC8SBj9O5J
RDJnmOkxWQ9Ru4058GH82+cSiCjnSFYAP6as6RCmD7NnMvVjJvyWZ0PFoG4ci3Ez
HgkcMzE0mGg3ahTV1dd777baMH0q5FfENQ3tCi9TMr8ncfDIM30fSxC7CdzRBjAR
gcixNjmfCV0K2Umn9vdIE+Yk55/lVUfSiSkibJAVQJ2wP8pDku7gHrDDCTX3lruK
3ava3KSZFre+qVm+Sh3FG5B9ZTjQeRWtsEB/pKcOtCOkE3UHLfP6lk826Z00+MyL
Dx4COlFUwOADZLzvjdSYfwDM7X1B0/MQ9oOkeKkm//gJC1//cvlZQ/3dk8vRPdSF
YVbKrfWpJJeACRf/uiBouAIRLCLAJ0IqVofyE+RuxiV8WO6wuQZSbjFmdLrMhSNm
DoUOK+tDfDBw60AXqRIRKPoLIknr6BTOoLWZyR3m+94GXDaQCqfsHLr9GH0vfIip
fSI8vsYvmDLnbnhwbjjhzuRONx+oRw+/xMOt3on7D1smnJK1hj9Koo+djWUewiiH
ShIc15muOoPmoj/WAXVkyQzgRDVUfspawxWb/5l3JJNmRYXG3Va9fWsQ0ye3Hk5N
RK9LDzbePhi3BSIl+jQ66FA7wmHWYPeOhGGO/YrPxYD8kQ7MMfO5M1eAiy/9YPGS
mgIeru6mljLnlROskSSXwhHLLXtLLDmV0l+Y1ifbGFCWw72TymxYyW7WwSTJAt4P
1vOO+fzOwQVr9IDowS/Ag+Ds2QRBFc8HgvwFoHaiUH5i5VyHWD+e9CJQQOTv4ApE
u3qAnWScagj/zPfi7txhpJ7KvgMQHG2mxMG2R8g+/hSb47MohU/FrPPM1sTs6pkg
zpCtBWS50zN5DRzTnarGM63+p4qwBFpSiRTe2eNUmtebB7MOfhPgnsaxNBRSwTHy
voWTCCJiVpTq7w6DL2NMZlIuZAY4kHigB77jwoUZZpPM9uQsGmHSF5WP5MY7r2m5
IH65jqE+i2+SZu2wma+1O6nuoyp1iArYoc8X1KZaf9MVX4odrM4DpAX/uonHwiHM
7Z7KnWCCN9IXgAkFvRaJTbpmLm4ZRTnFeIL2ynrUae7dnGvfhwoS8cKxUWUum6/a
pR6F8OvvWpfi88JBYwO05Z0a0poGImJ+PEdYdMmhu5NEEMi5NpYgi9QzCBVFhd5d
ac1lO4eWisA0/5kwKvScM2965XxGjArAcexPycpXhj4RWtka+BGTW8ZG1BoKZOSx
Bx27exTFhYsT0BFZQQG2L9qb7Gf+Wr8DrrVlPeCSD//kIisI+JSMAe1nFLIG2ssT
4J/rBu8+yMdGlsKxSYsp7u+m8Qk87XSzzK78JHpES1kjobUsAHKz8/Css2x2BZco
Mm9+dgf2DsIa+y60U1KqMNzs86mMx6f7JrsPFeoqSGA9o85R7WDWOeh1nj2i0Viy
+yFjoIU5C8QzV/YT38mt8wYlZJ9LUMy6JvhKnbCayHaEHVGrAqvb9fHQi61BAo4B
ys/yZPeo2z3JbaBz9dCUKGg3EB1Fq8gpapoKd2IADtvSfXcJnzgpPk9Jv2unqSMh
8cmO1eHwrCHG/a0ZcjYR2QwWpmGyhWtcaac7558aV3BHb9rAHUpMrIV6s0YnyXme
F5yK+w8eCVwLn+GqdI3nfAi0Y6B64qvEvOq7p4cL2+UXCLoo60wL619vvE1wL9eV
pvlmOL6gei6UDHDNBVZLxv+2DqDJe5aEEhZWSYs8FLfhHcUsnUWVtPKxUbRGqS7q
FzTrizhAAa017vaTH0IViRx1dFAsS74GW2npB3mTGrsvIqJJoxOmgbDwjkxaYZHr
IyylEJR4it20l+wMjaIFvWmp/Kysuv/+7fulwoCIlVZ3rJB6d3HanGb1zpXMN8p+
skf4h8NfYMSIWhzkVb5M63f2NIAUOkslwcQtH2X4xyRvfcfugECmuAk2tpT3E8p2
1mG5fDp5bWostdtgL+Lcrbb6wttnBVRgh6ByMXTy4+YBs7p35eqemLQNsdum6roL
SEI8UMyq2i0uTL93EyclVEdxKsiPVjPz67jSUobp0snIeimYMY9iFq5WK2jPav17
oYnMT6K43ZOGj28CeIH2YVafPb5xNVRVkGi5cmKFT0lb1qx4EfJ6ZruMsGLC0DT9
3Yxb7auxrzLL0292dYrf6FrGflkN+hYowUzIAXFSoPI+d1qG+UW7/h6XXJbQ7VP5
4ZtNJa+jBUv/cdpu0GdUe6fNvBSwOj6FIfkDeHLuzNG0wro+KCwVDFGiIf9hTtaK
ILtwXWUR+tQ0iCw4LQH6EwRK779QLZZAbe6UbsxgRetBx4Snht1fnpR94DzPm+7y
LFhIE6ygDJTmj4F6zYdt6K3PNRLodQ99LRm+3Wx9jFCFF01BEwqErNL7kb1/QBRr
ncMRc9hHkqEnk1U0AoA/DP6R+m1akP+JkL4cQGrqWwLP2jcHNtrl0M7xKflUUT5f
IOXLsvOeOi0sv8Q7k852v4I5luwGxTcAeHM8wvE/JhxQj/ezIORg8dCY/GU0ZXEl
4r9KhLKyCxJObmps+7wWdHn18tt04zXJMNwnIhFHHnd3P1F0Dw7qJuu/aJ4kvJjs
/WxtRXmoWBDaUdhStD27Bq2yG6l/vZjMOf/RgX9LUYP7Q9Q3LCamIJc7GQ/cDotn
p5OlR6Q/X9kBBCvRRHDrWE7Re4ZxC35IOE3J57ufMI5jCVDf/ivnRgGe3IAycKQB
cTIJ4H0KXFH3hXFkOogUt6IIBj6Ha1u29EC2SwrV1hFD9+UEOxL6kIsyA3BZqp36
c2Kp62ynCZZ9XbcGFweGog+IwBnzCRvaOi741HskRD6HzwJnhyCdzpVwXVzXrPio
VJHYvtgSpxMkt7J7zrJBSKPhB8+/z/Q7n11DjfXsH6RWakCQS2nwR8U4CbiK46EH
M6y1xth8Y7qT5CQyUa2SRbrI9lb99V/rPdAUDWAB7IiF//BzzhSnOTa/2J/LExgp
bVeMs798Fb2nTibXoPOAAPpPnyFh2jBoA1Jz/hDd0ItIiWpvll+mv44YIBJoskC3
+/uM2kzBdGX9J5jhCTP2WqRKSVKz0PQkCv2jUVugUsqge0YYq1guLbyvLyeZP5Hz
NlmMbYdrOHABFzLfT+eH/ypoXx1rgDHFnH5BctsIiceA6dXicQIdVH05WPF2ZTFa
ZUWZ1hrpUnQlDOMbcALfZ0m3O/lahdYYQiZohHr1Lyen+vpPlhlCiaW+w/zr5PSY
KbQI14xJV0noJTuDqUjeVVrU8ue8eqNQcrn00GRuwcdImlMV6cYiteQAb6y+xGjG
Wox27mJ48jskGm0SJFDRw9ebuItgD11F8EwqLhxs1VSmSd6qMQynamNd65sYJaKf
hWBFMd65DJRZ7gYht5eBSZfbJ2xl5oEXJze4065JFCvoBgqFvrmPlVga5MLNA/C0
zvj80OS6sWaaCeuArhrVakGGeTEuzZLpXegr22NC5l7xTxVfbKTZiRioSNXGjyPX
Of6p0ENwS0XVV/X0AWO2WZqdBQBuoNYh2vARZ2ZYUYMpLNpudKreFwFebBtOSaXr
b5yDV4DTl+l5VhrGKHmSOwYrUG1r9cFYG3IAOMHHqawQFsWthTzIdVC9i05rOnwU
XZQ6SJimXnO3fPgRyYYIWIWDUfK1fYeBDwcguBO3kOkgvr2BY3YfzQ6Hi3sYOYhr
oSGT3zVnfqprcCw5Ps7oAkDdBT6OvckerjJ1BJDlgYuqRWEaSVb1qGwP0/ACMrPN
044Uyga/3vA88lhPoz5V3PT+Zg6F8Xssyio2acgqv0Q39YEFOgdxnSTNnNkZJ/eU
jnaly0v30JEO+Pzbu+cGaH3XDVpKoJHmvtPTSyGjYhuh/62fa2NERCVpLoslnMlt
MGUrHINOR2E2cHEgh5HpYiKTr+R8UCFQWWUlEuZf9WsJXqHflafrRtnbcFGYilcW
TigBabYVP8aIjMxteGPRB7CZA7y60PGOiNZDez1FVyT9uY6feOBxf314fbhFZrxh
g4oqLhmBpNGUwt3faFpRDGT0ANeDgiar3objFjggi3yog4OIawKdV5aHMZ/aj8e7
Py2AWVlzwGv6MtCscYCfWB5Cq+igRGQTNPdXAPVh9/5JmL30IfeL0BR9DkIXT9+t
PUkSbPmKFy5S8Af0m4XQnRuktk+b/Kf5g/xZKwr0TbqIZyxfI7uu+NpIEX7GaP8J
4B0HgQ95dWJDR1KXo5iG0ZzlC5lPDQBaOOYYgiBNeDdix/OMM+BlBb7VIGTdkm6f
g2v/DFN4myR8AG8BD/uUTHGakWVbRBBTj4bjw0aF8xQzs0uWekQm6gR9Y8P0wmL6
ZE42B4n+yBonfF/aBXSnenwb0I5lnOG6YS0PJ4n+u4eCUJhUfbbSFaVxyRF+1gMe
zy4MXx/ifc5PoF+PW1R/PVPB01p9iV92KZH6uD+ssxN80QYGwxzM9uq7GnUvBtx5
/1zmUHXXdN2fujRLIadD7rsXEQeWsh8axag3sVzulTaePckFux/BcFnMhYiiJKrS
K43mdhEeEMZ596Y4K9LDpjeQSnNNQGGjHlRLA85cHeoIhDSaFZ6X87le/3Ib1cuE
pXNxxrqvXaxvbrc4x5BD8oT57viFtg9qVmeD9BBWw6k6uK6y29qrOy7FrkasY03O
JKrvUMRzZzoCe6k8zqRAW58nmuLEXTJqUUU+k6/3bVDMxxhWG2fZnLDrrt5kNcZt
HC0J6NCudwnfVs+lV5xG3Uc/NkRdKZMARHVym1E4fqiWULBb3+xmXcImJwlq9Pb9
Ar8MoK2maZK3K/I21VSzAxeysrE1G7z/E14p6jvd4ZGJH7rwydaTXe2qvE0OnMbL
PhIXRC/WpWZ9yb+k5bUTOm4DaFDBNk5az842KHqTS0GEkqJzJEGkVgzd4ccHjzPy
8qwbjj0gBqkOqbn9WSEU1Yb2qfw0vGnMg2rajYW4Oy/NQJA2xwQ1lBAmN9fO67y4
H9wwqKzBhCaFUgQCJ77mQw0NR3DtIzLYe/ZIUewEU/r/eGUj3Eq8dBtnU1fbJwK1
qjqw1Qf7v6d9BOSR54oMpBDiTmaqhi2gSLfYUtamGrNTstVpvpKRf5g/KusnndKz
KOuvU0ycgiHfMH6dr1N8y6Sz1cMx0oYJBlN7M0f6VxR8FN1t5UAsl3oo6wULLYA5
SOvOjpWstqGw//zkkI4ZLyhbB6O3NhuWagol/hTJCQvNnKhRyg99+GbsEbMmAqda
rIHtut3eYffLFJihK0LJTdRD1qdQjHO0OVQUlarNyzBYDOMnQpjAWSDUb6Jk96ij
KWKo0TTea49O81ZrEic9k7X0b9pXH8WB5uMttKYT4KTxmqPWWumKK2IgJ69oR03p
1YVOVchEZHOi1g32rZMZj7WagtQIJ2nDFBh21/3I+kevjr1CsORetRXc2M1Zwd7U
02cmn2NOGnCSvcQ5KgslA8FAFrjg0XANIMQ9atfHuzSDG7Iwwr5PYBS4G0nUgTdX
E+6hBiSzwvpVyPYY5/0xiyj7TTMnmzXpetuanWWCLK8tITxslESsoezRZKxqCsiq
UjVa9M2lx3uMMM4WxeRGcQVHtnPXsPoqEY8NgPE2yLmjkrildKRfYIolKbp1NhoB
I4QcWkwnWgdgnkboFYO2lv6VymHQNB3vmTozz9Mfltq+QBkrZOuVPCTPvpGsGwnw
vJubTirn8WrROdAx0sj103QiAthGTj2fRajvxTR3tHcMPqveS1ehwi1+91kHfG9p
FOWXYHi/UWEjYuOuqNXWYS8Cazg3gFz6nZKcCIT1WBZ7OYOXvwajVZk71XgDF18V
Ils1323ip0HzzajCzjAv53HUqqkbzifAGV8dxj7IknM+9kT0EtUaR/S7pdwh1kRf
RRCjmnlZm329hXMFj4n/Jjzkygd4EPbk8CTVi4ssWXuHEV6MeW9kIw9ClEkpUOZH
S88CS8F9xffe9LDXgwpITRGYgqWfIIKuPNezuaF15ewQ6qB3eZ8fqhUSKH1tCRu2
Ywe/0NXXyriBbeLE0LWUgLhFJZ8SmiAeCG0gHEqEjWldvoVeho4TbqOFn0PobZ6q
jyLE/lHIAF/ZN7kkQhFJ78kQR/2cEPgUXKJmqsHxFtV21qa5IPDUWURd0gSCu/5V
D/Psxbqb7cTSlKsVzA1CYpBLRd4hVbvmy4klpptRsenVxY8aKcq3nmmYh0wo4syf
aCw/joeAYtDf3QmlkWbQiwBh/5OyOEcpIaPGMtK+ldJkZ5Np4hzsW7Zt/mBj+aDM
ENks6rquXu/Te3gLxiuK4caG0EP0Di6wlmQaO8nRgSR5ijZeZW0dviilGrszKs0W
zSF15skTlv+hnKNwc6nR5cPs0UbXgttr0klUH6KNqQiaIX4yQr4IQfQ9zxOTOidE
jOZHoBXf9xjM6HlpxMlL+XrttJcNDrvbAUjAxQMl4ID21YhbVyAYPpyBCCbY9Vju
OcqWMwoIklWeUAKj0XZsKgjgkoE/UH62Wo1U4PiDtBXAJJ+xmSMLn+P7fQVtuvca
s4pvQ3STIHomFYh/2vggw28kgYDMJzRHYqlpiE2SLqNPCeHKnWS40ctjZd/2Q6Gb
Gz1OG6e0fri4UCxmyzultUlEP00HqLDuEilZzaUzvdBPV0TJOensSfM+IeOU3vsD
mzJIoCIgpc8vmi1eGm2U5G8NYvJyvWADr5SBZEYqN6zK+d6ilAS5hSYiJuTDYRwK
PHI3ntbr3WSdVS1KHwNnt1CeEQMDjvedDRZZe0MEQN/PvaN9G5w3C2ByLllijU5O
22mCEAb+F2XidjXKtE0uK/vDPGIK/qy8PvvqG2GZh9VuFk1qrgVJHds0vIDVQTBi
ZFtQhzpnwQd5Wq0bEiMGfvoRauGyMKDjUsVg8lhB7cnh+NHfLtr+iU0L1Vs9rgSD
JmY5NSkiR8Or8Ha4EVuYeiGAVlmjuNEoYarw2cdaMiqsVRyQ+8qg17zNnjL0eW+B
x4a7n/q0RWEZYsR9FkCFmcmeizMNkG5DEiiWq8O1Sh7sHmGjNM6gtdr1kPl78c5t
pTzY933gx0peUjsik+a8ofWPtQwtvLEgfTd1n7E1DGqnTZr3m5frI0lm97kN+Nf7
/gt7RaUhLeotCe7JDsSBIIPK6XE67Rqxh1ZXu3yP2ZBNn9E2dZHhLfVv+EcJMeWp
P9Qa7CFQwS1wszTWVfpzhYaS7pKJpJor8DjTbwPH52+GWkPET2ag3u6KjgK3XSaL
U9mjnefhJeLh2xJwBVWhqgqAhMtoCgP8Wlj1V38/iZrOnsNWPhc/66972CqFoSgI
M5yxqJ8ugq/c1hcvza+U1/XaZPG8pye3JyjUoFHhV6shpphn4INzidTYTo/Vc5Tn
433q9f5f22lQ59bYB8Og7vr+wEVJQUK8xehcviVuAoV6u8CY94MGkamBgJzXyumB
cnfwio0RnQPU+LDgsumryWdILRNpdZDbkRkbKyse+6DQoVODhbK2/IK+ylO/GSKC
XtRTGgwqqiDTEpBkeIpDF8wwEnsat2KNAyZAVBF6gI7wrrYeqTM/Le70GET5Fghc
NDWkoTMZgm9gDjbjJbjC2k/xEtAt5yI54967eZ8Q1PkYyhP//tUMP77a9tFNB+Pe
uzMKz7cwL3Bqz1IxjC3zN2IrQZ27eGhA4T8I5i4zFr21AnrinDty6q143ksf7WWp
hABPvq80N5s0RpcYzv0zrEQMFbs6+PAbzBpp+qAdsYjRr/228n8x50oXn/SgvrIO
oI/Ur25BSzgArKkWgyS0p2BQmYehXeinwwzq/5yYHcdy4O78h6+oiUGXegsSmLtz
6f9dwC/GcOs7khshngDimQAPeVe7qkPy42+7f24vc6zPcsD7onEvIWRgCfeXkFii
caCRVlc3930yR3DZHgEcyoqCTz6hPmHQvC3QLUB+CArlh0L3VGwrmwpoQ9rQitTA
EUMY8sFOuxnbdipe72rpsc5d5zFqD+jMY/bAInFSLizVTb78ZI6y8H1h8WfjKp/j
YLdo4aDkmc+g9OgEndhPHDYbFnmGLFLbb0YRzl6ovc+WYejBrnJIqKwnPnyZ0o6I
iJRj682zBR/KA0cGy6/fUwdITPl+/r/NgvIuRiHbqWWr3/RGdtcDoksthpdcjY0E
EmWU0gVR/f/mcOHmUpFBAG/ey3OJNwLuC2jQ18/VJSPCdHyNRpK1qugZd0QBvIj5
rOwPo6RQMB3oXu9/gmOAHrKTqIRonjUb0wIusAuLKzjbl0FZBgFQX1z0ystFjhiQ
JbO8jBKfoHVg6048gI9zfkLJUMtEBLz7HK6zRP3DxNQ8Gn2gdXYCBlhuoCx+Cr1R
gn9JbusWvn2y92hfXKr4b6tgfzH/OqGRVFoqLwg7BZPfxZiFdVVG0kVnrqmV0QiE
Vrfmr7fjvIn1dC3os3B+ymhTfPBpx84tHOBbcx+N9dbaUzSDJGyaigoZ8oTctehg
UYP69CgNgCsxoQNd0yDWqpb8wvgY7vRIgOEZ4K+UETIMoVSgutWqHmIfy87yRSA/
Ln7MzykiCKkMjxMmX+60+LHODcmyVHqPMv4uicLnANe9b5UEsxqeMdaKfxo3MaC9
Iv+9Twf66WZ69r9Qjhlghuy0jax1wfOcOadrl1XJbX/FiLeOzMuiYZw73dFJffUN
XdNRWkYFee3v6A5mD82PfR5yUH9OTbScZgaKrkznB+M4bKVqSYcbx1SXu9rUbeSm
sTIBn1/ZKlOBYrYcugh6s698PKiGXwQXDICA6/aR74yozMfcps3/mbH5uI4SZmlK
xOcCiKITBQh+d8xa/GWt2R4RZcIiLgF7KABY5z6MKVnZh+wEZ4x+5jH+G0RsgEY5
BfnuFwsNExpMqw+LY/ufQY2DW1bvyBai0URJ8p9CxJhHKTv2zatYh2Ea/GaOBQBq
zb8ZunnH9+sZXZvS5TRXjOfCXdoBDuHM88tEC8R/KOrTZHda98AWc1OpNBUsoaNd
XhJRWLPMOeaJvripANB5dfkj9f7kSKTCne22ScQu7lxcBDZ93i2gzxIiQVBlY32r
LuX3eOA8SQ5vxJkRVcgtfGdgBh74wxeVhWQRk/Xy9ZYg93Gh/QImM9IKHb6gTT/R
0I0je59gK+AtqOtFDhlaj2w2tEMwliO+ebaGTbYqB6sjzvMjcJlXYj3+Vb7sYiye
o1H9bISDbHJhO3BMUODZc7Z4M9A0SAv/muLb4GYX2O4aqKKtYIHA3bg72wYA+WUR
GTEGjIOpE8W+NdFEL1NIa6dGmCcMrS3WlG1p2JGUWWlLfhbYNZ1/m0AwCRnLzRL5
BlPYcYDDScxCQT2zYG7Wje722mawF0YnZHR5pkGNf7fc7f/4EdmQknK1Y2nAb/sk
t1MuYm3iQGGbuOTs3zOVQW8g4oVm9EQfA4v2/Whwi5b9Ic0L3VLC2WIjITSJ/dpu
/AUyqR202xcdsmfuXEfCtLz8qGhr2HHy/eTSWRaiYdcOvL5PsDfccNwUha5tHW4a
1qgJj0bWZT9s1n3Qxcvea7panghN1L7bWXrMqrvUGuUW0fKLu+gvJMwTfXOVVrfD
fo+fndiDrYsVOb+H0FDBeHiuSrRL8ewFGueV6CRCANYwEo4pfuRvSMKje/0hg91S
JWt68WRuhXZDZOP7ApQFBLgCwRnytkz9hshug+ogfZT80X7Ze+mishIUYjXuej1J
ejYcx08oP0uJdX1jsi4mIeBDSA2d4eLfn26W9uPAyhrjsodQwkIPpBETRuF//GpF
cipR3jZjG50jfZQgGQt6NW+xXBwBJxIc5ogQGt1ZqiN4uBoyftI/Sr/iIgJIN3Cy
BSZ9YDMBbf+veAC58zXQ4dQlDdS79F0C8+rwqLR4RA5g7WovS1/XzR3S335KkrwW
BME/SD4Rw0wqUa093WOaf0h52BpUoLijDiOuZxoI3oJHTBxng5UaKoh/RvFDXfIN
z9bcbstvLYcgUQaNvuLkw9OZVhhMcq9tKQwsPp+20F1QSE45mnowoO2/YerazHnm
AnTfBXu57B74DSvG5CDNzoINy5vjGI1zCoYn8Gy1KLG7gFWklLgRCRv3ORUTjWiV
D35rocoCjMmQxcTn6PpNTmYopGFB6Ei//Pg9B/lxMXWED8iuKiPOBRdw15lQw13L
MTDjmZGtcOf/fu/DUt1AA5L3kBtJLZWektXCF5Ey3fpAislMhWhctFBJxkKye5RZ
E5qZbWmtL6/mMVbjivAQpQXi/pcvVG0mG22PZB/PLXXGuO7hUNQY7aKYRJ91YnLs
q2cAMtGgqrWU8X8ScPVoxTZ3XzHnv/YRky6WKH7Ow/a4yGfumnrhC/AMf/GcbB54
/pRDOk907C15252my625SoC2DMcfvws3Wnxyx14yJ+RXEMdjDGoNKDOpcXIpi3EW
pQddu6G0qG8iou+NGJiDxzOw6eQH6ysvJdQWAER6TvGF7Ao8QuibMXsp6RMcEV3U
OR6oUuiEzrnMnoyxGaN88Ma+tIQcwGlG0vSogR3mHGiF1bSlG4d49AIB1DNY6Hmo
MKA8mUpZvvHSTUSfeKq//qlfTO61SESmxQh9cUFb2T1kIU3JqcP3uEDz/zosXvPX
ZJtkL1otiL8IqIzXcLrUGfabClwBQAIHKYpPfIUpYp9Pu5xmpxdtnTVh0lGJIZ/k
LQZYm3lUxpUgorSTxUsH8nzNWofecs4ChXkaAWJAc4M7BxmJXbm6HazKm6/t32so
N66jd96bQBXH4FSqR5xs7ZDOb4GvCOgGQrpQwY+9c8Sao5ONqBXaj/eTU8eLECJv
kr0ztm4DmMtn9c+v6XK3i2NxAQcKwPjaf5AWZESFwBQrMa76VKPOjuhtT1P5ALVv
61yujfwj0bPA+iJY0jMlOdyaWXmwk4rIlieHNFCq0lIWbbDYewRO9XcCWDgcUHMm
Evv9aLQq19cU0gMo3gaL9ZKXAAJXSnUCi57RmYSZqfXdcecCPJVOnbJ/zXk4EyKq
DmtMoOQ2JVOwBVmlYeETU9yc+HYqRhotePFp2d3Ec13lmRf11rl+WprgnfoIPrdd
M2Km2jGgM7CHL1TFlsAvOBNIZ7sTztVo+FeDCGhsaO9W2cJ/Ms6WqOoD1oY0yGpq
233AhcRJsC26kUssI+VDJDolhXBuD1+c7qHFWoajPqvwzBTN2tfCYGMVLofRvQsO
RUeHt+VdCKbLt0QDk2GNVuL3UDXOuqVLZg3Kwu0vIrGG1pIhakXjAw1N6XZW+KIT
JIHt3U71uPDvWHsahxaBXt59ZZQMErgQiTGV8eCXNCfJRZMPJlPsi4ymUhY3seXw
IVf2JZnsTzdRgqU+UGs/OLi36DJYhknHQQQEgToRFZBDHlRMJ6ZkclqZTa3tZC9l
F9ZUgZTpNaU5+HH/xPLc2tcLUVXW56yhS8ZOoCQxqD9ISS33ZtpLRh4UJz6BjJJP
lscsXsaX8rn5IEIL2MJsDaAJ4rQnKLXaZXPKZ1EYl8Nm05LdxdnCPLuSmX8BUi9N
p6Gg9wOSAmZWTGS5aD4ysqw9jmZWD5zDRt5X6DPWT6bSRl0Q3/E3k7dU0XRPTZvu
BCZXhv9eQdQ7mlY6j7MVJ6CecuWEUEAJ6V+muMQE5PGwHUxDBLQrJhXbvyEfk3JT
sgBBLxqTWaNDrSLHBqgqngbTGxtvht8Jd9Yrz/vlEL1TmDItdePv69AIgldTEk0a
RdIJ+mBCimUV+2rls6i/UP7LiXqByZj3Bec4+75mg/tCCKlnEuYEnfSdaJmw04Pl
WZ2WZruIZD5wDAj8aho1FHqPXrdDkaNHH6nqW6hq4nOS9yQxpEzirSI5x6nkQXz8
SENUVc1Vadk8GLsJiUj1r6ov+PuK2hDUAqua+VXb9BpCHYV5HRBMHO+4SXJqjFpq
MCSLozF46EaEvSzAtTKeEgnPecQxEM7ViUMi60fHQ/rOOhTXdkdiIZI4LjMtzwF5
23AiS78f3UoZvmC39Vmqm9wlUvd6dWuTBAkSD9Gyqn9BLKis8HE14qpw3w1Ep2Tb
bA5nPlJmqXEyNPFHfKfSSebAS9L7Pld87/8hU6kMzt/UoC986wwGI0IXmiq3KHwF
92R5D5/PmWdkCylXQDSb2Dlwf5zPxDi/LtIO7B2Q6Fm/oUCmc11LrCDbx1guF/Oq
N7K7NpuO2qHXSv88HYlkmp6xsgzycccMrTvPn4ItRU8r8PzUgkgd5kwpKLPzD4fM
fJmog6WHSkgzNzAygOwxjSVYKgRfs9M0k3vTwpGE3CDq8v5ASIaD//gq8FGfRN80
SzTKju9Lgwr7TIHP5jNDNhfLk66U7qLrow/8jvLtb+5k9hBnXYlq60QhEwhUNBE4
VVxDEsfIcf/4mP9sl1gKgypCbyZ8e8CuuDcKzbBihxtYMXa6BToAy4FgimQATuc/
11S2KXY4+FGCXif2Xr8Xdx5eJZ+3+7l569Wpr8XhmKSeeFqKochSHs6/Y/yH9/y5
NioPLADRQq6r7HOEtuLbhDqd3v+b+voIUvYy33eAkSR7VcN/aLORbmjsNBE9qPeC
elJW93cJ9xMmZKz4zy4TWN5gUriV8KHbCHByZNk73Ql+hRL12xw7jYSfgTqCW+3N
L9dfgqG/O5mrLZwiqkaNw7S7Pgr0puBIuTojZVot5un66/mQZN/PBTR7gKArYj/2
46KjeBD6hAItf2Daf59+JeqOMSCl7zXZ+PrC9nrXeigYAXrRnpKS/bXYXco8dfMe
q1P/5bKhjIHoKa4nRBnpSNQ1F4+Svjkyd/KW+ZJBE/D/5VsNg/zPMmfDFa6H6rlD
QHDxN62TTrNQD+Gi4NvptOVclEt1ynscpvMdOOSa/OWEiDDQinn/EIOzGlq54xa2
a8YDCSEDae3xVy00pCG3vpL07WoKX/oiro7CY4HspZNqr0WIAjYmL5yHJMZhPhEd
oaqH0eyl54epgKoa74518qKWZAt4htJSqP6aiGj1WAERgyrBCDKaCJXHn/zCAwzF
UNT1zQZchjW9uhJ7XD6/Bv5SyzxuEttPk1fA1GS239SyviRYSvSzZG+GK+k+gRZz
xnp3vvWssZmDvsZRtQXLxhRYCWljVYIqzMdl0brk9BFF2ZZTkm5GHbA1mDWUb3Cc
47M35jKcsKF4aB3aZjPhsUpwMKiVjGtIpR2FhLxAFYmeP3oCzrvtOGktfBwgcYGV
KTVJ47C0S8vY7UD78FWbIKrzhreGcQa4czzdqBvt+MIquG3m0EaBmPdkqM06uMR7
aAS5jCWFUSGcSmiWqUTNsQSHzyf6SCyusY1ZLIPEw6koZBjGocVgVFDLQDxIhg6V
Foe+gBNsqeZd9+l6+8leXeO07ZJZf8D3ucFdk3PWx8Px3zVdNGxtHfeKbv/54Wcb
gDqq4TpgKF7Ve4OkFbbxdx1Fmm72rEPVo+drWbqfoNXzMqflv/SNlzEK17TOlAqE
kgQdbX2tjOGghToUVgIKzPJU7OyoVW3e+U5vuFinsAJhZIdiBSCduvcN0AXSRnk2
rl6dczRJpEpd4cm9RcKA81Cymcu4FHzZjaoMjptgc8DncsZyjKhrwljpLEX970z1
T1nP3LApy9Q8Vo6TBlE7VXuP82eH2gSWoxKaNPwmHPvXim7HqRysIWyrZJ/AwRl0
fKOco6DG+BWTIEuWKMulBWL9SuDczOP/a2ooLIaAC0kytJwLfRIsTUUJVogO7ePU
dXVS5AGhmldAKVPdBw3T+ESPymekT4ZINBu1HnJ/MeCf3L2nPyc3dTAYW2oKlfAr
roJCaNNi3oX/MhBXMJJr5Bdt7F8Kc2KkItw5kmESWojHeIPscUol4e/rwI8T7LBO
6Iu9/Z1cMNqhv5OxrDDEv4C9qxImhPpWIYbJG6BdN86u8JYVM2LGUQaVOhlsWw1R
cvfUw39KQ3Kyu7SfHFE1mY0YddllWUuaZaJU+eOEx5bbfquWUV1ta64tGmjXg1pi
NG4S/ZfsNwo2GXnakpJZ6gqhEbxqxXyuwq3R+LEcV3ExbV9i0MLlz1vZlkBKt/Z1
YNGXIO7BJv57qaphOgyLHWjLg+IY5JJ4XsTohmVk42lBw6bMrXE4fwYYPIbmymfy
ctVlwzv991gK/lJAAKsKPF2G2P6DKuxw7p2xL5ehJlDqAbnBgpgPbBFEObblGQvR
4Fa35MyidhsXW35HEnIvTblTieQprDObth2027Tc6kvcQHmxVipc2k3AMN8Aj6bt
wEORIXxvCkfC4fkQLMvWKVZZcOqc6yL1o6NiWLINhviUIcA521gJEADMdsiREWnJ
tq+BdiXqjm42RK4ufWnS84ZJYorqPaUNUrF22mtDjFHcEvSaPVN8owK30h/kJiMa
WWUvGbncwKyP6eJmmyItQaLfUuPaycKVmaaaqD6vBJEqxlNqTezSKf+rcIBHVcRB
3otsmKIjEhQu62Np7zQs32towP1NOgv/KEV7ReH2jshAhF0ENBM9ZMXGOiDSW0Rs
/6EVelXHSXxZ83/t8BBOmoMjkpmHeb1wrW3HJyuK4us06youzcHxqwp3IN8Xp80u
IqIL6yyrPZk4Aq4KhLZTHkQoyv/iCIAfwKR3zB9tE6AR0sVXcANsRo8WFAUzCNLw
w8pPRdSJAydGBf/LIAi6veK9Hi/O9C6ZWl0hp++nGRt/DOd9lgu1EbWYKbnxsmOZ
Vyb3n3rCY+5UJyy4j4Lmx12oHpgUb4Ga9IcOmR7yweHUcJmuebIbkrRKa9lj7l/f
jPk91el4da5Mr8SWtm3SzvaEQ6yzmNlxfy0z0mK+aCryZRivGR1Y6k9+KkXOhuT2
soSH5ouqMiO3Prws00M6gExTBcGlwk1D8k1teLJq23iJ3/SoQLSw4eYyp/7vffph
bskW+CIPcWnHVhhQWl2vgnPc5KEqbs/xzYKKrN3fpF+ET4OJhcV0uo932BqAWAnn
LaWBiuEodkXTHmXmy+bxJeVBw3YsfnpAR0Bg/ptjvHbVBWUb1SLWsn3igeFcPIBV
TvwA1TTbzJzGlEE7s/ntm9lMN/EvcNs/ksoHM5XINAFgbcbYwKMkTTEl/H4rW38z
QEBvIWdTdJtKSAAghWGCMgEwUx+w6+2m4ANBM1lgOmKdBhPHghacUKjbXmQpJluO
jx+uZNLIzo3lI2S9mOWieUIvjoMMhH7N8hxufK5Kyme66tgdfTYX7WFJP58Ex7/b
qIr3r26hQJXgDeqsEPb6BMCaZY/GIDTLrOOy179U2IFHU3SfWSUqqL/oF2CFw4oG
tWIll80ppHZhUd56Sk4r0AcAawdTae0hvF5KobMlgmmK1ldqz8TVsEsrT5k2zszz
E3Wu+37CveXQhykpwHy8QbYuKO8Dmcep0Qa1mG6sZK9Q4wyjs2jVOBAopIusTVeQ
z0xrMU00bDG2IAU7O1SYhsBoHgJwKzCDvnDPeq5Pn4a0Jy7kSwevEa7cTDDwegdK
JCY/2yDXwek4uBnS5JcOtw4GAN4D2GoRXdlvndwosRiwSksUBPrCYlN7EsucLb2Z
Yruvs2hRpNOUwa5KH7ROMqdushHECusi9eUaacLkGISJzcyzVGfB5mlpxtd2Q+38
COVmg2EFW851W5Nmw+xcyHNwjvSEqFbfxzZVxiC0UGkKt2T3bDGYj5yBMwKUCrx2
lGO323fLzlIDg/CPL/4LxO5uzDNB4cXQD/idYd5bTwAxdsOS4lw7B3FUyQQgvTlQ
tD3DTyGRPjVjf1V5c2iK+ti+ubisLbcAxu+U1Oehw33YfLznUxopLkIiaTEzgN66
jGCyDNuTAvfWuTiEQCCMtgNPCF0Qz7pZv2mw2ykf63VvGYyZmhOTR8gZ9EGBFq8h
0Ugg2XuSogj/4egwqgE0hJkTGxxUj9BYK+TDp3IEfe//OfYzde9V0dp3qa3oX2LE
oamYkdH59zbuHN36NJY1GUDAb5aTk6jwe3favsX4s7nrIhB6DtzmerBmDlqI5N3G
NsIylrHDYdI0/mAuc1zRBFxigQVAHC5I/L9r5UhUTKU0WXrbzzmOAEz2tKv7kS3W
BzveimBHpMTvelY1rKLDwBujtYjJyKN9D5H7MZVuiBTAuBLW9+mGqcTfF0pzRfc1
jmzbNWfCI5DRZgZ/Y0tnzupT1ak7KwkSpDHYKt5cfNQ4nt7+FVsTnXRms1i2IOkO
OqK6K14g/YD3guTTFGnZ5VYQPnCvpDNZuQvDB7bQh+WeYmTl25gT9m/ngy/OUn3r
fC66hu1pfEdVx8a8DlvHPW8KSu4KHaeD72+pZGEf5NVq3o/ARsAsygQGpL6MlqAr
FvPgan43+eYsuoeN2gmLyLg7WQKJoH3/vjq2ryOWglcS7CwokQThYPJT5ipH1A/Z
HDvsd7yk5eDXzo0NA4bSOAhOF9REe1wUlDrOFiOdRlSWyhHs9T/XJiXthwsvxCvf
ItiX89OH0lK2zrvNeQ+VoAlYRvo3weUudlZ7z4/xboOklZWCWeH1qrAmRoO7jzdx
zO9w830GGiRx6GaqmDCFnNmWYMm7R5CYNbyao40Jj3plOEMAp5xpRLutlluCpkA4
wDIVqzkhnexBHjYgGQ8mmLDdgAAyj1mmU73P0h1h8ZBkqnnJTaLbRGsYiAgWvxw0
4yvAy64z4JTDBM2mOnuKFQqSFRpTB83B8tUAEXLdVFD1aH3tkhvg1eMJG+KLLfSa
YZ3aVEIblUNF34W3+KAU28J/t4qAURTrW6eD8+3pzwpZrfXAirEKOQ/rLlC83ecX
iAhhPdMfrmo/vU831jYFJQS1aJog5/x/7wFUsk5I4qBJq4PoC/SIDw9op6/LEUx4
4H+hhSG4iav/MMyD5mMua03qNpN1Aw3cKu0uDzJmyMqYkNmbPpKWkTPndmBTA0oV
MMQz85edEg3bFVUNOx9zgwDJfZvjPeo+WumB1EJVlgHSnxwHVIJ9u4DmQJoc0Uhk
Dfvnxccb4iqQ5pAtI0JzcbYdLN3Z+izFCR2utmlt/yPtK1evQA6K7dNyo3N5fSbu
6EMUQeFw2S3k6oo3DuR04Ij4/WhwpDjbkaUD/BW7H7kLhG/fP9/Kpuvz8ELTYRLt
viTWxdsjKosmVj6a4gQjOPEW6+uTuwYfI2eCha52kkGek9MVy+DLfRZmWxUlE8g9
wvi68SEhqTYj8gHKdQYAkq1LDlbhStIKa2ZrQ3ciS4bYfb1h7q/Kyww6/N760EFO
DiIgt3+9zk+s3U0i5Da7H9pzXmVyoQVDc+a92kBKy1KG7Ibmc/ylf1KPrmi9ESZO
TsoBLbEigcvH9rdmjsmOR4V6cocb/h/2YQPsNG1i9sMwIgVW/ktNqaLrG9TFMUE4
0/UbdayPIAANjntqAMhMiAHNf7X1hP4rDl31t7m1tnZNbRw/ZzZTHvOL9VtriUlp
g5/WLLI4++XLznH3kp4X2C3o0ghgD4aV3uwHZJGr5GQ4CGuLVAVjMVN/XKJdMdJV
tdAkXTfyAK9l2g+PgC/xWXe58wmJu75E3E0jMKk6htlYZuGwBjS8VI0QUA8IGTWg
HiRBGivOega9hDUuZY/PvJ1EtPV68upkQ5zflItwR0Zleq7uUXnpkDIU/4hNgoy4
Fc5bJjv3+eYeU9l/X5OX96teZ3MlbAtV/mbLTHTweGVw6NVqAp8d346TCbKtfoq+
UcZAQLU713ts1SpNkGc3HF8sh+W23uU1pzOPce8Us4mYCZRwhcb9HTHRxNl7NHqC
0cKClesj492yhJeVIlmoyZ4BieXFV49nwA+0X3JCqCzWHXKC90mr+EGSLEpYCwyj
iMQrsCWO7GFKeoE3d+JYOPQmknGkxZ1yYqdCcw05KJMe8iAZEZtcYvUIf5D4Nv5b
JSIMLj0u6YTl3RS4sRwlME24bR7kcexT7ytsuhMiBQswPG4xZhzvK/R5Q/1oGuqV
UJ8NY5LAP3sc7tjxwIDkRceEaK4Jvus+NC3hZ5ejjPX9xu3LcigMImhA2zC0nba9
PIl+zRvAktR5W9hx2WyHA9HvMViOI8EOzgMoQl1msc5gXkcH8BbU7ZSkHZ0TdPC3
xTFFVFGAg67C7dZcudI+BqaUD6fPL2f6SD5444rt4pKA9W/X1zcnLtS2HkaAP9Kn
xF+4LAVwEYh4kgJkOS4H2+C26fS7iI1XK/BU+ZVPNxMUjcmY02eLOaQv53RCN+39
KLYTDWa/oOsRtbj6zKL/RGExvrU39FkQOCoZxhgd4Rmwoos9BINvApqiRTd0nPX5
hsEsZ1i2oRILq/wCJYDo0Fhh2L17lsrcTiYA1Yw+g9WBOPbLD6BOrPFJF+Q4+4jL
QSztxW25F02rvP0+dapDWy9dPxpVE/fI2OgsAB9YFQjJdBmt39Fi1p5QGQvBuYEV
QsB4YKoAZP9E+5tybews0a9p1Xt80oNj5OtZOfx1Sp/0lknIbzDTtlsuqFEswnxn
Iv9XkblhgArlFrabx40X0BWHpoQatQt1iaMaoOYmzlhnYQ8olFxHPNgmjSYpkkeQ
7x5YIpugK8IH/T6+/zO9eP4Df9TnIfWgNoWfebwKEMy3uF0O1BTCQp5EHcJ/gfOc
Y/+ADgeOCvyEmWkeTBZc3KiUegs/4Epg6qVFqMOulDIo5Bh3TMEP8ktsSmV2Befn
bTGCLgXuVU/ZVZuqfjO+eQeCJ10nXvXEGdCkSKYA2ECISjqw3HhSz5FjhRnb40c9
SpnZeKE+ZyNwpUf8a8aZIH70pavvfsVdYpPnkABaAKkp43b0vzGmiVA7VzryDhP7
pi6H0LOoA5WNuaSJa2o6AQ10jUW74P1Ixp4s/vunxCfv79PaqhFZUOGUvv8hJEEo
nhUezVn7SqnDmXBGNSdpw7xwGu6MclT2qlqyWpTHVxse+9kEXSHmO4Sw3lLVHMFD
c8FplH0KIqrTGoyfljMwP3uMrKazxE3EE9/y3HP/tpVoyXf8GU4v4yhEDUHVFkt4
oxpdWtm3WaaYcjbMrvmSvW+C6YQPcYvljVH59/p1ToYB38zpzX/Mrl4xAzC6TlG0
rEKqMl2U/gP2s7pX30lOdGOPgH6jUIfyJzgCTMpPsi4Hlc5pPB4eURVppfq0Z2s9
ZNU+KdhzZuIFRkPMSCscLNsqAVObmH5zUVIxfTSnwPmBmaU3k8cAvo7pyo8xSSco
eVPnzvNEcoIfIW8Wmvlbzl+a446ESI4R+XfdFRd48/Q9VSuUmKY4i3nWvzGEZjLp
Qg3QNdcXv59YJCAHOoEwaoDMuU96sTw63p0u/rC4u32PBw/r4hKCDPgUetPnQGNw
xg/ZwbVyywcGi0uZCxq9uu4kmcaL27aeaEl059uapehnAok0ULwgAzu3r6EEdBTK
inPzuCIMXEkvJuPksepLRajkZzCrzggkdkOTTcHol4IRy5moUZ+f++tcdsbuKDDP
CHhDudZdcrURXYxKl67EYULEljR3drcPma+9HDrQUu0JmQR/U34e2J2ef+6RncZg
LZUItjWuZCNvcMxoH76Cml1je5vwzRQBcRUEWTjaqv258wc4Ie1GQUV7PJ3IOfSp
XI7qOnUu3cB/qTtfyz5vp32O2911bnI4l7ehE03DLP5Uog7FmuUS8fDdqByo1dsL
vx7ut4ZIaftX/yV9cLJ2fDpC5zqcE7sx48qDxOuLz4hjH8RXM/NvW4LUaIc8GmMH
CBGWSDWc2WcskdF88l+Z6ZcpZw4SrZomSW13VKfj98TaCo6Ic/nwjwc7cUi5g4Kk
M1DsrP86adiWQzxcSrAuxStFtaLizVMqjZrC+H56lt663OSMup0yRiR/1qAIukcs
dkPOnEXwWw8H7obKvVwufuAU1D1xpWbpUEi0ZrrlvSJ/0qdV6Vv5J9Fls1ljulZg
mZtmDnH3GYj8qrc7GZwmW7hgjks8zRYh+p45wdsi/oplvPf8S343LrzHKQgTdMaW
XkJrA4+AcHUH00K5dM+xvpoq8xx53mrTox4yHzgyzQELeK5F2t7uNtoTrzR1OLqP
YVWBeTAOcDoTouvu1htMWGcpNTOhjQNg8Ly5AuuFXmVD7KZlAMtoqYwFKwfb7R4W
z1h5GSATuuGop+5NSr1VL8AvqNi0Wi58yVzLc4fLvAMbVCjUY/t5AucvnCC+C5dK
7chi1VO50hgfe7a2fNa4v8CTczqCjnNZKqX/TX+5a8Mpgu/YWP5RgDU7359c4ChC
eyg7gz0cqhYFiVLFkCchK9+1mbEIOfmaOjmJTDEz6HtpDj1hca8oXXYNgzO1ZQTt
9Dc0egIpMoR9gjWvm0C2lVMQP0bv+HnTRVMXSCiNsByi4r0dLzwHwjbKAQ73ls+i
pWbJARizwUlBTmoKt1BJR+ryzSuHiYVkWZXOUhcqMVlZw6Rkzq0tcLIxOK0fVM8y
70G+AblwYV4E9CiKHhqQciCKfMMPd/BBgexDuQki6Qa1ziVO8JoraLthGZGN0T6z
iLJODQ46Tb2AU5nx+w3NBfHCvUPwDx6mUN1qKhAWCtwbsusYCjURdlvWQ9XVNS2q
JKN1UaMrp2ZYWlmq3i4YBsO/2RHd7yN+nhHCA34BAC4SeAc8fN/28cjUtHGiOetE
o+FaTBCuKVuvQ2rvWrUCU2LFx+sNGrNqSaZn48bo2M59YsA5c0yliA/79z+7awF8
/0VckiqupTGgo9HZarwA6b6xFBp+vnzS1z1R63h4VHT78MBTA8yyC6CKyKkAVRXC
HQAiIbBFPcX++Euy/IqT7CT/+T3jXxt8AWJyJr6qJVWT2duG9b5lRFYt6mV+4GaG
UmlThWazylreJanM8MkNtHkZLtCB/cvOgCwy+9YCrMLo7Lp1mbjGz4Ffm65FzJwf
lQaaPrsxv/WAAazLoRqSLfL6XQrI3xH+WZQpJcDVutMm05gTJT2WHYp3GYMg+t2T
FwSChi2wZc+t3NXrnUheGyZqrId0wDutSDmcSoWO1DkXc+OZAFHmpg+CtxCfBrLS
DXAf5v4NcOIDP+CO8aLzwWWl3UoWft2NiFwZZynSWugLzS7fiwyOcYh2Fn/RYmfY
cMMCatofwkqu0fIo8rpFdeXyXq3Vtbl1eL5+GVix302lvlQ5mW81eCQw1RNaxzCg
JHokWEg+kAUr0e7BDuJarNNJeTJmQBlzLZAoOddlPgTTnRBqMq1bTE8WrURZ1vqD
y2WepUBh8ttxiGsSwA+IhMeAOvRbaMIYKufci4ourI9l8GCbGu2nValfo6nZEmFL
pMKxhZTMejxcRMzsySIp/aOVdxa0FaiAnj9lFX58vFWxaOVU3vgbP+C4jOVFy6rB
UbfwTLC//M1zZZJTydeSuPWPpSkXfpf0JP1LUaJXH4v00YcFU+XKLedmChJyB+zE
LjMkSxXNrROuIaU94a8huV9j0k5uMNrG//eDQzdvMM2CPTij0F5VKpKGUL3Os0Gi
2dsJMYgCX+jT3A+3ydh9XJBt5V134bUwW2dQs8EUqilidJGxOH90ARw7D11NXWp0
urAPYcGjtqkaZ5BSvWvCL8i6MmP9KiQ+I91x5qlJ4goNznIOS8Qv/HlwbfXAVvxc
BWOQ+yqydwS7O2qrxyKTRvpsCyThKXEIWwCHfYY60gbbe0GMP5n2ZfuQf5TJbjBM
n8lwblX1EnRSKlt6SO9Kzl9iTJBP7JH1C3bqcM+TZcxE5OcbOmlD8vFby0Qwn7hy
rPKPFNPExgk8n8hM4xst8CZMmCC2PBZoTNmSxidZYNVxrbsUOk34sh09uRPkElVk
DoaaDmDDMknhidl1mCaU4b0H/zSAufM6A6zw0JDPDU5A9Ctn1WR7l0QrHL3CNYFN
U4/UFUx8dQX5cACV6EiVQuRObwqJT3owNpecxWo2QgiYi3RigR7Qx5PdEh4Tkc6l
uFRtovgM3PIgHI1iC0T3r5wZ7L8TvTPRkxa4ZlRsGShJ8CEjVWKH69T4a12XTqfF
c0PpJMINBcP1ssdE+7EPxGuO26YmhHyhJUep82+iNDbqVLPqPqKYgx9SlEaf9Nh2
D8GFC0fTupaSVNz0rdt/uLUUBGZA5sonToVzU6iIE8P/ywNpP6KpUFIUpFx6kSsv
vYZRtbdoEYuFN4mVFe5mQjdI7TOvzi+EWNoDJGkKrDgFGVq7L/dlnx7FuHRWGJ8E
WHHshkypFak08OFl4xSxMOmIiS7fqPOTivxon1lhjtWnZgV4IHuHquppKw1Ijj0D
akbGwe2f190DtNZWQVuH2fRIb8eIivjF0n7XCq0R9mAfyOvyNCnKdE1IFTjiOR31
/w+F7PCXuQm784GuKz3WrH/gnrOyCq1Hx8VnpvyFjaxCQJ/7zW15SSWKv6mcaOjd
kiRbbbTbf5aFH+6/zPqXcCgUe7HG90wgA1Jz4mMdWYxJKkE9zP/5wSpYm7RRUpYL
tpltd6z2HF7UfjgY2RMseWGEvyVSpZAQjyK2qEM+wiOWLbz6NyXri5JJiyOcv92F
8jZszxCrBQHh38PBnvzXRNQFPoqIyt3J+TPTo5YH7DTPK2R/w1fN6dsihg1IBrAq
c0pfnhMAc0uFnR9DexNXoxms3leMqdA2KoVJcZYsw36vN1HGcVNHCHYMVicEvHAm
Fnh/UU0ICgd4Mr0A8jZ6vdADR1304SxMMPtCccMJV+6iJDkyy7GyaisBksVpoxkq
KqmY5BC/JNoz8ZLceP7FQCS88oqxPj3UOpNKoPW3z/dfxoNESDV1x2iP3Fgd5dbi
or2yaLVRUoejVGSQ1GJtYGICCB3J5Ei9kRBw/DF3tEQdHY/hK/NKKSWK77OJY+D+
duBV7cVhSD/HQlkgHVh+yIQH9e7HWEIluLJxRzVkKP3ZImMTDJUcfJBG/F7EaP3u
2/AcheINQ7P5oybhzaYQY4N5r+wO8hDgV85cLalzVAsRSg9My0yAmGPnlbBniXa9
dLBVEUMiTb0NNAixkRMREAiWKnm6CszvRY1miYfXfwwoEw86m0X5mkSoOLNBPBfz
EeNdjkeHopHxVietkhjbT+4XCoy+ojp9Wmrbb07hc0NQmwuXs8jmbBJrTJiBWlwM
GrNMHua18cEBd6BGPvDmWlv5qfV28tMbefH660SUF+Y0+VFZhnsuQz4563pn1xCD
tNx0fpfZKopJF/KOiUREOX7u7ag/ZT573jpOMiPfgoygui/fBjYGgHudF6e1+A9E
Ya5FMc8EJW+mkFcUxLBdo9bTVWkcKJWme7lRtbmJxwfrCq7DKgvZVdcawESjVrkG
2UelmrRq5VjsjfJO+Wlg8rlclEFIGpBayk61slIYFmwSNyxlQJi/enIIOWhUfUP5
tYGoBwZVUiQWkTLFB5aAPuUMJ0A4cY6Y7nT6nmWP4g9So/8xyiC7FepeZQUyGqQW
aRSWrdQvLR0ljqy4ksSUpclOntr1zaIUnkSYLgH2wuEuBQ6TkFZkT9eNe5bwuqdn
b2igTP+rnUanok+Rv0ENJhNb7PkG1w3ZCThylwiHfdNEH9q1f+l4mWfgI6dfc+0o
6Wra614nU4TdT/JC3uIwc+1bKe/1lpIFkbD1WBfHqS9P2kJoTly8MdRbp/UiRKYx
7mtDBzyIWibF6nS0+zTFBGt7FX/FOdzJDLX0iuYvBqIYQrQK3ueZtvza4/vtRVlo
qMiYZi3vioL6nzDOBUUVEuS0SWdVpMP9fvjRMhSy0171wwf9DWQNc3vO3vEdw57W
KxfZ09JKWHWlAuUsFbL4W6Hj3/h8dOnoUiTWp5upe3GZWz7+wxwR4ERls7U0ubhZ
UhV1dOHWLC1RoijUxm2AaU/ZEsWB0bpwfQmZwnl9iGxwHo+kClcospRDxyD0UD4y
O4wtoP6HHKKm91ExlNzvEqAQwmZvsPKqx3bLvVjucZ5Abar3Q/zN3hdt5zWi/qj5
8cfnR+iWhjQpaYM3rU9Or9d1MGiMwm4y8jP0ZQdJI4ZorYAmKczEH0dgRX0/bG/i
jHf+jsC8kJoqLortr8qGcXCJXgqbNJKvazDzO/MyO42d+7OhXSp/vtfQVdfRffbu
+u5uGRHWcfuQfwgbrYN1c3rkxkEGSIekEuWjiv6IL/SR2PTNtjPsc6ffoSPtCPKY
it+AGc52Sn3qmqXJXM0DcPhVLuy2razlraWpFToszjfxtlQPmU9q+nzqQj2HQXxD
kBDLDQ4VoFPjL9ANvm0TP8GA1dHUgqLQXu11ML57dh0MHdhFqMlV4Do6DtQNBe7F
ufYCox1Dup2XYV8cprRT8FQoaNMreWDl/2odCc8ONTZpn25KKdmdwEGbfsP16rCv
1MjCzUL+9PaANGmKiMBnc1RsFshIsqG2ldwoK63pVtQsJFQavLweB7qk29LE9eW3
5Q2Gbs9IK/YWZPlKyN5VAzSKXA+6Onlf/1LA1+hHQFhu6z5eFMfvxgoVqIJOyCgB
5G966RfO12AfheUkn7QGqVt6RhdK0ysS2maLXx1DRbui43tQ7CQjpr1ftXxzxewE
CvR1NdBYSufXLQEx4AhvmAddlL4gbiSfl7krAlVuXAxGzhTJofg8mDAfkLsHRmyI
aA3N2LpG/N/wCXRaxPJzZ8GYrKrlSu2YgB6E/kLDC0rozvJdbR0ghNiPm0lMZXY0
qS3nkexJMWj8HlHa3Ui2sR9CYw6hIOtr9AMBXhEGjpOmcXdyBWIYQ9bB5R7Yhw6a
Day8iHriArKrvefOzYCb7rTfpmhBU092KolN+3qTWtWfiaUf8XUrSrkGWxaEL+tt
Ob997U1wVOCHEAjJAcV/pilBLzEkfPsVK00xk+P3+WVVhWPfRK2GMZfNoLGo3/Xc
a843DYEiXn7HAUU1t0qN+dquv2DTcJJ7BOGfSxyoj1rBN9du/dHYVj1EY5+HNXKY
HV2fbtj06Lkz+UQV04weSHMM0aC32CWzfAi9HoieBvOzK2DqWzhJjxGZfQtstAz1
QkYuz62Ur9i4ZORfm+VUqCDn9YBFrRYt+nJATX3JyT0cs9twWaRbu2HMv2HzPZef
iYyXOQQePiKJK2gznrKRj/ABUqsmeDIzx8bQ8QVckm+u+xMlzXJgJvAuro4KMzaa
/sbQ9/ykBbi75ijBNHUKC9zRR+rkO3h1KLphQuNZt+Q/yhNi+Us9r/kPDHERj5V0
sneKRMk6Z77y/SGzFJMrLR3u8GxXYTvJK6CDVPqqpjJr7BhOQkjZHmLtbVVp01VD
/h1MtnO4zw5cqPY4TvamtxZqvulr5CFk1Kb2IWv1jiEipR2p5amf9eWVd4+lt9at
xFB9bzfYjzytxhwTtK0nx7dBFAm4smeC7m5VioraDbKgZ30UsyW4Zk8pwli77a/1
ogH2txLH1IoWRDS8wsaeRFuabdQkzRjsr3YRsAVUMYtg0FQ2YIaa8LzUyjLnlFSZ
hvwaqq6QLCxN7lj/1NfyNTmahqkiwWwNWnHwbBfPzzkvzZSCf7xI/yHilQxTbjFX
azWP6sJ5HbLzfoWU4EwFv3at/mo/LC+ufhuWCUOC4QFCGGRerwrUkKWLH93KinZp
vXNX0j76Vf+uHEF6gCCkkRKX0ebMXdS/xYJkrUswlGlit6l0d45Ie5dRLBudWq4q
Mi2QW5fcUuZY/pxMNlwVOSmyEC6QAsmIj05ErG3XeuFMHlG9sUQIjYKUbE4yDbao
x30TB2Kmw9944rbVgb1orPfhrHw2kEIp86TkR2+tzJgr1xVIDTje4Ub1XaZfC9d6
zOToes+tL2l1O+x6/gNSD53Bz3udfQMqO5BasoIFogngu0gml5L32+VSRSzRKrsF
6Vxvvp7vzGzn/eVp++mDDBJz85eBjblqMw5BaSAIhOysuVyFAOVvpmv6d3nf9u1L
g+GzG6Mf2WmyHcw3LnIec/0rfBr6hhIJTrfF8R/tEAEclvtRd8z92D9EoJZ+EejQ
3Cph6Jn8g6CpwoQZxwEYjReb1FF98RkCFvEjMY1/m70o/zF5sT1lWrO2/fFzhWyL
g6bhVfXsazaiS8r4+joW5QGkU4taeiLYLV3M1HDPsIpoxhH0KbAOIivUKAgYzUhy
gY1QaOpJWs2htaZvs5bmZohjnHs5nwssKlM499tghYdyrkpAvx/DSCpKGZo81vOD
tsEu3O5/g19kTGZ2vWUDFaafChvKed9zdLXjVh5bBnBDb9xRQth1WL+3um43wUqw
OwG0alVXERWVVUmqUM/8gO6vr1D5YeT742HpX1ctNBFOolB6Jw3Bd4htxb8hBu7S
P4JxfHCKU6FANENmj+nGNMaw0x+0XnMBtO3F/7dLZpD7wkAMeJPxwlH/DXZdHOcq
PC1GOjSNJ8p9xZtGYs0Upn80DDK4Fsl210rmleWXulxPVAJNQ21KpJFg+89UmhB9
hXI0Ihr1zdJiMLA87uk8RwOi7radF8lTCScnMUVFTGReH5/zzkvy+oY977VzgaPH
xF4luk+JmFHOJa3QrEucC230IHktibglj3X+Uj72O/5aJ4DrTG/CtMmnN2LVFPhI
3u5ZH1OzGJ6ZtlafVjdnYYns2ytHkGGAi9x5j/na1S9tpD81b4SLezGuFpwK2p1V
pxxT2Tb6JxRe/b8/lpCbAef7AcQ+OTt5T1Tkq1/oXrr0TfAGOKSsGB2LLAfoGtmA
O2DNs3HpjGNtq0gDboslrXNLopcROU24LKntkVt4XTDrawkv0bqv/ljPoLVpIlUE
FzpF0i8O/EQnbh74XnlKGeWpHc9U77nOHIOu18C400jkIXDwWTqGYyaGmhrU4pfU
joZsd/qR5FCWzBNUbED1EVLZeE2Jhy1Lvjqb2jDDrydibYej2FzUSJ03sAWJhOnl
jpbczGb9AP8BubarwBT2EwyFlIqFQQbR5DcoZEERvj2kqR4lZG6yJSl8nFeMoB02
8PWEf6nxjcsFcnFTgQ7GOk/23pk4VRqMtOCwnI8DEGbZ6Gn0WKhQuNS4qIR4E+Oi
tMgqiLoj4tfSjeDjM6jifFqseX0v0MmeeUkBeWs7iuKUKSkJP4PFwKXLIvKl/aXR
MtkBMBv2jlQIhWWno0NYjm2LzProKwMbZ8+PJibKXWk4MruPnjhIaATy4yYt0htb
r+tZaEH4QLVMUYW+hzghBdEPAh+T2ysIRbIACf5wWtHWRNqDT+CDVMwW19B7clMa
/TMiZbtW4sqeA0AM725ar7g3q7u9lP7d/XL/vJ9r7PJqSwiUN0lGDNqA3D1nQKLb
DysrrSW6PzMVeSk6lYF+MFXBbYH5SYXHypuNYglxBvqiGqMxsb56eTwHnAwyU87I
wZfA4FL1eceVQO3Bu77g0dZUNR69sXVFqKsvKjmweXyn9eFAW0SuNXroEms9JXEO
0oKr8lL6LgpwgrNisK6Is233HHdd7c07e7otbeAaWsol3S+nuQyymJsrkyR8tSHt
F8H6QLuhuFLLzNkHQXIVADj7QlpIOV82vaicR/oqYVZizEPVMV1cml6XLDUG+Oo1
2O3YDT6ECwPJQQQkzrGSxLaWlxWgnqBQb/W6fVc6qH7ngRJmZHq7SdSrbFJLGjvN
W4ItwUeRDiYEMIrGmTQidG5O7rKy5YqoXHadhzaqkb9xyU7jFPtjGdjDx1ZBNc/f
92Ftfq637fSMQpG1hWAR7mXo2T6P8lU9XQFc6B2aWd+ZZ9V/K6JCjbVZ1IR41YOh
SDJWrK0Ywv5s+vH4RICR4hMpTpztWh7IF4KjJ54b6OeA5QHswEXomAzuet/k94fD
+8lQNpi1JbS61fp9XBFuufpHtjUPMlFR2Mel6aHrYcyRaqLDdFMb+1KfPZEV5OwL
UksJ59rD4yulfGDfZCcXgH7zWRwOu4wmO4fvbi6x7mhYZNOo3Nwc6nuROSvpsTRq
d6l7BrV5QuTfvFhiJhxxL1dW/bBaAITFBwLBK/LmhXm7xJ5t8QbwrKzck9YVhxzR
pEfb9rtBrj0gbN/cCcEI6tlBSipZcjOTfguNa/gC8Kb+5LNt7YV7zizF9+4N4D8x
X3cTTPCbjuoHcr6fZcFcEpE00Ukt+MuEit5yIjkAGp73VU7pjvziY3rGC4Y3j7Tb
P+EFQiFkntuvSOevn3t2mGaQVYTMW0dzrf6AfrgRNdB49pqv+ox4u+Zpnsby2Azk
7wsxlPHp3DixbNW3iCsYtYmoCnejhoYjBB90q5a17cAaYl4sbc+MiWOXPosQvjJq
Bw+mMEjCqcbabKhtlVc5+ChNSYbLI+HnFK0Wgfp3HOA9RaszizLBKrJbzmuBZaZE
7vVgDN+1cPmMpzgEi+sLA6lrwmTc9/x8LyPqyIS+84noKr27zmaNbhwmLVIDS0Uw
CjUbVz66uvsN/TmB5ydibm3Bob7WhXluwuRmDVSN6Nxjyrf2MoAuZEWR4vUBzQ6u
52c//QE+y3+K6izkCALe38xDJ3q0ddulNEKnhOsEC+0C1QC3UasF6N3SwSwAxDYX
21SGaLM6HXcAGLnj/sg6f/3gZRclHUpoSRNXppcOOHJ5uZCo64Vg804pBkOcbNBn
TZm5+5YzPdMPz0zXBkHN8w4TtljJ+REH69VrPf0HTmc6Czz3ooMlZKiGqehukMis
0Nw/UTqpVwj5I3UC11jBwAreL/cPw3aL7qgZNJUhm+KMXPXMqmFJoWiOLVFZ6r1d
yNQWCgBpj2vT7thGXPezHlkkkid1avNp1nmjQV0VryjNnpiZTuenv5A0l5gtDXYS
IMGHZ8rn4YezIru6Gp7TJjezWdDugYRwJVeJG9rPGLxpngmJHNNO/U56X6pTy00d
2d3c5Xnb3BtNh6bw9fmyNS3/3B3isC5RbSJH3QG9Y14HMUOUhY72QnKs9jJDVHtZ
RyQ0S2M+ugyVYf8PL+zlFUfLc1N1M0xdsiySua57654Qe7FAh8MPG2RTf6YQky2A
3jyOs1+xWwtZnidvQC7z6MVdtvK9GijnUAXA0SEb39wfqS3q0381jYFoUsSVUnvg
iKdAAwC6MbYB3LjOwKmBLrxOWGOz0u5e1nyczGSNuJosmfnrOng2syapO+IO7n9m
JRHLcSl7Sk+v5ydE5xuvfHBF5+ArevusjIx68oplRrqeSqqG/WKlcGnfYOaYLj9r
08Jvpa+024CGIxD1F1mVv/0lbizRdMRZo2VorqRLuNFAWjunnVpEZZIN88tz15nk
RXy/MuTEJJS0Q2NEZBBpaaYnezFiOj8IlljNufemlaOhoDVb1uDm4aM7kRt7XkZi
FRZntD3d6mVW5qvn51Eo6SdcGiS7E5lGmLlQ4hCKOTv/pDfRZ9+VRTFHbBHxHr11
oMwyYj0IXNXTNs9LgS1fRcftlaDJBM+bgU/Foddp/oY8VUZ7Mzg6AAFMmgxYk+2c
5NnSTZl4GHrnCuS5TrH009/NjOSp1wB4DquBDj0UE+8Wfid2dtGoqV3r5zfu0lT6
kmQt+s9PbPthLWisbF9KSi5v+S4A6+PhcT3A024J6meuIu0BeatRSb7sFQsT5RpJ
glC3J4n+m6GTJwahjcS5EhV3nOPsUVt7MkldFhEf3t2Bbhejx6RYIATCazJC7rGQ
yEj/O6vcmED4FSZ31/nqOCAUnHlt7TzjMMMsW3UlvfidUsmaKf0/8e91Fqf4h2ss
h4oCrtRGHVN56HLoCy5zH7iHOzPnY/kFIn5+eg0ygBIwEARgv9mGwV1fnVgys7AI
5R70ZVJhhGjL6FX4Sa2FvUmq/gQT1u3xdMZbU0okxVdBBNf1wac90qVmspZ48mi3
Lk6umSSdFdCFScOFzx1BdpJ6f5lXtTWULypG2dl48lkGOMSm9AuufH6MepemF0WG
MWOvizdMEWJu8OOE2h5VJu/2BATOOWvIfb6ovMQRkFAXv1D8kvRE0+knUB/zaBPN
okDOSgc7BXclkYN8XyncXZowYsSn9Cbe61XuU9qJmVSrW9/I0Un995anYpsBPp/U
pcYGk8mo2GlwSh3OBqLMKfuIUmtFTlop3vb08evThoyLqy7/BxVudnsEFYrAAYpN
ACyhvY1mlQ7UmgM2hYOL9hoCh0cmAHHx6+EWxmLpwR20+E8wmIQ5XS/UQ8I8CO9t
QEDouFgQvTwG5WECV5ARK98OlNfkKFilR6Qy8/W2cTeurxQ7JoCEVK173SFbbie5
ET4TAy28UsAg58SKVGVDrkZvkoLTkFgaTYPejZAwZ++rpMJsM3B2BSr3ae4Zu6s4
/tQAYj88KaCrhgK8z7iw2Ed5qKRjebxCBmi6G3csLwivKq35LE6W+Pj7Y2MZ7l9G
a24kPEFyzFLsfZD9Qlh7ph+hoxHmgHqaj1LKxCpa879yZYDN9FJAiwmrLDJNhTtq
TZqccOy/Tk3Y6hAlxVOGiVCmX5BpNsQG/izCMR9fGwHdL+VQFcK6CxhrlvTVsGF2
BH4wc4p2IlpY7al8DzyskS1SnBlm3JvuWdVBeya0Gqs+JXMaZ1e5RhK10P097RM1
R3el7BAxA9maUSAmOFVHo0YbS4yaG3mN4sWxTuDRxIXG7EIkwSO8OPfdgzpVnr7H
EtNfibSmod5vJhUAl8C+99AuiHqmrpJR9SuEMHgTtytKZTK2X44NTM+FL9IBt3Yl
54eZqFhxKMt1CFCFVgeu+fPBDIyGRtX7yFo/+6Ui0+CANLoTy51JS9lom1tm/QjH
CKunTc25Jr6zyyDzcaCzdcVm9YjaOnp7ETUurjnOZ51l3ma0KUy4V4tIf0ALjQ/X
4VnesU+mfr8C1qzwUwuAGLA2QYmloW5D5fv85wpQZNAkGiNLa186kzRJHIpUaxfv
XKhxQuSnz+DcsfM/zWu5V95Z907onfb8dyeCU+0UMl5z+7fzA3fwrbXd6syWq+8R
kedpzKiYe09F6H33I5aSqD2cv0ulC4w0+ni4tMysKUPkc+S2Qqiylox+2uy1WOeH
WCaGemEp9GIS6Oh5U/AirlS7dq7TZRddUNANygNq1aJ1KeiQM2QXPOoBsL6fF0ZW
9G2/aiQ8ZDIxIAYPdnwoDL4gGZYy+wUvgxdf8JdEWTESWbnqSiJG/QMySXRsmroO
MHJwx3OlMv//wg+Ds38wN+sj8GobzaC3aY+h4VS+2iyg9tVifIoMdz1N0oxEjog9
tnoPmUoNlq3N6FoEmEtdLSYjfd/QuV3aV1QRq9asMSg6MhoUPyk6Fj8SZvowkUhe
BZX7KmoO8/PILWBUefogUBAvkEYGTbwySjPgWfuaUoOxE96eLbFOzVB9aPSejC6U
zOkMAYRNH89BI8c09zWNuABnqMfPlMAv/7GEZQOpWCvir1MycCX3SlEc9iiZ/5KZ
2RZlMZxT6RSV5d9vFCMSLtZcLVVayKmderM/RricqHETYTnmbOWaCMnvF2e97YyF
/t0YfJoKtovzrr5subDX6gqRhpmH1zouyL1XVirIoV9kSZcDLxOonWIs2m7+e/K2
HJRHFlk8wJEJ+Aw9nOLTiC3rmEloX7ZKsXFtLl4FWOn7hFpEnCestzLV4e8MK7q0
jIEbgsGjyCC4bomPXS2CXpARwYb0JISmkhQVIXkUgQ2GIvxU8ionql2TJ/BrUGp/
3IUptlneimQjFPBtySeZDvBhJ8yfc4yvbOQUIWWtDxK2vbU0/ljmvs40sR9IrW8h
Pgi4uGteql2EeMjnxkGM5SnFclWEES9TP++gkkyBQV2ZNEN4h953+13h1YIMzADq
qIJ/j08MceAfqs6xNxdNSLJzdI5rtIs5lq+2eGiDLl1opaotr1d6ZNq9Ro7JNWX0
Gf37C4US1pQrZP2PU2P9c5rexoU0v04kapX/qf2YPLNF2BKd0exjYqF0IzVjKpbT
QRj76X0i6rUNDhFh6sj5bpE0nFXySt0VVkBPJr40SPZl1slfSn/WddWD4e2j8aed
2O+9SRgv30KwYvjVZZixc62iSIFwG93W/sktFzYo+Y2ZUd7ZDm9Petz8xjxGPdv+
8kL1PxHtgoqw5GV+//o2d93XguvwHNERtfL5zTIepn2xpkrafNCexp5SjvaXjLvw
SZHUa5pzfw2X5cF1pCD1ByIWy0iCQM6oHkjCSdWvM2ZHpr0fIgESc7dLhS0kUGA/
z6aDw2Sph0+FzRND0EmlCrEkcK3368+6cgGDkFh8IY/zqa3bhDccbJG3wmo+23ov
HPRpEBbqMqoLm4DfuO8Z0Dnl7OKwlNOroaMx+fuk6JBvr0QjzVW4RALCYjcmQumL
ojI6UygKLrzcqI2yOKnj0KyVwkzN1uX7qqv8xO48+SWJvcfpfDtYx+l2sW0Vevvm
bjZ/b/BuoKI6ZqKu1cOCmcseHnYkEZ5//5ZDQmFhGJjuedBZH/elWG6UzVahAmc8
rv1lhyScLYwZqLm0Dq06SjAh5sWZqTzF20C2JRUsbRtIv13hGoii5Xp/yKmthbZo
nY9hU8k2PqfS+hFSV0NsBlRj3gL0HaDBPzIxRcqYjk1YQ3yKXLNRcsOxx/h4Ve0S
ZnZVnqRAVObhpm7rA0nBbD9/Is4NugkFoA2L/Oru8NKBhtjhXLiJ2oujR531PUEW
vO9XdL77l4DhZZgwEgVEuuQzTzCIVWHAKME12lxO7q6vulWJ/LSzYZ9u/kJRdZuU
GpYh+AsVHX2cm9a7ZwxPKKsOhy5f3iPLbefKh4CLgfQD+gw/LAoyVSVAHNJjUS8U
7DFyj+px5LhCLaBxxYMeBpv0REw19K0WMJhTLSkmZdtVsw4SAQ147GiWysgzDkGx
Kp8oPIIVyjRgRlssLBbXmlvYNu4OljdY3zz/4Z1D4agDiB7DE79SSNXBAXYiX9pd
q8/BZoolOv6wZCnyNF2vf1EapwEAZG72cdrbYXK4/Xj/BZmj8yGOxLhwiPHA4jyE
VLEtoaIHsrRHZAODukmTJaYqxUgqUgUEJPWzGTVLY9L0kQQHjYLW5E7UW52l58HD
E6TbTTv5Qduhp01TmYGRlVhXY3rD7VOc5DovE/PtMQnNyFn3KP2BlfLbZd0JAMjY
4GTDZneT8Z7yRvZfPN1qrLXJTXXypXdrcBzpfF6Mk2qmNbIINGTEOxQMItEVo0Fx
0KIROW6b42yiEkpWd0S4Uvl2WdrPyMZ8jil+sW+HKJnOfUwM/FdoGjPvMadN3wjF
26ya3XH07UTK0tsjVuY5uZsXCW5XArin6G9E04d8cK6O7RoF9Yp3WyOhK2Friz+b
4JqUjn2l7AxpUXDJRZgAMOb83440Z1hy+dsUpOu8pTw3pCqVL2mzeGLUBmylmX11
6msQFeb2idoOsT8oCItMH3EBD9xwQvlou10X9QMbucBIeck/PXl7qmoP91a3TJZ0
yLO9KKsxiQ5Ff3FByIrPsyW8OASo8xqGaZOG9FArLDwra5zIDOUn2Kic/no5VYtS
jclNExU++QdnLSJ7rczBC8inx41gQHani53sKd8y7oAZ8E3d26JVPIRELpilQkrP
uO7thiVG4zQVoXGcLCAdLn1+1pPCiIAbO8xq8do45gfErQVQOCqakYwNjTDh9a/h
hHTFHNkIvddZQ7NPSriNSwnYMF3LBUEy6qajtpNOZgUKS/FhkenZF9zkT4GMiWGB
2g+tcLC+ByafS7wXRZuO/hsYWVi0Li0iPx3paycEFlxYC45DGPAmJEpf4+rIIsty
yTTl0dyxrLA7kp17hz2JbxSY8iihyRbbFYzZ3yLkqmuU2nxMzZaIJV1mmspvAjOT
wB3cGE2Wj0hxd4qfO8Cm+tqJFa5rDT8mWJBHfr2CIQr3Kasv9MFxtG6QRyX3cxpX
KoxYPvg2w2nqRMn4zoDXAAt51AKQGnEueRp9QV/QRsNkEQa2JOyx46F2a6KP58Nj
7xrBAesfQRub1JLfneVjBFQKRrY3sP3PxHTpDwz3ZrCSG1yQ91ZnsGzrZTLsuZnW
m3lC6666YFQxi/NJS0SOAF2q/v1SU+EDLHpHdeNy31qhN/fTZCd+bASABhsanP0V
3oV0CFt1My0dEZp1U6OlN+zJgUl1AZOrs1Iq4B/g47/l7Xt7PfQ26Tod0zbvJrsN
HMFfkn+wLCARuFmivUgh+RTuHj5Tw2YOV4GPLYvJZ+Og9tw2h5h4aASkn7LoC3A9
8R2/gKYWJO4ai2RXnEmHtMOHnesYkvc7Tpr/pDVYudfeAwit+eER9aJXgz1iJGpe
fdYcKhBKdDsWbenDGmU3R4Hlyv+2IY0O7+2fVR2khv3/ic7qT7KSluWb3+ODYuQQ
V8M6BGe+kl20KHnSt1GG8Nh4xiPLYbFslq3ZXewz/hy396/8Amp7XNKGvsY3xm7s
uIXDgTlKYua6ksfgkWGT0c9lfr0J9qi4tMpxqELhsQXVWLRjAGQ19wDXOnoEdpN7
yHoGFN/uAvgi7Q+GX1zkoICz1myks+yp/v7FZYRMdAhxjC9Eh0zo9zTW9FCmWjzk
nZLRBENtQHoDS81HIsgB60nt1lhpCYU8x+h98quGrHv2xoAtYkM1eOeT0+KvRnPU
KG6nKXZ/xyS8cK54WxI6YoH7esbJdpxa1wHfqE8ehCfuk5f3p+TPFAENurehs18I
T/CZaLLPmlqU/8o9a1gW4RrW8mHAfoBcrQMWWvghiGEGLeK+IrhJXOkyu1pUmsn/
bdqJUHw4RjjTYRjrJhcrNAOXTJgLdDyaX/ms3nXbyyNHIEQQsvPULJYHbozryZsJ
6GCav3VdahOJmusIuEE4fYVSFFulvWDZdbk77NEP2FZ0mQvA8L2hBRlV6a/SfwE+
cjiXmjhy17jH8Z74zdbzyM4YvUKDHeoA3IyJemFjfyofLBuOy2OuG+iAsBRVhs7o
2IR8HwUaLNxTEAU8ho4/5Tw3OFoHRfpVlmmIruzEwL6wZyc2oc9+KUuZVHiuQ73i
vhdmE88pJkRUudv13mrZdwXO+/fn9w/0DL7SVv0WlXFG0+y3/LoaACrjOkmFETsp
kr9SsVvUM/8e4p9Hx9cStjPzAfLcI1WKbv+lfPGcJoOKHd77TGP9RS2fFQqhCIcz
dqN+a8rfxXV4Xle3AH6T8oc95JlI1AYSS2kvgnOd32lKC69x6/Iffjfh+VxZdeNd
qnrkItdWxgptDBqbISi3KfRuwp6OSFsq0+8dT2ZbRd0jMkVVdHbd4ebLzIlZ4zO3
6eESjdSHoaWND4zyl6ZgUd5ekla8cvJAeRrPJwbpdqxSSq+Qckv35kCaXxwH93w/
8B7xeIywjzM/dC04aBjVf7VtJHO0flE6c7ZTjK31GVhp6iO4/kTen2ZmaEsdXR74
HIgGzIhFprIH5UtV5bC2rr3qwllVOOoWs0w5sUWlvgg8g/mwYrt3DXiAIHypbkFc
ZSiOZHlnud3Ll6E74olo8Wq/vCCThWTk/B0I1pzK0qkke0bBL63qOJqIkck4CRou
8KKWjVzzvgul9Jle+8blxxX/3RibL/88RCFxML2r9WXpm8GQtxrdGxCqT91XCeek
1qMSJ2v0EhuXE5T6LlI5VEH9cVI+5V7/d0oKJIjTlG+o+nsvLNM5H1DGN2SiSRXO
+DVQG81ma+9TkwhQISlVa+C/pq/kcS0RAlQ1ag83XxVyMvS+1BnF4rPH0NBHEUW5
Q+WWVBspLmVFuXimw4r7R7aCZN2fox2OX9hrDp92eaCutd8MYUiBnDdiI/ZcTEBb
NwxxpP1v6YTr8SWAXb49qWY9UyJLPoFc28oR6jF37yYD2v8pxdbMGYfFZoBIU8Cg
msSWr4X1113z/ZFdzdgMl4lg0TYQ9pywF13TvNXNUwqXf4jBDqfGm3MQog7//tWe
qiev6Qm3PNn1GRYJG+41UG9TYG+8Lkfg2kKjHqmMT7JdpOAWdJ94Sa8HKXJjzorF
8af3ba7Xl/4zk7+dctI4SHn3wnoHAZwR+hZ2K45vC+AG96vu76T2QjeoSFFa0HsI
dp+9z3j8eM7NDmi1vglllj2tzFqhLAeOnYYAtQQ1uDfQ22hnOHTQ84FqCA3V3d+5
HMNcdFhsjO1tbohtYLoJlom1VMGTZgbx+X7FW/LCQOOv5Fmbi4B7ulHcSvv04zNW
opQC/bc9HKdxlTv0RtsD+6sVDvMAt697s1EH9U6gBdbFx4FjCwHk2YlcFm0NJLGQ
uPvCYkqfKw5KhvX42ez0KZOUk6SC8O5Eszf2IQfOH3Uz6tA7OB1/aIfA2fq/T/1h
2YElYdu/00tORjmhNS+4fIOn3Kk2Uz4rghpOomnyoS46/m8pIGBNqORAhx7576/B
rauB5HlCowjE+RYJjhb3hMCf4CYIraeqrCDN7e2scXy1mwV7tWNAjFojXv2l4WBq
OGnrFhzMoi9/mH5OHMiZt8rt1Waxt4DzGCmhSyvsXM2wFkD0ucJQVIFKKmW4w7B+
YZQAi1XI6RMWdMsvEQMpteDfQfy5hg5KgOEsVKjaz40MAG0+yST8O69MblsKuGGH
MnBeJoKLRYtf3QYVya2vlmpCKggG2BE2zT60jot0lHx42SmeXp9xirIuJrvoH1gk
WjfRBm+jIAaTi0HavaiFhe+GOaVq43d3Jjn1sNnP+/JjpbyM4ua6tYbgTQEtHX3F
HpZBUxTjNTeQsf0hwNlv0ljWqr1wIoKgwA9AHGHjV2gIWTfjdsSyzUNqDFj4YJAj
oP9wkwLPs67t6fHHdlBClv1vsOKJmCiOju/2TpXWg6wPhxmat0ee4Q96OdUVGxlP
R4n1Q4C7tYJER4yjQSiiDnI2C0DtmZyYLjCKnFnVfOYN89Vb1j3xtfn2w6a9JUFJ
gWUrPkJ9ZTRL4gao7rzMqFP9C+/ACjv9SSPYWM0e2OTqdh+9SBtZ9cPrxqVBR9pt
912LBtms38SmC6PW1p/goEOxny1LFAKOnEX94Dsb6InJZvFAbaAxV4pGlTXtIh5u
EWx/nrgDAyu/oZIkBSm7VYy0f8oX3668yotBt57uGrDE/e1GCrGIu9dT02l82SYh
k0gX+IH4XV24DXSfHeJSA6vW/EKCs8UQpAljTTt60+GGemdERNkd4g3aCPCcEcrA
qhsLMcztDMHtx7rsUB4M22Y2NpT+Oex536V11tUvZyQMm3b2+kgojMLWnXYUuTLy
5R4+1RmlrU0tSDoVEwD9CRUGvw43kldZ1WV+x3az2vu9jfI7ic8sI/2h2e+LrpXF
A9rGWUHQAH4S0GOExFpdkezDJudadEaPxTEI2z8jGrja/vF0/omfq87STgTthOBf
e5OiKSMTGGwhQtTRZlFl6bHxBXm+IrPP0/w2cOl4WBmFRLxPnrXeXXRvWamoxhC4
/z92w49aTlk+fGh5ARXVAgNI6PC5OVgb+PzOOU25/u7TTHsFt8EMiAWGJxj3uWEV
kQ0+VU/Crr5Nx8OGkisBMraSrwO2Fg9zJv5eJJs1DLk5u88TvYi/HSoNobUKNM3Y
5NwiK73HWYy4pgHcK7OQkVUfqEanghmrQPki/VtmFH5uCJjq02fE1rVv/gQN08pk
IcNzX56iTYXbfGhrb6zrki7G6HPZBQIzmNZQfCvTDkfbzLpdO0ixFI01wugrObSV
Pk7eVDX7IphqgRiSGlEQlxDnZTIb5kfhi8qfcOZ0ttNuTqJQmFlr8t+uTG3eanet
2j6WYKUnLdABvyTC18wrizKvVVYA0d2y2EfOgGIhzbhNhNapAaA/JSP52tiVfpjN
4ETDT9OeS2sLi1xCH4GO6014C5M5bfEhzGsVg+tgw6+6/Pasxy18Vi1T+56jPyIK
hS9Bd0XuHMPhIiprMN7BKbyZwhpJeVPPWDzPHrAjmAcAu+DsamsHH3K23LCku5dC
39TyN9lG8UCYEqOsY6E/vomFizzc3Yh3I808Baiaaqeg6W6401jYkInoIuWeH7sp
ZKHgPwEIN+tqu3sePhZFHbYsvABPQCHVyL3bq6ftjHPmkWVIuBvFbjVDdXm26AWp
j22x4DrA42DKMhmyOmQiovqtbLC82jWFSO1SMMSONLAYANe2J70YwdS/NtGYnxLc
RbLg/xbxLm6cDbbNtBaxMslPgw9gQlKsFwZ0ljRkEFbogCxGv07+zqIupADZL65H
kgYOdy1yVYMyXJ5CEADUo6OEeKLyVfzumR9WEsLVZD+9V9GsSOVtbognjvzIyQgK
73Skme3nHafengHriFov90NMz9irg2/gP+tYspahHs9u10jGCwjQLzcyRpQcziqB
J1u+yRZKV54bEa2HHsAPCDK0IXTfFcvOn+lrDSLx3W0BGqbziidgPnvlRK4ZumX2
4Pbv1Nv6GLAc9L2TcwiAqB119i5Rh1Dp3SVZeGW2O4WYdiprxIYH/VeniZ+r/3/F
CF52D0LhSW2+6zJQyI/LPr8n6omi+TQMxEnxImxqkL0xQP7/B46PibNdVmun9SoH
s9r7hlwi7I3pxuKaPk8btSaEPiP4RoDD7djbxwNtD6sxVg2pQPNR6+jMUZI2KVqR
bjuznB6QLjCo1wL+dkZ0g9c/M+XZhMZ6dUgdUogfK8XkPzugyCLoNNLnILvcMJeS
1BbPK3xIMAeATrTAgZGpqn1kDwGA5VY3BCLj+CCYomLkI63StgbALxTtF0lDO7Zq
aEX0jvEWA4gd/4vlL4kGiwEOnDj6IL57E/rMkMqN99XhwQ1CS1wXnQ8jcn1Wf3bo
TRkDidWPrfepf82scYWsD9m0a55pmmitX4deyrhAaJ1oTSJiEFcpTz2m2c3hEiSD
phniHlC6HJpBKPFAo5SJuVcvmZt6xfRPw3ve8balTx4FfpfnyTxhhHLxBVYlPpbb
O+4kYcRCbz/Jlfie4N/DEh1IvV0crXQVoDGVmwsV+aZ+EF8VGF8hUUoIpdcj2rd2
sv9iNmBkQSqXmo5RSWK0gDKEYATPTynzTSqoVA2+qZbD9mH4y4HNfWER+l+OSD83
OWKYOQJCKStfJv2rZ/bhZhc8lMwwwRVluVsFkW6qI9Av40p9oE6oowWEtHaQe5ag
Z8UHBcLHi3ZBIssc76HshuLR3aTTf/Mp55PmnX284EsFEnwonOART3moRG7rbo0u
X2oElj64IKtDS/ndcIbsYKWbaw/EDnc9HWAf+s5OrZMCCQjEMzK8ai9zWGaeMsHu
ciEgaTx+BvYsZc2/1DpGaoMvgMgjerMjhy5cr7IH3S6PLruQsf2EYsHOvS0n27+F
/0D8nkXe2404Mqml0Kn4gfghboBGRAR2s7mi/KGx4cOApxyaquhTG/C2+/zBANLM
4tk//GaNFrMSaKDn6OATaJK6URbXYrY5vNtZQHq+P4LETOU6ujYLL/fVDeJp7euI
6qjAs8i7cfugsACAzQOmHoaiceSQ3AMPn/J0TGurqaWu0xdTjVQli0XGq2oiy8q4
tVgY/GowwuKvkq1yT77lRQGhTZetSurXwJaQCHCl0BnSpn29vRQ+ZXMwrabBHMjH
Y2ferABCOCNGvGmW5IEKT212hWvAxmcFyW8uqL13Y8XDO6jE6fKdbUqTZr83IeGt
P1DgD92z7MYy7E0HNnohx4k88TJlsHd8Fs1apFpS4c11HQV93usrThjxvwHxR2Qu
V3ambfd0Waj0pzu979X+vSHzdZhRaSkdMha1K1g9WQtAP0Ko/q9bWHC9jUT1mjKi
A5rdQIEZzDNNTwsTLJp9sSXdIdaNMefp8EAeLZvAD0IpecFEnxfd9K86xHtdO3lS
WGN38gC4lAWNDa99tZ3BreTUiI0g4jf7/Mr3TdYyDObfoO85p4wBQIozIPNI1X23
U9RxX330i1oaz9izkasOWvbxC7JcYziNSW3+KfmWesmNSevbow3AS1crKvwxwYmt
DbUBxDUGQfvVL5LsBDmf7uPlV9cQzLlYqTBjM316VrOKlPT7dVH0ZSzv+tglUqob
QRCdXGeENni6xdzqwtIdTR9O9j8zRgJf+7TN7ODAboGyXzLSBS+5E4F4oNOWk/bY
z04I5ZdpYIe7udqwjb6lb7lsa23N90D02eyXUoN9Q+DKMkhqozElpsy+56xHtw2d
+ukRU8XW24cGsNFSqKzDpICo4A0JwONjZKvMgciYwKqq5yRYT/IfA+g3ZyY+ncZ6
kTBK3vFWzwD5X9x5OdXb4tAfPyrzF/adPEy/aFtiS4h4XJVvfDY62FkXPy+pavIi
DVnUpJP0VIgbOL0kTnjfzQAxdWJ9sbYT2YSQC5nbbhO4F5gLsTK5wBF1ErBPLBfl
11peHUDWedUbe2lXvo1+MYKQUynO46XMCaPKC0vdHvxyl2t+q9zPBpWXr3gm1Qb1
dmCv0yEebBzBTA/iPbMEByA2ebmYSIrgpgIUKjuaXFK1tAIfz0RdC7F5rmGKv6ew
SYgs26Glsn51zPQ2OoBZ+UIvVz3ypBBfFRdiKACfXcvuqNsmEv/eqczPitxOl1pO
Er5QD0S1E0cnbAkSgXOYLC9KfBkhMWl2Vn9Lb2WpdNjW+/TXPtEAtLR/PYtPhUCV
JqRmMkqQHm1QR7rrWil3SPsC4jLMGCs/+2d9CiYMbz3q9z0dTbK9963UZNU3FN2o
pkH7rVNwFkeONpS21jNP5KwE89LQB8XNQS78+al5Zx4gkU9Sd5pKlkiPPapEbKeZ
gGemAsgpwEaYppo6q9YrKcyUb7dOhcNs2noQQ0tkrSCWijMM3mjJxFV9f5XchWxy
qB9eDxPtwnZjw8f49niBxmHxSOiVZqc8lsDfaotZZMpNjTnY1OjLlLxB4ETLPhEW
Zsn1Z6wrB1XPail9icPjoXyHoUrqG0VRCI7A/+5L8J8tMQ7r0XL/+yOFRo5vk7eg
srW9bXWpXH4lNjuBWe7YzQTphasJwgijpm2lbM9laGvZ0qv/ZfrPVAITCBqSdu5h
PCYmL+aAiy9XNtC8IGXI0wWx2m+3bhv0c4FMRVo/mbMvepogAqaXEXDPVzW9tc6R
xp23rgTeRK+f32ozkyA3PGNOXTUVFwCZtw6MbXTY9R7OLi5naObBxd4kRA1LJQ9m
ixOhQbYhHgP84KFF98Um8IixNXS3qcYo+lkR7sjnb9g7Hj1zZSuRdETApOOBLlal
Yl1VlCSCJebcXpg5N0ogKnxz7VN2gSpB2tFSj/sxZbZ6bKORP4E5q53EuXtTdfUo
MLeRem53+pKHT68hrBXH23jJm0JTwG6V/NmK2QRdLwn1k51Yy2EN6ZZoHUY2Hskf
SXEHXd2hoZZdtVa+Up1vDnf77Fqo8NcLWH090K574lzwD5RA7DMNgwRT4wFBxlVo
8GfpPJK2gYciT8H8DF3hP5KWNNzeZ83SJxgQGdBiQ7nfrB7EtOXQy77bmpGhUU2v
6iXTgHX9buF/zRX+9eT5K/RcpI0tZE2IXt2Vc3TfIxH0cG+/24VTZdiIfO8pnenq
FCCSu7ox6d4N4oR0lpHmje/MpHFFsEw9cnezsKu0Nd5tHcdaHEwJJURq1eAmNmJh
stjJAeCc3QWmh6Bp9sYB0mrwWxdXmqx61xKO628zgNvd+QyJQnxJ64wRDO7pqz25
sfxtu0ut//g8IX2ha3/E5E8tzwnuxMkksFp7/dg8DdgXLEfHzBj1rcAQ/9lScTaf
7Qac7ZPSLtaHfISeQPsOxd9AifwxatZXyY5jr6jy+yv2EQvHutfSsEBUSi8TITK0
3DsFJkOBk+rJY74zJ3ApJQ9hzCiPQKulVDBtNQN1nmBPDWa2olrUJ8nEmEmDEJ1D
JjhwoNqH2w+4bDck/QMCqbu8X1twquqYyYI8XPuuPDPQNDAvAQmYMho1Ut5n9OMM
Ey9TW3xHNJJa2q8fNxHEZrrgV8Z0XTnG9nPKQ9DrvowdEX3qCPtaE84wRAFAK5x0
PGj4jzi5gCpdvCFw3xAc+8vghHB/nmTlp66s4/eCfW6ES6Sd9DOcBBhlqHY79JkY
Ot2htU6SCZTITsZ3XJZ7PzMElvKN1nBNd75rvg6Q0iE5+fug80UrOGPuZGfe9ajq
JGp5FXMm4pcWeKvBhM6ADzm+0a1WGnjsrrYE6zqJyV5C/okuDFZBK2uNpWsbPFzh
6KZfzzdog8BRwXqn3Ij6wf3Os1Z/i5NoNrC3HY8wL3g4+EEzDxn0U+3HxQDpxU7H
fNwSg/oxg1iwi80aEM2JNOAn2pbFDOi8hBMdAThBfHtf63GaU1AXqFld0GiO8Vjm
GzuDrnim0xQ87Q2EIoeCCfrCtKkho5invIwQw4M4VMLV8p/5j0E5t8OD/cVr8wQY
2gXS+JZWL6Ch4eFXMSPu5hd5iEWiU6sNLftj5NXGX8Jvr7Kgn/Q5XbQkOhfcRsLu
wwAJzEQ507hmsBtC0XalZk8usQos/GAFytqAkUMffftGVlrw/mTVmvf96VIN6aAc
kGU/YBkGW3pbW23u1AMmQPdG1mjQEvEDxzpe3LXrF+sdsHoiMvgv8XDPA51lalPd
e2aF9mPiLpsQQCkQv3sK8v0ZN1FaPWJBepO3BbyjbFnKqW2DY7B2QZ8khWgEeBte
UHcDg4tTTyRi3aGH/8udv9eC96NrscjmqRxa94cvN4E+c3sdVkl01jkQKUcctbxt
echnQN4CzM2aPXznjzeKhg+vnT5XMdixK7PbaqUx2eMY0soFNT9UqWq48vQGCJS9
U/9llKke+7Rv/3SSSALyFItaj0fxkVVwlI/3mWzAkkXuYQ0P+BQAMYKRjGBtESS6
LB9T5VhMcValphUbtIcCmT3ivQABVQXNGB5WZ6RjmDrBAyFal6Ijrg+9DIK2qzi8
dQhazASK01xL3yI82X03KjkWNnprlNkkIik60xft8N3nu9ZZSuwMGsoBnxixPfYo
OCPtPkr5EtqNSDaCiKlegY3O4D9LYTBYw8A28RoAhuKqrK2fVhuzv/94KNcFDd/X
E/Lb2P54Fjvf+cUECTTM3XpjKuv2xXcjLa0qeAOf3ppxJTOVsa1TzBt3+akaHwxl
AWtlOCCIgdzMe27NT7KrzqSH0cHK+zdQmNqjb+dsLhQi+6FXBoqcpJp0Y1iNtIEt
k7WeC23m1aQIrAbTuHe59nhfUv5otZZ3qKdMiwbrwSCrLbMDFLD6Od4hPjM73jgz
AbrHbYA76539vRKTaaz3PaOzZsrkEt3BNS+QSxQtNiObRqOD83Bqkv3sm9JMUzO6
aW6T2IY1yi09AfZ3tCViPWtOIcD0kN6eawROgKoKxD5P3qkarnqeXWq9+Q3vAXnq
77XIz+qF8u22QlIKfA0/AF5ZMTkluS2yNvKsQnZRTDhja6Ous6oPU4FpI6KBv75R
ABtMUpArF10KUDavgRnkpmgEkp9d+nTd8WlTUXXLGPQTvKbkP4si2S3hMiIRMmm4
150Qe0YTxxFbWO4/SdIAdT8k+k2DcDhcwqk0vILSX18oQlRRkkpGookBf8cs83Xn
vs0NApweKTAXOfZ7GgpiwAMtfO75JqcwFilxyt1ylru9IHTjVmM9tR/gXRNeUO6w
ymSCTnx4il6FDSeOw1LHYvxyWMlPftDFiuVKxJprUKtxJAsZb+LxpgCb8Oop9WR9
ZK4vw8fLmT1AG59Pl4DNUSORvfTHJPi8mLIGO268lE3TNJupfPNX8Bcf08LiBlp6
leI895C1D6oZHtg9fFaWarn/54AILxUcUy0FDx7y4CqwVB+1VcgoJNuNtwx7rImF
GY4w0ZJEYEnJbSh4ujuEV+Lmrze7FKd3mPxKSd6RswAlfNmXYueXoD2kdsens3rv
RpOpNsEpJ/EkBcGNa3Fo8D/hMK2EkbY6TDxYrgOJ70E7aFRZWxwjxvoyPaeeVDli
JWIf8Envg7imhaVi3nT/+O/AzlFYUG/V1X5T+zovYTmVXUDYmt7ocqH801FuIhA4
qZ4QGqR0WJh0aAS8MVaX8ZZvA5O0FqCUkfMLKgeEq8SuaOMl4uunhpqC6R0TLLah
1S0i0MS7TZpLo6eGq7oHJDE8BUkEEvWWWXzQNYU6owOc8WcMYbX4XBdCpY4/3Fsv
1dpDUWvfFaIsQ+El2yQmLvij5x2V8gSk07r4pgqSnE27RmjozW2W//OJsZFoaU5d
eRrLMdmQoZVHD+1rslpfpjU7nH07WIz5w7FPABaEyU6uo9bPcGsSykgcU13itnyz
JbB8q42/zLbjvEI/Aox4e1grCOFj8LERXqaYwIf2+VRbxYXWvOSp7wU421EKKD8b
g4bOuo51PpqcrZw+wsOxtn1TRf3SkW0wTorW5bNeU5QP114SWzeAigCu4kKoJ7Qt
Nevmn4qc2pzs5VxzBLB+D0ySGCx/ZeFsL9Bw56KfVB0W5GjEdiKn7yACLkZKieQR
UJb836ERtFiKMnJw48/1RddgIXtGVEKGU7DUcCW9Ii0OnCSITG5NsFJXXeGmllSh
cvRO1S5DVtkbdVBXQtpkWrH7Ijx2ZAILh5ZKs9IuAmuAqBDzJFftp9h1FZeqcKT3
s/a9mhB5igDWYqNtLe9rA4xZ5wbZRE/aILT7KU2Zip+Cr9ymNzNeHCZhxF96CSXe
sDcTg/sFD773P7DXiFefp9cNCjhqrSPKlJWWdYIDUlqas4MHuf9Gx3QBBSdGY9ml
j1iYTNIfyC3O5stL/MEpa/xUqAhWg4JYytnhQoVaPvMDVVP4ybqWHpGPqanSurTZ
GDl7IN3hjuCOxbBLafIpTAW2qXFNvf844wZI8ZfllNACLoOk7DhuHh6EcEmuccqk
QlMceWEn2GECJWERvcazMgEsN0ztuKENbPKM0y+X8YUABEb5/zBZIywCgtnnPIkR
GKQQ3pjX8A7XJxJL+LLy4b++kgT+wE1/1yC4nM+u5sFGg9UfX3BgHh5mc/6rEfiO
/dsLkCUTA7jAXEjEbhA8zZGor5OMeetJ1bpAYEqq1aZAGpBdzt1zye9yj+svYJbX
TGbgChtbdUzYlFedIiLLwqZkBGciqgMA/mrA6tbFclSITqHM7SPPrlvb3UskjIGb
8rrsBo7CAWnaWqEZJy4np2KAMyVs9o3KmetZUTciPb8GOCSIIEpPftNlRkYeN1/0
xneW+3hhaU6/zRy22b0XdyqibVzscOjJ2+gmbmYK/cyk8Go2tpmZ3hhtet82yDx3
XnoRxu6W1KnMf0/afVLNhMRYXvF4IbcI4A//ZgfsVqBu+O9prj2CKdnEpNnPtSz0
PXqE5pmJrznfr7xWr94TAWzzRZuSToj47OnQVP8qo0nqTslr1H3h5UKaCo9SHpn8
Tk2ENy5oN4PJU+mRg4kuLfePufU0GREdU9fd2SQEgWeD5YnOjyzfYvDXgcz3k5Vs
WrGmFV8o5SArhCbZl84E2cSVMCKTTE9rsTf7g6lsQX5HzqYxEykLZ33Btc1PQQ3Z
a7UyP5NkA0SmTMYOt7MysDugcDNQd5xf4a5SKs/mDbXquHcwJ5lVrH+0oy1bs22d
BV+24JtqQ6ctv2QR4Kf/UQ5qyITZL6IGQ3m6IY8DMM71cIbf+Hgr7obnGjWML1+i
x/GsVCaQY5G7lOZc/leJeU+cKCO2iSD/H2aKHmkvAa7agcXZMgim7Rri1Jowt1s8
AJGVxd7cdcEkIs8UtCA6VCIoTkLuvPYihbxqA450cxm3Jlt/0x5E2lSb0aZ5U8ZU
yqdXsq7BGwrILuo2yHXCOddHl1a78Lu+4Pg236viEDQzJW+iNTx+K7UDsF7S2XT8
xnRPut1K7JRPQ5TSwl/OnTvJEaYltLbE3VA9hUIkJvbesAiXoqAqEz2gtg1qPNMv
cZq8Lk7Td+1DBch9mTna3eYpDn4uvNlpF3iPUkHhgTPI8GJbHD8KGbL2DGiqiWTq
oue8W5h+vg9BuAj64uS6BCGjuFc01d1F3tcN51bDbGOupQrMBwqoUOhkWii2ThNc
8VR83CBe5J30Geq5ji7ST6cBFe42CXm+1BLazBOSX/kRkvLFOZZ8ZyoT9byGxpw0
AskXxHqDZwIDYbWyUBHE+/JVDSLZiWSiA8yXVMIvUAnYy+a2Z+LKhEBsBorNkM/z
/mKpmCdq2mC1RWXGHzklOaA4vAodRfbPl+rpUUnRHJAF3BYZSlRiXjGVmbPIIMKa
Fg7omJU15vpYFZhKff0a/3fCehmQGpJGyvzyCgVssjB0QOIzUMDofUcuPgId2gY9
fv9pXJRXGjJfwj0KsagTbx8sB4WozcwpD28nS8MLHtiBhnWD3alPyeIi9nS1Hagh
TozaaL8YEu6ym18oLG0ybEegEj7WsLaWUTKCZT6f6TlvHIzd0t1lqCoCHmosHFXj
IpPzmYs7dLWyVxP7JJ/LJ0Ydz+T+n1rlwNygWojSPlUT/KjbDgdGHEAratHRHH95
/vGfcqLZVAi4DxQsDXfcT+WYmDjtfl48fRzLhrdFu0kVxGlwnLh0lpZxRqsJgoAZ
lzZLCqITpoKR6ypOLVjq9Z+Tls/5fsNhDUfDiWT8uF+UNt0e32+6rEUCrk/0HYM9
TF5P6JV8FSKfhqungCBWoQhFhu7evrSNCHymB4b0pCpekfJf5tKcWsRRDZssTlfM
zVB8vrEoEqtZB0ip1woqRJIMYcW6kSrjJ0OEF5YpW5eBCbQlStZOaR1hBccDIyGR
T/SbgfuMdIzRTNKOTQoCnIIjaRWUZEvQ/4whISdAMHiX6xxras8Pm/3v4eRWlvme
eXCkNQmBqj4l7WzomvUQflXpzlIFqCefWMUYLNOK9NdJzpACUzmBkcOPCRMgZJjc
TiKQfRB725PEtVH7zaxMI8Bvc/0qzx8JLIVwYqxDoRtyHNsZRLI5uw20IoLNzdYq
s2yMcyen35jXM4/vgggTUm4qRVhxKsmYNad84sbi/k7DtYGDt1RlbvDItYYK3pym
ZGWE2/iUcyePAewmznPfbjdmIZNIagHT8BWN5srZFII40WLShQ8HvXJSEXPINVJD
t5oMa+bJJyJerf9FRWXVJdYzLzVQbgplCEyf+oIoa8tA3wRq6tO41jYeYe09jmZ+
E/egfrEdQToDEbOk202VyVpJspsi1K11Rkvv2ztXnwz5z/e5nxI9lgniyyuYHySB
1Wl870YsBYABHSk7624VqEaZjSaageD1URD78SXtBafbHDcUbkIOuyjO+TAHk96C
W9j/gZ6T9N2+yPAFHE+nHYzyRCHtLxg8racurt1bD5gYMU4NtaqqrnFXiS9mmScp
ycQS3oSRlAFDRgSWKZhBs5ihLPmCkb4X/lkMNzwvpuzQ2YjbxrQAyyrhPYnQvCP8
W7RRTP+0roa9tLh28QoVl9oIVad/4bMtZh3tqos6ooVfQz4o9BP3BqU/KuHT39DK
CFhAGTH/S+0i36Tlb1ll6wEjQz4aZGfRXL9VAz9+q49Zv8978oBzBlWlxxeFRyUf
iGd85WTD/I/U/WHy6e/EEUn2L4SFbUtUHMOWGEZMlm8fEQp9kTo0YIzJh7wIDDpr
ZKckdDqH7Vjx7XRBw4/daXnztRtApMR8HQ7/mpM6zF67a0ODg41bPsu8/T8JWG05
155FV+MVp+ti3Hskhhnyev7uaFDqV2UIgECIPZ/68ZXyJJO9B5KqNWTsZVSyoZ8F
Roujs3gE6/nanAo55H11wjvyD6LTA8sBGE3QFFHQ3QbCEZr7u4Im6vjLvimCYnEt
oNUCzs05z/h+S9rhD33e1ILOlpBJnXCeJpn8UMf1F1yiX2N6nBP9QQCwDVjJ1VJd
4yS2BVxZT5UPDZcZCI1su21kg7jaSsEI65Odv7qMYz4UPVghk0fpBnWbVsSBhgKu
MQ2fMxrPcTnBnvMWcjBOUw/B4puFpUIZ+OdeRul47TQU+DkmujxlXTQJFbJLTapu
NQQrBzxhTt8nxDAf1dEUP6dzPq8km1HStuRqIdMrrHx/EG9gcvemlhDGP4+jA0+g
WE1Jxt8KQOum01lSzeivqCv3MbUe/fLnE0/MOup9l5vVxgPYTSnwGy6rrWg8suRI
TZ4Y8Y75FzpSVkknb785SiIoRooQ3IdXSnTv3x9vXZ2Yzs+eDgxdN5kQ5eMB+8Sd
EO6/98T/Zy1/+7a3lA5Rtqn4BHpiV9BLkKIu2Au54K2F9FXNZeb34+giekG4zcHi
JZPZoAIomg3dIgjoTNDAm7VRqWqzrbj9Icj8CYl5YUCEOTv87NfzrLkWlA3Zc/gH
Z0bLpRwXD8svnyRKIc/I1wHAe1622fz3i2s13Hom0bfqj8Mxq67ktXw8P+kkyjyS
XBvnYQ0Pkts04zjk7PA1aQ0CnYCqyI5Uuh1rS4ao0JdwacvEVa12qgxO9+8afFUV
qlLQzlZRPyl5ZWtWutvKS614orM+OjxNnncFi6lLQnDLtYHq+x4qn7o2l4AiUpbk
cnYS2qkswQ3eURu0Ls7nWr+GKEh/fC2FfdGtxHwLBC2Hj5J1Aj6H1FjRW9ZiIGzF
CjSyhEB/FDiWo/wVnqWF+79Yk0T6SuLvH0+J/i3He7H7WuHoetmEEhS0BbygbaQl
lQggpZVsJG4/dZJaphzaDoz8McC/uenI27gTb76P1sa+Tdh55xskvAAWExIhQlNW
ijF2VU7BQHCkeTIRAc6wEXdyRuqUMYTyLmNgB4Ou1iMjbDT3RXw7WNO4r5i4Ppiu
nPDBmyw998WHs7oNIYMl2esAL7gfbsBsIblC4rTt96ja3A0PPQ3lmP3AEwU4nFah
O2Oj20TNbcVkO1j+Rl88+BPeb7hYbzdn0z3/c9feAF1PxzZiFAs02o/le9qXESvX
sxRr4wr2o8j6rQJAwg1rYZJY5ghuYPd3QZedEqZI3tMQoB4BjyO0r/mODvstqZHH
CioHTgr/nwp1imXoAU98LRTgET6TXlDRGs3WmNoURNAexGQGdmhfD/ilwIzIlnhE
Yu1b3S3Yf5Bo5To9MSGaWHqZL9+MpRMtEF/2Th054vceY55RRVYwYrhSmaECEsIq
KJnfkqaYCK2GX7nhrEGMIf8ac4yqN72sVhe5PLPrwGiCOE6sT+LfdVb7HOG+04yO
fitOyhcE1y9Y8xRwkcYejFMjctECpcgLzvsdcDWDTuAciiVYSbaQg26nJMCMqtD/
hXLNwW+jw9soJNsfLW8D1U1lHmWuQHyjnTNEKLq243psGQjudeNqiWlkeulg+TRB
sE6Eo7ZpdblTKuH0oRQalR7Ex6sbdzIaRojmez6wMzFl3+ZJaJhalHeGpLHxQTGf
0RWv96HoxzMFWcPbSTr2QIMDC21O57bk1NltndA2TZxQWTlYnOF545O2Q9+ii/hS
BmzP8jfP1tF7ZdN1JFgJnilji9RQ/rDDjpQ6MKtLQfLuiH6IYjrSK9iIEK1q9HIE
+AHXALN2mEntXKcfC9wiORganDLne9UktUbA8HjVa4MTY+HumwdbOLjZJqFqTbBX
uZaj7t0ZS8zK5pJn+ZsiwwCiHKsjfipMl62WiZ/yG/jhcwnuM+/0M9IfXWAtdnhV
UmkJWSb8ICqc74XFoVBqpGvFWJ6LmTj4O7qGp/oxa9bmlwb+CaNhu+hEHRo8w14H
/03FzFSsZOsjVeGQqkkqI3J7PsKaVnQU/7V0r8j4ObXgJZduZsGliVV2+ZMG6k5y
B45fw3QpGBf5aVALES6MlaMHne+SeoRGIYkSlDEjcB9iiHIl1cP3rVpcZFwKuOe4
h1+o/L3uk2VFDxDgRV1bzhYTTz8TCONPiuiiNxmKvyvbkcL6ES02xTC27SIHbVcH
D7k/UAz+TsYSW3Tx2pbyXHrxvtW+dPRbD7KwEWkDgAGlAbdxLtO7ShmmHdH39yty
4+PWoaO74JkJjOpIgKaSq0Yy6jDwhbpiZUmNW42shIuHLmGAOkVqHaqJQKEELmLW
r0XGLfHiuEhQ/CFUsoy1iN+3z1q02fHg1u3cztTPUjTzJbF2Pgfhz3KeDh6cY+L9
G4o0jNVxb+0klIauPwVe64qeW/ILgCD0hBYRDF3ENq7DPcPTh5bX7nzjsm48GmUe
M9BVbUPgSnwdfS/ak7aKwUzlrybkgyvOqXXu6J1NSk632zzyHnUe00UPER0siFO7
OIkp5TOoYWYVzEA0xPIYuIAVaoRxOzDnsJak0lz9ka/59wvy24F+RQflaJ3+rKrF
Afq8HgupYabc2WQuIUgCHHi7ss8bio9v4wSkWgQa8VqnVoroahNbB5oixYtkaWYF
kUGXK+kr/TyVykY0tHDiKyPQx3tPvwUhVG9qlhhnElqD48qLym5qLXAmavIVhdFw
3GTJNYL83wp62Y2lQZT+5rAT2NI/kL9kih2miPNwOGUIIgGZyXgdN/iS2fXBv2uo
8hmP0LAIe93PW24/4g36a/OOqnoK38JaiLHq6gtcaCSEA31z0j7X7IlpYGYeectG
7mU1BUqYARPkqTKhetVFUEC9u2tOL6Q4O48OnXACrUzwFPPKOQ4ITx9HGSOj0stf
mgiJgsckFr+aKPrPDQ+cWwJoU91EfKbiNmdYr0GidJnUjB4/T1hRnAzlO0GMG6HZ
fyUoEx5KB4VShw39AGioOm4s5Agi7yUubgmXm3HX3qxPq7W6aHaP/k890CtJ9qnW
AsR4hMZ8WmIHNq+83JSN+/mrOofX8uDH6ImcF+/hT6SvaWxyAaVMx3fP2gpMzc7g
P3fqbd/zRXxEYOHys7R5GzZZb5xF1Drv85HUSEinCS46zqqi/Siy48ehbURUsMLr
cLGdv9h0KVs8f86khyLrne0Kda5oIcI5XJF4/wbaVU2xzg8gUCwAg9ANIdrCGQXT
02mGfYmLV1jDWTaOruQ/wNqGGLFS7Uw1uWC+Us0N1UvtQ6GcMNzihtyvFyhdsrrT
9ouKQ7aVoAeHML6F45UcEACnw3nbpmo+HdOVKUEDpnjjCubvyKjVDomGJCUrl4VE
CIhOFuTzwsz9e9vvdxgGAabf6iLJzS3p9pwl72ZRm12COPRKeL9obGFjAaTBgbn5
CfN2lHCjVmjPaOq1QjG6fZ+BFAxmw5Bb9+IEU68IN0md1gaxUNHMAbmeuuYz8DSe
6hPMcT4kzU9PIglTWEPg2jiL9rsxBmJXxeUDswBkUOqiq5GzyuRmNgAW/OL64lA7
9b3H3EyU9NuQ7bPMFmc+5sFq/tBfhiMup63/JOx3jjqCeFX3+Kc6gbEmQ3Vn9tyG
awOtRk8ALXhQojo/meDpMjvF9Hh4jSY3+PHj+m9wRHTDlHXvno4+gT4TBxzkjuuY
UqTGjewkmdNIQVNnZj6alpLg4FdI4Xdt/nFYqNyBuxbjH4KQWdG8LL62l1qjHhDT
IvzmvtN+cx/aX62VEa8a2T64YD2+B/VgzhVu8BP7auj74AnMKukNFJU8LhYm0oSw
VF4wkltaMULIrD+U2PWUlu4bmlxJm+Uo4SEklLMpy/wNgymlAfJ8gH/ReBYV6RWg
O9JCAwsol9ZWHHcv2YQ2Kuo53YqMg5KFr1BSgodWM+8blHCl1w8VdzzAf3pe8NXZ
vEGZp0FQljEVIia7U0i0121/SWT29Lq+YRJjSi68YNsBIGIcyI6QG/MFOUUKD3Rj
Z4dMQgtWEdNzkKhrZQP9vsHNPiodlrRUWItJdb4pkP/NZNYWhrJQ1IjzYsn8npwS
EcR7QErTQOgczHljyVlwbaBlcbnnZItcsZS7vvx8KM3ucHuPhRef6YoR6m1vkH6o
skHR9F2OeLwGYUl+r11lVjuOLLd/NsFbumT63FR3CIAV31kl3anVai6HEKaba4Eh
v29KvRo/9u99ybYRCyAG1aJGqQD1hoKCXPcTgB0BBgWHpCPAgANulzE54JcqMkay
mrdC18wsDcgY1TnpxfMqWmI00kjcfkQChyMN9+wpDyVRCxgCFzkrOFvUXAcwSwXQ
8RzbeGLvVLQR7COy7GTQOEtx7qxdrMBOYa24gGtOT2ETLjzRl/q+a/GPM8kOF5ja
Va5T9/MyR+Bb/vpb1/gm5FYWA+NyqWuhyw8ka6Q+pr0kLqn8YOUVCejy6Avx/jFr
3G8U3mdOTEXs/Y0Z32hYRDtk6NhLwrutW3NWQevDJAlTaGi6U1T8NXe9WOcBe9fD
Ufbhx/ljVBNJEshGenUucG8BPvshTpK4nfce2DeXkndkfDgjVt0y1C3XndP8VOO0
qMz9+vHEQofGZ7l3aZi8BaO3Rg7FtUrqBEb05gSbm9AfW8ohG+AqZOPJf42Zb+Wr
Vb/gQWUsDZxQsIZCkJ/1MQqyIlSUAwlZj6NByVklX0pbO4TMMcMAJDa+NQpsYhxG
J4GMdqpJSilwnbqg4d+kJERwIOr/gJnve0v2lC8+qusG0ZhsuWubvUzdaKJXjRWZ
oMoRFdoU6aoGzsuV/oHfpxcxB0C3ZVVbZt1h6zSZswQnJ6tG+xJJ05/wShhSjCmH
ey5OpMfgsfANFv1eUBbCv0u9WVHfPMwURWehYRs02SvBe1/TyRGdfknoLnv1QEiH
DarqsMB4q7aJtP1EzpCevdPMZMlCYu2xN94pW3RAJmrHIneGqVKb0GhdHL8kvi/d
E7LvVdYSvdXcI5SBLARFVajqyP8UeJ04OZLNMYl8QphiPiXVTLNqoXYPBM3vqHC0
smDV4GTbTFMl0oQtjTvSWF0ZezHFL022tEAZ+EzckEa0DiPanIs805nmRud76yVN
JvX26J+x4VzP62uKI0HO6O87o66XZfaZ+VGEL70qqWaMSuK5SUmf6JDByslovO6u
cj2zpOzl8anwVPzRJ3NS/crD/0zoQEye0Gx5P0k2Op7dZ/31Su26waqD6xuZpZut
nG2OpTKHbqh2oqDmvUK3v49o5YhFkUmls2Jm/3raQhzb0QkC9N+G4n8D6jXHphdb
4j2O4vkzNu9C+MQ9xSws7nS5NrM38T9cUO0oYy57IlBLdgmakJti9e9hRJrQ7RHN
wc+VhPwLQOzQ3zdObOXeGZ4HaCNjMb0/zzfmkXAPPK4ceSdwD/4NHSkboueA4tDK
2kEUn5KqOA72ciGKEwRtlordd1rOD9Q3ftIBypYwmbAaO9yTwSOLL8vXWNLarkIe
uu122T3h8QYVdw3RNxuNNLL3dG/BiJ3oTfZjbeHfA3owTvLnJBVih8JAs+XoCHxB
/yUu9dD3Jx5/LetG77/pRk1HM+a8JTkmH9TsS4I73HaOObOXi5BdUj1Oljd5IsqZ
+yt4gZnZAOUiaIvP78VKn4yw+9Qw3FfVh+ZO75gcsfkTadOhAMGHYqSRW5gLd1th
hqmUg9UqNb/aU2P1TKo5xIiHjH+KqoryGZnDnsLRM1dnG51oRj8hP3Q9RwWgHZp+
Z/9t8H7xlHhoIssiNMAUzNpFlxDZS6YGS+ciH81sL9Qj76EoaxPy2NR10RieYTGf
ZguLSUR344hDrIJS0NnCM03UGE3JIasTEEZ+3CUkSUgNgMG6Zz07Qa0ZaBPCpHV1
zminRJ6mwcJkK9KpkvK8Mb652BT2vQL5pDaQeErOmeSNoOth5d1uYevVr7bDAyh5
hnfGfmTsxIOVK7oLppSkfw+Hg3IWZBmwS3ZWpig6bXmwcwKmC1BlncfZuiTbIZYX
IQxExVfYx4NOyLgmLNdo1GnK5UFoSvXduJcSz9lqU4ZvK/HKLJcAkHjjGUw10nze
149iF6NdT71ogvAbpNxFKvNxnr12HL77yjX3EoDa24Uh9z5+3uqi9y8lIo9idw9v
oJHjl5IxDNg7Mvj3kaBghNPy42KP51mONqA7nyILBfZWQHgj/y0BDUOOMqffk5o6
SOPcf7B67ZlHmsJF8JmwMGr97d8zY/D0HUWXDXMQK+EewcgLfLBDvc6eVNht7vkz
Dgx7XtBbMJfdLlhKnsWexZSsyBI7zPIE37CGZhnwNvWzXoXv9MNn6DqsB3rwZEXe
2OIsGczZKmako/VN5SGkLlr2/U20hoTwUZ+q7XAZuzrXklBq2DiuVfVIZo9UgSl5
ThCTVf0I0W/vIlIyMVWjNRInlhiWUei0IjVHNH8Vr1frWyj/+c13Wu1MqiunksVh
0pyTvm1GmQ/xUDoXrUrrJzs5NPAJUKYnreFSAcD7QxT3x+24WErH3cy8xAJVJocI
0Ra0OVmvbQkV9bStq5tpNqpM8m33suKvolVJCGp5kWMwmoTFduun+1VjExEbBGht
SxRL4o0iK5eNnU2nhtookRyYAFFvuWY/qOJ15rZMlQdfkqawWB8LmAHwqlqyJRFt
VoeTnLph9jZ2/5h7vWxn6UlOYUPyrGexdM33wvokY9QLdZ/gA8F1L9agMdNHlnRl
DXx4QDF6+64G30YizQ1WUUvXCySNLHGk+7MkeANZ50J1M0u6JZzCBHdEFgarRV3q
eyjwGgP0oCD4NUDgoexCmlOFISHFQI/aIkhdgcdE0EXgAPqGqmgmw2ADrYHwjrLz
MM+NeyvhSwFnTUDfaQ//7Obkg7zzI9tColfSaffHDRslG7DlNzr0ww5ZuSZ1BntN
J43lj6CvZJg/4YkXRdLHC6qGMHc17BWYPNOc7yithSXaNylSbrEqkl4o3lB8OJj1
K5S26IxFTntLQkSTUtZuDoQ0ElHWUrxe9o5NlugCHJn/IhCGIMBq6j8d1MHT71N1
1bZS3MujadwGtbcSHPrY7bVD6urmvYRjsj9Ix7B7vUVHemKd0c01rpkTRlDiBsBv
R16Ir0hmKDOaWRrlxms29lxexnkmAh9ERpk4EW3anoVUilXNu4Ct3uDlWw6PaRSA
tr2/HHyIUS7b2dT3VjtHmEeBdSxAqB9wqNxBVE26VvbegwS9q/WjoYDNTKOliMll
c8UF+ZTm5vXFxyjrNYKAYK106fleLPuu7fJZtvdp+gbFPGdhZ5s/5T3Kv+k0YhT2
MD9awh4l1/9yeiHTw69ansyTRziGbUlsW7H7D1s3Ck30zSqV+JGynNKHXC278dRE
NIH+3vjh8bojAiFLVzVkdVrr5M4Xxh741keDgoHuK2PzZD52XVYPdvHxYdj2y8BO
V9l9ueM4Jd6CxAPXoL8+bXWNE5/IoDVRk5pJCrkrc64klZNs0AKC63hqX2EpdZeu
mYLAT3XokEiKQKRGU81Ffxx6XUFUBLa81YEs+Z/f47kOfdDq6HF6hkN2LmhfiOvH
JdDknMVxbswlJXyI51BedkPl/NtIiGbHehOWnmcwAZO06r/YsVv9hjUJC2ExLVMP
wYnO5YYnzV37LvEBKeRSF3nxt64IlKHU308e5KB1s0tBKfj0YsauTFWJ27UeUzs0
AymA0OosvLXvhIjbm9X74qcd5B88wdNkzCCN9yi9Dk9JYwHRAAqgqqfC1/ctE8H/
xZ5w0U/pyMrBdOr60RfzlhCqLYnI/SRfqi6FS6rUgFbHM24LVGbYu1tjlB/wBpYn
Y1FfwhadJUF5KPZe+cPse95YREoIQwiyUsKh8oIrTWS+dsUq9+MgH8tokBX0sQ/A
+YzUsy+XgGQ039OmSv/UoCzsgW7JNBWxP9e221lFumeuDLVXUh1Ow3a6iKsr/BIS
6oi9EukCq+FjfiYVPfuAObePvVFrhpZmmEB6wUI63PfEi+A5aCQT9szbUvfDib6s
16L5h+0xy4dutBUG7vmCA5A6dneYAI1lKLR7SwZjtwD7GisWMC2vjjYl973pdB1n
YfUMpBIf5+D4N0oaiTH3KREZBJVsJJ6MVjgQ4Shjt79rUJn+hCrY+XAtGMZ2NLD/
Or/4wSq1D3kjWDIMy9Vyx6ChxjmBqV4+6TR+Gc1nr3ofsA1xwqb0TohxHnLtkI0B
oDVrkfwZHz8phlp2K3+ZJsn9q4xNjzeobQSimtMLradu2m9suNmBT+aIBzZp3rEJ
dCEzl1LUsgSTWEWhR0Ixurcfvrszo8cOKyWbZBD6Hf09jU1umljd+6I2gLmLQIQB
Mb0IP7aCtg2UFJmOJQk/e/K6GTq7jB3u0R5yq3RJZR41iH7gOnWAQZ/q1mx37nwd
1/tYXwJEvJic+31nGm/CujWvL5dd0tuFF2N445GiClEhRek8wcT5VoeTCLzY403V
goFCpkxldvmNkvBMGgIByRIso/k+5kRsgku3krnHYEARsmQD6OT7a2ZSfqJsRoVP
Q7SBU7smjMvesW2ZPuslndV7p5EFOYOWU4GfpO79T8bK1SwnzJgsXgrukUdZhdYC
9/0s4s1d8ji6kzw43p9xDV4ZBnFbqLwnARoEKN9Njb1lOF3roNw97xpV5t4rjohD
DOBQJRrsxvHkUeDfocHbryfRp/f2EjSMTLBc7oRvLSw1e1+2+L4hzcEHrZ3b/3lO
2teco/4VTKMLQVy3vv5XxTH7SX1ryzq6BxuJDuaUKd3LSI2hbfrZMplO3SHWU4Fh
x1m3ZzUEuZj/uQ0BAhdWVmQEwYS5F9Y07+FpRrWKqYGAvWKZ0oPUMLjIJ8vc4fm5
RknfP/N6/xh7uL/yZORywpbMz93ymxEegYrBWG41gRfZo04DtFCAfc9L+4FY2WTg
h1d582ozqg2E4PDI1GS/S4JpIjdJgL5Qk2dEmk6dLiTqjz/LGOGcdXQYDrF1oPha
JyINZ2ijZfGmbnu68M3UH9FHPECfJe5Tp1xU+3RP6vrlyPxDkW/xTzFJXrAasyUE
0M+1QLkevbqQ8bDOTFIFJr0dXoMfs9MgBg7NiuwVNETbu8aciB3C+Yd5xzGsbHqK
b9Y89PC1hiDd4/orlR7ClCOk9XiT07uXkS3hfQx+GoXni6+7cGqhSxp0mwJT8XFn
ufCj1IubtHWcU293K4qSx018t822d3Y0rwYil5QfR4DM0dvkwLrUIuGqUOWS/nHI
HIkVrZGUyb8/xjRshBNNogOr/pxnRGN25wTTuUi+l6Rd875Pe+yo2xbMbheuvasP
ZnetnZr9ermEzsMo4Q8GDo6KrIceN6R7TnEO4W33/xeLUops/qLXO7pNTHyf2nx6
ziVK2atUz3DH64l1WhFJVA8XkanQIA+bWQczCyw2vmeQYj5IGSuiFZyTBCKIrL4/
OG5fmgBBFKET95yEMe4oS6cWSS+IrzW1JSEwA92eypTgFFVMY3r/bsNiZIJcWqvr
C7PVQpTsuE/KvVquWXf/sDXNxZxKihpZkRs8+MQZf4mng7RD6Wz38jznPmhf92dR
QlVMPmrDE1VuJE7HIE8t5jdAwd71IMh0FDgG1tGwC3rpeQet5rFtb6JpWGRoPqy/
n+OoD45aMJPQnYmhPlU+bV3NWee55yzMsngZuFy5LI3idZk0YSgyaua5nAoWD4ys
YJ/nUTndppKCiWBeMqeve685uo1Zhwnld2ICAKji+zn7CJugEQynNpxDQGKAxiK9
vFMM3Ca0xBRs7eia3473QGBJqdGtw0YdG3v3gUr15Pp7JGVlLnUt9pP4HRSFP12H
5mC/PBpZ/NhiOTk/2c/wcHRXK7peP6q2ki1dZcVdDKahdGKGBiCkZvPH10swsGF5
JGB3tOj7xvJV7fntcW1y5B92ONiwpo+2ZeF90Ow59F60XW/zy2Whiei5uZjSgoa+
b5XvWTqhDAmzbZD2usM7uPL61ih66C+Tc/6ictCXsNI0KZOXOINNsoDBPK/xpnca
dQluxSdEccrlLYfSX6eQLCp7N3D4nx6e96HilAyjmTRanDzsLMDZlYIDNBAGIg+I
KkgE3mGm6iLx/rAx0tTcg0ONIwx1B1hwDDWiYtJb+zSQqQGXYF8a/pyLrx3dD9eH
0jlzRp6OQ6Jl2M7HxVTvsUCrcmrUUafYavtAxN2gK5kMAstviVZzP6pz1ff5/q8o
IAwjDZGxkX4estzt1aSWfwvnPP0joPLMwEQQLXtn4hdBHqLMlbEkNlGWFB8rWmFg
D5f2ucP2MOc+2c+lAoPgPe6HuhGXNkU9IjXh2LKqnBvGIzOdbI657WWc1GcQrUFM
rphy4l6gi72HABYhP9eHnSXBcUrqybjSfbRgAFmWU90b66Bnm60yzc0IAu/O5Bd0
Oro+6L/Qx35WxcMdoelfLBwvjqP74XTJr1xqA/zkiFSI6/vzAkVNSs5prcdaOfQO
0TiWTdjf8aHrjjD4+a8cEypad94dvnf3+fxIImukQcZLOPIq+pKZ5zalIxeMFt7d
4DbF1WRkdu3EfcrGgx9dmNiLjitlFZRyvoSYKpuDDO2dsogKheo6eLzQs0gUGHx6
MCtahIYXp6YGx4tUOX5Jw+XBPBxMpyHAStOGsQCqyClt3j3YNSrSJz6byYM0pc8R
qSYQ3m15r/jxXVv8Yjva2Z168gtODlA56p32t+e0RMpa8JB7cdxLrqBLG/TBqesh
jhalkYSp5s0LzWt+Ckz3ZktiZxu3Rt+vfWxpM3CaI7Zd8L79NvXmC/7XH7XKkmnx
G5ftJnqzVOatAyltfyo/S1xHdxk3gNdmV/Y0TlwgJnx/We2DBtMfakWPV/lRwpd0
SWQRN2NyD9ivSSz3iip5/wv8O3BxuLQr4aa4PCCO3+Tq8O8ufAOaMuQdyZgPxFAW
po0VpfWQjGLVvB4jYsgZGPpsoYcvJ5LXFb0Gy0RajPob0T8WE2zf6frNx5fDXzxm
LoIwONAPF2eLo+zL5ApFN54J+zu0XG0Z/OtjwS2JU6c2BJ69M9c77rkZFwfgcRda
5M+n2ClkR37O5Mmhe8WcsOl2KbL8voVyZmHJB2m9qppy3LKbgLEAWKGYyfhodCDe
xlH8ZvMkd1ayQUJLQdIX2quYdhT95uh/s70xIMATUXy99BgzkdCrvDA6WPRjk0H/
ZqXgpr1XMQekybMxEe6U13ySo1BjyblVBSJ6U4Y557FC1j8xLCcKLOX+gltXADaj
HqnUHcWwBIo6Yciy22soeFyhTaVZdUxjcr8WlZbgxAO3fKj86nLfAUY8iyTJj3SJ
x8hh4TtqqxfwIllrd+cE3tux5gidnP/BODbJs7LPvLieoYiqzIyawIAPjIycsdg4
7eke/W1ZgRsxGybUII+B7rse/GfhuCWiOhnvvjdqwzDWqxvAhN0MJAQUka+FLVB8
ImuvRZyPaenpA3m+cMsSJ0lnwq6pgi7XjqV5alnB4ykpnChvdUbzyYQZDL0cdR1J
sF4VoP9WN3bh9qyHBDMgyjVXG06wCctDBc2uBW3cI5Dd2Kj0SmENQPNc7H64MS5p
Ncm4J4FvNybDZe6JO+o8aih+LFtEeHv3fW/GPhrjJQbVDU+0YZ5q1dfJhphGCKF8
PoYvuB5vhqKj2n0ng+PjQhpOwnjVcUJTlQi6c0VB/+iNjcDx1j+QJ2y6jAba3fgv
Jh+dpgXs7M/je1Q8CA2se3wzLZi7aTCbRVvn0wtUONfN0wnLBBzf5U9pUlJPMg/l
QhEjVuVZG0ApwP4mX4LNudnhPr6rDlIE9NGlMS3MShFQ7723LnkMi2fGacpMQ0gG
meJNcAlEFnvTAAX79vc09oOLDHkzz1EY491cWIcW5d+3fPUr8Yns8tHHlO21P8oe
SCnHqFs3Kp5dZzaVmdcp+uF+HRj+41c8ktPWvmLHrIhC7T3DYSxtUFyNhSh/M+jT
bxKAi/wBjPx+JTSdVI1ZQ7HAb3zmh7xWxh+XZELXZIPIaL8vetVQAPS/PsF9fCWv
Fbb3wjWirC9cnAkEE4fOAyFh7qPnFnIBodfvOaTUpqVELiEa5gvCcl/6hYr41E6e
HPhOgODEEDLQAmTcH/EXtpGzMS2X0Ia8p4JhKf1RLGipR1g2q3371tr1lcTWe3v1
AT1fJogtVphZYuTWzzMfYVCeC48izG1T7H0gTo8Jt6UU2UNnO+deWMfO+y9O+GN0
jmunnW1se0j3Yhn1qPBizYERL+SAOer0eGvkUkgW56slf4+YGYQ6ZEpBbjz3zSBC
cQqu48zlvvgh2pq+fxDqngsyig7+4/2fxa94ajY8Z3VE0i+7efZUyndahB1OCBI6
q35nCVad/gtpIpf18YSWo6kdid9jT+mwpZ5DcgTFqlP93He5CSF+qew1VVFjo+NZ
RI6lOBIC+79qUpVUzW4beN66U6oxtPkMDvX6TOBoh4ktCEmJZfm7GwOYdqOS191Q
asf8fj6nypplMJAFJqfNn1EjTrCadP1WQ5hL+ZGbPX7+BED3r6UBXkqYT3mtuPHx
a97lUNdBv7CUTYFgopXVmSGbu6t9y3yMrJJl3enTL20D9+ctonAWGlqgPhrHd7KE
fG/zCa7OhLnm0Qq2Ojw1xDow3pywBMXoI3Ie4BhaHmjppAtvsZ5PyT+3ZzZtKdQp
wWvJqG1ES1U5u4FvZIB1ZF9ujRn0rg7Rdcg6V2GsXEoSH4ROF6y1uJZUIa2icurv
VCKLO/NCN16Z6BQqnXUQYjngG0rZXSLqvz4OIBQYBLoc8ibodu4cR2YLApHzhsAG
AHGOJs0owGuOPmKNfSgq78t0GWV29vYKeVfrwKZBlYERbkT/D/YRV/TTZ/xvDso7
yo2K0AJeVZCGdGFvWzrbZLV/Y1zUIb0Bx/x//LZl7NacM6j4xk5JHINNeMebFRC9
9+2LpoweKKlvApjYNzrPuajUHw3Lv6bezH/OF7fFvdlJCcqvvjljLAepS/TyO1uC
G5TdGbRTAN2bQgUR9rC1/93rCzo5OCAmeRdtUBH85CD4M3DscAbXixKgTvJbiaix
uLSkeg/uUYEGVkrhAIq8+N4uu3OGVSPLiwQr707SYfMyVr/k/5PWPBIfabQTDHgO
47H2bHwQ5hfWoW4SfZwlT8WDdxf804ay/okWAd6cKkuT9zDQxUsN1owR++h2dd0v
AJTkOYZMa+vjqGAAdIp62/b0vWvAudAbKpm/o5eA4Q05sGrUVR078Bqezbvp83N/
/cxmpQod8ZzehNJUXI4++1fLbTg6ymyy6wEj8zQorEmBktHvONIYQ7xwzuNQBUgm
2v9Ja5HfIB9W6u/Dt7zM1wIWlC7MH5wvfQkwHrovoCC1hj441fLb3wjfdwx7fNix
eADAkPnKIPNlMpn2rLuBQ2JhWjLrVY3Rui90jT8yhZgZNL+ehhxN3gBKftVA3GZq
N5zkFEUNLpBtlZlPtZ7k5bTeF4jbMJy5KXHz5gnpZ6hREtwIUiEeXl325EzVVZ7B
tMubvvvCDYtWXdGDomeBhEvkrm+a2Eun0uXTKEcr3I8MBTP302ZN09nQTI83X0st
/5kasMVXPa6poZ7WWGwJIfxLTcGfKjt7Oya9N/Wn07EEtpuh0xnbR7IQJf3RZCvl
tfiJjfKtpw/WfMqhbUiNtcEFXvQeR07jX68M3BEAHj7JKGwQMmHo97BWlYpY9CAC
/L39y9Q7RPvibWxnsSB4N7v60k8cgNjZjbiHCrsX8/qJf4Pe5Lmmk2M/l01fCdkr
aqhIUMAjETM6vDDyr+TkB0Pv9kcc0vmAIDvbYkKf017PazmDSFJUx8FsRPkgCMFl
Y0Y81ZsXzRdThIOXh5NvcvwuCoeYVdHhFX5d4yLKYIJnyeuNwjI3SaukjeeTvteZ
cOHon9rIUNxU5NDYpg2VdlmSFl1EUjDj05fvHfJksLYGEn2GtazcHstNb+48E809
b8ofyTe9eKPUsjxw8ihwlMY3nR3u1LAF15zDud5meBS9rrI3gfLWSThn21OQTakE
gpNe649wEDxpW1FnKmQ3FGZaaujGb1rwf/k4uqjZMZ8QfnLq9OpNGGl1SDgK9Zer
90TK2XiNsmyKtYUEFoaegWHvwU+5HTxmqmh6L7Pvqbc/Zh8ktYdHH8NcHtZxRn7/
PtudloH341GJPOlUiUzjiLo+FtyoBI2+t0b/gogYSy8YR/YUpWEslnTRPnycpvNp
1GK6zf4AJ+0tbjasO58gD5zaJSGpT8Gk+y8X33FPfqwAr2TrtRKcYD16h/j9V61O
T0jL5fDU0akjzvKJPfUckFwo/AS8rpEPTVInFD+WcjNctKDci+Q/DwMvrPKzCmMX
VTVwcRzQvmHiCYj76z8y0NtDk0BZw0Nfbok4/SuTQk+TLxJciim8bObR5U5oDlXi
N+ZvmgATSw6wzNfUwGdlr55RHcjtRQrdQvUSsDEPnt+uEs9xxynMwdZvDSEzDRVp
yl03gLLA390PUm8tDFdtB8/q4bR+uMySZOt09OYxOxfllOGso2UN+0nSSIL0u6Lw
XYU4r+/nohn/blEpCCrJq2pvIdz5zsAQF7VDGJCTqw2GOVbPNjJayG7NgYrZN7lc
YhRhk13moGzsAaKPDSYFc+OM0boX2MnN0ZabyK5ylerKy4jzxRIO18SlC3QfDGdB
Js04whbHykmXqVW5CHHK3g1ZLyk0zNeobxgRsuG36g9I9Z3BKjh0jIuo1gvRrKYh
By1CM7rTgl1J6Be5JFEEXzBNfMUzRHq2SXWWG1uIQkPyIiOjRUQmvWywLGZivwL8
RKegh+YJYV33TK32OgEhsajh8bvWsNOg0dK27TLI3JBL65grX49+JHbRSSjpWmgx
pOwjaSNi6wypP6Wc6sJM2nJoLxezARtmG56Zg1kxMM40LcYZluCkBilrkulhj9r8
Gob0lGEPi3JSU5G1DjM5jlDCGp3GI3jGkJM5VL3yM1/m2YpKHrFH3yOMIUgbRPwU
3aKwkCSak4BiorGnPat/t2IYNpSHDwNsSD5A4r3Pi7N2huJu+eiTV906z5JkXqz2
wBEIQAnionu6j5P5bCAWOGO0FdLVYO1y5tQhHvr3gyuomyZ+p/EUwp/zL3mkcrlz
wQr96hXewuP4WAHEJMbBhvUH/BZSlS0c4pa7Q3RxtIt2prEgkvH8nnnke3VXpgd8
er2mJ/O4OTz4nzhkOwHt5RWz16Q/QCwEJBbm4zn6b39vKrOfnBV/yTocujGgepvQ
ZV5dYUzzNOMRBjEQ0B8bJaT9xZ7qsAtMxjrFSHt1fQ9dexhAQxKhr0ASYMEp0Q7g
+U/lwFH+ZYV2J7xm3o9iXidn3W3e0+yNwk9Vo79LdN/Eax2R/6P71NY06lDh60/+
0ZHJ2JBiX05D+3kkMcyTQjsDGfjvlYPw4tvmeE1JQmNua0QfIIi9ZVjyaHo7Kevh
GJZdABDwqeOAKXz0e+Rp06yy3G1JgeB4/gbqDQtGpUt0PgDoNwqJj0z6wYL/vMn+
ErTNrtW4iAlxq3YY9zXNo5TVGI5m95wPVXdFxFam/KWV0PULqm1zK/w/p16g9AZd
daonZUTOvUAD9dP7YBSu4H+9GRSa6610pUD9c5ZVCFJ7W24VtQIYJprUXwKujFw9
5ciIS2RGzlxVVIE0ouaD6ha4LDDXGTYQ7YFt/JcP+MPqso9RJZfGdrHeEpLmlA+O
XyCfwZx0qYsOVsgM5zqIe+R4ppWtU2kN2QrNrpslIVmybrKoVVSGOoitVrQBGOHw
nmvuLSB16fuZTyxxYekUzm2mz3K8osGLS/I3SBDVoP/DIQJ1/axfG0xUeha+QDjP
EzkrGYKtdcyOLMn+uQG3EJyq0Wa5GJ84h2XZZG2V4BKaSGRe1Q9+WS5p5JqSN5ui
cxWL3Rmz52tOXZerm9OBpucYL8+7MAXvOg8Y/ucY3IUlcBbBFCti4HsMGygaKUWL
mQSHo3EXn8Rnd3aDsGZoVxdDFmFMM0KqOfmgXRHV2AAO0ZiL8Zl+EY+1uRN26jw3
eIwaCntRYbV3CgqXHIQLkfwlLy+ZhrTcPc2EweSCF/0if2VMn0DIQ+Gr3LGrNTrs
xNSgQMJ8rNADfkF5EPhe33Vjlcu6lZSOV6KCjShJvHYzxcuINjKFl+PLZ6K1nkTl
4rDYtayWrafTXNq7OWbheDIHMdnLhMSzfFE++mvXEd8Popn8VbnucG4Wyfn+Bp7l
bKu3isCYMrKI0oolJbnrOPUlf5qZ8wKuza6J4jyMnZRPEb99ajAiegUBGAEBRp9H
5u9iE7MaNOSi6fezZB4jGw21lxoJ/DiU9eZyNVt2a8Yxqczi7uhxy5CxUBJYfIZM
XAI4C7MwIjbQm2ecNf58oDJlJjT+yoEHX1VfAK/fIY4cmdxA7JjdkLer7uDir+aP
qZhk94OvyiEOY7qQAH8x6p51niSlcPi6XMmBOdNcqMwHznfEn3aWjW9yqCVdoQua
AiF3obpxC/gxShzmcvh7eMoVgW3bRqWgcmVvxWNpQfQTleyHMWVjH+Ynm6C00lMu
40/j3j7ptLlSzEw8DO8+ajCwHQqnnSmA98hwCUcdK2peuVRI9QHGyBMC76IEq7Yy
ajYuCww5j4EqYb0xmCD4yXK/JqvgSvQdYkSKmCwoCjGofmMy/lhAUdFRyIsCHsj1
6BpfvrOIBr1GDyS8dH27gl5BxqrOFNeDeBCs00AAwI4LjMPnEaqSxwLZq1laergi
/SZWzNzkbYi6h8CkbYz2wJ5RXq/HL7j3Jj6WIfIgWaaLtLBXNkFzICtIAJDF7/7v
tqXsvvX6vYHg6jhzSpkCvnoQAaD+Bede6v4rf+NtiBF4dFhkjhkuzCHgQ35+xCNy
7uL7COil1ezk/F/fuSo6u9CFqHQr3E30AqAHvl5yevToOm8ofNJlrN5hxTqXG9Ef
qQyYXl8km6wZKYFHMw6b2lhHfWBu6d5rBLeXANW+qPgfIXOhfGKxbweoKFPojDIg
rTOST3gMslV6l1DOPjy+qTnOoDdKa+yPAwJzi/UOIC1leaEWSYOssCRmLXvbcju5
DnELkUatliaI5fFHKO4JAh3Bbs/VCFXtjn9jkMunnyZNfIJ2vcirU+dXZrtHbcHK
ecYHOV2Kd+TmdN/wMj51Dy25/9SPXqM/BPpNbyJ9ez6tl/PEPrGNaN4oXwVXW/oM
Eld+uagoB9gCUNNTnxcmf6GQ03H8QCLSKp1kZMqjUSGildQ26GFTYb8Wjk5Lqtgo
qJm4D/Vt7FdH+bt+VkFOs8+WZBTNytzrXZq1oSRh2mKpjEGSHhSy41Xhr9DzffxR
7NOL3UhrLztXBveHiK7kwp2rqpzpXpTMe+EBWv6ban4YW3mce++vycSMS5Ss7SJe
cmpw1N7oWvlmNokPOnkTncw73uIgNzFhP9Ob4F23Rm4k3EHqeSM0ckgyCW33M4Rw
KLkIdVNSKx2k6lGcumx1TgMVCPlhCyiKXa/K8IXStAHZ2Q41XEhMdBEe+1hWyJZu
T932n4qS/N1zRt2+AVl6kFB7O6my7Sz/wLMN7Pe3SHg3F8OtNaEV+zk2s1kTiwl3
Tqbv3iZSCymLbDnh2cnsn+dLnmE3ltjwxBMlR0f1rvh3gjbgxZUSErEikBywxf93
k1h0HPBWMhNsjsB2oP4Sx1I3UYn6wHE/8uZ2miC/VCEYx24ksMmlINVoWKfrrU+E
brNNyUTwxwby9/9xswGREvltSqtddmfjTIaesRPrX4H8+xN/qe40bWDrwH4O8WEj
qZ/MQvJssZj7gK9grIfu9nlPJ8fMVAcFoJdl2TqVcRyGUbgM+ANOgZWZhE2jxClp
gyFIY8kNduPxndCm5iI+yY+qfwMLnZW/7HXgVPRXMXNwrtc3K5hohL7xAi828tcC
xHgqDd1rMRauSmCTSCej2LRzilD09nH7eljwluyje81XoTYn9Kz1RKWuEwBrSODW
WEVl16xsRUjKhnsVWlFGV5JWjMZQtnbkbHKS250pjEef9JK8ZT0LJDVTRYAW1kMy
gp5/2pmEnwWUGGfmMufYcZiybLwnMfLTPElFGJrnWXOK8sxW3CSsYLPp7nWKEKit
v2bsnGIcQO0dnhnL5hJH4t60wZRibN622T9kuNYlSRfkd1EBOntl8/YZ0ixUoC3O
zfaDBp9zqVIhJJOVUGtZWR0RvSUsaMjZKGkRbauh0x3eLEhIQirtbor9/Q0yK3YX
gdBHyNgmSf28kmZF16Z1QX/XC+3LJVKD/t4L0Sta4pj9oj2GYnNwcfMLcOArOjHf
dnxTfOkmuv7LYTrd0GH6hTRE23hhQggkC26vLdZ3p8mOYUxKM675gaEVaisFtYro
Eiuk90Tz5KNVklwN7pm1I3H+NV8pFFjXP0j2Ko6YGK2ec/ithu2vxZMgFzuanQE/
F+q3BtQibS1ecTqmk3Vchv1/97SxYw9VFGhhcX8qUojReXeopU5KWC1+mpzIwi4p
zTiCQ290Tf6mWHVGxEFfXUDZZAD+0pDgbCTWqxMo3v/W9wfOcbkwiNH0nR9nDh69
9y+mF9syv98EnrrcmhHdRTGHqKH4UnOwfSK0Ub3i8CGlET74F3UXnflE7/AbHCPE
CXSVdClv8U0WECRcnGf5Fdeto0tD8kpEIwLhmI6vMFUt/69MQhuhMnYO9yeaUgK5
boAjl+a7VkXdDcKfAgBugGDFuvqvQF4nik9BHD5dWVAaGaHlDYKzQgbOB3eWJQNR
+ouUag1S3lgmu3ZvDrkQedZ6uQf3auELK2mKlVJ6cndHgXm3g4f+I0Pcx5eC/1yF
xmP9nrfme77syCpLJvhD2MqoLqc1PByjhdFJ8GV1h/rrv8Eupj9OUj0da+XSdDbx
WszvOsYhLMGRl1tHxJm4PX5wfGNenK8YoCGY1K881xV/laPnJN3yQiPfEDp6PrFT
LtbwOn7lWB8VqzvZWMd4RriVh0pmOPTN7w8U78IzpKnTam715aMqR4okkvC3/r3M
NhXPNDUQPITwV6mb4Zyl1o9kEAH7WIGZpt/gA8KR0AYyf6n0OupX8IL07gBMNCGN
mHCjyM/ldqnpFBcGJ/p79YDoMNhvX0Fwl2HzLLxS8colUvDyaPOzf79ZMy0m64Yx
oysXPCWOQVanQ3/v7GWf8bKh0EYjSeqUvBCaZf/9ugOaKvkJ/qPStxE7OirRHCzS
d+cHyCGPj02yjiALS/XsmJCjjIj1hb+g2GJIHYpZSxZHZ09TNeimxVDrfjwp5u/Q
5KHNfjjJ9bPWNcaM35/oB4O9W0osil2niRqQap79hgg8CnDBgGjiLcqYKNVjNUlS
aDZhgD9fylcuO7TX0bxen+nwKH7TiiRZlKrHnNTPH5+xwkLWawO/LEhtyJOGeF/a
0Y0uu+Rv67IYjceoWMM82tDbSup/+6QvbpFMPfFe6Um5mzPNy305cyjWiDQPBFBM
+e07+76gp731CX03C3wBh61IPcW+cRJAvcPSeil7SsjYufKfOOtZXBnV7Z6U+gh1
h+128Rkgld/iDuDcbMC1H7wPQDUu/5kVM2hAXeoDkCQ7Zr/2/0Ks9w4OFGH0TNeO
qQcrk1oSOV0mENBsN7iaYTxJiSOuVzCQ9mfFFzYY9+87EOwArWSkDwXayD7tvREP
ASyYqwzj9YVIAyuooHNnSK+Nhsz9bD8RGp8R+PheLeLH4yqTD4J3onWlKf2A1Kpl
+1meh6XgmKFB4XElPzwgYr/ASR/K61uMbusTucp5gE6koW/EUMd8CoadNeW5c9xc
ndR8KOHLiBnSx9ERCGNC61rUnWl8Usjwqpoep12rPGALazCvvVI7pQN14DZHrmgb
2b9K7k51dJgfzNb1CO6/6dVeJfB5InLLsEf5DiQ5y9nlaKd5qkgr/+LpFkpvatgm
XepkwAap6ZDkYICqhozhLOxBeAUP18dCZoZChokDH7cWOq1AJSMG077eBh3sOLXQ
+/Rae9rDn9rMfVhsBM8QDb+UXSxEegvSaYXn5mgfK6buBC5U/UmsBz9gDGr5eE2d
Icl2V5nFm8koTUQQJKxMIE7FPm6h8W+FAsiAYFTMPLASS9Y4SPlg4DG9uN//g1Ze
GNak8bGTCuguUKRlRWHVBAqs5PpbRhpypNlfqRCp3A/XBmdCooWQP1iAo7wH47WO
mxXa1tKD5fsRRfFXxLdasWQN/lRMdEreQJA7CThahVfgkuMSpHB/Zia3ER6cqG4X
h2DcQOz4gvf0l9+tKvw08WxAAge1xHFy59xSnrzzZm13yqFYSVA0+f6UbIOHtbRo
ljwjPpACbikQJOQkasnW+JEp253PJ+Z9JVVnB1HWzm+Dv9pPzqMyLIuyoFesIm0a
lTyV1zOpJy5YgxQRROvzYEPWm7X7Tr2lOzbQCPe9j9Xn57WUeCdDvKI4GIm8FnsY
JNBi3EIZBecw9z9CZBgUxMMRarekmfRb8XHtjobT60BBevMZM5YPzhu8bxXYhHwq
cE1gp0VTXO5kDZwKGAV4Szeky2m6Y9pefDFQnRVGpb7LSAlI3SeEFv9gCTHPBTNQ
V5V2DdcWwfXiSjAaE9epz/j99H3HUIggPxKAEWrPrmaNdmbQFjHZwon2KjI95lkd
A955RBT2DkRgemV/aozaLLQ4KK7kZXvwazZgSabM9Tp9QP6eJb/IJz5tex24CqGb
HmYN1M9c9KGVHJsLv2bLTX9/t5WPOfXGKLjBCyCZCb+gtToqdpEt7kZ+ZGlbTkj3
SUVuujQ6RxVTxgEOgTkAzvQQ0Gb4wjqM9ta0/KhfDXJzf+gEnDMchd/bbacMT+na
khx/dyZUUJZaU1QmC7bBVU6E+mnECkdVcNZ5BTYjtTslCwAJkspusNNAUXDNsIH0
6O9Iz1SupYHFDIIQb87eaTx3mEr1o02cr0DgKI09pSAGNPJ2KCDumBnb4i+C1NLm
kzoQqLNZUySdTV2u69CjmKJSjlCE5P9OhMLKwecE7FOJaPO4QF0AJJEAgCO7JwtC
WsyxIU9ofF5BM9YR7aAjBsUIvEUILIOAdJx319UZUNg5j4irY8OfzTLepryLYjfI
zzc63ubgl1UhKhxBdFfw7j2jL5mKkbCO88fz4SMdYBZu21+V+PZ3VkOthQ3SGvhK
7IiBa7EjxzECcCHjsxhz8rPvEbqMDIPSlNEz+YH8NWWGwxG6UrN4dkzueg++i6Eq
261NsdrrXnVNHRtUFSIIpmaGFqW71FH+iGn2FHM1oT3SJFuwQ8rtiXM15SaBp+I/
hmefOiLvrCTh03VQ4WwwaG2PBoT0UnDgVpkvksNm2/+H2X7q6t/3HcQ4/iL1w7u1
9QNry5YhvgGG5wCNNvx3szznR1oUGaTM4ZC54OWren1fA/g92pUCfhwUoLqtwpnn
wrskUJ4n9nHZbbfQHc+ahwjNV9p9n4At/fQLbVIt2Ljl1EzY3Q3jlYNQaIf4SbH/
ZyNx0CBt7TXVSeTjHVyTIf2P5VsLnlceg9Qx3RrHVR6nhxe8ojU3ubz6bA5RXL1c
y3SjA5vW67mDhSm9ndvtYgl2vBv2A+6Mro76/x0HIaTRYQf/CPtPDOhnAf1p/Qwz
zA9YlP9N6YYuGgRDjfXn5xhn+zi06r5jAwmkMoqPHDf6+BsezBmJPwFrRoHOHMTJ
/LN+XSjm6MmH0QZGFouL2gmYy0uzz8dBBK/tnmQljtXoUJ8Q/8YmrQPudO/LZ8IM
fzmyW6I9C50n/v4Rsy2piBvbrfVn0Ebqy71h1j++uH+5J6+WOQrqjxDwVY/gPAjN
5M6/tUz7Ly8MQjV9RSpnagykbjOzH0rHyCPkvJbUvUoqywRMPn7fWWQQYCL9dW5/
RiwJUevRNTk4WSMYdVmTFUcVB6BAlaSSFBBlp3wCp7ltbx3r07pGaiDZcHufl9fe
rOnyYH9YNo06sgnhxbxnZ3GVxHCWg0ZumrhpgS2M3iVQfGwbGSJEjZSsWTGgfCvp
Svqaiuj5Y7nBgcwCS0ptb2Tz3sLDn3vpIWz0EM5exMjLFec3LwdhOZRKyGbpgMoJ
g6y/0oRIbwK4RUgc1d44wUca9rbWPFH8pTK1f2lFl0l9UHAFbsBOrij54gDvQ1Ke
+92FijgaNGJWxWf1g9GsTPDuMA1G7NG3Str2fcRwunF72f+MhVplYuAoxkmLVqUs
Zc9VcsSihH9VmAqV21les6QJuGb+VTxXHsK1JS8BKnJekRfEuyGh+X538ubcL0uc
niBIVRW1pDW2Ed/Dj+1hn7riTf2MCfEqzbQ56bPFSzYJexRWjXe5HEcHyCxoKXUf
HndkBgUCOr9LFmLFnP+2FlhboXrzL/qjbdap3vx/NA/V9irp/Zhd6ZzwNlq1BzIo
2S4f3yHgWtlIF53MtYgLGmtswBpcsvDfUzEkw3NTa3bRdwInERasWLdAJph9+7S8
dL3R4vy3WRCUWoZq3cCTwKA1PtdkSadTMQCdwm7tvVT85yY9bsxWrbdA8mccTwH/
tvKgEvbi3VG0L4EVtdGm33pZKxdgDaTzQcYzUaezc2Ih+OM7V6+DHj714FIQkN8H
AN021aXq1+1kAB1IbhAxYsPsXm39NXp7kmUF98VNay9lJH6TTYDyfji++RM1VF4Q
HSEUuB38M20lYtfbEED9tJ6craoo8by9nKywdaq5VSCt1LUzIfGBUWp35h+jn6Qv
BPnEKw99O83WD+3WkD8YaQMmHJh4QUzqyiE4CLPoTvrD2028pLXzMnlJTs9J3AdT
5HAHAvWHlHUSz0V8YHjGeo0tuOxRTmKMleh9gIIcXC7zDyvOlJI0JjLbC28cesrK
QQnJNMyfK/UWl2FGJLKZPNfeZLg79zwe6BxYOWVS+TPPXJBBsyZ5+t4OokWi43y2
BQfgsNMkIMnlc34ePwSpyhi29uqSXNVmlJAI/Zb2LrR0y/sS7JHxJiyacHkCQLZu
lf7GJKBCgDF+miFgqI32LV2bmJ+8gWhtYVSM9DA4as46uGsPIuM8H3Ep/X9Di4kH
/as/wk8J/c1R0LotR6Ddvyy1W3N+9SkoeQo5mkLTOJi/3c6f1GxJqI4FkmexnDJz
uhCk9gPMDyY53qgN1b35bXvnn6KtuW+zuiqzy8RxNc87YI902vjE/HZVezyJx/ey
qTd/QkCtA2qSIVB0ZciFuqKRbSeoykwXK+WB0KoIYuiCkZ0NJpswfwHIHExN9BT8
78lQH0CdfSCQJ6V0VtvK7wR9wk8lLBdopCGoI273aiUQimKsp3YqFcos6hYkejFK
AdLZLj6eVUWCrlm/9dzX6IT/79OgvoC5oYag5ZqL8NP2GHGPKsEZNOy3yfSG1wgq
jiaQHNT71uRPwDhRp0PkLYsrFg473ifrGf4AGMRGQ84WUSShOwXYQNtsi3Ux9+BF
GO3LgTNUB8uyHx+N3x098WCH6WEkXwDLebnWNQSfSLqBWxLIG3mMXsAh91iA9F4r
DF/IiLMvWIUvr9g8jbBJElPiv4hBwDp10JvbxPgOut4jMSWIdbWJXQ9VXu+DJ03/
OJs7eXcSMmdu+QYoaxv3GnQUbdE1wEFjXdpCqS8W2rP7WiJBH3s07oFNhRgGHhUC
5dKRKtJ1SVjcYTqft9Tu80sT8Nww/U/gNStO9o9DVIcCLnMElFebHwheKD7mM7ZV
PqnmSoLAho4HrzKsmkl3LQxGmOwYhBZSU9HH6ct/N5yz8cFopMxrrOp0Y7o6R//3
aDftIQD995l2leWWdiPp/kXwVK9gLAQ4ThuFz5fl1Ro0v3CRF7z25qPopaE3YOIo
FQKrlmzdkp43JOdK+Qwexhf5l9x5ukL4ksEIqvjQVjPsrYzIgcVYDF1eVvpIAFi3
tVIkej0M7reDS1jMpR67GoL+r7/zxJT5xxtKuNq4EzPrk81yqwFFclbA/Q4/O59Z
emuOFSFDY5Z7cgbqWdM6zkChzigPYrOjIwisQlU2H8UYHofrlRx8qV4QkBG02X98
MfTghDyjpGxkVHylPHf1qpQohXZleDnglve1qnwdQbyf72Jul+P+qJ5RpraD+WiU
vajI/saoJVbooLYg0MIfcDT4jyeZnvdynF8S6yCjbkP9QSrlZ4lXfTweQbcm33Oa
/zEa2MVS+7VfThZD6o24gcvJ/K//zF8rsS20MNtHW9SjoYUqCCwxO8cln/cvcwXv
pn4s+2ouWRZvsXNisZOLnN9axRnTxiIoss19R7tYZ0gdcU3lAt1YVcJytREFnrlp
f1/jbAN8VqSkH4heVcpHax1qLz3uzeoTWcW1yX5sAEVtWqVfgyBduqNrMs/oTkBk
zhFebNpQALpMlKDn2t1rKBbCEw8LKi37mLYt4+qlPg6wasq743tQWggPgKx0Nv0v
rdKKX3+Xk08n67uqsF3KNOMg7P58mkK6fT54o9NOyIBpNWeiWwWV5+HWHagwfAUi
gUGm7SQMwZM0S8iLYQ+cniOst5S21iYI+rM3EjIOYq2oM6320vBiXqIBAYo3lioV
Y2K7aHPbku5OMsIW+9IJaeyPTOe8Nv9ScLXrYmn2OgVF+ShZZlEus/S2+pVJ9Oqw
soMdOt4u7T0HU0A3rZMWd+HfjZsKCCRV/gm9QMAeMTyMwhYkxEDCkSH5seioA4qC
c3+7AGMjQOmLdPgG5JEuMAQ5yYIEg3f4VBynAUqgOkaEusNpQyF6WR6dQ5u4Ts+H
1Abb633jI/oYeHhCDpkzPqq0Z/8GB1nkBXyKQH21ucd4AnY+ORkwcBMIjAcqQiFZ
hq/coq3ARMMA2D7Ah+BKJ63j2MubAuyOUlySA0IpdrEcIE0DJNteOtwAt014WwB7
VncYJhgyupmjbKHA4RCmFkT4czsMLY/7x6w3NX0hbUhsIlzAt/nxDdTwVYwCjIJB
dwo9xxL5emyQTqa1EQwF1cP6FfHYyb+kQrOafp+zjZ+xhmmVQNalsKaKUkUE0ejz
HzpRW8FMHLN3EvHYAF93EZFglPJ4GWHSrNbC3YkSogzPbcwMa0jpDyL4Fb/PDArg
lGA3xwfFxwr5nwwqgUX9ZhCdnL06IxZAfrGBaCKHNNlx+3VETk2djn8vNH8VOnTJ
5rEKQ0BeP6eai1HJewKlep1RJVi8Ydn1PggNTTxuA+X6kIMRxOim/aNyjOFVJ+3P
nsUwB7oK7qlHWMUm3gN08l+QP83sNtZpvntdo4kdi9YmqU4TbxuFPu2fQlq/0cA6
tAXOBGiYtiZhozd4qEOSjXBuVPRf+xUyBCvuGxraTitUwtCFsCMNS+3eT9XtyDr8
1PfK/iqezn2tenxlHCmklDECNQkrdJEHqBY2AmvOlN0mQMjHoQvmF67wXbdKarjX
aOfwEldEBVAStm1Wh8RobxrrKlxsKxb7rxeuCP6X66db0On350jtFZ2Y11uWJf3d
jQJ2Vw2ZKJJ+k4qr1ItwS1maj4mnmA6PAycYSA6qi10+GoDPlyj7b2PhGa1pTail
QUa71GQp/2+NMWeZA1vbxwXkzEGpk7s/xzO69ydak0l0GQl2Natx3Tw3okxr5m0S
yoDPfs6c8oOy9LCKaWghN3ZVe3c2jhs5eEwGG9SIqo34fW73IZe39sXNzW2KmO4P
sSNTAE1nWYYjJu7CrYdbp9UuBhmmUS+p88FNirjwaEl3YeHWBU1sw7/fAUwF6Cf3
5A6NvhrAKp4tMzR5B5TATJAG2NBJR2jFZUNKVrFHA3pODUYgB+jtN0SUsDbgGLA8
W+f0t134PoWRtgVn+yg+sGP2DEoLgBhZ8UDWiw5MVR26hc2hPR0ph9RJcTVxlhG1
ecCAT20g+tNTRkgJ3bYxvQtsEFd8vfyAY+TCXqgWjdzoUDyHaAPVmETsXywMdcjg
yE3DAaUOWUv6LY9F5DG0LCRG0LqH9CyLLUMj1MuTd2pb/PdYsYB8Zu/X7nzc6i1Y
C2k1EymKGPL1+buOChVv/7GZxvOvfaylbA7dLWW2ghoBGTAwK/uknnFTKG5qqXa3
ANxqVcj0Ydtv6FImMF/6H631VbwKfyiZGsH9B3KQ+/wvQAvS4a0hHPMFi5KDA531
oo/JdlMVc87d9/ickuarywgUQs1ExfIwwh8IAOB/N+XDrWrOvfvosWlIpD6MvLHq
1TfNRa57Z8V3qikHRIh6//SM8wRG34NKrr1ALPlPRkMVKCJuw7drjjyEvmMi4Iv7
15Ur4RiIT1yeERTwqD7S5Qp0W3p7idXGtKjhqCjg5PBPU2PsWf7wea3Mom02cFNl
RW740OTJYAAvY4x3B55bROJ0nsBkcyxEkR8xMsHuYmny7CQVscbmF4PcH/9+L0k+
WXl9GefbLUR41aYu8UAK9y3obm2x2ti3e1daCpRV8ERCJMdBxSi6Rycdr3b8xB74
RVclhQiFeM2sqEM/+9WaNR6hI7dnst6wS/DLuPsfaB6zoe0zCY0mHcwioKZOS+/H
vUVeNHpnCzaHYlIqfwatcTwOvtXEQ9fDrOeI2xD0z1Qy0MbTUdYZ8hwvHbSj5W1r
8TxP1Q4i+9MnVPH5qyHbsRhbMWFz6Uh2ieY05/djFiiVA0qv+hoXK3qw9oRpW4Ae
gxAzOXA6xFPAoRXbXsv5Jh+srg5vPweKuWyS47ZHaBJSkXa+UdIhT8y8DSwHtxr+
Cj/E1CUKVAgkUzgLVj0mWyg8PllnU+mOkrfToWSBTNcTJzu3K56mlMT4WQQEa/f4
pmceQ3pcxjpaHZaGRWEyEF8z6MgIir8NrZFrh3FKNoTs9jxsrB7J6n3wTwRes+mQ
XQm3awIcU6FAVc6sIyIkgAjCuPvRFhUCyoiVym4hE8Iv4Cw0NQv0dfWCo1r5JtQR
2fRqF+wTMUr6A6+Q8gfgp7Sr7XbPXQRvYXNVP/tfSW5vmLJVjGK2w/CX8mrlns4Y
cvDvKQAJB74qTKmmIMD0ySmTouK8NiKvJwDZXlb/I9A9yBsgJLEr6LwKeb6wUmzg
HtT2fa12HF36AG+WX8RXWCiv1FgY6IERrQp4UXzBKsJjij0deAVl3khgZVtzXevG
WTPn6gj3EWilRztfbtO3HarDz2D1YB80g7zdZL7YSHxoVLEsajlIzXxEFQD8mlLb
ChnDrel/0bJnL/L9ao4X8yu85FghWg7EslHeiabUoeA5i9a4bRLrxUAi3EN8Gw+q
Ex+o/CVmPRI//Kf//JtBB7vAU/de6+jWldyg/SOR7/8yOemuykyfXz+HTFPXJV3f
gn9DGYtLb9wAzruqxA9hVbOa0MHrgd+I3Lk/9ozxrnyhL2WRCxRvOTHfbz9bNcQn
QcDqXxWaBcruRzhFl0huvdqiwrO+JtHy+k0rd+PJcQwdEWIu76BQf52wJ7gB2/uX
6e5YBd2sKKqsI+VaPIrqTU5e93ES5qH1WhKgeR1erHakE9JzwjqMuO9b3Zzt/2kB
Lb27cEcNvjYlIUGHtRlsIXD4KjUU/8DVBU0vWvcNbcsNo01jO6eJbGfuoHwyltRy
W7dl8RERLK5yYykUGoh7rieks12fzMdXIkTG3xJ6cTV1vQhVXKRRew9MkXa3Q1g9
JrYwjQEm+hJJ3EBxF/1ZkiHllmnvWWERcDg0S10HccK0wEQfRRI0np9yckNgX27T
w+RfQTf/Omslrqu6OYY/kdFSxh+0LbP4tNTETGGYcg7t5FuHxCLF/YfW5FSN/sVy
DaSKPYOYpJ2pbfaKdcHuRICix8JfFK0UA7T2W0/If4uFjRQx2aiu+jSAnfXRjNwz
llFP08Hylb/nvT3rVyaluZVfyNDGKZqUN8kgLK+7vsT7nVisxTtTAhB+ZdXztGF0
jw89AAA823Odo/kpW3MWqZ2Zrj29zYkNiup0IquYwUea7c+BBpgwkV3wKpH9GVny
JXGP2A9lIQTVdnFzqE/lokV4dbT29lymE8Gguix7FCtrjD6KR1XBgdP72gqZe9ua
AMB0pDZBWAsrqBYW+LgCC4pUYCjCYPq/SwPBATmPDLudGDimwrtFZIMxm9JgutMg
Fid06v8G0IAZbsE57n9b566Dd2YBOpQzCUiv9IX1NR2k4A09AW8GZ1zTQIK2oenF
ARdIpb/5g8E279kZpcXr6JqDF1wPM8to5SybvsVUvwgstuAb1LT7mA3f9OvXvwIZ
qg5dMMq3/BLJRgrZD54Iy7IWVzhFV9K+joVEXYD90ZnpHYszqRArjVMfKlrsTO3Z
8FgGi5XJHwMAQb3TBMKGI5VwT41dJEZPW1pfQqwHYYy5AMXnt/ZW5Ck2E8qRSMvA
/LXfPVdHhEKtNNWKKFZrMrbxzcSjkJdAtk49i+SZD+eZoPa+9qoCfao4KIqEAlwa
MeDF+8nzPjxX54+K0H2djHZbrPoVsD0cd2ZH1ZGjJS/6qBG0P1QAo0W61lGKctuF
BZ8TGKd0qzxxkSvYg0hOK46pHcxCZUorNzKq7FvXC11ObI5+X6rNymFKnuGpi9bk
1QJO/qyDevvsMgAmmvzotdEcy7ff4w25cJvnPJSu7UfddTaCNn6jWQNumaXHkMn0
MvJPSgLyV17nQUOi5QzVTytbQZTcCUf0sEj6GALzF9E6K05YO0BzzkFQrvT6CBZ0
McH3eotMnvX8E9NBJs8gP7fYc5/Vo/JXFU35p/4SqR/VbowI+btCmlPM+/H0DNiR
s7o1hpR4xQSArKARly4J7Y9RaISO5NZKwvwGKCU+VurpaDRetCjdX2lmh5WYrsKM
wNdyMhSftAaOCQL13yaj0amuJPkQLOcbUkLRtyuHuOnrJb0NuGiuIEAQ4evFYr1W
1iNDco1xOlEwWhb6hq7vL4CNV3ps8vRrJQuAj7D57JEzTssH3NhpPH/CkBAs9pRR
GCSNJAMN1PnSO8cyd8gA9DdoOw+D+/bQ6HhMJ3OYP52jHk5yoF5njyLbhoNblheT
FGwQom2Poby1vv8tArZMUgMoujro3gokrkU7xbUIgG6MKUgxQYf6ROPh8J57F2Up
rtG/vL/11mP48rUsQtwS0QvEbSkNAzQuLgeJOD/b0osUKJ1GV6FxHt0wv1mvU0jK
36IZWxmeUoCo2bK/1gVsj8BOba3RCnpZAGeDGwnXXcPvxsS8XCZe07OC8CAYjveM
pD4Ry7/VIfOPAEAz8ygPPJyWkST/wS2X1QkrrMCRodU8DzB3Itzsc86eKQT6hL04
iMXGEHoC5Ru2x2i1pWUTizEhDKKVklCxuTSCi+nMnxVeLlI7/yTjqxS36fywcG/r
OZExmc0TyQn1Axrig1J6XqUspuXdAT44yzb4OKx+ki/e8d+sQ7QTSXILy06fFQqn
nSG/jMBKAx/oRs5YqOciVOCx/i7RSMmv504RwW0DixbC0cCkx20TaTOgSD8wDFc+
5Ks+6wr0ynVOAdDNxbPwzEjm3aro+D+FDXMWSFKhQXbKFdyHbgMdpJaJx5eAkFfk
MbL0DV+6UzxqvxziRjodw376Adq8K+Q5sEeFUpkl54JfOwQ2Oy4IHA7CFa1au7QN
Q7kbum2qXElnamx4E1m7I3Bu05HPwdRln6Wl9InQMfhPZj9kCxCVwimMM3hUF95Y
cO145iPwdvfY2Jly+StIgKKl9o7+0IKSCiwA08v4G+0NwVUwwmeTe+l74SLPV+oI
N6H/PwYWKFSo21Q6xWzT+jANrg1hq/PmoZ11aaNAM6lX5zKg5RRpk0A70uKYvomE
jpXM46500B54SaCliCE4cV33eAQAgexHx9ZRnu6rG2u/iyQlwzp2iiuaS2CUTANv
thgCiFMVQFtD76v1R41W/EettRbTn+c6Yn9BojSG1iEveNFsjvKqwosiAj1SK6fO
Qkuo9VNE7wvUfCbliurKV9a2QBOi9YCPngvXWTVpYDPvm0osXcRq6PC9+/NVH2EY
D23AcLU53PSO6vpnfvrsr0UfJOoKo3pYhhTt/hr5w/+ZDmo14N7QZkw4iYCOCB+z
9BpvnwjqIm13oB7aQvTwAwMvF4i1G1MKVjopBg3/GFo/QWETE6zUl8Jo/ElA+ima
tNzjbUGxOnMXKqdEL7uiqKzcWeMwTslQ+m81/lkIIFKmrkunFIyW1humf+H9GW0t
12yXlCyD0WIk05Ta2EXMcf3z5I09r2GX2MKoEg9mMEHMbc2hWnAK4Fn0Ru0ctDy2
oeDumVNXSfKtzqtuHJIK+1SqSkibudaUlBU65br5P3nZpdQHp/esMOBjRH1kGJe5
eRgbQd+dNUaocYMobjSrlBngD75zdqzFuEsOmf5tDZKUzk1inFks8ptSkRjiVNNb
DGVuXOqkf1UHgQf+1jRhtxweT25hUvNd4wVl5M37SkNdsp02txqUnoSo4zH+8mC/
b8w1zJIcCdiyRCP3UtT58YYZasOKzao8aW2b4+Nd9H5GX/ppSg2XHr9qJw6fLGfY
PxUsZNGAf/l9LGyrqORPisVs9wLDJGYdmxL2bwxq2DauP7IlMtgXPvKkxuW9jb8Z
NfMp3O8CBHg0lCmTDKBqWdSFFUPlGBrEjrC53WQQ9q2QbcI6x/5jrGZHDEhUvm+w
uCc/ED9VDojN/iHRa5ueLS0pc3rOyNl9EvLWbh+fe1eMla4E5UJN4sX0VBCi7koW
6SqZjj4i4uPySsWkvf5sDrcJF7p+n4CIS2t3AxVP1/C81UrqPXFHq4zZubR36iRA
5k9f5inK3bjkw8HZjG0tgn0ZDH+bNiDdS4HmnUuNQbEbBZRrSqhFvPo/XtVqRMzJ
PshY99wpFmL/Rv2SGp1yJADu9MS/EUKPHlk5A8SKRSa3j3+gl9imfbbAMePHO4cJ
ru/fn1AQVkHME27P46VAeor77pTXU2OmHV+fbX3DjnYZrcTcpKPWF/rmMLqacxb6
Ir5pmeKCoVKndQzqy39OgE7kts9h6hAKD9uKy9peYNgSLcUwprCJnVPgJnzrbTyS
AN1Wxos5MH+oskrcUT9lZ1adjO2qJk6Efnw/QqHeIq8XvZUy5Y9NTtJBvYT51ZUa
Ha8WHdD4SeMLN39Uq2pmMeBU3jWVH1OGS8BMFAejc/NUaomVjf2ioV4eeQIyyYvk
uYImQu4ExIt1iO1o0TDusBiYhLVNfoGld1sc1b3I6zI9/aYycgRynRsxzeyaAkvQ
DKw2zQuflnwTlysB/peUDbbWV4mDJgQySeL+nDi9X3HRqu6hApH+VVw2bQkTvNK/
l9vkS+AcDHhETPyxo0GPc1yg9vU57SmKQfr8lZs/QMrGbSgFhizQxD+p2E6QxBQY
eJBSjomN/koWGPAbIPAwF2EXFg76dS7Q+kvQXFy6FvSghAuoh/IsA/LsKoPYooQu
rUM99wPvQaUOZUU0ZVERmK8jdb8pT1K/uDzmiCpI+Br2MKSwhiI3jl3ILBQycACI
pGeFrJFqFQmGuDaM2U37+bvY+G0Wum+smvOtl6WNJSQ5NcGcGgK3jGHXHfgm3Hlc
ZPFQ5WZQOOlfnOKygQyaHQz9COMw7JymO0G1ow6gwvNF+gcOz0Zng1F0/AVubiB6
HTuevjNFTDUwQzatdB3aJDkuckMjf41fwIbmXixA8ELS2oz9XJs7D0vxWib6oJbg
pWjX6gQhxeGZFZPQ6anVnKmVJjlYDB8Myob8wC3ti/7om+QzYx0ct2gKOZl/jAxj
sUa/qCQczhzpEnqSlkCxoJ1glNNg531CbVpUD+SPdx1XCe9+ko3AnOk1wsPqRk5d
KltlUfZodGnyOWeYewG+edrXl1UrxEJrmIxWX0QZBryE4/ODtRCFzbs/52kXhxiy
3QItrox535NRl4UTOe8WtoHuRC7m/DiHVc/Y0lytTzcTfFABEBh+d57QkYaIRe2h
+ukjx6/fbLlz4nuYbPxCLCSaDqgZOhAy7d0bvtH1L+wBeH0fId88bDwn5uU8Fxk2
6MtGAlVV/Gpsb7OLJIYArQ1NRRXoOATV6YY234Agh4yMdHoSvp2j1vmCAjFvSmW1
SFty8fqCwB4uxaJvj2Cs89oUSstZzh7jSv6SZ0ARWWmarP5EPwFNz95zGSEr4MIL
N4mMaNJ4DrbdzSFl9L+aJDC4zV3YtIKNMc94Cp3R2VizmJBAQ+L2KRilC84kZUKt
K+pgikCdFJO1j50jfoyA5Pgmy29U26vXL2Or4OD0QXF/M1eyxkeR1hjnp8w4lhbU
iGSjlcpeh5NORgo+J/1EPtrAtlTbuvg+KjLItc6n5GP66nFNakN0oe96saYQJLXe
v/2p2QawyjLvgQswkxrYZ8drg7wMYlDKqrLkLq+TT53WU5NvtyF7/CDo0Yw8fIQX
BHS1nUhLjtMcM8ZHFzzpNc3WF6icFrCR4TGh7ZqwRx8Z3F0DbqBBveLO9WRj9Mxj
4bXahVxsMVFGmLqnXSUvis7TLRJuOZlQa/U2hImQTwZ51VuY8jI03kbqLFdF2l9V
yUyBRJWRBENM81/cBp6VtJgFkMqnEtbwIdOOu8Mkqy5nXwSKsgaqfWVUoxp4tIe+
boeuz/zJ3EfIslAT5kH/7WrEdqciiTcz3pwUHQp02jOg2+WK9BfGfWwBmnaySTvW
nr7ZauOwu1Upd0zKIGX2cGOuYidp3eqnuQOHnxpLu0wyQ57McUJMMj0KbOSWsnRu
WBnyGqIGP1eDSPW9eXauh67q3f8S0pZE8sRU24FwjsoJ5MOcVE2kVf/c4qqojV0x
Jt5MqxzuxQyxGTcil0tYZSagmqnMQz4Tu4sfIuPEDi/SC/Ed4OfqXnZSfYxgLuPc
xM0waK3KS9Zc7udAyo92UjjBuHEIuymv5J4OrhLOcYpmzZmF+cJlxvAhkejdAyOB
DYhK120hBB6lxSM8ZB4j+RdEZqYeQqPQ0/Fe/U3T/SSDiAyvv9DSOGVig/+ZPuyD
Z+uE8dKqdo/ZGoPXa3qGjYb77KYp88yIUV7z8ZdwmhEHD9zftjN3+6ypzhq/AhLf
v6ACK2nzub6ZRymnIOrMVNFWNtmxgoHWQ/CYFOeYSSfM+vYcVHMtnj7NyLfnrOID
o6TG4mY6CkshwjH2SGUIZLi+iVlpkvYUEtF1sgWEQMXA+fBTi6f5lnrSGtTe2uBy
wuxqlSieE/4qQUBI2K0rF4rJVzRiiBdctV85PDHbQdoQv/tyLB1EVs+6+ZcDYuvM
tQYi9RrNDItm3toFZS86pcfkGeuYyp4HWfFinh0W8y5C68ZvVbQVOQsYAgV3RDK0
2vdoeojRGQN7QAFhCfybKfnPLz7d7QFJXkhBMDxtpw9w47s9udJMIaHfOJ1OzCKi
B/mduHUpG6+4KH2yP1E3rlc63423ldgPfSTS4W9gUWjcyyQaBqjlTNrNwJDjhJob
l7FiSPbwVnBoEyY1ppFWkXGfB8NG1X0Kp3fgZVowyzZocCUzlg8kjGFbNHUUXv5E
bXumxbnztqSThlbZQg3xAUFbce5l47ZIaEsCnw+FpU0leqY9xbRVD+j7x8ko5FsP
xzjdedsWLdlio7sadKeGqVjvEC1N93n4wJ3k8PVHld3eAq6NkDUCd1O6VKyMqcoo
KFposV5ZoJ8SkOMUJZOHRn3MecY0gDXmN6/gi5EvNhTlehttIWL4jE2LlIiaVplB
V8ycFYr3eDW6qzo8/KnQzUluGNYDZOCehYGYHfj8sX/Czb6IdmIpO6IsDYVkSAmn
X8+DwE8KMa/PZWIMg8qXxsieDwEd//DmRAZFBob47V/2MzOBbb/z6aGMtsVa0d65
4qX8iekKFLWfjAdMVgYKTglu0gJT7J71TIZCLRaLnB2F1HZraL5uRggQkqY3yPAb
hUAr3/U7zEkajTu6KenzSWg2pz7KyWGuu+dJ8Np9+akqvUCK6or03gXNFz7c5iI0
tsg1+70aEG/6toDLytlu3WjewQkfPK7BqeJQV4C7HEmLWg7V5udPT0q49v6by/VX
OZd+Usn7kIVfmFUCB17rbbFufivCNdUK2ji3yj2hEOGyYjL/+MyyUyW2180wikpu
D0yQN8YK4g7/P5HlEDqjfO/6rtrmiHC5trzU3rDRk1qjDtc1jwsuNvop9l+C8DY8
/k0u33YMJerzOI5sAc3+9uATvX72NUJQw0oj6HyYomaG2OHbnp4yZSssT4ASL75T
/vS0tkKveMt4D6hm8rvlCxCCzW09fDw1l30tlAapRoG0/wG+ftUiLh02KtBZR4Ap
az5WLOeLEC6yzYNAtisoSlDhi44Hsg1bNY5aOKmwHig4C/WxuNDXqWDbKkl2nrKJ
G3yDeuY5mg1s7xihLqCrJCKMSWGvIIyOQ26qcW5pHpjWztXu1uVTybHsAofWhNcK
/BuDGg+0pbekZqGniDohI6Qm04+a06bojo5bnJRSVazw4uhSzahedAoNepzyrnBC
ON+CeufZdvljxTayA3FWOjPmGsiQsuVhzGxKGR325cJ96qjYCVJrp6da85hopvoy
m/Amt1fn0YM4cjrCxVKJoSUovGpZyqIESgf38sPUVWlvAmGx3TIZeB+u7GUF28+p
0CTW5NMfmZiPkCrQuRWqCQt0yoewcBHwOLQUV238GIQCkfdWyJMg8L60WqFMEfhN
JHIw0MbXJGweySq8W+mezCE+bpzFq+RAo+pNAtZbaDAgCvwiv3eSmaSqce+TKQfK
1ZWsnQccc+nWjx1GRtU63OM8yM6Or6UQQpLxd/elTmRgElL5lmI+k2BPU3MZTUxl
7TghtwcecbOeulXmIPqThXBWlQsk+XVk45GHboTtC9rWLQ/HA/71Nok82cOUVBJg
kLQa6TJaKfV5q6Vso3tqsPkOSd+K16kr5vk2WoZSxKKXTUdmi2rc1/Bp3tEKyl11
WEJl22fKJX9s4YFFmv5jEk0T+gzmJM5tBeyuGUWTCZD2MEIrgQ/cfJthRsMs+TGm
ogLa7UGnqQrZat4ZkZ7CxIkesFMTHg4bY6IbWq+1V51JaWwHACnufYvlDNQrgImi
1OT6sm4Evvm+k4IlBOjGpjTu2e2+H7jirAa3/tnCtQ5LEc6yLhu+C4GpEAmskkf8
2V0hLMLZCLK9rDS6EkIzPpGmLmOOw2kStbyZ6UQrdAgyU4GOAFN+J2uuXfXRB6bd
3v36EJcmYBmOWf86Nm+9HwtaoHbZcQwly0SmzFUii06IYjtGpAe22Tkt8eLGqaxV
Ogey0trIHlcbdW7couIVJzkHL37Iicaf2ayLlR7Cmwv+4W58VRQaFRDUlBFrUCzT
5aocUvdXF7iz5zjILLvgFcW0FS7xltOWMFqrTLpc+zn5E44Y+Sr1fgI+Uqf4C1si
0ZR2BdtJtWIZCnjbtXn1+PxWzmisFE6jNqKVrlgNtrU943n8BxLtFWR0kaY0GKQ5
bck1UWumCNUDfbkF1tb4nJs1SaqlsMQlRZvyMfZ7v0Nfc4rQgANTTLd7nj+KHUA6
bJHdiTsamGNFeM7jUVdbnfAOB1bwmcjq168FbjNW/fWkeWiwRgaHR6qEkLj3LI4D
bUn1wtLTmoFNnvg8/oFlNTgWTkPh/uerE4JU1+o25OW3v1RCPldJWw2eBZwbYHqW
UMSCk4umtGyKJc1FbiVWhTvRMrf9W7AoGMwixQr/iN+SPuLqkLzPtKan5pVa6kLd
m9KMx1E0e3sgiBxfkx6fu+b1LkteKoehbz8AbqL+hxw8a5jDADwUpM/sEsVxW9xN
gZMblpIleEvbkhg8RQo/tiA4108UkeEe3pt+g+fGLDffpe0LlTnvajWSh25w7ZHp
gaCdbfrEVc43sqMzRzXLOA7mOvjfOpNM+OdCPmbLqtXDtFjv4HFyzigTongwYelg
zFGJhIs+z/UtEf1AQfQmXMDVfFtgCDrDYdSiu9nyaccB8damUyBcMA/t9KV+eOzn
W+fEIxplMtQsT4Td7VGvsTbpxb7eQCPaTosFotPXinG5liHDuZxnkgSGY/VOtqUZ
4kAgSylsagBYrRuuO66cK4/6+1Qs3Y3w+RmripJlgBd1zXKVqZEAP/9pjCcfDJJI
gH+hYM//M9HJwvacPuZ6HEb2U4OHT5wHQ3xo37Ni8kORPxDG5sQW0MJrR0l3J9zc
sKWHD26mUZHN2Q7hSchM/+ALQRADT0n0lLTFy8NIHuZvXzHYjecBi8GIhclA/v96
/1yJ3Naz5fM5ej4IU+29OIG0Ub7OdRM1rvJtqSnMV30leN0N0ygMWp2DZeahfU3U
+l+hAfzVqRyMct003S/GE9zMUQxiW3LFqq7brkaZHNG7Y4wLa8lwyKC9K2MeNpsm
1OZ6hcIEGGgV+mTQUNbcR0URkhC6qq5oJ9SyjgVAPoIXecwOcA1hVvdaZAydHSe6
egu9fQ5+1RKJRui9zb1irUTU94LDiWyCyc6qshlpmrLHdNYV2NHjgf4ohl66WPP2
fAwMM4ernrt42X0cr7ZD6m98GreoXECuZKKXdAf7WYvYMTY6Bv/vq/6UHLhioR0Y
rAbDeFgQw/KmBh0zY/M+5mrFaW7r6fSARMOt79f7FJ1uRzsAlmv4eM6qp4EAG1NV
WYjIy0z5JGq2IoDbF1BYDHYy5OzvPYYxkTPdv/yLGRxtWRQcMXKKaxKZYDS5eqKx
p4/Pz0MS7uSf7/QvxmoK9/tBSk6yjeZ12Z3GABqFJPLiZvEoXkr2I1x/rPPSvlCW
M3WXTifZPbQamvRQZNRpgIEyiDZEmvVz1swRIQ/SSO9aYMfuMEmxPm5ySd9/+RYO
NoX210YQCiYcF+y/jCHl63/Pttod0B79MQ95L/siJh36tRdVXF90YZwvvFcsQhai
dFR8qFbzPSv18vuIAwo8QJY8SxNk1+CiPyU7kf9Jl86afbC3ZF+63R2YVuZeJsNp
MpPb2upPdG3u8tS1L+L7qti4l4+7GC0YbAXeFxF/a9DeGdD6SJ4jfRQXtqJfec4x
W2o4Y4Yu/y5Etpjkcc1n8SXjly866IXrbETicGzOdJosF/o9RDfI4TBOxzoM+fLF
IVTsG+2z4ucWqt4btVByDjLd04+nPXLBXoXyI/WefCGrO7w2Z7PQ2ImsY9zAoSRr
i4pxEcJvDXi5/wKE5Fnh92YK350hGpP8UaznnTofWmvAH3PZ8hz1qPsJW5k9LUZj
3NtbFB6oSaIZXrF94zrqsukr/32bU0gKYWx1zfFI0TuQ+RvVXtVabV/+5+BomOpd
+3eItJtqrXDZYJZnJCMJSC7TnQaE+aGigmBFsMEK7jCvEGYHvXKSia3IScqY1sLG
NNp/oJ0NNOCm183stLBJ4m0a5KBybWsSnB2i7/6Ej31KwX/H/dFnSveOqrc9kdgo
GMz4TQJb5up1hWcGgw+V9V3lAf2NfyRK/ZubhKsDT6FqqnVS/uz6HrcZmJfzSr91
xAy6GCWzMu9iXV7q1Ksb5sxvVjJlBSgZiRAetc/xRegIzWdQLdQN75b7RSUaYMgh
vECa//dgiR1w1w8mRsaBGvptObImWmZLSMda2AZWXf8DPxVAzNU4qEru7JLMYYgt
1bLxxFndwkOFIG+MQZXOjqzED3Y9PfevJ4JiHCYXFVjBLXFvwMuvdgAiw80GNMG+
iyGnOcqQ2fka8N7GIXhcMjUhkmA3y8g5hvbvYs2WcTungo8kpFhqAixqARTnqgSw
pAk+Mcg13I0X1RDlMGbxeUxFRv0zZC76r3UHGrEeofAsHskNrsbek49Ikdbu+lcr
aE5zxzOrpyzt5kkl/zfG7V0cPQZNs/UjDNChM77CMC/eRIpoAe9KJQ1MawRBWFae
pFb8Hf4V4kMFKwAMaM5lmoSU8iy0QE5/5ey8ie89llkieYPRspM2NKTRBsfnlNfa
+1JBB1d6AdXBUlws0YWnr9RzHZ2QVUN2IEnY30wLC5iEtZQCdBNP9l7yYdeducFg
1lu7i7PoG6skn4L/tp8MB3qv8SayOcDujydJ4vWF4hVvQ/dCPetoK/66GCAuMR6l
xXs3+sp+ShPmsLzMBsDij9iDtYyOdqCxTznDlTAW0mKuY5MWa/v8Ac/RtlFBT/3E
8rSWp1MIpUHkuhpUn6VOhIJmejQUH4GQFh04xoUSTjKODTA2NZmbJbi8Rkls53aV
0KhwqwzoXUeAyY5y7nwTCO1drLdxQC/vb0iyHgYGVzGmma7I0wRJNH/RlK8y5wNl
b9Zvlgx9Vbu9L/I/lolVCqtv2ffk3rrThPdR75JcIAVwDV0mrp6HKfBVHwnSUI6K
No6yR8FifUk6Jdj4lN2m7irzYsyDFBr94xIpF4M95apKf6xPXZs2ZFQT7roGxTi5
P07YkH26Hrfy8fEY4dZzAaTBXdEAKSgZ23rXkGTX2SB8azT49TJf7OVX8+u0sPiP
oM9kVWLSAhnvFwywjH7/6jLAZgfXZ8rB8rnHvyKWUCFMyKlP+dubXlLnUjtkhJ5d
1QtXO58XxbBkaomtB42TtxMvVB4CVmmT19KuVBbAg8vps863e6N8SYKtcIfj+LvK
8xUR32igRdTFby04DOqLu7u9llmYc+m72TBJgD4mY+ZDStuNtTX/APT8JnTT8lU4
pAMlgsHCqOuLR57zs6I6+Ymofe0Xk25U6048xvAg7Ty0I/BOFBLTJiu3YPOUC7p9
yMyXBsjWfwzBkyvXk5FR0FCjXtO+HXRCf1SXdoXJvD89y/lFzbh5Am3KzTuhnZ9R
IJLCSnrddyEvMb3URDByc74rNRHuWQMUf8g7NNdFJoPJDXGLRmiqaBXQmv7ObvZs
IUvnPfD2CatsJ6aTXHlzT8Zw7btAM0ofuMblp0WrkFNMIQitTd9WbIy6eV3r4SZ2
IwVPlLqVKMkUegiZ0Z2ph5AoiTmTCOssvL3C+JSVSjtOVZWuRR2ku3U20TGPhr1P
KwUzU5esY+Tvx4CXnaWPJKEJcCEz5GI/+lxru7laOceZJefOTaj+9RIu3/ZODTBO
c6MET3nQGZG4wq5ouWqmGa9ScRs9BN/KDQHljKvIbFG19uTq3rk6g2/y1x+tLAuQ
u68idtTSu9EUKNQNu0gByxyzitmFQVxuzysJiSM5Cf5L8F2cpCAmT866vvcuqYpJ
BUL8j5BzBMc/sU+WCO0/nwakg8xqWG+wcK+awDDrxCNCAzHR7KUENSZayzgqiXNQ
ZWc+Z6/wqZaoffWi+kv/k9Lmy48SdhyC5G66+apidajj180A5zqgvSmEIgEHdOg9
S/KmkpvST6dKKVkPiPnkXfdct0VdWVEPUW/VF7IBfDQLihNf1MqUH+xUVHqH46Us
NEkaCr1adBzWGBj6be3pRS+uL2sNmopvnEqJupdld0Vx1DNVDQmQE3berpLUs3Rg
O6uU+WW1DoTbMhkO1b9YE7k1xAYKjTbPiGV5UzjYiHwUAbxubUzyQBI07z+T7wXi
+d46tgdfLZcOBvgUrNYw5nmeGLZ6Deex3nwOXf0P/zrpD8WHcYMoVBP+4mBr8UFk
jzepobo6sLDVzL6rVoJhxK0xMi3t9Cm0XmfcQlGTUNVkPxGjctIHg0hNR7HQmX7i
WC55CUK+y+bHK4u3PGY5tmv4NE1yQ+lzN8NWp22IaJgXahSH283mlBWAUZeeIzdu
KCdZNnQEkB4hxh2k7hO/1svZNh7uLl3zXq0ttaK98MF4yT8opaSEsVMZT7w9RNbB
4JMNlwi4qVH5U/4qFv1kRTEowF2jRCQ7MXAdPZiVKW6ptBdeLwEET4vQDBMaresN
xiscWHI/NOoA4Pai8dXc/BTOUKyLLNhEG9wJi7G3TEs4RMcwfnucAKld35e5xs/A
OOuqlnv47RCubc/S0gs4iTrxhBhNAzIiSHfqnQq1A9E1xHfUeH/82ZSzOFaRR9Oc
EiEIctjn8eOA3PfkICEt6eRM3xvDFAyxxYMVLwoU6pFPF7Ptwsbatb0Fe1deC3Uv
wb1AKoh8LCHR1SB7Gqrn1NsbUzstTbWGwJfAuFBd1I+/Y3RmuysSZKTQQ2x9sn9K
HxOr1PJs5+h11ptTGtbRSBViglsIVh5ejvYQTaEZVunC19hgYOkZY5V1lsVsRha+
GheRCSySkZpM8ljeBY05E2KdAK5ZQ7tiuE6SMXXi/+A9uz5pbgOo98aj/F5kMnlB
QEthfzvuVsSrqFZSpx0sr/+1kH8gk463qiovmkPrwVKd6uh3wkvqPtnbmQEsIRrj
ADuzADcVpiVjTsSZalGTjdt7JeS1x/4RR4G3Er4YRP+hs91R93pHhBng4sumP0RR
N+SPu2RdxikERYzhppAHtysKGN/QCVui77jk03Bpdz9Awwtey/pLyeP3RErksmcN
VH1LLXT+9UDfP9gKJbDqkZkrst27gS9Ela26+XumuwIM5tLh3s5aBph+J/5pwDOB
7bYUs6CFWSsW0P31v2w76TdBB8qh52vG04Vic2aFxMCi1NeMIoRffAVA6uyOVQQt
N9tlRcjGvmutjbqsN/Uy1XawaC5v3wMToArZYbxR1KHPFW7eT5gWkEZrL3tOaZzs
phL70sxQSWygaIe7RP37073RVp4q3yDGghNquVA367dmNlFdiQHkEoytRmQd4v1E
GnMGIKsOEsCtooC88ARA1wwG0Ca9FdkTSGNlzoYeRlD3Y8ePJr2SmmeCWKuhg+HF
hxMGMNfxY3ALU4nswtl32uM2bennsYzQlA4+TCZk0S6WNLxYcu0mWVTLlzhU+ngM
0OEdRAMu4qd+OL+qZajIsVku1vr5QizStT4X0kELPXXmcaz4AH1VQuZe3TfyzTEy
Lik8pDQpZ49hG8v1xeEbkjMQ5LtZcL+mB8r+t7Zcc0s/9xszyqiXdUVjZhTHWbuy
hoxzepjK5ZK8nJXmbNyZAvxq5bsH0lMGwBD3KhJGl2pyuk4ZucazXvC00T+VMsfC
uGT7xGJv8dnqk3dXzODFhW5eRK+/JDGYFLNcySJx9hwgemgWslz6Ed+13o+MZlDV
YpiWqYzreMm0l+NwG+R0k1fePejg0+PNEdZX2FoBcZo8ljo2kWnSghOh8jWZeSAQ
chcErxC8W5WTipl84WUcxt6OycRsIVWr1/umfXt7FNVcFVEKkKsuat+E1KJ5j3lI
gJuXCkxmRAz3odY3sPrJzweQJfQPGSvuUPbA/ce/68PYjN/XZ97MGxwxc2OHvMCE
lm2tf4dZ1BDmkF16lMNuTdG/wawaK5jPMct4pV1AoqYVZoefWkKDlK2fa7X95VP8
5kVqF+ObwP+cOfiGj38yliBsMGWXqh7o++yleytyHc/buOHHMGUJ4Edqkt80x8RK
Lt1pkABiq+nw3NY0A1uv09vdiY57GxZMZtod0qmphUCgtL/tqixK71l4orMzT7I6
+avYrnULR0W0Qa8ICR6jn8DIdOFtFr5DGemYAYHUXzUCCI8cL9cRVbUNi8fSQIql
YYsrljLi55VuMu+/A/YrlZViPCxxha5WcVoi8iJsYHdcrry7XFKomxi6XnaDnVix
7zI1DVypFPmx1sGlPjw3McX84sqPXEUTirzyr6Tz4CoefUrVq2OIuSxlXuP4i/VF
vpr7kTQS7ySQGroRe3TjCSoR6oPzT7ndz/dTegFGnuAJjiNwHlPuOb+/tbghhqn4
JypTVtrtFTDVfY2ODWbmwP71KD4y5xcGzQ29DTdEgTrBI7w8NCB+9py8tQqkTTeS
wCtV9VXYNYZbU9hEzC1CWt53TPmINp6cLDvy/6hTo4BzFuu+hYi2y4rTF4Ae/nAa
4G1Qx8mb6JP8DjEi+2CU3PHSP4BYPYn3Q5hMU/9cUhDBlaqZbL9wX1d4Phc7YVFj
WUIzPkAreB4a/DbVFpBhMFWWdlURLHrpvfmktnZ/cmD1HA3QurzdbiajDOSdrVv2
QIlYcNJMK5uzGmITX1aWcOwCG9aF3ZkpiKYXGz8y4B86GTIUT0NK6GeVu1C8E4Br
2bI6fhWgYf2ImPrc9v4ylfpxUtlwIfqC/86IEgkScx7ysqfm/O6Hw5dmp4hHEreX
KE8bhFxZRMafomC1VNlfIhwYT8W8EkKZYkO7DU+ynOmBQRpdyXQuSYADauWMSfwO
ve85KE5/HGNbMkCYUHPJyavikCkH2P6rqyVwAxQRehF3J7SjVJLx2wXUEJqagq5f
ZTGxBJNkU9TAifn8qrEs5X/Z/p9tRUcKgZDW0LFDmTr95BnHXPVOGU6BXuFUcgGV
AMdTrhtDSPr2b9XmRIXinLiXhEgvg93bz5lGE32/JYutujH/7rLWBmH5nG1s2w8p
9TVzi5yIw0HR3YGvKiShxZGjIXCeofj/ZKbGZJSQSjBNR6fwbC32f3AlcE2l+NMf
7xZX/K6/fw/ck+1ro+bWnEL3eplrGVHGJYAZcHaWsrFOwmqOL/Tm1yKzL1Wyg6YL
lG/zUjmQcx6EeaY8qJF5CqoHBsNp+ZbF5bI2BHUZt0MYdLXUY0jT1pMbR/kTgfdY
vd88roVDFzi5ugG+abVdqDc9S6GnZWiDcj80hukXqHGtK/r2DnxhnKLPq2ryroB9
kX80UD0EUd6dirfPcdiZT7suW0fRbzg1LKT3xIuAmecJrBxeSRaHG8xyfCZt8ZQk
3iM3iE2/70XMx4Yeh2uZd0yBry9/TM9tYU7S2CM1eNzeUgfiBhka+8RtEEVgOM2C
yKzDzsVnJWoQXTFvJt+7UkKLpxuzDiIXB59cb2v6PyxkM4+ttUj0lryS332j+DNP
MFlbe5h6o1/l+1gMokMrfbeJM1mOZkXm9l13Yg1BjxrZ6XTczhwhHqVIhllKXNXa
kLm392ilJbB73fQvW9g+CT6AmJKyCdiUD6fmo0YJC097dFgkUwtaMUcgAeesBRvb
0HtcOZKJEoOm0VGmMEHt+DyG8YIdoH3123+TQ4u59X17ROHfFlmmRjca5+4LODup
j541fmbzExltt+gsYTSs81ahj9JhbxVWNSDlY+G8046tPinBlypxdULW3xFixrvY
kou1qjrMr73MO56505Cw+buoy+3pkhkCogwpBfg8WRSXGihO4mt8w81UU2Hj8GpQ
6L6ZVm/Ru5YlZtbxak6SgOXCHlHe3ZWWZ4V9N//Ho9JyH/E3ts50OE/QkNtwSWh/
I3CL7Kz7pmTOnovBNIgiAZh4GyqdwS/UoMTDnoXVLHfhEHDXL69fLaTY/Lk70SPO
zQj1acrZlMwYP6zBmn/bHDYk08B4PkuW77AuP6Ne6YQCU8Djy3IgTrlnt1/0B4Fk
edYKMGixgZZ8yYSmlYZChUD1DeJw0FSJFYf2Bi2e0uMXqK0ZlHvQwcSGb6GWU53S
CaYufIdWJto/v002pfiji/kOWzZTpgKAaIjMZlfMOahLC2SOY2w+N45JIyIFYLps
dxnF/M1wul014SRMNTAX6+ya3BKFhT42dxuhcGuR3jiMjVfFTkMEzZw/6N9QPizH
exxxM3d9kd1M05XhOVn3T7l+4g75xR72uwo61Z6vZbGmYUTBNNLqsc3yQ5fhYh0U
oUKajVsw/E4+Z6VysxJOrFDjOXmUWKWU0jME2CSRKhGaluPwWLoaNvB2Ok4HWQYw
9zh/ytNGv3Iwf1lY7As/8Qo6yPcrV8BR3VivUrG0f/YZH9ZZ43zAIbtdokxmUiYP
sw0sA/fUL9gSnGU84jY0h26pRtqabVeann4lrLD1KYg+fwINpip36CLTdOxvAhoe
kEMeE/pMa256AT9RqyZqkT/pEcFK+1dIaZRrzvhfb9DFsIRBxPCpzHcURvURXDIu
BPynlqyKbypKIUbW3DoiAH7G5LNtVz1Tjpa6PVW2OeGrgeLincdwAY2mR+VSfZdJ
R8gNeGv1ke8pB2LKOGjqtF76ms7Ldy0WuA1t0ERhdVXbDjwPaS69YZPLoYcwCYvt
bLKrXa7BuApvV2vMJkWa7It2DZsw0nMYmEhztP2tEtZdJmLTEtFdy6JbXJfn/wsl
57/WW4JNmy5LfY7AiLs2JVeDl5YwDhDxYtBmaHD7AIpL7+xP5m4jJFrfz9K3mUAv
T+sjDQuQhOc0dAkkh0U4VFxlQWyJ72F8QTZTn/uGYOz802vfS8/q4c++BRBSQG7+
zHYAQDGg5N+qWCgdHN3hk8CMAP45d6CKjDH8KrEa7brgOP2F5G5U3jmX1E28aYq7
WL9mWV9xXxq+3OZxC/aDze45hhC9E9/j785zViM++6faf97YlLg4e7FkN2WPb0ZZ
zzzYTrLpOterRthXdHCNAvStDwXnawinBlAlnft2Ls19EJBF7bvmkH80ExZpPHcy
V/852ROvWuwF3yK+pqLKJtOJmZygW1J5rs1YXa6MQnu7//z2zyxGzg05Prit0cvw
AcgKU53bCoWIF5qFrc2ledIYb/4tdl9hYSnvIKk7ELDS9gpcpifMxSgdHsJEHwcC
5Q5xvhC27L2RVsxWSc+OkUz1mNPXb5QZar6C9iYMhz90ssvXxjEO3Jm3k+adFgq6
yh01zXCZlofhNhWaLkl7pu2XCO9uVP7IibkwLqDne7CXTYHlyo+YHuFMPN3dz5jG
36za4tjizmeTjKg7zAq9H4NlqDSxPRG43XiQA2vdGcw61+k61FVrWs73eXprkvf0
Z6o/6VaVqto5YXIbnCjFa5FfrEq5PHkaHRYvjP2O+W/ZN5YUFCegoJXgv0Ko+S0P
a2gbiFeRBbAJtTpBYNGGZd8L9Dz+PuE+uM3vOikM4r/Hm2MaMPT7G6UIRhQgJvlF
gqoRzIO6L0d5tEQOw86oQ99DEsOZ9npFxWiIjVvW0MgPAhIFhaVprVcxr1Xm6vBe
Tfs73tZwRAGMkHBbeMErLVJzw24Qi9LB9ePA6dNKRSgM2wQ+ifwtzNHqt6CmtvSG
T0gvOhSnHc3cRErSrJe5BEB5o4dCquaKDwfpTcNLqxHNwzmMjSzVzOdlsnHqy27J
h8Jh52KPTODsRi19++7PHlJsssG8nnNwcGpJCzq8kcxfjGojgqMFsesLgt+x5w7q
6tC+Y3PIGmIH98m5SccALt8KKt6AgF7H+07i/KR9fXmG/GxCUZChFRMUwvqbX7Nu
r0GZxXPgY7A5tkbOv6iNe45GxK+61ZiV3cP62G/+NB73k66ISwTHpEXCHyfMf5DC
XXbzl5RwnPT24vIPrLOu4Z63kmKV0jz/budfcWsZv4zs/CXcD0T9FTBRQgCyXeh/
stdVoVNf0D/srV/I7xIUkJsZ7wT6Vw1ev4hKjnfprrQtlXjTnuQpx8x1xRqU2SJf
IfGUZnViyqzUe3S4HTkDZFzoCLMcE7qBXAr55sHHIWzwtvLGZJRCEGjdXv2wuW7u
UYBBuePwhJ/LhTH9zMxKkFPKou52dA+FlOqjkp7kJ3rHx9bCbX/KZVficKkzlgL5
iWTOuUnulJd8bjNgUB2Z6P7GMbGhYlpa7zoaG+mrKloaace957hqY2omjFYOoiOA
g3ndc7liTfk6lPQ1/BoCMh7mD2TJoJkcVzpvuqQUnEmbdCWwYnFdyuoPzTUZjkSF
6Vd8zTE1O/BkUU/fiSvJVnzFZeaHqg5sKK7z1bjwG3KJ6QejAtUDOG6p+PDoxNu0
2Q+7yzqr0NjfcDgmZ32MEGOeBu1lX56Ls4tMi1OcKT2Z+V4AbQ9LSqD+Cyhvhsq/
a1ZENwu9+JKpfEkElNuJFZSf6fmaWHjbWinGy5ZYSjwOwGB+WoFoko6i5vqjOZ9D
oLEP8grJTa6iYvaikpbZaC4uSdj5jX5tVImgFCFNJQWuIoknr7hUBGgjYpgxX4Sr
gIpcgDR0k/UC3NM+WkOVpGI+ngxisc+Upr74fUuHKc2Eq0MdbV+ihQTQizHxkb8w
Q50OZ5i1LYZC4exGLfjZ8yHPUEh9lVZ78RHsNhPbniDOwv7EvfLQRRW9zJcGDsep
CcVe+oY+ztHQafZQAB0tIv/3iwmlbVvQEldPnl2zdO99hS2bjqVtUiwmZ9vskQrU
E6+wXtE13/LGtpF0aoaJm1L8nyowht0H3pXbkwEYxCCBlh4TckvgFDOD80UDJIB/
vgWXSgfgVYLsnKqsA84vYxGIIgj6WjFT5diARwqsgo/NfQJ4eHDCI+hldXgeCT1z
QUwA3xgTKFT1wMMSNk4ZikSv0Vig7+ioSqwo74wyXiyyahIa+2ezJ/ggk9nWj3Lu
VJux8jpvg8P3B3gHvdX50W14x3zt8rtqbJXxy3mBRPIkk8puWLJ6oPsdAa4xNz9Q
R5wkFuRgbMgLqghOPwAmSJXqBPuqPHUaHo9jgjGBRThom9HfvZjR0j6qMfu6Z1vm
alOPCfnW56v77Nl+9j6jSlUk4o/4cMcimkOhAlHXHvgYn2nosHQT/6hoVonbkAZz
UmWKCaPHWCgEdskVOxIBTOWpHfoNDsjJrdzSnpILomE4Gw/zUikgHnhDjowuRpg4
UUNtmWpyjLa09k1VSwsseFEP+sSS1h8bpA4v2iwMuSp8Qtk2i/+GssOu+SvTg75h
wvJr3ueKTLHE3gGGkmBmTlRMLPCWFcL1xjdqtfHKzy3XsDyQFeXCV3IbARqwodW1
o2d7Ak+tO8dxDd5/51IiRR3pDnicb2PUMFb06T5SwnQYbGyUZ2tzZMjFShJrEKn1
UqR6Fdbu0shaagwVPJiSukCaJBd+CpLa5rZsatVXUbTZyPSzXMBDWKLaEYIyzeyh
R1u68WX/qo7r5DforPajuGkKdIMzg1NwLOok2HaO6Y4efdcMci/nIGhw7a2JVIK7
tU3fOuuZUMKCXK134M3cpsbRB1AcrMvMQOGs6iAnb26KRUe34u94ByvRHjN8yI2e
ujL+b/uo5Ubz36iS03RI4Ew58Byu/Ioc1SYxmk9V+6mLKit6KXMofIYDTGj5IwJD
pKfa1EDNMdlB9Uhd6qh/wvXDLdukcE4+Adbk7oSd04ZR7wLSg01UpyjkI0XglUxA
cL4CycpR+adZw662wOY4fhFruleLlWXZD7GuiEDsMrm81zz1ULHuTNmfhl4kKrBx
RDX30ZuJpcVo6Ui30b7PD+uaGtuRV0UCyMtNJI/eLQdAKIv/djLT/2XzZ30PU7TW
Pt0z0bh9ZqtAXf6egehM83Us+FAXufHfHCBp4NiDRK8EbuGt4SDbc961bawhE5+k
thBHJBJy4m0AHGHDDHL0UBbiuStzDNFyHTdQRCDoPxDrhlT4ARyC/lz/0UJVJrCZ
7SAusK46giRo6fJVKXvPMjBHpmWhFUorUPYD/8AOlqHRd4DpOmBGmz4wGPf8iAmx
h+4mWtagzhs1YoTkXGcA3I+Q1OcFLJkzMjs0vdDtmFKipcNb61m+5miXdjgb9ccZ
HScCQIAotyXibUppVAH1vPK0AoxWvuxNP4kuSgxmlRZjp863nw3tBu4H1CX8L2/w
B1OD9UMpYUVrpISoQqJmpbcgBX3ZDA05PO4igAlN5BlTJbb+EsuyiDbEjHsuwWny
b8C3YqCM1AcKjLgjD24Z81rnimgndpF2kmEILd6i1QbZ+YIIn2B6tHIm8QkHetYE
NzcK9dgSAvuNzGoXBnXmXUgPRmjjVAPYIHFx/g4AZ2Ly2xRgZ3XcwL8Wqfv6QjQT
mExU0633xQM3oY//89Vz/bnQoey+USmhTGZ8p2FLhDkz8/qQVicl5ftk1oPL+dnI
pFwrxUAMEKGh8uB0BVkS00k0N8c7O04s99i4DjjJ5JibOI8uEi3NZ9Pe1mGPCn/S
8Gv9LgbRugC5Q8x+WdhIHCY4gvDEkltggXNj99zBmEzXJRuZokMU+0nqtQPXVx8U
dZ75vTnNyxLQgn0bUxOeYvnuD48lWPOdtGZP8yNwHtdWDDf+r2+5nYrq2CONDzBm
0mE8jL7/IKrSqwA7pdfGJj8vRHUjTFDlBf6sgKlrHpdj8it/bp05ieGUAYFSPC5B
lO1gOE0yZxUmm8Gjg2WJcZoO0noS+w+f//KnK/0n82rYWu2z1d8N6Rdg7QP789e4
MfFlOAlO2W1/gh33Ls40Sr6FGzK0FnhifiHIfe3Vu3TOM3rkUJ22F2N/7wIM4HIa
rMLizK2ETU7260Wps55qR6ViOJ126Y539vI3JCJkG17BhNX+x132tEpdmT/C7fgQ
dA7t/NNYWLQcjoKYEd9SEzG2IQ54AwJ9jHZshm7B3OVnnF6pD8NnTBMbprFvZwnu
sLGJFBDsqb4Gcvl78MuY4AAlz5Sa8OZUFlIlHZu8STX2FL+p+s+REHHsKqJgeyyL
7FVObh7GLbqIPWcFR/01vwHvXvEiOmysllqRS/K9/XUksrI7HLRs8h8nmxPnecpG
4XTC6HimvpEwft+/uAnynRvOAqUC9ED2/DIyGs3GTWHylNaR7xFOryxlX8qo9+d0
AL7S5/XMmhM8YelNBIPkrfX62rNpWC0ioKLNqo9/g9ZeVlMdYBPT5tQqBsaCwiXp
TLK+hy46+fwIPXy10h9MxpSjxN/832TOiOhbliZNgJkpqYZhyextGYB8jCpu8pPx
//ycclIxzpTJTEDTyA7tNGEV4OvOB5Gb60B9OL6AzZ7Fp0VAFGyWSyQSouGFaVYg
rFwQKPRHDekGXSJiunMsK+AOxDaf5+/GXNtnlGFd6qP1LhnrN9+WVcHNdGNE8V5l
okQg+J8QuEzOWww/wei0UkTEVYFCGmFSVOyB127wLgVSjmr4VN4wxwzDIEVN6pbf
0IjZ0tIOhRACsQm6+gkBvSzhXfkjYeh35Z5eajfogw2vYxcaaCG0BkfO/ed2D8Ov
mF+7CWuIwdHILOW61LRPatpsnNp8rI1VtyQcKWfe7pCwpoJIPVqcprWzRqi4v4qX
utNU1S65x6ti81WcEFnDxhyRJtb5y0h13mALCxVdLDghHzREfm7z+wz7oB1u8/SN
TcFaeJwbXWWUr01TBUnEpNNNH0KUvmqJ8avnvapM0rRhW4khvyOdct04nDgGzLXh
a6OO5axGCpOeUwmp8TCxNPgA03tMD5zu/31Z2dNhnaE2xW9Qy8fkj7T2hmcHYvWX
mUzK0Kh9F4SuD9eNW83AgTJeeCAovQkYZbgF5hytA8Es7IQng3dzwNDx97M10+NP
KvdJaTbuXSsXHE0MKb30uFoDSRBvsUyM6Y18z1otS3gOVoflOm5Qyey7je7uFssD
Krat6fUd8KrYVAXkV6DpvYP9ncy46H9EjRM+KTIwGGAtoi/4EzbErNDafTQ/V7TM
ixNB4WZPK457cxZqHgWpA2dq2MlZF8L9OTqmg3sgjVPSz2AaywIOR6gJ9olLwdwH
+/Jnmw6VtP1Tesn1Wh0ssMelU9SnEReknJwKclD38ifDwT/Bkjg6JmbLVcZJBprI
BZYstN9k/tQ1TwSFghHanIvyG+jc9Pb9rlt5UnJFtw3cRZzd1WSiZPe/umi2RhSg
LdJy5mGj9FrVyY8Sai/3ChfWELUdswc7kimtVb5AnCtdlyQnnXs8ic+6Z5J7RIIy
vddtVytjq51dUYmYkdaaHEWSLDnpkbE8llbozaV0+0FinHzICle2LdTQufPzpLxb
PPWl+oNNDmCC+QE0w9MvnNKYFzlIyobGYTj8ZVXBLev0BNcWnx5KsRm9ii5g7xD0
lothes+V38oSAf40VeSo0Ipkz9FeM6KBBuapjMiK4QN8tdKH1eU6PepVi58TNrGV
YV+4C0x9Q7nniAyiMOv57kuSgaA1LzPPKRJPLypY2jrwr95ykKck/e02RnM30K5O
wVI/swajBXnuVDnYO5HpZmz6KDR5FoVJ1xV2+PGdtlWLNR7s3PuZ7++WC+CbIGrB
5ltqIgVCDMMl8k4yEdPYsLDbj6tfQBHZzEUTLd+kr4SBTTrC2RhZUrzRPGCFwd5T
OACtIXIbOdZDSYQAx4H0MBw1IlpiFI57E7j+bzGSZbp0BQJ9VetovqkuVhPt3y1W
mXcsFizxCbB52dxYO2okY3WKROHii0v4OLrbjcosKXE/kSSBj//0NEDyyVa/oHbc
bzfjNV9wr2JNgBeoGeNcs0vyi3mdWmLeQWh1EMMKSz06Qj8QlXVOMXuWX1nzuXZF
XTqMxLyD56jPDoQ+0Fzcx6VlfmILzMlZs1/4CGRWreO+NaA6400fnvKlwJuzXTyg
DwDxjBvdbKrl8JbatjvvedvkWpbAZx7cWp37iq9eOYWM+TZeBvDG794mkrh2Kue4
l0rzv3bMaBqh9aP2syJIBWvW3XB2VyI5nmrUbdaadafvxh52O4k4kJ33m1gJoO7t
p5B3h64svr20iBzQ3Qxjw0kvY9lJK6tQ2MInD6hAfKjweIdbcRxr3KC6/fXNyQOV
QWUrkBEf2GufGurgrBlMHYZh+Qji3kFBijiAJKpFf3g8QJBuXdVQlogLxkkF5yFf
YkQtop2/b5dKTf1uJ+SkrjmBIolNr0LDsZzMMC+hv5KqijE3+Ku0iVhUYfouDake
FCQU1LVxkWReVyP5zDXiQfeOH+H92mO0nY7x9ePTJwwNK5Hb2TJcg7L1rg6uWCnk
SH+lFaQrkd/RwD6iMAZhm60J+rZLj7auTcYEpwo+lcFhOftJiT8Xh38hTdB2Bl10
4oBcQQ6RczQ1AyLQq0roNOcb94DECCahg8Os9bSEWXsKgzZ8ZbgKAxdjGLL4nact
GSCRrBZe3OIZduRQBmWl60ttH/z09/8f9N5rLxZ4ZalNes0PjVdIpWK72o65wQ7E
G8xCrUCE0aSmVyED7/rpo1uD7kSjBcfq9l390Ai2g5FBI9RqGJqBs6bdVoDYvIJj
8B1gavDjScr75EegVvzm6CzqwduzT28Oe1fLhaXMET569soJG8o7ILG0WMtb49Ed
OwXB/nSJCBJXQ3yFwQn2vocSZrBvC2ck+WQ0gyY4CQviexb9xh+Vxh0z4iz11Hd1
BJ2F1Ogr7ILhGyY6O0FjUWtplfAjbgw80sE8WRPG+RGnrz3FFAvs9OdCtcL17pfl
7qi6v5gYcsAXh4yv8kkIbg7HHdFFWHc/oBeYjyH82mau1hDebjTEFwx//mYJwII7
7F/4RdBz9le9KX/Wi+OEgMW9ViGh/twXAFa7sFXQuPCHMTnZOaiuxmzvMkMc/c/P
6Ed4VwMsKD2RBSU4ueS8Vg+5aexlb5NADH6zz3ELAacsBeFCRBsMbBjeeJw68KBq
xqIM9Aea6nthsffvhnbXVYV0r3uMHTiioffz+l8qFCokhf9hboOmeuawCqQ5n5lZ
XpPw1Ljk6kO32SA5O0n+uIF+9fxkOpmh62VKtv+uEqNGAk7JjIPGJ5vn+SW4ff7G
msV+yIwFcWlPubrHS1mQF5ffhEjGX5zVsglc3eCWO1z+ZvEIQZIof8aFs74IzYk0
zX4xUs74xLVSCrnME/LW7iqoLb5bCVZEu4gx41bH0YWoeGdBUJOJZaCu8QGUSKpA
/4R6wpuYzR/OXH14gtLJPJhF+B2RZYGN7KV56M5VNcBOapiz51lwHIHCDzkPK1IN
s/3gVnaMOnK9AWALbhCklfyUCk6ukrFnJyZotzzPHERIKC0ICTIBJuv7Z+O3Rvti
H3w7iM041ncpKxk2ogL5DrWouU9t/EZfF990afHG0gPcXQBmA+dghNJOx8nc75M/
oboaB3MzUVoMguRt9CvkcmAxj3Mds8kA4w/f+137J6tuczn029sjA+5uFthfJb2S
n7sgT69KXXuMTS6samC9/h4MY9nR22l9BKnRfQHjUh/a6VOeUh02S5v84W0XaFTr
DSlleF1OCgVGSR3yeMUWNP0LZhJ4DoCwbXHeXjjufXyclTCeYEf7mUX98mUwSli4
VvfKlpTVPm8ekNUXh1VzeFHtyd25rKx2LvbdXutHq9Xb5rIhRPAYtVM3S2IxdL0u
ttek4P8lWSNbs+9iLEurg5Fjh87zJNikKvvrsy89tB+mVML9jQW8YBPK+BOAFysz
IaedW9HCxqQJgqKYy2+Y+5IfvJWBXTP7OHFX6AxUiWtkUP1NpZV+AFseTVB+MPMN
wpw5OdqVnaQVlapurKal/vanKx04P5SV8a0Nr6fOGI15kL5xseCgXDec9a1NY8br
BGgYfzcGNt7Gg4ZqkKTzGgjmtQny5oC+WO9S1IuGArkD5GSOTCZwStHqn4Erx5Vv
Dr1nvc6U9pH3LmRx+EdCbSWO24zTS6jOrffDOfkSbCuTX+rBirKpFepd/i4dgUAB
stYFRmEWO5/DUxYICaOGHac307tL3maC6nV7YXHpE8BPTrUJRrBw/UWPfGW/0mWX
4rCd/gtu+zuJcwaobLbz4e64sFhEXB5Ku09AeFBf45eplrN5G54RFhQB5JsReVTI
2QKKR7IVEtGs/os6Az6Sj4GLkUxFvt0c6+7fBrsncO07m1ukerFEaweiZUfPb18T
fkyRDvK02lOxXRROLT1NLzZmuPjcQVEGuK0tCBX/c/jJc3E2gK5ugKatA9MaTxWB
Yc1qZOYjxpXdeeHoutv0b1uy0clGm79NX+Ol6vodFESdU/oSM4RDsS5OfhDk0/e7
7ROoA8JmV7lxsY4/3rPTtJ4XaCUWh5vjpsQAEGtO2l+PDJ0mEZN71DZ5fcFPvwYI
14KvtZZ95w5GhyIzIx+rCaEh7242nR8VD+UKlNQN5W3BVQguWfaltqbAXcYD5+D+
VDLDaXa9XkWxR7tWoFJV/O9Ffr2cLzVEI32wO3A3qjIAUmLv3lofZDlBWoHUnJdd
Fj26gc8jgplyHuV4voayx85MnsfRREP7bsWTBPbIpeK89lhO3j/V0Opz9k7QROJq
ySTldsp6DPbEuUStLQ1pSfkyhzyAkEqe5b2cSO2UMnqodEz05m9L1QYCezUt+QUD
MyeAtXRmbYboLmPG2ZeNAyRFlIv5bIjjVvaxdUULSROrvRZV5UBheRYUyd7rlsvC
pU+1Ta8zefifdWQFjcBm61EQyfdzXru54aCqjVeWcdJiIqH+7LAuylMVHpmXStEN
/wn2G+kuZ8WKM3KvKi3EokL9Qrq6DVitqSE7ydOHSpE1sV+Todq3LmGhZpRkv+Zc
KlfFvaRZTa/QXEEjh5XWkMYZ3jd31HUqVV/QWbL8XJMPMd+o1ZttRyjrMKHD2jlP
r+kB1JQes5Y7KOiO3C0CLAZF0EH3JnwqU4og1+rtGQ78GfBDxlPY60genfpDbkGc
MZ4+VrmQhNeaHwtIPJ1ekWP2xadlOjVbllOz8rJveH885kJkfOU/TyNA9hIj7SXC
WdW2NoRCjTenU/EugfqvSpZnVSr3ron8Rp19EU0lan5FpI87BGlGq68CAMFke75O
rpib/L4izABRPN+OBg3X5+IlfOIVHiUX7V2G106AaRzqz3S00iDcmQTUwWfTk/dj
w/l7p7CTxpGMJpkDO/7rkia7DpPDpRDIKIssDDalJUiXCWDJXpdN0fmlb14mljia
VznlOA/xIX9nR1jXVHQQw/pkf3iRRZYC6Yf7L/tK7ariziZexLI2W1vbbm2IxA97
XGifcWVDbagasLvmOH15V03jZy13k+sCdguLqU7XKtWjP81ERTcCBKCvWWQU3TFj
oMe4+lugK2PYmqXHY8/xYuUEHihYl/U/SGO/QVw8wDTjH9TYp+xGQ01vXLHZjaMZ
gRAG/5z1npbO3cg0yhPiCShl1H9NKCuPQIAzvp1X5miyj97wOgqQRrkXi+hN1ato
WE3qtVjACA67gSa0fQz11w6oQP2kZPCc49dMo1lDFzxe8mkhfgYt7grP20V0CJ8j
KwzbXwQktLTqm6cupY3bUxkSh/8s4/pyJWWciNfmJPjtBkVQTYg0KstRsjn3cFTf
TEI4y7yLL0URGqbVvUHtPIuKZQ9pSFmYpqjBaexD8WEPa4nRpP/EdBNLvbnxtJOV
mleFvGy79jczEHpTrXvdv3+dSYojd/Kq8aCVqkuSNy0YYG5IN9ZYeLETaFFAqqRn
nMrq9Zb1kp+OvuYE2YgjOLAHx3sJf884be7srXbqFafgY+tS73F+XeMLw6G0suIQ
XHFv1ojl5tgPhnGYseYx+AbESH/bU5OG90P8/kIfr0c1fnYAyagvqZrZnv22cWoy
oPwWcA/zWHzzGBCb6FsUUfqNpujR2qb4ixYCTlJLdp6Ka0nIkBQQWWSK6ePq85ll
LlOTKeTT3FoqXkctWdc3EoeTLq1C8jRGLpTmIv4ozzBOdaUfua0WJHDVyZf0snST
HlEp7AwkJzcaxr6MZWtBpRosxuxGWZk9/kQla6DwhiplbdU2A3Z6feJZ7PiMe6tt
d8NEQLn6PY4KE/3lbfp1OQFEGNc/E3mJebchmD5J3OCZFF5T/ckuKqg4qAqnn1Gg
iDqUIpeISPXOAFLwqzgtTsPfp9AT+XO0wEkaWTS2KDkFxphBILV+KOVfal0kzIlp
7x/SOD77gINRdyvHZc5phQQmUEqbc5498xzdRf/O/mDnRiHnijv7G9jVs7SUbtvM
xHGNDN34IZO0xuaYfUqcCHKWu69GGSrfgSEYSNvkD3hhvCEZPhoYNGfBJAj+EflC
/zXa21XM+jg1Ka+a4mnpLYLzlDj/1E5hO+qVcOAMz5PEQV183JZRdVBIL8KFfNHH
7GmJ3i2vqsrwmrOn0B7Ig9iLru5IPstYytEMu1PvxY7u6ob91DzncJk6aJxQolZ8
T0mTib2lCHxq41d3/WvHPAqbto3rQRIgiAq0jab1bu6+Rx7RLDAd5b6kLS8eUbJQ
wveStr2f9wu7hz5GQN94zkuOdHE/bf2NJp8V4Sro2lVK9h5uc5MOBRGlLO5TJR3w
u4aLGA7gmXiGUVokHBGMHmae6W3YhRnXV3p+1LFBVVFO7ikVccwR8Bt/pOFJfCA+
micNY5oqXJCr7WEEuKtsXpRtHLu1QCMwM+lthVT3NgQROY2MhtDxUt/eAuS144Bh
DMReWJ+bV497tIlnmdC0ZNkLmH3EfIa2vAAy6e0SzvngpSGncv61839/e/i72uwN
rIJ1sOVIcSnT/W7ZvkQ3fHUaunTOng0gGh1+c6RoLVbNa85BDPAM7HM6qROe4aNX
uNBY4S8KgUOcB3O0FZZcbt0MjG7n2Ao32ZrVxpazdU8BTCxEXsCtb3rYr/kR2Ae6
LRY53IBFnfffci2aDCLstxcwq7qEXKFRLBBqYuUDBJApiRaeez5rmvq05tsRFW28
hu2+H1tyX3er7asknLXOcxeUvIqs+3Xshxi20YD9Oc0qbKAVjrX4QaTjJV/O1Q11
aF6R31A5S6nT4XjDtxrE8I3579XTlgDjT/zvL/cDZtygs4CDkfcNeAbG3jAPVUUZ
oHepTA52JzyD1C+QOl1fpeVv6ddEMPb+fjNybJrxHshZKX/TIaj6dXhlY7N4f4Di
sHyYaLNr1v9VH8XXpfWTwxk1x12lefs31qQcqL1e2Gdlf9CT4HVoTIpiJPadJBjn
h7VfGKpYRpxAhf6h9JD8kxi6dcXVXRgSzL064FPnnn0NKgH/YX1NqfFODpkeuaaN
91Q/3zIppSoa1w4LMSH8LX4H0JgNcU6P3V3bF8X96Yb2Uu55vS47N3s50A9+GQLI
H9Hk4u3kMmaFw/CicxO1bg7Ws3dhRDJ5vqQWTFjRyZXOYUVnVsbk4P7iZmfb/2uh
eN5kuEkNdwWKKE++Ch8ydQnj9BChbNnceUSV6b4FIebWedn0+JBDlloElAr4m4us
g6smIoUPjyJiQy959AtlUrDwJ1Tp+3Pxspy8Iu/F73jRXdr9K9KF3Q4xTqG4dbqR
eA9sXwHPo00r2OWlVp9RqSABmZFVhxGZOyDEL0Ltf7GDEOqKMweTyiAhwo7DfSKC
e0amkk0nQbKVrAx2p2ABtiVVy8DjHUmZ8/jqk9pwwgPIAZVnMhwP2opCsXlHQLMX
PLwixDtGzZoz++dVjSo7yFfZrNKchWeY8cR6hJj/AmKeaAq5XH9GhAJPZ20BvPy1
Ipsicq36d5VySZUj0DsOi9gdVntDSrasF3SRzW8nlq4PZHEps44wHItF51Ef4/Gl
2bZdtybUOjQ43AQa1g8vzcpjIoXgi8+YDVEPDryegbnP7OqeDKinjGw9U23x1vUX
5QJqBRU+f8bnhTCQgEYKUJj0z+JhIx3iMc0eUKVwp/ajdXDUHbcLL23fgznLGFNT
PdeZigbcOAut54nfNBh9ON8idt6zchg0qaxRuNfAvWCp2VMnRQTkEwotzbRzrMS5
Jmnh+EH2Zp2EZ70R6YDn2niZLifONHZAEeYCIPBDYcNSf+D/4otDtwt3H3lpEcWz
UH7aHjoW6P/FLgFw8WcRgxlWsHYp2dFuO+lsf80Oe4nsPgc/sU81WB01YjBiNrQx
PNpBXzX/bdKfDQcjlxR48bRRUChIqMP3CDQC3VIr6Kw/1T9SAGlbE3qeo+IaGQnH
l5nSs4AQnrdw/LyIRtTUjBD1VV/1IDbRDBeSJqIb26iQScErlz+Vl8p7vy+hXm2D
oXS1kzuT04AyxknGFhYiE5IFkEh+8JQDBknRsCigmvn4uWod0rveOJ+9lQT3S3Vh
oNZywaeFTq5k4nReS+vJIhWxkLoEkfAUYy3EEI5SVibe7tKEH1/AVbnfnKi8Q2C6
V7vq0iPsvSjsvDn4eFjWRBPgifrvwGN75z6JNhMiQGHAwcz+Pffkd5yAA7bDDNea
NUa7Kog9cJeKEDfm4oN8AiZZimTAzZ3XueKba6Dn1FOuqXhPPIBQ7/BUqEBp3EPs
M3ehZN11t1UDe+RU0DCll+J4l3Fy0QTfCP4C1QyfAgItTh4oFdCUEgKTHkrWoj1N
C2uuhvPShU0RGlhIXvhcPLHn/FCDv+yd9zY/Dqu2h4cDi5AUvi5PwFTQXg8JUO/a
zpJm/yV8xeBPph0Rn5ajYLvV6CjOfvRE9mXFFQ56eXQfQQtm7nKrBTErjD2+N8yJ
KDFgbIqj4Ntc/wTse5gyLHwdRCaWGbdJ8eQ7Yav3Vgy5HgCAC0FOpIkyI39tSH0M
IX8uNcmk8sM61qhn8t3SDqd5+hfmN3wZPiJbdrc85cZW6gLK4X6T1AweZnrT4yck
I3zF7j142xoHCZ3QfARXTasFoSyNUTgSn3tLwinecUpms/SuXzVY264+bygLtuSg
DyFYDyHrOidmNADehiYVGIzLzXdO6vg9IVLVZsfnFv3KMoBE2fqe8t0+xJSPSutn
RH83tLhbq1qs1wmSzLaF07ZE20U5mh98uyOm/HgkLXavMr92eIVUsJTd+PJuoHRN
VqIbm6bivqyYoCdSfFTDkV9za4HD6+sEo7gWTrXFsWV67NmelJYHNFooSVj7bK2T
0UlSi3nKrdHNyGY6NHI9M059MKGZhiHeOohb5uDHNZnwgsdN2vh39OGvo7t4XMpC
/wBh49NbmLDwr53+Cqjow+nsE+wo4m0zkQF7cVzIDeAiRlEq1ZIl4zrwuFWzaXrC
9FUPDXJSLPWa0UF/Ble2SCzugq4mqm0qzvFQrOjlv29UeTHZbilAHL3SykUGLI8L
2MltoqmZPEBeHJVHa/g5U5rFuMDWNdFQBjS9Khge3xZXvReS9OpafkD5I/j6fZmf
g5LTC/TgYS/pmCb+UXIjufj4GUdOfPmHo1k9eZuvSeoB8YW8aznffu6ACb3HtQ7K
RUPacuZOW+Hc3tHFnUip7pBhuRopxaIHcO8ei599HpXZnUWjSBfqWLV1F3j+Fwh0
RcbUOIMBvlmS9qiiQOlxx7TXh36U8PuFpyxOOYYQ4L4AKj/y07bKonfz/HTtqlMv
9TlEPxysZrS7hecs6TUMw31ZAkjdPGkbgP3raDBDN7PPmJlZ24y1HB9isNBzgO0o
u/sTwDyGGI5eVMtJWBQuqP9B0ZaOCj+PjwCrfgT0sw/oXsJer6++TJqtRrYHpyCh
/VSo889Fc4E7XmDFjn8SDGNPMYziZ8/zdX3LEIzZBKh8NuXpiDQsPe6lO9OqhrLw
Rkt1+uA2pqLpsxuJr6xIE6lfyY05pX+E7KMMo/d9ZGdYdtKpReONxZY0GoBk4CN0
JCc1WgLfIG6sZz8Ua9YJo4B+gK2BZD6jLZjn2myXxdCy1pAF8QznC3dmk2ovbIrr
/qhwK78IX6GaSTVpMB4iFQAg2CGurwyynB+F+ZiSudEuBkrz5UwuqWbsNLKKOy8s
3sJJ9mmDjElsQ1kG2eVBbMB+AHS2qVE8AGnOmrNYAZI++M/tmuKe/GA7ckBlApeo
GRGB58sti4MkdVZ0qg/JkVI4WGFLquZi3P32fN1ImvV5eerP79ZU2Zea1fXjJO/3
ZN+UT2MyTPrMNYnk2Jsjiqr8qlHH2im1IIIoKpzmlIHmrgRrVAAraWboaP/Wxnke
LeQ4jPofzIYd2ens6kfBpH08d8t8dI4eadhu5VKmPNc3gMB+FH7VJq/ZR9XFDvVx
n06z7nDDWI6x5hGn2CnasbclMaAQPO8QKtV2rPWvImXO5KXjILaWtAHzFr1o5Vd5
Q4+XUTKYd3QoSmKkzxOqowPEJo4PPmfr//M9xh5V8YxtcCsJCXo8zclcqmCL5wmh
09xt/GgZY+SAVb1FS/RFZxZVA+kGWVZYIaJUFK9Aq3xgmx117fcxl+XNCp+pVpTs
d1gFw52zvWerop2rYBaazN5kV2MvjDf/yp9tMw82h6nfPhdwTbIoJPV0WJuj5dSa
tHApxilb8jmVA/wNQmT1uA4NeQv4jORjgneqeJDxvc9vomrnHhX7fSaLhHURWl68
OuC+DoXFE+IBPoCMwijh1PLy+4lMRHVOETXrFTuvPjIuRobEUmBJvwUlOXySgd1x
J8Vt050jQ080PfIVNJcJ1d1RHkOhF7XiSYFNA+BC1w2fSZi4z9c5wIhA/BFGPpeP
Ozy3g+dlu4K7i5YraFTZWNfEC7nbZuiNdApaYjrmKMZu4uoB6YVVr+ajRRIM4+A5
SAw8romuO3p0RQVJMcR74EamSDKlit9lZeekPeqaz8hr/Ge8GtACilK1ciYH9CoX
fCAcnJRCGbstRZSRYpM24dLMWqUbyiD7Jd8gnpzSs5GNnorlt0fxTZCUtrkNDNhp
dbmXtVN9qEYIxr1SKJYWG58cwqfj2gOpktQ92TsMtN02/KNCtdOajXQi50do4J6L
bTbHJBq0sIbNIVjldo2BDW+2AgapbvcqEmQ90oLvJZ+fq4pdN3/ydN+oUcoZ8QC1
JM/jbtnMQIEASnW/2UeEvbBBHg/AmLjyVcQhBW9j85NBFIZ70MmeHsQJeKDEJwna
CGXQZtKvTSbaE+G5k201SoQS5//3Mca371ebQKwokInB14pMMQMNBCriSh7N53eF
1pC2eFbk171y7B+Pz1eFVp7ztNlLi1kauAPkocRMsIWIw3hhLDdJkUvfPNg9bGXm
bd9Kw7aWLfrJkj08bQGL88w9sk6mMcNTRMLQrP0uk1m+AnJsoF1sIzT5XM0z7fvI
Se7Y6rjgIUoowM8lREMJqiA6zKvfdeGHlbaNwAX5KLgIttWuZBGlhlmfiMIVbVFy
lcQU+z0GrNzsoy5LR/75y2JHtsSTYlO+043W8JEFhy6ViWqkoYUaMXQ8E2d5kX87
43lHqu3apVdeVuDeV4CSkh9INzgOeI2XKaQ7IG5M/HQXMJzPwxF+loM4ayprhLnG
unGTpJGECYlWMYaBPn03l9wS6OxLsRv56jCfHDimheGRxZfXSqcDRQW2FIA3D0bE
TcS5cKPODV6lkmnkaf95U5BdJmIxfdr7jhSQHTKdA68aHrTq6u6CEYhSOBaER1J2
fivZtaMMHr597C5p30QquJ8QQK2znJN+6dP0GrDpdA91EpTG5TWo0MhpHSl7aRra
An1tPrxzePqp48bovmClhX5I+z6+GN75UCeUrzjxfcUudyev9PaAVhdFgdmaMlb3
prb+7K9xyOYkzO0SXMKendCTGD7PWx0dQzU7AF5bGDbYxTeZf37RzDjEl/PY3HlQ
VIouAZRv0/uZyczXrnhJnNAiPZUphZMYEuzVuj4XsS/hRVqe02Y/AC7gmWe4C1ez
qkE7yw0+5ZKkLciZzIYwL1JX75xqbEYpjsarCxR7b8d/iAwJAWiVhb5b3k9v5OfZ
O+JvH95m3182CjqVSzLDHqezKCUPcQTj7s77FxwjbSsVXS4dqjTEdq+8I4M1Isce
YkUIO4oOotJEKmMkPkOU5x052oQAiEl+V/rHRf5FRHPeaBweFDlJpjkJqu7Xqp53
EIIY2Z2FDd8z07rxJ+WuoVZ8Pm8QpxIE856pHAFKr9Ka9EUvjDwbLQwxgEbTO7a+
zeRaaz8KSW+LwZjYqAPs4pCtvGjAM+qwdJnvmkuJNV3r/B64EZDKp1vuq4X09dCQ
Ugw/Or8xQdVcVAOL84LsPGa6FsXoLLT3V0qfaFxpyA1hSdGMu7t/4/nVU/hI5laN
Z5GyFlDL+4HCQT0hYcSzhNs4BV9GMCIlaXuUGF8qzLVomEhxqx9EyomUBG5GhLJl
yZhY7ls7Y0rx04Qk6ePm7KOumtpymAAsQMd1GhXuLYiDsbmhr8uIdn5uKjA1m9ox
ZKn0TH/i6I6mmbituL1MoUdj7z5fcfbOSD8W/24/dkrbHwErxHxBVhBRBLDQnJFw
98cHBtYZ4TIKe4zuCpzzqDLqUS9Z3RelAqlrv/VxVk/5uucQkoyCSLVeAVbBe+/g
bffLAs1RZai7Me+3/QVeF+T5v8ax7cF5ePwVpRK0bkmb4qJZeZ+D0QUrWHtU+L/t
0qTouZ5XUhj6aP1Tk+Lg7GGf7UEk+14P8GK61D+kfAZoT0Xh7MayZN+IQ4r7oKDi
92vi958vIEUKA96tRS++6aod3uvMczFsQ10cd+moJ3+1JOAFwAOY2xqMo4uOJ2YI
DUwhTcfHXo8Jof375VuWpD4vvPrTe+dpmfQdchhgCX2qmKXIjjAXWOk7ds8w7aHN
31whIMb10Z3mWERStQ27sd9he6pCjLvqXL7l2zM2H7H1B5HOslxG4I7vggGoQF+A
aFor3foxIHFQPZRZv/FlBMFT6IM+a6uVOp4RktZ++Gbe+o9OKZcSu8QgyFLV8ZuU
pEYQ5vrnnRxrgkpsx6Z54MeyK7usxECRenOrgGxSNBKHZAwHauT5aqWE3QYZoMHZ
khDBOv9+BSmfIp8xWX0RQB1KcaWDh6TWRMhENSul3f28OWVI96Po9He7874JMk6q
6ZB14L3QntL/ai4OoBuIXOomeqIZbM7qdU8FOv+xt9XWfBVBdwZ0+bp8gzKPNIn4
5BElHBuJplJKIDd/r+HOk6xZ2s4K9IBYtU9aREXVyb7KsGv2C3N8pxZWan8AWMtu
FE1s14fMEI87i6ATnVZyBhqit4mUhf8/fd6X6byq8d8VDX8RebAbM4xgRnjEtYTA
2iLPN7FHIRbvHH1+BZUOBZXBRKNRYYPY2ZQsnGihmxIo2RkHHJBa8wKoWFgAoQLi
HBhoUdhUoHhOFwPIiiJEgq06+zPaKe1Gm397fxmvV5aK3F1XiqK7l+JpmxUkpVXD
gEhJKni73ai4h6lxeZLjobTHXn3t1CXvaaZQntsIhSDemdf6Kr3VPTMOTDs8xS10
1IvrhuxWKkmvCCQATTtD1KyBsyABCBmaeqw2gd2pp8M22o5+OXm+vSgbfjHTlKXO
0Da7266dlVQAnIejoIhyIK/5GEtP+IZhUmZ3ex9SxO2fmIGVj0LF8iG4Y8vkg5bS
zCP2dSTX9xH/YwqyCYY7kZta+h28+u4GLg09ctIG9NRY0Ut52BuBhGezlUvqywQ2
ZOf46PJDSBZEjMOu31UmX0kfG4htF6ryYW6M/I9g8gANV8KhYEkIp0JwNZM2U768
TiPJ1TXBVnkfb4e5DHjMGVvdu5GokHHfiFo0MajeZGML6xi7hb8CSZyPgbzJkcwJ
YVfmjp2y4D5Dtt40OBt3KNa6oP/ucuyyhaHnmn65z+qIOQ1X1zmD6ZgBkIerwEyW
AYb1BE5/7F5VqShLzIpkP6JDzPOlTmpaKT36S1AVgDpmeFzDAY6hRQyqBXrEaxte
c4mXDEzsPlrlJIZeJDDe5r1HnxgG/oks/gh7msJ5JYBADeFMhodJnwKyj+Ipl3Ar
0cTVZjl1mJWLG1qvogeS3PuBP6hmBeDUF2biDMjAQwCsmYfjoxChMW3ZMaoym80V
K7XzQBLQrXcK6E1rWf8303dBjq/Dukx0D4sE88Qrf9wuXABXbU9gq6f5QsJefXIr
SriJQOXtZ5Sidw3YehHkzfx/A2GtIP+n49vOiPaGLNIMgRHflcUG2kEobT1D3Gai
+82hhmTbzReUehAWCTW7ykYb8mVkRWFyZYSXJLwIQq3HoEuJ8K71XXy3oRo5zSd1
5leuyl3Ycz/b+/FafFbL/ynuASRCw/fOJKo3DG5n+JyjOmo2GOk5MA1qt6Z8Grr5
fbC60SE6ttneKF9J/0ZGYZQ1MBcyx7hWHX7SPtnxUeoiTu44kbDCsO7q9R71NMbP
KUSjqzmehMKpnMvIrOqeFvGitOq2AI9DESIcfofGAJEnvozPytXdjHFYLmELs4da
O2EW4Q65uy64W7F9TNAosYcI1qFG3WwO86SQoJYNXePPaIgJhrbVG4XHIbO4SWnl
3haWsDJ3gmpxKg/SEX07iEPddhSRkcLKeHkryebgTL4ITx5QRDsyc5FQyCiDvk6I
VuEP1U/wSwzmtX+3cLQFu98Lhie21esYH4ekSbfyCZkG0ZQF5lNDUVdXutRRUAI6
+79ggPN1flldBEatxXM4t2Fz8tqhH8Uqn8qGKvK9iCbyy1zECmfKQylSh7QabKrG
eN6HaZF0BGle5JIRajp40e9xEhd/L1G4eSLwKfiq8iAEMtLhHToc/75Cg+B9JpX/
oBV1a7d10Lf4QGClicL9fIn7vE2xRybN0ogwS2gtkOlxmpQw56rigmVbPeWea+TH
jMDiIA0ksQlcnzP/ZAS/YXGufOcDNORPjA78JPXLtkpc7Ovu5qM7ulKtLTiliwLM
ZD42eDu+tbd5IxNet8kNY1AoSV2TJ8kWkmFFMYKI8wVydaLzH0PGLZfkOBtKukg6
i847TmaMjR8uLX/W8q6mCSCR0XLirlooPI8MC0Iv182oR6RGCym5cWxmJBokb6Oo
vHBWArIy51jQTgH1abg3wQM4iCxHQrSLbVsdjrdJfWNSZF0SoeVQZmqgBdxyi9kJ
wAYH601ogihLkZ25Mih+Q7y6c1SPSXL90OMziaNZiE6+ETGxVQcxBU8g0qIv98H+
F0xaXqgQr9L6SrMiDnZMSwZUS+sHQ/WJRBbo7ZFIAMAekA+pbNGIbFsp1psXUb3r
Jn7f+37WmlF9k4CtOFUJnzqVZq9f4oCHjK9bduOTB1itnh2XGm+XAPtmMiVjKhJR
tiDvK9/UEJcCOsDHcazqGGdSyyKcDii35GZVzqAkYOyNMuXFy/moIcTDXKNkoFjZ
yupj54T8S75s3zHhKqAvqZz+NPA3Frd5jZNFpKp+sL93wCxLgJHmZNJ8YLU82OXR
yctSSws3GBmdengi3IhD+KVO0f5RRnU7hGhW96hpz25BEk2zYhQ09Z9rwK4NhQjp
8AeKGlD/11PByvI2lnb8SaXboeNEmAnp0vJ2jT1yLx4Nak1SSnmnXJEnPtsqIOUR
iiQCL1ru+zTdfrpv52CVanqYOjoP+kQHt4RIkR4x5cLuwfuVNLL3qy6OSbaayXDm
FU4t+Yr0aZsKt6PZMZk3FIXrQjUFwsiOQBwjlhiJ55nZMJgbuPauYzAo/BSmTt14
qvWlxIhmiPDRPtpQQdLY/UExMu2g91BAc1u3T4ewS3UohQKoNSdqpEMxPJjT34AQ
GpUwZdxVtlSzYbEX2Y5faoIiJienKdn6VEwxeyjgMJzQb2TOamSCHHW8N7Jsgtvf
rVMCMfTtdBuDGIZ0gYJWUW3mFMBCRmqNi0VmDcDO/zWPzFbl0N5TxQxpoi+vs5x6
dNOVmt7qDfaVyKT3N4wnmw7EQz/xbmZWE9babezLhNh6jzO3GQjmQ1nG1Lv2dwqv
LjT3TOD6ZeP4lK07xYfr4gIwyd5A/hCuydJQRzFVv1dPSGwVH18H98ZURxNEyQau
VXZKe8hI0KtZWOk8aW1qGiGP99T1Ygbstyp2Kl4KWP80qqc1bIR96SjpmudCjr+L
HgeV6umKwf4o09PfcAcEZGCWOqfjYnFa3aggz9YkUFphIyb0ZacIyj1fa3wyx+3N
KB8JwtJ3Z8qKvS/gECibWo3bEIkFu2u8oxDx+JT9CpmTEcMgx7DIGPYZZRRzz4OP
n2l671aK7hEylq7CSzypN6JZVKowM7e1b8GKgpGlVuqPjZCiNuHrLQiUxrfz4qzj
D5fIPL+G7va4FIxmmglYPIL3+nveFuQKViXA02F5WWqaWr67deuIvOdt1i6aqelr
Fxk61qCX8gE16C1NSXCyRjOrf6LDXhncF/FG7IBOXqP0yxQ+4u91HjmK6Smf0LYh
kcmvXU1QinX88Dw3Ood5zZQCKH1fUrm4m9caTzGatNRHldOO/BCC3aAFSVEumdZd
D03Agq6H+cFXVcL8pef5dj6kUe6cg8Wy4P1D+udMY9KueTkAEyzFbFmWhERYi2y4
yVNIWEoLWNcBJzkiuqMRBe2xWZLngldViDc4Lyy9VKZy3985RLRaG5ZDB/h7FA3N
t0+ilZ4sRC72ejLF8XE83fEth8vzmVU7mtpeZPxYFh/M0ono7nscFBWBZsclKVad
Z6J2+66gbCkeBKI7X9X3mnQv4RNCmKnuZX1gG+ozLqEZv3snX0ZOqG9jAHBfMUu1
FYBYLCUO84feAZf/t+EeKFUw9uMu+YY0mw+DINmBvHqgMVxjwZf8Yid3rY6cTVmQ
wRuQt+I16+jR+dBEZqiUxo/obnk2hBXC/ZwLz6Alz5ggnpwnyrcb7Y/QQFZ+b625
xRpi+7wolnh+4t7Hc+ztgPqqWORLsK6/HSoehgy4NCg+OpI8MEx82ygC5f7h1+Ie
OoTSWy71Pl6qSFe0KGNuhpujpRuKmWdmXMUc6TXIBScnOhmUK6VWIcfITDf9jEcr
X291UYlQ855DatXySMPHUho88tgFPXA61LAEJqP+Z9gSKHFrlv85y9jcT2A71ljg
jV1wCqGDJymMVzBrQIxthHU7PxU9d0kaSBCWynPKlnDQX+yfCq/c3hcSx2SH3+vr
JAmllRD/uZM01cuaZctFghOAnx9KKl4bzFoA5bqUAq35LTja7sMHKjDkiC+Cbh3Y
Q+l0nmeY222pr4BcA+xMe6wEJ2VeF8ELDDm+A7AADSEuK/qypeskMTW2dl0MoegL
PrUVGKWnJvgz/zvTRy1jS4DWFHDyRUikZybmNm1WY9HnTIwOqwDpbGNnqrgw+6jf
zPVe0G969oyyID1EhhDdwKCqUC2wN+0JhxqcEsMUpnB3OHAF3Y4xeZliYpENSIWF
omv/hM+/XlEeVKeinCURz9+cxquobbhT2UGxA0vHJ8hxEpCe2AS4bGlJRZxz8sC9
dn+tyEQtGSgHyz3FQn1JQB1pC3V8XffIlNna1XN27vrrFHIxsDruHhcrIe5B9YDT
2jQ40sbxIEp0XtPQCjmynX8VB/Pnar6EpgFbozkzx3kJT7+HBQxbHPWXfmSUnzNk
cvcRn4LIA7NdniCfwQdASuTdRgHYMBBEJcblfnV1JeFzCgOaq0pOPUlS6vNWnKIp
Z0RJAo2VRofDRzUcBgFQ/qQ2sdHmFSDHQceWouHdFRPYO8AZ0mVd3udUOjezfaT6
Jf+8VNvJuorOIH+Cn5W+JXRTsM0IO/WxTCqoTHYdfFuxrCqlKMYnHNIb3qc1s+ks
+DPv3S2e78xfCW2gn9C3bUQUT+HE1zFBrVDIA1R8gknfOLyhJDNLTWbB1Gb3BUc5
b75P8ZYahTen88juyuTpZPftDD/zxY7PZ+1dmZoJF87ggYYLxykkUBfizUx2EsDu
62EPOZyI0XkqHHDCjqbR1A2e842AEbBh1x8RRM2cZJ3Mcihrwlsa6/o19SqKrIEf
HsdW5RAvj1irmcy93t7sWVjhmJ9HRxMWjzGCFxoHApXQvno/UaJlxRpxnS57+zTR
BpsDNDj1Kh5fBTc+ymqkgkW31hQ1WxzrxUlk/dXiN6VMo0/YHllPniht1EGkdYLM
GnScIPtKo0TI0HzWp1TATot31UNOghMZreXcoG+N6110X87kJ0ZryuSQOdrnf000
Rto6rkc0bqtBByDBCsHFA3DX4PxIyxWlGFYJ5/AZpL96XD40hrrEilWJbxZgs9x+
akWo7nxjk9o3usgD8xkJT1O2M4odfgPO0bM+nA3ZJVF+huZGhV5H+RJsr5Db4JR9
2Ylgz7a7YV56Qf42zB9qkvZGfuqBNAPkiJF4DDgcH77KKhi5KFVDAW7rGAQvB/N5
l7uY0L4t8KVrlm/whz2YFCyHSLpbPUt5PT6RrgL8R7JEiDL/P2QWoMVsyFtTs68l
d58UxZQcSXY8IXSWCE+HvjeidSgw3BSXPrGUdQ8zQptp7K82wydED3Jlhft4qzLB
Metm4GlQ+r/x6SBSU+OKcURuukYpbo2+kybeyJ+zxQ/mgJmLoYlxfmPCRv3RitpP
PmUFQ3saRcw1pUF4NFwNCqTXEAcZPx9ql1LwYT+0bCki7nqApeBQT4lUx6LTw69E
UsTPIN3pNtRfrQXEAOrfzc6/osO4gra/N+k2m8tN8Clr0LpDWfFsNaI5TYpBYSq5
EEzGUa0iWFORKHdN3VGUuRTPSqBYYvRchmmIH4KB5y0xHloKq0L6h//gGGbrcKII
5D6LJ80DDO4SXrj19eZHHS55kK0NrqkWeTMCCXoFyyim/Vo4avrT6qKjp5v3bFGx
ynnHCOILmSH2qy1tBT8v5NpLeOsTVZGRkKT7FWPmKo1hYPme7CsS2CthqVuow/3Z
+GZqQcCO746L5QWlri70Z9DDASsrtIk3ZOhwNHWe6ll1kap7skeQ3fGdD3uAnI2c
rOdcVmgoyKb3CoDbdjVlBnczOibP097HzLJczIo1mTD9Xtc7SknzKhsMcDIwOJ7U
Fa+VdD4NIs71N6tbcG6l6btRzlZVSHedYWakKI4DiJu1IrHHZt70+rz/rs7LLwje
EdDQ/VrN4WE6RZfz5/y0Q0JiQHOLQeSpeOKcCYWwISk0bSRS+JVN/wspc9fq9fKi
6iLQs9ZCJCuyhxhIpvdWt3JHvHjwujc/ygrcJyX1mQNXUX8+pjhisE57k8di8qiU
ylZaIC0BRocwBkco+PflmoGOxTkot7MSkHyl2gQ8lFFHzXCTKYRaLMNzX7yi2l5g
v2DeGHz3yiMaQxa24OduzYp3a1+M+FqPNH+RYSLDQn3ZEGTl4WYkJQqITl3n+7iP
kB4OE4VXP+BL9RCEXu8baG8fxNIW5SMwcz10ZDVMzI5REg2bkE6bADGuDAjSF1AD
HfAAaYwlUD3RIE3nTntP0HmvvIJ/r1m4GG8Osw9XkuHUk7OZp1P5lIkM0zMyOWMx
JZTn9R8vbDQhI8LGFLvKq1/4MTvcYvy3Lg3YqFAtauDxBtBiE3rKiks5KwxSVcZZ
sJbDSAZgJP8DB90vr+NIdkBFxNuBAPx+zezIwJ7pLOAGtJ8APB7O6wTZ5kYTHHzE
GXDLXjyfrpR40lQ/JFbK6HeUlrRhO+oWFTDPesHIqNlKMylapA0kYzgJw+YKWdn+
ByY29dWTkVWX5tCpkZUWYTfQKb70lGXFnQ4awPaCJRRKy6+OdVyqbwA05TQEs+6H
IEmCPU41l4NiqQxZOMP5QPWDM6gXigBdTJZzQy/eb/Yu2mpL8tdrKMVuTfBeHqTH
HtIwW5l36GQ8n7M6+A2O1YW5xFMXp0sLF6+JnpTWYNTqsklHuRWhv+GOqrLXfiVr
RK23NwVyMu/TRDiqa0zi9kS8mKNenwRSjY2f7YGxf/49mHK3py7wG4EGVR2X/dqN
6e41HYbynkB2JNXiK1tuyjOOZ2JuCIAkW2rKUs+RB3JrlBbIsRvBF5Mik1m1cE0b
S4a7vrVyDk3u1Dd24zy+ZymBZOO7r/rrIuEGbfDZHh0H8vIHFReGXhsnVWwQAjwq
G7dpuL2K9mvIpo/kI4XaT+qbX+nUhfaLIgB36Qv5SFLxO3ILmVz2MwP5kpt+qSMi
i6mRxfLwbjz4FRrYDiqagQK6rdFODO/lM2cdrwRAkwzYa8NihGFd3VgH8r16fEv5
ASvhI7e830E9q5qJlo1prJTu8/wVjXV7SaZcZ1COB/s/qgVZoUaSuMXt1Liy0HHd
XcPrUMNJrF5tf/wXXRDWSAYmFH7++puZLL0qdeCzsjQfIEQ61sNlUlCIErH3mWCE
F9kbBinz9m9c+9o5zdOA1PzS/RKSXenHoDFp3+nZeIqkavfYXGyDVlwuXnX4GbXd
tGRx1BmQ18wI3nIx2f3HyJhuxyjohOgZnytqYspBvaBrr/cHrJW+XEW9jK4OLdhn
6OY3Sy7FuisbdNHzFW/q3G3baGkN0WNl74WdZV2pxbROt5ZEsjg/DQgRd7GDAZ6j
rp+qmLgazS25bCE44az/OzuHoPB5c57dD3muZHlh8caOQdugFXarJ4zM1IpJLVoQ
UKM6LuI1ad5K+KR6FW80q8YYsJp7AuIzyiCcF/jZm1e5xw+lpnRGdkO/O6WO7lCp
pCBqLEgSmbn1fZsr+/0F5ZRjScoGGkqEmJBvnF5MoO7hXNAA2u12BZF06XwobyTZ
E3MNfNCIh1nfJ4yKI1BhDGmaDjhqdw74l9R/xcVw5UFBV4fNsR63/hB1CqibK+Et
g0hU0pDzhz5YMNVTIWpgMGyNZyIG7dOni1DAaqktr4o9bDJ6SyunyDkkMVeGr2Uj
U70XBJ8sS0lUZe4nqdb2hHRwKRCSQFEXxLWvi9nRq28h8lPec2G5MveOgpZBmTvx
rAlstGdjNTv0Wgf8gldTSucxamAQzY+U02pIwLoan+0bbq/LnT1/oXg2C33fY7oT
6rh+bNN06z7vYtRE5KkQ9tEZB7n7NIERroEDT4j9Y0gFvT9m4dIt8QLyghG+bHs9
tJq/rE9KNzabHAl2nUUAyeZbyT+kE0vm/6PRNBTwrDt/TEqmZ+L0FjdTEM8TjWZO
gfQgUAFNHh+6elqWKm6Os7SRghmYIqWf10hxUnA6zPW6hpFFB2iRo2YmuKhiWHOn
10MtfTs7iJEqHriRWGouVEqd8+6KnlOLwubNboxUK4Rc4cxc/BgNimhUQBw9ZAyw
AUb/QrDwwzxpyPOuHPdRIvABp4inQvuAhTfse9VjcaBM9PONcke4GqdT2rjNA7MO
h+cFUyk3oz9uMk166iXioBNccm7+Axm6U/LnQ8PFLcsPIez7gvm3X+jNhtXe2Q/3
3VuwDpN7LyT7SdRbGDgQ3CWRMNJ/Sfr3pmFEQj/iqDIGv/07bqAckV7CygZjWUKF
IuzG9atXPt/XwAMaMh6RuMPilSpyEZxsMkklkz5q/Fgg3uLu44+oIDaf/dwJh2xc
wx3r3S6B2ScsHITo1OjHG37tNJA94J9hE/8PQqVNrzKbITtG85Xbofqpg8k+kAFE
wPoeXCF2megkO9uAU/mWm/krZ7LX26VGA/csJgjn8zFkKJpR5KKZFymlUsIyh/JK
XJgRPJUrSGgZWm1tHKII0A39GkPbL3GhjlPCGn9ZBKmyvz2d/prLL9Qe/yipeh1l
MWSnt0/gkeBySjSPzfU1Cz5ai6rpyveiEWTeaYfoWWFa8ydBXf829TrwDFJpvQyE
etGtnauU3O3WyxsAWWVVyqs9yANVSMOaqSF2Gav+4pjxebBaR2f/0A3geXQf5gPC
TNq/zM3rSOlYooJH20L/B3U25vlXSBEKGDUQ+QwGzEtwuE4NcW5mEZZALrIvuzIc
dbYOI36Zv4sAfyjd2wnhn4uKnuILcy2+32Sr4ED0hGwe4BVnBWMUdRRYEaOMd1PC
KSDaoFptIIuPPCWH9zxpOhlh9OwFHFf/iPmabQ9DR2mGNHzFKuwzuGHT0apIByMQ
ZeqyGcz2Q32/8D71pLpYaKnyUnOo0n1vVtuQx3v5f37Sqwda/oeF53jhRb3CWkkN
msqcWx17uzY29qx13ytysZIWvk3obFzZlLPJmUytoG/lkgFl1q64OsDMva73gUpr
a2xQ2XD5utNceUsHMLetKEhljW/G3L5v1XihrrRvSbQQWG9J3eVrGEyuygXy/Prh
IQ4i2WVOMb0RuZzOgFbGPjPQizFGWA3T9qdjBTSoc8vsUrO8N7dGR4JjrAAdv8YZ
7MMSN1puJmArBf0dogG9GCmAZOOoh8rIaQQo6KIrXAkrKzu3KAmxE0gkABw1AKTe
HkYSTjGHcaWL+GoazDAeQUK1AaEdlmPdfjVC3gK6HlTuTTEULXLQdqy6bTlhdI4Y
LEQb0EwcPh5fwhgkPLEjvhz2Z7P5VeIapssa/saTKHlERV8xZj/ygoUhmtjD1r2P
m4ntga3Nz4pbqGsuMde8NJjYf17kSpzUm2+a+TKgo2i5P0KKAR1E937xh+9zmqTI
gEbctQFg33VWdtYB6gtISGoo7ZgClN2i6b80lhldp62+vXpofcqVpS5tsZt0sZve
HMh5nxeduM5/YfHFsgeeCjtG6oij92uZ+PLWfsaIDYAV3m0kSKBLDV2hX3YDa8BX
SrEbJXkbdQuHl6Ae0tc5tSmoyrkB8BF+Ddbn7Vu7EnsZ1fLHE19/WTdG6Z6/wyAj
HU3WNWPNCBN1XQd8FBbjZA6LJdtx9lf8IhxIU8ZF+WQvX8DGA02k1bMUGlYRslt/
NYL4e3tnn2UICj3F5z3SBTzgOTjaZFEbneETUYivY0LkdPCk4aqFijtTdnX+r72Y
VrJhARE0C0MSHEt2aLeT3nJ490SlokuK5qrr19oZHOPRNwURlsH31Y1R79ZsrR6s
WUHXrXSPvl3WmyFlYqarst6F7MAswV9VjNADQviiKzYPI2W2R9Jdm21S715Y/0jr
OwOS/gzmipberHUSre2mvEHRS/+XUo1SWFaKRAGenbCIJ/gEYYfOEIq84XBtW/Jt
UXMsvenc7qrBuApjAy/0J+1LER/WwweGHhHAn41M9rUAzA+w67mVJBJk9F6uwEV4
PU61Wgtqq+pIV5DUBLIGYxvRfuN71qaoeWzo/41Pj55cz8A24Fo1Ko9ByVuQM/Ms
2kKN40xyS/jQqtV6Cvo9t/vodH75CneXp8nDSI1WarvDaZwru/BbR8MwDRT3znny
Y8n9rgs4NQjAO5gQa4UYFA5T9EsgGacu4dN7rCaSE41Gk0g0dqWrzGP4Zhz0Je1G
rkp6t/NiLa99WaTpIzEkQ2F/Kja2vOTcasAZ5cbC1dT3CeIkvKQ42QEwyod+eb3h
04/TLnZMUz+3MXBVEmSrVY9cu3k/axGzxADobuX+dtHqaDmND2+yHHrwiM7ICVHo
xU1r7hvrPnumlDNR7YNTTm6mR45WsuZFjYmDCID60xWvQRGRWZVJqIkW0pXDiPGE
cCHJWdSSgShPDEicTawhwcU7/u2nul9G379MGEdkOTWAuBIxWbzs6miU8o36cqY8
ppVO6vIm5YdF8xJQQDUVjAlAF/I1Zh4W/iMjWkqMlRACmPdBi/oCJExWdZQzP6Vx
bX59PK5zC5odhp6LBPdPN46GsianaPb2P6LDN7YCUd+YyL+vyj2aEcp6TRXZhFK2
jbWA1hwCkBrqEgx6kHui8FWTodHcUEKJTEq8MZR1wSymM5djaV8PJerHvR9HD/Fp
ILMgFKSLgv1fBQVV5+v9dBCcNYFIqw3N3wyRbJyP9mBEWDcOddPSpTBdQaKnz1tS
+MCHXPT3rDaGGdaOQBPHz7YGbLFnV+PFaIvbQdyQGV0nULIaZDNtlcudKgd/sk9Q
8LD8nZS1KcoNKYjzTPpQE0AkbxhW2kNpZWXcPhyPV6iZo8yokLOCXBZQa9ro+G2A
fxpmNqjG/GZIEscLwCMsJWy+YVVbtpjRZXI+PlbpCSJG+f5n1yoRrFZ41JrYU5MF
GRm/w4y7F+1dFHBrhqtLjcFgjsRy3muhxtLRVtPP8v4Sj9xPNso652BTDrJ25OZI
/ilz2mxGT6k9M3ScDENgYYoUchSM7CmmejKZIiiNO0+TShIIu3ZxedtzLJosSbQH
a1WeHOhOhJQewSTLu2Z5XzIenD/x8ka3vkr8F9Dudep9k+oo3HyhG3jpAd7L/Hi1
USnuDhBiG4UuzqxitcdY/dvgxrXYnCnOS2C/2yKj+0MuBlQM26tW6XkZVcWTjRNG
B7ahogUZLjhKFQ6PpmT390SaoewgoCFoCRUi0wDwp8P6IFUthL1n40F/VxKjLv+s
gCTYJd/gXWwX13lDq3Vt8W5+MHP3oSrrfL/OZj08SGq4R6efBdufO4jSQGnL2hT6
lxhCi0yt1qvokM4RBXCuMR+o58rE6LPdwM+xUShDDMR4lA+L7GBebUBZxKvfXz/l
bFlbHud37tTbs+9+cwpRWBdbuRTfJBEioSb2LEzUucqQOsyx1S6WQcqcICu8o9sl
s/4ptUI/GVCETy8ReXMvbwnFbBltH8VOR6CCBR6zIlrvPpLYMyigFVmTRWVA71Ss
5sII3hxN+bqato3EC/c81McyQhdCdfCBbqGPPw7SvmT/x7uxm96uFISwS0nUqPOi
/Mb9gm8Zr88FU8/o9EE/nPoa+fzYmUtJSo1GWcfZOmWaTGE4EKVx3xW8+GInX0zE
N8/MedARY/tZA8VkYyX1dssMzk/KX5dwBSsEEIquKSzrHipf9uzrxtUBzKaaJsqQ
12fvC0vN34IJs16L8PCrqKX814m82SP+Jw+7P98tt9sTqDf/ydmsKPeWhMkghH90
77HkKy/LqYjFGTVDxMlOKBVuLZyEC61QnhVAv4EpEOkBx3A7m21e+p9RBQ3yeznq
OdbbAdtXCjbl5WmsvFymJ28j4jnZXTa67YTBL/rL1WvwWrQTCB3tmcZiB/lBPukW
VCVHIj2ZHW+PtONMdZIBTFym8Y3CEpnyLsleumWmop178YlI779bslRlhiMcTGJb
6Qr3rJP2fDvlddK/P5sSm+Gcj4/vNq55Y0pY/a7Kz7zd7StXo/SXl40QLBCuD9OZ
76CoMkPWTA3PaA7ZrgZEbiF6wCStUJH7Y90lRJnLvcj7wr0+I4UAm6f7G2rFBHoj
rW9YNbAY/7SvpTLWHf+iRIP2Tcku6p74vzt006PA4W9XlsrzCoeSoChhcVdEWTzv
SvvaIM1lVu1r0Aa1VIYl5FX6Lo9ifRQJYPgjyzXLHBjgLee+GVtTbICStT9LkrAr
XsM+leUAdMindukMkEmxm9CfUjcLWO/v4f6nKP87P3HzBvpWHDMhveVlh1FH2/KE
VKTuPOJTxj6sqlCTfD8gJTGUEXQUNvHNPvucRB7C+sC4WVIRgTHoqNgW9RFafSQe
Aoccros8c4e5faUbT8Vy0EnA7UOgh8QUuk+rB4dUc817fbBJKc5WrnKK6QVLdkYx
JB+4wYHYfEm64x3yfFan/ma7zMxTed3AGZfL0RQ8CZY3+MJ6X0d74BE5RGglfohU
nCxDBtyKPIS5qCXgcgqsFf7fF3c6cUkAQGlcI5ryfK0kEqw1Gi9emYuUAtaY3ERS
PpQ8NtNwz20VRL96Ur1o6Fq9BOnu28FyWTBeTwNdOlQeL4adI1H8BYeQkFP4eRRg
Ev+3BqLiJfiA+bQI5ebj+bgm8I4XJfZCwn85iH4sBb2bW7MGlg0C/l28oqxdkxvM
4HxHq1kPxX40prKX7UzEqPtjiXg1yJow5sDcKe5r5WGmiZIf2fOJdLTGincZTkU4
U1DlK3iRVCRqMjH0Q6hdhgCstxcZp8K5kexGAPwSHGT82TUL6FUqLFwfSDuDoI5r
hQlQO9gez5ClIRif/6+Vtjm0AhPglSOtJ3myDTWxQPfKL3QKSjwNVrsQoRyOi7Cl
bQWMduQF8qvaqnH8rDXPiH2uVjAXybSphQ3xECw+4mbU+jZ1BmgVOsCxelmeLRQm
GplGS7tEq7dkOy8gWoOrvAPpEzavVhORbx7Y69wKlL4NkK1FsCyaUEDJTxndq+Nh
M+HlFfZpMmH4EDO2rwBpqTvzwzlasPrAhoDpxDu4MQ2Kg8lEdw+V6OAs5f5BjZ1Q
RgCDkLW9+RAP5o/fbHisSmxGcZ1UA1H6ri8M4jRpbHDnBPj7fsNtg5QmnVVsIWR2
usiXFmrmDQ+09PJ/DWSIiV5SDq0GEnv1cUOWeI5asy4cpHsEknU76NAUCccXmp5x
E79MEbhYaGuAI9LXEFf8sUCrSMW5TZy2nTYaWcBcOwlEBDFETZyAk5sa3vF/EkBm
O+oIn5JWA3TjSKorNgToxMhNfQ8edySGrBftRoUF1p70rdpgEzgq7frEFSqMSt64
zX9Ya2fgg8Sx6i2DKwJeBqGP34vQFejKFFBcu6dZm4W65xfCvbAWCEReMV6hesAA
pFlmc4AZnM+07ltiLUEGl3yPQJpjVzqlbpvzLm4b4oAIwdRu4jNiJKSsWd8BrsHP
jkVNEPkWCcAaivLLc0y/n8HIYA3D6ayyatNNemQZMVvj9zw//Ly7ViVBgzAOhx+O
Ii33l99nUSX3wnFSW9z56cZjXXF/62YvpyPzGa27wZGpW1XwMOSQP787YBMk7COq
RkrYRuY5718qmPuKivfw8+xTbAQy8W/3aJJIKZL23+99RNcdcn34A7OQqI2A/xD3
zSnwUZ3brWXm4dC3N0hh1zXLNdekTxJiSHNSVXCcBwHsEi0xAYg0wS9BsOO3bh+h
gh6jMacb7INOEAIqUmBfUTv7sIrT/GNy8mgY9UqAKKaaz+e9q9rFoyjASzZ4U+Nc
o8DUP8U4Qn6C+H6vBeTRlnskdBGNWMMGtAtY/QjxrSJdHs2NDrtUB4pv/nCwa6ng
RlnWyHFwk4Nxcf61YvvaO1xusZ8KqffQwhyhWeTbdM9Rd338fCS9E5VOaFC1W7dE
J3KvEFwj9YHq/yKq9lHi/k0Jwf/xlTUuX9rjOnZYp9CnHXZGflUG9OzO1UQSVkfv
EWT6FTQSZ/PxLf85Ev/rszvt6u70tQ0fG/1glu4IZuV3yXEEexQ5CMyn7ewG0/Ds
mjMIf4ljsGDLDiNevemsUJHsEDz8ZwdQjIh4VPB4JAnFzffumUaCRv7zSMWtBLmi
MrZvbbbrlO2lsaLaAq9K1YWmfFjQayA1wvDYEK7a2AQlHBy9by/M9x1iMyDIaCNI
uxjxeP+XuiqUzPB/6H96GL3qgYq1etWXCamoR9kOi7hsPJPv2HdnSRFptZFSr6h/
lpcinZZaZNkgbvNscRjrJxsPM6c7snVeugQP5KQxdTxzdBAOJrSb9m6TipKxMl+C
F/XJpBndADTfRtJA44lFP3A8tYA5X6q2QvFVyz21n9WivGx0tutv8O8ksbahxPMB
0rXCiKqeIN7dWwKwBzMTuM8mxjIKhp8zsU3y1tLQP4HvV4p3rhsZwFWSr6CkrcnE
wJmIKWOY16JmQaV8u7YM6J68hR9YvVxVITVe+X40WWsiOcGbDcMPMJomSfvDKlSk
yHtOO3R2BJXtPI3XiwBbqVkn07NtAEPaZvMjzikxGBYQ8suMIkEaRA7dXFA72L/T
bzRaRUrbk3a3ZOTGbvTTgFbfcB4OGWFZydZW/6z8GIDykngqAi5PAmIWTnqx9WUx
hDX9UVzNIUWl11MV+rBaf0eq4MhWABEZ4ZKcRswxMws+YTlrYCTBEfrYN5H62lrt
pR1SPLz/Afi1IHLE4sroDMUSar0p7SHRlcO8OOPYBv9gZuaNiIk+EEKuUWtjUiZf
wkpC0645+ZTcGmJAxAOc5olfYpXI3tVAgMRX/UMC8bm4MADbQ6/xGxAKAIUKkd7z
iDqyzIWtNUxmIwA1ZeHKvrwgbccuG/EbCAQAgXASAdUa28Mrm+eIdW+Fi6J3C85G
ujgEMVKtyMOjR7hvSX7DHTTA0xnN2P7F6ew7Di8Q1WMqcvhXi2ffUYQvRj+PMtw0
ymMDKGaWpjlVN4joDM9ExuNVwOQiLQ+8oOIRD0m9QDwI/X5yAnOXcQ+lxrLLt6Ek
4ERnEUV0fjR21zV04DfzsKraRFpnmbw3Og+rSwURUZg789vzBsEQoFQbWEhp7P82
d/XaP3FM3J8p+dEzbiyFgLiUyK5TaJOyxflwUpr8D2fzGSWDwZpx44IkTVa5KE9I
+lMWIXxDCT1lLttUtdqcpf2OfA57s59T7reoSJ2IsVuPLFI/QV795PuWopQiVByk
bDRpPitb3o/88nOwDk7QdvBAaAO+J6E1iNpKpzXtdrp/Eh4ECwUo+fMjlbnKjrRp
KW6Vqa4E5Ew5vdzcmIqVF7OicWp4T8mlAe1U5rODg7tP3ZLp5Qu/LTOWUyOjURBw
Du6S5tpsSZCa7sooM7eTNnenfH8MQaELNh2JN1WxRKOWZJ3q0CnzOpKxKkY1y9R2
XubkLNEFoHohtoOrp2CJYRZdybtOBciecoG+ePmNIZi/ho23dtsqmPJmxK0whOR7
FTWMJHmu+UeRgmfgH5jVfduAJqZKow5MuxGfCyr3oYgDZVWSV5SnZkGbidBNRtn+
7GZ0FZl03J3truVHGk9ISyNbQok41LdQXPkFOvBNr8Y83IOKCjQnray872W5Hr+e
To1GWKlUa9fwcJwkc7E5CmoTvfW86sgTGYKAlaSXXbkdCeVAhbSv6740fDu75xrv
n6bT0j4jQvJCWvwo7/9/K/F+3xXxarguncIIlqL+4SPBhNvh7Tm0HMZ86YQoBy2X
8lSTQNJ5FvkzZ2NDsuazWLozCvpHxj1HokM+eQRG0mscejz30FT6flQW5X8YzkX/
EBV8ogb1M8YFJ8pQ3Z1tAs9M+2O4qwBY1BJXqrRozCQZhjksH+TMXHBqcnTJtwdS
Jnxbs6ShN1VN9vWNLauUHXUF3HhA82TX47U7rPoz/wsn7/OxBFdVjcRQZLOFTGRE
XPyDNvW/jlQwOJ7xQZ2f727L8Cy3g3LKZ1b278n6dcVJBOFQHC3r4KAMZKo4MhAY
Vrn638DZDZu75FBKXtsDqAMWmnlzXborOyXa4yzXNTG0UChrM3H5MYXaGkQp4ZkY
bppuajNuvKo3ZZnwkSJHz4znzXtRuDtzAIUBpOhMviI+8rfHuCbHHqPCG8bYneG4
jtL0CzspXV5j1YVhBmjzrmOxlFVACAwwYv5paqao7y/wSI/vQopTv0H+bqMPZtIc
2gMbE/DyMFNCWGvT6s8UYY6u4yJYxMPQhFPhD3CBTxbPm7Vfmy/SswsiggMHjNH3
aMus8zYqC/VP4ocS2ES0pHDlQbw20/cDyjfuh3qpX63V0rhtel560CB5Qo59WIec
DmRXIwTASc8vuY1NytIx+QDWYvfcwt3hQz3f/RfuZsva60Uw6GHjwalFBvgoG22J
hAlApNi0qVm7YHcJIJOHqw3of4PLe+VJL6BLGCk0Y9et4uwDqyuu0f5jgFdncSDs
0NN+VCBuIv0xZq+P+mWtUBbF40v7FPl+1AS7KOz3MMXrFK5RJEP4St8o488uzlz0
x55c0g0nFTpvSYqyp0lx1O3vP3mT5EGZQg9ZyswR4bCZI/dgHJr/ZqGTuBNpxoQA
/JxALLEffL7U2TuPxiC8wu+Wa/yn7FPGl62WyL8awsFqz3TiJpKejpAccC160vMY
npRzTC0h/bwxp01wJRzCLcGct6mi1A7tr+qqa8HajOgSWluIOY4lwMb5vo8AD47t
PA151o7Z3/fg4dwlGpnefI/JmATvY/8vjG2A/OFJVxI7DpVWjEsTg8YuAsFFwDAQ
Wuf5inAAHRhVOZ4F8W9JFuFhq7uEAIksvFuYx/XJdpq1LVFVDndq2PCjNwrNbBQK
JmME6zpPk6Wvyj721owQaUcGPmRWKqVp1ECwjjSl3Q1Ltg0W/7ZscPFOUwpELOvP
PhjyTkPv0roW0CZwPqTFfQg7sVYJ2WAt9WCgBYeKWsd8GKgw5NKDLMh+4KZ40OhB
WbbfZM7f8v7V5KBAoH1+U059CUee9ryldjbwvZ6BU40Dw6XDFtGCjr9pgOOjlEz3
vIVC+zNFPrETgKkdgDL4P2yWLGK05zKZdhfdmlbPti8bScD0388cVgr5bdxSKGas
ROxT+IlP6UkD5kv6QcB1Mf0LPbKXyODkKmE7rVB6XMd8rAfk+G+Zk+py9wUHsqgM
wiVGLLQXw1ufYJJKzTITUtpS/4E1SgYPGPywR3y6Jvt6ahJYMfnvTaBKEkLyUI0G
4yF9VbQCuv6e9D4Ds8kWFljRRtJD0fW0PzClD0hQY1ayuQ48/A9F9VS9XYjgZq3o
gEF6SjMXKeZ6bOppKk0deRvd/1PDl13VyWD2/8oRuXj4MzNKeRYqXZeKZPG5+Rq7
2fmi+nkCP1CNBiIyncBWBarU9Fpn+XINToBjfLapNCW6k1lyTDUsFjonV9yApmGs
MhKGLqdc/10AmAxbS4tRcwX8COHgFw1PuTkad1eOarT+psPhBNXb+GioLpd/AWMw
8TMtXsevmQm3sTvS6Irqc73XlguLyUOv4Gt+lFIW7QfKBLdi94GuPe2J6MfsJa+v
leSED0Z7CZ4nyVphlGPj6IE5K8UGb3vAYOCS10BjRTHMUwxybP1EYSSHC8V5Mb2q
84qPlMhlq/Y/c/njZzn0gnVfn8Swamgy8nnGkIpoM7W7kpQxIjRPvV0+xGRPcUQH
+L1uw17fFitiyTljQb5AVVNsl2ToNPuU6jjF9IJP/7QcHhAZGCULrB3ehk4tfZLU
lisfvW66qsBzHe5D6BahdUhPwILGRmq4iOX3K2PpUHUySty32gkeqJKbOhcFCaHF
GbsTphzMHUKohRiYBEJmFNwc+/04FumZhDbwD21D0ex3T1evtvupc9AaZ1GeNODQ
FwS7Csig6HYhAbn3Au2vmol1q0VKSJ0auuvmkSG28sBTfW0/OkwP4gt6WyIh/Vfy
PfCnnZzxtcccZrDv8POO63EII0eJEAq60g9hNW9oTedEl+ru7U7i11KC8DWtZnfl
vheSfrzf9vq98tq/N+25bfvrvKW4VdHa1uEkTYjFBhH1Lqz4DUDyYYLd/18C1rsJ
0EHZN1F1qtCwG8EPcNP6HZk69uT/lFmsCCA/QYWcx3yQXABdK0u2yd80DPDpliSL
R0vRJODB7jy25gw4ifTSf31lgrc6U5DQE92ychs3Ph3QjGpR1cUrFi94y2Gn7gaX
LqHX8Ud4DExoNYRaYWMutHJ2bFXpPN6Kx2oGW0HFVbVXqeJpjIHumyl/9aLEWjIi
sT9sXaR8dhTwk5p56wlQc1abM8r6/X0PBJDiXGm2tuUlEUDpNzrPBkZlrOneWr+8
qynKoJcCWDKNWG0nZVa+RolJzQeP8P2GzuYe51WeDO6981l/TtyA4fTBqPNwp37x
nKoOTKKEtVHTD1/zxEeBFftXXGa2YMnqPbU1ZS02OGwD5eD92McDHNWdMLT0EgEZ
eF6uET5fAR+x7TnHtcDxksuKRmjz78ggSNqariOOw5+U+pwScxhI0OUe5SbAxUUL
w2SADG0BotVra8T+XtmKvUmYb90Jhug4DcCxTbGms1GxENkjaOy948vcl1RGGI+7
CgZiRehBvP+zvGMOri9HvK6yCO5N7est9Bjl4z/51+JQaxKjlst7FyBu7RsBTIT8
pfolFyLnZWHqze+wB22KFgZqcOABlh3hBZUBzHhq7Ivdet5f/Bir2Hn3ouyXyt6Z
V++NVc7Y3XAPqHb1ThodQITRHr71peThH9TwDxXJjK01q/m9Lt6KUqXuiWe4VnXp
dwfn2DxnCN9tpxZEVgh2eQJl8vQfXqVKR5z+N8Xqfz6vpvYL8A5ZAEWImPiedRdY
j9posFTweuRIDs2EWnJjAnw0zXNuA5Kc/B/bNh7RI5RWj9bxzeIFNmngan4ndt2r
7xWnJvrH7GoStblXmpqURkyQAX/bPlh3AuTne9aA76BsUoIwz5z3SbzhS8TjeheO
+iLCreIx7d7zBLQ5+EN+ee4I7uzkp+miRYq1aO3CPUQUNlqRDrTtHZKRdEWE5xkC
F2IGd+5c05giyhOlbHQ2h9GVzcs3DQv/dIoQgWzFk9Bv7nxdqm7Hn194cl2VfkZf
aZX5jII7qgviSYrZMFhyMOTjuNSL1vugNr3asJX70OdNSjwAsnvBGYoSgAw/wd+z
ji3uy3u0CUh8jUdpnk/u9q9DMFMumnDKSFam6jjD0A6peaISc9su1jwjnWaSslFG
HBhDmnKhCnaReMbwXN6asnaFSuNJVLCgsc87EoF1S00CsgxpiJxWhwa2PpQxpTPR
xb4Akh8iOfOSpIQpkpL1wyzTQZsjXtFxsMWoE0R61/g4WfKiLCDkvUlntgPkMLHI
097N5SM1EZt9omdpaQEIU2Uz+gOskXliPq1Wc2j/PciaukOIonf7qoWQtKbcdNnw
lUkQorI5zGafFvUe6EqaDaLsjeTeGz3huQ04dEUtVQsVM8yRZ7YbUy8zzIXWgL+k
cx7dLmLescHMY2mVGM8rRImowT2RIwTUOzyHuz1EzxaqcnoqNay/3CfWfrU7agEU
iVbGofQBmvAdqcTTjyzZmOb3eAuIszuWCDbWrVErjA/WfzKUpOXJYUU8x70kqm2q
xL/kLe9X8U7sIZtK0h2fwFSWFv5ixdEjDXjcmVN2PAsgIKRY0ps9rjiD2D7O8xGj
O8GdRfQp2w8WfQ0zEDT+WFOYZxv2jyRVfI/Q59oD7MzKUnVLaMqmsU8Fd1jV+p3g
6FGxsnsmjR3EICKUs86ipeBKhJJGGE/Kb7z8TV86W1u92N7a9+YEln+oLsyVOZnw
SEikyDxFFbOJmRby+IuYud+YkFHSqwULS9sR41jmzhv51hnTyUHa0xS9BNq8juIF
puYasFJXfq6i3aFZgg2EX3O5UkHF/Gv1wwv/SCGXBFw0U0Kt0/Xf+YL8wMV5p9Wt
FPUtWOCsb6eHwj17Shrfo42bMiqPGI0x7VhErqrNVNywmoXLMlbebn/wDublzJZ+
rk9CaMjvFO8ESTgSr/mm05YDtvI9d4ZvGdf7BM7lRWV0i7vaNfgQbnCHawUEe4Cu
YKwM3KNRXVGOgZdjuFVzWBtt8rP7YPpPNyj+bwJ3IRYohHAMsbIkv8gD79JvDu47
5QzovUTwBODREjRHaq9uPTRtJPkltlZeGXNQ1O5Gsv+WFcd9olXlPRLXm/rk8B25
XCHikNEmXA5y8eNeceASU6R7UEJ3ZBeZ0cH86hpJBumlMifuNVrRapZHjvqwuZOH
HJsPX3CesUjGTdPmLc8hWMa4efqhRpsSeDzm15LMbWfiuLWhpQEQTgb9p3xlcmqJ
ywd2nXog7SQ3ojQSeyBzr9MxN1XosWMYySwE7yib2y9/mt/s54OIZAObipBHXbfM
bL4NaLflnI0fRBkfKZ3UPouZMUzp/unLHQNx9SW+eaamSwC5j/yvyW4VAb2fglha
VDg41VIBdyAubGBYFVm+Yr5LOvhWO3nioX9gy3J2qWr8TbKArtsXF4/h7h3dBK4K
5339AkS4ot1QjQcF0HR9lxYZd3ShkJ7rYTb3HYULyQ0nZQ+laUXCOtwD7b/XH6cu
PEaUoXXFhik2433Ntd+kONjRIVwsf7Ja8h9sWUquUjwggGU8/TtoA66P/4kAFhg/
WDrpaHTwiM5FUzTQL9JFMjg1+8I4+CQVU5+r6aEyEP9LfR+p6bzbK5bp6LLPm5RS
RFRehnrEbcpBrT0x09Hbl1n+gEPULttnnbiGwHbTnI4ZN1iUilKt2W5n+Uj0MsMv
YcOKjOZdPfMBAIm3dcHVo16yGfEGgKzIQTIDWLYqSN8w7IpDIgqTXTiPRYWJLC39
BIrUdR+CYMRDdOSvDKlr4q77pZ/Tq3qKv6/bs0RmdSpiJ9iI8jDhNkyVKeoj1s58
HaW9oJOyiHmNO/xjePRjffKB5JEw0Eyy/WBBZoEem/noncE/chv/AazzXBRnOjl8
krESEEDF3W7RXotXO93ZWm6bfPms/w9o0kZHuTeCGwsc1QthfV6fdNusCru5KHJ4
GvIXcMR73x7tF42EHx/KQtymklx8MYbNUlLWr9/JHZsWt/DXO0zHz4Zx9B8HO1MN
kxjDC62D8EWSJWH1PHN5ThpVObR5zcDY5FJ2kZnt82bBMuKH5ZdPpKl0kNoHf8E4
tFvvRf1eToMgJ5q9EJBQ/CytJvOptLzxy+3Q7iWrYi85BRZsq+g+HqJJoBpeMMqG
tHbrkaptjHmeude6j/yZsVCOs1Z3w0w9O190KjcchFpVM8xzXQ8aX05HT+90VbTY
WOxvmSodit4pjovfTwpgHMbAdXAxMtLVpkzLCSV7xpDGahzxfgJECtIbwbQb6hkT
bmlixCaIDlJJ5zJ5v8B8A0gNKfmkedRrOOgSQ2PnFwtBl2FZyyDvIY8xvNXTOpqC
Fm173jWgDtRaZ+K3bz0NyNiUfjnmwRijUHn8a+3ciyW09NkR6lyeUI15YyqQhmX6
5RDn5jHS7SIUVqlvxeiJ9y8fVN5SJGsjwjkV+LqkvRHOcXN/A1ZWLu8U5WkobreW
r7iJYvATzWe9DKUoAEDARDb95GCOxBggmmR0r+S+uue2jP4Ktjm2ABKWyTujqP8r
s7zLZE0Pskpx+SzGy89zl57KREgZ976JJmGrGRZZTSAs0liUhuJAGMmmD2hgSnot
kvX9YJdzIKGdwag8FkScDKUcEBax0aEwuvmDgSESgyhgq9B3pgMBvp2TmbmDSFfF
A8W5CBSwZL7fOFajY8nmtlLViwqlYEnEnU5o+mAjLMYUpohSTCOOv5vUVPJds5ym
EI1HSLCPA5xgEdYqzGwLc3STwyARQx8OwPeeBxDUT1oQoMwpGoOrkPWwe7tMzxtQ
RH8hup/8DLKqe3yMQQJLWXEXorUIdDfG02nZ8Vna5ICgRhcnXJf1DKJOyB3r+geQ
TvYrcZiKKH0yrxY/D39j0i4WNjsBWyPgn9hwXVUra70tqNb7O5JxQaJziS0YVixn
DfD6mj/hSUi/fDl3ytbSQ3Q/J9fyGrBBjyFpWEkztO9tO2fPRXE0tp6gfwm+caQ6
j8rlVIEvi4X13LPcFXNRfsp2ijIEKbYtgJUKZ8VtD6/fpbCpg+3/oOpt/hdUAZpl
prRh0k/zu6/fjQaWTeBNfeIOsVxleq3QHYOmOu9cuKxu12pw2rpxiHmKuGGwj0jl
FBlf0qL+H2i5yDfzGn0+sQZUlrqC/wVpWeVr3zm2pqgKi0l7vRmjeeCVpBr4G98K
HXpbMbGFo3XvlOYY7/XzU0NCtUXT6HsbF/Bjz6Eoj6vbk3jJiSeNcgGBCN0s9Fbt
e+nzAbr+2HqWC4nppYcXWrgqQe8qy0qvFcl42nKSZ06NR0vsaVqzok1W03NamJVN
/J4ySzo3mYH8PixxOlz3w34/epM4QAQFoOXoBeJw9uNWrGsExzJqO5p/4AyyCPAa
SW8gVtQb+GU8+NjByOhwZXZQBJF7PiuZapJPTmagqKWvfkW1mKt/UZONopRKm6sC
3dHnS9j4W0R5x/+e/tfn6kzV6g//I73CemdTrJuST3rac8XWDDVvPKV+Q3RPvYYK
y3Gb04aI1mHk+jUocTlCCbSpBrSaEU5V1KmITavwSi3kaphzejMasVpNxlto6H1K
F816tMfWLsYaCwBYZvV5jD7EQqVnLQEJCeM17aAI1Fpb0I3NABTIrLGUZnjik+y4
DuxPGe8cnh+mncbx5dEXhWgZBGBYit1/BCIKKEyWJ5kP94F9s5SpEX+xRo4JZVvw
NEwXtgoelhc8fDDRY8QZAlDCUilTcsOfYr2vJSM4+2lpgsI/pXsvRXtfmY0DpBH5
lVYV21SV3AT3IqmVOLe9eJRFi1etuNkGgtKjxOuGJwq46AGi7YuyMI0Z2oG9OGBW
26mq5fF/dwKH4TPfpO5XAJCeZyZPwF7f3eBuNPkuy0pM4vQpILHJOyF0/+vnyxME
xxYKvP+9dVgKiOLSGBnirwaMnb2tNqHlEkhLpZPRqOT3q/q9UcVVOFp7fstKXSO+
+qD2UtM8PtKCLPleVdx5S89mT89PzghBElamg1HEo/cfI2eFVGJxX0ZFT7npUFZ7
mGmRCMVIaomqYJS7gqmuWzoR8m04+HJFCzNcFA6LP9xJkXWnojJFARh4rv+sWdar
Cvo73vxAqVF3Y0vRCe/iE4Sqah7iecMsDp51va/4uoaJhRtV0n6EbtUMQt/GOydV
p/MsRtTNFYgyxlW51DiwiM67ENcTA5KxCGEkXOEH7uuz71B06mV5vFvfiNLv+fjm
4EMUCb/NhfhtRsB5ofwyBcqeuE4Gq+Kl7MprzOaOcmaMcE2Zpwd2nmhcs45yWvhJ
c48N6kqyQW54gtCLjqXYc0+xbK+D82sHVWDaKiSbOrmYUKDSM8vQD0ljuL+5SFc8
DNX21DHggvvIFO79pxgZWXVbATUdCQnw3FEZeaD9zTULTpI7Hl1dw0tuRV4M6L9K
xMX/UiocNvauyJ8eEEpAfMsNHzZTD/E/yMU2RCpfd/arDvPDVUfpFU4Lj0XCHRE+
lOWDueNMIglk2wxz54XfX9FhPtpSe0JT4w2yWJ0R0qrourHZuIHNNIz2Fd+dVjMc
+osBZCLX9knXrIS7eGUilMXIUdTQ9zViiiHtuIXOXJN5/rOgVf0Jqp/ufvPwFRVM
q6fpgR4ks2vMmhdMUtkQYAwXBgp78FjeAQWWUmTP8WnwPPKEsIXKarsOlAD2lVFx
z/q7+y/p0vjkYxb9l1B7VniUCmUAejkwDGrQ1DltenjacMcb1YWdg2OH/sviBCDm
B9bkQggc+0x9ZIhTfp6xj8XgJqxvSmr9HZcKayLrM/IDu1ZnnavA9mLewhePaQ8n
xp4159qswgcMisZTWcTbu2ycNSDRYVfxqm4VOiQkNZiuwOxKk7vB7z0PZGuGPyk2
Z+iXN7SSkynqIyfl7HisXKYWop+nIW+cbnzmndcCKznyUMM41V0L7yqW7N2yQqSr
HzYywBWaDNXa9ehYRcOGi2BkD9QaIRi0X8LwY6OAlZSdOtxQNRrymTIbboh3VHdi
FRUE7xndQygHXR6/l2q4eWO/qZh1lz+FigbCyXT0WQuEjU9Z0WWdeDRT4X9xr6iO
8BQPiGj0x+gMBj/RS2kvI2WFX2unrMD/KYsV09e+Giq0XToejc0clAQXNxM4ircx
n8HlphH04+YhYQN1vZrgPT0uBbtiwlnQPeT1uCGMONbZ2knpKUUyET2TRcr/e0gS
ZN2yr0rOgDu0xwNZNXT1fqOTD70aVw3908FrUA5u2FgBf7Rk8tVZRMUL2EGJOrwR
7H0FvpNJqwp1T8qdKzY8Fku+E15lmmjIv/sH0E5YKwaeVYUwEx4U/8g0Skkaw2lP
P85ygNR1essLlx9ht/PWVqqvkfGkXyOOjYSpesupGfsKa29TeOFBMEg1M1ZwZJGJ
1bNDcpBPzsGnTIAabNEo6FaD1cBEFFi7DXs991NQJPAKrPXZsV3gi20OCv6E2xae
VOdSbYntFVqDeAyG5gTANCCzjHDoQAN1UwrQHDeliVl+5BKjgzf1y7TSYQFodn6x
OocCqpsGcWfrypfd4VZfGrrpqIfO83WWLcBFZmddE5F/3NLBKm8ASR0t/7HCFRnJ
CMjLmflRX8umuSCFdOcH7sLfWOYFw/g4dIN6DFirYshDw9WDCIb4Z8CGlLZAiM/P
mPRbjskBj30/JXzFwlKPXqJtByURUnwCaw3aEpMBJMYiL1GrW6VvbtlA7GPw9WIC
sP26YanU4iAPPyPJk9Pw3/+q2rRfV4My4s9S9cSJZIk4KOxsnQTYnXflSNuOYmK7
v4EQP64eDlDFVyZwYh/9TcKIUiEnIZOwj7xdbmqK82/EE3+m3fVXl8DyBAUigWIa
meiV9W0QJt3co8kSi7o7Mmc8SlIOnPjskqCGCKqQ0+C92XCKwKPJvcmNg+haVLB5
GMdITDb4fWvrEIYel7StRZslLc/EbRjFrTGgn+SZBX9JOSpbg1NjgvVPXvJRbftz
fLkdYtuFrsn2qRUEguixAc7zzlBSRKi/eZv38h2JV+d2X3KAjiUqDtKwCvmlfLiW
saqCvRJvkf15sn8OF1BLBIZSZEg0M0dZj0qImNlicVhklCXEHMvDR0SgqE1w90sq
O56GaRhv3JXYCtpLl/p+UuX1RkpO2z/3VfMrR509WNTH0x6OMrslWUFQgskMVNUC
Hq18cCatM1l3rqUb0QfbKSYoo4yVLm0mwrwwTMFqGCLqsfi9/VoF4s5qkUO+U6VL
iqjg1powHgaDmrVk9zLwPjRkwpbLfcj61p4vt40VXyjUFHvTUsOk9GDcSZt2BT9a
Nsnqy843S6LWWm7YQSaxjAMinPVgaa+YHO1DRCpnPcj7Qj138e3bT+z/CY9GQbYi
86FS46iH0rwsTDn9e2m2Io0tpkZ2K2TYj36L/2GRYPba59nZ+vew30gyy1vGPvkg
Htsd03IUpdAThqzg3iMfJOvpyt7f5avechyAQM6xN+ZjmKBUDVgcFkROrjQMJRaL
ttxIwN2f8XNMxpm8r6tmcFUVZ4Quov4HjoxcfOniWPG89DokwWUWnnM4N+UaarNJ
arK28C5be//5aqFMxB3PME/LyWq6hNX4R5iMQj124xuyW0y8Sp9ZWhLZw3Kz6sgX
2Nb7HUc/EAZM/dypByIqUJ9+7sVXuI3VXbIptVbC8fYWgF1hJyzpBAUJYoHVIbqJ
Qqn6sHwiRO2BfrnufHw0aU0apt5aVFG2xkOIEjr9KtVnE4wo+QwvLE1Ic/Twgba+
RCgtyb4hKQDgjoIQpYooJW2KDQxs9b4Kb7Evz3PdV4spFFy3UY3qHvCJVlPk4Cp8
iOu5tZc4owR2AXjkqxk6PFYZaqM63Gm+v9YvuHdWAOi9/SfTBi/EWspW3tEkB3tx
Cd5mitjhim+VhbnWSbufezhXcpGLUJ0I05cdQ63mz52T2cGig+jXj1t0Lt13C7ZY
zFlsNwVXhqpR/vUmSbAU0IwQtTgsDTKTR2UW6sACDWfsjbytv4TPdnwZHaY7jGtZ
mJIdCsk2gFnSeiHOsxJEu99D6RiMEgHEfMhXA3GmYH7lO+6R6IGviiGYjfDtLz4j
hXPZOOWyLP1sHIjgQEQszJJdazGcgWjYRE4xPG4jtrUdVDsdlUAvx9irKie8E1IS
uqEcFkfdpbSh58X3VByWNAaK8pOpDb4NoBat228NoM+n1k76b4Mr+cAlNjD4iUVw
aJLqaPafEqErpSFclm4ghRNERoVrJs9rOUmqVCNlV7A3Ce/hwHqx6ISbTF5tVtVI
igLoPAINLBafQunyQpKFhZUYFO6xgWSsY6yuWVWbBzue55Hlk3O6hNWuvI1xv48d
YphUDuj0LZd5IV4VoSJg3OC94mKzjlu8u9nTmvrrhUBs/Pgg91n7xTRmYVUgLboj
s9trodl+hNSne2k+EeMvQ1mMd6z3jf8sAJyCIrsS28Dut+sRj2prTSzUKP3GGmkW
xh1vXW0h+eLedaF42pLw9v/ZJm470cqMu4xo2BVrY3V0IdmwWXWtF1HpaN7AwnJE
ocQI7w6E5NVqBLHkG+VEpMn3DQiZ7aFdHKyRmQlUvkaUiHbifrGXFHCrqrZ31cGa
ESQkRcZVQqY+vjOkPjQew/DkisJcsjzbL2fJ4EclXPiFkLaAcIQnmmmgnjI1FVOa
sOtm/oiHuoxSnskLFMHVHZ+fMZv5Pw0XFYhh8qWZnnP7Fxt7VITg7QVD1uDpHqxa
JfE6CgvYrnhoTTvZW9R2YlGoD5m5nJJ0GSAbIveZPQ2bbUI81zEnYRfvdAYXvyPJ
0qm5NQbVeM3FRMxSw6iIKztn+xzYqPvGRNg/eOedvTNN7PnRfF3MVAdJx9kodqkK
FZ8p7Z7xmozpGqxdVW42os0+i7mVkC9Pcf9a+xLvRnofdVX4j+w0Hr99LTdjkZgk
FGaLwQ5sVfrUR4xjtSmVyXtbLsYrGuEber+TMFiO+mCEA9lZUtClwX+S+ICce5Um
47wTjQWtXY4bfLkj1Qo+7bV5R8ByWXJ51zdRummB+jlqNSCDWtyLN2kOUvT6HfxJ
WSQ3ibyfeAd485OFkuSGwVaLcvpkL5MznRtCsk4E9OSTam2x5e0v55NyoQt5Q7kD
cWOXQKyL2zsreqSdMB8H6FfYJ7XY/7+O54dh7JMWZkDXYKshQ+9mi8QNtCm/Lpu7
WcK5LcCVU9iHFiOjshZJQ1NVGiez1IeLqVel1Ehk77RQ5av1jOdO/5GWcvi6o41M
zUoQn4DmEHpDN7LIWmgR685iOlOGcfyAAmWFLeSIa84o9VM6eocLThtf2iPpkDI4
TEE0FRd0Lj8a7W2YEbxN6Vy20w8Q8+xd7Qz6ta8pyFvP1Mfh0mgOtpqNHXFyZme7
d+lHLMagFTRb1Gx+zH94ZQEpstlBkoGkhpexzSP/4I6I6HG0rkf8p+IG+urjfVby
RUmWcbZzm2ByCm4XxogzHxvOS/E8bR/kgy56ZSaqjbq2OAEBOnnevwNE/UYpj6bm
45+3AiMTjyE7xg3kz2+DVrxyub5EHVujAPFtQ0teOoS94UE6QPD+WqT2ygLyDKOk
xsRf4PpyiwOadnOMzxnVc70XU7fvi0YxkwTop1WMn+2k4SYr1EmclQGM+733iftt
TgAZ4xdA9CXDm5XFX3t2l5xbtjEPlNQ2lThTeB84YgF2jAUq7wmN342byDafDttf
BYOLBCXNKPUanj4BIbCS4SeT108FKjU8LKTe9BqCfZELgXMufEt6P5Vsc0PHIhbX
UpaGbstEPq33Unt8Nc761q1qX7p9gfUqoEOP/l4F58VQHdRd6RRg2VPk/kJG/4e2
WgPXWG0+Zx4oZfjtT0Ugby8s9SnNvZx0oZ7ZoafeWEEmcbvvE3L6nEBzZLnBahg8
JFezMkwdI1AEXOsETXnkf/ES97uBMPLkx4bV9me96NZy70XxL/ETW8C8jX/K6G+a
Xcr63Vhqi0nHx+lJuRkovNx87Jvkqm7R0kznY1ThThCZ/Oudvb+gS2+TANqMuTVr
3ysZYaPDXQAsx1jGaUTTTWpRAy1qLzdySufNS1ft/A0T6GaQj73G11hFcvAp7soT
QBlc1crCvBnACYXJEq/hR27btRH0OxrcmdnMfD7wsLKGWvfikrNkQvh7DblYfFMy
WNZMxg/9jjKk3LruGvVLZbvVf60nud3Rnk1X7PO7cqBZILRa5HKsUjUH3klIfE1M
Mneis5v8Ud8u2bFV2gVMNR+zGVuavA2/knqDr92mHV7BjwZm7ARo0nAxf+ZQBoZh
kInN1rO34Xg2VR+Fr0AgostKlH67vOWmrS/YhgzN+MhqoOSdM2H3W2vFghnmNVgD
soVTaKbp7f+V1u/5pHkTf7ZA1wGj2/UYKLmjWxvXk+yBPFuxcbax8iJU9mVF6OKY
Qu+jXwfJmo+AmBHk9rwwRPejK6PP8AM08vFR5pFL3VjHZa971bFlXnLy2QqyiO4Y
tkCSutA3LWpQIpi6JmXOz3qK9wF/VWZHa1V8nirM3bZyC5trbm/PVTcN4BhU9jZn
ATyrDaJZgx69RgB4yHdrHOxY9M9y8Ib3jhAZr2bMR+FhKPwfeVTmXoGIrHpsznS7
+zQe7WnXCq22QxrooYGGAAmOq59xOhjpFttEP0TV2UREnmVVhXCQFQcYWJP8MPj7
GbeidV/iuK101S6Y5IKj1r4d0tdxzOTqsR+OTG3oNaNs7jqbKyWFICywaWinezKU
mG8qXLwf+3w26h4GWWxtoimialBmWJoW7I7RK3QO4QECVQhPT15dE4LwrpqpFzXA
6YOPWOogHSDXf3tl2V6D8bGIZpkrzGcAx/A+agc8F4s6rzxVyKHvLpr0Fyl9Ve2U
vLq+8XrLxIPSTHDX+K2RrvVzJ3mzW33HRxCF8oE50ivVEJc+1Lwk//uoGTGNZPsO
8TrG7NFsmsjZo9lT3Db1eaAxAlFQJlBfyrl7Zkezt3yai7ZC6WG3Aavk9ipW2cc+
JgYZrwhgSJ6e4qhqcQ60amFO8LZQnNIP9x3a8LulWGR59Ii7OfZFPMcZRPsH80q8
7BUMLYfXp0c96PmjZ3lq9LW0/sAcr3VHBnTm6pTGVwvfJZ3nWwuDi6j+FzdVSYYJ
Lhl+Fw2aIcN6jpzLkU2oOrtoE2s0U5sgQ8AAFu2vcNNJ7q2KD2FUBmgQ6PcDXD/f
COIeUkOTihvFEUIXK4MBEEBbpIHY8fApRVxdsm0nJCQA5NFQUmTJIYoWTpA+wDhj
2R5UIKJZdhZYTGXfbcUewCWbeEXxdMeUqyUmj0VaCsVohAV5MoRYWZjUva7Zwimg
0FkhzZ8DfpbS8orLZWCp4WjZLxV0hyg44+WIlOeMxB/UAHQTw8TGh1EEdE84EAEA
AyngawcAujRWQMRcLoMEtHyzhG925clJ1dz/oJxoly8t1BaAFQTlBBzTplr9+ZZ4
A7w+xYWcUwS72TfWUUe2P+g9SywP2RQGhpVOHPEGpNAcnNs3iYhr/ervYi0WXTIe
40mBbo6LvQk+vKu4hoj0+mUPAm6y09O+woxx4JXMd1NtwvpATZEDH0t0GlNEIyFr
1zjHzkmvI8u0flrBxz7KA0kDoTKbLsLc8A3ene3pRJ9hk2K9afPaaaHb2DC0GlpS
ysVeX1Dpefhk8Es8DqWrvF2kgLraaTGjcPTZev6RY0Hgaf5+kgw7HhU9w3GsXhzh
e2G3xsw56+ApJF1RssWBtggbEx76TJsY19/+elFmqpbeZrUsChd1jImd3x+9Odvl
ptFB+jnN/GXPRHQAClEVgOCreAW3+oFZi0gqihpu2HQew57s+oWvVGhyqE+CABVy
U6J4tKHRr45gvEbiRjiqAuWt6P0Rg+5NFNsq+OvA/eWWtJdBkqgGiuaFmEyDkCWv
nCBz/7WG/bRZJo4Tqx2i6CuvjrTW9UBzpGN1xBXHhj45Nmtq1dBZzstiin4ze0hG
SiBwx8JYAP8BBTuq18Ypsk/hZK2M9UhH4gjEasT1sx6yJhO1xPXMeuucVQ1v2RGy
tfeE4ZhUH5mpnOochSMrD6qbRr/08FkaB52M4ZXQsufjjiyXLn1klZ45CBeGLK9N
XMCwnQ9V+1+QQx9IL3ixEStbmg03Z2N7dK/51FjBlKL92mMiS3csg/jDeDu/Lyxl
lCHpwJ0y8ChJ3FyZbOipyOQWAF+W+70YwHCyY54fqhpI9EZp1S8n5wUWnTvO0Wt9
NyS5gzXDGU551zgxl8Sr5s4agOli7o3HPK5RPkJxQCEs3z0+6OE5R/e4fpk+KIcL
BVaRWsakWJYsxSvNnrN1R3vcNZ//RF585bdSEr6np8frb7sEWMWoPo2PLG7StTPJ
OGGeEZpzCOaToZmKN/dYOXCWkBxNpfA3eYAguF9gHHO86hFaAZLAoVHKaSOXx0oH
ENdnFb6O+O4G3lVSb0e9ghrMvsQk1iIMe+7+CuBRPZ+Fvpnzc6LAewT0jb+ZF5PA
UJm6SyiogQ3wCQBx0Z3oY9sRVmZQx4MMZzK2m7oRujN3JkejE7ob+zmqY5Y5mbqU
K1BL/qC5fPyiZMVQPJJgxkMK0PSsH3KOWR/vIUrMh+jMstZA9oAEd7AhGlV9D+AH
dAOtvwrtHf7VqFk9zp3XBwW6y6nwgEEb43N1DXrhHyao6xnNaee1wjC0ZwyfT//Z
mTVpYtabRrxEqZt/JwAtu0AK40rtr4YeYDitY7kLGg8c6paUwln6pbcLB1kmtCP2
vCTu3f37U8pMS12xD+BKt1uiTZTkpFIux+RmIgnTO3FiZiksf5bf9J2g9o+p8+sQ
KaRLjA+UH/uxMTsbkNbJGsJrlYA7rxgeIl2JZsbG0Tox9m8ILgZkO6G+1HNYM92E
YKDuW/9A+YWzedi4e+ugMPDeUXvkorx0aNZgzUEqO/eeOc+ylv/zZsv8vn+K7Cqr
nP9i/bIjmc07o5YAPV/QQTbe2fY7DsN2rCvelsXGFSLppqPcv04fQNd18UFbYD51
5wvLd2vVFKp24pfOz8xQPpQssT22XMgZATh+6Mx1e6fmfJJZPMa1Gl5EiwKp/NhT
Hi/646cQqsYvvPHlbpcFDAMcz8RfIXpsmwZhLrEweVtxC4wIma+8OF/TYldCm8j2
A0SJ7yBFQ60TQrCAvtOX2uUebBRRW+ld1s/4kmn+aEu3j+9woxOvt6Hf90mmzMDw
uzG5EWGeFuCl0uHXGhhyEMO/V0Wg5D+1dCbt44lmofC07cmwY4VKFhDhVSssKtvv
tYt2+iSV+HkECQhqH9oMhzR5uNiO+JtWOQoNIoe0Jwxb7RLLl7p7jDVhLGTqGv3s
SNoncJWB33s3FmdthxEmG9iaOEfcs+J7Q2gqP3dX31Zg0fWPRWRHmTdnEMjQpdl+
0RJ6RMMf2h8r+Wmm/SHni52jC4LcLh2Ix9yTqvkbql+bmxgHiimie5PdqR1EmhAO
/vC6If14kqWto20QhgLL9IyHJZhbvRvMacPOvNAssDr4XemAPiZ/S8vnG5w8GBGo
RgRl0zS/CHUF7/bbvApkCSXyVzeKwLgZkip78tAOiRZBbSy8NWHmMLyeCQJ66U51
9LNK8YYgf44ofOYGzIsaaUShz8LJXzTSa9rurAYS8ub22/ukYU+y6JXdP8HmMgnt
3UsJIsKgYAPFQJ/rw9VhD9hHzlGZiOlV8xqNjpCbUFwuJWlEQfnsQQLvjCeeeMV0
E8cyWgZ0yp6K7cotC16hg0TWu82hkpWCpw4G8iMTEbnFEZ7xd2ILoV3rTGlH6V6n
gIm6pdBOVj7XCB9gs7SohRclPgS5bnXvNAvUOmv3OO3OVAFPwoYv/XZ98KqhJOoj
33pbf1D9rYmO4G40uQxadi6zhL+S+z1d1c8j+sWlZkxgkBo/bNPmD6E/MK2vrnhV
FkYcKWVhCp462fJQN8iggqSQdkcc0GMStgIldUfKChZqX6cp7Fz/7iXdjL1pj8jL
vYsRWx0M/CasAnBZ3iRRVUgADghpNmpxJrSwtTbKuYR1SGdmpGhnVLrl8wSb1ZBf
CLG2F2B23SFIchO0nY7LzOM/WWbpbXWK708GMlY9fB0ChYORcFsuQOJDatLXm0cf
TzOEEbC/YEFkWtZ3NFciTu+wzzO5xwOxLwTtmSPwO/8kiMAAhTkKrrlQVRqugEA5
2CSirekFL3iGpbh79YkV6RrJj8LLi0YUmuM0Wc+Ishucr3PL0vM4AWKtfInPXgka
IhyXb5UMOIIRyeXn1qobXJ1mnPAn5cwi0MAtWq7nUagRVIA/n7KH5zh8GWeC57pt
UbqKHmVWjG2L7voQ3NnLpsd0EB0pChRzdI9/ad5hgCED+rEm64DWIbsEMMDm6Rcv
WfQM9ReJE53eWtjpZB+G1jHaMbt7iYXap9+GXSrNTZ0j6s3TDI8c/CqziBM08i3Z
d/nCzmDksBGd80ON/h6ZmYg2a1CYg86Z8YGj2NU8SLxiNpPsAdD12y18ynybqPUZ
PtVHS0tuSJLVPwP2Pwf8P1Qggx5FN6wkhLzfUy7NNDxaqYnjdHnaVij9iz7NiuWr
ROmPlFNvsWG1LCeLXOkWENv3IzBBlKFML/i04Jj65ZbrTXQW2jtE8pl6YdoHPnwj
z7JKb89wGQUYY6vIB0cV1nwxvF6RMAQKPd1FUTTOIfmoY1/bVmpe9jtoXj+dij86
juuAgXFq7xHer2V/6S5fWJDEt+bNalFO6nZPni7VInBQi51MgOrfV2BokliU02rr
gd+D1FyXVX4zrBjlQep4GZ++4BlDSeWAwaM52dYDaTDHJB5N6JsbcbudAFitSRNE
QVvO6HM/znLDQiDzlBe7rZIhNrNagjpJ4b0a7VXf/hNZN5uWMc3fGyqEiYJr5axY
DY+c+g81Vb926vX1pGeYstXUz0xTdCu/j10M5gzbRp8UBK4oeQmCWieLyTevIUE4
nKB6nvfxTtigZnk5dupDNyG7ZDwELqAxLZ9IUvJLPIsU+v/cJE6R+Ikj/pIuip+g
JN65UvZ/Ys2s1q5heF7tjERQCQJCR5Jg2SWoFp/ylLghQMXEtruKGHaop0c1URQX
n8OWwhmqo0l8Qb55HN+GGFakpPGBi16mrt3xBQ1bswq4F6f8y0Hfptkpv6dSwiTI
sl/IEp4nRert/sSp2ZsF7CkScHnMQlFHVhXOxKI/l/mI/H2rnan47THSFlQfU6VE
xThJsenJfOErebfsoEB4GVIXvHlNdyi4pPUkFnD+G136g2ro23TAZVNc8JTFSv7A
6hpoDT49MZLrZzK9LJvmKHqvKfSUqDC7RL6OSHdm8LQvGYhlR9OJ8V0G8ZsdWlCC
axfwjWufOiWC/mliEJZSBjxEzuTn6UlDEN+AatVVsgVCUb6S+kxYWygKA7cTirfe
RpayEELV3olkmDSWXhdgZsLIShI4WMVkK09YLzduIEa3OUn3I8VPy9e+nNOblWYH
DsGSWO4caJj2HnooXiPGpGl9mR4cnsEaNhUrQkq9ut7Jw5AAZn7QLTxSC+Yxcpp7
9fEzSGuS61e/eKM1wCCJ+GIdU5mgy5dkZpARy8pao7fPSxtWzNiSpYR+xxzWG2ie
WCP0t7Udvr4Sw0BBVyicBypENVA8LnKD0QtlQ6iVi+SZyHrDxbi3iSA12pSoCNIv
PAt730MOyyFdt7x1AZpt92J5OR6Ll/tG9gJQ6uCFEnuRWbJuJ17lRJyjPM35Qtg4
ZTU1KkH1fZqWzzPJrQWBSJ8OH/19b4+wIqAPDq5emGr9z50mBIOSiDo5tByJoNyX
BRhjbKMqNqb24rVv74T7ESXn0fO4xBRkBgGRRIPc2szHEhMPymLbmwEpQZ/z9LLS
QCgJ38zSaW/JqtDf8Uqu9JBiJAEcI9RanWIDfMCkRy68iOcEWUHOMawW5XyYXVtS
4X3kQ0H/jnGbpbJDl9FPuQqVRo2xvNawYOdwjDyhfnEMnyTCz6Tg61PxJHserqtL
UZxxMCnpQDU87sOh0XdfBZEiWD5KaiOkILaWapwBVRTl+0EP33ufXeBeJAJjDq/S
WZTdiMYe+HjU7AHphk1SR9i537b4Tqzx50y4qawzCAvnafKszAxUwnU0Kp72kvy0
s2lb/8G3msMqerZiJ34DhWiZf3cHTYX9YprDChgyuGCsa+WkGH/V8Ot2k7i2aOG+
XjQ6vIvCPIlFGpN/lfGj1nRzAIWn9iwj0DM/l2zzc6qY3TyR53ig04ZWi9gDdcLu
qpk5VlvuncLrtKc3vLdbgyoO/0BhPkcjyLw1ESEXOgtM9ZIcIP+zR2yv97NL0XWK
1fLItKrsaSMDIZ4JZnnEUpvFCSH+ZVT9EHZyOB6RbjaW4zIUM+HhuwfiP0z0yU/y
xfnr9e54v7+jhytwL1e85AVJD+9YciChDAvDpTyOPFUZpSuzEITAf/YBPpXYQ6Z8
8xV9N38ZX4OD6/j3CM+Kqo3EaZZEqMz9X0hlat57YGoZYcd7zTuOUG3xKn2jXM0J
0tjx5Ojj9d9Fkr5TqKoX1saK7ewkHNmiITW20uUf6pxJm3GsLeCkD+TMyTyNiThf
uXa7qP2xR7Ddxons7cZV+ZPFwFuFKSyV5LzVNVhW31qSYIC7Xm7KomYDDSt/7DbN
q3u97TYjOnYIg6j6Nz3GuJmgiw6koNXxhM//G2lxISqo5PCOAZe0JnrQbSDB5Fn1
lBdZnBmt6OJUeVgGu3quQIjvPALWR9dRhUo0HWIOohcLm8KL/Aa/puLq6VcBMxq6
rpfcZAXvqTQVNHLzQKXBdrXq5xLy0Xh9ItaR2em2DIa3CRMF+OqwZD15nbkpn/V5
+mOsGAnukVa6Za8UTMeB8URU1hT8ixO2w3sKFC7JWE3wDjobyoRjwZC4kVKBmG83
3WFBCyxKUA2oVa1as4kG1K8/omN5/FoWMofAQSvY5K/BXN4Ww6WUQQrBU62Tt3+B
dyekp7ZR8NeR/aQu445XhnYG5lBl4yoxFgBLIPP5iCTK2NiiW9yF23vGQU2CuJco
HULb9Xvzu/HX4X6tNGmjp3bWGR9vE7RJf/UGHRsq9tGHpYIRN1x7Il+ZFZF5k4a5
PSOYoTuYdsX3dhW6avhlQsptqOBzmy7gl6L5bqNmko810/zXAQp9aWo7hHKV1ENr
zZOXZJikgovRdqXU8gjwKGsCU6+oX5GCqMjo2tzqCyaIGw++GuNi86kpnbVYSO7/
4qc4v7JbhyyvGo7M1CWqsOsQh11Eo1q5CxM37XHzyLQ27gYAuck4sPig8tXYIzGx
M6As/X9y+MiEQPm2yoKfjXPYjpdpkcIzsa8hkEl7TMaWNUe/8Ssx1IESlehOs/AV
sQR9x5amzer00JQc9ZRFCmZMuRgKh395LTiXp9h6yTy5c4oAgI0Y7NTMQBWkXII2
rYKyOsYEuX4PNudn+NyY0DJmZVElI8kfrHVHK5FO2FS4CoH5h2+HcT9Bv/sbgfAP
73OFkD6eEUHHFS8hfb7dYiaOLm8ib4ycweQW2RESrqK1dO1DJ/SJU1N2p5dqw9FB
W+wjRPdcdvc20XgiDwwDdq6VxUbVldOStDBa60GI0pg/qnyJobWuwnBWeXi3w+zn
Ql0GiyEDw0QQFeqv0bJYMMl3SSczXcWe9SyzIkhzsObCe4lTU03K5RUmIVP4gKgX
WgOqV3hvJlvkP1zKauKIRIPNmH6pDDxWYPxQvPynExMMVMH+h89WKAA/42sWDukF
B7rDblMm9ATaGkunm99vqOgVGkjl1tBhnMqNpgn+K3N/Rfol9ZvOIX5MvAwRy99e
A/ZNXLMWEs/VEHChjyireA31ggjSoQkDvS4UVJH5cavB90rdcMpRpspwpdW9eFkr
PTK06jV3CEY/tGm4GSMycbiMqT8KKGTRmmtpgxPzamvFmyQzSWffhhfT6N/Bv/n4
I2+LLTY9pKJq9NpzcIMWI2r5VAUXRxZ9fvskXVeQcthfRsrXm0FKLX0iKUd7Mr1C
jCaPIHVvs9aHM2Sw7OrkEYdtDDMCiPKABj+ZI7GBI7GM3YJcCAV8/goXTapyuUAa
Esoyb5AMWtRewlb1sjYmq8Zc7a347aUk28AzVP9rBXE6P3eukPYGJtzK40dIfqIO
S35YtHvkd17HH1H4lAsiNkGBZHR/+2SB44+lg0/noZcsJ9uBiWrIBnQL1ZvBd1kK
Tyd3ZHxP2KlwS9GBO8/n3Y0Yd9385zmW1WwGZ/WZkFEeAC7iGuO0p5rzx+FhmuIZ
DFFtpURrED5DT1DBNIAwEnXjfZE5JRwnraT64jbyJzTsR1QrJ0KJYcJKNkgF8+Jk
WVLl712zWee7PDxMAZVC610/bmyHmuySKzunGV5w3EfqMST6174n48u98yZZ29t3
me4egF1ZoQkTkZ43Kdc3TE8lJVZYZ/4yrGPjUoqH8g068hHx5yMhNRz1c5RtbQIo
ewY+aCZMGVSlyMYkBVchLbu4rnLUiRLuItvJUYvtvFPmtCC4N+UeTN//5ON+wN3h
B/Ho0OiUL2enTr+6ubGzoF9RvVekfbJlCCRIqQIt4o0SZHVTiO56r6Rb/yyIbF4R
jH6DSYmogmcPyH13KwKDqKjctH98ogiNyVc+KjRT0cSc2xcGXB3rKyizcYiGi34z
4MxfWY2EDYkwrMUW2Ax5z/gb+SBcGndf4vAefZxNEzeojfOWuI+5leD0dafdzwq5
kqXEG4oWxnvz8nMGuluMwm+vp8eikst9A2CKgK9Tl2EDd2ODPHv0tkBumBPBLNYw
vxhwuAsYdfxKiRCjoG1tKCsXw+AbxklKCYKGHU7Ac7qGChPpqt5PIHfqR68P3iMV
g5KiN4lzu5V7iBL7gq8N3l7moCupOVGwFu6ZROCIWSg33RE2VJF/rpE2Drc7a5s0
ek0owUQ06aPDhxr9NQ0UlRGpRZCvDnJm3oMK2rjZY60ouGBp926/13wQ1npHxrgj
34bn38e+y3IUUMIWBWtp6X9BEvziv19gxKS93m5Oh7oV0to2iwFuxyVHsVkXfo54
N8MQAwgY8EHvmRp0j2nsHZMPWEGTNkhdo6P3a9WHvt25NiIHfoltH5aKV6Xr4aH9
LTnNqKYk/1vnzcbYj5yjYckWk9rNGjx+k2OGfmYeCXTdRhJY0l5ANdUc54Kd5q4I
6RU75OsJsQ3OLgBjMQ5RK7kBqvb1X0fu8sspcFr56tRQNb5Rt7oXRqkjjyshEHLn
lfptbsPY7hDgaUNK56/Uzed0smR60O0+XFD9F+r8YT4aD+9+vKt0P5tHP0eTkhBe
vd+OJ8+MMAgfWOGlLwtLFWlMrfKUe/NU+FNt1vls9+AltrIG+6sPW9TSTaCutAbb
/TD+FQKMr3hKS7RSobKA8ojDWGktkQT2KJoBYRMVCysFOi77JfMI/TwljInrO1OH
AMGW6eJAJMQLIRmO+0DpDop6J4MAW44YiAFtYlF7vBkGjVuk/YAIc5ovYRfW3IOv
VG7PgrXVQCwgaV7EQmi0MqRS0SE/ItThoits82xgiJVQ1juUoOrtd+yOG0WhKXb4
kycfywsxJgslz+WQA4KehL5Ggtt/bPB+32sTlJtAf7KaMDUScQqabWw3rd41MmU6
bhvv9q7lSIm4heWv4GJE+0SIaIk2wSArb7VeZlOdG1t42t7HNe39VnR1btUdVQvT
YwTfVE0Tkm9PZcgSHj0Tgos36TpZZNCScsdGjtNlaJG7jT0fDARJB2o2JDRIFz6v
1+veP/MsKaZn7hgB0m8Rqfx+/B/SAJuUG/4LHAybK2c8JiCB6ieTStlA/17BqB6L
2Oxcx6EJ83v5+lk5hQaSMi7Gsk+apm3PUfGum1W4khin8YzKKKiM02UCkuZPaSLT
F3OoZA1FfaEwXcELSiPDaY+eNjFs7gU97SdmP4BUxbe6DU5Gj04vNq+oqS/kU30z
s/TCmHql7I1a3p20HbNxEtBMQI/l+toWDQDr7WNJky2zkXIF/NfjHcfu2wlIQ8y6
5aBSiHh5PtNpekyGZnegyxHIYEqvX1yB3NQX/SDy8akvsxAS5yjfp4Tuj5PRkxQJ
FWeWPwvbP6rlL5ptUl7UNHykcHhD5FAmsSnVoEdg1s767ijeHWu+bKmofEoQFpx6
8/ZcJkkkXs12KaNMig++b739RCqRGXt4jdOJh4Ow6VVZFvyln9HKA6MjgddKUcOq
7MY4Qt1LrTZXbqjbKTcS1V+6VjsLH/3k0wFChFNQRYMATF7l06IQl4UN3JEWjklw
r1uj1VhCNvIJYBBxZPhUf/gZ2a4gsl4HKHSGRCDWXVVO1jEfdmYD5vosP0bLlVq1
jJTFRdvQ0IlFDwE/V6s50+3Qcg76sMOatnMAFYXSVW3RasRbfv0y23fVEtOGhsgJ
O13ZjbdJ81vng1vDugp6CGLocLZyUn9OJE9X180dCBa4z252QSqpTPcUkBlBRWmY
RIBcGBmYxzZJIISYe0FAGwzI1Os8BMM0ULPlJFETQ2AYHBNk+Ca7UYJyWA2eBVau
UPjDtcVIil0cJNbDuE1vDyd3qj/6E7fr4v9NuPr0BkEAH7QHYSlpo7YxhuZdFMvu
7VmjS9MBenKMkyoo8cDNn2O4H/MDFwmAa0E7bUof6/VOv5Ux/0GabEMZKgNCy4W9
ZX5KQWcOUirKELrvxPcNGd27fhCkC+8BbWMxcpaAnuuk5/N+twG3p8NGEk+klESf
gwDJ5B3q2kR4EUhMkv4FpIZLJz7wKfpfMGsX29Csp3RVZc5vsACfweRn1gqUlNf8
cMyktAkJzVD5Quk9fxJ3VKdsfYo1wnBWYwdEf0R6Tj/qdumiut7JgcXtut856ddx
Ndxnifrd01Tv2WJvfAqDjU6l/JQy5+A6JhOIvfz2p5JaFU9aMJ1aFYKrU9eqOEEo
0BAsZLJLpL/JBSvfeb0knSFlFAd3xnRbwlY77tmmnulQEC2AQJ+ZTHktG6f4uagy
nuLyCt1fUsh4gRb4bS/RpoQ0kPgmII4bpMC7PEGCLu3mP6Rz06+ecTc4llJQLJR2
0Oox1mb61bgOA/CE8yjxyQ3h7ymbD/IOtrzHMMbdl5i0YJJM1vvA/QIylAEaJGzQ
qoGT2WY/Fw53gd9HYp1x5VBGu2BHqpxRgWfJuYeuUZd/iS9YWM23TPbaDLYB9cJK
3xomzId+/+05NkCW30GEtDisiodpzJUj3oObslm/aoH9jfA8XhYs9q1Qq+xHp5Zu
U9DwIHObR3/bctFK1hYa/4dEoeAvP/s76jU5waAoGfBhptir5qIfrYrmrdpa2+ZZ
09bTY2TlIDqtnwVfFvDUIm1qXq0nHPSedS/fS5bJuwlKGPlnNG4WfXQCfPy1gJYu
CFqBJyd3W1jUQWcKld5lP2Ss5jnlHN6DidbWZb07lzF6KNL7K4hn+QDrQgujBKbS
gINny3BCsaaqlpoHptRRyuZxz1JIF0wuXCU3Qx8gewBvwMX25ixcMju314guIER6
+3XexgFiqnVC55eaISVhnCIkXy9UhPgZhjxYUDH5zWKQEPE7afSYQLgPM3vonc2t
gt9GrjsvSdtC6Ln+dNhqc+bZw/DkHN94v5c+ZOU4YPaHOS6uNWeT/yUX203YsVQz
y7/uu/OVCO8hnRgqfbYP3/LeNsdAk2ACHSkSxtO6HOk2kWblW/wSp3Zph6DUPvGV
B2WkmSNe/O08NHynQQJ5twKaY/p4xYc3YeUVulPBBDdiyKkZB1VWST0/z+hKDCBa
tiYI5OTdJp29iZdRiL4cohJIKbJGv6ZhHyCW1jfQfgV/pGODu903YnFcQefoZIk9
OwrjALWlgbE9tR/vIU6Nm7jaqYZEz6qD2GtrRs6pjn1vNkhry1cN9rRv+H5t5a9a
AirlGzyktYAJmDrVwyxGBePTNbL8YkSyhEW81JRaAuyHUkTPm/tZayXSAe/X2hmv
Pp9IQL12aaTMtg5kwjhOR6ekzDE7dVrwTgJmn8VJ25AfQBYwOjmRBLmyS8YrpSKC
z47cAlTbLQATvrr6J+e+L+OU0eid43MbSMaMGAUR46TrkwMphI8eKNY2uEwxw4Th
HYIDdCvTMoVZQ8U/DAyx+cgym9P/Tzz7NnuUzOQJoCabo4VCkTxMyX4pwDh4HdFG
T+soQYyqy4uzwsZNId0dTS+rBzf+x8gBie2QHw425bfgjRU/q68iDN00HJC7mI03
FFidfmvQ7VRczlV60QztZ4FiY6OklgPnsH0+XcWipx5HNLM9eonb7R7BrU8GiSgv
TRY3rkCXZeXzwNsClDEyDJjhj80WDIqUdTVAraBOPh7zLrt9ZudSCdQEU6jIW9Ls
xDYIV1H4MYnG5NwP7n40eSgae6WFY/rV/vdl7UUztoWR8rO1GSRbV8Dx+RLtZh40
Pan8i+PJo3/MC8wqqKlK8SSzSyo+qhY2O+65PbgP05d1SjHuw+IsW7pI4PgpRs2z
wokW7agONS0oHQKj8H8Z1fw+BOyy5zfVIaXdWdkOc0zo8tL10y/a0zOvZCrBYa+K
3ln+vAS+LijMQicR1HmabWjYvh46gsQQH/NdYU0ljDCJdJ/tBg3qg8cxXzySLyq2
X+FYmwV0nakXazOJhXAzUEJJjm/bowo/kedVaRlxuGFj596H18iCXhT6vEeUkgcV
7pRMUWzoiuV/vAG6iE4HIDdtSjK9BeBfbm6fjrvfjxn/+LM7Sl5PAjMy5qgkzEtE
s0jG56VQTX1v17hXWWdhKffdPCka+PiIAqGUjk0OLJfI0ER0+oZNTc1MRW6uLjtA
sTjl9kqdzGiLi3nG6augAdorAta6Ano//+CKnIvLdADz9db9uClTR6cE5ZBquEy1
1aNwHCfLUsH3FUv+J0Lo2cvvdmI89OgT0oe3Alt4eRoF16RQh8z0MdwWjmk2/X3B
cZ2jVfzoIW3LIRjMMIkEZjda/1vWiCZvrUpEnxR2YAdpzFjSls0mqsl8n2evPzJK
hEAiQxyK4kSeHPTeMr4UMUMDV3BLOvm00IDPIdNnZt5xCJ9ar2v+61mY36hKss3U
04hWOPaO9jjm2dTRDI0AxyPahbQUQs8RNnhko2mzJmmdFfUPklxVbXouhBxMMRhW
MfBZPYKpRFfB923tyDMSrRppwFv0sUJ2Uy2Y5Og5TmOaVZUYn77X8JvnOXl9S9yf
SdliBno331+/Em2QXI/g9CxyGjr6RT5OIW7yFtGZX9vv0CfbVIMQGYKkk7kaGnhn
SDCokyD7Ba0gVN0QHys2syj/pbmYimj86B45pJtMHEH2MxXwz5xDmfna6fqpQpYH
K9alQUEacQz3+4rE1MXWub4XQj+lhzlWY0dEwt4guAfxS+Xm7yi/cN0HDuTJmEsu
Eu3roVCiwgIx7FyIAI5UyQovzlZcpfCYTY3I55Tzlh/rL2JsPOpcCRVYj6SLVx4b
fSSlAx13rkoyaqX/CPn3cWcysOZTgfvRGWQ7gxaqfzsN4pvlqVxgT3xrT16nq1B6
sWejo2d693Cvr/SLaXqKLM+xlBpi5/LaSbTDhCBKj0GdsOJzU0DCfPoeEddupnQm
tDGEeUkUaZG+iF3UaBtuM15cCIzQO62zxZtCPY9/aXzjigVanleDML8L7NapdqPr
WwbsGs8hVQY0RpRCP39O1vOAqLpb9N7IiIhxEBbBDHUdjNYyq2a2DsBeVZIUnzH1
VZUjBaLXURo5A9VhuGWVUV3T3PrfR2lsrb+3wgXoalMhK9UN4Mrls/IV3dGWIYwQ
h4z+wmqb5i7T1ZF68CdwpEC3bX6zSFQDDAPfCzseXcNEuKu50qhwmB4WStjhCgy6
U8urUPkhDuNc1Gt0HxedJnqOT7vMh5ZZqrZS0R2S/J18mfB53/rAC5d42oUzBCcn
0LjJ/TzOi+y9ow7ATTpTt4aCp+xb1KCVGXWh2ryfBmxGWM6k8tbTi/jPgRKlQBK5
1+Agplzaa+LI1g9SEMPGZw6ZQxWvIU3lUAT2myNBZNCf88ze30h1CpQuarOY7oQ0
/rCuO0UutsGQA0dkaE3RUlbtk3Ad2Sri21qVPli5mBoY0h6VkCCFGTYDvnfZW7rW
wbKHWdtZiKFUHGI4/pNL6DEaHOMU/dAjZy+XDT9XW8a9/cAnN6U/GHoS9FbSYV4f
xPJIQvYkc8xvQEGcWnAuGNQ+D+0THErQsPiNpwKXLKKxJfsxvOJvPLp2kuLqqYnU
QzeXSiI5ECKYM/Slr9ogxeVZ5ZycoLvSoZl9BvsMgoJQjfDD3ytsNFbpFnmWR3o/
VavFO4JEJ1Q3HVCxFltdOUrUhMlTuMxj5vShPgfWJfiwflVQde5HecZh5AAUc0CO
7ksK20oM9Tk/AqRA27dK2JxHD/o15T9Lbjj4lEcj4jkxNCCS/ZpUhBKDwXJY09/2
/RoJ47nMjO2l7j2h12gyKdgd2uGQpecmtCi5V5rKPus56RrD7CHhetmAB+wkDc/w
2mGdxwgOOi7A4jAqOcZvTWQMu6ObZOXbdBnZxCTQKLWKL3C0qrNFo7PUcdjSO/lG
NXWIY+9OffIP5qkQCMYqZ99iKuoRdSFI6r+3Ttcjt/jEiIu7IKCJ5JGRotRr+gpj
ZQJF5VCRZwY3zETc9BOSuBjbVKg5jakWdYCBjN20gWi5b526r5AIvFChwvzaRHfB
k2ZKLFQgw9V4N/shiwQe9CMag9f4g/n8Fs5D3n3I6xz2pl9VwaZZMtprkVY+RdOy
3ay+beRFBlRempkRDeYpLxw3MKWK2hq23VUPNhHm0bfmo5OebN4uziZwfqyT83/k
ISqWqLQUYj4bpQbFmMuixkinVEQ5eEAZxiXHyQc3hVdXB+0OahrQvnstsiWTtm6+
bQkYqqOmL3n3rWW3L9KuqnaLguCdX30aXOhwFCTliz7nAfGmRog/zjkcOYVapbfl
VL83B5ZxcUxrXALeVcqBjUWo9nJygXMazm4Al0rYjXtEOp3ZcEy9GjfTs7uqFhCk
NXXbOQLjjQBjBC9pTcVYht2jopQZg4v/mjrRGivAbUtzKNaejQnw4EoRM504ypk9
v/guHkZF6z8URTXxq/qWcq43qYAHdRuxi2mBJfe++Qk9sn4UhWlH2QJT04CUxHmP
KXvnQtHJQjaTl3EyT/CIKjVnv8/hM0yFS6Jw5OHuVw6O/m6HxzDdXttjZlxBR2nI
zlerR58LBuqAgaTtiit3gueJxGAJj1Mrlpw2/TYmZsg+6Ut2xQp9FYCjt05UfA34
7n3uwtu0TTnkOz/74IbSiZE1hjfdTMmSgWRqSZ6gtWQ1iY75hnzIq9juzR7xziFk
rYeo02+6Tg4gZuqya13wkL78PyuGRF8KB1NoWoEMdmRXRE6znmyRPgUQEBQfKKkM
etFPKMZYwKiZ7zGuRCJ48wp2ao/Z82Lhb9XyU8YYw3v/vFEhMC7t8KfccniNPnKj
AWtF0W0TsjKUUgwIQdKQfGNoBNYu5T9BkC5e1dbWbp0gT3utpd8MbL6bh8gCZjOG
XR9BPoWc2qeo5JjasVxzw9Cl5mPhW4IWkzxenXkK8kADx9a9E0iZsiS9Cs+9d1AQ
sTiBaPjaDoDACz8YPsy4nSJN1o8wbI5Mx+sRP9DWO73obgqQNBG22Kil9NZHYkeS
L0J8vRJCxO8nYJRGAB5iYUC05/MsCv8Vdi4hD6vMfZcE8H2u0EHxbo0bcYzZPGEh
mqjPTWN7X4pgJhYV8fiaQAVJ3nDiVkTun9YIq6qlPT3LBUc9TYLTwC0exrXLS4ED
d8HeGuYR05O1felRIxB414yez5zW0YqrB2OVQByDkeemSC9CSW6gHFr/DKc1tffq
gce4z6YR1yZKxlszVD7rUeQkjZh/5WLUB+CDaMz0wi0z81wHfBS9AdCtps8h3pxt
oPZRD3weLWuzN6nYw5iNmi8bdHEOsu24rEm2BXWZ2zjn1UPu+spm+ksYPty1DFRv
CeM+JGGtusNP6aoaghfFYmyS3ATNwMomArLbtMxk+5Sem2VvE6EMLuiQkpQsyWMf
4538r0PmCRYG6aS6f5aThjenE4O35IcY4mCecUCne6C6IXx5X6/PzciUEpCvsGuH
EA8O6+Kugk/rs4t+ZzOmbPQsdLeUnIuvwtj68jKMY0Qp7ZkUFERMZzIEIxC/CXfL
o3qEDrYrcvt8h9jEVZoCiLVDXI025/cIwalMUJZeAj7N5yvbE3zcTY9oWbDiOfNd
C7PwvVr3yxLOQAr4XtfxU6zhlfwjchLjoVxh+TnZ8oTk2tGMcA0PPCjZ+C0oTPP1
ip7dQ+6sAK3FA4An2YnRZnkMfho7Ju72OuQ17xea3iHNo7nwA3RGzPGI/Oq569VI
/1i/JJVuVa+yEC8Eu+usgfttkwSUAEVtzGFIXE58GPDAV3dBJQ9TIllJewcbYm3B
csUVxv4zoA5y2WS3WFziIhu1Mlq8tZfu8aky3f71edeb8V5XdrNAQNcYMtPyxL3q
fhL3OyuCfm0kMAHB19iAxT2ZFEpisbC6LYzo+58OSVaysZWmNIpWpVvUEpfyP1TO
8BSlVxaXv5/LhtfX6hk9aiyA1EKRXzPoCZpWs0s8l+qY7aQZVLb+yiFFGAjYmQ2T
mysTN/5nfQ9d7WujazYTSfMIzMypUd/HXp5Js8JuHvo34ao6b4zaFoFUycPqtmyl
CXA8/cPVpxMpXhfomY5K6F/djPt+2D+T7ZcCb1YiUAol51oMOtGc25VR5Aqyxlor
pzG6cUBI7RV3FZNZOqWzGtRz2zrBlXAnF7OBTVF0CGTu3hw0AjmqAS+xUq7CHgmm
brhJUMV2MZT+8l8Iil+ItJfus8YNA+3PN7ltnQhWAWiuTAOlK12zr/9XK3SenigO
PGl9OAboV098ENJ/brCJ4pwhreWn2QXjn+1MtfqrFePWfGwyfifDeJV/1csWd1+i
pnAm7id7LEW5k1l5eySFdP2N4GWg0tLd5E/nc24tVp5ibm4tystxV+0bz6jgfd7G
sSN3YgsjaIX2IaumWpCbGA4eNWQE64qoO9XYn+NL+jqem7k59yOX7BT7r3B3RuPg
AmjiQ1kTZ+sAqAvSzpXzSIyoLg4+bwZEvmAnPpft6zLOay2UAeChy8QAzYdchTWL
6QKLPc1d1m0MFe32t596S0opfUoIfxlkXvak+1idc5DGGLU05weHTyrHU7q/D+VK
PHA4VZAYMmxWIISdJRRbwm5d5Rk/UJhzcykdxWoN0yUt3+98gY2Mo++Apyzpe2H+
8WxZElDSmQqPnflJw95X1eEJh2Dm3ReQWEg5KPfUjmTQNeW+IeJjcUUCW4UdmF9c
sSYMdB3Pw6tEo1euc1fqTVULxv62NhwaGFDUac+ACY91eLiZ0LMbMgU5VyzB9R23
oeuWI+vXPvZCS8RqevYcldU65SyT7xwY4ZNYBERTuwODUcyZEeze6NmJ99YK/RR4
HAaWcMLcqKTQPO+uicFgip+L+/4o0qt2QMOYi4sI5r5aWRCLpxyLZhtU3e++xu1X
pvsmJ+AZC/tgqhaYNnNpf3RnWUg0dfb7joFtO6Ow7+/d5fknp9RFemWgmjvWslYB
eldnaTZF34AdgSklY21wO5znSgOo0YFc6n83OY/cma8RAVZRyUd+JveAOkQEYCjX
wiCdf5Ces9zjL7IIeRzlzj2Ze/ag9XV/DOO1B1t28hQJds74k2C3apKQgef6mp9n
qaIJ84xMizhybPmfgCIHW9L5ZuKEzWXTqPCo86E4TOmBr1GpEBLX5k2Ppuetn3WH
Rxg3k2wSFARDmcBtABXYFDoPzm6UHy3OAGr0tFzko3fSEfgcDXohN/ueToC8o7DU
Otyjri+vR99RjhVyuBMKrqMIz28e+GQLseV3JbUii1ZOZfuBCHNDxjbn7CmBb4rv
VwxKmQVNG77ayzVC69zsff4w6xC6TRWWXoNhgVb5tdTo7DlRe0T+tHGvP/oOEcUU
v4eg3cTvH03h7hpBFdvCPt/K7RKkvjG4jdStLxbB+BoD52YVWq4QlUp5TZvGAyzY
VDrHygiART3OgPipPuoB8PT3OZiLfP/IilVMhDztm+lbq748Hf25LbJtacTDD1C+
/YmhhTXN/9pxnXbJrXMlKzllZBU5/qelHU9lDV8q/nSep0wqh4H060AQS8Bo6STA
sTGGtMpq8dlw/hP+SgEO0gxwOIzQyEx9FF49ijmTJCYnD3aNA/r4h43lYC4PfzBG
9hjNytbcUI3m79l9+NbHRFRpLjNrg3QdLpyYT4p89tKchNMoNYg2ZRe3zlC4aHOS
HMa6sUHeLzbSRdvCFC+S6jGQr8dVP+stDsgl1tR1Ea+ksuDMqYy7b8+eYSmEerLI
AQUitzXWwJkqFqqd8R3r6tqNszvdEbJxEodL2sQnp9Fj08uPnYrRQZxlyPH2z3CB
QAiedvbLtoTS4WMsT0jXjhIx2ad7s4/E2BPAj7OY/yhbTNEzq8dMqjUllIRu5N3q
4jZIBsWJIzoad2PjdykcSAANqG4uRBA5FNFBvJFHfDlFawesed5/dIm4mtKoRjy5
MihyHbuUpf5RuFYJ6ny1HcW4g0/bwrnjUnq+dEFRK80GrrUH3jI0s1nohD2sSgab
9BKSq2oqJK2Xt6HWwLlgE47rC0cirqIeGFzRwAZxZBxsfzOhinzoXDoqrvURCT7y
O9DbRaXcITM95mDEYd9yq3tTJLF+dt02pGS+yeaQrc8yLdsYRaYJU0lzYjcHz5yz
w1AqGH5REAkFaGSQK8AX/xO85W6uJrFmpduV80p+PfQN+jp0I3ieBXf14Md/Vjbx
+doTn1pQU+hG82PYuzpdO4av2ZL8j6nQGsKKySR5LOsfnM0MMstNz/R6WUmsVCud
3YF+YahinTSl3F6wv9HNm2dmUhlZpIVbUc8rpaC0QSebNwCfY7Gh7r1tgqFaBzaf
bJfQwSks1BObqIdlYcUszL55PL5Jrj2fBXF/7scJeoCm7s4OXLDigknszt3jHsdn
WGVF5TeuzxLZV4yReaIV8vscaellDRZvsqea4RiCaw+UPQEWvv2TxiiMZqRcg1ZU
3YvhGYvFq8jzPG0oTKx/T67F7rWFDyYVOCqNuoIa4njuWo2kFY2njVeDHzap7R5H
zL+YIhTiOvkFTEGPb5Bi73oUIRLxOnPPxFvxbP2tGxYUaRViH9y7qzApftlMJhSh
Csg20+O0N2lqtZx5FpvwK0MKZUHOImEJj1hnMy2HY4nnKTUdfRMo1hqg4LZtpbu0
xzQTyUI2SUL1XkU24oct6TVoSh7AQvoHi+Om1Mqj6wkk6PgE/ebAILZgCgTMuV53
yQzWzpycv9LUnku6ZaVRRV7jj1n+owVhRWXtyLkVVBfa66vsnn2ZYfkvpNZ57fFQ
w7uz0PT4eUuPPArw9GXqzMSy40pT8QM6vpAizBNadfUCJN+l5SjfJT1Bc+7lqOfs
XNaqmUd0oFbAFvSD+/yPzwezOLo/5EpGFN3QSDIKKBuuq+I7Pf+CSvc/hU/vjXeG
6cjLAkKGlE18msPwNl06JUa5a81VUnlqrMyzW9KHNM9Spa/3UQzGKCi3zyDsk13z
FhEfFPvqS5A+8p1r2+y85wf2QhnyJD2H4pteOuJVgAXua+Ark9iplwQIAaxqPfud
gdircpWaHoM6QSEJqQkOpdf6Xte98TajSOoyasbVFjI3Ab++6ya1Lji6z5rSrbSD
2w/7nZwnTOKO/uwy6gJMQnDKCWtOwCqUrA1+4DCmCmvp9wpg3OVNnR264HWKQAt4
bJOBaeR+GfiVQYVgMLKBkz5p6N+JQmYfO0xaNPKgCoBC/Wa56OuUDzAcB1C7P5AJ
J0tsQy9tgSL52Bjtb7Jg1/OetSj577Pns+nStq/UiCaIp3AkevbjLJQaRMy6KdVm
nuPcwi/UTNQZZS2WSxl+zNj26p0WBbUbVbqnTPgNS/d9V67RcPyxKldhcmh25Qlq
UXXbROWIUfVC3B6XVyG5o1huxuTzakdBXvvMAhDGNEdtkceIo1rkTlvCwH8ke25q
i3n/25s+1uH8bwF8xsTfEjreLn4ovAt5CpS87plkT1eGsgQHPEDKpzvdHB4219Vd
2uyeuvhPovRIDa4RaT52FQQUW2NfRSUuHicRHPtQvk9Txz7npIYbGolLHtvXMFMt
lPb+9xc65C1T11zykLjZTMtUQAcyUFZt0xphtryYZOLA7Fcbabp/8Wt5td+PyL4J
TTnNJc07eW+shHQel+sg3FOM8PcW8JWgoC839zXDjJhkwbVo3G+I0hp0HTLBofyO
ks36FO5yMbP0aKrpnD57Ia/kBk8luJxJPItLsXIxo4Hdv56vQphiPBnNVSearROk
2iIqad0U68bL700PJ6gHgEe0B8PlvooY1eKJAcrd4rYvktebAZceMxiwDugmGKzX
5iY/ORPhyXze1nNObxEYpcc//SuSGDiI+pD2S1eK9eGpTAqtyeySObjwvwzGNxMw
QsKEHL5lGvoex4u9oun/EuBTLk47a1bO1Z3FcHDDOfwTWCiBEj3ahGXKZHAOKkTu
gJpfClsoeLdffFVxjxmxXx7LUytM6gpZMX58361MiJ4/p4SrfYM4RAlxBt2lDhyf
B53f9AnB5qIX1K0Ag8WWnDI81LPZWkjgE7Zloawr2AnGgTje9pEVEINxMkl7iFsz
KIuzd4XMBaPfWCBbaaJbJtG+JdWz4vVV5LFn38uCdtdSsLY/lOg6CrnGbJr8tIKK
HmgN/gZPfRmclYjmJLesZ6qkPHb2LQU9IkRry/7IlNSN0y/9+rc81bEUyw4e85Co
WImDkms4CqTPKIklPEsMnzCYeQJnRDTqNmLrPCMXvk8uRaSS6SC3oPjQYI3+c2g0
mBTQmaMbEF8ri1um4q92pmVjEqOiuBJxgEdQXSX33cYg+AkaA2zA4jHDlRiiIDzZ
nRaOteZfDMJ12ddSoxZZmyDjUGlY9yRq1o2RZoFOg0iB2soRs/SXi5rvd8uARC7v
9VrM7SqxGSl00OQrG0D5MnoeZmrHb0huSIXyd0CueRmLWulFQNLNVPMElWDzp+Hs
oe1mtG7jinEP37az5vd4gDfiFfcdajPzpUsVqu5GNnyjzLMGNjyPzqCM2eldeEOD
FAj0Ro5suAW3XH1bDVziZwncKmqwa7Fz7Mpz44mAeLEl6Pg6I7HJe2YNgxFUKb48
W2HE+ifF0yD7BxyjLGgOncjg3VJ7q9A6SYuDbDIygLGNE6V00+DqFQ/QBtVZVU3k
jfphs4lRDbaJaCcLqQCcSCq4mLFyJuX7p02jq5+mT5N9g8uE2WkrT9sW42KHaZvK
bZDhjbiqfGlR4wW2BEMLmk0q8SAgin30/fpMg+oNFY94xun8MVuKuHPE9aP/vk+l
JdU/Uw9v85TclD35LELJI+ugdtxFE8I0RGb97Fgf8nraMm5wmR6g/FMCNXT7znmV
D/wCOGL4iKlYhIEiCX9glIj4utFkXmyeehqOXkUJ3fGsRqReX6UYOXoy5e5hGfDS
KSrLUu+5Plt4cqCYXYpPJUpbc/zvJ7obRTk5aoRY0faCcjhQOtO+V+u3HmzWKHZN
5ZoFvZ6RIoGX/f4cWfxiDLBJ287+32VTnkf7W09cC3eGYvpSqU0BL91AypKjsKZg
DjjePPLxWPF/MQ4eAngLlRKqO38l6H9+cQdfyQ2q5QKxYMUJJUrrU0SoHgxS0ZkI
gu1E3qrlEzRdTMWF0y55o1Id7zEhZkStRxA8PkRWuE6eH8FO3MfmD2csXp5gh+Sg
5CalTlROz7l2N46m92cMmFM0aLKfich/Ybv6BX4i2HgcPJuH8dCfKvW24+q0zz4t
XuZSZB1xk7uJHa+E8/I7KKBFov+h9UEVeJqRmP6bhzW/pjMnn+KcyPlstuzBzmZH
jR7MH+V4fYsDywzuB1OfqoHnTxYDgbWPucNuqtrt6pQzuBx+Pu80Bl8s3NhhS/Ja
lB86rg51I7OCUP4SVPrJC3Cg6SulE8NJz6grpGQutdEK/XEuZqTW8S+uOoMYdXzp
B4iftkiLMWfoENzg3snTnEZJWzTUfqACVxRECWgU/ZkSYiqqD7m18f0CDfQ60tYW
wCAlo9KAvY2zgSkJvmkw1BChfncWOkv1oJdoF2qBwTV5aaV7YLt0Zc9fswaZUEkF
aIfoMNlDFoUg4YLjdTvNIbHeIxfragJgTOydIcMcFqWDPjVHeu9hsLEuBsIXalyA
m3IdEy8DFjeJS8F69Y7hd/MfSbinQfV9nrw5atM5RjBJyUXyk1XfsVelhDDFtsMU
yZOFykBlQaN6B7hkXoubQ9KUU6U3K/71XTBb3jQFWQvELedwu671aUO30TsA9Trn
ZPPEjtkvbbr2nwRdDpCfiFOuBmLT0YwmYTngpxKPIXy6lVJhbm2Hrium3vXe+4z9
4NeEJbno3C+/ZE0bTOR+zBDrdYVXsCq/y6hpjMT1az6aCJURb0/+5rwmqv+NsgOQ
rkdV8NrtF0nrSnWFzU2bkabeMLpSFF239r1RS5TlgIeIyuOIIIuQ0VDEw+h+STMw
cHb3kSPUkHqbks/4l5noY+yuVQ3kPoKuEQNhSswdbFdRRWzAHyaH1ETW3f8kUM5U
2mce+Paqq0QR0JwW2BqRpd4UdtIVISDv4uOis6qveFIB3YSdI+RYmc8Z3eL+YV4w
P9uPeU0pSJuQiRtpqoRjJ1PfOGZhdLCQwMQ3AnCFhd7cS12Ko1oeIj0jJbeccDHJ
nb34k/ZFB7761URLCe6uNEomjAcRPPaufyheeocPXNK1jVe7/M/tA7nqjInpRl2s
CfqzRBTxAM2DQC8nnDxXFyNgw2zKijAJoNKlPYirgJEvwDwIGxdda0K/EiELYJrj
bmSk46v6WNksyRwpcSoKv18ihC3UhJjVO1iqmbHGJbx5FD0AaXRxRdQ8NtiPOpZM
nazwhCsiWPl1jTSxFK86NIWlph+P8u2P5kPUikw1Av1d+sWP8qMRgaAJMvpiVzqA
1W0SGk95XR9eqFWdOfkiNed4xtS6GK3HUrjvoZwHXpBVSV1XK71mOF5OhToEBANm
N8z6Qngi+YS2ChN3XQjCTzwO9iFxhLUbrbzWvpKVngY8A353RYK0uHgvMxrhcoEn
FdcTcQbBDz9rZvdkX4mntClRh/m2+14ZGRlqaMIqTb6BV/dkCXCuaDkIpoGh0aKe
MWSoI09XU3XoYDezc65YErWZQsdWOAdBcWt5tQKydvj0C670FZ1LdD7mQrLtrpM7
iRA2bprGwaxkHlaW2pNCOGe7Fg5tzQt0lDaACwNxGJs2K3i0MRmr8QyxGH4zQKrI
CZurqW9gRxc8+9Bn6Ki+nTusnXDYBzZ0+8CrY7oKmKbSrqr3a2GUJPyu8a4roG6H
ba6RQcR0DZAime3PlbYFVZ0xR9ito6rbhXHnp+R6efP7mJY5ojDqV7yzVGeOrTEB
Uaxa+YS4OWmBgBFXXb2Upozs4Q+Po+G///l/xEl3kCz86QwhQo5xBuRN6x5XDnr2
jPF6pT6gAyw774/SR7sNELY/6bopH6QkDFE4xw7JFPiW1lFpJZYdYJ8dCcKMBk/v
uUwRvhtN9TVm07bvgiqIeIIK9rC63T8YEdAbbxdobQMrX+eITyGnUY6nUeoaLtti
GGeCcgKMIXIwOt47eaYfI1egDWvk3EL/GQlGH+1rfULsZuKlBjxwbA1L18O7ItwP
sEjOEJlHoCNBy5JnTP9ox1HE0Oa9W/pdoVeHxqJNU2ZkktO80n4a2IU/7EYTtikw
aLXgmRowoRlc1L3ArQSBsKDF5q78YYq7QJWD6l5Z7A+uYBQVPmvU6LupC+enPnpo
J25gaRCahPMmi0vt+QrbgyVTTq4n+UaKrwuNSz7douSdzZyz8cNVuJ9N2mEBSUhA
6Ts73NLfZCrMv3J/4TJvEzpRqN4MymdaWcIy78rg3M7ryRBJfXR5ugiIhKqb3vks
cSsyxEIHC/bkIEZUzGwWXl3g3xT6gsTN2VS+dBM+I7g7jnQxN5AGDUXWHqMA5/l9
p2Jdfrll4aLXUA+Km3Bb575rUgysYHF9gicjzt2wYOt9dKs5ms0iJuudyySFkVyU
hWjzBed5y5LHtoKQXFCPTtRPNZ12HoLIwyBxi4WOKlLNsAMNjeXYMb947sYIY1I1
qzpN0EL40STnWn8pC3YyUfDC8sakqIXPw/U40MwYtgMWBH+0UtPazzCSHdqJRqxw
FFP45B8U5EIXu9PcTbRc2A5mM29kKX/Qu+fi0YC6Le5E19OIAMYOYnR5H5zKEB0k
nKLGXP04Ejw+KADRgoVle/FAZt9z9I2rnEn8KSJ8NPLF4arMyO3PJxF/OWMz8s9V
shDZyZTqSlIdc1ofws8jTWqxdQiA7r6h+GoSCEikfG/6mq8Bed0nH/EsciLcDw2b
2leytBuIFYEaFtYqE0sili8bbYLS2UuaB8MOY/BZBqkHvhvoYUSvXXey37hQq0nZ
RSV/EfmJ9aC4c29nqLOrUBFrHxGr9/qlA3gGP8Ra3PCPjKtUfWK93yepuIvrtKkP
BQAVe73DAwVLEKVyHwrWPTXM/sSrTLiZQA4IW3kaDArGf5T6ikGxp1cdPVH+h6Ey
0Ckd+knsfefoEfRAsrvOddgfgyoHayaHZX+Q8yEEIeMep0P6cSmUO/Bh559Csa70
rpTVDJ9J9tYQ/MRg9DVngAL3tv7gw8INLHNh/EYHEu7DcNaq+NVc8Ls6Px4sIHtw
yQf3KKvlsxGBdjQx7G+ne3O6atkEcPmLSVm39a4hzDssC+F775l9lpjfJzCtlxas
zQxySWWTNBy9ic8j+ZFxL/fuK0EfzQ01pyU8IlNoHxE4vUADQU75FqIeOXGHiW4l
3p2/FaOnpepmYBrGMsVnJZHD5ODpe0b0LswNXuz0Qg1z2PIp2YxXEKB8kKGu4YLi
IS+vbWYoP9SzLuBqcoOw1idXUkWCWQ/oQL5G7Xm9xUkheITzT1NnNVE8nAd5zjln
kdhRZQpsw87v4MGe3VbBS8odzc/xpinBaRsv1JlVZRCK5qljCyNzbb+hsiFTH8n1
tUXP351HKtVau8PKjneivtvtUzE7+jYElH+ikFh/1vUMQxZuCc3IgjY31HutVOYs
BWD2WS1+/a24nYiDOsF2NYQw3nyWKcGYcGUma1bFp42cz5WU7wMqQoF00g5rGH1T
6xzHxJjQmwaJTiERU2aVCwawiOEzpMNcOKCdSl/3H/ehepMK6EgMBuU4sdtNR00O
woGv4FsUKBuEVPb7+0A8Lx+AORRTuesodpfUWrP5+j8+eo9+Zc2Z6+QxpZjPgut5
X7Rix+fC/BHiqRow6I7jv4a0EqaOtY/wEEYApFt8jz/Uf5zeh90FLDF/DTVhBuOS
6Da1MJnFzQBHIct3TZNW8Dlg2ewYtrsmY3pLlVDcD8yao5KJjmnYkvoZJ1RpPwqp
ilUTH+x6wCA/5rkd90EAOZPS/vsd61Fv+1c9Owr7DLWkgByjEtF10yQaNMj+eTty
ZYZbosVIpu73Q7xJas1zmMDqtUhGbBBzQWLEPGaFC9rI9twdO6VnUHaW80TvBvU4
Y7DV72kGMgjj+a0SCEmHFpquVX5vEYfSx7dXBLw83uXRFd0mafnVRRh2fWgOuaD8
ikIdqAnt+R73uIJg2q+HDYS+oXufbCkUjJQaW2EGCwhIMV0+1truYNP61xtN3gYp
myBe9HNZi5YTJJjmjahMhsMk45eEPAtVKNETa8isrhHICeocdslzdASzZ7/zHiqC
JSDi3sQC1Q6sXY4SM0HQwSqaM10tGmGidvKINVA7W+2X+ZZ0lnYCoUdqY6fDtz+7
BqXT9jRbCEAK6z6adgIYgi0oJgxOaZnnwF+7RyiE1yqU/tb/7tLTvmKJfPAkOQ/9
xf8eYLyBO/++vIPa+m8AFsQG0RJn+0zpZ5QkSd0qrUel/uvmq6hlbYf+mXjgg3jM
VaMoBrcc077fwSRSlJWLBqVbxGh79A0m2q24wroDKzHezGGEMgU3b1Cw5jEy8nxt
QRWk77UonMU2IhapZm3ji3s1Lf+o5Ip1M3cLT2kKAyNiN8cLm0sLiBcZfDPfFU4v
etPIUBVf+PTfk/En/HWfdf3DoVAA6h4hKGk9141+fDOo2sG85UsUcZhfsOQcoqPC
PbGsEukmzhcao4jGhkd2Fpj9ha8CM6QKLi61zNgalVDWXb8YACBOXoSsXPKULs7C
knXQZR3++UNKnplUoK/YUgQckCJ7PlOr/HqjOlwi4gtf68tOwyeXzvdYET+VJQy3
saSAmMQl5CMjIsROXC9Oa/ipqaYQCd2FRxOQphfc27s7xz/ZLKt+mTDrEMePXTwD
rL1pfKaX/koE0FMucb0/eBZZ37txVPTtUro2uFOXC4Fh2PZ0AFifN1DdPshx4Kpt
7coCyNqqZe2Q4rPvhQL0fYBlNwRf7jwDOBxIPqLCuvQb9VZqcOxhvPG662OVGG+N
hw1ArpJGJd7IuvTQcoB7YblwB8B4n+501CCmXteUYUpP6k+A8CUcaDIrJkkGWPC3
qUmm/rrsHRkHA3WdtV3Jaz6FNNPGdE2BEgofhFtoaRrUaWw8bTxTMmIi9Md89ie7
C3pC89VlH3Kd6GUFd+76xSmr8gVCYeTNU/WytIyWL1c462RSidvisEP6V3yJyC3M
oMIlZlKpd+wP1TAkKPvgYyD9BmLq3wWtc0uB5AzWQ5+KU/XzFaowvfakIvWJfvWn
MoYGc8522vxwlp88v4BsucrNKsrEgSvPGgvpQsL+K3XCqfn7vZCdMECQDWo0pS7x
0F49ZAHkOIXekZZSCo4+C6oB82y6wlhQYdvm2IPLE4XjgJktAcP89hPINpmNbs43
THeU9MrK1H8SS/2BG872pgWc9qHiu/vvMCjvz3h4DYn5Ua/qZgJpeZ8vHM9wlZEf
djGY3InwUYxzewbuRg02OXLGWvA8kGzftbf6HobS8Wja+pzGdlPfHEjuej6RA6Ae
k/y9RIW3WAAVMyfoX4Z925TWcupdMsU1t/5XlYPfRi7DJ34/NmkWUIywljOt2+Vv
34MlS8BX2WdWaitOkzifiiZuLXYlSpr84UG3C9FV2oIouFwAbljFAXHJ2ilmt2XG
xE63TjxqUmMT6vm8BdYoCPeuDsxCbBItE3W0R4FPDtBghXs9n3jeQjfsN1negn+w
l6rnz7NVOlnYLXJ2bZCpLp4aY48nUwV2yqU5/J6daOHuZ/fI+We56bDAJxp/7HQ0
whkN6STUxGwdb9U/jW6IkEIgw5b8yhHQghk09O2sO0cFw0k4jq4zUjbN7OtY80oW
nfhq5yAUTYn4grAia+YxHjNzlIREfxzFtcaR0oBemyRYy3hk/2KiGGnZYCeKW9MQ
qbiwUSAA014a+rj6Prgt11crtJKwaxwUDnX5REguYFEJTTSSJmmba04FGlMIMpQ2
ZUYBhZN0ziuBrecDun+0tI9pfRT2gpz2i+s1dqdTwDpP1Xpr+PaVmpVJ5FGHBZ/l
Uzyzr4Gm49t6sXwQEZi7+4xuVu9lZXX2z5NUWOBOPv+zf31LGbkBA9cL5aXp9OcK
BKv0PxtgWnzDlk+e6GsbLHH6znhU2XUo01gzrEERnPRUy2L7hx/NFrVIdQMuDGlu
XWfi7PONFVm/1P3mji/j+0pFMNOaQB1NWthmUOF5N67Axw0JFV+y+2lkl/VVlaum
QhJciYh6ygtcH8xTbcbSjo4QPgLcmsyECQbUefMDB4Yy3Wlk1KW36LU8X9F/T4pF
Bpv6KzOpttt6NZA7gtjZzwjmepmJycIvvr+aXPZAh20lwriaiF8+ljFP8KDNyVze
yQwjZBluPuiRGBJrrXwCb+DJ+b1E1HOeBd8x8tWMw1xyoB2FVDB3Sn5fufwYFsX6
BlBVPav6R0dHNZY4/7NXACkXCCzwb+lAChmDqNwQbqhIPd0kqLMVosFN998Tbt99
Kph+iz/zkMTL2RArJfkUZywwNpXOuZRXtfUCjZ/lbXHc2fdNq8rJPuMSm47HNGem
tlZ/yJNaYn8HCIZKIemVfHMwVv63KnSijrMdH38P+yRX/gATaafNxsvQE0abZvjk
tr6SWNT1lQNPDFAMYRIYN8blDxTVtB+gtZtz2QaziXCoNf99rb+kJuEElupHokG9
mXqzuD6E/9IVkw+fKNQG59PVCA9OaGJF0PQ4gqk308qVIQeKpP9yJv93T/JWexQu
BhFCllhYeY2nIwxTcVD6EoWbXySgN1MwnIMgP6C5/RcjsBiuthiLp2Va71VyEvzM
Vc+Q/IEiU2LvGfffIanYOj5j0rnxVWLIX5byd82AvSkeJ8vZZEWg8mBU5sr20S4T
l1K1Ql8D94toY9gJy8oifYOzFuDTf0jZeYaWuddKksJ0t2WHcsO21RLqgRf9BIB0
V2d3gcJqG+5oxldchfw0MhvgQwHc11CAYZgXkh0e803gT9kwkcHHTpCvUX93pkJV
g9ex+PAvNMA/TZPgUhWBtiXEOwsqTmY8U4Oyp3sqfId0eb+NWN/7YQZ/mGEg6A96
Oin8zq+XnewLu30r/A6KrDEUj7N8qKRc7uy2r5UxbcOX4HN87JAvgyJY+BKEZJVR
Oo0fkprrYJ6UgJfD3SAcqIhH1PzY8NzcCRStru/1bRXYMogdo4kznBQESmtjDV82
UCz8iBi5YOMrYPENf3GaQCqSOdxtVEVWtNt0Aof4AqkNHBbxorGAHjztgPRcRWsk
6SSEYtLrkUt4K3wXYOsAQtMWXQsCBywX/1+WdufY54k0zi1oBii0O7IQy94yiqwX
WNf9DHqxgNik9liHSST87a5d55ZFTuFhaVO9106dq5w0lz4Ql9jlyNhzEmuZiYF+
BpVS0GUlRRraVwMG3jgM5gcW2QujSzJNXsH5PYniS10dQbtzv4GfJzWwekfep9Rf
pW9fE7+ys6aFgpnN+R88MfRRbUFmjZ2wpD4G74UyzAzEwVZClzlQ3kByDJ/xVxA7
zualqsIWgBi5Q3MybL6vr5A92TueA/aZWPQv0MSdgW7NV0zMz5a124FTzT2WNnG7
yeA2i340g/KSKkD5EVvaNklUlDh/p/NV88h/If6LeMNgs8zIiIP9VbooEgGn3li3
2j14MVFdt/iw8v3iDdC35ZCtEb3Rpdr/fnoMnWeYvpH5gVEJr7WxeGkFkqaS4Sga
98V6u5K4m2K+GWg3imXsLdPRqNb2KjGfz2/M3+dn7RMyfuzcARD0OO/zRwUBjZnC
VP63I9vOiqek0GvlteSNLTy2vOIVijrgE2mf3wPlApyofho0YoHeDd3KMigRiLOf
bLE6TgzrwFONeeDeugH2sDIWP1ZH7PXahiApXfirRYumVCAozWN38d7pQh+dYCAO
6tjp/mctwdhF56W2Btyy8w+UHk1J1i2J4+AnnMTV454Mxsb+5nXVK+aWYeAuehCB
sJ7XSMm0zUiqBKjPeEXGV0BZyyffWjwV+48yX+SraZwAucY/Ltsx/nsPUsLrmg3q
KTOwOPyLwXJ8wy4MvBPY5O6aX29ko1DUcWI1PhKO8qRUXqAatWt5jpvVxU5LBWZX
v2x/e++Jlb0nyfunZcv2ksn+Y4J9hUZUFqfdhi49xoPX8rqY1cN7AbmJJCLtUvV2
06DY/aZTy6RGv4fIUZY2tcAXtUFQOpPEd75J/w2oN7oSWdBfV0kOgGpsLEaQ4GQx
8n3U2I8a6QRblYHJG4xKkzso059QIZLjlLnYB9fXtXR83cWFHks8LmQlO6PJH8lD
oMNT1uGZnKMkR0lx+SJPPuRdGnFE1IzVibIbUYD1r+gINImbEs+VtOgx84Hx8/uI
0XxxARq/43ACxnokmsJotKZXqlDNuHeGzp49c1Sve3VpSWSP5Jk6RxmJ0sN24azf
FNuzitm83oHj5joI0tHUf0OI9gNFogiYaADavmsyM0KE5gJ7qZmGPdXBfAXNu6So
tBI7R79xujOOjtWPGSd3ltZeVXj+u0lt0uQ21lKgcUGVqvE83uFbzSs4EpUJhePY
tXWAkMbpMH/CTn8vBpjrFkToZzC+f15tJ06QtEAUCZy+K+m49FbSZe1CXoawyOKa
G1+Wo87N+pslREhww9dSxeCJMloZJSpOonWYlIJY91aKHcvO+bRz0/ijrTuprpwm
8N51c6RjRkYHTdnbOb4m4gVudI7YeB5Rc4bheobVhs4sXHlxArKCwtUA5G0jA4hJ
mD4VVMPLzu4JW3/Mh2C41lC0x+zIc4bFVXy3AmZi7Al5mfYiSF+t3UtFgRga6UrJ
ee1X9x3BUMveTeL0fvkRfzM9NmLrC9eVks1FN41i53RVxtVKA7y/MujflMccPXlD
ChXtL9evk4w/ckwqv8yxRfMOVm3MWfSp/47P2E7ovNBXWO31b16hsKxsbW1PHuUE
Xo3fFMPh9m4CqrozRveicg3VkZdNas6oEN/PYAvLdFwhebItIxIROWfxrFmbYKl/
Y659zBkfFSwceISEsZmx+ovNp19cTHYw5g+jKNQjaQ91QFxpRZWRBgaauiN5zWod
YbX05zZeHiaXEFYb+oUpI9YiDZ7hV3DfdCi3zxazhxCJHe6Ft/7cAtNhR/236Y4U
xSz9F/hq0BLbq7Woj+v4sywhGytKD1Z8tbPfnxQiu7Y6UMArIC9qU1/QoUcIbRhB
PboMtO+HqT3zurghfCnNyYBVbFVpElRLJ8oVTl6x/anib/dN1SXvTZvvJby2kLEb
b0WbomyF8ydWNEwbJCm201PelUj8QCXMrcjdMSBlGNxI4LXcNMsCFNVyNGH23uZf
MrygaF7o4N6TtRpEsGZI6mRU8tGQbA5K90VrptqGAcKJG1i5RHPuECQ9oqy92q7Q
74X8XOY6b6u3cqnuzutu0DfyWxpRSQfOVec/oRFTpEX39Ddb+FoYM7jUeKS7+yt0
gbxDX4kNss9Xc2VJpLF3Eve3htwjDIIBDN37VZ2/2OTVTy8hcqR03hN0xyOWROc+
AXlnG4vLQuKe62eiSwHNQ3wWJZ5HqpTNT+CrrJyHfNryi4jojK/lWs/pYApKtZCo
OTyq0JkJir1f4cR/4zpYtbDmSy88KxSrY34GYds6zfmveyZ22c9TeH919u2f89yj
PLIICE/LafUUCIILk1sVZPEUMvHX0P/KDkZSMwFQkP5M3vCZ3a03oLTanU1MABkY
USPBctrCddDw0yejniQ+6KMHRPsVRgdjP79y+uV6R1CUHbgM1AY5adtbp7thdD8H
BCluHG8cqqWascERM7wTzqbJgGkaAJXa9CcTP7yWFP8kz3rOqDF6Y7bj2hYPJdqs
41IYXFFPpnacE5gb97sLkMBuaT7g4aO0HuSrxI8JvC1zrFFn6SQRS1RGnd+Fhci2
9jvbo7DNXIeCnmDVYryF4eIPTkxnkTA8L0ECeOgeBaMIP6Fw23djQd9Wp3AaWzt+
g407bH6wtzz/AsVMM71n3cTnPXySkIbIU5XP00JMv9iX72u4FtO/G/R5UDJEHw+L
qo3D6XFjvjI9KOzCgbTMHcDuZ8lrrm4jgw9JsNJiLLC5W92kQIC6VyAjRua+2ezX
k/AzRqIdCPzpk57LQEkXLb+uIHCn7yEV2aI2dDVlMB72jx1TgGBkGcTOQyWUOWri
lo5HqRcxi9L0M1eyL3+xXRn2Eh+a0x0xRwCE7XLshz0IJkvTH9MSI2YJ2iiZvc4m
SQ0Rh+7bGyiBhCqvLiDrN0mZJoRd5B153hFAfp+XRlv4J7c8cM7BILZcD73bKQOm
tDa6TpvG8DR+w9q1asDRboeNk7qdV/50jASDH16L8UNc/MZ8T2A0F4ffeWi08qUu
cZc0gesDNC4XbHnkBI6nGhiA9xd144xbhsLm1jZJCiteScNIFSR+NINB2mQLWyv2
BXRbqorgZJyWvMu4HvotPfw5gh41klSfOxy8mjxeVhTuYeFISCeXKqrL0aKs62om
wYmJvnYd+D9mB+uEWr5yuDFSa9/FIfBhxypY3nTrTIkFXNtp+W26DXd0m6CrPMg9
8nX8K2/m5vaIFlWYqiDFKHSbpapb1G6GBiyjfJhj413qoS9oEuTFPGaZIXDc+tJz
IeqaxlD+og6lGZgHjEefE9kldpMUOECXj3E09+ABr7hpnbArCnPa/NsoX2KU7zG2
NrSuNVZsMbGtgqGHE+LlYH8ottP8i3eWFOQ1ljkGhVu+OqyeE8SY8Fwtd9Y0HE5S
8YhoIwrB9Mk5Q3k1H+HlVTqKtN1VrCCjDeBov5OWmhE6O248UW8DARW6VcxVhDt3
cnzK8878uzFHVjLUZLBf5Y0mqPoYn/irn9xc1cHAP5b32X0XxrHmshDIDKTdnD5m
ToIn1S7BIcmq999+8G0LdTHp8Z+MnTlyN7UpZbwCQu8zG8h8CEBbbH7qS+vd5mND
IMC7NbyDY/OSLnV/4JnhtMUJ8+OixmmZAiejS7BmwW5yvvFbN0Jn9a5PVFYgYnop
BZQCrIuXOIPlv+24WFYpBqaNn+A1CU+C5gp6tcjzM0iVPY9hii+sWKH10x5JF1mn
DLEk7XRUt5cVT/f+Ie+0oHRIg2AHjYEgEx9VLFXWSw5qeEa6LxCx/naXfdYe2kgP
P4TieW2W80A7IIniqY2g5ZFV6wmL9qICF+6avOMCWD1uC1FRuKNcMmWdqPJGtw17
PJzwfOcHflD+WBTaGCs/V2MNq7AS3BJTOAjtjN238tGrdrX8SQBz9egCZKptOoqC
dZzEqjLaGKxUatIXy3cnBEdwJ4qJ2lnM6qPKP3O1hA60BY4RGaXfOUaVSlWj7c1F
8SsjZS6lKc8UhnUwfXRo08Qg80LDMVR02DSrmRjGDVNcMZfSC3joGUziDIG6AO/L
sA5OCQ9NgVAyUr+FLEWZ4JtwQ+Ufsqty5pORywstL+bab+ckf95b8xckjU3a/PhC
Sj/7vEvB/K9eX/HUPd1Y+bpYVUolGKUFJxHGWf8s9QNzKg0zKil5vU0ImxHH4Hp1
LdHE821+ApMvkV1cdY10UXAOOGjimaP0hL8o1ya58gMqoUBVvBSc68PiCojemvKs
uCFyA65jL8Hf1sIflNi8PhoeSKhOU9jqzus4xKDAulGP/lsKV//dVNaAWEeJ3QQI
NTHJAetXxtHga9NPizZYtSTAgp9tULrlc5HLHQkMrfZ9nMaSrxVWY9pwXxPG8RPS
ldGSaoLD85uRU6hZ168yx+YKfml+f11FluGTEKopOnxhdz1KBK6amsWKeB4AO2Do
WWufOa8tEvfQvYQz0KEC3k6UwWMZNnjuY0x77A85vizQsWdnFcpX8YntNbCihzai
JOaT87iov4vKYPJC3jMgmB07RemsIdtwoBefbcIR3s8+QkfE0tg7yEhdUbNZiArL
ak2T6HeB53uBVFvKZjMvVam5eBbvodMUNcv7a1SnUvm1KxSMcwu+mAHHKPPsYWMi
Gqs++GHGWla56QuZWaQlxVxKd1T8kztMqIAJm40I7zh3X4PgEpFX2rmradlX0H4D
R2nQFMVOGGk/yv6AXANzWGx4VHLD0VfjypaTnkYrY4+oAtX8d0psKXPvGTiPO3a1
pCru5HIrNTvESrmfJfEBty+pGsKpOwgqpxzdcbjtNSM8KGdHFJxJcrHWoansNgYx
CB3SwYNahY7A9Hfdy1QC1NfW04XLwZ/qEoNd5IxtMNdyzL9u28VyHY7Z1yiOHnHN
XpJ2UT8pccOX5+aqvwj+1O9LQaryLOIPG0gd3qJo2YzDnCmYQL/s11s0YAoGWCBm
ca+Cslb6WBtJoPEO/he0erlEdVODGClPy4YLQXroo2PU60FvsMKKpAaRsGZX9644
P3hRkradvzKPZh2/KJ0O+sajMn31N6mpYZIGFIiswTgGIgNHu4nnrZIBHxuYG7Uq
cKnso+y9UZofiv81mC1ayS651w/o/wx3gapBfSd7mJNUOuukaGYzAIqVt7MirWWz
kVSA/+PVsVlhTmyWw+RN5IevWYSps5rEi9A8fExi94SPU0KgvLULvMteaopzX9ec
ZOgNWNXeDZofxlfzxztNMlGC+zuP1QDDeMixPt4ydpu0u3RRwCyDKr2fBnVQbox4
JfzYcS70IPu7ICDyBgmp/iDpfzXq6R2eF0DLO/gtgW17h9/htYzA6NdZGdXbnwQQ
Wlm6r059t4826epNUPQQvTaIOZmDPYK2biEtHFFpYjBjJxBWlgPJFQ6aPZw3+SMp
03lX/JXJ4IK6vZ+fz+KdMIpeM7tQliVRv/Y6F1IjXBaDaCFUofo90ZxkFbHhID+G
VzzCQk8s3lUAaUc1Txqen7Z16QIkYOr5W/nn7spjnM5ojUM5dEFVxi1Nfs8vADo3
mxeh2ZZFZz4Jtd1btKOPG8Jt3Zr0Yj4orxS3FWXLhbqRSyBZTmSfkLKFp8v26MVu
TNUrhk75y3fllqiATgoX8ZlAaKNEg9CyuNrsckU3GtifMSUyCk05St2Qg8pJ3LCY
FsoZLnB37G7sBVxSpCHx2aCHUp14elnlxDH6jtDXsCnn4ZFSNKmoR+5wcIFmfOqa
l7o95DadVR6K925aVEQOcApEHxzlt76rfXZ+obbi+u/R662/bHWGedrD+ImyDpnS
hOglaN69vnM5eNQ+eryyO9h7dSXsHlQa4tlzj/0OM8K7AxsU//KHjkg6D0S49e5X
um0+Jbyj4RmLf7voWTz/KiNU26gEkCvN+9GINp9iD0vLeQv1ESUUy+Yd/ygzmYP2
2Bywt9SqKy3Gv3gcqVW4ydArb7x4/G7QbofAFWaXqNe2RBkoiaTopQ6EdB/Y5RfP
ui82j3nLtLnjxTCY8bChAx739+fo4zl4Q4d76CZrUWvnJuqURabPR/OSVDEW5GYG
1i6jJOkhFA3SCcZtmbOsP7Mfe1N+00QXBZNuHJcEjEgWxTnzWYVDuwuY975+U/I8
hcBW8+V4pm7ephuux34j3FgqGQPpux+J6pOZa2puMLYpw8St9U/QQL+RDqsttCJ1
IfZ3QYdEoXeYiRv6HR644g3AhInu59WvvcuMGP5LKSbQKC6EnXIUFIX3xT4xNeFE
FfhZve0MDr1dN6O/quSMMjQRB7In7fYcciN4eGPz4tZWCri8jrz4LGUDIWKL1mTj
DDaNvtRU1Qa3Hg3bTybv5rrH55JSkBdBSwF8APxmnDbHbaqQhXIbz607aKuNVgiB
NgXTtdH9wLj4tlyJtnlTGvOvlv9tRCUwejbfR2bEyyT+VBe6NQHNk29EtyAFYNPf
neGC3BjwnUuUUjRAmCmBXoP2zhH7tJr1xN6Lgr0JH2N9rnENs6e7+kWYY3sb5crs
gFC7LXJa92C5uMHLlHnk5L13jX8qksL7w3QgGOYBtORsq4Lzp9MaCmqPDAA/XvY/
mIt3vf+nXogRdzjJ/o5bAMd3o8PlnGa40Hd35pjXntxP8MUqaWSBgGRpKYrexHeT
xXXtxKgE77vmh53QFtDeTU9GNng6fhmw8xIKi86gfOx+COQkECIJvcVWemcF+LGH
2fRwbuHpzup3ZKgpNKBRbJs5XagdRb6c7uXN8/Q3kAB+UzG6NSZ/FxU31ELwYquG
d16z+q6RIHK+AqkjWkSAESDwXlqXwkr1x0VxwCqjyiqkJqwu+HymyOwqwH9pXnP/
AT+1aCPbNALE6D2OSKq0Orjglf1okRs21t+dbvIQDWphpOkdPAitpFMa0UaXDsRn
7Y1FK/GbAk2Y00CXjfBDPIwIa9e6JNYyJlzzOIquH69WmYpUw8IBIJVA4RWy4frq
RkRppco0vxeOgAklwlv+UfiQzDiXBsG/0DKkPCrCELdlPvJu3l0ACTrdB5dWJ3R3
TV+kjrPx1Mb+c3Gx8RQ/RzeUM/lQeT+K71ezW+iP9GJ+s5qR2VhJ+GjvBixabukq
CMQh+33U36VYNP0R5uyoMKT/Mw3dMI0fcPNAC4302urDfWdBBXFNr1cl6LRgjdPk
6ou2Bqx9GP6pIgpy/fATZC9WsxOpkv33Vp5MLgn2NNLn0oPmpAEtp6aDqsU6+yVV
JrXFWixBSr/d4uPQ/8FuPPSShOahyyGMB8mzlboeB46rU3M/6IwW581uoP1pzMvn
BlyZZhh0SCY3GaiK1dptNdwktme/qgffea43AmjH41LZ9j+Crn0jwr+MtRfnkX5L
uE8wQtPnJ7QH1wCbFGsCIv/k5PyMrKl58ZOxjqbtRvo8EoWeEVzalq8z0wArnc14
z9VCmmBRssL7eTTRH30XrDixYRbfNhogvC0KZii/lmorldy5MaZKa9YEwz1bZJCF
Nm3uAWzoDF2rDv9BJmo6dtXWoOVf1ECdj8DNR/QA2U3qqTOWlvCpfvog7U0003Vu
l+hYr/wmnOJj0Cai1unsGMHllOfBmgrUoNkT8kbyEe1PjEr73vZCQBcckERzWCpQ
7ob9ChDxM4xE3q3PrUY9SFODRDPe7IiRGFnvF7gODwnXxOulT5fRFr2zyBphMaQd
pc5o8aoeHwwHPF9gGS+Mcq+LXKuRW/Tj3Kf0I6Bt4CiG4Zv1H/7bBpauJfTa7Mgk
I0idcOgCEWSqD2LSiL4ApLx3JawEylv0r0TvAqlqrobKP/lsm1/octmpW65mFb96
jESdRynG9HTnYxJwpBtRhsntx5QPfiUST7fTXVl0EFQVJVcKFayxr9/UPnyKSI4u
74otfcumMOI+89SbzKPyV3mBBDcOiwViKtHJNwSmDO4mI0YkeKpsEBPFhCEOLdmU
Z/vevClQPk0lYjS/qRZYsrvhFoMBEkJueEVnMNm1DYj3LODyzjmxKqCFsEqOUrNx
c25IA15gCKAOLjhYw/MUfAM4YG04a8tYMZSNhrihCUCcAI9nkQP31xshBOYRKU/S
3zrm/7FaszyoFomkK0++SnAjWS/yutfr++gm9Lgj4wMopaGJSwLSgg7ZFvhmgleF
mQ9MKltjNmGvKknjYM/VQvuEOHggVUOWxObljLfts33T1ZKwydsCf85Zeh7ot/E5
JgXROAwRhPq74ZvmIQnX/HnuZ6XloawGn7kyfvoOeLBpinvdnS/1tFjR7K/QyryD
8oTTVL/SOmC0Jix7KJgROOpa1F2+gD23ZwRniYKTo+4+r23Z2C6/NgdCEwcJvBpQ
DQ6lN6Kn2xO78Z8j3R9FmdkgsGiJroBsIVdldFEma79vg09t/5AXT6+lwohCsUfj
JPzVEXgq9mOdJYr10P07ptOsLeKKgmG3AYwvfxNj92k2LHDfbyEIKxV48Ntrrgxs
nwg79+05M9QjrvaLBw0LMD8+hIEItyTuvy5pnGrqaX1kfNZWss2eUFHAqKMs18AS
cTJAwfcQQB7J1732aW2MGkQx4yWkkET3MdO8qyl8ufv6dz1b7kV9PPfkSMeSilp5
neAcDiMhazM+UCFHl/pm3URTxDEH79WK1IFZExW7kp8HWvT1diDTheAPCbtpc3g2
560m1RlnxFL49ov7pIPAP+pa6ddgIh5pxBtNPvn3DXOjjNDQl8ZJzxpcHKgWHCGl
B0aEAhWZxkUz+MHOP+CFU5gQNN65ZOBjKqMTTPDhzc4lH9xh9bD7YXoBvnRvAgbz
lizNnYoiqX7G+Di4FEKD4Kp3eFP6DVwBh7n2FniyUIvHpEPR9JXs2rucr8cS+81F
/WNcloE8RaP72jAAayXPM9Te8ea7bV2HNpje44J5fADRZ/48HsZJqtZc+VNfXkFM
TFw1KKcStqTW6/Ce5OSc5kbNnOTTX3Afd2XLT2S4FzZIMRfM9cEfOxoD2xM1UgCs
guGtM6AX4SE9GyDwBnGNkBaFTUisM5HJ6Az0mSq30s3FA4CB2J+KUwWSp18FAnTu
hNXH8dVyFhMIq4P/oPI8FagADXHAXrqzrTFwSjh3YHn0fjwhLOz1Zjq7Z2TedGHk
rsXkHehOr6LeizoHS4Rtgpz4fMoQTayzLEPOGFDJPY0mBrsq/fJJoOPqs++DCzKV
E2Orl+2GhR50CmF6Vd247D7BZRoGcyryQz7AexIcBsHkf12+WwyTEIfL7YxBPuMe
Bwh+MLM9+kNINJsCZtIPNTdYrlelpconXq1pITH1RVS4yEhjDCrBeM4XpsIYFwbQ
+aa0+rU9dEeNdb0DlJZiFXpbhaAxMNcmV3CE1RBHp/4cGGxE3QFNgCmJLMKKgHZu
UCtNIjZMgMIqEqHG0HUzAPvcP0gFOtIXa2HdFjlKmAGfaKN11jJ8jM4osGwIKnCr
XbKegK3p4OBIX5fhijXdf2Pg0SykszAATsSDJIFGQGHhVuootOCj74UOyPC7kYVF
O/js+ZsvRsj+qzjJ2AJEhWIZ3T48GG0/376AdB1b7zcXk3nv5WuUIwVZP8c2grb8
yimdPF4LApE+D2RKERE8vbXGHmQKEP/JlX8EoGXmnfQwirihf9Ejl0KcJK8J7wPt
QxnTNLXArXjiPX2zax64KpdRZbMdxr02Sb9SOGeXlHO5tiLN7Ip2vKHdSvoZioX/
+QxoEzpmegtoduPAZ6fWEfIFkecu0E4Yg38B7tizT+xwE3TcC5nRmpCf3L8iEMmb
jyRaVxi52NspvEbsF88PY0tqcMNd9bIrrwa+7Jxy2losMGH43VKOLoblproihoUr
L1iFdzst/MWirWSpLgr872HJSVOmDhhDOz79/k5TKnTWyS8U42HoU7HKjSDxQWXm
QKssBz3mPaCnLmPjiffyhla4FbkR7faYlBXefCTFdH4QllWaqKaewyJVw166LOuu
IkY/TVNEksAEJRZwfKHaXQVLublEc1WYooxzBXX7vERI8RqXJ+YpIqtQ0hfH4Mun
kHYWRtKaHGF1XiY+1bDaLd9HS11NY5/XlChTx5k8/yq7CzqHwNccY0PVb3xzDV9q
pw2E7eSGFU6WYzvRn5c4yE3cjdlAKM1Oj8jPDINZkDjdOHCSDECunoQbsrgw8a+o
Ui6STltWafl1NDLd4rQgAirSB6tZWuZUH6GCk9DhLu/23/7cmxmMhpuPwe3kPhtd
hKWUBJ5oXvGFIAln6S2qkyEmLoY24QCaBZaZCG/uC887SFS/pc1v7wRkfYgd1vMX
VM8hPFt5Xwy6NYJVqxSuA9uOgbDKWfE6C2YexQxxogXQE9GqPXA2jU/CmRTe0Cer
Z1IGos/4rjeihYkclu8xEzcoNLEicePfL8YqXNSIM87AXx3Mojmn5x5oCbEgvMdd
hJ6xB7XTy6jB8otpfUAX+jPiJXquYRwV+sf03QvGir78cYmvhIkDuCTyocutmdQS
EVZBn7YHRhIs6DwyY9EoPd8l0v6XF3/z8B+R6VTIbutkqDWQZq0peWkl97rg6/mc
HQHStuZv+qa5SktGCjPdWml444shPwLDuXOP46Uva2CrhiUZNGXSWN5uCFESurnP
fp/TvzZ1vL2DqPC3q+coXKe71bwObOanPCVUQQnBRbaIN5TXNxZdCLeCiJlSIjCa
deLyPwF19Cptr9/d06t2jRpkXT8OOFttygRrtnHB+ox9OgLMrkgqak+fM5DtaMS7
xFvgfiyf/xGLhn7LKajcvwnKDYP4q2aXRW1PsJP/17zM+ozm4bIcK6o9tgc1ToeP
fdzIF9Fz/NUYippTgYNVVOByexXl3Y7jpIaB0amfXLREG/xxp29SKArmqkjIXV73
Mj32VV10EflXnr84NLv3Tt3Lx+qw0Sz4lEJ6xF+Iy0Qzz2dMW/79jEUSmaoO7Ptr
x30kjua7svzfQoCYPLBZws+douZlER06YN4UzY7T/FezAv+KUzkT8StlEPGNA72Q
ZFFUjoWCtlHp/GjRzFHaiPU6zPp5Rqw3e6fOP1IpPYRsO6z5JT8qiOA/qqEwfy+i
h9rokoluie9gvQg2a8QnGeyOdeVPkrx+2dBuoQ2IIT0OZSY9Y6T5zk8GynnToaCY
YIIBGYzJLmI4q17TktvAhZUWjkX9c4ljMrgTXn3U8RbKpXwn8q8glMPBOtOCXotl
VjW12sLILb8qoEq3OdMnqKvqX1ZlwHefNfTTIGkfgZv+wcDug7SbnFJQOasqXusU
tS3sSs4RA7kzuHOZjGdL1ppm+2/iv0Jj8P1H4gHzlE+oMwwWYFG0bG6TYwZtIrQR
MBQ4vQ8x6w7c6Tp4ylBvBssRuzAbaAUKVKYzw/RoZY73nBIV/FqklktFcJPTgony
JmMBOX7SMZjwNxqckua5oLRmfNz9XJRvr2fw1EXSAoofFV1F8meCdfjGucGB9ZG0
tawaYQZ1KFhfRTdnFfO0XwEcpBGU7ydQM1i/HHoOMqaBWng+5peZ5ZTrRan4xGPo
mVKgpiYwnGllLHz74pP/zwoTWvIcwEtTlJcd/7hukYCd4DQcmV9NTjjm1c89B+nS
s9BDQ+Epgj+HCdzBqZf0mqfz4QVAVv5FgMBJnSwf1VsUe7rX4xgsHHTIjvRi96BJ
nTrjniX/V1Y3UnFrhOUrd9eyTTzVU9rbdwNblG4dnXhGsPdipI7dYRsV6jvHFN1a
oLqhiTzVYvsxxHMBrPj0c8bHu2PnvdM3AHnsh8gaV9fY1wZTGd0EdckrrWCX3nfa
wFPZWpwhm9S/2i0sQgg43vJDYmc7iWiIqOXyFaddUgnmuaZ4phZWlIswUCusE1MF
DkRZEMHWEUUjTMoSR9xVqtmawDao0Ddr8wGhSeSsUWCEJqDxmXNtyoCQToUv2ehd
Ao3mk9NJeiXiP6Lem0YEsZg7NMPtttM/k/sIMBsBWfKw9ouSXQAh5qVDzHzVSCr3
Yzz0RcVfIV43HXA5Jru2Mr9+BB3wsO/w/HbO/X1NBcW4b2CFYNCCMSnghQwQfPpS
xgcKmc1HBmloigIkb9wP0FjsqeeR0pUH+sWXG9Zn3eqeK8ZORzcxqp2cpmR8zJo6
rFIVpsJiqFYwy7roXDUvzVbOvC7APV448V+qk5FLU+4+ZT0qa4b/pNj54XiUirVL
6NMZskKcQLni65vA9qba72Gk2/m5MvqBStynz7xhx2fRuZ4V9RWZ/OpYL0LYNNYo
nwKRh4MNZ1BrQD6egfoAn96vM2IyEhmjQbcfxVb0WJLtR58RosED1qh2UECZ46r9
JtQW6P7EoCPoV1n7StSVsLP2RzWpNcPVezdKZZmxya5Jba6s0FyZtPDPaKI3fD6b
EBCBRYRsRJj1DHMFPgkYtzsU2s4nFvRU4BdxJZmM1boSlQX76cQRuaRu5UM5sp+e
w471EvPyDpKwXw8dNd+IZLMef4we85TC23+QtJzmMBSz3GkkAZiPRYJWw9YqynR5
0a38ZlpqU6DNjS7C2EsEKxtILPTLBSJuOc+KMng9akjBiXUKelkRD7UJgp34oKus
HjMlzvRhU6F+ebZb4TYw9uI9kR0CkwkbP7tNzgoWImlJ2J5huV53/8TzQTV83gvX
5BD5+37znc+NzPHJMV+NbnvRkQ6dBGaCKmAZngqNJhjUdB+TjQJDTg1Ro5QXWA+0
dV0s0iMzj0fqfEZ9xJxmonqB2myv8KjXQINwMlUurqgkgm5KHOIPDPzAbzB1cO6L
3/Fh5AMN4Va6IkK4HAMgH/maBf1XM7Kp6ol+K8sHTQi8Yj7gKdw/pI3R2bENPIfo
IgxCEqMtDJXgEAN1HfWgNEPsJe4SUCnZM/uHvNGkGDL73qpStGBwjfCKnfZI/i3s
3X0oGKHlc6D4Qd+gKWRkffG4J9IOLvyP+OIbzzCAYWps6B4LwtF9UufcTmXAWKhI
pHd3xF1O2PtfL+DvbWocYkhZP/tKD/wsU1PQpvOyH1nPO2q8D+MADFPUemQfijvy
8hcc1zZpWI2v902x91uR/meHbO0IzfTTBnmYPbiwwwmN+7j2KeQxGW95H2S1JSWz
f4zA9hmTwlya4KeVx9Y04Hm3VQnaZkrnc/6K0qlJShPyXpbYsLS6JmLaTZRWkeX3
zfwqcOqNVfaENT2Shn2nM8b0u8YBSnUrWyLbKzVmCFYgz33d4OfXT4KknfQR7wZE
qCwtgY7jePgS2KqVtEIejdlCXn1zZ/wo3nsSdVU5sQHgtBCRN5IjnbhIg84ksxHT
SzIYIY/ig2l4LzB7F9NaRAhDJtHeR5kodWRibUDIz8S0k3AOpMPodT7DNopaWh+U
H5OZXoxZsyKwG2dt+boWlaG0EuQRvuAV0mT3sszdNcaSaLMmBMMVQeV9bwePI3sn
iRIcotAjjhkZ/q1yyDEctVUrZJNHoqkM8tFx73IMhII4hOP/aLRaUDW5hj05JSUK
Siu3ao/kBLGTsiRn1Pj4/mTa3pcH0fyIyA9yylPQjt2Aw1KVMq2PJn98QNIq5PnZ
AduNLLba7slkAuZysfD6kht1+IXzziMDNMKplyIJL90kgYMBOwuT6PukjjYu2g9M
cNOB8Li1Y04eglksq+emr2PKSGEcrAz4JFO5th8KKH2Shp2yPdMxFokFFpYW1HAM
D9tCLl9QIR9SJzGXCJOUWE6P5v89Ugkjiyit1Cq6FeKWUmrO0Q/Y0o+MZciXGxWa
S8NQYAim/E83aX5veQ2C5X9UNsoD8zKYUHCtIuIpq8+vS0snpcuFUcimVo5BsnKx
49fl2eclnNB2dkEnxw6lK/gwx6ZVwUCTxSVcSkoEb/Gy6478QDg5IZohc45iaOYl
zMHqXBkcndgR9NE85ovQ+7becGwuKmHM4b//6ZLmDzQxZP7qymYcazRrR+nCD6u+
57OcMyFxy8GSvRI3joMpjGLCGFIDlPI/RyZ6s82axh6wvPXO903004zzeFrGYxdf
sqKlJVzR+Eyc9AHUdN2e3jYT6S7/UIuKl2hlqxBnGgMxRfVll2V+P9sF0zlkKDXe
KoV4neCPs7MeMdRCtfIU7Rdr2Gmol7v0PkF6Cl9X6yaNLXDs6XivfeTiwLjPFbSw
xVHu7xCj1+hWYosowl6+6/CaXbTRE9VfKUvKcFjl2wL9fGwXYd8dzxHCekLaSWKe
T2H/X2tWQvHW8gg/EsZFdGXXucRSdfvQoBpqueKcBUc/QMSi3HZWFeHQryaQ9VPK
PXlUmWAF83Ybm+Oo69c/fancWdoLZTQlqIgiv03Nl6C4IAtrjMTlWPIQo3U4WTBe
XVDdt7dZ9zIb5rO7pn1mBu/GsIAmXVHl6m/P+qdaf9ql4aWbNIs+ch9dmrOx1FAc
oevLuKSLk5FjaQ8gW0+V71+q701vv2FSNdPi41T5Fe4UNFkM7KkDXquWoGBUpjpj
2S8xoxmh87dWwQ6zOBiE1RapVy7v5aFjtClHnZKvLiB/4IJ4lcI2/Zt+GiZkyckh
D6QK6OOpN6mGA2zGqvGtZ7uALacsVQ/XHsmNAIzUbwbYJ0NfV3DQXJsVeNiywhYD
N9j7+51XDG3TDdvSedSWkX4T9Zr/KtJJ9nEVA7DH4zBixNrdFU9raBOpY89t/d0L
1wwFz5kab6V60aOgvGqynVozBG9PQYjKTPVJbXxQNKSE5xgVwa1SewMfgwRUdXIn
4f7NYuZDQiMKCOijZIBI7A9k/bpfIVnn1apXcEhUCmiA4cWchF6hXsaZ8jhWlmzh
6FGFSqulj2Vt21nGiC3qzIo+gkqdM57r8CJMvqA+IT0BY6B3HN606o+mdFi+BX7A
9nKz4R0CHYhtP232y5nHsnlsZU20uYvPWtW2si53gNmEw+dnHU8V4DVK7iMqfjuu
FKuq4abn6ghAWsi12Vk+72ZsUBVExGPQT7senmcM6Edk0jLykJrTBN5JkK6dJ18P
tYhWR/E/p86u8QA5fywyWg21/AhujJ7HwUydZ1IpoFZ+/F+A+Q2msLFwjsHIAIK7
Fg/NDGckML+OcJOYC8xNJ54n1UAY+3RvHTKqIz2UNAM87BJDiywTLodT1+RKz8Wx
5lHfsLlZjRcE4DmsLX5iqtYV3tp9vOGvdUug5TFup5ArXrkyEIt820zv4t62ZyVA
9ggV/vtf07m8es/ySoQar6o9eRhreMFckBvBYg2uGCIIHFnGuBuEJdkBBqeK7M7l
t6G/9aW4igakmaOIwRH6/xi9LsqWWyL86r+sDu3ygAGe6yhd3uWnlnJuYR/Gc+yE
NBU71Q+M7j2np52naMxUGRS/JUJy2QMd8qrtxAEbDH4Cem5xEBtMi7KgXo+/W7QJ
7Ak9+eWulp2Td2/9mpH6e06bSYCmR4uNqsawj8uBzZXC/v0uGkFyw4Id9FdINhMm
Q9ns7nM9HhhOJf+zM4ptCmunJQznoYvDDp4pk9bw0KvWWyZwP0uf/EU1MbFiiNTN
xD8sRUcyoLiKYAKSJ63vyu6USkzj2pdKL9VFZ54ygx046qfr+w6KbXo9/QTXbaPX
3VC/Nxp0KxXOzIa+VODxteJGfhyzb/2ib3XUUqF7McYzrF3V753XKmVDTgHu8NQm
9obXCIMSCtL364n5WN2PhXanYmfGhkqY7TarfX60oLmvbhH1cesfEr4MzRhmFcMQ
vsQoinoFTCs4tlGlUekbCk9aw2zo+anUGixWKzwQL9bbOBSYi90FA1pHIvIa/AfG
t99QAUSmtYJj2Cy7pVJ+QSgmix1In2lD5kDH7r0h+hGrkDX8OZw66TosziqUq+Bp
GHRoHXgDk+B0uBYGECanB+VbNORFSFC2CqBz7JomxMhAxdqzw9QSUEkDehjvwsZb
TaTnh+EJlOTizHP/QL5vmJwxZ4WncBbZ2IarVRXtBYngbq75Isfg0GqwtsXWCgxM
GsfmqNbsB4Yc+rSxmvshPReYBYEvkm6S/Bgzmi5t/iodYESoF2221s3pvaNqdAKN
v6rqPmicvXNCfhGOb7nJ0Z+LCmUpZyt7RA7LWzXdCcxsow7YAMwjmnz6xcfDpCJa
QS0dKy5peuWvQJz/MY65dTiCKoyk0nlQct53och2gGbO5uChxNVx6AWwNaqrKbJ/
bgt44uaxZkd9YD+n+0Fh9j7+rkjMdf52wVHPD12DFzkXmTHaoDpBiXLYTV2jG3DK
ZIg/tVB2wTuIwfh1rf1cy0ZMAjMmcmPXZCSxs8j9L/A7eyRWPRcr8928YQLjhL7M
LC08Z1sDyKSLWXtDhfalLGMXIR5kN657LycpZKi7+1061cD75HZ652Rh+DfgxFHb
+dSBQF/hDgd6z4HbKdbSWS2ZBlXV0nQoT0wKUqM52lkv+ccWDIuDmSKHDZ6q+6Md
l+nXJLE/8ccbDe5Eumjr2+Q2Yc8CZh+ocLXtSjqNZJFfMKUBuPmQtOTfReupt3Fn
Sxskye54XPW3I3F0UYroJLrkkbIA0a+n9FbUSzKf0nzPpVJNOS70mOieqW4fIWOA
aNCVynQlhLGYVpArxjbA+hFM6PLB1MbCZ2PVfwt6+sg5xHKEjd75QXwYeGK1BKUx
xJoKWCrVmwHSkT5xV/IbnzQkXK6KjXCLh/cVDGXM3SIO8qWR+WMLzjOQKtxWnkQ3
5Tp1+plILA6kSoalHlL177Yj3Xz6XwPo/426r4yq6Rvii62+cbE0zN+aa41C3aUe
e1AbKuAvK8pPZs+ep1JFXfQSqnq9G5sGgyy4Xd22slaU2JhuX+YC//fe35aarHVY
b8OCxNa43RooYOpMhmjnKYK+z5B0mj0iG6PulyQ58DvY6kZaATUc2E2TWweinvMC
ua2E7WJxVoOvkBOZH2W6T4y43WKZldW0JOxeg1xz8nMt3Gaizrn3XFBIIJXdwqXH
Yp7MRKKkNDSJ8W73Cam/QNfGO7+LYx61OXfMrAVGLb5QI2UoDjioFXxV27+Xp/8L
fzl7mjnMJWII/koeb0LPpmPp1blebWtk3e+mEw1VQbqx95QY+yKHPuC7k/rkndji
5pKh5I9G1J6X5cLH+wY4Qhuguyu66dkiCb+OxBOtF6quVa2EvvlsLfmOjfYb8vmy
WS2gytbK4I61gdwxhtkvL69SRWUnl4taz7z2PY8ozo34FtayJUykbSuGvdGZuQWH
zUmi9jnmH8gUXSKq9bYy5bfhWVK6detReOU0cUQBcDLC/rTqrRmeLZCVsB6pp1yh
OyX0LH4R+ggG5q9LKzsajm/ctIlfnZOA9+FcjJi0L6Py0Xop0tz/2zikzlV5CWV4
u8HUnKvPMxz9gja2OoqV4/MQDSYwo1mjEcM446gxeDy97oV48KVl2P18dq/2EN9z
MrkaG7wcPZszOlvh733ui6xoiPk5Af5zbcxW253VcwAaw6CTT8WHQmb6t1Kl/+gO
60LQFys+CN3GO/alAk+VmnhRheh/ipSku+YhYVEk5oLQMp7/9gtuI5Pg+xeipPVQ
2WJE06SoEl0I5cg2O47k0O9Vscu2A8c+yn6kZIm/6bxkDdJT+Jyrr62FIusYnyRE
yULRq78xpJIda+fbhqiYofD0ty07bdKognjZAn0LJy+FR+KcqIZWRzmwdrnJbIz/
a+ADqWm38QtpYAOgTdKa8BW/lAgEheNCwrs1xRNjE6yKDfTwBqus3yxiBp+sKs+8
Kvdc60K2wUTlAHNB6y49/f0EwCLt04LF1D94KepBQqpVCg30vMva6Vr8r4XypxnF
jy7AfB8nJKLMkXO95UqEFdEwJqOEThfQ5rU+KYdS2cQlbJi9n2LXvwYjsqBfL+ke
ucIey/11JV9jHbHKCzGgLYK1nNha3qg5wJ7gKl450i2S3PgvX+W4o3XXBfctg1A3
facWYILnc2xn4NAzxOYDoqPBuoWD6iwmUltfm0OO+oAkSfuTvm9MQ0BCuIm6eJU8
cgL46bGEM7hVL4rlogQP0mpe1M9qUfFiLaZh8iAVgj+IkyhVzuzQZYkF7plenj0c
KBymvbC37H24XCHghSS+SO5JRwzBVUX0rHdAJb0avd3/n5iotoxgXO0cPhvyaDZl
FGwHAsJlKEqw+GSsApLjduTuFsrh2BSZqlLkjUiCeeBaI2PlRTTQwUCP3anvMSk3
ND6EdQ0kI+3KoCe1Drmh5Ubqo5mho+k+y1yh9LCjagYQtrTaYlPbogKFm0tnoh11
W4qy8G+UF42UfqzJS0EeqgntTudm2fPIDuZg0yQBYemBsIAQRGKEjzKmXQ06d5G+
reahmX52lCWSGGebGkM9v+9c3XJPzWn7AAt80hP0gbq0uPKEStvam7u3DhBRZ3hk
JHGU6SNPBRQCKBVuiG1eSA1yyWo5YKWh5eDBl7dNcqnEhbdqS+GNx7TkrD2dgYs2
+bbnArfXf6iMjqk/6HrNl7WW9istIQ2juhi1qXgs+kio1vToO6GmOXh1JrqC7q+n
Jx+8Owd00dkaC4G6jPd2pAFJP2SnCa80P8oMrqfADGvgUxL7QdKCQ+OB4fbAjFUf
ijtCY42NKOjpnhpqp2V31lbhp7N/JzvPyMc4qz4882OI7l8aiEmTH3JksWeBRGwy
BvFTQXEK7WhdsVIH2HbqSRgAgaZid5a6okTuO6SK/pWUDPxpQpBb3pJJ+gfcbZF1
2jcShhH7mq1he+B4pdWEsOgXutDZimcluguP3xTKm3rljYqNKhfJ5mBXAkZPInMM
FS1kf23dwmEIMqXGlV6m37gEjifJINzrMkVIQPN0EGM5xlgXT2wLpFejg45aOKaW
koLkxWy0s8XgAH3vq/x2hfXwVqfgqhyRbZ0+gLQ2NDURppDR4wywrXRaIMWOP9iw
zJf2sGlPAZdTnJ0ep7MdTboh0KYQlZgNlWoX38n+NdnDhkzgpNZFwG7RsPvRzIJr
B/7IU9reWqWwF/Y4jiep+eEF508Q7CqULfoKaVzxikuKj+AiVuskUB0sLDmgzd7n
g7EYZOo/sqpDcrFEPm2SvYK6aPAL9YoNC5cp4Jxn8NKBQQk7QoYKq2q9yaeAhlMG
Q8a2x1EtolsZsRY8hVzit6RUhEDxns91QE7BlRmQvhAGKD0JNk0oxK4yZubzzp8z
KZOa/P5r0rtvSNVWPyuytlYcDMCo8dvHsxizRM1GTa0dScEvZ8NI1GkY8X/ltjH9
yERpCStirfchPSutIEQIHU3syCEqWxbJBC5aSAbf/q7gEdKkL9r87Qf/KuO3/55e
9tC8bx/pqwmm40VRQ4hhI4t6IqS+ryjFXRnpyZl0pKmgwUqKn4h7v+TM2X3Ilv2p
HCWLvnsbSpzs6P8YSywWJAOPqGjFlDJN/AVRBu5clIjtVhsNa8Roya8H7n/1drQx
ub7iKg7/6TJcixa2+YqmRXQivs/9d3Q3VoKwFWG+MsZDt85yKu3hFVuvYCNC2QR1
hYaGwYHU/xM3vwgWMqV7q8GhPHokSc5TP0qUn2vaEtMoY0XUwM5TR3cjJZWNPm6m
1mVsnb8V4Y5o1pAr+fnWrWW6Jc+BCNfW9XWTEtyEKEdXx7BxY6xD/dbJteiKOvDq
D871QJ5zYpIcnwEs/NLshbhlItb6MSvUkisFFScJEPO3zsIf8Ix0kWE99eQT6zlr
/0xi1CSvL++Weoff3dB5pT4TaQBEuwGzNr1jdGuBvKs8mDpZ/gvOvm43vkNArSH9
yg93nOcEGAZxhm/UW2QxFvYZmP08qUUJpstMaxnR0mJjVWxLDf7zKfk3iDKrMJFL
pmQZB76ySIvE+1KBjzwrAZ2naDxuoZAgk58+0WmXhrcneeZveDWuZW4vFXzy2bkj
OnKtZh6m5/5arlqyyc6Gk6dEOz+6BHsjXa84/gQyQTEqqFn3fp38QLA7+TRg2l4z
T5QuJCelU/fvfmdmArRWYQxe2EOzeWa6CUOgxrjUkdwx3ZD4cW2CqB0YLt4uIAdN
4fMPl29yBzDskajovVMifSkGhR2EPbZ6MlJ5j2u2C+t0cdBdfQp75AT+Rq35OJBz
vDMwExderwwd5ixxXqhyVOakdSnnMg1sFxt1/FYFLGk5cSFp5WiQSIech94TH6SS
EA+Ceo/NEYUmJ3gIGMyVtcIHYL7Ie3jG7P78rFbdidvekjZKEj4A9yvA109bAMTA
Lhl1y6/36CXh3uy/0WhA2H0YyUkCNyC0jHbMfRQX6lEinWH5DHT2PbsgAXRN5Tw1
xktY3Jaz5LWJWzDp1eCka+fS/ltw9ZoJK2c9NDfjW3U7Wgj6rUFnmt2Sukd878/K
PwVdwLJuhVJ1jaEjz0Z6xWIrxwKOkAaxZNTnxfJoKnm4aXVuQWGvOt4RmhK+vWdn
0bjFkDivLXnO3pkqv5uIynpw7j8XE+nGzuddMRuUFZUc5ebC4x/SB7T+9ZWJjk4l
WYIJurP7WUaxXGVDiRHg/dHQi4SMinazA0Xs102bBh+MGPxRLtufldHn6L/cEKit
1dOTvHkhbiiCbaeKGkyLuADfCk6vwInC16q+xAXpP6+PQhA/9mSdjGGpZwju5GKI
AUihVsBzvD98yf60/NTjWPB4sipIJTwvPvSB9EWhkmi2bfaA530NyPYEcE6h8lq+
PcBJqPIWhIqp9oRqjsXgHjV2v8gcdMO2MNg+PoJirwnhkDAnuIDpSIRybRa9yWSN
uAUeWGzdaVzZYVlxPzoJq9ME2oHqYjExmo5ESOB9ID0DJsYNnhayrO60zPF60/iR
bbidZ8uU2stt7T0gpC5spFDki6r/syh/HvebetA0iTkgDGfcn2tQO9psTRjYEH+K
9MSFDp10NIGZZYgodO24yVzPhLNjzSj4UcrGSiBfWgovuvqZHg9Yste3TpWEWIBt
4aiZxwcjDNTY9++AzqM9lFTlq5JYplgtMTh6Q0HVymOoaPPXsi0qKPrRcoaryPuR
YY+6LfLzNHNJRanV7e8M/OMng2+UKROg+wBfaLUYeo9zGZnfVP02/WtEo0bKbEep
WrF4bNpmUhWjg3fJBd1YvqDiQUdJTrrdxRFZH5O3yt/TfaZGfnVgA77F2Oa4CJHB
Y1SeBf7+qeAgsv3xUrSw20Dk21hX32IR/I/RO3c1jx1kalZ2uH2JMMiAJ9g4AmSV
SsOObWg7rSMRwYRI/7xLtRisyvkbBXn00Pj++LBgsQchA4bqClDOPNJhoBUiXZbC
IEy2i8I4/S05wKpVPthWp9HKvBO6CPo9i5lqsHisanGHNxnHt2Ydk49EUWMbOb3S
tXKHKK/IUi2RHIb2H6prA9owSigmmqcKq5oU9z4MNP6E4GZ4ROcUXZhdAvk/3Qvs
Nk049A/n1ljZYPGR8t6VJXZa63+VE5YQSW+uL7EgeWDh0lkUgYvHs/RMFg7jTvK7
qopAUTULFyC9bin9g2J1TjaHCwnAKAgFIviRrqu0de1wjNYk6EZDFwXz6Wf/M5cf
Zm6QCIrEPAZCs+SaKjYqKefCIg7nd0fJ8VXuBy+csCfvDylNiBDQSeR9qojT+o3s
cCoqFwitUxfy+9IhZN9Qho2zeKFaUFvndw+UJlqddQqI0J2FFgBzUOmPsRqod8LC
HB1rFrrVDGPfmXpvYFuwlEkaIa1N9rkwddGtw7cA95eBbRo3h74iyIK2kU8XHQzG
avClp9xDPZeZtG2BmVrTjdkAunZ+IBrsd0LhOK1P+epWKm48JCQcYo6GZGZgpptJ
KM4ycBTalcKh1Y4DJ2+ptbVZ0t9ia7URfAkxNViYO1SwDMpnbUOywyY+rhe6P902
fIeVut3Lyla2qYDoK/2D/ZuCJ8K5+MAxo0+Dyzv9drXdrMYxLQC81SpSx7LfqW4F
rk6bt2QR9zUecxPigQhFJoUE4maANptoACg3RYzKKnOZIw8pmhcCU9dDEmXkRNNN
ux8zh+3sHo8d/mX7WHR03O4s9GvIyw2zSydGhDhq7mZXw8LXRjuKWWlqt1ns4QOV
/px4QcV7JKt9iny01AWCqxcIHN0hgJaQMtJQekgxw1gCB1shEviaFP4hKHqPZWa6
Fk4fp4gkCjOt9J5kYoj5zsv/ait/Dal0XlfCZ/cdlx/WEff3o5XtIM2XQk9/LKh6
rVaBVn6oK92QLbqJWvDNN8OPRZDTVe+myxi7V9OibKIrNovwvAWhpRI22CUOb1wR
9NpRadES18y3/a/Rgi4bkCk3GX7gkk7raKWYdB3nOVrt2BHCTdFnDM/AvDUaciKu
TfN0p4oMe9yoUd9SkE4bnOczci/QRdh1jlyAIKEl5F6OqemquQio2CafetdwW9Aj
J7FTq7Qhqh9FZEY65Bovm820HKO/KYcxI3A7+A4b7s+ApyzIEJ0QOVwFnqghUHio
Aiu6Yq6QJN+RN8iaTTwR10I/t7cFUZlxv1hXFhjl2Mls3XHQbds+Ou/8/F50WQ5E
eo7BvSDLcr/bIqaQ71JtiIT1iOFE8oJ+AHx23TqfbAnXgARzqGvez4RMtXUbKsKa
yB19yL7vNcmyQN6z3/0S9u8ikjVl6KavvJgs5xVvdx04rLxLLYu0ABbPmaCBBblR
/fomX96vwHzF0PUM1aF470OdSqJz9aFG612nABnuASukkhWavX+ZkbU0Vd03/8h/
kdTv7gufuF4TFiAPGj7CpJOqmzeoCLJMu5sKWPCmfWvYeRhfYEij/whBtDp0JD4O
9FTo11aGGWvveIeGY92on9evYBi7fLLg3sr1UfbUMmMk0lWSwX4fs24VoNb71SFm
DtbHpDgo8Zipmqsipb+4JPUSYjQpWu9iT/ekF6gCWXEY1Uzmi+y8Iw8a1kZJdbX+
AWdf7E0K1GlOOpF3CIaJSl3eQ2tAvCxpAC3xCA3puoUR+CeqvTh3VSn/EF2wPe45
P6suwWmvtGex/Vz6NZiGHGL7sk/0K11rY7N5sKolxSE+Y837spMaSrzryqnb3P8I
QCpnZ7MGcuIsjdofdsUQXKh5pCF/2Gtw1oWq29ITN2hwyuvtfpLayODS9wpGurmm
Ir521uBxb/17zDzQMAFmZFAgv8i8vf9WfE+iBTOgeQ/BGkUXoKTT4UdJ+n8WtGeW
mItalmQO/xNqyYXsOV13Gv0xD22N1t9DzGpZkHY83XZLQPPxHmPneRObpAG9e7b9
9GPctBECA4dg40ad71oorKSHIP4oyyrGcPXtw6dasvc98TSg9vV1LkkomSMomNbV
pgvcF5j8ZDaELdyD/SUcybv3t19RJMlAbVphtFgjGI/wwqjQKrJQP7B8c4TmN33g
f6H6VamyeYk8uB6MOHRZ4wk7wrAY0vB/M2TThFTtz7zIJKPIk+9vZuRR7jZy3NxF
+WfdqbH1DENOuSVmi4Ja+3TsM2F2BeiIgasG9+VMzmcUaS4+17Hq9pRn/G6UIsCp
WRts1XhvgSyWh2tuY8S3H4wWjTZCFu+gsV0GrTBdGdlktCn/OVNG3Hd5mNnGiZrT
9zRxlMU1MDD18gdJA+knj3gr2NcLjNGMZQiBU/ntMOkKD5XqpDB4d9UfDpfPmw8+
zNBHD9Bel35zSVxBqOKpO3Vrn1aqcbT3xgJTJOD6PX5OdnGaVZWbdF/mGpbEZL57
dAw1KyYsjCwdS0s0jtop20zPibLd/aqcSNu6HBSSskxC0JSpLnOLxc3f5kaEGCo6
lXR38i1CzYJyCW2yan79iKH4kdHw4eixGzvVZCmKhpJ0z9HVryWljbhlBWn9jRh6
l40t09ZI938Oo0T4f50ZY3EB4O/9es2Lw15i2vynFydAD/wymwjQxLRWrpuQovEW
4m/8iRuehWJHQ1LEXp+3tAAQp2e7ZlH34HGRlKzb1P4oIova++3sg6tB9Sodl/5+
AI2n6NvshZi+wbtLeaN0LBbOgEh0SUPtmETgLvbinfGBPvrFHOcP74qJFU5WBFhb
thicdVlQS04ZSkAyHYOdYw2Ta1B1vXuvMtsVN/93ObatgGadk8QfjFiwzfjLJGPN
wxchwBOzwHE08h6fzoaxzVNAS001byGaMS0QmV/CPAAP9We+O+Qs2VtG++xr4Brw
nLntNbAPl4NeHq7AyGG1pcy6uvyVXZEKRXKCb+mEZu01O54yQH2Fuanf6+F6ciqK
s4IyoTDp8MUxU9bpvDl/3YHAZ/jNgXfFnyr7ElH4fYhMWKZClBeB6xUdKfohj0vi
CkAGemSPPEA0lrXHdpM9n1DiBF5NJfYndTMUffFM0r6rCP7hXi9ZJ1ED30mAw90w
UJb8oeaV0FtnknJBeWryajV3PebbyzR+pHcwPskQFhn4evW2LuPK77QOQQY0w+ng
jMFW4vC7ZjK0TNyD4QHKFrf3GbtPzKYf0o3JX+wnGeqC/yShZ939bsgNit+//cMU
A0EIW5D5Jlp1z4fAr9GHVFMauozB6KTv9M3NeaiksEdwdjYEfUSotkbEUlKRfwCC
FJ1wwHUr30ur4TQNmZr6OB7O5xyzCc88lCu3ma7UxrHDyJc400+XF5T0Gt8cVPR7
t+tvCK2t8FHAVTubgR/aTPBJozvAccGxu7EzTQb4U3qe8aOxV7VkhGZDYIPZFvGB
8EvIW70dXgQzNpIu+2kq0H/pOCGvG51T4ibQOyohuXMIXXHq3rN5lYzJae2vuXK0
Gt4BDgOxrlFot28DAoyXFyLji4eVeX3FvS07azOpAJOj3k97j6EiqY4fB6m+5LTB
ZYMdIAQUTXpLpS/WfYYJNcMn1jXM/9jT6X64BmRiJJxOlXlVEq8COXje+P0E7b+l
GDV4pVAghHyBKqJPxwuEseY1jQZHuwcNmPq+npYzRhqKg+472lQ516SkSy3aUvtY
NUlBLake/vKH7lvV8Mpsbk7cHOa/uYDYplwrU+Q7Zq/s4X1DKJ9OwxCbeRn4WMXI
NvrtK2zGAR1L+lHrZQ+evrF09Ec9jodZM2OYm65xkmE725PMKiuf5qBdmutc/Jh9
6TBjm2OMQ8sn9x/314jFyre6YYFzJKviLm5swo/0bAYNzgUsgDHixbw5Prkm12CW
ZFhpM+Y1+wxvuc5mL/khpIRG0RG++kOpFJdDJh3AS4026zZlx5THzdtCMrcFHNOh
s2DCNgl+JiLnnVDSvwdv408tWBh6y5UWagT5/ZQQPYME+UFVfqv+BjaBA2qymLx3
t001ind0fxkOw0YOagWL8aN37diD3n4mQPloUrzDzZrzJJ+sJ8NiiIYhqdRQ3V05
/FSHHqnW39V/5lIDPd3S76FJwrJHYfsPxU9HNQs652Vd9hAXpMy54nDZtvh3fXUm
MUxeUJ4hQ+Kt0o9XXgKk0fVODyWR94Ez4Wz1ve++zKesCvJLIYkhHHEaQbzTtiFU
Jy2mo9+G8z2GPUTErV4HH8LljkWPyOBnFHw7qfvUlRH6qtkqDUD3pC9XjDLCbTVV
G0HG6Ogrxth3oFQtEphtJH9Qk2a6sH9mP368rFCr3KIjMhHKfjdzlhN3QjWs9qkQ
PsgBVUTPcXOLPvmLjjg2EZAeIgVE7JNglyoHFdUhiydxfqdvpZnaf30iHfkvdU0Z
TRus4tsWqtEAoezfYHrEvUKiX3RDADEERmZOgmGj/ga8vYbOpHpcN9UIAw6C+NdC
YVFYdEpWrQuGzLse71X4eHfHVmJF2mWPnOlxJ9abMw1yoICURwcni7bLhVAciB0W
0K1zSjrErCvFwUxFmHvdl8Q4jKO2QBQ8dOMDQaZjUoZ1sweIINd95Zo97tPx1juu
KcONIweHX1ilkKnQut1tgNUJ942lIK0RTKRjqkpme7ULNm6rmo9Wb2CcNBw1uyHO
4MOAEPTsc3UiTXhXArBZHTH5ksi/RrmEUXoJnVvfzBc+ojN/RmELe9buBSzUhdgt
+J6UBI6pU2eSwLh4EkNWAx10U76YJcMa7AYUTp9MEgSRNxCvpKeSJA1NBTUWzA+m
LwdpkouRjS5eD2KPX2WBSRX7BpyNz4NB3gf91uyNK6pycoXOLsA7kDQYspdDXyll
9H9o7Jir6T7S7KO9mtQNBiUp3xwbD7K2oCrwckrtbNSOe9+934NFrKNVBcBaRb0v
oEAcw/qW0VXdqOMqnSNQNocNmTOrphcQKJ4LDut+APgIPZO3FNrTwqtKqc11N7bp
1wsMqoxFnyOR+0WCh9nzpB3jZxOUUmsxJKC5GsEvmxdJTltEh9D/ufipE+LMBQ+z
DBMMOD8t4vdPPIxlWmrI7EXaFVny1Hg1HH1T1fIAc1idJuN5dtF6eOLte41K5A+S
JTzsZ+rHNlyQ0ThLoQWkAqsCGjdepXvZXqTZqx5arLXwz4JojCtNYBemM3BoKdcT
eLoVlStuSBHKZLQO/gwgGwSuptMgxeYNwBFoJQDW1ZUugBoF7ODVyD/1XO7NlHxg
yl0ZteA/L8tN4IH7yA7J00um70iTe+z8MN/82P5wGWdJsjpXBReAHJtHflFRd8Yf
Fn5DpxM3vWg/MS/grg46/tOTlxfJG1P+aZLZq1PBP0bMhXr+FzL3d5dPVx94EgE6
cQ33Yb3xs9dh67AHzuzoicV99REoPX0jLz366/OrztOKJzXAqsmSU1gcI0a9ka6l
q37xlsvUabzLtKziSHbmYmAF3oaeslQ5YscGScN8zMInGyB7bSI+q9s1FfsHX9ut
375hWL9ity8F9IHWtXAPRwcvMI8b7ELksTZxz7dcV8SvVmGrmrPmZHhP1N26jm0x
+8dwQauIDNy1vpoacUVOVWLy0D7Y/ts+N1Av8rfRs1YGT44a34TDqXfh8v3PHKX/
aL06hdJ9HWbJNL7PK4xmkVghu+bdhK1l5Jwo9bxyI1JOm3ZhbFcHNc5WxI33ui21
hrL4RiMsIGNXKTX8UD2A5luY0MAqbnf8+FNfE2rZJf+Y3abu9lC1ZldQK7VbdrDv
+A3Czl9ONJwRnMwrx6oPg9j5koq6qYzIBdy1FkUj1bRxJrDSXSNL+wGdifAhlK9l
7+h594cGmIPBqqZ0Im74cvnhbYvMKjCMtLmSJ3R0ItUxZ36wNL58a/NHWN61wzk/
pVJ2EnLx17dlLTdF+y4ZZz07umUoEhtb+O/CDoKMEyW7jF3d2SIDIveZ69/tHGrY
So2E7wI1+yhioWfllP7ciDbGRHeaCoHWdc5ToZ4ASJVf2G/7nEdDSy/Pgszcq6ZD
KI4bfOkez6m+yn8tRQyrS4LyKB/clmFqHyhEJplIY3zbHeXjnNJjU0EFXbbos7yF
90MQHL07NcVKZWp2ddAZC5Drawz5yZdPHf12ZZOl72HItou0cIqgaMXigq9PbeSV
bpCP7TcKaQkTWPOPdHsAFUG4Qu5WGFslqPb6jIp8CyRkIxtG5pCDgHY7k3WFNoJL
sKwDh5ERC/28fWzC2CRVPsk09VDVLOZrY1TesCSlhS7kegKcfNhmK2IO2Gvh9QCo
uCEzXAvl2PgqSWp43V/X4ELSGichh4mhgswZsU0P/uiw3odf8WnxY2ztZrNnVwR2
2o+h3GzvxXS0hxrn7XuklmCQa4m11FilwHO6c+DPTeN6KbMlh4ZZKvyZkfbl3aEC
yFv3/9xWvAKGa9Hgq8mVxs453kU/KIJEYoyhvWhT9/FlnG+ibyUTL+tsUujcouzM
FTT6UXb1d1AJ/Blrpw5g17md7CEKLBuDTRfwu3RrYetPCj2ggeqLxemCj+3xR1Me
VdeU93j53WsNd9DcESPXB/0o4EcOJamrNWFkhrcWK0LyPNPOya6tCz1eztrLmJR/
WnWoU46tiyh6IpP2Bw+fNBNX7gZHsFPp518VRzDK2QGmvmrbTV+Ge1rL6aFugJSQ
AWhBRNOQsJVlPYQQ3TDpxas1PDYvpMLJ7YCP+y+kNjxz+gvwxDMacpZBFYn8F75c
VVNYa95M8uQauq3sH/eBUlXV/AvJEIekkhVxT1iSmgOpKuLeBnl33xV5vyQqIUf7
3wQZkH4JeNSPGbqo/9cNg+muX4CH/QFxcFzWzImoPv70UzTWhQfq1I7DGKdQXF1t
VUmwBs6llDcwAxDsrnKYCIo/8vlObYDxXMa3e4LZGiTyIxJi7zfMKGSa0eL3dmYB
oAzDbNTA+9xrHOviojNjSLtiIMkKwxE9XRZg4X/GhISRClAhaIEoUt4FQVFIVhs4
SZd9L5meE0IkRCSZrMB5O/F8epViF70SxBEwdGa/ggcx++m29ACpNMNNPaXOZtrf
3y24qJooTRs14VzhjXqp98uOm15E8w28qBlOpRL+QBr4+iwJixL7mcXxn/wr7jUx
wPkEIEuLKQ76kZC36GsdCjkfAc01AEtWlnjxze8YzttVVVdrAnxWnpJcrFUFBRmA
hDfkDes6bxcEKRxSEIJQYTjCLsVvK0BKRPOcRUqWwRoB/TzDxYa+Tc53QFI5D9TX
DJIa3IqzOKmRDSUk3e9Dr0U1TFspUpYg03iep6/QdHOc38FiUYi56HBDvnT/EjmR
7LR8XXM/g3LXqHbEo5E179Uzs+ekQo9C0RPvSOJqh1f54zzNb5LLFJakPNLk3kHj
0hKav32Yu2aX6IDNS+5krh3tcF1r+OKdrkVCArOz5k6b4m+RpgfYve9v37SUeBO2
9emn4Pr9sM3XOuH1dF5VcqG0Jf5ZACfFMi/a6zHq5iO/UHoYouya3eMn/w8Mf9AZ
uj6nQF80RY/BvP5BkJd8nK/mmMgSa/lvzt7Qj3/WLAhxdK2yc8oya4GdbUfkxSkk
ywfffFE4xtwPmaSds5XEPuoS2GXyNLOALBHz2WAonWmLE3BvdNl3EtBsqoq/yXKa
kkHpNAltTHHHsMsmhCQoBvvGMUsc45EUxbTf03dh+EH3VBJfEI52vdcpYhhpfxpo
erWcbhkrptCwl6Ik+mbnjXc/wsC2+lrdZbW7dcVNLepw+4g2Mx0Jdabl0Lq08qhg
AxznZ21iirtpTSl5FmdvbJW7VO/iPV2DRan8NwxNEFbOdLGK4VGi5TDPssHWhU80
t3lHEYSmK/ZitcZpnWQXqFd1HLB6d/f6bnE6DVj5ePixTh3odXH1Z6XNS6SHUct7
tKIhOciVlLVqAmE7wUPTQ5MO+0U01ENobPWKBRbQlg+HwMyWBwQuiiult/U0J/Ek
krSyO1HPdmX+8aaA7xkEaGfc4TtLBoyCwW81UqWt8b49YXT0bDfVSujTVs4wmk9k
M17JHAnIcl5FgNkOjZ3b6WPWwHWMWq9uyNcNPFPnM3SvFP23Na2O9hPBKXxtf4S4
oixf8H9vom5Xof2QKfXzsaSCiCZc0a6+pYOtpQnWgItVy3GKlvkIddRSWwggj29a
Z1vWJB4Rho1i6sZm1A0DZRvZwJOlhKlv4Hx41gXQUZXD9ycI+rccgc07WgePOu8Y
HWJOL6NM/wk8EYmZUH0xU3j3WmBnvyAE7CMiAdvsgCa6iEGQmGcNcCtQYScGKJIL
RoZNRbWKBkCwhuotzup8m+RmptCk26DvuEmbb23OonRDvK4qqniW8qj5+buzVCOe
itARQs2pfpU1jS6iBjp76eq8z8T+sdKtdgTCsF+BF5lADNaOw6/+25YDFIUf7CQq
fM8OjBJdxKw30f5iXN2ubcwR5x6QWmW0MdePZuquuB3tteYIUab1zzhfgZzb7lwf
+OaOg8yYhksb7S+yCJD3RFkpKdDz8v+aUkC/grCmsIcEqd/zLe6sPpaDX5/CpTdT
zpDd4vnoscLcm3mac0Y/sds+kKXJ09drsfkAZDPvswisK6KbZ5HZ4UYJqB+bDf4b
DbNkaPlu1OECz9HaoaAe68kNoqnAIgD7D0bojm/2ug/booP1B6rTOxxGDW2UiM3F
ANqxl+rUDCoYSrszlazg8ynDCVl8LFfTwmWVwscpKpIJaGsXUzFESBXoenTyukRO
RVdEA9J7ZbsFHo06a+Csn27UsR62SQQg3USXHdrMFn3hXEGrkTfDATHRsr+5/DOq
2QojDK616qixzNARhL9WjIMlhh2KaQXS77vGNe5cvlN57TUZj0O7eMjj0pjxncKN
S9F/jOzgrTWvVx+jMZ4f25a5vp9vRKk6YitYVCm5f9MHUjBton0BSXcmrIGRfm/D
RygbGfmtE6S7l5TLPPiIDX5Yr3SEKYmX9a6CFgMKo6O9weezzVx8zigCayHtdoB0
c335U+kxgg5kuJypxsbjZR698z5q5rXPsivgm/ywm7uwaGfN7e+yBb8kebq7wts6
zh+CQtRjB26QLYUk9l3xQB6bPJA9DU/zbg2prZZNLFX2LENFIjuKbu+OLKTmY/wf
d8u8F7mDUdnHOFFV7R7qF5apPUuKBfkprz7I9N+RC0eoQfpcOT9qmRxT+4cSwnir
pJPeqhFGuEh84shSX+cCab+p8ARnnf7lo1kNHWKyZDdxUZ9PsKkc7jDHzO3AbL44
4GfiT9mZzqyOFuwYdtdIFoAERGTNbDadnc8I3vdwNgrP8KWPApd7wNpCR4HQM9iC
Wf9HezqSgOtoZB+XgdvsHoZF9xQ7WJ4R81pV1Agzh6QC3AR59LC5KMSdICwCJbbs
zyJnZWDjwi4wyb9+W7+HEJH26eLV4UtemZdDmxwj1Ta76oAIVG0lePJzqXZ0Nnfk
C0aVbIm+1Q3gW3dmcPLEMbvWRQ0LqejRBge4STKHkBJVgHvdNFlLgJMTMgbDScTh
Im04abD7IyOvjzfhZFvOqUNyPKhNtFu7yas5b13IkJ36/9ZJ5shs24+Det0BuyVU
NDjUNb627Kf4/N+ZATW2XhSrMlwhTs3fLEOWT3dBQuxqz4TJAnjIK3u9/krlICiq
QrcqyCYVOzK308QoxqM6F6cNWJulCAGxtn/jR5R+UiY/tez9amyr+UBcWNCade0C
6Yqz+fyHlszJOlROl4H/MQJMsTcfbchNAxrQPF/yFZUTC9gU0d96+bupiE5mE7aW
MVGoIAtXL2m3G8ZJlYAAM/bBVnQn4T4RCMLv2JxJiUdj8fwkrSeTN9EAClSbPFNb
oNpmbeLCjO9DcxCDmdYJYWSJNyaoIuqCrEV5Z9au82vGEZH2hNUeLs7mPMup1x8W
WDAgjX5WjobrK+eyDZ2lpBCbdxhpbMc4eRU9NIxZNWdgiuFOz+GZ8tqTykWXgb5T
7xZR5K2SzkIBafezf/2lhOrOyfUbiyeigMH9xHsjZkwOw6Bg0b8i3rXzhDGv4xU2
vp75bGG/cgp1txeqZn7mg+m512CfKcA/ID5CDWtqnVtB7jks5Kx+uWyhnD2UYLON
D2TcMwberOYrl2w//G7WKbXV3V/3S/y4omcdVfwTNK01KbPSFYH+JrQHWzKzD8RM
qakalLdhjXDRob3DtmuH4cSGK1W+w1O0DVTw1lgLaDi1LNaHOIPCMDhWw+OT0tsR
7pB3Xe51q6HvzverJrMm31lmd4Si5Cr47NLRSH6Fd4GdARoN1J/5ts+I60DXRwSd
xsdnN0jGRKA7kQ/yu7aL5ygYx7W2c/e7n7aIaKiitkAaGv4In5D8zGNnuLHGi4RR
H/yinUrv8LWzD/lFpz7QDvO0WoHNqpqDonaVADDFqs8MagD/3KeVijwgDaIqjcqv
0/hLRGgPTH3t1tUIm7S/mJpNtqx8L7fRjqEyCLszV+AcTZ4K8KgRaSx42jzij/wb
G+WdUFyjuVec6vmhP2jj5LgRhjXHHa4Z4yoiAcRHfu1+vY4oFTlpmK1S98pMZp0D
WxDGXgCaNlkB570k+vblef8oVmsZM1miY/nRgcRS6EvbC3qeUDmd54JgGvBeIuKa
aGQhq6d72FicMOAqJPND6CQ4AB7+sAijhhZTK6OBhgMj+LBwQ298icn+pZxjUGyQ
GBhvCZSn+g0uLeTy4eG9+rTnQKNLnOdClFxT5tfByWaW2ZsI90y2yAiO3uyopASO
7IvwfZtK/B+ksA0pkFYNkoblSD3TEfTfNhgz6O91vKaJPWEQcTXOGJo7lz6jZQOs
Yn9GHyTLhgjkQothIHcX0Yi9oHPLA3M1IplpUr8MT3ExgPF0ZbN49XYJ70inO5rg
8YOfflZb1sSi2uueiPAmH2XQGTtfxHnF2Myl6kSo6IJt+kqexO3lvgxHQHY2xTiW
Bl8H8kWVtuKWkW5arGSThgQBIPjFKnEiQf7wpTR1Whl/qr+ctBkOJvkBkAYWyDfv
5ZvGMrnW3lYEIeJgYs+oIEGgoOM2iPLK2C7K3k2cN8J7fRgsNg7JyCHnz7pMINTG
G9HzHvu/HKXGYIdVGlo11K/R6QVch55XHWat6NTXNRmwGALk3d7VE1ob1PayluXu
o9Cf03GLzmxCKS7PP8gRLn55+DVCHbPSPsVLqF0hpczxwJHlhYBRkcvUyK0Msyd7
3x0myaeoSfz6G6OfARTqyjVBzulDIK36d5OrSHXd86EyIpeqm9Y+IqbRqD8GniC+
Yhpr+68wc3XbWHYJGRHzQ0lqcAHFRUrxfBg0b4yUY7le8BjB3OVnsW1b1yB+3ax3
h/KbYw40XQbcyHJHhMFtpX6UWubOw1BLZgO3PxKtevVUlBQ0eisvI7i/SuGvBOq9
acV0UCBWkScKQxY2sA+SSuPlWt5a+0Kg1Zup9A2XbRokwFF9BGkbjohMyJ1TODZr
BseNJ1rhL4euSoGGxTzNKIK12+TpdzCoT3u2c9FC+Q4SxJmtTVqd4NK0UMk9usQY
d4WBp8KKE0vDy3gNL9XDvwfUpPa0dn9kckGpNl+jd7GMz0ywcDwY+FSS5kuGwvKQ
qFmoqVWTAouJJRsuJ8fcVTosO4ZiM5dCEpk6RQNze258MuaFGS2SAUh22EfVWLXL
oHxmF3zv/2sDa349yhplFEE7Ik7g7Pvtt2B750JWkTaHv95BD4NoJD36GBeAvtoZ
J2sLAAdyyBFQMSuV12pm79WSso9dlC/qU9/J5om433VHqNOVBKlS607hBoJ9BwM/
t1sFzIMNhTkm441+bHkWgvITHjOeYcQ5s3mYZsWKbtRHvcX9tIyYIOv9tieG9ztt
BNOfBE4QuDbH3XhpucQg8c77l8J8EME/IMpz2E7VbpTu9nJUjjqLviyqnQn+oXmN
p5EYTXrhS6TJWvV9H+VcG1RMFY2C19/eQk2W3h17IzzHmgb+JveEwv/RXoAWoYkb
SYeIVf3g67Gf6JPsR+tTQPqhzv0g69cRP0gXn+t9OBxYWe82R2vlbg5/AAVYMxe1
K9VAAC9mWNNjpo0nJ7KCOxspGj2KlCteIafhrft/yRTzFY3LDn342i19UJxZ4Ykl
YP5W6qc+yr8iJyi1tT/AvbKNmBDBWytnG/AHze7IW1WAc22Od4RlgDLoZRmP7IdO
BtVXJlvYKLIgD90Sircmnm/e3AzbqjXFXAAs9WlWsYD6FlAjWn4zUKouF9R8ufh4
/8MYwindAa4JpT+YtrvORitJf+yJOf9nArhipRw4BF6XVGA+mjCKY+Juc9DHoGPx
N7OgdTmqwUyaXOLM59Y7qsXDZoePVGbopCFZpL7wNIRqPL265k4dOy6uI72K8euC
t1k3FJyEPy3FCxDRE0nmE6g4WPjfzqFnKpaSwFz/Qn8/5/4tcELt/UZnxl0Jfsih
SWPC4fO2tIvlVjvDotpJMVBY74NQHMcBj7bPAopUuRpjoXaDccaWe+wxo2xZLUlK
nnDWSrV0lBE3yaKy0eQPzeZdtl4PUsKa/IOeAmayliiku/CzMaeujOrW9uGGZgoE
L9g61sVzmuAGMuHzFB5+POvKS3/W2WacEdhrK+xrSJvk6na8+JCNlBBtxbJj6Y1U
CG+xZ++e1iifvAAhfECMiROogtEHpHhbkaJ945XEg9RZFw1EAVBxuGuO0xrfVzZE
IufgYx+IgW+7ZZMQTz7phRsBvuNjI+J2FVYe16okiLf0a6Zwq4C9cy2bDGr0Upmh
TWog2jVE7a/y8JFUIIVs6HioRvuwZIMtTGnbvzF9NxHWdS0AJ1RG+9XXtY4lbdqJ
R+mJTc7HjPNOZ6E56JmDREYftwHpzl2nI7tZ8NzWqT5RH6UpBiQfInB+a4i3rqPo
Vxeht+N3iH4GU8MGwvxecszOuDqP8TgzwMahwJDzg5fqnTdUuX1PKRNMPqBoRuuy
vdwFjNvS8mpG9R+0RhZ5BJkjlgPh+jgaI1vsbIDWCyDcFH6ceLhau8kVt7WSP00S
VztOjg9pWi29iwrWcDMSCyqyH+uqzlBjRuHS+o+Jhagl6kqqJbObC7iaihNe7+9F
hG6VAC9067ZpzbaKdGS98mhUroVxXJbPhU7KOv3Fhc803FhItbqPfxuCnw+Mv+ey
j35EbdaPCn4fUb8ud2B1ehLFdH8WfDQ1/hrf8q+8iWoJ9KnHe/aXeakDb+/KJM4h
e8PZU4FQk6+ItlTf230ZfNWuUXMqFPXYSkG+IbGgtbYTHe23YQuyQb3Lk61C40yR
NrF/sUwjnsspoVqLzt2egWw4GvusFiRZB/dn0Kr6dwqIHCNPXhkIHsKCHidYevk+
BhAK56D7DIrxzEZdILwCltrTrNATZnj2XXU2t/h/6FCjc88j1eT2xEa+0o489ZzF
2j+ZSFArxNDft36Q0PxmFuAjP/2qiUXolbIvi5wEZobfWiIBIbYME6kdyXMcmAF0
JQvSYs5sOFXCvrVdK1lKI9+TbJka8o1alSvvJjEqLnsfNsrmFS0lVgJ1glaDoTVw
IDW4QyDyrpaj2Icc/wyEKJ3mG9G9ALbO3cDgOkZDznS7bMrX4gRgKAZYa4sQZnHZ
t3MUWSOWS6NTfbNqeS0aRPTkD9QkcjSkWmR0dOTXzJPw5kXzKZeMSLEKv2/3tgy9
/HlaS9Mpzva3F6xzg2d/5uFr4cbfYuuEweLkc5qwIU+w9EMU4c5b4ElIcgPRWF8X
7q2ssMdQYkaiYm3GJ8j0CT2T6nloONnGrWizmmHa5XghA1oX5R9UYFdjHSqqW96v
Ij6+tVTbXKj67jS7V/LafAZIrevHPTMgvhewLFCLCokNHjMEz1oHPMpAgLUh1475
Je96FH3a4Z2rp0/GiBAo+Smm9dVKaj/n/hnPYj18MaQeqYK17lFscMxKLbGBTOjh
mOX7oi8qa3neKq5kFJN5h9CTkt0QCr1PzWvyFa1BeQhkNYrHSsy1vSsup3kdI7TF
Y8JlLqCNmj0PBYVcSS7NJuUlHVx0iSxEL2FLnysB/4a73NZ6LG9anOPOQ5wZvDI/
IAd0DV9W4+nC18SUU2NBdU0l563KAda10ChRsWFpxitj8UKIa3z0XJGXwiSwchLy
ubL1iAcqOWI9UH5kwZwNRJ4zm8lGOQ1H2VAWTAOZ7l+8D6ERajLJwEJpQsH7FXec
5yPNpq03pOa1WhYaHDntVfAIglTvk3t9jW6M7J8fTepc3wNgZP4+dnAajm/cz+IX
FIfhmjsOne3ZNWpbx/8X5oCSwzcJEJ1hDNBJMT2zEWZrAx96vaKEy8wxnNleSQEx
kTQ2t7QfYoSj9E27dCNmkqc9FA3hrSENhYEuHPnY9IAMsV9MEDX67kDEMKojUy+B
7SZp27G1LXV7y0XOtwSiojsog2Nm0Ld3bVbkW58uDEDvIeJxOWC8sF4m0193b6UA
lUQXKV/Q6tRww9Ej/RLLEagWg18sY3i4QqnJ12cdRacVAJb6UbaXeYLq4nEpONlZ
oMp9CqZbJTxo+yasWHWZ5X2UdJcUmUzzjQ78q/JCSAHHSQmBKd/f4Gi3EWd22757
KjJ0dpfzu1+dbda7R0kx+2LzC/Ed7dX/ruqk0671VXRrCxLiLr0PfVQz+8b1KTjK
4gFsdKgAp5wJxeLcasV9FHqqqALC9ZU2gBO04zA912eUN2nPXxjDXBG3Hd9+4yf8
FvLMrKnJgnqXAVTFIAS2BM44cUyK4GDbKcrS4xlCe6PK710RDyXp/fG1OmRNmeQr
bXFLUy5jatAeQSDkKXE4F+IehhEznaW1Dp67ZDRLDjgpmJ0PmgN7eq+JCESY+pUw
f3Id60FHHJBVEtHDZ3YHFkWc1tF331gEIC/IN5RH2uqfz3nTbKh8uoU4a+HnInnr
Tau0d236J4Sf8sWreEaG8oAiNFUY1SHY5Pac5tfr4kO+7Jh1Cz1nSCZMDudrRdin
DFaD8Z57YqoYu8+ZxlxdxMesGnKK3CRMesi+HumctiYPCcpGzU8LntJ0aJzAeSed
BN3zjOUdjTMr7eQ6kOogBcf6VB9NTdn26bO7VzTQWLAxkVTNR0qGfoSY2qVxwwYt
C7/sxvHMXMmfUDrOWJx6oo+hZgZYJCQKkaQ9Pr0ZFt5wB+iCo8QEvnZ01qwrU7O1
q0z/YywptVEvHbkUxlDQkmk0r+pXhz6VeoMpWftURkfEymdU2wNKQqiB7EL5kfIR
p6Qp0KSg+ApFvPy2mbUuIUGdcSifsel+fR65hVRDr7o3U+DConW5mpRK4xFVOxai
/r7yb3DheZ+v2TPJiGMBcu4QYgKgulN5tFNceNHm6XT5gU/DuyctPMym4XVzSVWf
s3KSDfCff0w4IYD4HW5yB3tIO28hc9YpVz0sBpfGra+3lx5IBuZER1OadRB6LsED
yvaNau6poCMRyLrp3J9Vai6dm4ifiaBceN6jtqVZqpdX9voaqr2qeWEiYNXPhb7U
K+DsYuSOBFH1YPXhkTZ21qDFU/nPFXSQo++ixCBHTJlu+YmT2EzokH0NTAjf0uHX
7rSnxg9Yx6rK0U//vQGm19gQ0QsdabZ8x/DAM7+VT48LDf14Anzb0lklwIyl0+9c
EzMhrt46IPTLStYiylytCqqhuP2bRlBiIHiDkDATwvPTy9Rr25YZJEn1DSQTAV4d
KTMolQgPwj2+Lr0ESw7kxLTfBmwFW4/is2OtQj21q8mKfljC+CpUX53vg9Vssn4K
sx/xHypJfE65aIgBMWGhRgw4O+5xUIw08D3QWEbq9XeAERWiWCYyjwm5hcnYRa9t
A0SC7P0Gg4LnUPMkmkXKQLPIIC8LSKOE9XORWEWqhH/+HKsHW5Xb2FbWBhAHosVG
ujmsEvj+EzYIEnQZBmz6d9t6HjYWF/vll69o3Aw0LxO9wXmv7IMffh7g4ZiadwXq
SHULAYbBXEANGHvbgE0n2Zl+c8/aS6bZ9MKmMdqadVsw1Bx6ub2e2CxU1eB1pI8Z
+o2ky80bo5ztWO3xbOOQLn9yVBo0d2JvdTdoap+uStUcHMXEUpU7LjnHuMx4RUbf
jkneEGWqjuSf6y1HT0xLx2QVZ91s1jIednH9vlcXE8Wu9SuGej0m1CT5GPS6KFz+
MmBbJGjCbRDkC/LEPITtxSnXItrwZi+GbKGoVJgIc1sDcx9cZUGufaj1E9qr+2v5
1hEPSDiy7N/BjHdyJe/nUx1KjylMxZOdiggRv8BeHkA6scnLR9hMl/kaQyxjnUiP
A2SR5aFHCyLrwPb+XEA6RT2JGTmyMkq87tcACqDuXNzDv62feekwd3hADAutCXAI
twWC719oyBThSr1o5v9qlWQzenU8KXBLHp4nH+tQ85LyR7UwsOLDD7nk950L4RKg
5YquqPd4+JZ3T8Rlvr/rToO/G3tFN1tB0xlfQQ5PlnzGl78GpgKAkeZ/BfvkFIjh
9cYjyouTQHu07GSewMRq23mkkezKYVv6YO/3l9pNBG/2rSwtTc81CLkqSZCxWEfL
yBKiPUF615BID+3i3YWxla8cuovoQWSRoP2SfmRt+4yF9WgybLvpoQ1sXpsD3Qk+
o71qa9i4tOyxkKhy5rINtUGMqwI3CflzYv2mHenbnp2H4QmvwlLan08BOjQA0Qdz
Md+C20h79DehRd3Iv9Mfo0SpWlbZxqh1AhvJmoIRP8NQkuntyp/x/ZE7PaRGmGtD
biMj2pP52DaFGfoy6WADM/yQcdQ/AA0Y0vHIP4VSmUCOuPskaQ1U/OPzvFPH7RsL
FfBG1JYoXtNMUqi/c6Mry4esmg9en6f/oZutnom6XgqaAF89sPCpzaSqd/SqGS3s
0/UsVfLynPt7lxF/M74F7YdsM5+RxV/w3nD6zkAaXYDHnyjiD7P9pTay36n1RUPb
bzzhYllWj3ugwJNRa3V5RaN7hJXUSg8FVxrbFfT6cPH1rh+bqUh8zvVKA8qSmIrK
qXxrtkA/iSn5txK2Jc6+sgFVuW0s9cyQmj30e7TWTPNRkMwAQik+rsZ1zNc62ejP
4X3LzL5tQYVelPUDoPoZxCNrwZHpeDDjkCyjE4825XA2e++YhgBaBdbt7iGdSLKR
juazKZP9lmDcqPafhWpwKEib+EdGubnLXyJ/ev5XYPe2DAAtrFbyKNgNSLJdUvRG
qUQs01vt4r1HhcRgOVGaP+rGBcn3tbSI+jxIQ/+yNQlBhUk9O51dPdo6QWeEiUQG
ZLM697bCkkDnsgfD6YxQBr7FA67T8Bofgq1iUERT1VRNT0go5xJMhgwjCDRLVhot
NGzz2isFUm7AVPl9nIibY/Pxy2l1M0WYMV7MrhDCftQC0fAdHTJednyUpBSsQnyV
hdnwvoUvpJGXJi3OJ3f3WsQLlvA6ddIteGZyMQ+mO1mWa0BrSFnbPZl2vs2p8pjs
zn4Iy3oJGowDOZwQPbjyBWFV0o6tUd/1WSV7ogFd949FJ851fqf784Djcajr5u4g
SJ0FYBpGe4qHioTMixk/5Ip0+1rbhSD9DpkayXROdEwpnBvUg0KN2ezZBGBGFYvu
HLkzJMt2ot7B+YtxJ2TP3ECyWhnduQ478A0z57MA9rLOzYg3dkm8CZbfwXzUKmal
OSYTfKSAlqVYDfq3O1cGoOVWKqGNg5N9QeDAfq6oldp6TW/0WrCWH7VbBRsVw74V
ndw/jZGqzCsvuszHgfjJqQz0sLHo2PEaUZs3YVZmwf97H/O2R1Q0ROoH53aJOD86
txF+U1jravpj7KehmQoy6XQGd0o6W6qANQpti1WzrZbgF1z77bGkCE5voKAXP/92
DssgvlTL3jFb0e+5kzBAWNJuPtCM5s2pG/TIIuQ+PCrG7uO2ChuscOz/FWgglNEf
tNHHXGXloN5j0XA7+COlzxYJG8eLb6I+BHeogMO/T6vDF9X48308zoBqx+Ki7jzE
8Q5y0ewlbKo3hbX1dEaTTBUzsIuIhlh3dIilaHq3SzaEjMRsiw0EgWJdr9cm6JYW
UJk4dq2Yyw4A1QUIOADJFXik7QQYySxEbYem7zPOSK6k972UhLvKvIfE7f4rlUtL
yrFgiLYMdwWJIOAKHTJLmzb7Jd+2JFX8sdIrsxTGUUPDMi6MsM5CPALoa6Q8tHjY
BYdtsBdq6WjCr4RzHJMqNiL6BGqaFOL8g3hzZS8GYxsuKNVWczHag24YsI5dhTxT
9UOIiISaRkZRnlShkT8AT6q9FZpUlCRbEDDx+WWYAhscMtozyh7S70XXCpRkOPFM
Zj0EnuTVUkPL0puI2tMVMwFimq7mbbF7o6lWYruFjw5gqng84ibun2gyMRBHbX6R
//B3FGBOyb21s0pBQYLgG2dvMrQBqjWunPYvfZRoAmP6EjkLyctiOuYZ0sikJPcu
DWNrKqcYbAPh2WbAd8GQFQepCgFf8E3AvB07tHQx97n/oOUmQS2HfdY3uiPPw4SF
v7ec54X7A3nyM36p5rYJ6doHewWxGEf6PfLP/TgkbSMhREHCWiwh5T+sfCKoukzv
RlHz0F5VKdbHLNE2lZAkoON6HLwZHxD8fxi0t3s1JqW7wFpuYsNYFiAAQiq1Mg5s
riVwoPx1LyoVRrp2qPT0nrvI5ocQHzWeUxggamnriQAR/kDVMEHTFi+PYQwk1q5j
2uwVvCeFv7MLR1HU/i0kp7Fp1/q43Lz95YXb8alAKloSwAtDVeWsIU5W+5pDU38f
Ks6QY/x1v6FNhx3Cu4qID2ZTtzT1KSSfke/WZe1J0wPgoSlgrbf1ni/L9t29QqnX
Uj2qMWbEBVfjzTXvr0aKdqfEbYHYBY6w/gPG24zMQkiMjdu85XkM+zPCCmURtppv
ra7qzrRQ2isvLZmA3STo965MaFYWhKStJjgy7duif0I4Di5JtmPEhQaJDQKht9Ew
zJ7ZTkZdDqQqseKWkuZT01EUG15+Sm915HudwVaMnGZXF6VQ1n61YHA7eS+qygjl
0XxYK1QqC7IAgVe4xanXGtN3OtwiITRDD+p+3k7ecGoBMnImDU0tOKF6r+j0vjG7
yvhOZeffRjfdjBaUoUn6z3N+uHa0yNyb6/DiuDW/lrr+eU4e/mO+1ECNnQoz8jrj
sr1bkMJa3Z1d1+OsT88/m7Rfy+6NXYxb2DWm5+7tYAQ2Rn3FyIapyk9+ySLd1gVT
63vY6c2gjdb9l6vaKE422ICli+zeZCfEnUeofYqkyoawoptNnssP+rJFY9TRhjVw
ZE4+ki9bD6lkr9Gk+Rj8CB+VVLdt8V/tGpsOIrwcb3/aIQi8qga/HrT2eZ1IXGQO
J2dukT7NLsX5F4ez/P681W+awZPYNU0+sxcSBtCjvb1SjWcCiUYJwQa/RQkvo/9d
Lmh/vmRL3hcxah8LaEyeGfMEy2PM7IzZsM9tfHABPGZpl8m4HGjP1JtK1UKixuoD
YWPMwakD1KdkgRCbJOuvvbWgJiDWTEkhv+M0QQqW6AycNACiXw2OTx5MBBqa5fRh
u/fIkGA2NMQSs7BTWQyhEYZxKPNlaTXF7cx71g50PETd98KKdd+jUJ2rAogbWglq
utu2pA0+VT6fLxyiEOaAXoMk0Kj3ftAZqoh4n985H15M9lAPyU0BmvP1i9P0iYh+
JN5Wk8ByQQVC0WPZGPR70xsQb6u0fWaLzMenoC7uMJD1QYuHm6JMd/IKI8q1MKaX
78YmutocUiRpy27480qbnnZ1qBocVditylX3Z+6SdjPSB1N5QOl66c6vb65Ymvq0
apDzud5OdwLhVMp/n3nJorDQrd/yJzfJw5X126yovIn5V8c3yWeVcGrwnT38YQr9
8RpO6DigVP4O1R3ZZAbpFY+FRicEICjI6K+g+Ar9+aIBtZb7ApiLhDS5g7FxM1Wf
QDloyPTkcaZoMWciEFDi6y6qun6crf3RV/JXHCBwjHTHbQEOPdYOaTkyoMzWoZj/
AqUQxwjUTX6WW74oFHoNGjqfz7yq8cfWZYKEhHi8IfBb4Th6mxEXo0OCGZK3UgK2
RB1A7dJrcqYs9zdoi/bbTYWl6d0k4V4GJkN7oGwruTRKunHq2j8OG9WeEjVSD6ZI
OZAbuIHc4wQuYMkAmNk5occ9dVHSPF6j2J+WfruBNbzYcBZwMKQcmyvHeEle9j0q
2Y/dgo29REimo39GgrM6eagwwjbin/1jvzdnEhBS1DG/dyaGD/f81sn8e4K0xu3S
1FSSjHKIzv0NQyBgx+jhWDXSVVZtXioF3QUjO2mAXH8m4qYlTe0jt0znitJB7R34
uXUPZRRcgMEKY5Z4wsEzMU73FocfhQzksucSHBhASZBwXSDQbpGN1xEnYg3CYkbf
5yBX37dU92H2SiiTOt25eOIb2Kzg3otyC3Y37aNQF9aa1mbLTYsL5CPI93NIaDv4
hXWQaHQaL+NAKG6du7ocSTUd/iodUiVPBs0YhWWRHihF7+6gd5f/TQyN0kaP+wmh
bvdOg2HB3I/kaHSsxDH5qBspkrJEoEYeXfHn21eNIypKvgO3VMlnzWQMfLcINwUy
1VO+YndhVOcv2BTbBwbJ0BW1pUV+GyeOsA+Hmb5XSNC5iUf8467gJldv0zYa1WCM
IBXwbnQMSWoAdkQ6EAbgQyK/WWG0Kwewew5CtrEb/EsUk+ndfKvJi0DEyG0BbjwK
J6YGoPc6Tthg+pn8jPcYAWdy2U1hA0WuvwaZyOf1qEilDEiyFHkojrWeFfo1x8Wl
2Mm25OiusBnv2Thtbdrxm7XLDiF/E4uQ4H/+jJUlT/zl3zWlxYi7gd95p99RRMrb
JpwFcRNXqWF3MjwPX4N1Wii0ko6lTpwStDPf69mZA5aT145Eyh34YrHQlzSVtSoN
Gumn2MeEIgIoDuQwNd3SnhxtcXQff4wKa17sEN9P/LC0fnrwj9Lsc7LNiYYEi6HZ
regkpb4U2NVY0wHzvBLGzY/Qw29joRdcKwQ3DOjuMDhJ1FB9oZhytvYLBrULgi0d
nT1CX1ihrF0Tsnicn1WO/xlcIOBrl5xUvdFVBVVi9rxQ6q38/mkQ4G8nNtFTS/eP
xyPTNOdwu7ENnRnlL7kZ8crhM2Hw8R4IfO6fhJPCLcSZYRKtFYjh77+d+ZMrkixC
2LcBtJWYslNdpOP6EuFZLwyXokwdKJ1T7h+4BW/Y5Tj7SIn0Fwa6NjCZpvWVBmeb
qywbFobGfou/zSQspc6dvGsSXwnMYn6tL9Eh9tXFD3dURD/PQwpeosILEKEFmPi4
swzfEpoFbMDfpxcR+SgqOBYcw7EyQfVvuM+r0cSDoY5QhK8970Ps0U4MwmpZxyH+
hg3w2lbZFf0TY+hlTZfaCFV8yFaTyrlpRj9k4TtFbyt96/fSv3ycl2c8amm4JKcu
afDo5HnYeKL+Ukf3bZ3owci1wxI4RO2qfzRhgecq7sVuG+PV3AjsRGxW1KMUBA4r
hzqef73IWe1HlZD2CCDWjCOkExhz9ol+jL1E8qOFyit5fgEgmWv1f/n0A7c/lCe8
h5Q3EK61KvZi2Nzpssno6iS/6SGKmwhCColQnToWjU1FWHIjQMnIVpj7aOIT/B4Z
2LKKAS2n9Y24nCDoCpefFCDTTWFFPqzwdC+CJWiw6lK5mMwvcZmfwRDuzWEDETPs
9dR0DLkXWf1YEpV+hoFmkP7hEWnlED8N59nF8k17ZmBbmrgC7EQ94xFywW2SMlrV
fCLdJtFNddvdxEA+14V7NpWifuBv7Vlr6mLyY3WenyYZff6/SBCSiZCgFcXC86p5
dz/3aXf5/PDww47ngVP16fU4OFRQjKOag7r8WzT9Y0fd8S1D91IBveCRmufBrNw0
LJnQXOntFUaUGanxhbGQKOAgi/QBz2xacrLjuQ9bbTq7lIfI8k2EdgLb0uWuP4FO
UgrDsOKrR3FB5IL+PmPoZGVEXCExHLqrAqpF66eQW1Om2aUKRW6drdOViH2Zyral
eK79gECLvFnN7SxeJ5G6oSlPXQVXDtdMTIDd2SY/Pee14ZrZG53XGeGJmazUppbR
JUf5SszO9EcVLu3orNelHfB5um/75Aszq2BETcAxAveeZesiYCLwsHUI4DTmfZ86
Y9A6BPoKWLutlIlC4NT1p4PfQ0OkRKhEex+KltvdwbMZEJLeRIAmhky4ZWg6rCWh
mVR0Cc9t6kLtOH2+Ug97CyEywBjI6V6t22GoB1CAtD+2ecvM7SkArOMnT3rmvzV+
S4NwzrVqzAC3uhRFDpieJQQvU+CLhI0ew5eVIQf96goJjmCjjknLDKXPmVJnVMDX
TwAWEUHEZn2YDU1tPjK7RXu9+OvYVLREDrXug0DIxW57pDy+layd4uTwQvwDqWrr
46dfGOSxWrsyME4htzoI1MhaBNAGSsQQZ67XTzYTkBbQLxK7qiP3FBdTRfunR9n+
KlTda3Rr4vWK2NsEgfyVUiB1iUO0zdGg9TRQjMxICYU4RUwFTOVYXBe3rCCv5QXz
tOJ6jdoc1KIlJ3k0XskO3V5PQHAwU6HYqJdPrKMPF2XAPaCyXjXGrr9QoScYy4hh
66+evKGCUoUsWAeBvBoMXXJPnFieeZkLpCBb1/hdwo5KPJ9rlc3RMQx+yp8ibV8y
1HQROGd+8H/EucwxvKvdvU9lD+BNcE7k0Fr/+TbFmZhF2yO7cMpRXwKH7ZnQqVaV
nOeK44ITPk7aQ87fnlgt+23r4kmOJD0StE8uMUNFBc2dQHtNTT3JciVGg1KInifF
vZ0A3Lc5SJo9m8gBd4g6tZMi8ihtMI9/1c2gOfHFzXx/CmdR8+8DRGSM7BwLBmoW
w89rcOOLZAyMufh1sbOBZyBDkMrhGl5Ysrc+ZRepofwbf7ktBriSmr+nYyqjuboS
JDFvfzT7CZ9xzz6w1fTIYdO/z5uoZiOGhtRJAL0L8URVGEsaB+wg1QATbLXOAKcv
318KAxwUDAqndh5NmlMwG+4aZwMNNXw2zWYmEV/OpCZOhDpZfs2fn05kFv4LYfs0
j0jjeeuGxH0jzUIHl4MB+Dik7WSvLiVvTUbmq0dP5ZNSqP2hOlyy6j0WPD3f/5mr
oX77QT31/isznH3c5Go6aUTYg+VBNeDEMGDISXqtjhtli5/BsHXYArEKwLZtZC3K
snvHJ8okQeZdCou1bGL7pJdrKRPSJDNS/0jzM4RBRcG5M0ZD1GVZ+Ag9Ye4iJHh7
XyU2irItRTQRkVhd/PWXNJJgAiMJ4l2Q9LWvVA7ezu9JgM1Xd4fSqoNE4DMiGmPL
tdnMwyDx7J/oJX/zN5mSSgHnhoSVjQYqh9ifXo+KWvB213CubW8thhbhPRPAH5Kn
9UmB1l1ups5zbRQbFcUuv3O8L3a3mcHQw8Ywy5BwgkFILQ2b5jGNw/flgPuQaAGl
7gj//7/5/LiT5+laR6jnGgvRfHRV4zrQi7LMROL+xuQoawS0pJ+TobJH73ZSdtW5
R1W3To29qpO4zEIi1Z9+dbzRN7GAEIpiIkXMXUokOa1VFAM0D8W/XnVa45i/HbJZ
qbZSGqTn9BlM88QjG7WjXSKIiavcLwy+jfCzMLL2kkDcTdc+WD/ni+ZXenTTxzjP
FFS6nPuwOt3kj/mswOMcpo0c9K4OH8ZW+b1iY049EtBVonr+xcq4+QpIShjfkdta
gdKuLgqWam6YYffB/lv1jeTuJjLaqUGd4FShcRsVUNx9BR/l5ernkhr+ewbIgfyK
MqBrE32ux5ADS41arjRd1Yj5KTdPTjAUOoKVrE86ubPheD/pkSmCESx0d15rcaUB
EE0AQ6/96i/2xIth7yVS6FGnlb+7ViFWGEyJzGs9pxPXtkuur+N1rqRDhTLoUl/f
EnUV7ewoABEYTfwnF3G0UFHai3IheAGjL9n9SA1P41/5UC1GnrzZlFKtsreGao4M
QxCW6qQEJo5uPISVkl2FjBUbtbMKAcHIDb9d+WMoIaCSQw1DX3GjenTI63V/LYF5
T6r4sQ3KFwmxLCLI+Tt8xmuLuJUgc07kMZVxpWLTc//NqQjtavYlbor9luzQDi/t
CdRTI32dHv5uuilH3kkICyaxJmgdqDz5KqU1OK/bQw+94cMofS/WORHNjdihhsBO
73RsrXMmKFmRFvwkTj/FeW1y5bXitK+lwq1Nouci2sswiG2rzR9W1zz3X/CAU27i
ykAzlqRmljGaQ//iW7eyErwk1kXIbpsOEc7q9Pe8K2scTcTMbRyOxz0okWCg1KBM
mTVnlb5CoMWzesY7xSS5qE6oSVdAiYn0WAemZWenWonAPUFyGTH9ktcG0J/ShPo4
aW1znk32bK8vW6fhwDBTI9V36qt6pdSBVWKsSXKtHnDGqO2Fpzj+MCtIIwbLJYYX
FMJ96k15/qWiWF57OkKGRJt13G5muANITVOTYWux54KWIC5L178bsF+mOwQcHV5V
27JwtaAj44h+r3U3ZuZsPxWmZ+OqPqxgNkHLMPXzSzKpYZs9X/3GhoQrpUzH/ynp
WQI4+Ypq/vNMhaMTd2biYxXuJwTG4rQukI37GIn7Ywx7pgD5rbpoA4Ofkx7NSgf5
JzuSprzi3Tqyb2Q3fk1jDQXceQQ1N4O+upbYOHHN/8fCswGuKxy/awmdObPu9T3f
9NbSdyi7LkME5g8djMgIRpYEAfElR3LmX+noVbnZ0Swg4Vd/vAC4zwJ7qHco0UPL
D2nNjoDuYvy6WyxLQcw0PY1F/FfQjp9fwQzFSaBrDWf0UAzYmdMdD5uCm7mQW203
ImU+DTU8+LI6CVUwagjDMEB9oNJpENNUdW7Nx0znPZ6KadTh81292cOneMXeMSXM
1pAbPh4uHO/Fj8/M9hwBuzT4HJiemLnLShCHHqXXlATsxbH2w7jlEtrHk/M3o8nU
BrS9WdkeiigceTFIbACWi+K5BkKVo+pGp5EsUNIh0gyPATsApXVXP87+PG93LXhb
NFFQFytuquxP5GeSbqFMe7cdJHX6A9bqs9NpPhzsQASLEDGHol41W02KdK0zLAlv
VTVRG9f7hMwV0RSLku3GInTd2a452FtDPFZwzB5W8W2LD9QgnvrG7g7wVa8w7oKV
lUQ1mrFpKfhBBM6gJq1MehXarF7Z/g6HJaHDD0T5Hua+D6h7h7hpCMkV3Kb2A+fI
T3VxZYHw95tRRlj6V2fBJAkq0PmyTI5ZCxLoZj7BGYqJGXIxwngUTG4LP148HTHF
ruNgCFSxgBKqRmoFGBwtmChjdM2umv1BLcg33XabCieaLEQnU1z0o5t5hIBJZdJp
vWQlLdpKdK3QOA9yoMaohDaf9REwlTbeu5Xs1SGwvLCMVCqKI3amKZhuSwnObJgI
NdL2zcGfOw3kc6q5GlY6skiC1HA+LweBjRV7wO8yaeB+pTAIZqrUD/eSdza/BGRK
AqUsKMDAEfodZQ6PI0gnTXE40RwkYszunnVmKQr/JI/hU+uqpA80I5e7NPRjldkr
G8sFG1C/6+ePEPuntCu6+nwYSXE2FZCmPe1LE7nbTL9lY52QCAr/9GvZxSyL1pJT
4c2L5GOpX44i0BIYgHEdqZoxl9XvGy+s6YFD5OcBmNmdJQ4e8QDopPmkuovezRgM
J6HpLaIbrauXEDtCuakL6kBK44jI3IQVSr5GWhxEKb4fJKNXOVw1O8T2xmOrgd/q
eCLskETUbVDo827fflVYurkk3qK58fxzoSkVUF0LY17xIT3NRazUrVE/9F7T9jT3
h4tRprbtDNKiLY5DCZDM0k1hI9uK63vXiQtCDzUar3ppYbWpzIPtGPzuXxTU2Y7y
HSuBXGzhmCJ0dR1BkQaJgPyeY2xfLo4nM4XQeNdY6Ki6MvH7hKSBbwTEtk7yYGTl
Jak5KHobWiBHq/EbN3RIt62kr6JMKPM2LVRj5cTiGHRfh/NoLryQcseUrmqh15Md
qRbag0jorWW6dII5/dJPzo6tJJMJskeQH2XYsh77QDD0eNOWl2x21i5Wf3pW5shy
4m1gQ39nCyY2LH3ishGVtyUtSjXxdpav1iuJZ8k9MctD4gxxxeTWpNBN2RuEMA3m
Qtd31rhYlFPahCDAioZSCLt4fV3ktGM7IyqMxIof8V4RJ2RxuXjZIlrz19s7I+4+
h4I95aXPi8txWLgw089xBxa58i4bjwXGdgy+eMtiogu9l/fwRLEyHo7H+qL3/daV
gtfBq6glZQ4DenD/y2hTGZsImsqjDhKB+Q94wWLZFN0w7WjV1okeVzP40RkfAPYl
AIooyjVVjst1nM33n5ZDeXNFAgEVKZ13EZ9DdGlTTGJaqBZJTI29WnejsxD7G4zF
HulLAhXI4LRtxjVHztDypgE3gf5JeOw5liCMWU7mq2UR/twkSyB3QgIcmMSy2aRf
zjIJDL7eDJ1izHx0HRF4qS4hZ9VAhKx7L2kI2dSqBBXbEvtM/U4YAgyfHjGHe7bP
gmoehSUhMFMDZPOtii+lSYkXGUdbQij13MaMmlrUnio1cQMv4z2ZY/qa+CPzss4z
rKWwMek9nDeokkY7YimCVCcNMI0G8wz4GHVmGi9Ck6BVmhpO4CdaylR+SHq+yANo
vatBUQzAKuos27ZBIPO2eXc1+rApJmPNAnlFOCnWweyy+UK6FFqIzXp7HWoL9vKr
FmfNcFkVfSeR05v1t48dPunJFPIW+vwb13KsOGphUR9pyDNaN1fqzib4hvpSvjgQ
ypV6HIzP6vfSYLUOz73bLSOP5slpczdsZJsjMQBxMKAwp5bKhFXeupI8aBuKQuKD
jkP4bt1nBysR11RFJ2wADktFyfBq7QMxKQBoRbg0L9tG9xdCpdQEvWDw8tujK4Hj
xZcSpcPY1R1XzROYOnzKZ40dfldgaU67pty9z9TdMaWJhb8Z0rBM30NjTuxZBixe
uF0K+1HFgN6ojd9Q7/8w0dCWJ8o4LsgSbEp/p4cxKI7RAj2jJnK4eJ0qmk43fhD/
fRkdriidfc4IEUtl9ObcmHWI3zDrTxwO0AQ66JOPsF2oV+mv4pYaVTI9DaX+d7+D
TYg7W76u5E/xZmVrObix36PZXkaMy96vM8IqetjdC1wzOuRSL44PeeIkX2KSAOgY
Tp/s8afQkglQ3/eIi2Xh/0KGvkjvnngedsZcqnJkxg270nRdR/C127qrEtZmyjK1
7mlhbfnynwPGn8ffizh/tf+SHXcXUHOBSXGvp6y9U/mBqqdwvjHwPiuCTgNrFJ+q
RjkJJguHZrPbmwaZC/DsJ0IXJ4dZecb3WGTumP6TGeHewXrKDNgbcGVKsmAaxT2T
ADmA191k3tTdJBw2IMmqYxd5gHrZj5fPbSh8Pjh3u7xjCEn7nCelolGIpxmDoi9X
OqAdYDEV+cZmtPsO0HPP8amJc+IZ4PYnRi+dOmH4Z9ouWFQbeDwX6IwCh9xzs9Sl
itrIBMlI0uah5dlX3fvM/Gvotxtrv+k8aSRnQrxhm8QnTjjm4vSxzCD/pvZUl7XS
KTuSbuAMwEe1OsP5PHgkU0nBC72iMPmMcAAJudOJqyyBErSRNT9JqPC0X8hysrFN
+RytCUi4cww2RIVdQ1HZ/rNyAQKRqvDoDTcbHR6fLTpnUgEDbDlyshFvqFJfV036
ATKZFBhNh2BLqrxIwugJOtY9mQckvthrDkDjVPoAi+78cvhjL5QScAeB5L02IhRX
rX6JtWCylObzyjTkytpnuIBoJXZzR3iVD9Y4beM9MiXfDmpRVweM2QSEy7wXKCWo
J5b0ml6GZtn9P5WDKKzgG7etzGR4qVbNhNJs4Sly/eLNUXHISxSjxMcooLE097KG
efN42q1XTf4qUpYpI+S0Y5ldPvASZ8pUfcKFZ3MVLocNdXHfp9a+Z0aozp4SqcSj
UV4iRjqr3ARJwiGTl3ksJXpDq+y2vygT1pmS/7u26RuRpgh2WL0TzrldMlH6iY90
vAZcxs+ITWL9Re4oxkeCfnuYPWHgmGssdWqXRCWQdSzvgXlDYHkohQLbv/uBWiC4
VmUSm8G66O6qHmPrQTXLd18lfNzo3HFq9cHHvEKPAMw6D+YbECZG/9biXEghd6Ob
nGQCkvSK7OiErlLepJjLX/UYwd2nRqDVHL0MuowSlLin6jMBFzoZ14oATJDLT2HQ
9cQsAzbhu7W8oB0c+6zDZRGN4TzGclaDQ2/89leKexAwId+jgnPGrJhNB9uVCnOu
lnPwH8s43GPWmFG1jrJDxY2AZnyfGTFFgMNFdSb6TJv3hXYDflpTfGgljNWHMik5
VIPM7UHj4i8i6PVWPOzhpMEE4/lg0dPVj/E49MpFC/OGPSn5kO4rK8xaYiS2chh/
pIOM/pt//IHmQ1VYylrbsh5eMAX5QdYAKX5vIDNO8Eaq8tRae0JibnWTLyx1wv92
towb+do8GobaHIya1eIHHhwhQPlU5dJUH3V+Ap06zqtDVwgRnXmZ2TPRW38gq0Mj
y7Ul7JAwtol87UojDn6Ic3XqLoYxHywzj4IWxGazECTibmvT6MnfIXIJ447hCh1K
v/5/ZYpss47Vqzq4hjAsTLM5v1lhGl8aEd7uIDG0xB7FmXSEEvwyrJCeU5qqOYWz
fjL/wWRtbm6r1RzsXBcRPkBgh2ufmIkUXIs/VBLc4q8Hh7hbb7YE5GzKhjQo4PC3
wNxkTICzdPauAdvHTx/MwG1HWvWt+K/xcAkxq+NxjatwskdxYTrOU5n+YftKEJyp
sCQgkWrpT9C49+VYkj5WbRpmfazARjmi/RyvppSkvwvRRvN89zuhM7xLSa2a7uub
KSyS1ete9o+WXZocvdORAOYO2u3aepS1/N4dmI/BA26iWqj1lUikw86D+2JDG22b
WbPgXAJBs4CtVOQbKjKhomG34ts/9PLuw8+eCkNRgX8XLCk8N6hu0iYrVYdoOQGs
Kzy/cWotHuuf1YeArHw9kD5RL9CCqCrTUUNGJU+C717wgeYaa0z2RidwwdosCXT5
kpXUqWCNCwvZPxiLY1w4iRYZjnmqupe5rrwe3xxG7gMwT18E2LSzMkEOT2z4E7AS
OxA6nJTq02k5WIujBVJvM1oPVtETaL9IqYOTAlla0VXLhXmF1sTGLuThAAbud2f+
RdlsMx5PmWUcPEdpKm9aC76ojgQ+uPoO5XafZwEUFBXOR2BkeIDk18jRLW5Tnz9f
gsjUQGtRgPLhrL0zH5qneZhAJOnMy38O4LySx7TvXE62SgGlRmhGdqIqlvkpEIpY
weqQQ5nFc+N7GsFCOaZyKgj5Eu4BbGDQcyDM25t9rK9qoMsMHSJJ0TTtzNNofN4+
IZZ6KdFIp8uC7Nor8nTabPwb6ZvGv3nFtM3MH5y/ONHuZVZqPDlGXUUXzglH+Qi6
Gi2YahBJZk1mhBAqB8wJeYSEE6rtOwj/gT3w8DEormjm2V1P9iqn+r6+pxtFtIuR
4wVuxU2aCWxSFA4+c2pY3hC+c/arUerXqJlPsWcz0OUfz4BPocz8jg4t/0WAg5ME
sfKDGMFGh6oJnSF6/hNbp8GrIWH7etZMz2n8TK8237wTSz9ixAyOg+gCCmQ/h5Ws
wLRCw1uaYXpY1Rm1tViP5nB0SyydBBiQF6cNXY56OONjN3/P85J3f3AT7XT78id0
t8xzxoQdjMQCw+1uR+TqZkfQ9yDqUjvhSDzIjbsNcoQmm4hJGwwyEhlB5OaHAfFo
U9rBquwE8A4uewBXbHxhb1Akp4ca3sUwLl6GxcsE6VTjQ5248vvh+RO7+y6WI2YW
D+6aT8puiLdi97B/yR7AwNZ1Nww+h5JLO9uK/jMT/hQMuWxteklszy4Xgx3hOdPr
b22GIPM//DjZ9CU5bIhk8SvT7qDYaVj/OTACp6s7eqeZ/R6v93MrKLi3inX7LMQb
7fcG9s7f4RyDOE5ggP0a2H7PwWKnS5wywWb9kY6q9NoMFzG16i5jyQS+Z2Ja/774
pFiGXeV4SNjbf8QOcJ2xWEWKwN4YXA6DXpdTgnBJPQGyBjrKulbwe0C1tnEnxZUD
VqkelxALE+59Xrkm+TgyoL5Xv0mFjUhVBoWjIsDf/5VswVz8l2yQ3Jtlw6jmpPeY
O3uNe2qrllbLm1mjRP6AuVOZiG2dAoPhOz+dsU/7GGCM4iudQb7wKnUumij6HqjA
l9jxj0widPKF6daQl4Q1ZU7yxpHopi8eq5a+LnedBx9AjmVRD4L2OJVBBgJPYNgy
9ARD1CerW05LFxNSu99V+1h+55m+5BcQjedsN21YFlXekuS83fmoeUYxJP0uwAVB
Llx6r65W4Z3pBeW65ctzSvaA9XXWNtriygJOaR99eyYgO7OelrzOOrcsfFgxJ9Ag
nQM3EROyH5WtKotuF+vnX7qndw0rvgkQYflutOQhSN2VOHE+oJBE6OnO/UMgJsxs
9Z6lUFGe4d1nHyV7ZBpWgrh23TJXPIORHq+KwrWGyogZirBcsbCiNdyy3wn6myES
MSvaOlfJ3Te3ukWgs/mn5T3iJIUOk1TmCL6MCuzwLjeVaSD0yWnlKyox7fvEe50r
YiZD1BuwjiE0s/7U8BqDiCi++wNGS6AjudkDkWdCM8/wDy4cO3iNPt1MHAknraYb
ICodC2EwmyeyiClNmV7/e0zSZ128eIylKtKO+GNOZEJZ4qfz2+hB4Rqnqoiy+Lap
BUg4VI1Tl+UmmrpSkvmLdKIm8uCULICcnwxfHLTv3WVXnVZHV9RBuZ/4lKbiwQ6p
WsEyINjuSVbzLK5b7/iyRq+ChxiC28KGDryqEi7EkqryoDr+tTgnIm+630GUqRqG
Jg/KkO1QSO0Of0Q5d8PiGI7ULL3FZaAYAa/IDhJVWkXr5kefmy8GhAgCL4YvzLT4
F2jzWVKu41pPRY28TzNiOClhfgQMQ4yXo9cRPe5cM/t8Fd1yeFtBlFsj2L8OZfFs
WSPjhsaDv9lsmrbu2W3iIyc0j6Xto/xDOqVb3t226q+eCbokQiLUgQrkMvZgzOwW
RQSwh4fP79TfrK/lFxq0oP/AMCQVhnGmiMnXGbKqiVISRhP4sSpYcCOd8PIjOKTK
yyisvccK73Gtk+m7aN3N/YM3s7l+exgpyYTUp00CfBIpUXIfiRvoovAyxkdoXsuS
9zC17icZI3WIlatxswnh4gPPxn5aQjgbMp8hXzmRdPPfbK9dLKD7Uf3Mf47pikiG
CPtkjpHf8Muhgi55t6HvDZ1VwXFdRjsa6YuSn2qD6jydBYNptXOTMicIb+xmxtX1
ZIDahuuZYTak2Htdvr5bBmL5RnMB9wEeU5KWhMbJh8A8aj5oLJTmm+bNBB8V1Q19
mFyaFH8GWVTzp7LwmF/uWQ8keh0MLS4wCFaeBeDIzWQpaDsD/qFf2y7QB29Hyoqk
NPUbMIQMNnVZ6dcZ0NXmPnM4U5YpP3zanpPoziYdKuIoqYf6urK2Thr7BGVEOdc6
K3AKLSRPDZnITHAPGm1gyyfF6qOJVWaTuJwkCbF0/f0SAstvv+shD0+8FA0AfGcy
Lu7Tvbd/fqxJQCiBU/QTEvfB3VoVs8o5vp2Yx9B8+d0xWzh2Aa1n8R/GixeNohhv
NwYVfeQSos4tIUWEfmeoR02l6ZMy7acEXmvIlifmZNKPxtA2kT6d1guAagHuY4po
cGdHBFiAIoMCMfkUMtOPjX6AJ4g1bC6MXqS16zk5X4ZO22Zq+adtFVLaodt9MJHI
zffKfTMzc5xDgRgtV8ky8SCS+c77LUJRCmrHDWiM0Hjao1bR7cFTCg50vc/RtsOA
pfn1WakC/Ls/Mt6aBA9e2BqWNYRUpoiRiE+vKlIxi/UVPPSKM9Yrb+KnYPX6OxPu
o9nROyDdomoDkwSjf90PKvsdScNMBkt0ScSoNMtIe29wMECSZWM08Kx6eb+hERE6
YIQM3p/Wq5aIxr4tuZHItbZZaKPON89hLCAo8CK8L7e3RcOev4mQ7go/3bqea4fx
JJp2Lvs+5qx1vuG9zDRUR8Xi3PJylg1XKkIsqtp1pGUn7OD4AqFTHvDPv4FkcYJj
/9EWQOd/Gheq1TdQYlXsHXPTvpoOdFOAgx8wA6CmOZH7i71f81pm2YRwUMAtl2tT
geCQREDjnyqZXk94hr5VI3S5/x+iA78p28p2Y65z94oZddpGWHN8h5axhVZr9rI+
NY8RHCs3aL7TnwkLMMT0F4BbfHWhFCuHh0wkji/K4NNuN12nGKBOjwlb7Cd0YFkC
uATBlb6MxG9rdg89epOgJx/lOsnzzdm+ZZIjGCtHqM2VYq6PVj5ofyTVhrUC68LP
EXcULYnl406unobof7rY0VoOgKMZF5GS6UbPQxZA8tS8k+iDIi6JrxJcYLxwMTsv
43stkLGO8TOq4HSLtgCDqQfbElgJ8BL+j9UkO6JRm+T1hRwWfwXMiuBagwLFh0sn
MUwsRk3pF2aLOVmLaquJgZ1JRjOkHEEpeslvhpUudq6Qx0Tip06FbmJTwgLtDbwh
KPDT5SM0bIp0HHg+/PfSj6xikerVLsS2ZQR0TJ5QY/g1zuTGldQz5Kp3ZkVaDMHR
xv28U2j7MsQX3bMYzY4cNv56UNUNWs7GBRy3P0VRcS4QoY68It+TjKg3PrMZeaXA
lJuzIuQIaNS/9qlOZRKGhmBw/yqY9CegoM2SHwuk+vmk/oTTIfgVD6LX8E7nDmpY
QpW/B/4GLpjoz7wjEs7kFXwnGrOg7XquI/JdTNC6f0JGpEuUzYoExQgl87PafBw0
W4cA1wKZ9zx0xhQVstKGnH20GiN6n9fIIuGeu0Ve1So5zrH6/iSQakQYsSsm5E7G
6CZz92izXKoZ7JY6MngvH8d5HXu0F1FuOw0HCyOdu5BKVSOJ8lmez40BowFARCBd
G+EpOy2h95qddFwWuobfzqk7qbXQVMdEd+AxmK2Wxx5oViftWmlZC8+wfXPdRh8T
Sxhy40GV8ACRxU+qielny3Dp/bfEAWjLwEnap6tecSZZBKvWTZo1I3VYheRK7HnZ
RVieMKmVt/daYoQaW5zj6vjdYG0R0TnMPk8M+RdwMQ5vpT6S+djEW9fZpP/6+9/0
P58uCdD7kqtG7i3QXpeIhtwfxMqITI1Zx648Ul6jZblBh1tAPG5JG/TGU/NYzUx7
xNYN8Vzrw+4D4BbieJvd0UR54H/bWFqgxsNO3FU1bZb+Np5szolW5LvPmDMKh4xd
Xigr4xH7EkBll9lRz2q4ZdaSgH8Y5TjtQC9B/gud2y6YYwiTr7q6LOl3666cmHrZ
0Pd4w3BxHfQLL6y1xj2UWfxsVQNgyZjfTikRkwrYczKb5fUjsgRLGssos4vuwRo7
JT0rHFzhLysKIM8bkg2hZo7/kO5LOnSulDqR1OLbBYoSBS0d1P58IlJvmWJvsp8w
PhbHJWe8bakpioEUJ0qqe7NCHDPK1QzLyfQghkPRQvGtCQrR+9/NyH094hKBKFGZ
GJpsBSr8Q1c00okSIN0MxPMOgmjU7sjCU/kAe6jcOD6NGTAAc7wDJzq1mk9CTbWd
eNjcqlxVwYvgL09CcH4MYxMYIqAu5y5RqpOIcnhsLVU4KqGfrNU+sSkKVRFKvW/J
KeG8Nz35sQ0t/3JIHw6NDoiD893DIZKeU/xttK17IJhTU7ZBIZo7fPMMm+CCqIwz
HdymWjKLVCVh04OpDnXyFPvzWCFQE8FK69OfM9raajjT7ogE6fVMp5yQspOonZOq
3O2zOM+0eVBK+YJ/cyO+5A75jMKFyHy1ngcfxNYfKkDsvgZoL6aqKWQgQ8QX+fsU
6J/mrGYxK2NuygY0lSKoTtzLBz7fVELI/yRDeKpTWbhSwBZIu6p0D8rGwFCcQaeK
4w0zVmrFJV8A64fBjK6K2BZEsauWIz7Ia3+Hn92wX6y0IPVYYnHQxv+/61EI4AJp
j0xy1lkc/Qw3OWEmBJnvKpzqidDuDh2+tK+auKLLd5I9Owy24efSdgMYbB7vtTeW
TAUgKSImucdN/QH0Nc8xBg0lPRvmGjSQkf2a++QQFnv22UATPyCpU3f/x68cn9Gj
pr8c/cvq8f8nVC4PC/iOWt7XyLoBV7Nhd52bsngqs59akWgw2NRRgjrpSM+e+izf
4Mohs12Tl/9KePIDRBj0Jn+L8GH8rcmsi1EB4WwG7vJZrRIEGcekAQIYeicfNZMD
ClFJ/08pvH5BP4PjC8pvATfZkPanfjesAwf1idFd6jX9Bwju5frsFTq1+R4MzXUz
WO2kErfY/hHLFN2X9mYQARGhZDAY1jLibXEsWXvMMGIW4Ovg5tUvI7IkNGk2f8Af
Yj5pkwoGnWZjdFBELsHJ7i1dJxzkRWoiJW/gBSOQBxrm6XA7uKHQrRvqD94j6dR/
5CgJXFUQ+qlLJ9/WGZW8Quje/xt/omRaLxiHtrTNpewPt83b6dj2Jq1rLoB2nBMW
tHZssXAX0s7Sv6/2G32uVsNLi4L3EtQl0qKrHwCV6ajMxnvCYNCWLAc+Xtq4VzMg
e2ossuP2TUeCnbrhZJqhb9yfnIaPSqXH/2Z2jAX1yAwwezuuLXN9ZOPf3G0ISZ2K
sKJL3uhw4WO4wNA4NFEQJcMdUiknllxaZJ+4a2XpO4P7Qo6mmGuhirRF6DrIEPuy
n8AN0jhwTvGOnrrHyS056WBCRnXsjbaNla9Lnc6/7AlOVvzgp5/MSxWx9pJ5U5Of
D2lXtnIAemWl5/Z3zD5kGP0MxmOckfHaEHOOhyhkuSXMOz5jx4DCaddSb72TP3m3
Mq7niQCeS47O1/wNny2p+zXI7rMPbEQssYb26nM7jbUoUv5uhNh44LLziwtY50Xv
0qvjSawsLg7rY2zQkP6PHNzIO+hXw03sT+Slemg1J9kYNZu+Ll9rN/QC2aFADPBn
HTN+Hy+V4P7Kcg5T2r6sH9vi/4jzAPEePUKDLJyfVN/5mwJfiz0Yu+1Pk9wfvdZl
nMtWCJGqgR9L9pBvJgnlFRZVrUgPOYz9qZAh6XnafJmkKP+S/HWZxh/YDUkUkA3s
riP8nShsLpzaabYrXn7ypw7qCYXeQ6GCUS3d20dsfGu7uurayBg0D8Y7p8D6tGMb
TvDDYX/AS6pAUYU70Boh1AK4lPLRZvRN+3r3JogDtX98fG604Vx5laotAHpbvY7I
rM8WGzN0C1vgadqaArvc6liTiT7A2AJotKossq6yWBB3reCRiHvQXUc1jlwfFm7+
ItwsA9N67N3ONuKVNDLid2228RO29xKFqmsvCjpRQfiYXu+yGU8Jn7Rw1IkZyuWL
rkUzOxOIF+cGb/3VcDlI9QIJ4KzQBrI2kAe1dGjSnVojrPji5++va2MuMwCWGDuM
xaqYvgdXGFszEgEQx4aaQpco7B32csXZGmbhzODLQpXETMddJTACQ5jhZ/yU1PJ9
aYiyjLeHY6K9mS0iWilzb3aeFmqbHNA6rvQRJLm9dq2G0O7PXO98aaRW5D/RUfLy
rDYbmUGwWOBfXh8wH2CuANXqoSWbkJuoOVN5tnMtN/YtO1uIMSBbA3M9x7QLrzLv
wcQZneKZvY3RUtcY52D3N+X7Xhu5TIflysi2vefxoJZRpwt394Q0BCKgX5YQAuDl
1xq143gOxjNOXToi2f/htklPxdTuKnaHn+h6py8cs80f5B2+0/2aUaIahsLnJa/p
t/iuHrFN7ZjHs+vgh/6m7W7ZPTfgT0CKBxUOW151Hq+u2VgO4ZFNYqnsDx42hm/W
oAQw0JCAUrfALC4PzEV1Nlhwfos76WkDHVV7JlZl9EPIj2fUf4kQtEkk6AE/UrtW
WNw3TOcYjuzZsrwT/Y3SUKbIp0Z+Iw0JJEh71CINGZ+0cSqOw/uaNkKPR9NwlSd0
JO46BJ69GVey9rpILFQYO9qqrXhmOb/4tqACUOjh+dhG/g3mjWEfaVn00zf6+ab0
oy0ZKB0UMe7roi+AvW/V9vA8i6NxtjK7/FcLV4cDn0E2YO1NhSZTglyMdlm6xXvl
idWJkR3EWzWJh8LTYfBu5OF4WgoK3R3/J8uXE3Ht9O1gSS8i9/lQLSxaewecPPwy
ULdYPlAnJpwi8dMUkaYOIOmvO27r+iei+LBKVAzjJVzvlanJDoJfP1l4oNRZXb/o
iwU2V31IBMOD7UgM8WByHFSDKL42hfgOJYOtNcIWs8scpHYQo8raGla8OWxHKmsu
cZm9xkcEDAcHJ3od7qQ3radDZNiCaTghP7yYp3Ynr2tNle1b9II430amcCF5o3Qh
cpyBVj6rzmuXvHrELriegccNO7LWpuGEoSj/LiAsaB/+7u0MkBBAGiQIVkxh6OY2
1AS3AgRV5UGnQ3uEYaOGpJsutV77xsjweoGDXY/O75DL+hHrYxsatH77wjeDoaX2
jOVvMXJS0l71pauOFS+JNstUqCkmBtJHwurgj3Bemt+ooHItbC4o6O4vfPygiCWl
+EtsnfnzA4+3XbZuukbkaYKYB6rvme00XdD1oE2VbS/U1w2nAfODJR1I4AdIa03Y
lk8BWDqUzdAtPauumehlsJnJM03OOQ6Lv6RiP1bTrvqu27e5AdP4Vrtz0eK2mvrz
3sGT2ldkGNrlSqimBnCd3LNPoDAG4raoJL91+POb6E68Ht8ZJkxNf+mrKEJ+HnEt
oIpG8YPtv/LUOP3jBD5Wlp0t6patamNfaRQ9V0atoXp8k6pCnFZPkaE+mnRII3fJ
rC0xCZ8/DzGFhIRjx2SXsNIcidW4MlEW6VEVDf9/FKyBoYs9XTlXdNjG6FBP2qUr
zDV0QpTcb2tG0ddUP4UygmxMxeuOW2hWYUsR3MUffx4kYWtHS2cTMV5fqg4eXq1c
dq6W5SjH12w7X8k015+WfTTSyjTMSapRRPxk+Aoh5mFCdUZ/vCFQYXLmBbKT5Ita
9ZlCzp4jPsHCpNBJK550W9PUB9ga3BateFbAA9vcLSXqcihwg9zrLZuFqljR0my2
vbYFxqe2fb94b8a3mgKNB/YaVnBWLPNNPFLyUtZm1q7fwqbwxc3U8wmq313NwroK
7rQ35Ql3czX/gT7GNpq2kXgGQ/vXh4d5Dr1/Hn+IWNCQFQkdF6tkercaB0j7eOAc
y3wK7jmno2LIEg8UnhwA1GjERhSNvL0I6mGSWIAT4D6RFKViItud6mGo84tEnVkX
YYoiemoMgb9RdEzE7Bn6vR0pYUtC1EzU/H9xgr5rnfmXcuBz7eCJ3JSVkZwlpY1q
BVDQGTRqkTi5d+s/AbIOCrY7Rvp5g06CkEmfJpFKSqm5yuWOHj3hm5SbOfelnvEf
hNTfzCxc6mS+KDu69kizRRL9SMgU5g2FNNZT0KnZrsAv+Do+ardntPJlicXicdWR
+3knK17CcCRAZk0aAY69LBGVegEz3DUjG0Lycpeh57rlRfBLHwQpvlFUz1Cgl83X
09QS72atJHuY96oa7UXtVM8ZJSkgY7spyP6jk8V8CXsE1iCxvdXJUO+7qda2rvWi
let6IoWmEO8RyQUwjq0BJ9HoI2SlimzAlMk/PxVY0G7LjW/o2D+h5VY1eCwEguY+
Ogn/fxU2FaZoyZRwTDlF0i7t+xLt/crQmPx4hhyIcLzpNjP5+NJF9LEZ0Wh3uUvA
N5Ob5wYZyRYs45FPIY846SbzHAnU5Jmkpyajx5AYXII3/hHzG1SpDILeY7DSTBr9
zYw4CqufLih5icNvWHtHT2Rig4fG97bmVpRKmN7butSPgoHCpbUmRedNdOSk7o3K
k2M8V53AdfiUYZYkx/ST70PajMPvcKfNhG47liEBc94EBDDrqauBVt9rPZKb/DB4
2QnmiyMCdgRD+h75ODM8NwqbVFBwa8FxUlrmg4K6kX59iknyYmsDRiWABURFX6Ur
FO6Mbvtxf3ljdwBWR2a05vWB1DalKLn+wTHkrsCFdz0zjieIgWfExGrk7WIGTqaD
aLAfO24RPjF4Xn9Eynq0gi/EXrMDnd9wnkY3ha2Cd29dPuFgdVmgHTzZVEhRWT3k
sEs+OOs9X7mQPnEE+eM1nWb2y3FKoQ/Y+50JAActPfJeS6aR6EgULDbVC+CPVqsd
jBtmbImlHd+kU/U/x3mi7n5AUJYwJrj944btiFMDGhJ0H2gVxYzsKAtgogcZYJrm
HZ28Uec3IXVV7gP1NYKjWn7kdzOB+v1Rt+F+b179cATOxv3xeGWnAAXbjL6u8Mat
1MgR/RQ0R8M5zZICnc9SO4cf26TEX6dIDq9MJfsUPCXaujMwQlWhCfHveEtFMPsB
0fsZlm9zRIh1C6vFLcqPfcv/v+3UEElWV8sM4W9jiVu/owNq5FqvIu3twYfIp/YG
9zom+rO+UvDdlCyOmg3Rno0woluz6Hy2IfCX4lHxu/7Gt5QGfuABCUCwrftoVh2N
D+e5D2zUVMCgJPHfYgksFSl0nafk1ad1i8g6urK/VSGbJj0ZZwXZW3EP3T15zQdM
XGJHGdPb4xNAjmL81YnMPUdploXvn4zC/InMutQL0L+UxIQFzbmxpzLGuC2rfmF1
niF0na/By71RJSXY3scLqAvn9bSKQOteXT/DcfRNi/L/9tCVBpiswpHceDqXXULu
4R94ZOUT1U5aJHFnV9MMmaBXiZ8/in9h8w7qcsgToRCXmHqcJqKfJhrCZvJZFnr2
0t66rYZCJTxEFXyQNCiUUKxVb8mxyV/0kRTnLXfUbQrOqJCdyayQLBAp08d6RPzY
lbHOvX+Qsl5O8CWvc2pNyi/X1Q3MrFmDTgnvu3fKb/6aVPZF0RCg6TrAbvtCp4Uw
ZsUNbLdy7F4XXNwoIw82rGvBywKtJG1EOkqlQBTZi7rCGcOyfvqbUi5WxXQ2DqSY
S4rs/xu/wU4iSLOh+f4tBl2mj0C65SHqVE5bgHd3eiR5E1IrQuPpPT1OWlNigvFP
bBzF9sJ0v2TGtD9OOczRjrFSI6cP+KOEODAxVRXmvNd/JqRfEyYO5ueDIY1X3yGe
SkXH/jnIcGMkjR9g5uxmq8UZ3jHZ2rhTP+J0YrSWuHBvIgAMPjXszD+9d0KXNQ2O
F8Yk5KFAryY42uhII8knzM3m97Lc1tkwBfURnogjD6OEu4AAB+p1UiyqZF4wnoeR
SVDeh85ONPcAR89x3j5AnpoavYYyudEFSwA5llt7hupx5fq3H3253HUCjecxuT52
oO4vWtuyERuvHCRDDHis7ujrtLwL6ZJZ+F0hCd19cLslb5FRWVPgnac6Pq0M8amO
TWT2pEFl1kSp4gFYzLWV/1IyNN0fqIn1jmQNISSgwik94x9SVMMoNn8DIjojc55L
rIZYMvdOMZsnSFDXUK7VCBuRlMYy1eocx4qroHHdCvYgbBk1+cX85G3T43FYNShY
hKiuhDuNfeI1j9jL5RoZSlRGrKcjd40rUEmSO1gQ+AMWK1EIvNJi1D6WEvGpmtYi
BHpqWda2rPWT2gqij1G2lpNIwzNFtQMViMDziUgaXcw6ktZ3VJcfHwX8zlxsW2WE
yMnKpGCoEldG3zmeZKUEO2Z1WBkNCbCRYxkXkXCDYIESEZ5lGbB1Q4rlY7gqzfpU
AxZfQplkOg3qujdOKNFW8tkRcybIKMoGXNcAdGVvIXPigqpUMfQGyza5uyI/woqw
AbjC3sCkM5eg2peAHFh2ixsWOGjLyeb9t1EhrM+xNtusaCrPT/mAJqIuj9nDY8zz
Ue9ziEUGWXd9/PU/aGeZytAp+I97uQC2lebRCVhHzZh6GhTObkGGIet7QegoHthr
y25NJ7z8hzO1XJU9UOVL2G7eoy2VyJwffWrjcV9jJag5QMA0j3VwQG08Hpw+93PO
X/eyr1TKkRge+BL+MZFQyuNihfa3y2qgFXrSXmo3QcloNnsprbEIRwsLVQIC/7F4
XtWC3l0kio6yvZgKyLS2lr4/F8pR3gO4kbzLV53R9OrsJFOvLFKqdApw2pHFp3AJ
qOnWxGt8mKQKjN492Cgv4T0SWC5A/TMG6sUYBkxUO/7DK0L+U1CDpOKUK0oNBXyZ
IAjWcSoAOZDSg9H300IF3OUmGRy0A7/vWDFmU8jVz+l1WbAM4H4YceYQWbZFKS5N
nc2wX7TajjKyBlBdUP4TzkdNBo+k4eLf72H0L7dNohDEbl7vyTnNwF6ds8qKll1J
pD/99DNKAfbIuz7MckwMEHih8tgURzKWVDaN1PyXG3q58p6nVV/f+6AeN+lXALVO
Qok3QKEowFa5H+JFAhxMcg07coe7a18zmTXNnWW6Rd5syw4GE3RcoAD+3PK75Ccn
9yk+Eu3dSmR80COMhgVAVdL0YYEPE01yxb40K43fiv0JY9gsx1M88pIgLeiHEWzM
CWMGJ6ubIXpsiWpOdBTdYeTavp/pcE/UurTQ8T5KWz70UJCdTv/ZJN3K51mCE2af
UDWSMGYG/Xyz9fpU/fPFRneis5RMQhjKPliQnBCOggZDPPi9Vg+UIhGw7UXGUXnE
Go6cPzk3EXftvN/43ESEkw4oruJVwKLzCgRdr4QtjkMIHgzInQOrG8l1vE9eKipU
mgZt65u9xm7SNxeXNuzFTF6pIEuksMPMnYAKiDuvntJTV60iXjxh4L+AMRMhinZg
jh8WHC8kwMPxKR9F+HgXZ3bvxYPBxBw3vqJuG6x7zaar3EJFQ/gAQrE6vIRfuaT1
bNghwnyT2KPbvwtANbW27eV487BM4lnou3GUF8vJbYhp0XRz0IN0N4hB8dMad/Dv
r5sUSLZEZzgO7UF6uqRo01HvqAtFm8l9ftrGtWIVaB/1X+HSaaObBOH5ovOyAm2Z
Hk50eqxBr1EiHnXnHT0YKCCkqgaVlBV/ECYUlh4XgW9PQzFfe8b73zBtzwoffCsm
b1hU0UKHMDkkHU/Z7ND8SFABFTgVsdCW/T/ggkf4UJXVjNrZ/oOpvR0kHPUbbeJd
I/RRkmI1uqv9V0q9ETsaT7jPoHEl04oTmQ/eNwJexu141ut1JTWwsGmI0KtlXR3m
DHEsfoAPohQdzi+03zyXdmEqGkAvok46YjpwvqLwORMfYbmaMPHl1ItJYP+Hpr3S
jysGB8Lt/VcjpRORRVHUdTFogAxA3v7WQY9n/cN5Lyt5+VsLwytB6y5GKrT5nDB7
4oOf1UKwjwCodi/o7U5i93QH6xyEqlE1ZAQrABAWZBsYPvdwvfbSLP/+r+bVDVJd
QqYdRQ+ezk1MSiBPo1BYupR7YMbaxORAgOB7jWRHarxKV9vVKD7oQPcPIejTAMyg
cW+kmWYGckFYjR+eqNLIMIHaz0v8f+0dLOXLFiLS8JnMI9UmxENxqEN71tBy2CJQ
o7b+Zx09vOQstv1Q2USBukcNNJgS7IpZ8czQ2CahBIjnOVFK9ApsYSdTXZuKiJjK
EGMAwiBCZHujXOmmERefoUHh1NX9Ye3llQMIZkwCmN/9wLcb8Y/qte6axdMzs8y7
Yjf4O+VOtYUUqbWh1gi+otsk0qmVh4OIFtJCfU/4uBBEvFyvhWShPLlMvrLYdHEh
kUGWKLqhPaRlLBhq8lv37gct15EDY0Qo/EWS0bBMTMaVtEXEdohriR4kNCJi0Sah
Xsu0G0syIYagxfWBz8RyLl9aCbA2OnbJvlH/iqWAkHHpFHrpb7zm30CocXW+P19o
QJvhJr6EI+oi2GFvwX+1noJkaMhDPtt5QogmfVGe6hv6yfbIzUAJZwunL9txXeJL
u54dzYK8PO80bIz6NVWdDD7BDUCkcu/SXgM1ROG+wH/BREFHcz58fpWbPvTkZ2Cn
lHZGhmIy2+PHBfYGQSpBEnmVVxcOXaFQg2WbjPsoLu4mLw8FsAY4VdIpq561Rii4
chXHBSTNVkWm0sQdb5pl+5DLADpCmDeyp6R/tU/Nv0OxGPV2ohB6ao/WRy56aJsk
XHDHtb/mjRdtEb71WDncg1cLdQqNlv+z9sdyZQKn2g3RsTQiPaPW12wDj0SuhICl
UydgyWKMlxYU5cxVaBCV8K14Lp3MB+W7pTk3ehas+/NytCqLms5cYmV50KdlV8Pv
uP92QHNHRwsEb5T9UAuJeQ5KROoOjbMsguOzTqvVyO6Y1L9fZxoDPgzhTdkklIlw
itK7yVQaZmtqCmpVwJ4XjMpgtgqOOriCVAud8KGbiGH1VvloRvowryXaEJ5+QrUl
x/JEb66mCPPUD06Tf62UDyS+J59c/iXXWz8966W1BxyPfdNPvfkKj2IuuoTkNFNs
BaH3RUaev+52eaGqICZmvyxuueergM8LKNt4s1S5M6K0Rq534G+k4vBanOTUhNMs
31G8bAFPwmie7v2LnNIjMb975YMfJMpswsAYGHlXf1QdygNHj46sQifXow9Emz97
V4beqv/j94J5gXRuRo5Avmp3IMpDll3K4fMAAFBjoKMXA+70q5UMw+xeA+Mdc7zg
AhJIqV8Kx2G6n0t6XVRlvjVV0SKNfkcDFndsKEqt7SF+VkFUfRlR7MELFXA0eT49
76h6rTu5+5mMXPwed1VYRSlbKMQerLZ7OB5glaLww9uTZ7NZtKiubPYhMWRQ+hdw
tm3PMJGGMGxWAC2zIDNxVxIyeX3c2/gQM5eKgAJNY0TDdFjF4fPo6v+hH03EnQZr
C1SdYzjvlpopFG6kDHc8TmbSDXQCJSiah7rk3tBCjQNeSdwm5jmRRc4YKM0MaLHO
Y933S1wtMrszVXt36NOcG/SCLCdSsWuD1dFPvYGSyHeHoHYkSlZ1XlhWdMTtkfPo
TgInBzGYlGi+oMMe6Ga+AEmBbR4vSns3o9LXIMkc7H9ZVLjT+qmsETPI3gcje1ar
dSDNIwc6XmwOv71mX7zhnaBtxX8x5YkyTnznzrBwYbZxOkUElpSC2mAq0unwwuSi
IGp2Z/n2I4pbjjppS8l2zJSXHvbFU+/ZCHQlvYhSAhqGI+HGzoJa/DyhuCmKGw3B
o4mlO8VyneBHZ5L+fQmSf5Fx0jLnzGD7ygr2vPDP9P0mbo42DaXnQYXyWckF+I1R
QMgt74RXtzo7NuWUGiSwzGq12BG+qzer2r7MLyXDUmlhOaAznZmvl4oO3mYA67Xn
LrnGAjpP/xFszOqZ93we21vNe7wnDK74fH8qv+/gTdqcJkSsXNwHuU2RDCCMVom0
Qnr9qjfv2Tp6cpFvU4+WDYk+crdooJt+r0Q76Ak5k3BV0iguriomvYGdj0BHz4C+
ussIjeuv2iyJ4JLSOasrjPNN/b/VjL0JC9EB0Aaiu3CcKDCipa04QaD+vfxjj1w8
Xyl583a29+CViPfoT3I+otHk6J4iMoZ/v46xWuJT0NDkYGH8kUWA93U74zBvzocm
Y7ZEO1jwlaBJqxHaPVn8xx0VP1AfsEOmsOA2sPkPeqight/fgxEn8WvJi7DKeIPK
9M+j5i3z8wHhmWOSpNdADPqgS/dcG3j76UGi712wKqmr7ItGWLCOVEG53rfftVd3
4oF7VTbwnc2IVinLHFkTwzhsMdOqL/4q/UDeHLc7znhjLxTb9UaMKPA2K124Ousy
fgbpc0eqV6Bsl04VF+3HZWJuqenlEbrHXLSwY4Hb0Xq5iE0xGOamySIpzRYR9N1l
rz39uMfHRpdHZr7XV3LxcJapElCqygpxUjFOwK7BiNoCBNjq/mUKSBFQ/pzVx2Fe
lVEILqE9m5qhXqoHeY2HQDXX0OfiXI0owqPfJVmCUTvWr49BsrPp2dy2FRlGyE2T
K3uBeFnZDa0WwOddmCH18BlMNJqFPfFCmRXeNOrIffCkHTZx1lK1OthdPYB83MT6
AVLgGXvnZBau7LsVHg+RrGRgcr+QBM05AP/ka3X9sbCT5oyfegTWW0tsiuGj1Dcf
lm5LQkHo7bBYBQ2TQaLFFGWXz2nhlumGlJsSUXcmgctcyw7DzL4MCdSydYuk8RN8
UlW6imnWoZ7fpDw/4G0ljV0ss0yuzJlqVUv4wTKN4LyQz8fTj569ZwYJfm0i0r2A
uPW/ny++eZZI6QBJZnN2+hqFHmUPuC0am2FaauOSlyDGVxxlg8IPFlz7f+DuGDCR
pfbQGtmhUw7HPREpYboS0Yx/VBNe5JzKg1wRJ54AKIzGzimsy98gMN/B8HWyEM4m
nkxHSoWbdLFA2/03TRuX8eE3vWoQB+NJwbH/4gDJkGF4Z/z2jmTc1GcOWNUppf4J
135ClaNJNND7LXklcQl4JLy4z5L333GljirNuqM2576JssXOlLi5S3KgYfA+Nste
wG4KJnXJK32kcxIWigYbM2DVWWKZT5YXYkmLHvTs0S9ZxCiP40q+VgNk88xNwq1E
IoouSrGnwuh68E8zgyCSJbBe0dKjjHGJprU7w8Fr9RAb3xoLQ+BKx6KNmnym6GDw
x7B0yaYys4n+3dDjW3KrJmyUpwjaRt9Ea23FvmLoedMvxYSZTxSCl6kHmXmZP4m9
kWHhxiT9i4xI9FhvBSNswx683ASrNkDllDHlrEW0xFYxlG2BFJOZenUPtdgmSZm2
CVxcOx5X+n4THvotfjVaCmSjmyb6weFFSHAlpxYXirH4fEh0NEGPpj3TT6jWVL4/
4PwTrSlbAEAPMxg4Sy2OJJx/s9xzDfnT4ZfpWNxmj9gadvlvUP0VNPWlZ0IOsoKH
yZaY6Ke08JP7MNXbY7m72W1eabgD4lZFdsiZKuGESdznlK061m+lfcgXEPIMz2UH
ctMQdOklWjHTmNB0yRzWxM65zZF2xkxgKo/DQk7CMNtXyzszjhffYlVCMEWWdpT2
laDeaTydRdSvwrNe1fsKGY2TDYacp+VUNV+8J0IPzZrwvmmLL0cyMRL7y+CM4jKi
OtUuhhtyWHGziRXow8QKXXS6xihYk2/iZRrNZ7WSw08Pv9GpqHE8AGRXhRvAY2cQ
98GkEUfT8xHscxaiw1a4N7gUkLzdVHJ+w4v6jLhA1nMRO7CgIdX/kS7lIBvr/VOc
XX4H9eQD39zRBQxDEj87nuirqiJ20sbSFvovBBvgdbVaVrcrWKEHFLmLTzM9Ykdg
3LokuccyzqDBqdL5ZaJpj+vdmq+x3/D2ukrR6jQwrLJ+q5vvCdKh/pzb6J3CGkft
tykKf0TFKY6D14An+CyoQSPe8VE12nhAFKvnBh4AedDcrVRoa0d6WnANEtyLMaba
kxQO1/J7su/CKRDP/hzcLMAqviu3U3iLg63/cdwUCZ2t8aGKyPFjyte9b/cbamz+
oaSzgnaVCXLYPezLOAm4UsxO+F0HKK/ItJ65Nito3LQGSof2f4tP7EobS2rd1S6W
DNoRXayz50XbPFq75UbEO1WyFELEFi3jQycDnNrtZVYnCZtfJHi/EwWIm2z+wAMN
yPQWg6RrLmCzSlHawoBAWSOeeYUXXtPXVXzgwZPpjK/J3/grPIj9lBholTW759jK
gh6MVAuOlSj+D48rVe5o8GmQR0bVV2mIwaDqyXh65FLq8xVlYekZ9kZXn9MX82dj
7JbKPu2mZS+SobYCxDOdhIFQoIatEVLKH4KalTnHmgm6XFlF/8kbN62mzWH1ADoL
eis89HLTaO1uBrowNxVABWYtHUMLa3JGZ3FpehWuRrgg8beKsVf5tw0s0KYKl4O1
YK1/U9UEbX83a66UAYNvOxq73K8ToaOG/SvTb8hCd6W2Upeo+heFUzHrJQkuzCQg
2V9ezB6zHVd4nynUDHJIAsAVmX86nfEjgK9k7FoFfLWun2cYdquQVeE+sNJLzvzj
fDXHbgd2DTJjdkPf2vtsZv2Pjla7xw4mjkd3aiZkERxcqcM4quAtqL8YEv3XvUvH
J6skf7gw24NCO0ABpN7VPegIkFaQ4Fc4Z3+CTGeMywCKKpR+wZeZtNHwHX24QrL+
VxruIzqbY7cR8uZutkzdcWkhhSfu56ROlQBYHakSzNmWcVt8GCBTmH+wxusi+S/a
wG5o8QkJJkOX7+nP4FbzP2gpTktPgNPJo3HlNit31cYZ4JFkYwQl8AlNsAK7wXMa
j+1tg+xjV6Na2B3cdcPckSxT8yPhrWzpvokZJLoRsd5JKL1rSlspAospnkarO9NA
a6QCjtFyeejtoGqsMHBBQvd44slO2CYtoS9Mavrt948wBravR5QmY/Ybq5DVAq+G
81VeRe5s6/KoDGK+BBsCGG7+dVP0yGmYjX2ox2ueCP+Ly2rXNPCNxFoB0NsXG0if
THvjatQJteBZ9rosZ01LCYf3wXzJyEGVzOPMAuwivl9M4dPYlkjc3ZKw0o4c7+DV
yqWislhmZcMtJvI6wGiSYPwb5M0LIKyZAVzE7lxdpiNFSQaF4aef/FlFdiI0/s88
TuQNHusUgZInLoUsGsGpFEjJc5BZR/PRernCmv2v/qOYgYCh3blbxUXLYo+QAGjj
SRUraAOga/D2dPOxDn8I932P8CcFvkHx1BzjjeJFLgksOc6+DMGh8gs1bcsT6bSk
q7awwR8kiod4mr3ESBaHjulbzhmMlYaQna2Kg4PAx0KuJs2XC15XBKQNLyVRjilH
t9fuv0eRFquKb92L6NzT1wFdVHZcoxAxQNyKvaLU13Wjtgy5/EMJrBBA2iysT1ic
tpFukH00IiWUVdc9fgYbN4IzLisAarQt5Sg4lIOUn/GZZxKI5IhISViNycUcah70
D+StLdtGH8sHyhcWLFf75aeROCo9ebDeE889w/FX139Asu9nx0G/6+R7H6HWU+Te
Xocf8858yWest3tslIsWa5hVglCExLflIAnAr1cVTcBQy/UqsjHspm+4B2PdRcoA
nsrEivqcHtiquBqQMukz9wXuE+tkmkc1UlFNUveai92/11FxCXylu1JRFpViTJwN
dYA/RN+OqDm8wqQMAuCitsakCZkR/z15nT1bmodrzkagQoJK3bXbfyzNjnZS+bh0
ccnbnekelDc6BMmwmlECgePCTIZtUFBm7JuQuP4JYTUhT1lYuPfNq/pJ74U7Z8T5
DGd1m6tztWMChR7A8bT+WvyD5iKVbU1cOXDlhoP3hODaQ0mHkIRVJ1jBFAebemxL
AobOAoKCuGMxi1oPqvUuMBUHWEHQcoyzLCE0OvtdyDnXTu96g8aEbth98hRcpVJp
rx2dg/FOwuzhKBA8FuSzetLpTcPMAwGiDw61ghvHuq+IjC7yqDHKMlIQTTLnCYe1
Vj1495tFYKxuxLGHbenO1U49xx6QnTyN/6AgA1a64p5/253XqWvLNRAC4MZw4K8z
DIzcxbI244dqbdsTvmj00iyMCYagf1FwprESnL5MjoXo0EC3anrBABFSTIweoEbk
x+rI4LV+Dk9Ov09JSot3HhZvFZi2y9ORKngUR5t33ib7cCam9Lizj4gwBT87OsIR
gCt1i/cJRsnxHvbgt9aqcHXuK1+UitTQ/A8Td05SUp0yOHTW4rVk67wGLGqAJpx8
euHg3J2Yh8blSVuT4vCFiiuoQWbyM2CA215wHVg0DI2VgzB7VUOToBOywKl3CV1m
zARvU3rHTqrpOmutxpQrCyqaNy2nDcylEGW6TEzeGYILq/+jJx9oayct9ziL3ukV
s5t4Ic0vW5qQStvO6jw/5qNHZBJ4FfdYbQt7DUCqp+1eAGYo42C7utGQWVjvVhzD
1gI3ErprDaMFHQFXDF6IVcSWMdwY5ymkxZ/cFroe3BIbYOS77GCXSqBC/GHYPR6k
tKGdhgKfP1HuV1U63SiJArWOhgacDOYS1/9SAIGzy6AhZjcdaMSGSw26pNdVuOg8
LZHS4IkqzNdYrRx2Xzgf9Le3x80k6e1iBeDUc/Zy+2pzhIVTLFt23/i2/EYBXjGq
FenGPm6ucQtS42UCLsskyRK2MWXwsvvv25SO9Y6DajCWBFimiP3aALPHwwN58F+o
uaFIet/Rtb/LFojBm4OyhcgufLKQtrfTcBuh7hftMMOhh9Wl1/bh5QxByxCC4Mw5
NUSyAwRCps2LsD/8B0xZJmiMQeQVE2IaoKoWTUqcwOxgPJe7WPT3cVsqb4HG1O/t
JkEFOgCmukL/oIVJw0T7EVaztc5MF0YG6wA6fny8WcgmVDJ1jUL+/C2bYGnczZ1T
YwSf/DPFFvvqCn3y9OHF6cBH2/Sx2C1FYFcu7Ti+tdv3PFVID4ZcZsJNZIkD17hU
JkEoRZrHHjdDVrehIMiLxVbBhvUwLIaAtXhCMxUwGnPKhe/q0CR7aKQfI+uy7OQt
aGYqppy5noK68F+nZJVD1YvQYy50w8a3zjkPCX0AxyV/OyAUQ3z04vkvyMtjjTLw
xrPutW1PSECN4WgujDi44ZN6OIhXdBw99FNswv7gP4zqK6XxGud7wc/mjkVZq163
ZU0qa36pnc1rmlNxpFKDEWkx6Kho8n/sHRCt9PhnbKKmalT66UthBZemgNzOzeBw
bbrhcNE68GsO2uSqbWeYvWdFe1D7BvoBoo3jT49UKq6vud3Tk85wScIDhACiBaHx
zV7mqjjOkX0Yzjeyj7lTtfWdPPivldqStbsgcjuyCh/elauU/o9C67DuGXaHQ1Qa
cFWaZOZ57r+jrCWvz1+2SOPFOGc5N/OAAi4CAmS+dnRSFNCk/Pt8N4Q+Xt+WFz8m
r7mWTH/shmml6bMqbcM66suxPHSdNiAor6m3QdFg7DQcjRlu+p/6zY7W9ymT3TRj
kOS5hCg0liWxzYgkKgVOF8oibNSEMkDfWlQEKqHR2LloRgxk9EBUUPJr1whxR+iO
wAjPDHI68Z2n5rysY0GIOvSRygFmTxMM8EKLzdUMy/SImoS2EO7yiej8xy0R2lAL
yeoVT4+dlzM5XHndS1yv7c3OqQm0yJ9/tVbB4UGu9/tdAKZJeB4JdGUOmNMwtfd+
of47SjEC3NvYfl8L5oyWiTmfi1C2kBcHRQG+dzYw6ILEfSMoh/543tn6Zz0Id7vG
u4P41WSWHdLjzoxbuXWPtt3YTtJvimdXN6A43OLJPq8DUPDxD+abSWkZlfCVQwEU
lWtbXPhYPII0bymecgpMYqINpQ1qnR1SKE+y+Fo6lkknrRCn9qy7T1Mc6PJiVJmr
rJM5CrZ3QI7nE69isgUm4lH6dloG0DfmRJHj3aRScMBHbal/i/apCnGmUPlD2DgC
g2/FIvhPb/ibD1Urs7EqjQPhXo4lgEDNSRAl7s2rHnadn5pOFrJulO4ZVUtmMgzp
lrRrk0G6C3JWkx4LizggzQyyF3kdJpSPUjW36QELY9PUzQHwpFBYUQdSrKSVcztg
fZ2xSBJUPOHPy5P+GsxzfnobZNoz+OlQI9J6QVVrS6IeMA8tosL8jjJPAaKxuIly
2pjoaqjOcYD+H1UUGlaxMmXnWQfTV7TXFX4EvJBUfdvPZBDobTO42eJmFO7jYt7v
h7+ZtzkBsGk3bqraqbN8HG9pPq4e6On9rJy+dOWCQXWrNP5WiEvVYj+/56r6aIS7
EMVLsuJvoBXKojrKYkNRys+hq9XSpw6LxWzi0S7ZYyEDZbrb0rF+MLEcjGZOrSEq
j/F4krTWXvfCLgeZCkWhGL8uq24a8L85WAC7OKfTiRR4k2Hj7peDUrKJvCHzLG8t
T1QsCgnjq8EpgckUS1zy8ROzWf6uL4FWTmjTFDqSCDQ3UReHS5J2w9+1S5+brXs/
3MRgL0gRmCyEIU/GGRIQ2R+Ym8c8BdpjMN3c2MZ+LrlMu/nYYPeNqeDbXIMgHjZG
4T7FCH+oRKW0Gu/R8x6GMJUBEfAuXntKnyVcF5yYw/Ah5ckGyzKRxbwb8q3A4vSb
sH+zU78qGfHk8Eb/hupmcRba0mQLBXHiyj/5Z6qk3IFoO52FFGMz+VSNWjW3A2io
eqlHECd9QDsoOI+4hManmk8nH6VW6y759z+lbrJ20ro13hNTNuJKs1EcPdVRKn4M
qC5lyIZHQInk+R3YXFnjiDTFoMP7+nuLeEUI6pNmjUjtiv1vu0pvPCjEE5yuNMLt
tw23++UckmUG5FDy6bZQcp68ji3K+U7pC3wAkLTO14vdWHBd4FawU7EMZyE5xzDg
RKF51PM8RR/NYtKbhsnl/UYDapBlidvDBxFLPv8eFtQX6/uscwfYmwcFjQeCfYqJ
wG6ykmh+thCdHwR/KTnjkFjHCxgrbFS9wGmYRSssmokiynmpOHMVDGgOPdafgmNo
cbJNtjP77dO1UYqSNLLAuiVoB44R2yWyZmB5CVaiaJZBVOx7XybRrIEymjQ9D7qG
Rxbjjqyh3vOk3xT1eOI4+rA6AXSQ6mt3mSC7pWuJuzIoNlQfR3BOw/pLHImSL58z
5SSrb2nb0tVE91CRDIKx1V77NXlfH0awq8iKGSNdM9pWlMOh7NnPSh5cUZlAYNgF
0WW7Uh14jJ7yuFvnmMJIuAyi62j0Oaau7R0oCFHq36ARPmnHnrpQDg0xWgP9zfnM
sV3tuCgVOLR9tQCWR6JsgkJcBiqVhrIMkdqPbmHNUXcohihvvvTTRBKuZF1T3rHb
e+MeEOSetccsFQP1bxVulm5gVgL6BvlyrEiY5urPcllXpajONtRqMXzlbyc86DvM
vJCR/FcX0nDdGRRDxa0jl0pEGVSWH82EVcnt6Ol85s8kV2DkXc747LQgAuVC6A+m
3Wub/XcPDUU0Pa3yfaGg/nQVwDSMYsiYoG97IVV428vFhkCS7Uc3oFZbMa9He6zZ
/Vc08nwh4LB1MOybBJfvtWqA6a/hTWcTH0UDXk6GGr0YHuoZCLtSa7pVC4BQWoRx
J6RdyL40XTD0qBiLig0uqjaVdWC9UZrgbV5xddCu0IVx/AsjJL/zSJB53YYhbXxd
JHeFW3dzkSoI8slExwigr2nucfpEyObRE6eZJcFt3OF149tnrlJKlzEcbNEJv8VU
YvJmlzrAGnWuF+7dkhTu2qCFYuaqZC9J/eH6IKuu1L8mlN+M8Y4em014E6MjzL/3
457J0tMh1aQwSOu4iNWLeHmQAJbA43+hDubTEkXRGUDcEqeTGxHdKVSWlQLZRs9J
FrDW3+NNTq8/enBPsIV6eOltZV8FyHiugTH0qFv2n0uOc6LoHlwPLvq4a85xAIUB
o8iEkkoPJf1eIP7AKKPR2r8OOF2l2FhZEYs2y7v4OfbhOzSdeG+I2zs3dYmSrwFt
wtFGm/gn+ig8XyKbkv/AQNBItRDlOcnFfyckYI2A+ZZmXWmPkZ7lDzQaTBgpSg0q
aYIV+NcNTJFeSEeqJeJgvchS2Hw4smvJbRhE0WGjuwMcxMPei5vr8m4RgMf6vDCx
kTLsgXZEk5QAVHfuAUDrVLa6Sd3hVOZPCKlg5ErZ7RR7XyxIRPD1LJOfJyyOeAj8
iQje4O2G5vOtD5XwxUMFnjIBIPLHOVNUazD+d4x/4O0fHqHwzk3YCmo2vGxcT5O+
SllwjA6z/8R5kOGYBvXrBEBlJyzMAu+2AOxtjKdXOG/Xbcifaprf+IrHquztn18e
cHedYYrtj9ECQoFcL8F08uOZSZa3QDvcCj+LEfdQ5lfGeRrQOQdFZjagyyvpZeTx
mpbIaCaNbJGNL+OLEZviCtgDROmCRfoRu3YZ2r96TJ49ROWAGg6SEX4WdUozqiO5
Jzw2RYZexDQA+jePaw5rPOdxkMgcuI0ez37/c4UyC1ixUOKA66Sh5WOpM+kecPEk
TKaJzh/a8jdcD0dV9a5c3GZkIMzU7PsrlcNaDruQNbkmkn7JKthh0/Qg9En11bL8
tYZ5zCe25Q47gq77WjlgrgLTU/5ciiQ4UfOAwTNQmO2SZXGbNvgDmOlcPOTQnUKE
dsg26pbx1VDMSX5x8SCwJA7J8BqNkCIyyPBKLCVQYUd1NmureMmMo12atR4yup5k
gXhND5rjM9Rw32S2bl8pi/nK2oC7f0RMA43T3Hu7JD6G14iWhmf07tmFYOC0IY8Y
ZT3GJdkdV7LCcH628QZtDInCcTJ59go3ictQg2mjobq82Wa8/7jTkraktcFDdGa1
OSP2XsrtUOum9v88bRwkh0PX+q0t//mQ7hLYjyZN2R/CC1m/obAwZnUeFZdyHsG9
fDjGINTfWR4WMchoFFhIvZLXEMrMiWojBDeFlhndAaX95S55alm1/R5yIumWRc35
M12OF74HOO2Sj1hoY6yv2Wg7WzhLPWAOTACOBROnken3S340IZtIq5wdZHNFB72a
5/pPk9uqCbcuchS18jRZpMZB6068iu2aYrBZOu51pdoldupdXN6lShmPu5YFZDfe
JcjvRlJMJJAfRMy/pAch40REorC1ZFRA6FRXhvHMEMkvGnBS8RbawEc3noJF1wjJ
WUS5W6f894KYRJMyzxcmRFY9N389UZg5fe22afxaz1/Va8RHOGDwiz8M4bQyuOcm
4aXJgrefmUjlkUeg/1D6U1X7S39q54raaE3//cngi1ZITLtVDe0anv8pUeOmccXU
XCWMA2iAh28nLJllItSM4kCwn0ROsQc8uWH4Vv2LU1UYkTd98jDovXsr5g/B8TWL
Dt4Da30JXuaHlVTa/LEfzWPskYs/WI/2TAfigiUYuLeGtWWouELXurNnXx1I3pmu
i72e/O6gu/NTiXOJeDXZ7BBos17sBs33xcAUU8xXe0Kril5mUpDRFpFz0o/wMW+0
1kQnknTBlltEyjYDk267+eSSzS5Jov1k2xKYS/aSds/LlZ+DuQkcwP8yil9nuGoW
QBN7UeAHfYpn5LPrfmLC0UtCSXh8A22PnaUbMUEak8DAy4rBVOYe+5/jsEkCU/IZ
hPrlGOmENV520vp2xM+jtbdBxuYk82yTNI5jbOaVRNgfIqxAUgOIfe5Q/KaOwZ4y
HjdK+QDcMT+fm1f8bXT9dEGzYBOmOXYI+dEZBmmpkTozZr8ZJGNOKrPNgBIl5Zqg
qzu05qAPRkv6WaDhsB8LGx26Y+zhwlrjFsgmK17fT8LJFJ0Zvrs8Hfm12wpiGl6r
nz/SZkCGzoNJSXLkFPj/B7nbslMqzBjzyCpFmfqkVNf2cQvqD+wnnCelCQ4TV25X
qfYFb7dx4zGQced27Wr6wCATfXe/l4fHcQdEja/3FY47hQ9hqzjKaZY1wwUVKCMn
zsXU61g7P98+6i5qaEpdQbjyORsBWy5bR7nskT3su0hRkp3+dwIb3/zO7RPYvVaA
xYy/toMsUa3GuG2vGwtBI4ctsOD82AoDkJqU5ztOwukY64Qx+WpD/OpQaAAM+XJ6
PseyjSuBLx7Niymjjj9wXmdpo+AH8Fqp6/NAGzAvbXWoV8GTkqraoJuLp4kyjsMJ
JZWw1IDhu3apKsMiX5EONLXTD+g1laQxsHU1eZXltCyPIiw0qP24v1r/hfzl1BFs
UTgyfnrNcP0uil7jOefX1yhUvTdCmUvdADgmijYURikI0QbzLu+nOz689TFypX52
QrwqWjsWYOXVsiEYw9wTL8fF4QFhQ3XqGLa0MOD+kzJKueISAx9abvJ2ESdo2wFi
ATTc1ShUa0oLFSVB7eKS+mja7HN+eW0wX+fnAvGvXOGoG1fpynkEy5tAv1ovaHnW
sPzouC7lTMj9T8HVIjsZApaSLQKYy+S4pzH3T9QMbkZvn4hgOeA8gyQDRScvakJS
O56j1LouDrxB68ITeOvPSr9uAs4KV5hBXeh87MxQ5ySioVsRDXhVQ1LOuUXq1UK8
YYzJYk0/Me3fjdu9egSwCqM8sX2u8xV6nbVx4jQF92Bl5DM8XSVzwmRm7pX8PJ2V
CmqYh3P92+ynPBvz1cxq893Xk+PxpcA1Kzd130P0kWhAonA7qF5Ws/VhiMCRarVd
UBS9PP+1CODzzNPiRkUZaAPMPAmzGCgAEZ0dh5TIriv/pNE8nFcuUXOxOhP7ULgq
Vsj+hEINFKv4fNZ66fCx7SLYLi16XHQZfue9IzQmOMSFlSusyHXqkpCOppAe+mpN
nUofo43eaxOh3WN2qaXmr5X2pRzhP8OV4W0c3GyNVRTpSTrAlKgzjWvZVayROW2t
Ns/BLdNTj+r/GgI9dkEFEKZBs6Uoi5spD68ib7vvZA65YiZt0o1CejHLKLltJttR
UhO+5Zd5cfrkjpnillENlZR+B+ppP5hP3aWQSaZwgxieQmGIgwVF8d11FynO2lRf
KSSpXWC7CVstJuhldmmluA9Hg0L6aRXnz9UumnbhP5hKsNRwxq5AdsIKh2/Vy6rY
rLWtMClpSwm6HJ7akEnltBXCItN4+r/nMgXZAoIcfMXDhv249Ld4tR4FC15+n3Lh
2XcsGYiZ5ZeGnThWgqGMkEsHAP3qwBR2WJtWSt0cJA6vmkoRxdxZKey8pssHGF9V
7VZobd2fK5/JncL3sZZeF/v/rXTy9znPOl849+elEfQTJGxOPyMdDJR7mMEhVj3l
DKqnpXFtxUPDy2vJV2mkegRBKB+SxQzEy1e+Lv/t9fjeaoYcJynh61VacbSkuOwj
pKVbO8fLo63eGZIwES2g4+Lz0Q+sSXmvnb4gm5hIu1DIisWuDo31RPzUJOo0y5qB
doqikZIXUxT5NkhNFh09EduCtRAS2MrhBDtxGqh9yQrplJYCtvpcXV6MRUYPXW83
EYZewUH2QimD9GTCEtHeXiggYf57wQ31tXi5Fl96AwGZansiECzEkBfcPLo2s1C/
PuLR3H/vZGl0iHO8gtQIPmWRPAgV6CdqcBDFQafdX2r3Mal0qc0YKqNKRlFYy1fB
pbaOVkAcdoiHtCd0s4sHq/HVe8xOwO5edCJ1W54K7eqA4cdeIXnaGQJxkLpRmlWp
mDQ5J4IjDUBx1pxVv4ahmjXC8/tfeId8zpX3p68dbHTVZumC3Gy/Q6lrZnQfK7Uh
xGaS4MelBOMBqXgfNvlW2MKxE+iyV2NHYIT78HUKshUDSJu9pd0ONWaFi0e17rSS
gMFZAf+1Eg5B2dvZI/X9GX1bb85/Zc9KyR9ZBW28kPo23z9fCdG8kgcqsxoClBo+
ioX3ZriRqQdquHp1G7mwSuRHNEJ9g3uRPnBNrQrCaE+WaY2o3UXcKfDh9I5+/HFg
VyfjmnAua+Aqo6zlbPKdDkJnjEDshKWH6AYPQMePul0Y9t1z6h8F05zaKftTiGDG
x0WmuuRR2Cr3V/Trp1TUXWmepJRkYy0sDuTuXG7GD2FJykFVrGc8FJHgn2/pY/RG
PHJSdtRiU8HZi7ZWuSyEr1DAG30eOAcpAwx9psxEVdhbUvf8Z5OymFlTjhSFLYXm
o1FZvVvf+5/YFpRTbOKzHLA0J8kvefneRaQaxPLUBSlqvrfLWAvc+oS/LzgmzX/s
80G5Kyyb0qTQCxRVUUtgXC3E8mGTcRW67gDJ3vXX9C9iANhdSW5mrI7WUIUP4xhw
G1Y61G1HyGJfrn41MtpyDRH2EhnCf3wgG9CIHtu45zgX2cinGTjOYHNuy+O7qSIr
sVTTMNqOcFZGnPEcwpauJY6fGYTl+IlyitF7VHCOLt+W0+kP0bx6XfDZVc/aumWR
hsYtXSkRtCcfT8Z9PvEKaHEVXppczqgmmyKIuXj4GOX5QIb217FUuVqTlVs15HfT
LN3O3ERsDDNrXjxKQYqqpcyTtFX6lNa8iaEO1aNhbeyzAW9seFHwrnWtv9sHYJZk
rukgIHPOdoVv8sFVpIbkUNneIasRA8qsNdSt4p7kV81NWi8nfXN7RA5lTxEn4e7/
Vc3In8C9h+sdBBlKCWr9CMj03HUzgORm2YLAsIjPWYWApONTP65nxo5hhn/rhw3/
Rym6kT4u4A+MFHKhtslvLwqZn1oD0lFlmEBbgxL1BNn6OuLjvB28Jbe0a00U/CzB
SJmIoVvQEYFQc5nEq511u/afHM7KBbWaPZ+ZEZ+WmZz8EyYkrziOJZBiehZ9rXJh
6FeP606PfLvphheE55+Q+W4JBMAjC6+I8PAc3fQJKcl7OzlcCXFrnhG5w9s6kLrn
S1hutinFxE9My7r4AwdR/5uMcwHKGiE4GpCZpkbsnhLM+pNTg2tctYp0cp4sr+CO
4AG505K/LKdwZ5ncEvsflEs/RFQ2ZdeM+jHyulZzS0iwPt1F1qqRIC+WWi0DUmhS
1taU7faYOdIi0D3vhFpToxd+OZR9Wm0cz5OqoNw0j95C3QNK1QV8/IA0vDzUBMNN
KkaLtGJsJ5dgqorxCCxxAlZ4pv9tsIJrgRh93jx5dfdILJSPG5JFEgyi1mojtqRr
dXT+FzEBLldcbrSBeNriqxxsWldH04nul5UVBem9kv/0rSeD5FCYcDd++GCD5H6g
wmmBBKRpCfg3gEFswm6kdP0Qd01U/OOBwoCsoDGfxyyOvAW3ZNTi0OEvA+rKyXOc
nY+mDCr3Ok2DUuGFOtOIHJuIZ3osdytVgm8n4dfx8xzfvABe5+vBcrno58ZoP4yH
XOy0YPKnB+fOHbEpvCO/ZWSno0uN6lcFkaIAauT/0Zxqe86jes/WyBFfRzcozQhY
A1i7qZzP7MzsTNf10mxDof056/BZZ4Ni6Mtvl9qq/Gn/SskL0L13GSirVhTuGeKA
dbwGZcp3jAeKHDie3J/l/nDBR2s+la7JDTLY9vobuNadKaW+N/NjKGWehckZ/EfK
rGJzGDkBj9mIP5a8vDxaTwmhxijxSf1POOGh3wxNYkWbgYHH5QYDILXCW36cP1iS
JJAFaFE2O7APXuen2Z8RpWvq4y4/BC6KiP3A1wWgrjfblQvn2S/WnkpPNT1BkL3F
QcySFyXeJqvL8teN0mKy7hGuoBg48oLW3xL+PWlPqfcqghpRodDT57iVCJoFKZnk
VSzMe7NFk7OM9lB5dP22ZCbWdi0FR8EOAwrXnns/cRhp310ogbMaRMWoto2VNeKV
I3df0AoPgwTGrUMqvHow7vxeKG9g5r0VXBEwwPtDgHnqkTixMHUxSEx8MUqW91zU
ltnIKuRXHMjlDDvSROrS3+DHrRXqdXpUvptRqbHDs2PdKUeMQvo2XRISdSUkyOoa
CX/4I1FD4YTyRTf/5vvvqEjxmtRJIZrwBv46FEC0E+2CeN7xbmxhZDaad90Dt4db
FGEUE6PIQoXfmfAJWEL/jTYB0Ysx9Hr6u+QSoiSfKvZlUEtSMcb9zePtWs3ereQU
h6H9U+Nw45Cn5VYYdwjbfbof8UOnB/jtLD5iYdHnJqd88y+qQfJ31ydtRsH6tDOs
Bji6QtWk+LUwyc3LOlj/mj9WLVjfjN2srhBxPtHyqRpXJNYpgYlzBdvXXnWuwnbd
xHUjYNCKA1ic0pb7ZKIZULOnYpaqVsfTK/jVSpEx87uTnYIM+ZRypMPfeRU/hCkN
6Wl+xA2KWBn5IzDVaZoI5OLCRYLosmAuZS/Vuvqc+/37+EsbOkOcA/qbgoMRqdAY
gMQFVRK1XEuMDI+m2RD5yd6ghR9cxF38K2Up6mtq+ob+GLBcnWe22drJkAKNRhwd
PBTwAlYYAq/ZfRb+m/jniJhtLOxxKzGr7bEHatTKlcQkC/u9dGWNbFAHUY3cNslN
U0mEsh6PE92a24wfBIfYosFnPAhEU3AbKxBHArpdcm2ogVoxYkfz6VFYT4g2uC2u
VP5WENy3GEiKhEXPKGnH52P/AzRAyuNS2URFxixfq6LeG4KlSFMxMzPkn+LSf7nT
fn8mHIGpNJXxtdBz6lGybuBDU38neLX+BnRfhMrNPF59lS9aCJtp2KR3NsqXESCJ
NxY1ddRtzl2Or/81w9CNINFNujaJzw7xvL1RxPsapFqW0TIdN8yttS+TlUaBQt4g
iHdfprhMLw56m9Up5TLsDOsM5Bf0J2HpYfvh/ZCHxmLWaF3GShggISuZbO2KIHnV
0E8z75sD1Ur4V7uYjEGChC/V1qAM9C4JH4e9tlAQ480cPQDaaRbABC8VKTMtaxkC
biof3VzP29JPnX/6oBvN7XFdMngoSyfoB/wMSqk5N4/LdJhM1r5OPwhlcxgk5ed9
y7oAhFYcdSutus8tpxDXE/trdqksWi/xiB1pDxZgoiLsr+COffNyCnpYWawzAK8d
WQJFIthO0PASHuiF7cqRHdxBz5z0fehapPQioEvfrXcTzsmZHU6BxfQGwxvDGvc5
jtLoqyYbhniUQiR0THSrUfHytdikf4nNUX3Ij6r+E1TDaRCRnt1zX95oIdtUZoSG
1jGn8Y5mPKVQedXMv6YMg3BUo2QWZFSD7XYO9Fpz3PuN+ByRp57u1v48O3Mwvy+N
U47po22RLy29Aqro7t7ibVFUi35mELO5GsN8by8rzjBNX7pg/bVYEgUH++v9gj/k
9+LVwARU/XMBrtnFumG52TFx2JB1eQrsUmPmaQ6yiv/VrxPl/uxHewY+SZKWkvUp
BO3UB2Asjp4jVCTvpEdTh6Na/jio1wh53hsgrhATYeOzUniJe1tRsX0fTPtIkZjZ
m1UoAcplKIzWZ+rbQXBXqwaWZmTXcV3/v3Z0PubNvnPfaVxG5Dk4V2JbFdvIxXgH
sTe/Gs5YiLP0vQyrpj4mtBuf9yEiKbC8XGePUz0HpVXJC0T5BHg6UGNqFYPwK2rc
1ZZ+LsXOn3sNnnRjIs174LBOk0JifyBnlNTZcvE2funVUTK5BklVc5Csz/sVCeVc
T3uzTrbr2ULI28WGieNoYAr5BatLK0ZjW4VtHl7u2V3Uji6h+IkyL+0Sgclecnge
Nz+awB5mA7uT/+zK8JwaXoECvh2fppU27a3EFLvl1gQOvCnGSeRg3/4qn2cC/0gJ
JGs7v5nrACj7ipLy3YhB5Ew6XiRtWQu5FAAjbP3ahLDlhvH+fg7WemNxayOT1Wx0
iyNn/Q/V9gA3sgRCTanfb1WfhSt2Ngm/xyDn7KXHFhAr1flp5454+YZzti72obqu
mQOefL/sXW4WjhJYdbic0D1sZ2ty5ZnXle/JddXS1WIrz5O38/WMSXEYW/15pira
Zh67BJEOcOiI6Wyn/OIfWL7B47z+ZzWeCGASzOoWYBCZ/5pNUjAV6/LRswuzxqTn
biD4/QhArBgJX2RtoAdyE5NdgOaFaxIo72Yz4lYCnQLRq1JC3+PMZp580lehS6xr
fdMlrkCzlFo8PWrr2eXiVD4Xg9p2nuh6oh3KvuDaqLwwptGpoFn/mFPj7Q4rhccB
hnYRkrfOXodtrW/SDbQBizlSfCvqrLXeksnt2q5BqPnc6JyXkzQNSL58jqkTHV5g
W4W1zJM4ML9DXF+RdPojF8HTeQ6JxpBIMPZ2S7EFxz8FqTxkphn9v/zN9X+WHTJj
orMPme89XZTGldiItlMnOqn+tSddmYB143tfNkg8xj9FpV6I1sDJcewPyEsdjWRu
JvigS2VE8Gm+JoHgM+DSQTi98Na0ddf/5HKVCStfRSReLOX7EmMsuQW43UuAyA4e
kWs7IYbMenNyqRWNU6mS3AoeeEo00NCjuOEJvOiPCAJOXwx6voawPNHkq4/km/63
HFDyARt8dgWrMst+/NKnunaJcC2ZglfxmTU72PGgjgvHWAVSBAVanFSyGB5R2lu+
NxvkX5LMp4TCxxbCrgSky0OnsXFFozJgR4yDkauk0Vzzpo1oamNroP5eqPFwAY5f
bbi+OVZYb1gFEmSwrLVxypf5RGS0Fh84jGL8HZCjyLwR45RogbWl8UvPPklIkt9i
Kem5hDoT0DGdLWnTmU3LmiEWRlgTzieWw0oz0pgV+Euih/lHwgzri+QCLis8aBol
vbAqjwGAiPnagtRUl01ypfRA5ZygErCyehKApzjt7WKUk79yt1pxCQ9hpJ2Vi0wl
YBk5bFNs1WnPv3OPVsxwa04oJCa+sttXCIcRCVjAI1l8fxi8EuWhK7K/Ek0jkGbX
lNmw4tMKUmdoL/INydKeUFymLM34l/sgrG1eVrtVNPOLwsxxlFVYLdgRGuCqerdB
E9e6ZZbQ+UEzIR0jVnz28U0G9uHeDUPtA5NU5Ts58MLm/rvU86wNdeRuSd3nLIz3
JwrVaEMkjh/HamCfXCG8qY58NrEFQVaTr8im1cmVdLFzrhdu6XiRlw39q94onwY8
TpYbp2cUqB3I+WqOtTInrfKGAMYB7Ct7dUXG/nxYsV3/mSPO3LfjoWAImu7dim+6
xCq1qZn6i4WyHlAqdQKl3IDXv9angb5KN0qYS/bwu3cyJbQMDLLo5PA3Vu/Fi7Bd
qq++04E91sNJrrln9/YUHu3hc47clIGMO4seEYzWApcUdTtqsOAQOxg4CH5pBHZ5
NWxRZI9VJ5QzKD4y8mtcQmXvmOl1AhOs7IEki5oucRTXDJNRWE0EJz1DBAyOsT7H
1922VD8qQtJXhDaS3UZA901YIupHsFWvAS+en5c3elnfQzdK4D7yVOox8Nfs5Pf6
DhYpwbe1SwZvIxUn8dOBm0JVXEVR1OHoCtsy9blbyW64X0u77kWTq4ZwfjprM4KE
1rOH3iYQrydGPROVRdWLVJR3QpDbq5nLLvdri13f8AP4KwoyLqTs7CQ35PUmX+4G
UxQ9+SHNfKO5kU+XPqSiAyagxqH71ouoqyaWd3BbEyo4V9niNoCMJuz9JCEeaE/c
TJTOGiaAZ0ExDjn9IDUk+MeGcjWCRTc61tfmHC2OD7bkO6NuucXze/Y4cCvzHf/N
D+1Mt/bBK7xj1OoqEYIm5fjDyGkXA3SjzZ8EyiWyUvotGAns6TXuUQDPDSkbyngS
hhn4t9fcAEcklqq+xt8cP8fkw7ZEZjuduhtW1tMWgbmPw0h4/9vJBIUhtWpXRBxn
a/U2+evMIFUkycTHXo/bpk21CXJsNwBFKB4Junvo57rS+75kqjTYr9NcqM1CD1eh
t9L4JWaWpGOxntAxlCDoOXtspcbx5b0bEbImVXMUWRHS87F5q2F+aBd2QGgNTULH
Ol9xMWKNlkOykh6J3uzzI4GgCK0tJv46Z0t+OXF2vt2JpfbwHRUphjVS/dpQi3nQ
JFUy7oEeVD01/IP9jScBOEK2MkTMwjXZgUJgL2u/ICRzxvqEck8zcCWxRhnKGhNf
Okt7dgnEh/kLgi9usWgcSBTTSFzO9pqbn3j30wVsZBqsKTmJpcJXL7ffLO4eFb6+
TLlhG1Dioz47InmCWTn2Zfu/VlBNrG17olfZ+ZceTP8rSsxsXTjHThxtfi5+FgC0
snSneDAKcnG1w1OXARBqqkYiNWb2Dnh4dbWrYIhWkcIWl6T8xkg50xBdFDekxOMP
u/BNXC2G3tIVtiS5hmC0q/JM65m6oPfqNLhXEiTTOkFI8WohCU66YUZGoEm6VCDW
rgFXYoh2h4AcrLlx1ClJQm7owqNjWOfSw8PKl/sdy0LuK/6UsTLPSWo3dQ/+1I9Z
eeczmBZ5nolmghQLRVNLSCjU+fzqmRbsFdvSBOkTVMK+9DR/GPpJgzgJjwjrRzK/
pJDCNpsRi9fTeNxUYu5ETtcgBdWRBZ0seJnQHxdWW/RILeR3/Hb3gqR1NW8QjtHK
kS5/K/rjWL7GSEV2Fd+zXniVx1OnScpNV/5hdp8GzXCMRpYlbNhT8S/s3xxAv2+z
grI1nEJnaj8+Z4JR+dKwVqK9tPkNjPJDOzZlJ6PVZpFujBK2N6kVHMwrJb9ch78P
h/YMEGFj7jleE8JSOnychkpCGyQ1sId4/sF1TJkzPqW9KLkW2gaoJOeEQZMl1L+C
E/aweOdWLNZVITWFed08lJpuLR1cS6hDD3tF3nZkdMCwEFlcsGWpSrCRWrnRv1M7
3aghI2P+j9mHgC2Xd/TL1o15Kl0YS6Paw2xiRKJ2iy5CrMCYDDLNYfVnB8h2Hz1k
jCKJaGQxitEBH9dZ0szaLGGmxk8RD6oHRJicO/c7IqzpW/D0K5p88mUPvcXmjL0D
c8jhDXcWxS5n4WwHZJjJaUaYIm7RmqvYVw08Pw7FSFzzUwx9YZPg2WlcIDF8EYSl
rrdvDWamj5M0lUKAqXjCWXyRn4W5qQxrZeOaK5ug/ral19+s6Gc6Q+la9AiuEgCe
idhxhwxc25/17Gy07bv0EFNBKwDCK7UTusOyl9fJY9ACDowq+DqK0y2M9eFigICC
gz48wGKLhuVgGWUV9db08HQ9YLS0RbLSgny0j/SSUK9ANZNIwfLg/a8vDl9NmnO4
W9bQtcYwhKgtVCiAvy9hOqULeKrvv3ulAEwr/bEf7tv2xFDfOgRbvufeRsqcE65c
H7K8WNZYCFs+x7nz3/cY1L+kaGjlGHQviLr0sVi4y2eZSgtW3ii0pIP+Lu/bYJx7
rT43YUnB6ipAAu06BBHyrNYJiYMMfYjUmiQBnlRpVUXCm75iCumk18xeIpUxbwbA
/ynLoicIy6K8Pzz/EfQ01G5CPZjYVrcOcRO7IcRW7OVcLXtDtKgmNNNNZsS3Jl1H
zqh6A1bdRqxbnC08VC9M+j1xToEZv55c76k+O3EH3+djOMjT6En3Y0L5fEOu5V73
m+mVD9UL9TOABindB4IqDyg+WXnS6GyjMqW3UP9ojBn6tcXoWtQxf/XyqqkskQ8E
xKiZTO0A6Pm2d/BhnoX35lE614IQ7r3ObQjV9DQeROc8HSctTVMk67ql5x/+vMZy
MBT+BiRIQrtzFSu/1aBoZMqDyJFYdYF56RsQwu9VYzf8tIRxX2d5JPFBF+T74/jK
pdksIxybQu+uch3OsPQFyGCTSZBI1m/qBy3dUOwRt2bdB2OEqoS+Ak4DW4KzEsXt
/hIou2utYlVi2emyXTfsQpeqy1pvPwq4hCssf6V7Fic0RU5rjRfdxh/sEm7rTv77
JUOnP0sJOog/9VzeMnlNgqZxoxNg8FF4T4QUjS2GFuOHtSVtR2oRLqL/YnER08Tb
oTNFJAkgkwXa5T2tBrf6nQYgGfnffjNyUbnD4k5fNEJffOu5SOj2dm5/sVFCEd+g
aIjh2/evVJh0/3B2EawjwLZdIRE2jNZW4Qq+WrvZsfnWdJubHI0ra4oKNpuLYkYQ
LwEaK1i3KRRhNJ3+HoBjNwGM6f7QvAAtHNSBGe3IfWNEjQJx0tmQsssDsGP7gzi7
zN1Fg5+RksRrNzCxYQcLsLShqkDQu3VEwrYuxGoY+PwgfxsiwJAI2t66HWP934KK
7bqmUAT77RNmfSOAvyonucDcV6bV244l1BFJ03E/1aAXBHaGaT0Zoq4Ve8feyMHk
i+TOrko72SiwUfknln5k0WgBQ7xoHSYTn3gTBnYFZWQHQXRsFfhxqziZ5PPZtYUe
ZhgUF53ME0AF1Y4FeD+oiRx/0NIFB14movdJw1adH6qBV1AXOcp5gciXQoUXEpK1
R6XwgF3tvCoENC2LMo0yMcqhHo4T5TwsZ40BUR/07o5lO0G16LH+dPktfSwsP51M
u09D68vo47nrhNcpsJ+SP9N/uNVTgOd3xjkpVNwPtFlZgW+GGDQL4zTaDACcuYle
ZfIj1Od71+g909DA+Q/s1+K63s4zjzNfXtIWGy831aCD4Z6sXmH6fkGSAjuRJP6q
I5w7YFSfLaGFA2edAfkPoIW0sNhpiTehu//J5AwCKJtFGn28dU2vee9RY4ES8rDz
NpthQ4Bh5JXGyFJmsER3+J0HAR7ryTazB2vEtqiGVQMWlqcSuTTJJE2STKo9HyqG
Kv8pPJRpLPR+gWWMfBVs4PuS7Tx48e4M9IYIa5w8oEXXORbd5OlTFwCtmbGOW/G4
zQXqktwamgHji0t5GQLvKjYP1Gh3gSkzTrEvEDE1+jrnnQVpUOXBpbTXpRmx+YmN
93WyN7MxqdHWYLbX+3szSmn+anYbz90jLWQMHKWnXw6oYwYGsD3QPwxU9qem8xYv
LyXyuBNyctEwxE5nUxf32342PPpQYhlLepCx+F1KPS6Q9JNS1fT0sqiajv35HS6U
ojaGplSbK8dYlIn1KcRTJbpoHcU7iMfJyMw2V1KvwD+coG2IT0y4c1PVMTFqa4Dt
Rd2oOYapZAC/m8O/uv64svOBkVhfOf30wNFjqyCjay2cG1SxESquBM51kYss7Q7w
wgtTcyN4sfv3I7ukjF7LanwFtNl1qonTF4SliuvLKP9mG9+3xUHXh1RIP4e6pywG
PncrPKO3iD2fN+jNqWIlujp2ZjibYEHnNfyMyU2pClW3R4gZYITReHccttp/N4xm
CqjwskGsHupn14T00ECHS5QyOA/3YgCDaAlWf3JoKIWTU9LMCc1FoK1Mhm5wUyN0
+dEISB7dEaKbxWezgB67pbByBMPPZjnWSgh3Vc6aoawQmARWk7yNKJGyP4ackw7s
Elp2po3zHNSVRE3+m6+IOt2eI8tUu12Hibc1U3XJWKOIeFINpEQFlz6+EHqoWzxb
NqjkJ7IviMK+iFbuIUhJl6kHl1iSkj9mhmpKF22K8BybDM+TIUP9JZPC7+4PDVug
0sSjqDRm4rsdO/z95dPr7toBBLbYTETzF8/6wgTyN20g9uaxH8la99AqrrCpBGp2
hZVscKqcCKjE7lPZ9lWIwYqKE55QODKqILvWEFf4xcp9+KO1Dmloa2q//H9igi1w
+aGydUGlRJgX1NT5sfXz6/fVJ/PIEVT0q6O5hEypMNwLfjI9eUmcoN0uA2Z2zA3j
rv5B3GYlAHNDVA+XX1ZuEPLi8CXT1OH/2XlbB2qWYknOJuemPgIZKMUmfxVFrF1q
qpRms9pftGUgY3pUEC/c/n+wTCNZ+xhlGZxsRCmIn/Q2zbyLCE6QsMTQa3eJl1Rg
Mv5SSBrtiPWbi+7UvISvZksQC2GwFR05tVXSYs5GtZ1KbHxtQQvF3Ci0w7qFtFfI
CWRw7T4IJNrIvf7/gei3KKPI6nDSnEO8cz+GdvOazSTE63cAwUcAIokHTGl1Iqu/
up05G2b9tyUNvrxCGIuZktfTnTStSLdVIehvHwZ9Dzcs5/u8zXhslORyf0nEPktW
GUJUz+oueZa9vF4+ZajT6scPAqHFyI09HtuXvOXt3+940aibNb3SsBTM/zmiA+Or
GfJS1wOHJuo2OdbohJ7mCHCEDA6M1rUIdVzNHMtF+BfvoOs6FTQHpe7ns4MJRDeT
YRjrmiDf1KOsPsr4Q2K1XM9q0N5/OyHax2XjxsOmGiL5WOTdnuMOcPCcjw2tVPs7
57U2G/GOGeFl5rbc3HfAEt7M3pDa/51pETsTQRxQicTTDorX3XdX1KJoKad8kBd1
/PBPgHL4yJ1tx3QgQ0KGLexjiyMBAmMAENRG746oiCmVU4CeeKbGixmZqoju8iXe
hrnSJKUNaaszTCGHo8PrO3Xww9WEyFM1AibqzjqimxECnqm9lSrSlL2HDPlfwcym
en3eS9sv2vwm5QozlwoDhX30HnxyOEeTCeao25hxhDfQEY1BJc/5uS2UB6xX/zCP
qrKhbvN9xanqY7Yyidjmnm3+W07gnK60tW3mIg3XwcES6trKV9Gp4NYM6cfdlZuu
D1pkdJGRQgNfC/TYYzrhBsL22P5Og8mAPNmtY98vJ8RvIB4PTVxLTICBdak1Q3Y/
AMN0lWeaww0RX6em7cn1m/IyxvAPLcVkSbhj6fRtdMF3teoUaOs4f3aBIowYbT36
StHSU4On+2bVbNQ87EuBSiu64fgrRK7t4goVyrwUMqIpGf1RfTtX3Hakht2u5Vm5
sLYnKpTFoWzJImB1+LnNn14xfKu6tMa65fZc1teGoiC5pwd1AU9ttEt+5KIANAbU
SpGXswmN1Oc7dLYIKMQUh7G7DTR48RkdZs5vSqURQLXWNTCUATRdbDdRR9ejY/N4
v6yKOdM/NhiDBlZctwbFJvRn6XaemC2dO7LyDZ4/K+FhAlaLeU21E5Ky2Mapx0kw
FpUzWCVpQ2rt9Nzji+/TlXvFTdLpkt9ZW66FtJam0e0QawuumV6Bavt5m/7l1mOd
bLZ50EAECGs9n3XWJFZCm3YFoKFsJwdQoUIiV/g0GCnITUVNT8+luGQf6nalEhEi
kuyzkyhNgqpLMwC61slaPCJSwuiAugraWEJ2BE3Btjk8eiHWbCZ2xly2zcjcBVIp
gbm/zjFSICwzUXvgf2SqPAAqbFBnOZQNuj+Wuqn5XM+uSYusRHP+Jece75vr0Azp
0LC3C6ko0hsE3Th68AFTpvl0WKEwjuqBMxYNeIuTgD/dD2FpkWlIgUNJzxyNPGYz
w9zXYUwwxeRnkQup+KpYlevWPrYnp7+pgPKdnIb75fTfGSBUcTZ0oHurBwM3eIhn
UKOyO2T5PcReAGn8t0UpxMdYIg0VkH90+8nsJZQ0XtjQREhQsupn90+/fa+YF82h
Q9uSQ3ZMDGxxkPViorug0VS+CBBOG/nVo9ep1mKBYci/iIER7TN0VjONeL0j7sNv
CwTAERAaa4vBCgwqfjotOS0lXSzkp3zhFmStq10F9NV3896nWafurPRGEXmyd7nr
IHRJuH8wbyEY4r+CEwHWheDMV1mm49ZVWVE8tCbMC3dguHGkN92Li+KT5ahm3+2f
4XVvKbHDC5elvmynUFg26Fi3GejF8HJpdjsLpnHAmWV4bWtfIfxwi1G6F5j5yv4I
sXErZTr67FpJ1+2/AFAvCYhcY1bvdj2wn6St9BLt6N3UCU5Q5e1uTgtJwb06dt6+
X9AChH1YTudzCiZa3gmJEsOSkGc7U/nUuU0ogAnTzGlio2JGX1HkQOjQuzElih+Z
9KfSU2y5iK8yysGQYH15kLFckjRgALPqAbejQZ8udQtmMtKgMx70x4xq6vaOdHKK
y2mRMa7wqyH/xtc/dohXyuvZl4OUAclCQBo6VsI+JlYv8bY8sAlDA0SfJ78B7Mfp
fCzo+TsP4LNz6O4ryY1m6SbY5HhpbjdbgLt1IFcXm3yp+qiPc4LPIlgetDtDYqKY
sLMq734NrRVH9p5PqC/SvNeeJJrLzHkHiiLsfXb+hzfwxcIs2/n5dMjvBLGEgtpg
5KzgAk9Udjskf3DsYmnUybL4s7CHpyEZhnpz5sUl1onhZoLACtsK21/tIMqAcoNG
13kpuLhRlFPIet2kzrjG5NRBMZqPotcU9sdfw5/aLfKcwl4C9P9NbT+4iFSNQk9K
GDeMOTxltpRCcxfFFlzdZEh8HkHFt5l0moS5ghgxFMHdLYAkis2JuDkdkFig2HGQ
X1I/r2tHT80dnQK8t14Xx1LJ9jWnP7NJXx3P3wx/hSEPIjx/80sMDTtbxZJcU7tF
wL3KcRiDj+tnd2BF7PAAOfSgUeTLg/t8rkjkIkfK2VNAiglKNEKmJTJxgeyuHHwB
AVGGymqxzfpFpdUAo6DKi/naYdZMzEyrk0gGfNHUOpeOBDSIR+COpeEHP2iqi21q
N23J1UY58DdDM147oBw8WMrb5IWZqpKLYmgE2U/Zw9orYuHcdPynh1NJ52IA1X6L
kNU9Q3uNd82LfkQNdg2soRpDo+sifJ6aTorVJHiIR1lBrU33JG67nqv5H+pZjkGx
NDo0pQ3/0rvme3TG3EZGLTRwKidjRpTAwMqcf+v7etQv5Wo4x4Vw5tbVj+pXIVhg
G3/4CLWJLeGgkzdYHkmlugABLt5C8e84Sd68NQIoX6R7kEEBIiRA81exrLmc72bB
gtguqOhGuebtIBP68yxn/C7Ki2igBwi4tslmFSAhX6NmV6XrMeMpxS+OhW4ErSml
RbRI2YrK7HVompAtNxGdGOVhsN0TNlkTuHUWt4AI0fWcTlu3DHqodZRQqtNsOrho
Wa2fCCBfsbER9TehJnSnTVupHNfuMCP1aHMDLyikC2fqD516WMn6+Er2glcjrz00
7mZRk0Y4fFMdGYXi2kGUeLvHjSLXK7zaTIGPwDyzyGI7wvQ1xtus2Cif7+Q9Wv7L
WXTRbmKZTYKxOfaM/3KgRgXwtA61TGMtApkeCrcVbGH7Z48wIjOBkbcH1bBoEAFa
RQcL+dE7h1JAb+e4JzYq4hLpVXwT64QwbIjVs1O010p0SuBWp4N9RT53D0P09yjt
xLt+PC/Jo6FZRaNOcXiKhfw3vylDat2e/mnL5aLkC1Z0X5cEIrZ477M8kFw9wW9c
TQF0xg2e9CpfRy45Tl5hY6Gy9dnZ+5yWDCi0hIbj5JGcm/vhWS6x6JC5vikupqbL
ySsnjSw95tuUp6M8Z54BYimCA7o8Rnd4Y+hHzAXDzQN/Jq8qxlQMViEW7/oNPR5S
q7eKDNK56I8MGeedjCzTR4LUbw4/R7SN8cVyRldN7PXabG30Kt+m3FP1/4+Ecre3
Pe0Um+uivTblNIhSRmngsqMFnFsFJHgSh4DLO0+K7xVYnC7eR1DMO/8BXh96vahR
bLR5TnTufmERuI7g8E5FByaS7SgEEDexee1yIFTTuRwBt4iPkSsqCLEQqk9q997r
/T2KdsuTpzm0AdYn2Hcf2OJSKuD9+nH9o3FYXKlojvmyJ1jBeEJa6+Uvzl4mJ6rZ
Ou2udeGUEs5fUSSyhVIZT3DbmpMYnNrKPG+A7STD4CCCXrQ1nMbdFlCMVmMYhFeK
5OVrcqxsIxzb0kp06EaCToVy0yinIKyG5arjdM40IxK4dTlaEvJjUcHBYT/KLaKT
UTlh9r6ZafO9HOpa58g0NhkvIE6rufHfo0CKiWLssWykfzzJxs/TUcZio7iXdt0m
JIzLOL4iocmXcq883sqaFuHCiSwrrP6Qy3KoLCjO05lM1f3nRuMxuFIn2rTiwEfR
MWszCq6rzHSSEsFF39VRyrV+krF0EKTenb0e3duZyMeSyV2ma7kmtsGyDQYPRiO9
yTPI/liloagZEjexNyl1h0w5VOmP8WcIBeawxQNV7FZMo0Kf2AMhgumnmmPRnM/i
bqrJXZCsxieq1MEMpnv1mvZ5NmBMYFdb3ozlxhfx0WV9pjkdXSv8Y45nZgcfiZCU
yLB9w7Zq0WBaOyrEzUBWdgqOK+WI2h2IvxnywT3aZ3tAZFpiWaR3E2FJfZc9yYM2
cqOKdtqbHkcHeGAjv3oFhjLZyHfPGblw3DDcUTpqOOQPt9uRjNfeb3CGj6y/8AIL
KWFiqt5TEmzyM72RuyIASwkTt8+L9ompOx6/OlzJsapR6DgerxzOR8GFs8o5IEBs
+dr/1PBBf1/BmO6MKTMzuATVyRX677R4yzJ0s7jcGfCDU4W9bzxOfTafrZxPfkZN
1drfG6dvV34Ohvw+BXsyHB01ZXmAjVpoqhozGasZcLHyPodqV9T5iDkMrFuz5wYn
wtFAqEGcqwKtKxzrNHKxFfNjdXx+nITFJ9p+uuqDlNF6JnQPosRtqnhkKRAVwgMj
kQkQV3lR6/iouCgCD8tykjw3Dq44vTa+aWmaXTV/Tjq9HVrLUvBBeWxBfOwe9u0c
RzzXavWRHupqumISBISMqehu53gc/WJ7EwTf65C405Q128xa0VzFgwbK92rh7mj+
liZNk2AnMAF5zKiI4NHlhtlCGfqJaBYVuZ8sVdOMgubc0V2PMiOEg3kJ60R/f0/4
b7aZdyhtEieMx2XCZdavec0beBobVmU113vLGObPpkCqUdcqd8jndr0hGlXQ5O1a
sz8XQx5F66dOknOLjMQU1TRs/XxXrtQNrPsmj2ycD8tOEpzUIbgHQm/h/PX0Act/
0rpsINc7TAqoY5F5YrjpM9+UhvZgJf8N51DnOfxnaL2BAxO74i8MMn26AfbSd2+Q
TkeSFe0HzFMsaV5TYqwOK2/3V4cxZI0iU9/lHa7kjN/ucv9k2NyvZQ0wUjp4e9Kz
oAqW0/BekrfOvCQ9UZM/CSSRe0JiEzknnPFF7l478UogQqLgywrjRdhhtG3zNcU5
GDpca1JI6ZIJcx7VXhVnX80DrxHDzjHWNtvRn2Zl4dcUcAT4P6ZC6GCY7gSsXfGp
TxpZk585oDa9wbiYTnsBnd2GJ0qVGZgPOzqK4zqYI2VzGeT6s8NfUBLXex0sSq9I
lcTSTeWp6hQ1TT3a/9Rs7nB+SuDYuVE8CmYuU4v/ToaRzGlg9Yf5sbIYauSpQyn/
Tbu0KJtlzE8Ay+q9Ocj+0UYiA7kUyvlaJ0FZ5nRioBypG9BD+MKx9wHWqN5gXv3W
DjSMvs4Zw+Bygy3MNanbrglbT5W50hEOgBrHvgahRH/PJ8dm4uZdJ1WSyj6/xxNd
U6ypLoDlBKUfMmHBqmXKatY9GKtVqwJUNULmYAve5TR4FMt4gwuR2CRHGgiq1JcR
iFvzFJSGDnCRU6WTaUPCDSLy7EyxRLZ4wz0EeGbTlBWZrO9Qd/RjIMyiowSp2PtR
tgMNRmOapPBD5eqQ7HbZ1JlZPtcEZwFRNgynHrLDV16ixSFu9E5vahAZeORLM/jf
dAS6wthoX6yHyAOGPzz7IcWAPk/7zzXA0E28S8yAnYDQfyPuvOHUtTmsMr6K3anL
m1BnUWEqB6UNl83bND/ws5BZOb7clIbyEvDmtL1htmwnxGMs3yLY9SixYfT6Evir
mM408i+o2XL+ZC/HdHGaYmQmkNbpClgT+2omo95hs/llyRh29KF71WaKUPKrngpc
sqkxiBznB8xSS+vu1nSq8G8CDn+YT9FWvjmiw6K30Y/6evW9/MmG4O4PV0Ra83fQ
ZHSApp5iwuGgjC2A4h6wfPeBt81HT4/AG/I441WSL1lyL0Qckw6Xg3dIorg5cOJi
9RLO9LZ55rrBNV0A0cVphL3uS15yi3eb4LrZFsQGxiyMwiojUXICRPzmf5W5J5o2
sIloqgNmjHiBdEDRi8Rba8AKFOXGDiixIfxXY0wWQVdPl+XhwYjLHcuuEW9FZTzb
dTSEbH5rFrlCdfGHBgCVXOwesXWy2ZBaHCRxMoQQZH9/n3IiB90Eb1/1Xl+FwXIX
ICXHQGgYBviMDD1n+Xlc/KfSI0MV+JsFkqxqCXAYniwIJA978TzlT/SvC6gmrYlS
WdBCKMeTbrtx/jjfgr02qR42uAZ+XdwC4RIWtTcXpjn0MpzeBQKpCdsS+Sanxw9N
YN0SCAxTmMxU9ms4LEHIfw1G1Sd8/kYCq6Pg6ZOy36D+KBeIH/9PfODuwL87B6OH
qHVfc1KmxUWeQevd0b9HJefw9RlzzrduxhspOhtJ5TQtrsvMO7CIc3SbdHnqrLGJ
X9TvMbPEW4gnEPhFFGgztAoU67x3z0UwwKlhAlscR8ZPpgKWspdCzjnzw+lQV0Q6
WLKV94plhBmuoQ+YQ2sWlNo+/NWpduuNzzN4MduyjJyb8nMUIUplz+RG9SZlFj/r
n3QQ+16Kp8uAGKPwHpuYHl3Vqq6tE+mP6CPeCFsEhFqrtQzrPnpD2Ku3qYXBvqhM
jZvft1LFbs6v9u+4EvzA188X/GkzX9v/Eh+ixJNXtEwPjxyDCKDzPVxZvOc7WZNn
XJNryjetXrghCJ2Y4t50DO5Alu9RW8mt0NyCcrmjdONgeEdfeNIkWzHCejfQIVDa
vn0PpolQEnqx7HgH+bpRpTIgMqY6+pWSU6eXMe6PzX2obEmGR+HzNe3gLlcV3GKQ
GxEWtf9W1JSg/b6q0XMikJ12UJQh/wW9O0CYDWOd8ufZI8ywuiY/DlcYXHoj+Jar
FVfxB7T3as/zFyNz49oIXQPVZk4lkkvo3XaCEX/btXNjMuPipkFF6EudBYrTjPU6
M2trvUd5k9Z+FSK9zKFE6j72ajhgBylQYi/zPq9SS7r4w76IS1gbQbay3OJflKAQ
lQ/QQu+rYsfSmka/LaLtqP1lWiTouelLu0Kc+9UivrRbBzZccWNdC0nE44MttmA1
T0cDzTvlvvoamBXnjcVReHpVYQX5bBIKfD2cQ8tCWUNqYeTmk/uolhVyYW9eHY5e
g+cB1AF5JVELgiZNZ0JD2dDdiUYZPeq1QODKkxKKpGBiZw0duKi2SyyC/aZrGa/8
xy/GYAckjcJvP5bLzcNd4nDgw2SK3nUmDsQlqa/V0KHc7hePWLCdusEiCGpYOgpn
1AQq+5CIecgwfI3pl5VSydHS6etsMhgkO3dNsNGy1B5w2RqtZ/qNkkET4d17gw0q
XKxsbWhXWLYFwh1TSV0VXyZ0kOJA8J/xTDOvYSn7FoJKB2BK4iV0agqwViw5m4MA
6pLJAH3fz5Io/PUMOdf1RIPIrw4+rcSQXR0XJjuW2BEo0+KlNHSUwefhY9S2yfQL
gsx1JJudZgMnn8/TrMN6OQnyyzduVZAYZrtK9RI9MshCBBz2JvFcKdAMHum7+9ik
50DsXpu1YIlHl65xDaJW8xJWbPMtNIIm6WZEX6Bni94HBEPE41B3Z89zBURzGNvL
R9xwmi/nexhye4juL4xUn1pIefuhlftbn1eFJIumudAtc+DuLTy5X9hlESyXMXnX
2YHrzIxpT46zSb4UlLpHFDxsXYcZNJFCRNo/RecLcdz7NeZw5VOkVSQJjmCv4Xn5
+gp6Up+oddSzCdwYr7BqKAcDSHdzb+NLO8WbD+WyGLhOgV0TH8BtAtHhcXRvWHIP
xIs1ftAx4+fpN3ONwZSb/PFQem7c4cHtm6Xt3u44X8z8mglHcRI/K9UfsRuGko5o
CEfvgkV5YOq9dDv2do/Gm8gw5lvFp9AyZodmuOnGK6F7gQ6df74bJRQ39VFtRUAs
ohidigJSCR3+JUIknj+zUcMnrvt4hbwio677D4TyuHpcDx+WS0wjYOxveB72zBDP
GCN6KatK5Kuyq8JNnUaODxqmG1P//L71LQsM6d8qWYR1HFD+GJpeCR6XD4c+Xb1t
azXWLp7QKGIxWvsRDHlcQnVN87uc3JTHJqOKgE9jvu1WvAoz0vzXGSyH9Lksa1/0
FJKBNkFiRHqBYw6EuBJ5VJ/h7aD1Vt+MnBXGxhtsxDCEGzcVhMakULQgVKznpkd9
CEE6T5Da2ZLE82bh2Xm2OhV6v8lHgG+BK7k2X+OAZds2NI4Ywq+eWMdHilcT3fpp
b+lM4AaNLqDSkThLGWPvLKndmFiMqVeweUvLqSfXz0vEAmI9mDiBX+rvdtA9qNMx
/lY6VeAwcseZtZcPuj8jnabIsQPnrY1o2yKum9HeFfBb3V4ah0hlqXQ6EZrZHYio
E4tT4Lr+e6UP7/tcv6LZ1oZdFfvL8PHyQcMxX+u2B7g3m9QwLu+JfQREN5NihYE0
ODMrg/OAFGKk8V3MIW+1lqFR7VUkM2AZrOVS4HZVeld/j4lKGEEjyscimCTr/uyC
lgt65fyMHIc9127dHRx6zdsjayo1HrFsT0IvJmzYVgeX2URH7eKzVlullxJXBb9h
KqfBudMDjeDgIRKse03loqaKl9PjGgK3NW+8NEtRdFsRD7nWz7CF+SX0u1q+rwub
bGazT90AWsORV4Cxi27aNw3QuIJbhN+Hjq/qlOD62ZOm1yuUBC1be3mQzMCXJOQp
ESXf9NV0KcTdbt0HFNvWJo2hxSIToYLTzEU4FllS5Vdw70ehaR8SsAwFJckuWoYP
jCoOEMRSUIsCiJ3j+UJYkKWYBHLD/341Ozj7aL1oU3llSFJeA9P8Bl4kwD4DaSnf
PysZvpyyb3M45eGq9zVM/WJKRUevVqv3LkmPRn0MkbctKhXNwVtc+z8gUjckdAt8
pvYW3+MILeKolFkqbjgdV/IVwzOy6d0AvZv0BbropiggGmFq2fgzH96TUJgAWa2q
LybNfeGzpdhR+gt87gP3yAJpa2Aegqy48pzb2qjDt+rO6mcz059V5IvURGmjK0Ul
QrLzwx79yczapqPbcjYGShFYke5/wGFd7cPeeK+AE+R1Ewe8E/sLuLc5Ze44qGcX
QCxfnj6DHOnIvIaeoQML9Gt9fsqJGaNIs7VANFhJYmOmD2uRjpaFOHaAzQ+JezoV
aowL3M+lbq6r0007Tl4Ue/GgsVpux4hLkBfAHNU8QswNGoYOVvAQDIptxOOobDRf
lLOcEbpYdlvDlnwEDJZ+p4WafiwFk96i1UFpjV/2ZvpkRiaJ1oN2l7f5p1FLvmD2
Eq8AAdg6uwrQ4YPjFslqO7b3z8HeG+/opHlUxuAI2uKNeHKffXf3Ji2l036AnJy0
u7sEJdOkC9EHUsvd5tKxcKAyc5IQU1kS7YQwku9p7ohfCIbfdylfT1ZBFB1PGvWa
KC4AhAFW0Srmp8ZVVMbLOZjVrHaB8EH3eGqgiiSP+zxtojaVrfyw1O2KXsG895iS
1NGm7pNWokmA1wtdvqAoXhW1yskarAEryrIvMxLojFNiRI4nM4khAam5SdF/Sylz
J0r//kCHWepASFDlsTbEd8dZFpF16SSui8L7uT/jMj7eLmEfsE8XE35a45Gs7WSN
pzdT4N/3YMIMX7YF0PNG47yMzJlGyzsmEqdQQzq+6lWbBcK3Qa4JYdXOpYPSSp5W
D6h4odCAX4mr0K3VFE5DraBgmPzN+/RsPSZ+EBeOf8AKVBvhkxDz3AWhFd55mdXQ
iwPnwv+zK4mzK6+KJy+GnjSYZi73I2k+UJbTLEVkxW4ihKxcHfwUCylm6wghqCib
4s4Ax9N+DS7a1Uxt4ytTnagaaaVdh70M80l50g2WbEkOvti1qnUTyY5V5e0CccRw
8Zyj0xiZ+6/WL9W8DeCYYumGcodsS4n16l5V38ywZxP3Acgmj7zDCa4qzzFXOCWN
NVSuOsHJcHAcb5KX0hMHeZ4+UZC4AlKkfIiHAw9i8QJoC2EBkwXVkf3v20Ua+Bg8
dsXM2+KWSZcjkBVLTzoyIVTXOLDR783dDo51Jq8stLMNbXV1UDSgYmDslcr2/J6+
yzRstQwne+cKYQrSk/cicC0r/+bpWUti1iOHWlIejjqGdQ+zuyMPF7F5Gdyvwq1k
Bd8V4zaQf7HypLPJN9pMLdYHpmzH++FHf6bQW8niD2mJk538hMIEgsoQUXgAvh/Q
Djv6LHku5qQNBCn4DB4/gMOoac6wpPKr1IYzEL/NSKjdWEXSF4MFNen6njCTOiRP
0ZFT8oLkdcoappUA9Yzr2aZI/NXVzOwgIBP66U9sB1AMKSLy+JtBiokZuMZ0xT/Z
jqTutUvj4YFnaaeT9z74ZgYT0apGTeyWIu2pX6gKlkqIfrZDFKpfCiNMoTs4H8M5
OdazpDX/M0cnfZ0ZCGGk2LFsVe3chUCMSOIhWIlkS7s6X5w3DUtOLxvf7k0gwhuX
DN6uzj3TNsxQt0ChOyRkXTCkYEGWpiSZpuKRWS61ZXIRHnbfO+fF8CDIDuQopumC
+QjWxejZ7j2aJRHpVssq87EQ6Jd7vN7xu0Z9xeoIQqyjjV/BFt/AMPjXl4h1hKSm
lWouWb95a/te0VMIOJ5381kj2+vg8Zo5Uce1+gKTfLE3vzBNnkcUkDK5as4WY/SN
4qYiovcqj9OWrgrI8Xkw8SVwMHelUUT8m+Yuh6yduGw8xEEAcFePYFj23rWEm0Nc
9aS7hLgJZErAkXxzpcPvDCQAuPlAShwYwvTZsy2SwA7lwEyk4UnoaRVa/VcCkJOS
luAY0iKAfEXqxTTiTUDz/GAepeZ+jU5DPy10DNj/vxwhdC8VNLD3oCDdaheKFKGO
Xx58xRfErDqYFRn5nP98aJJdDFlcf4HnZGiwFZ4Pv7WYMGaWeDxtntvMgPDrho4M
dHpWth33ytk5CE8+bFlA9fBYsSN8whTmm0/0/k7ttm8e3QXEuiCDm4gYXjV2EIcE
JSr3Q8q4cXSGJHAPHIzl7iujJ0/5+mI1Fy6XGFvv+Mzm4rlHFRJkVQKPppqny5A9
NPUY4CHpQV9aj/2mCSJ8T2cE0CMp+MiB6pzg1Zwf3v+swTcgxiMIIIAx/gB6LnJ3
IOOc2unJdcrtKxI8NxnQ66jbmOQhZtGO0uQz20/0736hPhMOLaILBNAsp/lpXgUM
Gmf87VNCDkCDf51X/UdcySLcN2uw+0gkdmiUE9D50qHaOALT/IT5MKEcpygJcpQr
dBKmQsNoYqfVZF1sQnH3H7xFNYL6XynEDunSDCoG9m4OgVbhpHtvm5Q3f2pxyU58
byinH/6ylvrHXtjbR/Cu+34nSv1XkzuN3odU7WDKXVRMiL/1I3B4LOufCVnRS7Rt
axPthVBxAjqEDmasraq8FK5dqlIPfpp3MivOAR5O4YY2u1KJiTlGgAd8sUmFgUjf
fUlmeftBGhwfdYNqmjRq17QiJqeHFquY6lh+rZae1fNE44ShF04MkoYU3VnNiEgT
9/qIgiMug5Bo3EZVhKvLWadcYJMxMLjHsC4wf5hXXh5oFomPiENt0ELmtOqIi6LV
mHYUn6mJYJTygHi4DtB1YyTHT1WRSy0RevfeIy0rGV2p3j08KZSfaeYIqBKhLWFO
KunC0z9GlGSCSqYCLSc6dArVEgY8KjfTXeKFtm0coTlHeZnv4eNiqzmH6uhqhgA3
YSFW55ZDHNHluNpkjAjT96oJ8RvHCvTz2BNXpNu8CxAunknU9g0L3AghvqEDx6ad
Y1o1mahsXNZZ1a0TfYATP6zWcmN6897xMiMFELSFkv/cWs7CWjhbRBfcT13D+GDz
gGhilinmzTI5dASTCFBTOIBb5VeNAVwpDp+3pZDCjSyMemKJZ26Ir84O2FK5j8ts
78MLPjzpVs8dioEz5sI+FO8dyASa1+OdpbjGE/xZ379xw/tU8XX/PKRxA8n6753d
qDoBSILMHxl7WiAUPpya84loUMONAA55oQR7jIyPuqA1oTS6pAWdRsi52Zv4wLXS
EQT3DlFSsDW/J24n/IRvgcrOhBb1xwY3kW2k+8L9q3A5Qyt/G1dBKFUY9tT5FGUj
Sdhd081F1qenMwAGyhiFsu8EeAtrOosfRn+8kXISMu/+eRXcFPDmQ+4Y/AjLtYAq
weE9bZ8OfbAnk1yh+5LKDlcFBGoqhUH4A8pgrB5nEw/aWCHB/wX792qDjRZ83AMz
VIilJHLxIGZkA7zS53MwYO3Vr4teMvkbYcNhpKoLWniGd6R7MibvwSF0zqwu9oA7
w1w3hYc+lVQsxkYD6hB/SruRXojQ9pCiLMcbuvUhfQKENhPPyDAgYWWGHC8nebiG
sQNlU4uGTc74S5hCwLDAEZq05DUIAD4qqWrLeXq3gutyQhQtyR2aqYDLrengF2hd
TUU8mSh4GMS8Xhb7ZO+u0gjuzySBwpfP8fPQ4n2ik7Ws51ZbFIu+uEMkpRaR4hSZ
VTTjxAJ9X9Ec8pOtag/qKdZioPxIaaKzNBh1E89WjRqMhCUVkvCVe6XuR/8r7zk2
eBk/nLVtcV2U3NWr8N3A/Kizy9yfMTwclOc9CTTvP6JsD5hVXhtkxvO2LO/fa/vW
YmdQ3Y2vkhu4hy4gE5TMqhnL6CJMLm52KhIUSytl1FBQAFfyxaiaHZo/yV1yJpf9
bfy8LOWkN9ymv4qBUEHOR3QRdx0tuV1WeW/9OClsi0rlo/e1C04Io2+ubmAvGB62
+0PDPJenTC0O277jeJELSDZvoaWfugJrFo3d+mc3nMA36ILkYq25e4bVhzwY4hae
nVnhzg7EPEEufqbuR8vC8YQidNzVUP6tO5NJKaQ149fPNQxqvshaoGenuRK1WOqO
PmqNT0AWw86piJuAi7DAiyptGV6GxtCL5YWBfK+Wo9PePrzqYaoUQptJYByeG/wt
zv9KFksLiAfzyr3fiZRbYtIIn7k8zh9EGaR+BMfXroQMvtPwysX/vuHUMJFWXVFQ
+iFVl8kgmpsLVVGfTxoXoS/jmY7Kby2DmTffFGJbStyum/lRL9gr3FS9fMRaBG/E
NJ5SRRMy9yV9IpQ0jaeR/0FZTvOezxc3RRBEkeViLEkCfabinEQhXGpEDKfKbyQz
blT9zjOVbnCcj4KfZfYBa6mxTnpyTgD4qObUluHdhnlT9kCb8vCWF8jLgppzD3Ac
VzTrMcZgPOTR4YuR68NNbJFTuv/GTo7QpBvr2GsNn/kHN517te0XACcgHcp2lxow
GKhCrkyavUz8cNn+LGA52n+Ai7XN7G7PfoZZsl2RGbTN8+SiqTiDhdS4nbHOCkQv
S8da07sb3JHnk/lViTKEOk5TVkHPIQKqleiHzYOssEVBFkDBAmz3UxZAcUMLFAQM
XA6/TMGCeqbxg48+cJq8XPbIB9BnSYhdGID1hVsUMko4Gezc+fOyMN1gyn6m33sv
aLvSv12sv3HT0P7tN2F0qiComSDtvYdnzVx5qS2N8xP1Njj72NS1yYeCNXy3MB4Q
6NrUg1JJqklE0PGnAC/QOc8wfeMBFm44oMxHMNP33EC4ij8suRCOVPM0qiyJtT3u
74lbL6ALHDGldObY9mqN6WavTH7kgMV71CUtaf1bAX3Ogo90qu0fwU0rFrpbz18I
VrI86a3T6IeKxzw12Y8Q5Ab4Wa57dm0YHEhVE+ENzG0TyA6a+6N0V+INn1gD9r49
gZaoOZ2f+RR4QHTsShX2bVMbZyNpGFuQNL14w09By1oV0AE72KVVGD6kz3r8f9GQ
RYqpU9Na3IDmWffOH1GvwY6jggy37RiWRv6vw+PbI1Wo/L4VROS94CYlIdPHzV/2
7+8+lFT8eIHA1kL35hZmwbdYaDDsaRC3sQNVoE0iLaZqsDoRGt5sEPqe0oEVrZxJ
5JNgvvont0hqUAG3SwuV6zUnuciIrEAvnGI/ABA1Y16wOg1tfDQMxYe10cmRZ7V4
HOQZi9a4z+p/zU6NjUl9gs4RopTOd6TsYFSvQap+TjDctX1JgrpvEbtf1dTenT4R
/ZPq8d4iqXxPIPeDGTsSX/SycBJJWIvA476ZdY2cUpMcEACJHXKwW7WS3u8JW5gG
Vn2mTu+5GXEMrp8rbQSiz2dhl0AMxPq1dlqsTGufYsT5wNpnvp701KDomiPLIl4I
r2oUAN/mBCEdUb2FE3bAjJDE12kaOpkaZbMG5zEeWnqDeVqeiDRph1xRhARfuQG3
mCcNsN0iKWvWQVREt6G7+KbgySZNj14nhN7Bv7L8atroJ5R0mZJeKtuko7pw2P/p
4n33vTAIda237ZC8N9gQiwjedxza9kKMMYLID88wlsZozdBqhvNEUwD7B0er0vws
5gBHHEdY9BETLOmdbt9g/wFkq5cfuHRMMpQs+CZNxenhRjTG5xmp/0GvsAMDI1zV
tv0RiDyffaKxPP/f9ySdcK3922zUqA4lTv1emb0XQ15UcBYWPnhCTx69NJW0yMGJ
k1XBxYjvBvn/H1x4OdBjoNSr/It5DRocuu9tYCo6rqZWammzNYM/9kdRrK0mlh/m
+y/DldKhfAK78tnG6y00dOglGZg4ZO2QVN5HvfivxCqkCaT8oefLOEqkWkWIrsEu
Xvor3xLpkD0l4b6YlE9H1MZCEsgW9G8JW43lkrWSeafB+hwtaddNW0kiPqUxYEqi
c7tlrPYj3ipivWQi4Bues4buYoCoI3xwQgnVsLzKhPNs06utFFK7u/NWFY8KYYdI
n3A7z7ZHIGQRHddzYnVRqAX61+pkHClyNC/2QlDSX+0UVFiQf75mxbDVVp58L+a2
WGhUXI3G185ELNMONpkMApeyi21vspU+UcMi1Xf7iYTrf6cClieJKByLLdgM6aFT
E6iiGy7bgomGu3TTgqr/0tCjhdsZMZks7cIDVD9FeHOpVWb5MsQWsgt4jzSI0IOP
xeukHxMDWew2JYzlOtbrDQmGmYlH/YtM1BppG+iIGJZ+DJOSqDLS/9qIvK7jjvsd
+YvodHx3nAKKWi2MWdcfuNBH22toCRRrR4AXYoDUHlzMes3xhqRzYh/IvZwb62RF
cK9LqsUokKaBDQE/zqlvvKwsaIa71aLp02zWBM/PY31b5VMf3acYrPA1tAVpHdCE
5wwweRUB0sTyhuvDt2KqX63BgOWL3BX5f+Bk+4n+UyUvm7SrMo5/DtugKEEM5F15
FRKXrtMLQe94yRFXMzc+zgQOhTRwrPXxH3QTJAkl0TC0y4+O+A64zV8XrFBjFenL
cpuwdrmjuhdQ+XKHpqJ6IYnZpOgwZcWdcyatfQaB2aR193/t73DN1mKkpXrJgHhj
SoB6E+c4pRWXr+RX5h+IqybiXt2ebq7Za1hDqPqkRwrvcF68sjVVb1h750uRMTa6
vPqmTKIFKGsEoPhvR0aPHGG68Aia/WsLto7+H/bvHzpIvKt+N7SpviPa4T1mdorm
GbwhAXbnoMMJHxk6fJ2QOjdN8zWuwQ1mexEk3h5RChSJdChMjHKAZoxtIEWf2Ec8
TvAj7OJfDofyO7u0qrc5OdmWI0YLE3Iq+YmnXdfNhooUiqeerC+vHhESIRyJlv6s
g8C4JdOUXcSwrcKjswKnkgmKCFyla+y3rF/pKbjrhzudRkl4UbypbiR93Nqiev3n
8xH7DjA71NqI1q1G/DGMOTfxOcl4tAktxQoqILxAjoMDK1RzsbttdjmYge2zB8aw
ASSdivMvsZjdPeMurU4D8RnYw8i5Cm/C+yrhMm8cpoI3TrWWA9oHTlI9+weCdY5Z
3LWt6ERHE3q2edlibnrlpWVSjf3JtSkGyxAB6hPE0QTjjKwdzS/qiCKHk8D/Bt1M
+q/A86sSEk7isFfJW19QxoZZYVQDrZVB1cHgQ1q4Kx8R83ZvLNS8rs/gtwinbAzu
GzEaAWju86f2PIG7rkuJf1Fofp2a3MlJspORmOU29nENr/GSxja+MsU6fhwOeJCV
EK/5kmFCdASCtXWPjSBOCD8Lr/Kylm6OF6GCbwmH40XbdQgOD4UUel2wiyOFmZcV
RuotLLpG/ccWroQ7uXXLhZ4YS6rEBiWwhrJ1e8oX04y6sZqBZTONAVjS/s+Ld0n1
eNxEVrM16cRhceNMeZhzxTM4MgxqTSXb/vT3zm1IfiajIYmMniSnwm/KQzaBMz9X
KhVKYRNHxX72HI3ge+mKWSQvL/yjS0OW3GyCiCvN0We7a5X7f/g5CDLoIAUpac6t
aUUOS6qbrPY6u6XQ1kLQe6ygXwzowjdRrv2LH0MafVcH7RXlHgoZGEGDuD+zv1nz
IC0SF+X9Xufc359lmK/395wXRPhjcWZbYYTrdzumLci9/di0vsbXpOmZnbPNT5Ro
nG2wh15qAxAjcFYm0wHG9x2oiVDsJ880a92ITU2pw3s4wJlrq+/iw4rHubsIJwe5
0r4rU+lom1vgYAtPqgfxCvQQhl0EWfwL/6a3qFenH5My+2KDDdM7HpY/ZwHlKAjB
GAQGr45TEu0FLBjxmxAPyvTJXHZJGjDkB9Py06f8n4ThP8oFsOSynsmjdQW4Edkw
9NEd32wmMcuAwKoHcgsmUvX54PgCTCuYC7RsmpXNtGfsPNjpBvMkDcyJJGHAz15q
p2LLPMQssLmVE65hBZf/2jU8U52czqg5VfjummpMJVlA+2TXudGmXTFsZPoWVoy/
dTOdgawtMjAYLrwCt8Wr4aGhS85wVM4bM4U5Qqh3XtOBArIVuWp3RzomeRN6nTCL
U4Ccn2EwUGWCMM2BsPH3alWUEGJnVi/RmTbW8yfuJer/iSQ92DuhfPoRYIkvJNEc
hfqd3VHLN5GY1Fc4QLy2NQCO9aZJXck0F4MHzaJDQZoOtqWhHz9OKffVbWeMDHuq
YC+ts8NbF2xiDB/HvjX9bkTvUEXbObxuBlWUUAglTLKAqIzj5Sp52du2RNGkrl3N
P/rdeERq1zhPHR8YR5vQCPxfo8TD4T1w4gdOkcw8wrcsdjMpMJHZhZjkyafzxjGk
PB5MIwrA1mS6N6O7jmpw9JF7XsnkrS3kyrdGdc3mqtJcG+YPw8vKw8WsDJDj7JE6
CWBDHfJxKnw1yRR0B9xPcbPK9jTIdqMCzA3lW6RtGk3Zl4k7qlLXPV6yuD0K9rcK
y1oE+OJn8jep8fSfhs0Mj1n0D2+KsnuUPoOkrAqPjwqYPd+xVeLjwlbypscA8iT9
2v6SF25bUfOf8NCMduzR442xviTJX1ITqyPEl87Ev00984jYLL7vt9sIRwl/ugkV
RftE0Mejkjayx/lak7xt8IeuQc+F6W6ekpMi2HtZP2iryRCx5PP9AT+toYa8N4ye
EpfUnH69n9ZPerYpuhXHkxzTD2I0439xwpKH3eEPSSjQ74ztErA5i+EhrVgeCko6
XHC/y5JPggq3xNCVBtqiEtpfkYMaygrEjNCldo49xEgx8vx/Zmrv1qDQ7np8TTya
owh3ljYhtZ4FbesEH7FQXagr0Bdqi7tphoIlWs814PN8M4PhUsJIC7P8QXhqAhgf
qmSubmV6Ej0pP5lqT52+aHDy3GxBJBeDIoZxBtL8l231/2TsFWcofhiyvNIJy6yP
zHH2ESZNJzmUUzI8df2cDIM06mNf8TBXv6aDU3En+qColpjaxy40CpF5NytWTNFB
U3Z99lKp08wg++EcX0n88p7Asj5PTUVkC3igRzh4xPlum1mLh7HUnQQDV5fcrcpV
JkN73yYbobmG60pqYexCIP/U6FCyXSaN/zCGNbpQyKtu/WxT959iiSsQMSK9mStC
9YKPn4m/6C8lH/9JuWiLLkZtovBaIszBF7Mej5ajBon2b5dFFRbMxForo04nXZRH
CvuRHjx66jhVXkgrTQhRCywvO4sWmkLesb4SJTvbEK4U6fAZDcOp+eKliTGXZ6rl
c4dCAAeKKJze6aOnJWNhGw8ZH6TRGrzdjVgCSfY3mZl8sKeBQ+Po0LXOHDSsknO6
X8zKqhloTB4gWqf91K6iDk2urKwKCYPVpj5Ab+DjUMf/TmA8rzrIj4XC/EEXs1K8
HpdK/kgivrXFhbDa0dHeVbKg/lRxmyNg23kG4YV3Ke3jEitWdJbGXeiyhnUHdZRQ
HcykxCqRogKQm9JfFGvIGsDxeQn3QEOv/kXQhx0ovN13n4A+ViUqbvHpUde8PGv9
qBlWRhvBal890nacJNkSnnv7uQcjxbDn1kv6BX+88LdF4cVZZyb2XqkMJ+rQPpuK
6kfMgqsKt8Q0DhtlSsJT7I7z2RwGne+Rcj9FGo3lgK97D/kyTu7MUWqsD3rtQ5I7
xPZIhgF+JqgJnVIzoEJ1piVzm5XF9JB/DQYISC3IraahsVSB9qfDWDJ3LSySpHxr
8tGjcvhCLhWSKw+ZzavAWxyTZlPiNDzBMFErkuWWNlLkZ79l3qqePvt04OzpZHj4
PhJ9rmZnjeqngPjUZ+cvFfjkuj4QUswwOVqpAgvhAybfHUcpU+RUWH/jsrYsO1f9
jqr05xvHK6HJP93cfmoKdlnUVJLMffCDFNBO5q6a+pszDoF2jcLgETlLc16mJLcH
glxpNZrPXWUkkO08fN9KzoEbiip88P27OuvBwAiKLb7SrgsAnpKSjponTbT3QnDe
JPn4+yZAP2JiDUqXAUbDk9VKrbZ/CFVr6cWthjZgKSZ6l1fwy8JqVmsKXaAbw+iD
/X8ndfnZZ7o5mJnC0qz0EdIVDMgf/YbaksOhCYc1mt9JtMEcU/HR/YPxOtYAYKBt
VioYJt9RkTTCHxTUYtwulp1htvTVxg4gbJXoT+ccMfbAuAIekjwvW3JPpVbMXReh
+RcnlGKKWA4r0JHT2BDcRSpeyxdq/f9QMVVDpr5sYbLfHIufxW511smb/dPnJKm0
mQoGcOGtxikq6FDvEOzs5rLBNTeYOHP5Ug+cdyDuwHRqx0IwdIRJsP1zw4lTiFOE
nuJmGEznGQt6ch6ZwfCnTx37G7B6LEKhVXo/wA0p8zFt1Yhu+6IXRToNkDJtT4Od
rT8B8fecaUcLoDaXi6H7G34qTrIRapEG1vFSXI+a1hvHh9GkagQqhUPFCLvszlOF
tj076A9xBFYoh/5anZJ3focFzFbvOBV4OmJ451OwdfWnZ7ur1Vmjjhgykj0uSrhF
Oyig012ktbEFtkCoxN3k+pMRhJbnZNiLgBfgmxnrBIUPGj76mWlDln8tTfC/QsX3
lfmhWdomk/ObdkGqNFDxEeY1tvD9pXJE/tF9XJpKm5ZcVdCTsUwCCuUYJCo4Bum0
BRqo+4J+GsEXmRQ9Y1hxEDb3u5KqVrUCU6oZACDFcRdSRiwTKS6CVy9KK63XFZaS
1Py/gdHcjn1gy0CXrnJO6NajJfFgKd/ZxyoTjR8/G/vMSQahrRHfnacqnZHaj9eN
Ttwg03YZqV9SUi3eqG8+H06g/EjB/5yeIdXebsKE5Y6Oso+d4zLbuCE1mRKzWH+7
W20ny70a2csfpiog8hcZ+BMkbn2J08toVxXbPs+yNsQrQPktmIJ+abG3IWHKtjFE
fz4HipQqwCAyaYMGDVRHde3vjAFGHfrKOfKp6gzxj2hONi43aB64dIJwd63PCSEU
Rsib6+vGdEe/UKdS1xlpwkeE5FqS9KqTBjQuZTAFwHxBd4bjT17S7mJ/FqbTUC3/
Z6cn0b8SXG0W7nkfdzgmQTBaPUcXvmJHaB6716NpXkEZXNpe65oGYed0k4V9o+sV
aksvxcvbbGkqpqQRQZhzHTjc/24VipZUFyoE+QZDBltEkQ8PNufkbH1mXvEBHf/Z
ZJKnz5dXpnVL6EYBc+X5SwvQdm5CPJMgw5nOSmYz7qAU0xIyPmcP0ETHpBQ0ah6o
C6VX7BrBWji+7UqyMYcxurT60lmiIM+FcA1LxyqtcR606HR9K4OVLQBuUloAwY91
v+mYoYxb72WtyrdrSqxzvgvmnk3hnhxro7p7f/g5utipeewIHO538lzdjGp6IJso
KJ8QqPV8j072QaX0pcpFCn00bWWYoLVB8KvJZSGNIBU34l4Sz5ROhBHxmeVWU6X8
32v71ZXyYn+IZCj+tgERKgerTW7fqouFRhop4YCEgIGmRJOlNRftiNxXdJ7dMpQv
ViixQ0bknwrGT1/Q9wU/XqpiY4UPOty/wSW2++DU8vYXKk9eRHwN9URbN2jzDU5m
nYwKdskEkmCyVO8lzVotHcQfJMdbjFSDMf1TuHbLPm/k2XN8R0fHs7P1hcQ6ZYvH
3QnWl1ZO/pxZvuvQSPvOhQ6rO3vC365HhDbE77/dK25GUZtVmibaUXYQ572KQ3Zf
WTWqYDU1lGlZ1kbwXxBHGVubFr97NdS5anVpIjNZszN1jR3zWlO/tT3ZMDFHyPdE
UPG2XxD/jy7iebzpo7JZ8Ss8EeXTuDp+hZP75cfhG9MHmUSDT3PGoxt9gnvFzt73
i2I5/DwrTutn3VMxQKhOEZFCcACZ3HrJou2JlFAXBFbwfWg0FRt1jmFeexTlNZqB
TTX6xZs8fKbFVovJCLkh/pdVfnwqXuAzeEK/Vsg3s/wJPlNCS5JpvV3/BgnQ7F5v
0AqYPtU6poULmCUPp05/dFXI9bfJbIuBZWn25cJ7uGeyllnwngiJWuOpFXnAiox7
CSN3cgfjAav7ER3xlGH6UfNfVONNA3ZcfxZksNkBcolYAPk15K5GJgvArh6nG2X/
/CmBwHW92QanXAxOx4B33d+JrM1LO7DTjy6WSdvHZCm4Dvkd2JRrgKCCMEtbDkgo
G6KCgycry+pJKTS28s5/8X/s2NcCHvx14n6pFcBBdYBLR3GbS1F4l52YZOQ1Kh+l
T+PkY6w7+Cb4y10o1t1fG/PEZ1JbfNtpc3XcvLyMmtVBqgXjYq7M0S6qYECwO7g+
I1gIl+FZ3HFeOyT3ikB7m6XfGidAojbHNINtTdz2jpZgVQhKwLLNFba/Wv29NFU/
j6kUetQKhElSb1Ofasw3f74DzKFx5liWRrSWzLMZPtDYvVWEJshyxwFS+4gho1iK
lfDLRE/RCYbwL4aR4/ZwB7zWPBb3sRfWtKdF2MIZgzRKKjy8doJ6/7vqvsbNUPls
Ucgz4khGpFQ0S3BGhhwT+Z9PWNyHfS39ls9OI9OGAuBsjh2OSIEuX7CrJFE+3iLV
/GUJMDmcb0szQML6Qw5+DDOVOfETdv4WsNzDrYWfezZdjmPOoerVu2ymzjvR4fJo
5oRarqgaVqXwdZdr+RHGCMaVSyy1r1xSuq0d1FQS6iMPxgdGpY76KStxkeYVznJT
jVILQVHR1EmqRMCRtdsoksFZjt4GpweKuFHiBLiqO4tJRCyUVDOnucrom/K5ymWJ
Fly/HUZNId68zCd56X3Quf6Yv78beeYy2j2rtrbnJSRko/7TS1VbPXH8Tz7ZpPoT
McYvCgQPth2DYEr8+K7QqpnTWqNwYFt5/LB7IFuDs9fZT4NnbUs4PVW0ptX1Te/v
z9FGS2ZQYwXjo3sFYm5UWQFMFAoCJ2Qq7VM9pb+ysjqQ5cE4Y4yxig5grTEOlhIJ
hDrDQndqJyzqa5Mc+gpTg6toILJheRCtJz3eaeWzDTPpakE/alTy5DFDHHL6QPcG
eb6KOQcB36j86/hyJXjlvJI0IVJiMGyCPDNUog4l07V4DODG0jYjs89TU00yGPBQ
OEcKGb1Z9utgrCubgpEPa9a6vDzUqNlkbNF32jNqIJ9tLJpl5jJWeCGEvX/DVpbG
+Dh6Rxqp9YiUltXRAVmZDlV9EbxPySfp46EtlKJvSjo1ST4MMZMljTkBefjiH6KN
OQWUPO1LxlJdV9I9W0o8H3jgYzY7vJ74+ZyLR0QzaaKo8MioO9bCmKgLJmuXV9pY
ETHsWUCZu80Kg5lOBPpc09irbiK0JQNuoh1mkM7AugKVtrYxscjkh0MpIL4biSIs
DFG4dKChVTfWgo5qXXH9ySmc3OODEWa/2aCgrNiaWDeQMzDoT0Bg+V0i9iJUy4Pm
yhfqfobStIYXjWTV6nGj+lALLT+YlwZsRhqxnVtfv+e4fLH8EjiryP/LSEik33h8
k+yuGzfVdHc1HkJg0qYbbyobQHUBIj035bPv6bLhHrckYkG1e7rOsctWlardgfbe
Y6N9GUHTquuWLrsRIt35cmgGtVHDJk74GZXRT2qHKzObNTUK5a3+8RyYuLOAfWnk
u9Y2uoFXSI8YNB0EDJ8GN25AVD0zQa55iF6At2sFZ/CNrirBh2Ejt55iZ4dUYo68
izNpqI9v9eCtCK+6NMg07FB0bSpk9cSQr3+Xd96lvZ2Q0z2XXowdAa2u8WIAz9Vl
GsQmXnioUnOX4AiJ/rNeT0VKxXGqw6joZUVwArzTsV+hZwL72+nNy9HpEV+F8a6M
cQNpVqgT3D6I1RlUIswm3+9IRHOjR4kxET7GSmlldiw6OzAdpbsIwDiQmqp+nWC/
vHHNNEiKt9k4FL3MFYKb2GVxhkHNqp6mOerwWt1g6FChNQQKNTtwMAxc2FMwVzOv
rP38wxmncH8ptag4+H15naBUJKCk69FO//cLfJIKScnuXmbGCB2H6dOhvxMr4TQB
Ic9dptS8+yicSTOGh8H3oyM9ofayK22x9z+UbZGaA1cvEQh4of21v/9UV7pMLlgf
B3yTEj6Y+4HyavdejzitLieWl0OCBQlHu7q0NFYLAGhR4QgC7IK8iqMfAchuXjzs
UI8matH30yrpC86yD9gvrkXbIHopEUZtWqZvisTNLF4OfH4LgMDC1wnGMM+sHJS7
fftLbDpYVFAhCJ4G7TECNl6pJ0E+x7nVQvVNUTXsfjm+6O74BbuSeaIQKI/3ZyTU
tVQrMaMvxqCJK1xsL1IRfz2l92VlJiQsG6ZG6WZwr1tuyh/Mx1y1OrzaqM39/+ub
uER19ZY0AIqtKg90sG1LTv5dUO/8AX96zMYcke8oVtq8agtyAQBN9IHEmFz30rEv
DRypvpVFdAdL9zfJw3G/c0/1nWfVoQJeavOIy3gEay43AeLlzoD5tkBu8lxr4zlX
70Z9I9hVyFKEGimyrjATGmPq/hDdGWc6gt5p4qH81YuRownp3+P7SEYDbMqs2X2d
UKdA+xMiNeCbQJ5pmZpHjtYdpoCABgTQxBdViUDaM/OTlbEn5jkDjUy+Fj7gfWyE
fEjo0vNS6a3NIS8+xqqwr/HmIJSuRpufpTXZNpl5FJdZod6eK5X0S/374abGFUpW
77blnLw3ko1BiArF6rY/RYaJI/vWIaPJXfEQYi1CMVtdRrDwJB8tF3yELx4Nrxvg
d1FRHk6JkMaOS/EXLAjF2Wzz8huk+U4T8i6EGy780XwUuezP13s3ORXZmT2k/b+7
iX/Wl29JABi/DuLkSCJwkMQ60EIJ5teHVeegXFaW1ePpOHoCUHRwsBxyiosSOzLh
XgaDQY+OHAGhI/Mv17WSeTZKcBKHPWokEvj481WfROVk7Gz9iZWid/qCZcYBGnB8
awovsW5McxP/7Asr/dmMy1qOpWhJ2EjiIH4Xw5W19AnvcR+sjHrg3jdPW8ya6GZu
N+oa3gYpJWfWjQ6aj8BCBi0LDJGG1w8Mijugvvmc4dcou6srhTyscVs490aaQD2W
L4Gy2D/3ecgbnsGEeFnu7y21Wm5RQdz5H7jCLI3S91yHunKnirbvjbbPKCaMhDaI
nIfSTPoZmG3AgKMaHMqaayYmk9vWenp63I7NvlmICOzcqwRito/qXS3FEu87QUe5
MB+axJkkJEyErL7nqZwxDzT3HUP1A93xORm4oq7f4qTh0pvN9if4FHY7gX9/7hF4
4bZU07SPuMAkD+MctVsOcVGRwPlpWQCkghxXAU8wN/fXKtybG4QXuDEgZznpzP9a
e6tLx0xufnE6gH5+sUxSJe0T9q7eCfkChNSfFXVgzoud4++uLjAc8Hn9CaRyPoWo
oo6Niv5O2/eIerSBR5kEd4lSIsMpFI/LoRRQ0tczzGFsghqUfv/Q8AfbVnQ8uhXB
BWSl+WwuoAKug3yVlWNs993MZo9/z/BErG+rT4FU6bgi/No0wr7afrnfX9g3fFME
UbQatdMUE9ggYLTwJBulzwDGkngbCPGvlsuKPU1u4ghG3NspgHluWt71+pHv2/sg
BTb6QGTJlgGcM0b/kyI8gGghF+gddQdclqdeIWVcgdGLuz2MftRwYjc3uos56kxO
rAH5W83HfrgHFO32/vFgiCacewgWDVsJqE5hSK1Do+dfWY+BPBsDEQQTmh+tTdFP
ufbOvGvv4vG1xvAjeasgD8zHtknLEHH26f9qHqa0kl/40iECFVEEOyDy2tjv6sML
MnjCm28zQedMFYC8JeW3vgtTh4zJgD+CuSpWacy72iRm14xLYSytva6Ms7X3XCEt
OZtniwDgSr3YQbtPrwtqHyps5mq7qC7Hf1l6JS+HhvbzJEn6MMqTX/cihQq57oEv
/CyVz6PHbL5xbR/YRxff8Mywpmcv905o+RDFmr0fAfrg3KXhEzxMNFdMZnkyewVV
0DfF1qS+0/QddNSf6C/YhOchrVaDml5HlteAcxrWFZRW4/IuBSvXR8ez1NRiXVr5
8H2TQUL/LeNo3HJr+eR+SGplcMERRVbNbkCAFhCMW8xQ5jni0G5otJiQ9DKMwD5F
3Kt8c8tSGd8rD8ejHYZ71nGt/J3wnLduvIq55J8IccRme4ZXtoTfc+5G5MrCh96b
uJuxJ0O1JZrIzLFCWWQBg3/WanAEoVp2MRZbRk6sTjCOpQ1GxcoXLIxTdno874Ow
cdILaxoRzwjU44PBSMP80nFkqrrU/5iPWVZbqyWcbRuG4e4hqHB7JL0Le/zj/QgK
nm4frtRC4/83oE9/wj2gC+t6v0CWVBmJGXQb9cqhVjt7nXNMp7eqqRTpoyKES8pJ
lDn2/O4P+jaxGtNoOW8bdwx18r5K6mgA3Y8End4pGyibIThINTm83INOcabqlLI5
dBUaGyLHvYdHHCYhwhtIvQggVye0ANyLIor+PjRx0j/OreGSCfUCJ/pZFKKDSrI/
qEqLhzSYjJEGNFa9RoNyi0SZ16hhpmCyhjydqqJycFdyaGnWZR1L2u5DFU8CJ1RR
wMc9XQ1xh9VH0E8tNb0BPkq8UHZ+le5H5Srx/0/UhjjQXj7Tg0Yp1q626xr3t89m
EgX8UcudvZwqHnoijUwxCKc2vZju/LAsp8H9y8qqRpMrNyBWNEDYXJF3juNpawuA
5vaHJzZRuFT16Jm6kLMVTJJfx9jM2WtB6F6xNeRRgpEIqjridXbCX056UXhEY8ZN
NUrtPbqR12qA7Ws9G67a2w/RFGQsnyGWe2MyH1wldbrGMxixpswU4zwvt4UcixLL
yqMn7AKvW/gTDoNieK0US+6b7o8xKGoJMESoLm+EXTtgFbshwg2odXumEkQgoTHP
IVoIUoVXV3E2qj/lS0o+43SzMgQ9eJURfv7zl764YAgNTkQLZQeyjQne7scBPlR9
y4nX8Ik7lPjdhbBtWAIxBD1Cq3yGYOU9RoSCdCWC89a6VFsHuBwkYAUBHsX4mizr
Jc7O8Lvwb+5kIHkBKAhr5xzSEkowDT/9QtkJE7VkxQztWSkKCwlRMEg2NWsNkheZ
cjDKFtx3z3Crp+27iDFv4UNBsB4oU2T0jYIu3xFiT64k1pnPeulD2HuDoq9dY+mF
ifdAE+a5Fhr70HSq4ZGQBk7ezrlNWnGgLhc9WNKARonsKxXbeEA7Fvbt3+izDhcl
BaDZyOPMIPwqDkm41nWQ7fHLmY5HlNAcO4JG3TUShVUrnWb8m2/kDNgm/QpUDx1l
Spl0Uax29549fL40dmA5pC8wzAnbm83/5mIe9Rw066CrgG4/duWG+keIx5yVDf2M
6d8ziFkUAcqggRoAAi9NLvD1zjCWtitL8t6CqA2RIxkynRBYLuF/A7PnczamnZfX
5k5yZoD/NcbD52s6fq5MuxX5owJXnBng92Ef6B+gC8Mo8h1ntmpGK9aiGhgA5GNF
2txtBncOJsje/XY3WlthXpZejQ41wVYPROw6ji03XgQxb4qqeeR8Gpsjy+dyqFdG
fUBqp8zNsqbG1oNAN0ly37hPiOtpTGU3JIKHGx83FlQo8Kj1gDsMYglBvgHByeKC
aSUUETGxp7o0Pc83+Hs6LyI9SW11dn0tgYBZkxCeRgNcd/vavFxWHBt8oALIsXxI
Xe7yxTrfs43SgH8X7vImIh2rLvj0qzRkjmG0jUBAl4vIi6DiLmfbjn2gF0djNHRr
uochYVXCWQcdDn2hpY2Ss3DS9vN1av0SVB9ZFZQ67I6n2qdlFn/tRH0GVe10yFiI
e0QGGgreWbSEtm/gvYMcKZhCCqgK9Tu+T+LMMLGhn2Irvwyz7ChmqtbtayPTgAqa
uOJCo4tJVQw2NJiSEfMaOrzRuYYix5Iqp7XEwivd0Ge5x+lOky+J7b/0QomW6wYO
wu7oZxEbdAsBBnEUd+mZCGUoBPu8YXIpMBf8Zi/aeJcOgtYHEZM8OW1EZf5ymLDL
uVDbQ602QkTVJTksFN4ZZfFX4oqRpliwuXCHiXLWmRuUwRcfgqTdbxzDNAP7Lyfj
rns9DGT/omInu8q1kk3y9jQnwVzZPlwHBXYZn/paWqPu2/exeeEcBBWWzOE6xGvV
rNsknwONViivDMg29kboy4FmHYlPQjF24ylLBNXTrbqVhN+37BzP0kU8jbtuobN7
Fro8J3ALHDeiXeVmdRQM4DXjUslAWzqGAMfsh4jlCvppaJMEWyvHWshqFyYQxvGv
JF8BHml4ONMdxGbq7m6Sbxvx1E056U5Nlb0MAHeW6c/fwFnuQwld3fTzZHw5UpeP
XcG0581blgF5jHegsZS5ylTDXQ3/c4H3qpapZ/UL8hwu/bRij32SPK258hHQr5ek
ghEP3/44JncQN3+ntfcME/T1sd+Aq0jgJArWNccYh31BUtsKcATH7S1n7q++VUd4
n6m+34VR4ZQpO5jM+ddOU1yDtB0Pa7GZfZ7hBi8/2lFHUb8xp0tJISDsmAVvRXJb
Ut5U5o9uIEACrXTnutVGFysrILezfChtMOJDF7dKhAwV1XK/Cy7Cyi9UpO6VbChi
IxedKwokLTZoRlnO2GBZxJa8S3ENiQmk1hsNtNlfk0FOffJtOjlE7TMBOXDPl38z
PLnUevBNkJshm+SrDzxwPoOyiAqHyxvwhF3DpoaF1vFvNlY6FDj8qT2ztk7+ZqaQ
cNaslMbsCTHTXvF2NduOs0sdqZrrgytCTpFfeJ/Hg8eGD4gabaHwdE6cuwNpvHq4
aOaJe6EYdF6B6jhIrt0r0Q0mKyOo1IRfZldApi7WfedcrI1lcsY0bjMc62brLkYs
SGVhMRmJh61OWDDy6gLjc4AGZ2fSCfwyNi2JDLvUiF5WZXlxwwfWM/zdxWKk9in7
DpMrPOCUNBLfeRfUwMo4Psh2sIHyLnKvwG375uBqvx3H92r6zlOoE8X+LAHUAwzW
g3K9YqB4n8toPbCQ0orAcUKC2+UaFc5/LB9/yHCG0SNEXE4B2LtaRi6HFr/i6UNh
x0cA6gc6/A/L0cNhsDRcgA+Ti2+IMgjJqbvp2jfywpMDhIIYFZ4r+sZMXgJRIlU2
a+Ln+HIwgq2ct/m7lgz11bNoYgcITv09nljqYwmGp4SHt82jaCXia+bHi4NQ/esp
RaDivPIvgdjglQiOMjkeMchMG+5K/DvNJsJiNoZfD6vp79EFVDzYdjivuiyUBxPc
uEvHDxN+qHHqPA9qkKSbbusnJ9+l2vmLkRfR5zSLpEk2+qwA36/zuTY1ClnZqii9
r12AYQiF5/6CkMySfZOEHipZKR6H7vmpTzJ48i51uGOfHvBH301YCGrNvCZ/75eS
vldwfkzn327s8g089kntpuWjppDBbzh8q9aGDV/3X+yAis/xoZ8EVykzCfsUU3jS
/JrRAgiz7BCJpoZoRoGbpHny7rYg7uZJJJkhTR5lhrAWDMtZ6Tzge+RDgdwaHeGD
2+mghjR3gYYhbSO26PRLSviEa+S3udxm7plkvmlSF2+nMpcwba0ivIm01BgBmyQ3
/bjCrLOV6WyNHvFGUvJmbJWdlYz7gDBS5WNu3gDs2koAqxLTYmq7pMHTn6OKFY/D
whFPBMxxiy3vqjSXNGf7rCb2ozv2+Q5CxRykq/9v+OKM6KQm/E8JZSabJ94RDNes
eumYGdkHcP6NiGcUe2Jk13ScIbdF+RcwseVu9MDAXJl5EGa/d7HT3FReXiGdqcMb
1v4mLpgVewgcqIU1FMarHPoA9jZ9gCtcNR8Sup/hQorN08mZiCsfp/RtdHqei6lx
jP+BMx8D74DE7Npp/ZnKHQpNoxeY9OjewMg1yVsaC8tYJaDk+4DDr6fGIznvxVdS
9/sU7tXSwyWpqsfZivNhbzpu60yXV25QmBemR9U0wHf5QXKSrYOY6CKuspeiCFXW
D6N9wrlKYhEdENWuhnN2hwVO6q+TdSsb1kIXgHYAyPMOGTruHCgKO/r0OsEIex6s
UPxAX3swRj3GgVvzpVAlEcZiLRyJbwTfIpwdsk0E6V0oAmbWWPp/zADpmDh4pC50
ewjFs9nHvqfWnac497u65BZ2Eeky2nwIJV9vo2/AjtoHxwKCAzdVfkiq286Wmk3n
8lrDFW2Fk+1wO+U+Z7ahbNkn4p6yySc4Nc3mr+9d8N9o7QxwwS6SVQA2ogvaiE7n
5LVyx2uRXJ/12dblAJ+Q2EgfciCWytmCDFmMYvkgcc8vcjp54aZWScdlpkCrThJG
8OSqOFTJM3l5dZQLxdKanO/+vxF6ZWnfln99c7cKcL/UjCYuNM58IvYAktVXVe8L
HL9iEPjwid0oFCFgoB8QWWYA135gckm2mV026S5nyjnP69VdDbVt3Zb+jPZP4l8y
aaurtvHNhzG71B6O+cZFAIibcHihrVq8qpalqNBrMAX31fNtIEpQou+yhbFGhZuI
62H6E2avGaGWAKbXUsalTCttfZXcEQkaQC+2LnWPvD7jPqoOS9aGVr5Johg0k3Ha
Wz5tCmbRgdv4wmKa6qIWQ3WrVVRHVVUlEWdj6CELf7NBYPUY25Fh54DtZEM2atTB
YqKTnLwL4qR3jfoAr7hk+mr0Gojm/qjXVthALUu/0bYZgGwUI6fjjcTUiaZjrLsd
yQyHU8qEzouXjrJ6XW84xIwPidnWKrVQOq9wUto35Z1DZvWcWy7a2uiIA4OS0ZV2
IpW/JyYSuzz+QWnbxWdVz9T/2r22ma0cJqngF5ZSkZ0TNpvmjftGcqOSs3XB8TRV
RfoI2Lj4aazydKz6TwwjRl4uJEe9TktfA8TUZ0jVm57ONrViVRJQXv3/SGz7jg3j
iT5ZEoMPX++MirQkHz+Pa13eM5ZqMsF5ZUSAbV5rbVu94H+QQgEnreHNeq98STm1
hHdctuwZRH+LNAicRPtEleybOa/gFfeuwEvR8vL2xS9Z1bth/DGhjffCxtbSEe9g
UITAeyFuj+XQXiu3wLmT28eRZcUqYgqrRD+TNTSIeLfDhSdZUHOUepAXmdHN+Qtx
dKu1DIvnz6LFVVWv8cFFn3OJRC/TGRVISlyrzGKEB39JFmPkTtqEawsTNl/7P/iP
iGzGn7A9hhzkxcYPL2UyCpew8xOkA84anQ7fsZ/g/waToBx5rxVFkqzAP62+ipFQ
gAbcYUDHvp5CK/a25IMfs2PEo9EvsNj67lLjhk9nfRmav9Iclo9/6wZOhmweOiYO
0NjIV3mcPi5D/qZdL74kLwkddL/8L58yrFnqH4yHZ99Bj6WgdRNhsDF2HhM98eQa
T5PalUY+F5osAX97oLahpMPh2dFLaDeQjlxw20BhhAceUQpjqv7uoA0il2lAFxem
PM10WmYsQD4f/IVeKEEOY9V4hpbsMbT/m0p5wF66dx9Q+gN9ZnbMsJBELdjO8qu3
iQ72An61XWrQXjEPe4G3/V9at6WHcwPmwO/JLyodduWnpbb9przqForoBWrz1jHd
nQV5s1Zymfl7Hpj5ROZLInNe7MYX4nGgVK2sqYy1jJ+Esz6pCKhpH4VGvfzxuAJR
KoroJMQd+6Ma9LZPRAykBqbvQXvbN12zcDTq8wkQ0qNtSoDI0gBCnor2daEnM7HG
6EqFNeteh+pW/Vg66gEPiwgroDjYaIdEH324nmtSju5XQPhe9wqSTwh2OZgziPYD
8jU1lQVG1tExRb0EGzNDZQdKWg3YGUIC+sJbi6k8Si9Of6EGKCS11tT9fcQuT/cE
U1yKd/HJsMg6zzTY51zN/rNAAIPe7SmMsEuugLutysBihEmF9acs+/WNW7bG8JIS
7iItA7thGVQePCead9aqqtEYdZiPEfFhHuE88QGsbuuDTn6wDDSevlwPEj8nzrLa
gxbebIBdHN+MBYBniG1x1a8TIh0Js75WnHrIxs2Zl8yfonH4cbUcTZd7xes5H+qN
l4WK1C2FWnbxIoPQFxoEcArKPWFAItzPQBg9CDoOPCNF5hRNY5SLZhNKtbWegTqc
xAO067WYQybJ7LIu/nwrt5Ue/GuzkCvI/kmggkfjgw05G3Sy14krveoG4U5YZ2Ik
j/lpHS3NoPMjA1lys+TERotmrFrz2plNZnMSbPUR/v7yWGpcVx5GoRCFNG7tbWT4
AudiFtTTdL0LnHNGCJibw8RdnLjg/buPX2sNvNdoTYoarFoZLcU3Iyv+YG0sZMez
7NwFIP0e787MWObgL5Urn+ESm3cAWqKUzdK+dJdUprCy8Rd2rLhthl4rEcErmG2k
pVQ/UswD6++aC3m4ciAtMg3a6ukXBq9CGXKbSo/A6wpETTawz+5WMk82Q59ukJaU
QnPjuDeU41Z8MC26qRE8IWzrQTESL1BPJZcjLhvD8vJrQPuxE+LVkfWrp/VjNzA7
NU6C6GBQUM1QfAb2QFcb6MQ76AN+DrgIwz6DNZD8MqVh9HYco6Lee3s9PgMQQCBB
yi+DUAekEVu5Wv8eC5SHAvHjHyjd4O8ZJXjiYLt1Rb9rEFL402a4YddOqBvE5udz
DLR83JcZpO0ix24zN/72xYOGELcaKabltceZNsc7FEHCLIf0bMdb/vpY2DlEQ9Q8
TJ7B/VVc2ES1oedA4Q8nfs4Easif5SFQn0rO3qP+n8XuKHu44emKm6yJA64vFPRN
2V/3pQtcYdRnBsl3HtG0pmOHlfHre/TAIeR6ZlRf1Rd8I8ONN7y0fxgWIAq6ZD7p
JHwsU51yp7P0i3VLzfkTzdq5P3ImtTu8sm0+N3H1OtaTNOSRnUigzLndDnyzDzE4
FmCoeSkaexv9CE2SpcLmTeUTY4zxgHM9BdD0hkmmJjC8eSWngRYIorrAeGZ+ZFQ4
oS1eWxLcNKy8Ky0k1ilztOjbDg/a6h8ZC06qFWCO1aQN4kwzC50g34nN6FMyclOl
BDgzSdy123EZV1hIjsWesYfMUS/aWNyd0+1b4aoXwl2RKqt6ZSjSOlZqlRf39a4d
94UHzpwVZdr56hgXVRkVHo16GrjODk2NXKnYWC+uH34Tl0PJYpDWektA+idXtyTf
csmTl1W2hKw+/se+b6xEKDCGcq+UronB6vk/BpFnzqQh+8bgH9EwgGth7YqZ30gK
DjLBmmFugmMK7jHYF47fyJgcPuelLvcKWQqbtg+IGPCUzmjS5fad++hnzmvIkXeQ
6xCdYbaDJAW7nDIqpGrmHGodqRvAbCx5NEk0RXRTzbziK7y5yyeeMdzoVzNfdl6a
WYbS80L1XrjwyVzU7p2FM0mIogt7+NX5vI5r5Mym3uQpcyZgiuPpSfMFxp40UJt8
kTr3AfC1RTCTuLTT2psjuyHNicmxDlKlyphB2gKgElOK3W4KSkhOpeK+w7LYo4DN
/7wi6GmuyvQi0V77hswmXsIDSAFbLGUOOHIIrGlOzMUtrILSjDElFTERu+8olQ6o
29fLx6tHmWmWnTE8B23b89tft/jdQX5qymZEWJ86SZ5tm7iztHQryZVY/xht5Kxa
orrFyuFvSvqqyxH6DQ8oYB5EgLdsMG6qc6AyPB7Wi6+Oik2nQG+Yw1leABTPMAJm
XCpO/8T6ex4fuoYNPLA/XhWRt/jlLN/VxOPCHyr+lHVHXGcBzkeKTqYh9LiqoGDI
sWvXHS8fOKaq6WyNOo6W9FYKc7MFj6fxc27MiWFjbJeBA2WZvucri6pxaz+Q1rqp
iWNiBfoz+sXDrqiB7wqg00+KkC4GcGBPAkj6qOdGnRdkn5T25aLJ1SGC1LeYSxtG
zbvT9Dp8DmRVr2iPWueywmVwxfBXQ+zLyQB/nLyLG/raqqP9OsDF1o80tl0h1IEC
+TquMtm1hWptzv0OlBzTOHN3+GtcuO/scSBkeoTU6pf+RZh7AFMWGjUjz0fkwpY3
37Uwz0QJ2Y49cq7UTAY7TlRm2UvRXKXizLUXT77pSbIwYaDRK/rBUC2r6R4dP3l3
1bLjQGOaipiAzUexxtI1EPA+PFVLwdX4yX+g6Yqud+uSjjRn1U0F6BOHLIp7BiRm
ZcXCJTBRdGoozL6pXZtB+75zn9/WoGPJmTs50BcUKyle3WCzDKiZKo0ml2YQSK5T
iXwfyCAQy0Wf9D9yDA0jabgVl0E5vykBDx7PNUYjKHJ+FZVWIB9ghQRvGTzynAGo
C2FLgF7d8myr4g9fA242WP+55uipirgmODd4LblEDjmXMiuWhFy+/GePD7DddJf2
mBftJSUdmRs+3cx6R8drH0O2+NkSnhJYuR8X97zMR6VepVkPzsJVwJ174/RSNZ22
8GP9tDhuL19z0aOba2w6d9pPuERvyBZqKjajd/U3MO+RwSpX+CgO5X+HjsMnAmVy
2IdaAkif1gfQ1YDcQ0cf0BGQcr1NyMm+wfFWYmCeT6kNZYU/4z3DUWbvbgQKm9pl
MdiYeyeQ7mQVPfUhcjn1ysUcp5ke8Oy7u1Ih85CN4vRZ9sgc+5m63iLvshcNvGZ3
+SwluVz5xtpY+1YsTdKr3I012i0+EajjqWeLXJVD12rwTe02rDVgNsf2aFNAg0sI
L1gB82r+gbdANfkpemsgYx9Ydt/5I+UTvdeAr88PhsWcNv4kMUuRFtlSyGssxq0q
W0XfFgNsq36Y/2bYPA0v8/qwAUd+/+ZN7U7PVrnTU6GRfp2q9Hvvk6KUH2AISpe+
hcOkTbNsxnUgRsLGP+mf7BC0Q9t2OkPWILS2L5zk+oPIFfjb4tIKhxJHxresCw2n
zEbkEGhvrL2RDUfGXn6IyCvOp7A1P57/7GLqr5U4HQk3MOpqF51LiymMsvuPjCng
pgZqQf+dJC5ZdvKEXafj4i7Wi2asdiXJbxE5lh2P9OetYkNkjgosPdLeMGkXGOJR
9UHlJUErDYLrXGIzmiQZeQ90uR/i7bBIxNha9dNGvVt2Nlrwg12AtFWD3OaCHsBK
h8uM3Y+J6aarLRGwN5LYGfQiN5zh7wmBmMyPmMHyKAatA5r/Hrj4nygtmItovZ+F
hGK8fdPiV00SWYWorU+JA0pP09HRuScAw+NfzdjVwAwcgptUtEPupAc+MsFRMdKn
RXr/1EfYW/+SlwMBDSJAHqkU+c2H5HIVZXmu0h4GC0ipMeZjfKTDjuWWc33KI38p
XWx8Y9mTAkYY2bTWK1bN01YNHApDzZtmXdCw9602kKDWwHfoLkhWfhyeBPVOZN8D
T1sU84F2cqOqVZA0qrpdxVhHUHVb95jB74LsykF/zr4y1thaKaFbtRgWJ8Ib84EZ
5ayPG+XFh9Jeu5hqZ9AT0aNz7LOeSab8omQG1kSNQbEcZ61Srit7qDrK2/ZuRg4m
itcK8pOtYYC3PxKS4S4IOwb8rBTT+7rMJCWe79sy1VrEMThN8JA9p8rHHbfCZrOy
xchRACGzQs3YYYMQ9sIrYIM/rHHuXj5dBERiWWCZFaPq6eXK5fWK+SBTcL0zWMSY
nLRBRKUqBzZyGP0ubq198XwTzKOWYQ2OtDm4ai2I21uubL/h1iXicfZfaeBK0R1u
jLag/Pb/UYq617nxxIg2jZsi91ofGP6EgorBWBt+TibwQ/ccmhuMwN1YjrkSaIqa
2/f9d7cvglvIz7dOMxcPsyidv+zs/6TqF20+JpkhfS4YfMo7IzW0JJPCDbpfRilW
Nmi5lE5a0S3kCj78w4q9QlXczMJPz77JzJQJqtU8nMWAJildoW3FoH9X4jH1TbSk
QTUFeIr03y0Xin7i+HFrClf/OYbQ4XR3ikXEYW6HGMm6hAa8EVZbUwoeleBxvlB9
wAksAdvJ68qKp4weIDQFZdpJAX8VHINt/yUakmy4onCAB/KAp/gjHAflzUD3WYES
CHyijCEe5egW2QjsJp7quLHV2kz06/teFRrD3yNQSM+CadeRn18pSl9T3dG/ZN6D
JOCNwPjBYV8Qmp2XcMYRT3qoCYKAV4XDwaqrE8lr3UkEkfRF6IlrKnVxGP4B4LzF
ByrkMVQiJWcTmlTz+RSnbFHwHp2mthkqiQEE9jWH0yTtD8qNY2DIZzhEQ5twlViM
y9G0v5V/sv5y8ITwRPcfbdZGVJQFcPB94+jiDLX57KG74VZk4wxPbPf8QtR1HA5r
ENBP/wK5CY1bGX6OtE0SABzjuUcndOCVOMcVQgouge94/gAdU8Voh2SRBawRoQKx
p9BUBaU4dIEgAldinNwXGL3hzVeniDC3EbbEE+eQR0jjsvZ6DIX4hlUU+SzFp/Q8
2klgOcQPX7Mzik/ElN392bVgbD+trAhStZBrARijZK5WNBcGJ53wtsmnTnjGWlvr
bJ4GRKDGZsdp/R6NkZ48rLgkU05wb890U70j+wWZ6xtRo23+dYNIRtJ6QLVXG9wM
DPatmkRy2Ml/fVAsLl1XSJRrJrYpmujrrfhIsHs3T4CkEsDaSp+Y1OkTxdVrG7Mq
RlvwhKvwpjwgsCZGUM31jpfwCYjNU8TDc4H7sfkYWdMViaZex/Jh1aTxUnOi7bWf
qa9/hvgdFqoqjvW/FwmrsITSDacv8Z9rR+yP6FrNkBTSxbbVdCPoGP3NalWHiGQS
QKCWaZFJNQbE4kNTrV7s7hQ2+we/MCo3l8u0wEg8TuTuTuT1Ps/InHBNVFmkixu0
K3eb+R5KyVfrc8h/hE0me81vMe5icctKAQu0627oOonDYOmH1drljOdxGqNCn6JH
dNqZmmsiQ5Hz/x7UjnzGMGuM9/R7z/n6bOAXJJKJvo0CCzegmRmUTVd8pPcBOpnc
9BuBjPJaQSSHs+yN5jUK9u9jb6GhTDnVxPBBw4RC1Z2PoBv/6Ju0cwJMHaIUX4ne
cpLjBDThTygZROvebljHgTqgr7i1uNLzldICObGiW16m8nzVSrLSqGlZvtdwXA7V
rdRtKzfNuiNBZ5OKvCFlgPGQ6R5RbdPQ0Mi+U0G3/1gtGKLgxD89iZLcbrsP+tLD
fG1R5m3cDtkqjczW1Rk4225TTLJDbHdnQr9E/+rCOoKN6Tv2vCYVAjgZXy8pelhH
nDNCZsWqLxjYwwwAdjEZ15jm0c5GnJiCeIYsveom2dSF7bryYuryM2x+XNl26fV6
JMuuFSlbsqF/FKPKdsjZri0ntVEiBgwBbLJ8HCOuG0A/0PwMrlR4QA1bXZ+ECm2a
b7yLva+5dxJodcdgEnQ5R4pFwg0Jfaffu0UuND0yDBn35ckUf5ORYMd6dvVZhnqb
EBTHkGLPSZ+i6nlhHmpKsYt7UQFBzMlwCZvJbTtU0TdiDEYx3DAnAVz+lxJrBhbF
+IE/uUK8UxGzLBib621ij9t8e/kwKFx/AC9tYLvhXyxnoqNelx1fitJVe6YXx54w
QvD76IDA8/Dix5gxPYzAHTemOiaMcBYFqtWwgnmyrYoZcCvqez6nliEbcv+x3AFr
saRSRmOjI9YvWyAUiyzRyIjAjX20NtRES+TvAcE6+2qFG6auCiTb/TfK1PI/Ze52
oG3aoQ50TcBle8zVNmJsbqOIZDHdj6A/3v1kx7ehkRFc3vpdb68qKLNy7sKiIOSg
BcteyyKnFzJz+qpbGujL8mCVJ74I9IzwfoHnHmrKaAmzMDVaYBfiJgQGM4YD0fH0
Hn/r5ksHkJOG532KvzihdQD+gwzM7jEatt9FRq9HvdLdueqF476S1kEqCcyaCJif
3yGLKDm1Fw6jYTWGEr6BMlUoXiCnh3KaKw3zGDyWE+jrMtHMBIcQIUkouFO4M1Gc
HPv4nri2gSP3mQNu/Re+aaLve0HgIVmAyIQIkZLYB+zk5K6/9LC3kYB8B3rCbPaQ
ZOgSSlbdTj+ncTvubhbElvpo9kT6CLxV8GcmbiHP/K78sAsBCZmacHtzJR9zao8/
uUzMRyAAyWthARyTvEZUWriExro+jYMelmrsY+le7Hqj8dXhXXf/AcNIxfG+49Fu
lWFPk2+Ry6dlZcPeFy21ZTgaCcSnP5WSreJV20bUYFr3fT0H2I+Vgx4ZqfUqQgtW
zoYxPeJCPb5tXS4f7Ys4Xs1YGPKCgja45BiUMNnWM7sebX6IZoOVsCXhJ5hV7/NX
WJbn18GrWA3+gC+iN44gGAYWzqWGAPDytak0V+wsoaP68ovBwAc9VAp4H55a65GK
wjZ6mkogRg3wU6jWJVo10mTc44BSpteNJ1+5HM4XNIca7LpEtlCRr+4+Bi+93ZsL
13hDiU6r1r+4m2amYZx4ziz//ZwIz9z3WHXbyeNWJ2D2ZlxPKBJs150EQ9R3zVCn
QDs12Fq/ZPdedqySb7nPJdoQuDhXf01qhi5EyvA9c7eXOlJeHr4qjcFs1ungH9+E
Y7xuUP7pZ8ChInBIwDoWZsGM79Sl09TS5gERPnwKaFwQI8yVh2++bnfkA4jO7evg
EIzGJFLVqA+NK2pPPPNzhGobVk0ZxgbzGxzVeKdIESHuWB7ALtTRPDYRXzuvbyke
LKqwLWRnfI5Un4/uP7y4Fh4Fo20CSqrTUHf/4WbZD9NlVSqRwUgnApvPWpSegYhT
1RNAXuaZ0TmWfORlJbIV/ZF/OzOhvq96ORemD3Mpw7kGt7PLg7XUYYiLqzHRqYzz
s/Xs5NfnWzQUtrsMaw+7+Wtgumpu6h9jOe4/wWwc80ZdDwOKZzylZU6soUvVfaNm
f11yERmgVpe5bQFJtgVTEF/ntlBHq+USmZVC7M3wBS4N5u2NJPciJ9/XA+22Dldg
NO2PfiVTA+lJZVsjatfNLNz1wrJZ8HyfBLnD9+tvoSucyQtUs09o6uulSi3J4YLh
2X/9B6LwAs3MTFYycWfx4ebP8vhuS+U7iWLQEl7I053WvCvw2YY42xxnMIpBi3b8
xPQB9E9C0+JDyI4sQkB6y9spo3wNu0p5OzQzrk0o7NcMfj1zbDu/d8cIXZr9KYTU
Lbvy5xb91bTKaiJKIn9dB8srdzNrVbyFKblBMSzupN58kBflfzYfmLOhQtHkxq9w
41oIRDp9u0XFLpUR481jCuFIuuXsqIqrww12Tr9ZhJosHT4Y7xVF3Z7fxHw54enS
/qpKMSYC89Kzf3DmrfMXdB7Dm4DtLJTPN/rMazIWN/zdop/66snlfI1pTOIHjqq8
M/o8J0g8LY2dy5vAA3KcZmPlzRCtUXwls/clDJNeZpZvBz6L1qZ144OhAubVmyKQ
O5NXLkwI4r5BD3bk42QdvUQtQBRuXSN7w2sKMwGDhu9pFMYvwZuhcQ/ZCK2nUWpc
UvnwG7l+Pf/8UxlE1Vg99P7XCCcCQGkzIosUPq4qogYJoTlHIwzSLj9CUunYaojo
qI0m5Koqpjf0TEX8j5eV90Ev+C6+dxpnNa2wrQSqrwdz6YZmS3WMkm13clA4FqYa
2T6Cfs5OqpirPbxe3A7WMsBc6Lr2WI222kNXJ0E63i0HuZwsNj3wb1luuTPjR9GS
JQERHt+ZOxX0DHwCT+pY4BokBbC7oPHhYy2UHIWWpCiHIunXLxbIowiw+IkkNNFP
uvS7edDvEGfnyqzpi+92TJJHe6tIbZwJWjfWwnfXkdQqOmsTzAla1hD3pSzWCL5t
9GNU5CcJQMqT1f1tuaklSnBKaXtfTwXdiC2EAH2lEjYeVdCVJNHgBSKoCBFzJ38r
lC3OwZaUppzRfIUIkMoidvbhcW3Bg+Qx2MOTAKA+Z9R1YBxhvdiDhV8dbT9KK9LR
b0qpii65tTMAlo97XzSbJv5Q4QDk2VCQIE9jQDnQ1wW47sLhIoFa+QK+VyPMqGUE
qnAClBfnGVVduq5R9dVPPoeWe+QkMxrOOv9e+/IIC7r+H0W53fmOB9c9xmjk31vf
M7MgtUqaMB1qvuSJ3kQEO2ts5sQxqGn8Sg7DJy5oTtqxST2BTZD/ePqa7i32UHwF
UBi6VSzwBnjww5cE//GBL4wqZ2kydkaJxZWfYJIzA17CJusUUaJdUOrXIGGus5Zf
gDyNDgSYvW9ojl51iF9sNtpQwPit1rmK3wwwyp1HdRiy/5AuuGLk+qP7+hxSzIjn
sTOusngmQ/QPouAev9AAwlFI2RfRdq2SDwdDE7VKd2SA9PomCieMAChpcoaLRJ8D
4jywTgg7OiMKjiVARxyrjeLbwKfTjpoeKTgx7DxWQwgwR9ZU+1xovxZAhgWS2uEx
tW17zcnIoweY5XuAYHMq0bFmpv5LfgqYPgVJ5EKD1lhfCV7JJ/NCfrAM7P0KrCPR
2BygswqIZMDgYcpTG2eblNlcwCBSVoORzIf/mi2XjKRuBDIeZEwUuAlmwEO2h32u
6jn7X5FO6GuI3aHnkPhiL8/KZXTDGZeO/LRJPXTIKTlYhGrTYhh9+yquxGS/N8to
E3h1WTz14JPhbmXACwDYlYWQbqCPhmZTSMTszfC4UoFyYVGBTfJwPp/xQRGnjmyY
4ufsZvPuz1oCK9PyokrsFoTgB8MsXfD407k/VxexARpJl874sF/WupAS33rjN+Nh
dQ9img9ryPIBN7LrNIV+e1D1WVGJfwBEWqqkI0ZONlC8KG9sJRmj87xXBae+IXrG
RZ8fQzjJIKbrwEg/Tis8rOA9Ct/7M+qkJoLgCiHbupab/wI0Udv4fD86QzDcerVs
odD2/QpxyxtG/FfCtdy/v0QovTow7GrO1uAcZqmFoSehgmXvzfp5nhEoEySi2PKw
1VyIJzUTfOn/h/oKtLxA0dQbggX2ChVBuhTZhX1+gPHI3gcmQaMcGIljaHr3UAM5
AKi/8wqa6AlppNP7QCKU/addWnAJaBXaeiVq3e0s20dX+5jneICmU40SXKbTyG8b
U7BG/u9HZIcFPMwROxFNGSFMSMnYAurBM7Tc+XnlF1M53jG3MstU36ubXPc6cwI2
qt1wsNHBz/vSVzwJxWcerk2ynkEoFaU1fSUwy10h6Uto2E0a75L4YYMxY86AS2UK
rTxEs12fJLZH6ql52nXyXKpNTEpA5fKJdAcfMRRsfLOX2XzSpNru8zvjZYxPlBHJ
vx62DarL+tq8YfCEETznEglgOjQDXaUeYnJ5kdxdbhPv0fPeBPLBHGt4TbQ8TDzl
gNKfT46PyRffxcfCqPD0vQWqygiR0quscgavF45D33Nu5Fi8PzVxwXGtyHrj9B2d
UkLzw2Va3DfyIr6hPBIJqqs17RbhfxETcPGaLHOSeomVC+pqDZjw6j4lEJguKGKy
mUmhY+fUE6ZCKaomtZ9ZHqyA6cNLPjOkJKcorx2CZYSX4cTkRnO567XPmiBBZzsB
oTpLGoQDgSsjgQ43/qqdhu3TrqSiHPeB4aiYeLHyAuQXA8NYbbSJxRQuCDDwghV+
ER8O10J2VYPdPzxYaFrJ9PggHEBzMNCW9ShHB5zS4hXLR9l+l55vAitL20EwuJuf
oNQYqnAYkQTGqJyOGuUX76v1GaOAr4+SYnZksPFtYTAn4x2k9+m96PE9WLlbLpDw
EulX7AiTJdhDi8YzGo9/FIlLs3c2f7EtxahHT6nnJo+Mk3mhO9rF97czwdTocsTo
chdyUmuhwQHqDn02E67RfO+il9XhExsYBF4InWjoN9kJNlMsdMmLk/Sw+lp4YR2r
+boCG6dW0UsXbJ0J4OUeN6UzyhcX8OAixGwjpXdPS1DeyZzxNC2NaYzW9NolhuPx
/bZuBYC3L1xV9WD31u13qw7Of3vIs4+VhdfFnqQisdjVIRsZbUws8VbIp5/DRkwM
g+vAgNk8M2bs5K1z+rnxFUnDtOe5D/u1oBoAuEzGrTcIcGTVfUIA34R10jVUr//9
EU8XXzFVqoCqhdS4TqLVmrSvpGFdBB1fiW8sn78jZ9EawFvsor4v13UIkg8hGlRG
ie6VzcChOUBcYjgx7Z7T3Lb2YP1hk3z8lyfTp9KCJYoywqGO1WEie4IgdD9oxRSW
6trOkLg18zGW7bVdF+23NE6qp4XtIn/PClSfeTI97K0mhcrx+HmfenLvMohn2o/n
jXrz+CXLkWVgQRvib3HGLija52NHQgYo8Lc7QGWxGJsz/eNNg3Mbf/1uObLFrEu6
zKGaQiKnGQcEUC/E4XoH77DE7aX9PLSnMhOu+ZqrhHbhxh9eQ/c2GUKb+/llDfbr
k6UKI/U/itIXW7BF51Rt7qKl0N40JJZOiJVS2cHA2vPaGrHyfc1yESnfHvwYHlAB
uZEp+mp9cauqUEroXC35RIb7CLQU1YEbZJ2pMEwYrKnO6FQl1w+HFZ/KmreJCpVa
qoiF5Ar5FgakelhY7SNDoFEvJsOvuITlZY72vZiXTuwL7ZSkqmscE3XCeJ2EdRWf
0mWfnWmbUi/BE7lxoWxY16kJlPJ6uYv6RgXVG4BKcB2JSScGRTITpwd6ZUnHixhf
HTbTKlU8o/afFmuGGe2ZRqyo9W6Bx8My4pLB4wWMhOGjbXakugq8EaQ7tszybt50
nyVE/rOcjmVpzAg6bC7YydxVghjs0q3hnDw1WbdbzuCLTdoUdws9HibFAQ/DjRE7
Ly7nJgyIzgLOyb7VaF90v+guN4LMlG/qSBmgPjyVwrB2/9vChzFk9cDJLEuCNMXg
9V1KjV7tWgQU0uxIDetJ0BhdibC/mVvVGVzzkhK1vlrDopcyKsX+ennBXFHkC3oY
iVMPF4RtUqu6yfLFMnHpj4WzEZXeVGfeaklRbXwicFcPzPksZSd9irP/HSKoOM4X
u4UyOXbNkQB+kRNg/GooNrYfe33qu6f18v9mNUceycuXs19ayB1hITAVks3+z9Dc
GXULPjUyJJ8vLa9uPkrunitAPa6A9kn0Nktu1CbcyMMTb+ff1HRxovlcM/i6ifoI
vUTDmBNepDLpg9Fg4Mm1VnE64V5dstrEZ6H8+3AQKx4b9K5Ky+nNHZWZ8zQvM3pz
n2F+VtJ3SOkiDzj+Mpm/4jb0uKVjHCMA25V7/bwMlRPRhQFCgmqCEFWXEcEKpA7E
N/O4+7uZB+eVNFLOqXRglB9YmbsPa6HCZV7MjJVkWLgiSzh4A0fUFaTIOYrCX8D1
Jinaji+bQJT7wiy+qD3PUjTeusVO5AGoMeqCjnmVwNxAxAUuU4dB5yU6uUe69Aj9
Ng0ie8Ze0WAUGcRqw5SujK73nvT6xO2byaugDg9RhloBD932/W5lzmtcY/8x4z5l
K1AudBCna7DcqFypecZtJ2Bq/gBNK1/S/OiZf6LZbo2wPyRaxF1TxS/+lAzhKgJc
7pC4uR6DU+X1ZV4zuzLsbs/3Eu0LQGVTt9N9hxYKSl6RaO10I7ZPdj7AzqRfceR8
rjfscSwAeRl+8ltOC6tEqDsDKi7B1bKuU5vdqPXdGaWcJQaGnWIqCgH5X6nSWzC8
RM8w8haYq6hLqklsl/3wvaYcwlPf5tw7FeyP4HKUszsopLe+WT1FaAcGacH2X630
wEBuWTp85+5M9LqzWPR2uzlpeRAh0DBv4InNi9BjkW73kFLICvEBQXwmLfNIE5Nj
cCJiu0z+VGCbTx40r2wiBtP1rGXOwij7w3HEBU0ap5w0o6tjgCb/+O+CbsnRZK2x
Vrw/J48CLgZ2SJnaVN7MBasBjbQzDNVM0b1yi4XU/uko96ubSlJO0qxHUIhxEP0k
yzJnI+Lt82MEIhBFQMkhZZocULEeI9OauaSyi9S/bdcv29YTGB6zB4j7BoxU1wPq
B5aLLdindfmooHfPEkRe91mHvjnwE26nEdXibBTyV7ocmb0CGVBmCLgAjkRkUGxz
3cAkOC5WHf8GorScFWj7+kSwCKsB0vboSu6jG2knCWWVg0FpX1xA0luLUdruY1Sc
0wRaXueevzntA2Q+A9OlmA6Szkc90sW15LET7F6ZLBltNjlbW8BK6nnTsBMLGg7x
ECxMZ+JYtqndTIilbuxlNmbMYil9aJsBwWxyt1fSeiEZ5867vGl+v0nyRIenaLqa
jRdFkEWY4bN+9qCWbowP2kt9/neEJg4sm7wA3jEyNZZZm4xLgyQ46hC/16mRZWSm
i7isjxoGIf1WErp1PEKwg2iA6EBM44Qp3Ri7bTjqlm4B3jqOW0iAES0fWu5C6ICT
sYi2Yfp4NWv1lTOgifOh+u+HiHlN9/3MplP4b8VVltOL65bDtnDIlB+/Ph/Pgpq0
4U+qJWhxp2/twoqUPq6iaRHe5Yuq+cirjP8u65vhCWhCxQsjKdTEhgwCJzreKGeC
rvOjhCH4Eoa9TOvuZt1TLCAEZkbMZintP+3OZWoRNBlXkGQco/JCvF+VhKX9/KYu
B0gBysQDEjPKDt+4EjYxGxHAQMZYSwMvC5tEY943L4Nw2JPZ0cSh44oj0gzKlrKz
1aUUbE4gITOWTlBkAqmFB9GhsbKUi5vBNkdXpBfDxaZddSNUA281A+ZlqE2DmsNW
ZNrUZo3yK6z6BUIGOoQRj/j4Z0GovO5lR7GdypKs8CzWnwWJZr4wKhhP0czgdm7y
6k+s6ph3GmjMzvZzPNfT29jt/jgj28+b3maR40zp/EbgLGHj7tBHyxYwXZyzUUWK
Yg1Ljk9o0F69iSl2aC/UqudJUgKmyZ/tT8rZnlOwru5I+JFTD+pt0oU9nOKXN6WL
AL7FeBmgF81N876W4mct0QmCrqgepxeIeC2vuKyO92TDhSLey6l3/8nwd9XDjpWr
GikCFWQGQAL3kTu7GP3htZYCtKsaOLDU895pDR6RxeZfeV5QkNPBSrB4OgwwdaAZ
IgwyVEaSm0icHabMfxpOj075yfMo3akCApVse6prnOTAiM3HULO3ANx20UA2mfL0
8TlJUvtOZdF6gzQeSSxKOp22R+/6QjXBRP59DLAYzaZPSVXS1bVuEfvmIOnyVaUg
/iYAsBHy2/RJRT8THXJuf6dp/Zckt6y8I3ZyUhYY4bDbTmHvPGpmNfDL8QlD4s2i
ab1oHE4ZzmwtO8RZZ9gjJS8T+i37XLT/lU3itkL0xn5zuN9dS5fqJzPGWt1tM7SN
rt1hKFmyPJQRMLtIM8MaIvyCH/ARFxE9fdsyYczS8bECW/3RboA47qE11HuQq2dn
o/UouWwTxlLNnJ5PvG9wX+QJ3KF2YAEJVQnDO1fSfJLIdiExl6q4BSqJWDm7v/9X
KBKzYACGb8rnSQexN5sNDunD+B4k0l6gLZBMiVuCVXdSgEW/4/HQlDuWnrCkJL9L
IphkV4dTiPq+LHI03NjBtAJvl/QW6eb+4SFHm3f5KVfcISsbz1V9EreblDF0sTjE
ZkRbR+HkLOXfjbfgVHx40JAbYXMcFL/FIKP4CYfFYc7VMldxr/12hyvgXm5ZJ1fr
vsgEfpb/ujXt3NixXmMVvPZoTKYMWwt7tRu8D56xj29quUWlhfwLbFT8T643ib3M
3gmlhfxrvsypq4XRr0OvR31eb0vi6Wt07r1dW2GsJ14LZ6SoIZHwdgZS+rG5Qvtb
Qs6DKIphZZTUjtEpr1MgD3E8AVB8cZchzLcMRNztsITHzTsbcdRfxwNlCrdshy54
VdeaGc2jFaC5OUfWM6h1ys7/FODrMi35venmPaQI7FJXN+p687Va1bESdv5ZVhar
CUswE38Uf+EMq0ZfJ94maxk5orBPL/4Sal2p7gOPn2ZJDzIjC2pjkgbAvcAIKKvs
M1d3n6Kwg+WuXhcWzchWguNR9oRGygWOzfR5mtvjhO/ZJ0FVUVncefBnaYIT6oE0
apUSYx+oAk9vGvJ03YSBnw/qRKbDnQtaKbaeHDgn/VGXCtuyAcT2ZOCbos5kXsiA
sNTSDo4zbjAtmG26bQfnU17cKay/Q03UpN83Xv4nEVt704IQWWKf3re90puc6cMw
T8LyPz18aLT8fu8H1Ct/XOVvpkLGzV47+wgh4Ffn60vX7AZsEw/m+ZPykWlUPTf0
CigzrPMlcayV3Nh8wQ1ogAE6wASy0bTANk2PCwqJzBdZiUBI3kho+uYRfVYfs3ed
HRCMQns4wCMlkRCVTHDw0+t9r2XK1f4SnJZqQQaRjrYIZsZyfabn3k1BJuljGjnz
Pb+hIdBucUfSuyRQipxa8IeFz3dJLXOEVPyISl9/57o1Beys3affKS91QA2Rzdtj
WzPsS1E07kRNCLl67MrcIcc2j7+U6wNrjDhNodH8+aZLbUwt6rBAdARVRtMQHl8J
Z+xMmqLbXT/4APxnLk8UvU6oDilfSYgBAZ3AyFEcCS9woQTeidqPZSZ0/rHdMmoD
OtO5HfjnEwlhG7QQMlsTvsTp1w9tH9zac5Z3Vug8wfyvO8hEh7AJ7EdCukQ63M9L
84QeH76rFvwdoMkZiYQ2ku2EBpHARvcAlmoWf1aQHJVc1PU0vpH5YPYkg4lhB/4L
i6Jr9s56W4jJEbDttsVaS7ieMvjgXllBtTUZfNuLnxCEJVNqRJaQ3RR6LoMozCy+
y5M/9Bg3/mri2tlyg5LBEyUiNRoURYaKwxVGDTQPcnkzZeI2Cb+wCeg9ghjcjORu
+xatFvdZEN/4tpBE1aoMJUoZ8k3IqNf5D/tNveo/VH+Zegrt9Wzs+jEuRPNz2KBR
D2vCRunpzTXQg4GXkognuOcakMtnb4E/sWY6P3434kp80buC9ySxRffpuGfOztfU
KmnQ3Y+GlCosTybWzpNTeAA1y0flt0x+3ri6qPDUlblHT4loaIQaWGRDTrZjKvnE
kHqOdHjVIwiXpSdalPvI1xugTUkjCN7nF6qo1/H0e5re/cgURmmI4Z0GaBEX7s/p
y9fktVm0Cdv5vHExd5zPYHsFyRDlnrP+GmtcRl9OYST1/tGJfgEWinFZTf7zM8La
YiP9dDvoS6PeJ/RLfm/6Cz14HKp4kbjX/yCId6RLkCrgSTJKywx9uHKVlpApPzlV
oS99HUj7wn4Kr41oKi8TrVDu/73a/sFuB06sn1Bllwifc/BQ5A5lNZbQAMXpNzsR
F+6HNhznqMmucKY2aZZj90xAINNibsC4RIjLuGMMqPL2Y9aAXm4OomPpaMVJXmHG
1IXzDFMQ52HLbYmWSZ1oN4VMDjwPKuOAIkB8VA6qTwXXGgXeup9ZUEi5xUfAVvvb
L7/4OLO3ZF3PQD3ExSD3YX8y4sC8g9xQhQxExLQzaP3i4mUkV1Eidm33qzbKlwcn
d7Y35fT2QekDROyY99yVOajHlXs6k3vbQjDz0P6iS7V27eoqjMcF/6zT3RdytnhZ
Za5qGWOTwNT0IQsm5kUEySuoFi9l5E+ZSEmewRtUhXQTXFTuES/Wg/1RF11/mrvS
N5Summ/bd4QQjySpeKDkF2BpWYmDzbzGwOcjCQ75oIS+5sQBI1SR+Glc2plwOZc7
D78UR6zBMKmFQeruPXCHaNha+NGeqSwOYOA1RiJEB0ppvuBg4Sa4OVpAJTQv/Zcw
2cOJr1YIVGmvLdMG3AF18ityZ1SrmSsO6ZWvJ86GwfaVipIQ2eZAAPevMKtqApRQ
tg6VP2/S0CxskIvCES+iZWpnp6qakM67WRkT601N8f413pNO6rGWJvYmcYkN3GT6
07fEqnNdZgk/1CFXFNqMxniR0Wj0aW6aZ+USbiAtxiQemjPlPM+OXx1dWIny1SUL
UdokBcSRI30nMaFjQahnM9Qs2zWfe+7PdGOeDt7TdD+U01A1P235wpzDHW/PGTic
F1DLgGLAhpSqs/LiY2099ZoCPrV1k6XjdOkiZ5CtFAiLbsx5y19J8zZUnEp15yaP
17o4fYBGdnP1Dc4j00gKhHCmYRFbTTIpamyfVxVP8DxL+fyfbqN3bGCXkoZCnrGs
8OGpePSLYVxZnXdRES+qJtUw8WFkuH8S+uZZij5Tcbk15uM9t4a2a6erIMIqxTBK
ke0FoxYF3SCA/7iBSZ7qkkqiVExror7ZL6l4+T3/PkG5JtongiJPQVKn6cxxBBrm
wMkZZ3T4q/Opm3G7ISXuTWvCXFrEPmmBzR1idqmbtnxX404jh10yOh4Wx2AQfdRH
fYvOhPZ2vDZVXTt/cI0zgx2LVRdoubK6cEhsUNlZGUGjUXe+h5QtkHl38I6WJkt8
nLbNTDEzcPgel739QnO31N7R2/CWMH50bYW/FwqeIbDQ5XSEmvrSjGurm4+1rZ4B
t/si7YHUiYdpBm2kygT9pJwbmOmVMpnDNqS99Lc3d4az4svIvR1ymL4MaWsH+/3X
Ma5dzKh29+DLFxW42MQ4xcJLAvcaFHDyCYpxelketM2Fyb5rn+o33VmwK0te7oM2
S8Ob8IE6+5AIyKp4hw9o2GQyeAC6S7gBwyDhiKN+qY3omA8QHa+PtKcUOI3HJPRq
nVAKDoADMjTgyYvJt2Ntn1683yWUZTXzvE2a6tDW+lF6THHSqj39dQtIC17HMDr1
3zkvgrfzwKT4/DIo2V7qJKWpDu0pCCDbaE7ML+bDNuFa4TCQlp9hePkXyyaDGtYc
0tCBLRr/JsFCjH9nCpQQw5M3sfQEV5JoKMFkdUSudQktb4H107hsWynl8YKDtQ/L
FZjxwNFczvfonIc0LMFBsjhtdl7onD2HtvFBlsfdQU83srdhlvFJbfOsVsRZIWSQ
fXCxT9tudYeSkzKBh+JtGWbqUZzz4979leZyOyTdg/iP3o3T/yV/6LhPB0j9qpoP
+57j2SRRuPiqWehZb/NWHtLuBF3BownnLSmlrPArMqDUN7pc6W3lbNvTvHhOgsR4
6/LSwS6BSSjMcvDoehkH7Cs7H37nT+bqn/pjlco2PiOijuY7r4FidyoovOvk0mN1
xT4gwdKzPDeJm/ww+pHiPlWra9hdQFuZwJ300qxPhBeMQtTNuONBSOAvzSPDewUC
HBummyZzQcBOKzSMJCJIuW2+zhLbV+y6k1VlCw+cG1Mh6+brq81sjSxukSwYLApg
q9Lmv+9eF4sELUqD5vL3kRiFDmm1JVkM+65Z/EEmmWjVhwodVGM7iWbfhIceHNAC
zYtq+WjW1+mZC2l39dj9jWd22nvJL6DZt5RS7GSKezTs3PtM7K0TZX3OvPG00qk9
YcQvaclv4bcklhvrxYCa8yw0OEHVp6dT6LRwhQRTBOLrYSwfg5nTdQM/iDdV50ec
/gcl1bZSgqDsKj2TD/egDLNFFZJUTw0Gtp7Hy6RRXDO/gghoyFCmhf+Mx87epXGo
FD+WsATDBA+k4ACX/7ehf1XyhNK+7QoAEedzWlUDrj77NvickHywRit0Q3hnGVq+
qWwMURgEBDfModMQg/wmldgJZNeN9HrHM8sZVvNZuEZGeEKKbURm3nrtX5+988vO
SEWMtBOF9NfHbBI3i0cQUXBLGpInmp65fVzrd0gJd3GD/WjV/l7gsMgN5DDhlXXp
N8VqN3wT+ha/cLQnSFL6i+MjS85K/EYzoykJrsZy4Mb/weaauHFeIlQPXG9NUEvF
3qFZPYRV3nxUVCFafW6kPLYr5KBCwd8b/rIwbAN7bZMzgczfH89752lB3IXxNhqx
d4Qeb8TlVEBKiStHn67xRcGFjiiXvv4p/aewBJYcg0tKafH7OsSCz9JgXhiO2pgk
sB9c/Keg3oY87Whh9N+knULxi19OcqVCIBOZmg2Ru/RyYk6yyyNSRpLVKG0yfUZI
O3UcQU8ZJfNu/mztQZiLq6iOB2RYTFrHKDj4rziKFL4QsEHYba9jjrcGKogLsJzs
2abBygEaIS9atvVYxnBVroeT5TgCV2+PuK33eKlidz0YJ4OBhzg5MIY8aoNLkjun
9ztKY1bBqbhv8XE2o0AJc84R71n7raI9pPOMB/4UQYC376CrTuteUARfR6FjIQJX
8pOGAgYb1I8zOUNSD/pYGOnk3apm7cT6PhVd9sUYS4ecRfRoHgEmHf3OKPwtlvBj
2m7z3HzXEOx8fzOVAYY12YbIoEK8kgpCW+5euwbYLmai9O8X/+X3hGLrh2kw0HUv
CzJEa1Es8ReKlSKNUvRx6nfToiSkqRrY1NJgs1P1Gcq3nqkppYYJdtROYLPcSX+P
zlIwppGGnRmtn1sHIJ7a3KxsaQpOdPFUUjci2CGKMWSs4Idd0y4wRLP/gwtze9/G
PaeVZl/sqwRzojEG91TtgAO+Y5uycBuxHQduPskIc0Bc5o71Rj0QV6SAb/bB8Qsd
laW3A+EvAJflCPttKoD4ObJr5l8hC1R1X1kXQtdKVwjAHr8G+4XTEbKQZP3jJV8J
Z6IX+78FKti03INuuYpkXRhYhxeA3DonR06j8GP31YrKtzkH/BKSlv1CZfjNqvNx
xpmrC9JsRRV/Jd5ezTQr3BtETbGdhWYSXPbYY2TIn/pJDOwYAC5WqBUc6KNV5frf
v+qE+yoKNjSQiwMjsZSSzoaCIr87ln538OUc3B2C7bVFh7YNZ7Hz1PAe3AJS5swu
Ff6zzm5yDXcNCoGMnQn+zhsOlp2JIZPVvPwHWFyV6dSZraDlWWrG4ykAceCsvqaJ
BeQ6XfAXXd24JzlLD9CvTNsj2DRTlUKbJFbDkmf/DqruGu9J7jCpdviQEa5HuXIh
TFU5VTBcVx/YwZwIE7l4+LmrOx1vYc4egPh4ZS2PyIo3CZLwy1ZsxGErxIPz/vR5
wliuCnKtiXz6nITZAiO/1brd0BV21xykGBslthmn9XF2NHz/D571uG6GHY2eQKBS
MNN6XcRUyiGLNHyGD/BbwOlxr6aROi3heCGoJAhHTubD5a+ZA2pvsLHo6eUCRvN2
rusCYytCLzwH5SyqHW7kbxrsN+irjCGGDdglYzPLWw6UKGE9eBjSK4Jqno9Hb+IT
XOJUhMULtFehVXwsT6QgFkCPuUMlzxOtgTf5xlpZHf1bL7AzkpJ+UZWwP0uaSBi8
UG1my3CtQhPPYDpZOEIZ1tBPZMnv6a8koECYYFS4NuqMvpK/AbQRiFOTWwGElZ9T
YLNx0+ZZlQp3PRDT8NkRm7YEqDZR1HHRIRCb2GPOSp+VTIuO49vglanLX13H+eIn
rYWdswEiIqpXhFZBEOHayF8q1r02hYI0/fIY6SQ8UzTvPKrQOJdeq3BAu4QFORty
qgy3mhHKnCU7RPTGGKQOJKENeG+GGcLDlaqskmmzpuDowpk6HXRGeBPr11gYYNr2
P/PG3RJJQOPu9tLgzcZ3WQ6ibG7v2L6wZSzkurS7+mwaMynAD7KL3lNxEVuf7aGf
jlNmgck4Cyggi11Eaav3AxlmaAhfdcL6Tw0MZVq4qkhwcfvt6N1/wMyJPywtQn1T
ZokmsImLN6FeRZVtjmNx0+8Nvw4mymxnby2b8yn0r1u+vffPir610RmCCkuSTk9M
vQmCZ7urdojq+GsgZWWJz6DDHrWjs1s9cY94AfWHD8i8Onzv2En9u2dH8oSErgGs
c4yU4zhybVkwat4zQ7hZtuJ3NY43mLJsIlUFP2xjGd5Gr0fUZJDmpgVp9klwdH0v
fhu8QotYgNId5d2qL2jx1kNbMKvzemv7aLnbUmYeaWpoKiudDpDvKS2cstTxDS6j
uvbvNMddV8/KeRyuS4d8h7sX3qMng5PoI8MNcYVaHf9NqLdxueRf9t4Q0SM8vuiu
YTukt2EUjRNe3K2yrBC2q9uJWlfy/4qis9XrYdr8K31O53Fq5oa7HJzbyOPX0lte
eNGlQTs1ovs9QbOSx3SVyZ2p9YehJuWDzME1RYUMIYfN5cR/u/TtggNlsKbmz3UX
OAO7RVwa9AikHTYXmbgglG4ps5bjgnZt63rThokVDz8pQCbq+uzaBD0Z+KArAYVQ
pbPa5kln6FuLH3EGj+iiUg66anXkblErlLnYSgd0y48eaMKE9pUGpj/UZfbq9wMV
in/D3fipnsbsdUIhXKciPXVF9rs7Ag2pwQai3kshxZSym6QKjOxQQATui2rrfuqK
Dt/aC5ZUImQb56TESG2H1wUPCmoGd7qIU1Cr9oMYMqm3p4ZAcucwSfkPmOoYMIsW
F0E11VwT5HPZT0luENm/JemXLHvD2XPt33JdznAkxX6XHw55ejx8ix4ru8Srg07Q
ceG2OrbBmDlPmfyHk+Ws6hrTFXw1YSpA/4SsTQVBlqlDyFOOnZ/lyeCjXDxHPCYX
U4zQxBQyedN+cpniLHT5GyM3CftReffKW0/X+EsneU2mu4eGjln04dvtCJuXXxiy
0UbxXKFteDOaPSy4qarXg3ENQR38uz/KZp76UT3+csvqxel30yggTqFcKCrP3L/k
rvpqtN8TnIH7DOlJbuVc/sGnWNri8rvLOvgvY36rNJO4D9pESuW+eyzSwaq982e+
9CbuRAlpdIc0LSX49cP3FZRXc2zS5IhEL5QlT6KmJvZHsunVg4vIFI1ElM09KH/w
n338eKHkSjdnw58HNc6ivUtiFrpnjsR0PeTmhTZyRtAMaVKf11QVcuX8sda0CxQg
/4XX6xwKJCpSlvqqRNbBqph8ExCVvkdivfzhSMfqdFsVqmeqm4SxeXzqOlLJKqR7
Pm2369xQFtPszi7L/ftr9n4/UMHlQGcQM9ZxMRGC+VGAoGXDOTlW1hncprR+bndD
3870CdMpdfRZNuSdZk06Zm5wKQzixPcXWNJhs5Gna1Tax4TSkBKX5kVHNYY6JZEC
wmpPXg9GVgwKuQxV4sucuot06o11LHlYAwEEKS0au8kPkaFhD6fbQYdJmQbhK6mv
0osyAoJuO4iviAans/pmyusG7bBivxusWjACy+SE8spGDKTayNNFtNFAK10PqB2y
zzOZ8qpKyshjIgdiNCXlTzKxH1qDH5TpQypwQkX14Z9zjJH+SmZHv4tI9rHPJJ0W
K4a3BMQVt1ez/XF4cnJEUWulHsyM7Ihv7aMolvxa2ICY+29RVyGDr/oXACloCv2Q
mjORk3TIVUBHNMpMd2NDn8pC07rhPzF9PshYTW9aQxxoLP3ADLAsPcvRjbk5ojzK
FRUzSmewzop2R6epID8f/dUjrG/pZ/kXXsHL4hriC7/+xC3BfsBwU+OpgBwO8J8s
//NTeFL//bdOV3sanM3IX0QF3WGTvWo2noD8RyUoj60NNC4oSfQ8L8bpwvC68ERC
xyvwf4F68smLxGhfEW38N48EzqRuQevvQWO6Z1Rfo466YrjG8ypEHfq1zdFAgXZi
bBDUp0ubsDGNHViCEwa0YQHB6tp8xV5bCSKJIEZVcScuf7eoePvJdvh9CBba6G9m
ihmHrPYTr732SlWh6jXIXXXOsP4mtZy60zS1cDv4NJYv6N2GD0zVPKussyOdaxGX
+dfqyxfFqq+qG4UG8MWOhT3r+BpdXzPeMmvoaExf1Bq0X/H0NZOM+r8A8mDLYyOC
UTF8isuwgY1KWRnErA/+EPrzYmJQgOWcSQKfXjL17l+oE+DaxlUuYtg9W4ltfbV5
M8X2lEsQ3z7GrzZ0oxX/f/45zk69+6BKysSCJbD5t4MwSrQc9cb5isjSwr0R2Q6W
AutbSHm0dRrehVRObo5xYxvtLzGaHuytKBCLbjXyAG/uLyGX8y9d7n93S1XRbjmI
OqTwsdBMxj+Rm18Ir33C6VMs4bZ3JtTIASQnK+fnnZHPKYnx/Ow3WR/0UnTCBLP6
fs1nUQLlwGBuf0DB0T+OtiWuvrUNJ4jP6yYxoCS7awFOopWk9+aq/FZdJcHsa4NC
gMGQZIJMvBN1NDuGXby23AYtUKfUN/d72FuDNyxZysT2Vd+XedclTWrwyCMjvhYW
4r2hNYteBCDTIFd0fuFh5h2vxkbbMBDJoLt9SaGWI0AMHzyP4c38SAwN8EwC2Yk/
bviBG4m1ji8+CltpnvUGpphe8wheUCH2bg8Fx8nIH7q1RK+3Q0WONeBy/ZmUENAQ
+tQaj2YTL86lEp3/QuFvc1HYaspFtkR9VWZNBunXr8w4i9a130+lQQLTBIgjdqUc
/fBOvUhqbiyLhjoUuowrDuBgliU3On2U4htEialQ0KI3ldnLcteP3DIP5+cluxvz
aQ54YEslUl+/tp1GIgtDLsWmO2yk4V6uTxqv6UVpsKdoHVwwfrZEoKrHFFn/nIVk
qpHubQHrHCS8np3nFOErKbasLQlxPRPh2gS39H8By0HR2USjctfP+bwd8fGVAxgB
3WaYCAvuUriRv4IyKs/gBzVxDZIEHbrRg1a+qIzLYtvGeP43/aw8HeO6njVxcqgd
6vDqp68F5Z3GiHQjXtc93y2QtjiK0VEHRSNf+SJYrlAFdwzFmS79xNlRJ9picN+2
1iuIVvDmtoD+WDJ8fj4d8nFlW/QfwtZfdyJXZgXZq6MMzUyWyifxhBCrA8Jq/D60
LAE5wWJSo6igo9+Ya8eAcNVarP8SuXKodO8HSqLiV3+XEFesgbOuUR1RMEWqUxKe
xxse+vSsfKlQ7O78jhnF7POaRKYDYozQNXU6DGsnBM0fvlq51wFUJ2ecdUjWDx9r
PYguCjpEgUbR7Dld9KASJ394DAT/tyDK1cEDuzrZKN9U8IT5MIINL/L4N9SQSqHz
sam4dPW4S2U0VY+Lb+don8ciCoz2jkaVNg0uf30pmzx78FIRjlhdhnd1MXQs+KGv
ZzVpYV9VYVlfCThJtY3vkSSi5HxxQrpIMpJ2NBEfr081Nvdf3raTxzH4fJ7WGv7g
+hCHAqY5eaZelWzs+E6UrzWWrjDnbuZeHloVPZuaFcCWxjZ4VeA3xc1KrtwI2HNC
70pv4XmjPN3EO7tLMqilaMVXQ82Gp/uDcFzs4JOtdsqFnh0T7elQDiYkbMa2JkbQ
OkjNNSu/HQGF340j0M09HV+v1Yaks7wvC64tgjK/07ZG5xFgEHCm/hKLZBb4F7Ml
/oyHhq17myqk/0/lBxgwrQMjAsbU1X4Wf19se3YIEA5L6/6Hmqxf4bizjTEPMZYw
5Ai3cFWYJWhKJT94JaUybtfzfLLd/Cdd3cM/PWZIeDOmnmlC5nu4hkhsGEv08SUf
1KV7y2ZZ0+IX7o7AMaJu4zXjlhj0DQIy3u3eRlD3Rhea7R9xQxppqdD2Ab30mMRQ
U8PNSbNHCuL+NTLXz5zKnsm41PzHK4qUyCewKSI0dJp70bi8tpv3vNJ70QGRFvTi
7Vau60NOWxPzLUdim8sMneqPPOE2qi7othpBmEXyCnF+9ucb1FLPNFkFfYs1MuEL
PyA4CWLtcxn905TRd25o5pRtC3C+R0Dh6gtuvRo2A66ML4e6fB/CUgHYteIlqvLl
7/Qew5tFVzUheMItyTLAzKXdPJkdPU3ehdzzo8xHYaOarRpEnlZHi5XmwPtI2PYX
0gb9dzxnQeIyzomalL2L+ohVU9ay4Sb1uw7kKgYZxPsTZSvx0IFhnhAC1Gm8l1zi
HGM6UbXAuUN9+Lsbfj5WOFYTi7Xz8+WuaPF7SUmyYFH9PAXMgddHvTmPlCnyYPrZ
u8CR3rlCOiRp8YWHP+x6oWpNAU3NuwyWdU4/g6Uv+pRU99GuaRoG6mE+Yj8pciGX
A+lDr54BmJ88I0Ahh0/5E2MHq0omHrNPgOplbuy6NsWVZ8ggSkdBfnEBaMX1EcCh
wFI91YOvKnt2iGshJTJDYh6j8sjqtsgZThJjeWKe0aPoWqAfi2lPaFJEt6GddP3C
J/wL2TKOLWcL0coYipThMzrC2hbsusSIl0Z3e2yv2G8wK6YNEMLXBN6DRvvoQMdh
x8w7qLUuaUhy3e2znCzE5lw11geEag6xF0X2Wm+VE9BcrJyAL6958CNktzcjqf8+
SZ4ftz829nr+bsqjzNt60Lidwv+ZycMNFH8HpSuTmo4vQbPi9x02pt0CHuXaAapZ
GkcZ4olowB09B2JMaW6eRp91Z6Ru/IUpiBTsJvLToDrLjQUX388/KLXZFpZ0uBX6
RMZQrvf0SDto/yegP9apEC/FExxtMpnwRqvjFbeeZ97v8WVV2Km0tWhBS9JPpM9d
/j3b2EdYqkPiCKPXlOmPhGHC/HH8eYAqoWotpH3pxooNtVW1ZorwmAfWeL2N5MjN
ffxYEu4Ajit0PEa5zIuXlF6IDpgabnD39C5h5gxFi0c4x20QwnsSXDZaJP4eT8h8
Y/tXtUVut5v7w2YQftDSe1mjq9dkNTwhAAr/L7j/46629p7htGGjlBZzidqlcBk3
HP2bJoXdsy+1vo3ZoWkddunqX78Oilh+ekA31pGUGTOvP9j9buexLiBD7cvezcEa
GN0oCy5s2zo3MOOZVxI8Yv91vlat6xHxUA4maapPIlcs2BTL5CHwRNRpb8gq95uR
aMda2Esjb/8Tjsyxio8AWW0ZefwxJqkwLEa4Uoiww3QtnQNfBmGz+TYm4G8L7ZFD
boW+JmSKajVjr2/AJWSX8SZJskMnp4TeEo04PmnfbvHRomS9sted2nEDZ5XqYRhB
u6zpOKz+sMysD6adeUrWmwhL+YWx6dRIPnWB9fENidk7Gh8YhWLs/KKdXfpZ1zXc
gCwdyOCMvQEHVP8QqjGCtzKtsRHYf0GOXiADgswojOXRDXcogP5+0pBOtc0mMn1E
ee/qwR+POPBTTgfAe2IKKJAzwMJPi465sUtiyxhlGq6yQCudy9g+lR6gwkXkKKmY
P99IAFqZUEiJ+fJOpGhUUm1LQ07kUOgk7uBp4j6ysGJDVGtZzpTk0KqHbea7E7pc
/hU1cdTmX4zIuPSjTLyf9z0n3huRtXVzJtei93uwByxTVoeylg3ErZbtLHHX0gH9
RD8CiH6RA3QMaKBUfB6yzZDvGe3HiB7LpI1jCk1WKfcod9rk5SKXgm68RRNdeB/t
2dAU4/UpDBpX1W3JTxWvdhqwdj1vQhAl8WS/kUJ2TCtyhiRigIaZBWYjgOdbqUfG
jE4hBYaYE0lIz8vefc/y7KiJmpd01QkbS3/3Jf81EYljaVXKR6lllaz/ALPMOgiL
AaKSrEkrmctwjcsJBMgUHXVAD6QriGKlgkMV4oNY5vu+Om6hxRYDk5+tV4GaT0wf
EhToZJ13b0Plm51w22id5I9O2iOjdIPcWR72dTcs+MFGIiZFKHPAl5uRLhD+G9jt
DXNVBDc8vU6owuSXSGxtDEtqm/Td8N7Ap8LEz1Up3IAHEOYCDV1xkQsfjFbcvlm6
37tuIRP9fXlAWnKkXXH9OcCUN+hOm//d/worTVoxzNxHILP2RgD6w86dwhGaoPY8
LMy8L8RJy+4Nt5eYrstgUoPXx+xOPzaD70D3P2DZqYq2N4WXNg+awvfXITaHy3vA
0cVhtkfKBDi4acDXaoMchCNWYsenYZ2SLYbQ4H4hMpDcXDFuTrDUptBMYVKSYmWR
FNOA7ghMPoAV19nh7rhCjkHR8cEoAdLPxJ6EwXyPxYE4Lpv6iu4GCrowpr9uD/LH
/PQTub0IEcmK/I0GQvEZL3y0d3IRgq7mIiWNCZg8OH8E/9G8yFq4D6aOMbJeqlur
g2U0KKmikHZ0ICaJgn+J1V5EmJDf5iuLXFIJ4zrMWUcvb3uc1uqZPjUOabkSVUnn
QQV/UohiYOQCNkXx8lsTHywSx2upv4ARQa6JkYHiKA3/GPiR1vTGx2nZyjjz5lf2
NzDOJSUGtNtN1Tlm/BX0jOumXSc8vwD9S7nhdb8P9hM8hoI5s9Fly39iNTXGShLt
YKUwXPNVvc2pRvwc1bSGByaAzxKaz7kfhOYdq6d05tBTXAogpUL3VlodcGPXV4ih
bTr4E3NgaD58UZtXsbMDMobOP6O9WaIW7KXfjFI7IFHoC483h/n5E8APJ8UfZC41
jkGgCGJPm1+OD6jkgxaVflMfmQpncKi1FUbT3UZLkXfmszuCALzv7c8c+KNe9mw7
lKs97I+2f57oIJ1bmKsY9+xLljt2tlMJM7ODP3YnKVGa0KrBZh3lf5N1A6KO4rvC
fdjqPWpmdHXb7KGLz+WMgvnX7EDf5BuNyNGFsOMgOOnmEIV8cKWBbQGFlccGmjY7
nU0Ijw95byv/cDrWo+ZITU2oOd3Uoa86EnhfETzqWCt0gqfYtoFeQ8HiPPduckfC
SnN1S0jVZb7vFmT3zp0wohwJ7I5yoi0W8/BSR8J5Wt1zlbnqTcV67+EturP5QpvP
KNHeS/v5/EVZeKKWOCis9jR30BnV9QIwul1SZgl1YJ7JCMKnBXcwfYfccsbVEotz
OnZHbv5etKNWe7tzX3AxOufetDIe9CBei0gVnjZDPCu6jR+H9YWkyiiZFmtU7OvB
nxXdxkWf9mLuIwiELfujjP/MmQMfKF3YLNT9B9hcjm8dknTSeWkGUMfV7udrwuWK
9FWw+ov14hLd48Yp3+NOuM9OTrI3H5CJdXDT8pq1xHx60nJ39pZaUHOJLcPOsPqE
QkyhonMqmODBT+SaazPhJfn+q4Zf+2HstahmV6TyW2ewaxviqDVf2+owRMpxcPEr
JuCZriVHW9+wak/taWVNXsry69O9U3q11Exs5SBduIRahO6HUwv1JKQeAKTbwNwS
QDL9pwpBd0NgxSZDFeaKyuWWMBBOgek2dAZg1LGePMTnFcXcjg9R94JMms2Fnw0Q
xCtYAxL97vT/IeWXnkO6f4r5fNUJJ2uZDJd+u9kIrV+96tsX0PcfzCJvnqNhq5DS
CqBTKZWsf9/M19eZ3Um3PPwflH2NEbUj+oMTBhm0QPfBkNcJrWCpvWapQROgi1yV
66WNzkMiahZabCXYwwMhJE4qSUDxvVp0rPJGdyrUndgakWlhrSHQIGLkJmiZeN5Q
1LOs7ERUdJR9WKzVKDgWm38nWZPnvcDJBTuT78OqI+XXLuAXKKzNCa4tnh7kjAec
KE80cYX+7eC0s4nQP/ZkEtoc2ct4vCy0nwGL0ZrUFmAl1U0P6EfyrqKxzmro76xq
zRdkuXRyKDhKrMEfPGpg8ZXLCZ8viM/n+ePONfF8LEfp/C5rSLkl6J2CRxXlvOgy
5BFKQPQvihRwQa2NkewCeHGWFShMADG7Qwp0qXHksM47De4oQWIoseFMqxDE566P
Eal7H3lT+h1uLiy3Ovv63hGRKrBbAPG2sHgwcOXlVqh32vovGOosMcJ/Y++QYQm5
/3dy5LAkLi5hhgHZ+7XmqJDbUfK48BKUBi0wOMgpZM3bPiEg61UUS5wjBKcV5nUx
EyLsax/7lCSFKtRuZdHHW2fOiuSECWGLEGdVI5FlcmuYUnt4Cesx8R4TzfVNFZ5K
QjLvb6J28XeQrqMYsdNyTWb5XL5bfLutjTN5mRVqRPG4QIpwAz74KIoD0X0VlfJh
c9MiXx1D6xsW6XLisdOVEmQa3qSEDsuef9rJw0qpTalZuUFWNe1yBZiVpUkC0IY3
rkMzzI8PeXiOvx/cr5mSNf3+4ignBMT7K0Ka8rm2yjAoyWTZys97aTI/vmzqp1aU
zeeK867Hkz+qhEB2dtQehwitkz9/7HaOa2iNjdsA96GP7BW2z4I16WJmNUqynwOm
lRFs0aP7yyJuJzBHCBqdym6/usHr1OcMm3NnSJfZ/lEySWYSRT6WT6cq7z2jcTjI
H9UF/xRalRpTa5iAcd/x4zTvPwwDmVqwZkSV85/XWA9bTt+3fAuXJdOc5Kzy7XPj
HqOdK10XqZ8hq9EirAc1w5GEwIb/1BE2xpIEKqAzPlv8/3FcIfKqGWvGKWVsarOW
N9d9j9V2u+kmkIPmZx1oBVfaR2hS44NCPLqFgRo539ioW7C3Ub9BjcMpZioFsfCv
PvrKPdZ0mQXWNRApwu0RlMn06pDJBDfkTxCORvTCU4E7UAfPbSqL0fcPxvK9WxJR
DUEEv/OKL2ix1xUrLSv9Fm+H7rLPDKFnfeXghTjluyYqIQwLUMCpgY1EzT5wu4R3
4B8/cUEGVHVud1SAvg2hH6D0cSAC9j9d/8KKO5+d6qUQ17mtpWCHjSiBJl91kzHS
Iv7DzlsS9XPU96n0WF9mVsPpp0pU8IC1Io2MCNvBp3WX5etemRiFc4iwaCv+339G
ADouZmYZbAQJtzQDna+Pxzlk8c1rXpGDKXSWik6DeXNlwPRaW+2O6BF+lizlayIf
ma6FdWuoSH2/SN0HeJcWJ13xNPJRUTdio3b/rkzexC4oqv4d2Rj7cc4YTl4euW1n
Ovghz8OtGO0PGq8U69lT6SVh7I0cMaItSzzBzAwNUeo9Mb3tSb46daVK6b2RXCDn
5JkO8Rh2Qm+wgLB64XRC5GlRGFeroZbtMGz8Rss1XdJnOVjNcchdBL33TLMzqId1
qf+gdq548dKdVbpRwOVWXBNSDY0Nf1oj8E779GYzVt1KVqAOQSaIGeFSMQIv/+mq
jJexRdfV8nb0oQqSN2k4eXrP8pkjQ6iOslYjCQX5sFvLwkBcdhFCxDST/g68r4X5
yEitn2eTRyaiLMG96jUyVD9iMRPMimNXsCIB2X15Owgb541LwmiMXFAhSn1aPw2q
d6LeZ0XWJmqZ9394mgmsNkfdvpL3E6V/qCFsLtYUG9vUMPTuaagXO5L2sIgjKa5L
WrZ+01erysngP+TqNQ6dy2yiy0HWRq9kZjdit2wPfg7NV4o+vT7BU5+Mv4O4btGR
3Eh577PATyDYdTSNcVWqtJdBip80gB5baArp8035th8amfrihroqAbkrrCHmCEB0
TtUxVl44BD8PabIXkDk9doraFoBPJrZLyCIOFusj1yPDWfgbXd8CkTbLZwCkk95o
5sVUCukhqLqC8J6nX9oEj/lg0uepujW80c92h5EpGdMkRdahTPvEO7HIHzBovLx6
Cu6IzLrWAXQWehMibfIoEaicRf0IJkb7Dh2k19MeUK44Z9NHp4K3JDIsX6EKriLp
Gs5MEu9UEwBzlU2g0p2oavI5/vXcLwXl1vylytEuvwo7uHKDvdHqMpZa3piOWQNs
942vVd3Vr69mKYs34UUTgsjXBWIWBGkhL4ZGXNr2bW6H7rtdyBJYyFyxwVaMOLKs
fmF1sfTtiMtsm1gPnM5GsVtFNTt3vTYai8v4QbPpzU6Z4Z7BNH3IGQ+zgEfOgNka
vrTPybQ4qeYYE76Gsnozh1nDr88HzQ25KpkpIQJbVyJcgbBwWUPbWF5g9fsDSRcN
MGZZCSkt790VEHBaBZV/jgQTJ5XCugDd2SinRKRRTo6sHDlshmYYW+V55WSCPHp4
J5si3x40+oFBP6XFLspibMGo2RZPLFTzo+IisTS2lI8iyob5odGcTGzuFSXRCBSy
kc0GShSyTS/6YyrIZcKN6j2UYEoZUMT7JZUxz/jafJrkuDDVomzWN/poMM7RSbJQ
Ar+N4pN8uqz3xRcnr1uOxZVE/WJrmo7duAcydM33rCVAISAyW0K32gk8cKXqdzbG
RNKQmrB31Xac/wLr9teR5g/0EcIV3eEmCdyizYZNa6rn2Uur2E/s+s1V/kvm2uvN
ZUhLXjcOhcVkYeLdDL4j3uqFmQYZL/sYCtN5TYacV7MM5uhiGz/i6GrfLeB97ta+
IJI8s14fqONEszCPsov90lVuQKk4WvLSBGwVHIJlcEm6VUHO8wOZvNcs6uIajYOp
g2+K8dAOmncOla1CswDVQH9u5DGuOnraFDiUOCBUWvze+bFrX1/4E/GObQl06pCf
4jYDw5TzQVjJw0l9DIDA+UHrdQVvE2SovopYoHJMzq5vbgsAF6BlYyXA+2aESccN
wP4ymRjdp7iS15hj8E8eEC1hbFr+ScjhSRDMWYyfxUyNTR5Rw1lzSlpxNOqnxbyg
0Wh9F9vtBEH02tp8gqgmtVkvhthj7CinHi10aa+YgAIxyWd/nRdK9bhZVMhBDzCY
33EyNrvbfB6GHjWWUj8HJxFpSnqIbG98mwGfgbnDov5NEbt1JbXhrUWE79Bj13LZ
oM8uIvf6amPhyt+Tev334V/aW2kL1fSdtG5OcfxI7LW2pRWmTriyd0Cn+zjRYaBq
o5//R2znGcAxXxFNNZRtN+Oy+Biz0Zbq0Q/uzYelBdkbbqzG+Q+s99izV4kuGjH4
ZUc/HnvV/iskkZPZ0z1tFisv0b/jI3huu6UqEz2JG8zGscdspMwWsjT2UFc/u6xB
G1jJRiU85G33qxWN7LA8TmIrxnRyh+ENjl7ik1ISvjsWpHLbZ6gxSVMVyssgqt14
jIY9oydfm7vCmEADSt7IbeI9NBdKiUb6nDESMsqnRShofGU3GGma4XED0Y+552jh
66NZ8ReUh7QyqP3EF1Ro9YINvxp0my8fiAd2RorAIstXsBLVR3TZ0hKIYg4srzkD
5YjJVQd0Mkp/cprO5P7sFgvPc2U7v9qs29WShn8DQv9m89JsyHrHPchKgjRRt2sh
7lzAtIoDwqq9uASHoN1TUU+MKXugm0nb8XUW1fKosfuc0mMBmcxk5aStHLG6aC+G
Cqx2RrlA/0AzFFothLxhpC4fZxXQli6Z24i0q2TcSCSA4zYzJLk3awS63Zq8R+qk
QptIFBENwhXdAzIov8QiYHctFunhXeEgFH5Pr0DrU0vnNOKtjWmZ6c7xxaGB3heF
vjD7eNZLImxJ6XxUnKemH1Pia0JRzqr1lnQAMrzNwIvlLmeven+dF/YG9LsHB+2J
wm2sB3pu7C4V33v5J0cghvj9Bfm0j9PgXXqrFBI6AyRRArlBwSgKtzcqKOV1av1B
l3HsrmkTCwIjJA41qPLPyGDN/6mGXqsAvGwp5COI1VrSp7fAAGLacurRsUZdHKUV
FTkgOBXD/HoPfBpZbXWdUVGipErs6/9bgSHtB9goZN3cuHUV1M2hZcK1Y5paVDGE
/Sg+iIDnfNfD/jjbCYQoz37g3QXZGeTvIN7STT8H+8uGXXNr0mUiCJYKAmSb/qUR
Z0NWdPZxrmmcgQossS5zqdWc9zIB+nQjHdjXlNPpGhnMQ1IyNdl1fvHjoyI93ZU7
aDtXV9x7ShLF5bWCCYPzlV7ewgHy/kMkayrIs0onYdJQQHrGPV4KloEhKcqfP1+4
G+yylOWiiWxfDDP1tN2y1y/1ghh6a3TV3E+Jp4Wt+XBc4ESOGeWCH8CFMl9J1PV0
zXKpbOa5EPzCt+2nIG+AxhGrGAjBukVg9nhKXG7heSFpyo3fJeLnYs7r3I7jMVo3
+oNFeY1ZNXN3Z1vBs8mQTvwpTfixbryjMD4A/DKV6hGNgP2uJbV9blAeQZ+YAIf6
uMydm8C0tqTnjpKt4L3f1kH/7r5JuWhPXu/1UYafkyu077+tlqxtPEjynHUs5dgy
PqlAD4QyawVBv3lpfBVI0K+9eblNmvRc+vqL+/+0DSJeXWMgDYtDtWx+TPHvLsVa
PM+Pdp1GB+k4P6A3/+RSMk9JsFQtkPKaJ0gPmIi6jvWGObs0rplp77qjDw0B6Otd
tDRBk6Hl1DTwnB/rXMJoqoUC280rrndtfgp88YAGy0nSWej2DtgvVz4EtUESH9lp
uF2zLRFhwShz+MgLqynsODvH8yroMCHD+kB6VlsnNCZR8qvskExCkrFzFNKKcA4C
Q2BNlm5e4O1Q4TePA74varFLSaGelXJ/Oz+MOQL7DXSDKIIq/ad/Y0NtsCduQSvy
9Kcv9YobwLfQ8zrhx9SJ8sdvg5uzx245yT1vJQT6WS1BN2YV07phk/b7Ml3WrkLU
/lsOO9Gns+CeBeXX+HlpmRS6pfaa9QO9cNdwsAmapO69z85tw1FCsSRZrKg5yi2e
Xcnvr9Fq7w7Q0lOj9YoybiB8X76gZwcETJnnvkmp6ynKvIb7cwpTwgQs2Jm8CJAy
afmvJrkBGszjyna5Rtrt6M1m9qEi+KEHPN3luDcKxt7lRxiX2gCKLpK43VOmtC81
pnurt8QI8qMS7regDN1HQZ6oJyvtt3dbEkb1OIzNyz+mIsb65V259zM5ROB2iJsI
IiXgDaPJrkACOR7FZ/ZxZ8pZpwiLb5LaoGhpZO7JNp3p8ThgJ6FB27b4t0+22JOR
S1CPHqIlljz2qmxJrYTH2qeODL1riyXIsf30dyJjv91z3dyzjEYyxphcy7Tk57rm
+wFiGKG7+sXVBJD1yf2jJKItwiHAUXdhKtvLm6wSkxcsHCnL1SZf7KdDDrdyQ2Mb
KE+ZsqNwAk4Dz7B0g1wXhc+Ws7196hRyWbfmRfS5wvS0zrO8P5yy68qpEyGT4mhJ
QXqAESB0yl7HvbkSCgmSp4HcA2RMD/P7DhgrNgbpdZ10Q4B8IpLbviL1UflBxUHA
PP4bzZZFP1L8ywGMWjvINY787MxEVfm6NC51ZyUVT/am/s4rxczHULNcnjh0dzl+
k/KkcFh4bOR5oTHnw6BtET7k/Lwlkr58yBv+/SQObmPRP7dzAApuqTpJGrFyHP5a
1CnxSWRJaLEONYTofqInCgJsJxz7JeJDdtgIWb8VSmU90SG/XqZKqyAYz6X3EXup
imz8HK3/9zp1TUzZlik1fcvoJQlHQ5OgOmjw0pQyQG26zyZvE9PrK0vxNpp5kguw
BvyWt5usNRMh/2DPsuu1W5McHHWnU9AnOp0fJiwR/AsXdAMBg6aVkP+gBKsTDvyc
GTHhlCubiJmCKW1jXaoIrNqmd652w9PDtZics56aCRCIUteV0RvNsiwazokex5Cz
+3HfV2xWcoXY3a94GisW+0FYPsclu4KJAkjOtFQSbBkgJrf5Bu4eokHfFkV+rJFy
7cH/VFrnAiN44G92IUsKBMS/FfOyTJ6/IIPY1YOAov7o8HzSW2Qdpevx7AIh+8+6
vFEBJVamSVdhuM5XSD+YJWB4wyq5CHBwmuQYwDaMJXcl0OZvBxwuAcRGdX4wV5m1
0i/hopu1kmoDxRFOJKBjbQOMg6upVvTXY6Q/ihYzcs1JIntdt0sxTLb2e3rzN0Vb
hm6I49znOMJeIQhj+Nw8QNX+bTx3sLT9EeYcVYDeawytBthm+/cOB1SLKcFWT7XN
rtLXldvr8nKcVBu3+3yxPX47SbcY4F4kUcVdFjkaoJU10ec70xVsn0LG3PITCOrt
OtXn/R4dTf8mDj1E7K4bwVkHf8DUFcObdM1EyB8IM+b0p/K5gauu2HgaJbOHUDWu
F+jL0qdOj2ql6yuW175ZpLe1EVnsow1PdKuZ0p7CzmVAhBnZkW3wIDvDVGiXazQu
vbgAcBcyScVduf/v/Tao4FWb3B+mXhmyX+BckDIKnTMPWMw4af7xYfWp6nRofUqO
fyCtw3SnELrtniNnhTqobRfNS/EkYBXyn5jqjn04HKr1hherp1jcrFUGmcIoA0Hr
mEmT/mnGNnIQL56F4l3hub3Y9urb+RtuSItqp5kRtjX4t0y1QsqsWMkGZ7ckSJ/p
KO6YvfPj3yTVEINUgQwtCx5bIdpsMY5myIU5hDmO3+ABMugKMVSwCZI/9pZKEhmR
2H0OJLcZ4Pz1ZKRlUbBtxoJeMI5PQMRy/WEcImLLF8dRjJ+DJ+4bJufvIrspP5+w
8Rb6WjbYwVw5G4/pLZ2v9lmnD8aLeCPX3qMHUwp0gaMdQL39Zu7o3rQi0Z1g3n3X
/4uOCKXNgf32YdaCeDTIOdqk11snvhp26VR+TJPq+AyUmsOZapbvtAlIzJ/9NyDl
XNgx/xkr8Q1ZHl4oPGuceIF2x2Qd4MSbswW2R1f7gV9oNQhqbkHKWPEJDNA8D7nZ
eIBB0p+1AT/SoHUq5JSzGOEJ6kdYZpJSzz1MwhC68o9tO+R5l7WADg/B61rTXlN/
JfWrkDWPXFkcbcy3q6ncmZ77jsszbQtR8S0ABBefYGz5JmoF6ssLPckiR6emMRPW
iW5wUdqtmqO/2WuOHrzU3Sa20JHM/HotSLvLigCts60JGkteOzwlVbTajOpTEUUX
QEErXXQb0xBMqR7QuRKN9y4RLgShU2aUbNKP8xNyJLtbgmvi9X2bRRbQZRrtouGy
ThCcfNpjYm0oclNjEPx1HVKtWs1V1IjYss6uLaTzEVjR/lTrEZRQj13cjfE/Xvu+
bsamO63NeMqqWCcHdDrAYBT6jBj5qGvJk+LrUSGSGIN++Gqr7nh4jgrrzFVo+Kvq
TPmJpYIakyKZ1o0RIR87bbzIgfW7SDOztG7e+IH5KlkXqauPPujigh3RChHhxeLW
BSYivjcTpGXnRcm98frMGAWK/VvwB231m2RJbAtpo7bGpdBSmnun4w0ecgQMiFfy
8DlkLCN+ZIA5MmHKgTaIyHMWY5LelTEec5cqhH/io+yIkC4YhmUHZH0bhj60B1UQ
xeMr2ZY3q1I+1e/vCfqiV/M8xkumO/BhDzyz7H4cHImbELlP3mOujfzd7QNfolM8
bwk7tvJJ8OkeAXyDbKPoTkeCSRUxTb1PRX6DAE63ON8DZ9dNFidrxNfhlp+zy2/9
349+LRu3C3LdrJAL/cyEu3qbN5tNps1IWoyh0CCIWd0kGP9MIy9wkQhxNimIQdp1
fjptEJS68bLQ2BvG+ThOyMKSm9pH85ozrVMGgD5IVN810BSaMq2wvCeTNONuwYB4
1senrGW8RvvpBjmG2qCWFlcdKXZ7hc92JnAOsgrUZGaYm7ZUIIhmh/u4rE5O+/l2
aXjzQ8Y8j4BllfI2a83MNoA/YeffV2VgO7XdsUj/dVWkW2RsZJZI1Ea6RC5fMpLM
X85rqaUyVuMPwTyZIAasPYXhUNbcdpHgmkSbAgRXsuuV4oz/d8QavStdu9HHVkwK
uHrXHGxLM5gcPpeyi5h4t41VRKbciKytgsoVWZJ+ZS1QQUBCswHpUQso2Zuh8/Rz
80PXUK5pc2GlSm60fVS9kyT8/NBjHU3o5Je/yiWEcY8JNxx4DR9nEV9H98LFXa8t
MTMQrScHKka7WY6Kd0Ep/atKnxHXHKSTQBNpDDKAdlpiJ0Vi5HLEPz9wJ5uSZi1x
28/1Um38NS2zbzYgpMg0WvPCzNhNb/plaAn2l0ie0wf8Yn750k9BG+qNUeG4KQuR
gclg3v7f81Vyvp4Duc5J0fUIJhYrdaCX84+x2EUivUbk0ABKb1JPKDwKb1+vUJCo
eVOYlhgjRVxjCDZydGs2l7wDkT7O3jNc+y/ZE18F5ywUzeZHPgYTrG8WsJf73o1H
WAcFLKmoZn3gc64hVXQFYekmCt9saj1D9lvqPQgN5ku2Ydcl3GvaGZoLjRylWhUb
4oWJInl1kDaFzglk/RlHkfLL6VfxS60JjY8Fvw1wDYSMQ0yk/YVLOUmCLDb+6UZs
7S67+N3/kqkNNL3zMycKZJk7JG6TXdT6Mu/ErI0OPFAvJM5cBUcFPItxJkM1cE6s
Zp47mA4hXSJIwHpTAQynKgnUPoRTo/wv0awcrwcnVUNZxxDfaIZENiFATlGNfyFp
BYJkreLyfUFLQMfw30Dp3DI//wGoDeJeLB9MBTAgz9Jznq2K+axm1pqvV0POsqE7
kCP4L1Ri7cqd1/izXYw3Dn3sCNdL75Gef1Z1otFFx2tVMQEQWuFPpATuKOutYEbq
oZon4Mv5axvoezFNqkvsPAQa8PIcQGhmAM7JunwKLZmJjQYxuzINRd8DFu+lLPO7
kY7TJ2FHjSi+2N8edU9erksT8kEC7Xr0Y7PhHL40tenbtXmlfEFQ4igIiip4hHc9
Wl/PToRDCGFUKBmjm1JKteK56Vk3g7CD+rYCTBjF3ZSr2OsIZzAJJ9D2vYHxeqGt
UrUzxCX6YC3PHORdgGrIE4lZviFCoIdLza8hDAJi3SNH1y/o2enhRvKOiDoNyJka
j+4MjVLE1vPeCgSvaHWxGRkIVZq5o5oYOaYLZxODOTyYqAKAVyP7rfKOJxfNe7XV
oL2Ar3WK6vCI1/unqEs+YPe1uqDtmFL0zToE6SDRD6f8MpyuSKy3UoTjGYSv8nu5
zIMljEftNrEUSt4CWGkjniejYkRhv8phwbDMLtozcxQ0NTEwvKfwavVI0IgVELrE
ISzZ/BKcDi8jFq/KN/cLOS4XXyuZDWNci+so8Qts0fsiLGRc0auxgttSIukdHZj3
vwXSICoWIKy3nAAbqDiKt7MmBEBktfXcGpTYTHwLXSZaH3DI3YJyAMsqDxs3JR6i
XZrzg6GuN80e9oYY9de25cE6js9HNexso1jjG4MaiKlk9HVvZF7y0XHiz+ppV/ld
SHR4DMr8kGnqow02CRJ3WHwDHTY0kr4ByabOzrPtxco1XkspZI07ocP5L7n7ttmW
wb7PpW9IEC7FMSo8N6A9+aW4UAmefxJfHGAIu+/CR/EJzhucZjoPwcbKK2qqOdx6
qGKsTDyyLnBnFRxn2pLCbRnm4mR8oMBmAsrhI7BiEWkfRufZfKfwSipWoZhtKZwS
aQNpNwji7d0hCTa7C30Dx97PZ5MxXALINOXpAWrqTyb8fg12IdptXOhmkIoGQ1CQ
zRwIjuZV/w+QqjkxMXkNJnQR9QHzPaONhjo4KI0+EZBmzYV4zbdaKwQjFTETVssR
vst4F7mIvr58tjkQ9Mo4xO3KRuRZbInrLltn0qOaSELikwJWcK4Y/MhUttbKD58I
lHHfaJbk2BuM5kgX9od/OSJf+FfbeSjToxm2yTOdUru4C9I8dGW9ZhWqag2t/ZyK
91cYiF+F4buN+1ivVTTRJHZk3L9x2i/Oh54VRBBHMyz84WkpWsJ0R26yE10nslyd
iR1X//fdCMP4ii7Rg05JfIo6WCGs/WvLa410pGAUQOnfZJJ9FAeS+R4PIjrPeVXS
9bVzVzcBjcYT+U7TNBJbl9Y9iziDF7q/owG1fAUDIRxJ1aYRyi7RlM2RATvhfkPg
ODeuIYhNjvDqEESPQj/M17Hm37iEJi9H7wAG9z3JhBP/FDDdB5l7oS2Fo1PyzbEl
CWUZBbnEng+Y02D/X7SIWLeCEF4jJ4KNTdNQGIMHx3jWxgzK7IditOUszB+NiTQB
6Yw9amGSQdP6TcnfUt2DZ1sXMQoWg2ZWjL+DsVrzW180TLmck8Nc3tQDYK0ckGUw
37qSnLZoacNK6BzgsKhVP4kJZaJWA3TlauPQRHRvBBN56j3vLZ0IGVSBP7SzrE8t
sRlFDf9xNdKUXzx72qBHuTQO6ymOESaUmbEnEQbVdJmSG9XPdmuulDKNeHTykC8D
tf9/52+vza4ysZbasudnfLZh6M9i9HZzg8xeygjO+HmOfyQeCDwVcdwPW8PciRtI
jKUC5QGv5ZmDEFfjoJcVdCn9K2NtL7oa/3pysKkV+kgE9OwnQuRfxTH37fQH5Rye
UahlHrO9DJ2Yu0sqqal8VfGwgXgAMrYMR8NpG4CQycU2GcHuxUiTL2FfBOD51KWl
XKdV3yMfzP5Gf/SwVcEJYcO7TwkbyKh+bpZ9oZXyyt7ZsW8czVNyesZcSmAkPuiP
iiYgMEIozmabIyXr9vgdV5wBzmNcc6yyKdzZHLyR9+/Agh5rC+d2TtCjTttPVn/W
gHqiWXHbbTddoMa5ilTY3ghKD/y+lJxx9wlsvVYUxEuBPCzqjbEex1Mwh3r8cu4F
FXmb7rsCqKHObsE40MiSGbPSveG/ZPEF89gp0uwhutiZ/+nLnMoePFjRoS2YMKGB
Jprur2ea56ntH6Tafj9eP33otZAoec2ZFLWTIC9jQ1P3jTrDPXaBGnnDpE2Ix/Qh
0+4i0gEuuOMUa0hqWDutk2/QHqXFn4b46xzSI1DF4Bf2otvu2dneUoUZAYemQ/Cl
A4Iro+MO/IRcz7u4HfYMe9y6dCNJb678F50G3jeg3yMEqqOMq239HfGJljzITKT/
3Gj7z42wFAZ2mSOg7k2Wy+vj16zeSQGXeUannedMoVcWOL6PZtweJkrr9fD1AgK/
7QZCKTt3McEbpTfb3L13uLdrWV/Ey/JxGDldSQtK/DDJFEzaAGBN2Ed5VvaPoqOc
x0/PuQr1AZanFmK9omHfIjmjYdbRjqO1R5prGrXWzGL8R50M65KO3cUuu4WEddaZ
P4qWynXxQ3BzGv2OQmU7b6feCR6cv8spk1AE6XtsG7YrGwEttZP0vhHlfp5TFGfa
AY8YkoF8weKR+ZrEvjz4sw+56mgMBVM30TVhEKd2M9rBOfSlPOMEYSSFC8AOP37k
tUblAhpYFN7us7ZoAldN539ICJM4Nqd8e7UUd5qYQSH6cHy1Zct8QkW5CgyErQzb
zE0RF5VbNI42kMiKnVypk8HKsXAkmVT6dDU7xFq8zJ/umD2XbnAtCud1l6Id2jQ5
fKHfQU3MI0T1OZFQr4CL7h86jO4aS/6DIDzY4ed0oeNKvhjUOVJiHvdarq2emJOR
EEKtlVU6QH6QFMkGYRxx0Lpp2Rh6dvp8u4CU/2anBhSdvOSEJQNGihP5C85ZFgap
tKZuvQaHCm2pLgNO9jscRKAdCUs9c+mgl5cFL1o7J7iaIJEkDLRFpeRLwsXRjdKv
B+AriJV/MzQj+eQYzXj0HrPNVDqx2/kM/uyGh8UzKwb9FYmcM4rIfZBniC1aetUU
9Cek2iP3yVpXZ542mPV4QjKmF2Mg8loxFKs2ZQQo3CPiSTA2WKVkN97rViZmc3ox
FRsjfno2Ea+/RfKhXj2n4P9PwsZZyVX96+9mp3vyQStJVWDVwFkl67s2Zvd1HFp/
KZ9KUPN94oJjttl8F/L47ALqCG348eTs143uIHPnNFQCggyxjBNyzjgqzGcIKGiM
xg+4xzBuSft9ZlVqVQeYRf1mwyTPLKJYmOCoip2Dr32xiNfDRNCtPPsq5j9PeHB5
hOZYVCdAjjRK90+yQlot/sWLnhKTVWEL0fXe4Vpt/XC6YGxbuQCiQ+6QULoTGIQQ
ScYoiL4AnpdYt1eLyOXmcLhpj7jLGkue3bUmb3e4MyDxWvfUIxciXSUk9TbyDNYM
VwMI4e3eDYwoqfm8SzxNUVvZuIdV0LUF8rR/+xq7Clg7vuYrWK/JvjW5vQsKsje7
T8hIq4TsYQMkJmDkqjQ61AOHn9WCvvJ/1biFi4eIt0TvBFSTjlI3w9GkYpvbbgqX
AyMX5NfgG1cZsfZa9t3a/hsVVLaC0Y56/v5pjjQ9X8nVXEckdIVn2S2JnA56GU9N
YzcGkafsRqHbuC8jNULS3GbocOmyN9ItPw1i9T5f2SRKxj8iTlA6yMgwHhf3DJ61
0HJ7HnNeTjz0Dqr9EQ9aUslR14fZ1D0vlSq6NzzC4/sdACV231Ww9y2ecXSslyEH
F/wM29Ipig9IwDecnmbZBf3b+Jq6xVdZ2IukVAmfFvnE2ccWi+RgpdZ9Zf04Hf7h
85f2IBqadAKARH/i0ST5Qj3Zf1iY80vO85PtUXMnvwPfOpI6hmh2eREBnRKsUxOJ
TZMN9V3yE87s+2Rzb48IKhhOPblGnImK15HaFjkvPLJ6QuW0shqZoCDKxmebRKwM
jh1rjeKSCcwFCR5FTcfFVhCC5tf/hbJnq/IAKpOI9DGjAvKKpXShas2QAxMFjKaX
R55dKoMd7PkDIcBkJy2LFaY6SVqbE5pK3K79C/xRwEeNWJvOjJtEzx6nxUlj3rGe
NHT6uH/hbOE/7eYd9FWFhNZTEMIfYDXCa4JBNaxY9+DG52Poz52Zl9Vrhlv/0C4j
F7n81BK/LSv+I6K0S2jTFgnmSWebKiPKAjaXo+DStKjxSGUTDXypG/RnlhL3Pxs8
2dEKfXzEAH0kLqiAnRLtaAW0cy1VUEwMtI9aJATwePhYpwny0wG5TQNHHH2GP6rk
6zgURFxkgRY9NISNHsJORNW2GyJP7bLQh9u0UgTJ2Tq8zdOcyGMAZUUnjp0tY64M
YAbE58FqyA8qw/kOCRnxUTD8HEpCVTsvlapZ51RZetDdcj1MEwebL+ZLdrNCtdTm
3DqEBq0qWkMbIqlfYDXfE3a72K7aNGOsYv6ewsn4PgiNVKZtVatoET44aczDRy81
mNx5xtrdY8aJHhis3Hx9pu9g0CwqMpA3ZnXkyIy/DMiqrvXU7cxTuGARB6cABmGr
kNlZm2TFLgDeRpN/hvfBkH41qiGhclxM4MHkYg/2r87/ktYaC61l1+Z3ksjQK8v0
coWgtyU7QWUzWYOqKmuBOHIJjYUZLFy81i1JzwgQObH2SWSJ1a0juxHSMDCrQC4n
b3AABOxAdsCoHirjVvsgHZ4DDGIcXtWrMg/LOMkQ4oG7ftfyy5a5bs/Ml1PDTQOT
E3bBl8WKDEm/Q38UlNAdyFZ7MLNecFVNNP417x4pn6DAe5rl5v5ktp0zUsgK49t2
Trr530gn3b7k2ZlvS0biGa7E3ZtJT73UyuMtnkdbMpYXrNQiAe4uz/7WHKAnxRXH
k1JEjnwgf6Rn2eVCrQSqvDSbxOq9SQc/AxTOGluqvPfqWQKaS8U58hsKVEssbHib
bgWgCbSj1CvI41NuLT8WSOb2VwCQgdOYsjmHe3HIslZgHV8GvevmmxtvdDo0ulFU
A+F8O3Xr5mOvTXwDjO9EZqreHwPJQpWgNUCLhXz94w1P2Jvt3RYarxUvuNQ6P3sQ
C8y09MjBCRVUQ0JDdfuEIs68vnAfPLgVo7hySmSYE/jkh0riEJ/6cw/45t+d/MgC
JXdTclckpYQFgdCzxovGAIy5cH61c2DrF2FWpYDWQaojWYHJ+XbqtVIc6rhuGNae
ijLH37ScjCuIghsv5eqBvsFkgKx2rFbtkuuh8SuRsVtcTe4h67GNUBYvMA4/W9Ub
u6jt+qeYzGNot8yJH9tqnfY9Hxf3k18ElkC6VtX5mlIj/wknqfzbE5gMZqzx17JG
1uZ+JiWnftwv61n91jDoBFXkmY02EFqKaH6jwkTYHcUusqFy3M1trzRZZTL18OtL
eyVIZm6DKIi/fRWvjdZNsu0gaASHvhK6Bo0PnUzv+K1NUyOCYJQYIonHJI0kOOHR
V6USIpVdJVv2QgOsxSX8Ws1yJDc/Mgmxzgc9E30rDcCI8Ztt7unNiRYnLlpOFt9h
OrEt4pUP6oSggaweU6goQ5LiiqXZQ0CGET1dStE9oun6epwo/1caLX6Y1MPqth4V
RWrwq1k64Qi/LXCCuSkv3EpuYi8injRfrdzLN5dJe9zyWBO+ht3a5Z4m3WcurIdX
1Q9HlV3PmyvmE5n0ECYjJcRsgyuN6YaarqDCUHtUT4+iX54z7o1h8tiu7n3TrEFZ
gT71nzViha440OJ1gIrYmUcd4nXjYXf1wc3jq58q+sYb/O8kDK4KxmJbuOLlhPhi
KDskb0zGxaSUJc5R8m9VZgnEN91sdWlpvMr0ApzCvXj6ftcxqClUYMOwFx+98tKu
7xfk6PhLy2I9UszmnbpD6roo6cgPv4zQs1Pzdv8xA3vnwaZFlYW+r/3NvnIKzKiT
iz9qpLMEtm8gjzAvwxv6MxZCfg2RrkxA7ikL285SebipJZF3qmfvNEaNBSJthitQ
uQ8AB9t6t7QfUJiNyMTeacypj8mhUrVH/1VA9H29nOTVJcCvk6gEJn4JZH11vd2B
8KvgksZhgUPJAEWqI9mHCAItJ4JemXn7wjC3HOdXxvpb6hsrXNrA4xJnivdtQ4j+
TmYVw/h2ZHX9BWQpgfBWGj7KLUr/B+dgA21O/3jiWA8lZr/ZL7WsnXmRo7s5gSI4
ZCARWdK1dPbC0HhMfYfW3qG4LDk9OFeDWE+Ni2PhKV9wM6tCedHgyfA9izgt/nZ3
vAj3KhQvuTM0is6MTc0NmDViKXjF1qbD7H6R1shS3RJI+/NtcGy6ISpR9wwS5gdr
2VLktxgzmA92t/pWpAZhfFTQQeZMzgHslKf4R/uNJZ6FsbGdxQ1meESTE/j73Eot
0NElrw6sPAbtvEpT8EFPRutWgnfuAj0FTXWpevcWWTI+RoEKyno39tBInjFeeXlp
5epWv6/YePY15/7SYkxJOvKS8+IiHH+Gc9zaHKtfwBXBYwxX9/zn6Xp/U3VUvt39
wnjsPolLUX2Qdygjh4NZmW6Ae7JG2STejcotPKmPDBp2pHuwOmAg1U+hHhYOrb6M
Bd3UIcRpcZ2lzZPfBkc1OO8X0+BN4ag2ztKyHgPV4/BUZ7HrBpd22jOaNJG7tUM3
rAIb3eWXQU4QSU8P15Xf0ghTKbqpqALYfkJklN6iYWpnobm1KdN5h/h1zADYqGwM
UVaeN51aGoJ0aOPt0akoQlgp7z631imh+H6aHmiqgVNshpio6l/m7c38iOdzn9RM
mb/kwUx2JKesWK+MElt/pAFMfPseEEWMJoyBRBueWH3t5yLvUdr9iFl6mDaYYr41
5CpGB4G0ehPNDlzMQ+B0VwQ2tkjs8Pgj5mR+v+oLkhveXrz/XF83imdMo+hD15cG
7HM34nzbyUvGKZb45PbXKgSO5dajg+MAQhnu1F1hI2uDsKa+n4k2T5Kwzl1g4UXc
C6AomrB+7ZzsOYZCTcKTajHqWfODXApJObQmpGijlO0AOtVDz5QXvuem3W3XwqgL
iXfNO0aWGwiu+Stn/3vH2+rOOz08jyW0LWLx0npc16E2WL9hxPLboJcVkxLcFKm0
ZF0MCjVQmf5D+jAXw9YjQvgF3mUg81nj4XS117lRDDaiLwXb+tDAnInBGYnk5wH/
GzQ81GZroznvQ1UQQu+WW6yY2M0cwKCUX99ZUx0BxRBA/aLExqh+xZJPDRF7ufI4
QWY+ZNgpPbkAyLb9LVweIemt01KZJm7WaD5tZIwK7ICICtX6fc+PdWG/fwFQKrKU
e55ngfNNmmYPWhC1ZxS4zqwrK+czFCpAFCRpB6WhDCIPHbq+GDl+Lql+AwomzCxI
HOF9JD1rWlxodWp3jfOqkNjOojf2j702YdMBhtsd9vD63Ayh/Bezu31Xnox8jAfR
s1BocVCA3pCh91SSXsNZir0eaK0H2O3p+gsoL6y9m2SZlngp2YkjBABWn3FwzoA/
uHfgwrA/UnQVtygH91Kg07yJRa2O3AKErdh2/jqnJOIxHj4IF4Gipr06otW4ztL1
lQdH0Zk6XmaFxCoPEs1UKof88r2DMbfvc+/ztS8PAHeg+5mrYi3W2QrsADwiiRum
UyYeOlm3o37ZkPLwUhOn1/xd2ihMk96AWD44b5AqtfJT7+yALVYh+FwCr1aen8pz
EaTykhO0SWy0Ibv1NjpMMuHBZj3yqmyHMfEHwmebx9t5oTGCh/r0XblPaoy45m8b
lscukX1DRe4K4dhDkeEh4jThc+3UlitAQaVzWltEvY0RVHzdQPJG+4f46SWRMeqz
497Ll/7uvBKs2SMlgCG/oaHmRtj/ccxBuSkMf6a5HtuN9ShwCqcccFr3JMuaxruq
ubLe0RCsxTcPeV+AsRSB/AY0H43oDjdf80sXSEMPZ4cJg3F2kzKcQRieSV+QD9DZ
xMXt9umDj+pFYvLd0ibrUcF7Tq8J+T3VqXbDQ10eXmLgL4Hz47Qt62eY3SaJtnkI
kMLqRkz8lm3Ome8e+q6hR1pvbrPWxCTVZxXy2t0As31xNxJunWiubSiYWakZqF7n
/S6qyNo6vE1cDTTCU7tOxotE+k1lEChYMfoFgDOER37rJC0tVo2TZASPH6obhfGR
rmia9xClUzDFsn7qbt2kek7ElMEiG/+e7vo+Fdj2Z0J/MHpjnT419R2P1FIOf3NE
oW9PPVdAYwK6nV9feyBXver++I44fC0sKYM/0pwVtdsZC2oKJmcZhYXxXnZ/Rf9R
j5aGwfBjnLXSLOQPbw1utJvxL2GnV4+bqSe7RyZrhAPnqDjaV6BhcKIUqGy8vvCe
dpP4HF4vRD0sTBFvaqc//340j/2OipHa9AIl/PBiFXQ+PL0Q0ofRPFFTY7EFOlgV
wu7XA2s1ZTI9mfHxEZRAYWsre65o68dUXchLNwSNjMJc2o4abmMKAOa2AMXbeBr9
j9ZNwN7eg5XJghQYTzF2UqZ+h5RAXn5cQAIi5txhqP0UauRgVuN7S4qH+HbWqOgu
ARlt6jOUUB4JJ5yGrjz9axzJTkwftN12DpNmqe6UaulnlzElrD3ZNvC7O10d+/qD
xJgBFp6vgjs6CuAA0OCu4O9te4dh2MfnhI3wjL1jXvEQdcy9TCB0lLDuJy6/DbEm
TzKfw089HXcbOZ13xOQxwguQmhSAizhQJAIvJ1elOZnECJztMk9QmeVr2gu5KSTi
S00/VniR3MPaq0rrIkXyrRdLKKkEsoD29RFAt22bTMGjdvr+JbZNSfRElJYY4sKn
MDrxAiSqCbTYvDhGZbK8Ax9JpyR1FUv/+fzjK6U4OWAC5h/Lvms+xOpkXLCFBpNH
Qr+CIw/dn4tEAdWWqcHQIbeFyzBOaDR2RALCsdsUTTnV8lbkTwAKbfgVK92Q9q7P
9JD6U38HP0THZ7UcR2OacI3MdZkGFhncOkmZ8SZVmXbW0O4KORfxaJCGe+/Qduqi
269K1bJsm+oDW1PUpAD+3SVY4GmsI1BdHOEvcr2JIYra3pQx6MOk5VQyV91G+HPL
Ds0Q984OwaocCn1mHOTmI6bx7a6XldvOmQXOvrtxyo36PRpYrE0Yk0CYLfmdtgq4
9mwfA6jfJPPqWoB5dHB1JBpfMBiMfnyL2NSrhp3lF0oMQwBV6TFCJe6cI4prozPz
DG6K8UZQCmDc0H1bwxnq9zF6xLagU0O3Sy9fLu+9F+4hx+zyLDbd1/esHgxPRI2K
2BVZa7WUya57Ohcqd0G6J+QXcvaFxOVSH8Gc2skdMIfi5GFa/2b+/g3GkgQ0e9si
l/dh8E52mEJhWPDvyHi0Qrq/tYLz9aThKTvVE4Xee7jnPp3rRe2ABpZwWpu0i6Ix
zVxVu8bNhmGjIm8BH9Ubh7oXhhD37YTyOVtPaJE89Lf26kto5JztInfEYNsPFLOG
TUJpeCZIgO/rp8kyNSzmMiM/nPtENFP/lBmMnZknlWEU+bHyjLmHNovq3CPpaN75
WWDzfXrWha88f3F/Ma7sFMe9i6bFVVIqySsbgI+FRyYrGDzg8x39yVQGcb2FYUtv
j43UUVD96ejPVKA6gE/8wC7+3SDTfMPDS6N+m6ulEkjfVkQmevRSD2UEgU2sOKYC
jMnPKvqIpMrpTgdFWcGnFMUQ1YBixNRdzmPKn/QG+55wlQkvhe93akUsnbuBwX1r
R5iLB3PEEaYDDtgtjATahsN3tCDaWIUDoHf3q3z5buAikI8OUbLFy/kLVlAljw4w
zmWOgvIdn3NxAsBJdRjJo70iTxB2hl8Bv/kq8rg2adWWkq5H+8DMKltVuJXgjddW
qdVHLjDlbEnBwxmThivVxJRrT8OXgBO3lz6PCy7p2a9OYtaEsFAWtf0GWUd9vdlJ
zYirNRn0shFx12Z1eE2GJh0UZWDvWjpSzWgY9InMXLr8pdlDJ/At9HNUj93Ze7EW
2STc3Ue1jWTDrRRb0Bgv3QlN+/U6ZNX9J4gfYAozyVDVQr95cehR04unvEWlqr9b
1iL0Jk+pDKn4ORhEfWTF5ALAD8c0iIr5cH1FbVVAgErxkl+SF3f7K8UdqtmNvuLU
n0xms2thtUaOi4ByWvXMMc3zU/tk2Cf5vSCzblyKFhl2tnq9GSzIJY+2NS+qLssk
v/k1ee9nR/d8Ob5/uMkcJvJgNX+H0BqR7sae4Dj7GxoG3Fv/tZXhJE3r56L/Q2Nz
axLU0bL9E5f/lTonPz0O3951XhmTPNLeO+tRvwyWf1q0hRkROfSg+zZrrullVuCx
fR8V9O1fkdEURyPnzxrVJYSi/io72cvcBYa0m1XDD1v7aLrU/rHdqRXjdZAgxohv
yJMVnu2+3IOF4zgcSIJm8HNydC/XS4UaqZFmKBaKdTugOhTWDMJVdw7kAktN08Uk
65VVCaSuFzTxjgILzcMpgoCApuoWUanVq9Q/OwX4ccIrvRRhY/QSnwwPGPbO15aw
coxbkaigahO4GDjbys2HtLvOb/RItt+trKacvbr8Pt9FqlPKrgMo3ypSAmd0k8Tp
sN/qL5Kfrpl9ibCipr9HY8HaPAReGq3Kx4nlnfxlOp/pxd+uooDIs080DnFhYbg3
J5kkRKal5+Oy0945UKYXEhNzE1FJ41ujKdgnNO/Uh3uK/fI54XSEjAeSdwYRDsaL
DFpV6DKuFzUpIC8EYjSfYxHdkAqGNTKMPjzXSiXaCC8xSh/XO257ELt4Olkm7h0g
Qzyi/VUQn3RzosseymEFnzh0UuZ/Gy0Dd6qkgWUT8xHko0/bdBrW+GBDqCwo5GoK
legPqBhqA3y/Z2/bCDsRNUtTXHAm229Fz3vRX/S97v+HFw1UFsczQzXxXf0yvK9e
/6pGF5aLOtNcBSjyQ4mlWUIATqrxNW3vpyXvoRanRFNhzR8n1lswHBaxLBr1FM5V
iuZY4JqlRT9TTVoex+napTaKO5GUa2oFaB5D7Emk6ed+nfjgJNLqczIeU5ZPPjPJ
31Vh77xGhSIsiVvXPU0/SUXxz8L75Vivw8WjtDtNdDnvBhB7uWnRA8ZHct0ufwdW
NJWUTNpLSch60eyuxNYS3VhyniuvE7bN8+bfk/5n54/ClBY90s42r96/63O+aqoD
UffC1+KsEXB3QOO/FPQZjcYHUWi8SkpuS01VHZCzob4EqQWzOGSlLiNO4bGPtJMw
ri7vFQWhyAR52GiTR1TOcInsMJ4qIqYdPb0aGUAZVaU0GSq6aM0UAmARmnVutLKE
mb+FahnKOBa6J2CwWufUKocLqOiWYZAN+ztVVvPMr5Hvvs84RoLROcU1vO1kvyCn
2w5MXFPTIYORw5NUWsX977eR17l31GAui+Hk4ZMjq4f6wY74yJ1i7e+5KAJ3+xyf
ds3GQCeJWKw10qKP7MCK69E3C0zEC73glR8EXOUDg/p0ZWso/ULenpr45tKSZUSa
qpsfFK7E2WVWodsCnKijF/2v8TNZUAkjryWuMFC4LvOeHAl+VaF6I3ig7M09cLYa
4P56aFXyj95liDq9807fs7zRKBjZneFPwTzQ6A4+wzoCMZ+S1V5VARFIJzXkzvKT
JdX7KfSCLeUvHr775CoEhFCMff454pW5+ZiOhxmpQ0FqJCMy6XJBPGjx+XGOegXY
8Mq7J49iwrx3h+TcR4FfkvygV48JpHBcjmtSMkdiMhu2aT/zUPThFlxlI69/Q+zk
IHPrBAwUgb07inmgIRq1crTup7rkePOZ88YSqdCU/cYHr9WOhUfwbqRqxjtJ/0q4
3hcWJw/ZCB4BISXijVFypW+lhfnoP+RFOWjeSgUQSG/fjlwMYu/bn1tb/A01NYo6
rw2xJhpT4u9oo6wrwULInQUA7cVmjJD1lPN2Dx9CI5DyS/x1xnkV6qM+zc/xupoz
z9EUoXTu4A2x5xdNQIcw2+t6OodMSG4w5cX3ytbpRitVsLZQMk+gQB4KcVLu7xci
qq8gggrO48gSNa4dUTcsXYMx3PP422JQfFXE3M5Ilavu6Xh8CVgh7Vdl5jnGTrcK
2JUmz3iXnB7pAZ3IVlCZtX3W3qXvMxBlyGI55YHte2SIsQvcCl6kZGW9aFkqAPmW
kz8qi3CgBJKo+ev3rIMVgIqIFvlwD5A+7MbwMYymALE6OV+Lj8ZKu0XgVnTdseGe
VF5NGhR0PEwuWawkCtisOpk6+pVcKidsXJ4ZwfSI7RWCvkss0CtIJf3+BMJQcMup
7mThTWahQzoxsMFHAV5LRqosU4a3a2VpCWjo4znhRpZaLsCSlg9u+LAb4tLaYhOR
lqm4MRqVIxaUJ4yuOZVIlS0Jg+G+ztNMdejJOR3o0HmKx9+nzR5A/A1aF0XYSaKv
ooThRN9eddA87BEv3hPxQfjA/7tzP/LtWIu9yLWmHX4PtNa7Emxtrq0nxZb1iFB0
hS5WaFXcs3SNNJOkf8YpZ55CLQhzuBE+vqQ5N1MjX8xQ8TCzpzXiaXWeyxYXabCG
jmo7Ad/3osoSPgTRgZUWuoROlf6zZh+jvnVMsSZP2EzJPbI8SAE9uL4U6SlSdw85
MTxFE3MBm0b0C0dr6YnHg1xWWaZDLkYl1U9cLAu69AQ0SljT4c1BwGTNrFjD8OHY
VPwnjSvml2hSgyAqgVN9lqJ2lfg7P9QhMvgwhjWhAVqDHBdNakqV0gU6moJ2/IYf
U4Boxrjxpf5pt28P6SLP6MdGk/7xGpyUs+wp7leMcMEkhraBH/+t0VXBd1U0vYbJ
Foedabpnfh1BXmN2ra6KCjme2jJHsyeei+73vHB9GoabKoLwVNlJMR3q6PPuN7oj
rR/y4g+bgDnX5slB7eSjlAH/d15+hu54wxvzisucnBrvEtb9v7BVLPQvV66ucikw
6kfaHtpqsffICX/jTtwVhn3YuqrVFAgeVLCWEnxqhS4AXQZxUBvaPv+4vIgL2gLI
6hLLajAzmyzxW514DZF2dDBaQ5/i9r4fR6WoYFnUYcZ9XUAP7cdRs1N0mUBlfbCe
2RoL+UKixS1bgu+XKb6A95B3adOHUopC77rrxWGR2FLcr3rrJUxD4L6L4rRqIUvb
O463EcM40N6I2QjrkrTO/GdNSRTkI61gqFvUFFTDVChJRm8NLsv6QfncRnzPB+Cv
sEeqPL8tZOc6IO7SiB01lyXJQrB6LTopyNUAy21f77NsY/zPsb7CtvgYj+gX3IXR
jDGupcIw8Zl0KCi45elrg+8tGXDoGB5CUVi/C5zX3GXKpxs1FDhSnUM5kKGFFMlu
T4ohfsBG8euZcobwN0HjRx3wKx6Ff9mP6EbE8HbpGzHe/Bp6mnhYpcWuVloIoLRQ
l/kAoEWL6kF5HJc9UbIPnouq8bSlHg+2/UKMBhrvxC5gZawRu6BamPun6WBeQ/Wp
dqUhfTtHboKwX4XOVKAJbPLsPBHyrFqE6SMTooiqo/Cft68IRX7t3jDp758NyPJy
Kwq0hasliB+6X1GH5QR1YU2+AlVks265qkiQSy/Y0XZsvW05Rd5UhTAZ57+MdzSj
rrp7E/7+9wiva+7eq/jN5eUaP38x0+MBxA6dxcl0zg0yHy0r8Zh/GqWJ22eXZfbG
FVTRljtIccGJXRJqrlQWu7madw16IbOs6YpUY8PfHwZ7HoBzLLE5vtyrXrWIdkfP
PrYMQ8v28OsfUzlmHDWFsPmipEDnxcxV6kzWXEMMU4cPwDnPanDcbwzVJZMK8Uk8
nIEa3/BpRGM6g7VRyDzWThk7jgQ9UKEv7iFuHv7EyJaGYAMYkqpLlACpK1zGg2Od
tJJt8UGdOvEjMO6vmurs+G8myRJtEP43N2k2hiaJZNb7Kht3lOGeOjW1YwhnnNyq
kQ4x7yGwCIaeST7TucgUdJET/sc3RitK+Dt/Zn6eStyMHQLUILxQGvSYz7Pags+Q
2YtbKUnaef4ydHJI3gHE+gW6rR/n2JHXHiXpL8UkhWGdhaQpJXiVNMc8hAymjpiA
BET/mYuGr4EaFA5Fus5O5cZ+AXkrd8zD2m2698bSH1VRe+SsOgfABrg3fNPzab9s
vYV+zv21OxBKfTmH9TRrn4xpeTc5596auc9HjWDEhFOVT/nO4EQq4WtDCCw62S/4
Zq9VPBsE0wFLcdWEr/GUnT+PIXGEhdtGLFRRzh1+XIheKMWyjvd1edYfjhEyLrjI
8ilStl4QZhF3S9MvUYcgEx8/6lxDc5hGdRlVkt4jesQRDlgvYburuITp6vtLOS8N
wBvcdgMwX2+sUk1vG8Rtg1fjfgxMxg6bcYo7/5Z8fL73AcjtchvADhOmcOZprkUo
haMovoYjgjCU3upNIlEdrVMtN1A3wz4A0NnRoBLZh7Ay34IJE1+kH1hPYa5hTMtf
BwrHzOQ+YXAXuqcPWg31DIxr0UJwgCk3DeR1PSA/3pMFokiNnL/vHc+msNNUCDWe
kCa77T1z4REz8xy6QXo+CiT6jCpU/dj5Es9aZWRytjUyzRXYgfeOb5gMion7KlVw
0cRNFVB85p4Ge+Y/CNt/TLuUxBs3EjLOYGJOTXGYYXVFm63RamKCJHKY8PXlSbhy
4BXo6VXEWbgxMKD/VNinKCYBFhwTbga4yDblA6jPqGZ3C1WvucSa7BpCgsVKZ3uu
3xNaFBeSEyn+VaEOERqfUfc+qFagdM+T+LFfhKvdHLqxrZGIjkjUZnulKkun4GsA
EYwltD9zWgEI1qCBFRDl9QwIDCfP8K5UxZYg567MYfA8UEavqWOWZM6wTm6xrq4w
D87XtK0oxbRwGz+wG+CFtX7YIXBOqKZxy0fqe2EDkTlz1TsyXZmHlk0XvfyJFxpD
o5WevPn6uuVmN2auvpqK9LoqEKoOXB8oHXanHxadK83/hnp0UooeEerOlXCPstsw
IFLur3OL1A2QwymNkxeZUIYNC2B/GWql81VglUfgV/xA33RMmTj+VRaXOCu38CF5
6rMIn0uGYesmIkF0lanpRjxjlo9eHtIM0uKAx6Blj+p0C1cp+eG48rruRL9Dy6T1
5ENKEfEHgJxhQc7oWHLdWmU+r1DCvlOmPwVH+hqS4l1OevAhzE0CoXmQnav8/xK1
pXfmacxvJfinQmHefuUIUT4PICgKwoLMcp8B4Qll3y4+IqnQvJedPmtMHLaRdnGJ
nmI0E78x51bJRsveg6tKJpXWObJ+15OE3EDu2Tpb+htl469goBNOxy2Prq/VwF1J
4w2vZxwKU7ELSkZyc4bZ+xUkz0+1Q4Wp7MXxA2PHI9BDH6V6x/8KABPqXmqjQNZf
NL7N27QCEL7TUjAHzpUbL0b+tluDuTmJkGkwP1Z6Dqpn6w0v6PrmLc18xukNygri
MJi02teLQ4YrcM/Vub91HQK9MXDh/uAMxoPUlmjZ6jrvMjOQiuiLRG9/QFZm4Qe0
q2FYOn8htCgZzzQJBYR8+DllMGsEam/nIx9rSrbzNMC0R+cYpbSnUlv9sxvrScYG
TjP16ibBCiqQYr88nPeMLQ/JuJOM1uv/S/mn5Mj3A3Zz6Dxr0ZW3Awme78VVApvA
1xaPzV90K6JSxWMkfMZJPQFh3/sbhyIekSsJVcyx2NVIoDi/n5tePo2BWdN1w4dO
Chk0IJb2wunpF6WxNKfBhKV4HLuWp29ZVvOoh/95+AkxYrOo8Ji4ck+KrqUy4oRO
gLab/pJu0z7XA4RfWHwo4Hj+rUc18Dzez9RMnTYSf4ZMQUUrlNUlit4i5bhzfaao
ECZK1lfKkpd+ZE1OkMsjgzsyekuXD+pI7Dy9ioRhDSI5nhkMWT00xWV+a8HGeQsD
Sld9adIZ/Q24ekqvHSwUeBJPi/EFK74GsGOvi8HpXBUisOGVLc4yQR/JlxsrUzgs
2iABFZRInM/VwmBiYwN3syDihr5bdESrvtcGTCb6Ma4gybw62QPYNeYqNfIZnISa
99mPcK06VKZ9cwbjIVmDMdFJjqqqD8nu81ecvM1qrZU4ffRAGNtA/blQ6OCvccbh
LpWkaWcP0KzbfHjUdKvuFS1WcvxkJsVIc0i+uO6Ec678uviTBpYhGbeudJjLdCrX
u/eBz7t7dA6ZCVxFecce/5gY8ltrgA/yxVkj8KOUA4eHaIbRhteZXcMYJKe3Rv1A
QrIdvsTJ9r1YW6alp07/TkbgYBkcleFIV3Gnb9zc70wGwYc726w57Xdobf55Ica/
HAY/DtwjVSt3AzU8sjwFMpw+A/UFT1afCacAJd0L/Kn438BLsGfHgl3LWPcRTiHx
6ZhGP+pOAeLUT6xbeFXCqFq/rj1tQt2XVwjcjKmRu7OY4nG+fzRKcX1uZoJOTX74
bZpgEBjU/YF0yJC+P7YEbhl04dbqVpluPirrLKQAyAn3A9IF6lElQ/vdLVxhiTGV
oOn/nFYKqBXfFeMoKighjmvnP8a9Zb34b3CY/51FcavB5gA3xoPsSbwSX4z3vPPL
bZ/siE4JMh5WXinjq5ARFS9mgsuIuieuPghsnEWbbWvzITSd5/9lg5yTsaMikOn3
41cORPzFN9r94rS+OiC+NCI+YgPHtBaRsPdh+xrmRELkuG7fI1tuM2FJbC9+l0W6
asLDtn4PH1s8KiK1Rlsu303RnG2N7WZ3QFeIdlezzl7uiqBsx6hD5YOiDAs1pNaI
ILgCFHyy5b1F9Ic32pI3SZUSilvyyuEg0R8HDZSaMyFu77ew0n7KCaZoG7hqKRyj
GPIcMPvHtXQK7Y0xE1ysIPTB18GZL7uIdt5gZ5ftbExGBjahJkmjL3OZueGXWxuO
k+9PRrDR7c/ShS6icKlkD6eIXqCAlTi42SABtrRcP/HjdDdVNCQZhNjMcD4QkJeb
3+F6XkJBI3lSoStwQ1woyDdMp3lhcdX9Tl7iutu/E3Tj+NJbQlaq8a4MqR2L1Smg
KjW8S17IUS2cMzaPbIlZw1lsoOKasakx97pTeFUWuHDqWiBjSYNbTvnKDse+pva6
Po94kySuhMkfBRDC/7pbukt0UZnKCx4z68aIEVz5KWzH/5fclhasFK49vHOy1Hbd
sVy1uXENknORmVTKbrR7rOudT94Y0328+SIhb/CmV6oLheMr8U79gDoCkewVHyRO
eyoj0hfsuUDIdidHLKeydBJOMeBqekUa62QR71VqPh8GDwV19ZcPZ8ADifIykNos
2tk6CW7IGCLb7SyyZi1xPVn3hpkHonM9yMAvOQOyt1LU2oexILgRcdjYmSR1PEZB
FCvGDU6OzqmZyZZmn2lD67CX5KeHuObUYmWorSmHheScr4sq8/dgyJmM80wlessy
hQewKyw4edzjNXFwh+SzHpQ4DC52dMiQ5FzlSApKQDzT3v8MVbprd+F0g5AuCAFF
f6sfvnh6QsSC5tdudi1jnkrxutfokOjnJt/FbrYByiKMilXjM+BOJxnsO6EhJig/
uApuYVbXazYwDfUBRfWsHNl3PJ+E8KNzHD09yDsfg39QNPikPG8zkWYv8PHcXQ4F
J0cmVPjuwzllWe+DmpMF8Lh3YfymEGKhoVLphMM9SBCbQrElrFeMxXMNw4HFpRUK
UpAIQf7lgM3OAiRmwJCB/6cPKe180H/V/SqnVXSOfe08xREL/IdBL2J8wV7zaqgX
oQAHc3Xjhtf3VyqMXANtsPCVpzy3jiahc0huQTCtVjZUycGrZ6+SFb6InMcHm3vd
IODZl2bSk7sYMUJRazG08gU7goZPrDfLzGN6lQx5EJIVzir5dSECs1flqzgqPm8A
2jkX9qvBcSBwxLfxlAOeKaaftPu7e2dx6waB5HD3DxdCt1p2xQoFi5lfvYLSrAk9
PcEkso7DBghm5+XAD/hilODzCabXYcPAF5upzy1vgrCscLa3k1V0T+2A2QgUY2rG
b9wESbbcyiyFMZKn+vwvexd/JoCXSnjuGB2GY0GqFNyd5eMxMu2A5GTceaOERfBy
VYk6g1uq28bT9GTzJouElRM9RinPSOxi2uoNEz4Ii8BuFozyNRYlMW6h3CU4xhrf
m7+/crYR2IUwSlZkpM/M0v3Wwp4tsgR6W6a/m+K+2rS8xQFsmNs/3y4Vz75mABtD
hQ/vkdWD7G5cVJEnvi7dhBsEHPczJHFfm0MtiL3MJCinoMl+on0BR08GDcaTZs5V
3FQk32VTFxmycQJxHl0uQGtdShCPCA8PaqZ+jboyurGfOM/A7zVrak+9oiSemEpR
cwTj3VA+nXCBWQuzMevm/Pj6cp9mnTVVaxERgb9Rf3DTvFDOyqAvv5UF+BhpJn4A
PDcu42xuUTlvYq1KAgNADDB6Rbs7ZSxEIBL8Nld8UfLi/gWCjXqbW8GBTIZVKHqg
XJT4rDpqoVc2CuEODSL9EivdTHuD1QC9N+P7PpHR6rUG/hiHPjLiguTF/jHZJn4E
4tTX4AUlV0EtDtUx0qsh1V+2t9ORCiH6S6NcXkn2T42C6mf/k0AsQrbR4KBzf3+/
CbmJYyrCM3jzFUPKCsifHosKej3A2YuK26XOHS+bTf0xKlS0iOufHCRS6mFy+eGR
Sj48TuMpVUoAvr+6bLO97xFl66qhWoOrwygbw3cwE13ibDXe2XFoqm8ufTrGUBEG
He4Urqp5SfbYrRYOAlNcU3q1nYf+WyluUOgaWjgeJIzk/La6H7/1W+WPilABhkF9
PKHMAOiqMlhDlATnYUGjochGaqi/w+MNqAgWZdkXvzXk0uw+qB3s5zwarrYsflYP
OFAG4HgST5x1+zkyCmX1Ub2AZ5uJTp9ardzyZLaPCU36nmI3RVfagxPggds8PjE6
dPWW9bO4NEcjkXIcqM+Ajz5VrJVfVP2MY8vf7I1oo8NcqpX6TkLBRBA3nFvYZBOZ
UkGI7NO9rq852302evJDPgBqefhNyW5jiVimndQmm76a04l/vkF+HXJGZeQnZzIQ
efIQeSMOX0OKI9ctMQQ1AFhr4JUHtbzUD5hpICO1YnoSSDj3zDTwB2SNsmiuLmvR
Ol+ajDLhUc8K0pZnMTntyGJNlCZPXG/lTKArZ544TZTxDemBcIc8YMVzv3pZw2nx
DSRsvlwWxDForgrVd3nUQvk/02VeMg1dZ/LQrDbGt/mfLBxG47oW15oOXfiw5oZp
L/R0i0YJOmN8KePb6BtnZSEU4Mssq7dwftl1tRGhVMDOQ4i8pzT1xwYe4+C2Slz7
M91MMgLihE5zXL7KdNhw9IvOc2/jqTRWcwU0q6Zs9WZ8XfFds0MoF7IW5YkPJLc8
egFvJENflUKvU5IFbmTGaYipomDvMFcAFx4CKB2yRu244ZJtOSSKn8ov0u+PtIxD
/Y6HTmZvzQZZAQZFCBVTWNqbuMT0EGJZTS7bsl0T32T0VTKzN1svuJDuMx6yW33X
pzFbv6l2QpwIIPj0DGykH3NPR9wUqR4hRKojEl7j73yrUitMJjxLxOwwrOmxWa8y
SWqU2GBVr53+lPlmxZHbPS5omlep2kuw2E+GbOLGAuX3/VJ6NBwysPCNnAleLNYM
80italgtTct5fJIoNBqYLpC7fVSK8DYOy6s4rtdYL+fmjuCnkLII9OL/IVNSfs6U
UKkFJYAQZRCCFfCNdxRPTQ/xb1gj1zEeOQVpT6UvAjX5A0/HMcnHqrgQtjuLSHvN
TLwpHCYqOjvChXhY/mE6dom4m56QYipS9wnGBbzlzwEgqy37dLG8XOvw2pAGSik+
UFLo7aW2CVhzVGT9twFW0Arekq1yD9Wss2xCGw861acL75vjv3Y3Nc/ug2B4SeoT
vYj7Mdr8ngY5Dl05EZHVopgPBGPQsPSJ+8bSV/4I+fY9weEiVU40MWcDvLacs5s3
A3oYjQT84TBoO0a8vlUHCnaaN/kstnu0KtsBLHph25XUNOz3M1WV3WBvjrWMWZdy
yjAuHH4iUsEu8s/gHmseVMkOpMcitjlV36OZvkRaXkbQQTXI2K4py1bO/XU2yFoa
Rys/JXm9qCmCiuM4w+9n+xHy3dDTD0kO1xAVUIjcAc24V4xmk6e6Ua3fynUL8lbI
QWf4K41ge+jDme8pASzgmQJB6bF4WCkpbJZjE7LXSJtyjGsrLInvJ++U6aner4Yy
6o0ubIUy/rHejZNGOUumpp96bnLHBZiUB/PaiiZEnlGJZs2I0NY8ISCzGGc21WzO
/45TV9Fg2az8kZpugWfQ6nK8h9P2KXO19EY9nfQzsIbG83q1gdXAQHu0rysdyfKj
rSacnYL0OqRq0n/NOuOUUGSt0tvaUDh+lkZcOaHfcT0ZtpRCiLeDY85XXwD8Px5D
7ryC0d14dmRJSZoWoJ+cLsli5xtLdwZHtcjFcA0d4TQxwJyu02drS9t+ez4ooG2Z
v5JmxrRFBSfiWXmi9gVmlbU/vuueNj6BQNCOR0BYQtg33RVCKv3S7QN1AgxZV2QY
vByMv6ZOoUqIxDve7PBDfxHn4cjaiPHx3vBU52oAE80xr5zln12TAE8sBZ4DF1wv
fdMXfXqxvGSM9qn9jeGurqPWboKdgzdGykzzGKlH4FMbxHPUANV/pqTLM3F3fqmS
18PQaR0LnpzAU088SbvQPPmvPnBpsPRebKzmRV9nzmVvY0egItdjLhBC+vO9vZR6
8QFJkAC8QVZ0YFYI6C0XRTuxwTueOUyZ5d6aTbafasB4mhYiZqk5nt5GZz3hLzS0
c2Dbj2QVAETwjt+ZUc54myIp+LijtrQb1R3fd0IUHC80KmcWphnRmHJCX8YyQW3x
8XVSZ3biRubdLriLT9qLL1i3VFYAP3scaKooB7k/bKEWIxFsFabukRDrrnmW/Rwe
iQigABbO4u4KmnNOt31964TOEn8WuAcHIGWUWnQUnnAzZfNG2rnNnenlye5Sq9rQ
GFMOmlZUn/1TMh/TdlBBq0Txi0Z6zar+t0FxOsDYdxq4QI2psjE7JZ1BLeHCUmR/
8A16Ftd4TDPrYweJHsnmhY5r2C/jp46wwn/cGyCKlLAZlfN/eyiuAXYArP8lvF0s
imlSOrP8mvjOf/IXSHR9YO38QsajlCRIZx+uS4s6m/HHu2pTO5qqfqLZp/ZY7ipC
y4B/UZNzHV5ioiRs5eenExIQp7u62wMC6fasvQ6gqQqZSZGQ4vPHYRDkeNZXgq2S
0gdrBWCoCmbmXrKkeJ1ZxZtSwQ1O0Cz1/NLG4Z66HL9crJycA9ni94N9Qt1zRbtz
YdUs2Acq6wjrRiJTy64iJ8Uc5YrDXLQLy4DpzHpsYUzISJHM6a1f21E90Z/nciwZ
b1IQ1WvHr2T9EMOlAPetLVviZGHpU+2gHOOH8nWoUBP3xN4oPsveNNfSiPiJ2ceD
/qVPGUQb3osb/9NHffhab/fSyj6qnIHw2dzYMqnvj7K6K8IGWnb6ATeGB3a/YTKT
CddPOzbEhuJ7PWZefmEnhVtbLaNwD03PalHj8LX/nTepFFhGOzRy+IBZr+GgCRvd
YiyLNEk0pTUqHasOUGW7KS7w87GBP8ASEpZzbWq9dF5l7hs8BEa+hN9Y1tewwWdA
bIXYh9nelDTCMZOUYR1OK/Xj/z5XsZExfRC9SdhNNXb0gO8kpOR7B8bbnvALxcbo
gCuod6rupYilKJVfdoYAt3kDHNRM4rVjyLMO2krk7eQaTuu/ocHp5EKPnYbe37/y
xtaDCFrcKTgJSB6Ov34J7WlXtaLb4Lz//aLKXbh+GP2mf7+0xMn0Ka4AfWXHGzje
oOMWO9rFqiKyXDwLeHpUKut1UWn9JaL5/mHWh3LI/+sCKKXiBDgdfRWxjwgEWkUp
vDPu351VhepjlC2roD5/NlYK+9W9Yguql6Vl+iHY+4hcfZR59gj2JpJuVirZ0KvP
7/gg4SAdsc616JpsBwzQuD/uCeLR/RjHsQ3WZPvTc5O66v65NynlgPvzlu9CSpgR
xOnEkPhxMuZIr+7puMlKSsHxB+2ZxbZOKFuymJqx3eINZRK37bdbfL7nWzD7iFpv
p04Fz5uU/1w3qT7EyZjZzYspYMg5hnCRrlaQjqoN7ptoXQuTk65YdKnRicSMU/8F
Q1as1jUU9SdVy1aimj9bOX8r/Xt3SHPa3n9oKbG559ls+bLJ7BQiYR6P/9fSOKh9
g/Y8HcZSSeRi5pM3UqEGGyt0O1vqWtbF0sBvvpyJRyA4ebTIZh3xmNMAL5sPsObU
iuMu+VjGq84eXephvn9h7ByClD+h1BmL2nTrgLehuyjOLtgGPq41Ac14bpZ/y5VX
SFpRD5l7B9ZGekngEEZ3v2wSRAkICaFIKsZLa8gMI4qh834GT08cTXeAiM377Q5x
2aYbzQhk4wf7k+UsWAJyhfQEcIJHFk1czThgNcLtXFabhQBum865NF4gZ/u+TcFh
XvY2Poxs5LOAMzryyTQ6hgNYCKM9wFwDBB2qnPNhP6Zcpv8sxAKKGP7jrWxxGVE+
QRxEkC+ZwewejOE+AurEpAPulWKTOs6d0r+URQR73pI8fZaCUAAe9r88o2bloPFL
/xLuzKftob8l+ZnI3HXesUYrK/G2yismcUTQXtiqrCyJiESFtXqkkrohLQHZHpOB
/NbtscsD14FBp9mjQm4CgMWGft4yRNDTzSIy7HSgrhHs5FiRum50RCAOadUMHQYD
4CwUUuni4pIGiuiHPJVVadCnEMt1wirRfiNPrpYHb7Tyg6T6hWGX+rnbsJdTpYXs
Ff+wzSlOCcYZxoQwrvd1PNmtrJKD5Pnijcdzp/XKWpWB/Kznqqpwe6aqKz5HunNC
YrkR5c/iDKi/S+eNN5p3GQ2Hnp6FVROUIvfrkmK3yTu5hJbnWcis8pbqQhbo1HOU
J6lfVBs2O11S19IM+s6n7sSbzsoFcXy5LJOL9hwSmFEgwE2KUbEAurHG2fSRFm3O
ueIcAIIN/1K/EUWwhudeG1SRDLWqPq6/emO0nUNQx8K1Mcmpz8WqrmTG0dCMfqQL
ZLcQgbmNuxXl2SykYj3OW7otFJyFtodKzpTeiuI1Et3WBC34E2AMQkkSSW2EkVDS
hgoqndg4+QdSkaJzJ6gdmvzra2Fy5pTOmhc9yaA8cNaWlrSSGuHFruFkuL8DU8Q/
O3t/SG4YdEDLFnj3PiRtRaLsAqXukjj3kdw6ID5kNRkFBCnWLnYJ7dG9EIkTp9C7
4s/DOh/gFDGzO5kH2p4ainua6v0iFzA6fKF0sOxmix/bWBCCWlLgbYb96sNI6Bxo
SB2uVsSFc9uVUQ6VzzamKaWtbPE7ubY1hiGlyQZP8QougsHemOr8K3UYp8zS8Slz
Rjg0AtD4kafIAismP7cDlI/ZkA/6M4ty0/jQ4YU9Qt/SEiEq+brcQW/kHSLY2dPJ
6u7AOJiLgNIuCuctb8TyfdoUPtid8v6UuQiCw+aAnqV9qfVsUAHfWZkLYK/IdBd8
JYvJShTBGh70jt/UEokEnQyFwKz+ynooCoeJ9bccyctyPUqeZCmouQDA34Ftipzw
usZ4OmmcaIfgag/qMkXvwzT9cGHbWgTsoka1PM72iD1doR3zwVQXQgxcFh28+RCN
Un2kMNqO4Y05xcmvxYr8fvEznAOw76Bo8puOWPpAzIyf9THZvKYI0/2GScCQtz8Q
2gaHpY2TzQfw1RaZNkMLPFWchm6v3FUCPdV1sAiSwexEsLSX1DfycRzrhml0D5Qp
jR4reMHF9K1F2itBlR0mJci46slWrqHVPSRfVZ0uDFSJJ5hlaMObVV34xJQx9O/Z
CVMK8oOdXODqpOpKRmeeCcCDtv6SJoutAB2AIWz5Wn488xXCkiEIm/SoEVW57jLA
TTxl7SqCsCDe1fedaUTv6OiDxNcveM93zFsAo/Qs6O0ksKXqHOEtHC9flL0NJQM+
ainMfvPxOgGDG7/ZTQQ2PyONOHEpbLRyfiNS/A/lbd8S39HQeW1UI/AAVJ94Uq1m
lXkzjYaheIEjCfO12J7F9I8IiWSwi0nD3mOO/H7uGUB1DDG6r0Wj9K3mIaXU/vlK
GNhQ+6FvBP0Ig3Z7D7X++YT44UFqujHRF3/73wvSzu6pLwDEtyVnWTPnXaC4L0z5
6JmaCxlSzzJG3yjeh49r1uOSEVy/s2yLc+d/NaXAq0lLotsLnWDydfGKSYonZMta
+6koeHu24OK3wD7t6PWCSuMqtVTqEtLsS66DyzKXGQVHCVQbQOGUo8G29kyRL/Un
fIRMV4xLPu0W80dr8ypHWSzJL6sI3JvNrvO4Daf9kIOYM4hWgb8LLbkfO6zhW9o7
P0FLn7zwjInFpuHt6Bi32HJxi4ntgMgl3RsqVKdSc9TtOsNAr7YJ39xtoxxokvWJ
2qkMJFthugkFCLK8SXJCosYQ7e0NB3pxgUi0a4J438jiqnBwa/FlhZbTABxeuDsa
EMObNhP4RNNc+XZojqtRWRfy1BQaY81Tjl86TY35k32fsGDt+g1A7WEARgOlQGTO
0k7gg2USoi32OD87AdrQpqOVGXPtlMxMRWR7KfcOE2T9nf6JnDzQTmTSTLncJXoj
45PI5/+7WEkC6i+F1+oP7ZS6o0zTaRhkXDFrp51r0mx/9Dtgr35oxi/DvwHmfqpz
gjYM6l9RLolHTts49KEoqVnu6GdTRSAZCYvP0a/xx/3mt5CIePz6EwhYoL8vtIWf
U6jHj2sl+UmY2jdV+M3G94caMXtMaD78T1vptmdbp2N/O0Rv/NEPsni5ZQdc9jVj
V1bz21TABWCWjxRXiArKL5vVvqTR/o29dpEcQIW/jdM9kPf2srM5GlufhcpnArmz
oBxKFu5rhMKPckljROLOss7oO9R4zMo3vpyOUt4H60yLKjHmTPwfr099nlrybkUr
XIYPmAsec6rmEcdbDu32gKRidGRZ2/HvtUUy313gvmqEsRqewJ30SLSEFEFuURGM
SnDexS8n3kfOvKSXvYe36xyhFBe0S3V8AJuI1A/tW4335mnQBmtIReZKBibf8OOm
SauTL9xcUlr9qM5y+vUnhKjlPEVCEUSWLM8jAJRcGAc3iMjKgZ//D47qKpe3JLvx
UXmTx7lfypgfqqhZnTpjOOgLQwhsfjCi63o80QflqrhOd7d5i4ag2WJ2hRtYFEXQ
C9CFNirfCPdRmI4mzhsHOC8vPw1/ngY94T72vHRWVxE3wNF2aUkOemsknrxOKNt5
zthhARBCuh/s73yC8ron33QRVqLeu134gl4nKwm4YY76j2pLnBZxm0Ld6qob1GJK
5tOf4AzOJFRYBdEExS/ED5h9NyFkplGyImWMhiK27PLixlfpCAWX/ZU1xRzRcS9i
pUdH5uVI8ZhhG/dTcQf531ju1pX1b968tLLR2s/xCMJs/eNW/1wnnf1Bt7YBGqnI
FliIT7OfmIZXC4g4b9L8k5cxkSQdCo5mULOAM89xtGiI3dRg4jhQQxG6USZEnP18
BoqHQtZBXJtnH8jPtmquZfvlSZwwjzsDlmw0EQzFGbFs05W6uMRo6/Y1nkJQrgtR
CA71/jw5uqK+/ZrV8Eb8nCSF4UFrB1JuvOQiBSe7W0XCii964KexV5y08IaQTaOg
6dyguM2Z1bWiHQ5hdf5Om7P7eylc18uusY4Nqm4R5IFMDPI497Cdt3wz2OOlh0gB
0L4P0R0eDF8cWkh5+ubTEIYRNZ9+VOsZcQlves5xg32w8cd3ZapN7YWTb1h4xlVq
D6+QrL8d9ucbhYyjuoglWV68ZTTB/yqRbejCv8bLcxeSGj7nGIGPxMR90A2FZkJk
TwGQkpeMa1kZwy8fLIxZ2xrvGg+JXspF8AXLEPjIJjpMdO4f2vpH0jjV+SDAtufL
Rfs0VAd/7584DTQ3WX29anAAKtBZK6tPFtBC8oPg2Tj4GkHfVCc9awo1WAUUjXce
kMwjp/RWfiXSC0zrAULZMaYYn2SwwDDnTDm8F2Grl0nVB02A8jU3O27jrpayRgNV
q3xvAABOOHkVHQxP/QBLvXXex3q0ZerY4vcv4mjpuqyqhz3QK+nwgZbV4lxjymBW
Po/evnKLLOjJSxCNJqn3nZmc48jz7V0DmSOqzQiFIA5x+galNiF9K2PD8TF54VoV
58Oeu3KBsIYg5Ru+++yR2TB+6Bjq+ju6cqIaHbQNurNeKGQhMSi5IU1nsvygT2k+
cR6qk+zGO2dlDX976QG9ZsyhVNaTpr3Q+F9e2sVyPEbldNIChHXkgnAmvUuNWDMf
WXB3fVipwGGW4CLcMbTDnoBH/gGl1RzhtDS1Uy9QhbDeQGonogH8AD7vn9qwkE0Q
N1fV2A8SC4qrJb4kfMpLbqlcFfdppSCQdCJvHYYJ6YXqZarNqrxcUwCdjiczalGp
FvytkR7nzmU2YgigCiG72uzpgUUDsNQ42Oz/LxvyYAvqddCnhoH6KC+U7iDC9maT
djPD238SswVi7TJn2zXYehTbsf0FN82I0+x2a5g4roUMA+2TT3tnoWUZJ9cEnzXb
uJAhwX2T2TMy5uwTAQjylFD9QxD9V8yO7ess2x93Mg7hTEAFt/MrVclC33OVMX8E
Mdw+f9PJ8btTro7IwmuiPV2CUVaToXLSxcwC78tZX5xdYI+B8Uz3MxeuStteagSN
OT5SELOZm6w8H+ScWTU3pFB7f0+4SRO0ssr6ug4iDEyX3QtMgN2YaGonK2+K7fFU
iRIdKPA/dO5oQFMmYDyeMZzLlK/nPqRXhOQskk6298khxCJJeKEjrpE1wuM57psv
B6pZix4Qe9KRTvHOq4AKwZafKvjn5CSyYIqeBrdAEC6A/GQS+Y53neHTGt+11oRC
3499pCN7EDdyy4tf8yCOe0q9F6PVNT6O3loGDuNmsLxI7H+hUP20rj+lR7fGlB1V
pWtZ9vhBqBHFcfA8WN4ahHLb80mJnZPmQfA/nAVj5wTPw8otk3j1BuWxVjk+fETb
tLZVlqsRBuRJllNVuRnTZzWyuuuS2fjszKOlg5HgSjk+4PtSTZsciXmWnLtYNwaF
ZOa92dZyP9N9r4jHcoO6cYn0QCfij6e0o/Ix6LRRdbc0ansSVYD6p5TRfaJaxYuo
rm3XXiIZf5AxsatJCyiNNNgz3CDH8uWr4S/FyLEbwOu03VoOWSzGiwqzBBwTr1ij
hnrSwnUl+H1VTB+lmXoPK2mUzQBRw4N8oroHN7z614Gxl7qoKCFmBKEeGlu7zSNI
BWalAj/DeYDg0dPi0MEXvTmIrZAbtbzLK4T9vL552pwqYcT4asVeC6IBjqn+zBr8
999Qhno8F+YpJhe0AbB5usF2T+vcZWzk7eqhIbO6n3CQxOazAQM/cx9kKX9h49K1
rsV7OG+nRa6TQZort2Z+FQuZx6ksUOnIlVrzZOibIjWlGnwg+Z/dnsoVemedlCgF
e1RpwApPN0Ai2mvpeU3xZPAxS19xv67BLL9tZn6WsYKjwW9ZnYljQi0DKYE+u4bv
EKjjTIGgwnsiFfYBJQXfUz0guRmk/iRjUnSI3D/RPmd6ijAy9oBHBEWDwgImVpxZ
tG3EuzEYc0CtML+ktMyI/qtGObyLmdH55NGvp2yYJsTK3fq/FIGgwwnIOVG5qKEA
n7hWc1W/3rfQAxYzSr+HAiiaXV6xfo9eb2GvThCncOktp1Aa/+lxATGPwZra0rP6
0YlyXC/vO5DRw3q3oi4zdzaY6VO2Enl+9TT5JNDXzSOYcviziq2AeA5E1Tf6disk
MyZNd/VEshTETNyiW5eaOY27fkOUK+UlAF3ocKXBpskidrGseL4ZE8J2gtygRfU8
jHQ+fykAR4XlBpgviQ2zT2gStYSSIato01zsT/K9NyULvP7uBpNsTnUJIW68Qum8
YO4nIOqIROBCFR0ndzu2HjamP7cdq2h+FGmgaX1IFYBSREl87x1m0gseTGQlxJGC
avfXKBCydnB4iaMypcUJfEwrUIKymcQJghk2nvMGu0yNGEh/94RodAKC5jePHIki
IaQjUXJpXRT1/ez8GCGtXhkBAA3nJ3+a2z3KHEO4uFj5yhcMT90RC5Mk5NLGekzx
iOAluhZWInVYbQkgozopydmSyQQRF8O1xRB2kCTWDtu4siC+R3982Uk/wBDZpFye
XJSoZyZyDJZWrsuTcPNuBGug6biZDymiLS3YBeKJL2wCu8E67xv5xeGPxHzeyk+7
vH6RjRmP5N53vpUFrQD2jft6Jlvc42lycEtWxqU1wbbh4igdQJW1+ovDLrPvzQyC
c3THGjIowwIVxAtC+CzqjyDVhA1AYFU8ZcUdpocHujxA2zl+8O0oESRGuie4rqsg
7iqpFJW76vFIHodYepjxlR874c8zvSdM3ppkmmuLh9/P9xftbnNH3N2OUMrzdLJs
1LzJ5mB12L9QyUQevqBb5N1TwUFh7GtsK8j/oXhCwyinSOP/+Z9ClOz3c2/7z3cE
HBU1MSS2Lym/+OufDtnZOUanaBTy8dMGjWXIzATGSNU03kGoZPO4onAP4xmgQdTa
s1i69aStOXP7+ChZeOrv+oscAwAJApr/cZv90ek1Xp4lZK0cIBzmWFoYTo5b+oMe
2vhixH6l/5d3ZlwMjSe5klZqcVu8Qarglqdw2KKKl0Ru2nQFhAOn0LSRIwzqE1dA
HsXwb2uNKU/ECxABcSdlPZUuOH+YyO16tZXP8lEiu5Bll4ixtPies/lj8KtP5KY/
9Yij06tYGAICKA6/US9t/eFApHYGM6N2i/HBJIjpi45i6Db6rPei6B90GjZ+7Ug8
vPRt+pILFFwl6n/h76Rjx2tk+2orqpindkZW8yox5YqLxceTCpFfN7xA5GVvG/SA
wA267NfG7KkYat5vIOOzy1i4f14BVZFsaq89u0F56fpEH7ty92TwCxacA63zJ5ZE
Bo2v9VoEQrbuhebFLdvxhm8r9+p+fES1CXV9GVgaCNnJOvoM7O2kZEb91pp7ASqn
4doofTrWMAURqm2ZbrizS2f26AnK3bnmweahOvSQ2X6fbltSWfm9fjzr6w66nCSZ
TjqWvC5jey+3JAPLSNIfauzDSm6JD7uE82sJaVHUV/To2pArdiwfHrcdpZzidrUS
IYDxQ0HGFO6TZS/3pYoQ76BdWPMnGmXgXJX7uwjNJ545DzN8vqiJUdaW1VbTKVBX
xf4/5rnl48av3mldQZl6WEE9EDK+pUuk5xdiVVrl2vefF6I92QzRSNeBfn7pHaNQ
6cNIq9q5DAvdlo+/NGbt7YDL69uodM7dZpUZpkzej302QeX3M43g16kZ9/68lw/6
va3yYV7rrGR5KxJZHX/Iwu+EgmT70EW44wmysEDZa6H7MzKMAVG86uTfOc7jWcUj
V/gyCnb1m/pR0B8VIgh4uVldB53qxZOY+n6qpfYaPxde7Wq0DqW4BwBIWXJvDY65
F1h20hlomMTRmCxqC+a7ra978PBTkaSmeo54/2ZmUeGEdPttqDK1WlBklhjcneOT
D5mJVRx4FxPCS4IB7B9VhNsVivCLMRo9VrG9GWkcipOtfTIXrqm4ZH+1O9K1Mu/9
qleq+civRvog5cHWgKKBz1K8jsl2AqABbDIoCMI2lKsL3j7FFdqAayCWDt3R2mnP
gkLRS1dMNlJ42yh8ajW+n5WUgcbHpjKPYYjnjwhLq8x7P3MsWlxDr9W6LcnjwwZr
dqBEroOsAILdzq3nMDU88un7D17499KhUP6+rvukdn81DNd5Sfs1wGHCejHGH0Zb
SK/m0S1kjHSoKj2jLjFzvtV5SWtemsUgJMPn/MHSYeo0GRd3zcacrVxZIrFyAy4h
5NU8CyrjstGmOqJ0RwyhctzOOumW2haJzQoxlvY1IXIowoHNfwHMmfS+OgWXe5Wl
3s4ttVrFF5+nQUVTXxul1AEjjQC321o77XvbbomvzAxV679NeiTbvLHYEzM3+Z1G
OYd0XzJDRtIAl6+EBiEg/E0Qx5+woq5LZVSTcndxN/wxfPif8hkQX0b5FdSC0bQ2
9AHIuUyr5rCCTa6fxi7jPjAycEHo8cjTOAvxZoUGsuTGUM3BGSPXDWHt77nqDlBL
B04ird0tYHHDS9fWT3KE0xkdILSRPCGEix/6FznL83ZQ7pzLQnenZInIc2okBNf0
hC7aBOZVoQN+nbYg71esRKGockWcUst+7Qa3WyAaMIz6ce+ar0ldG529+yjmVX+m
lgBRXARg6aCE9O+9O9d71cWJq4a3DSEumcni+m2FD6ZHmFGqzSwCBfnE0jM9PFqf
7Zwe1FzRM6nBQf4uViS9+G+aO7K5BvmgB75SNkhLxkqt60b9AnfCAnM9gi2xiq7D
xi8FF7r+4W8doWhCExHfcH4/LfdzJgqX+T6iLKZYpkYJfKn4PoAXYWts3TO7uuIx
X9wigq3McRilvcByHqEVwcrbGdH16i3psvCnzQsb8SclETCITnsd8OMm9CcleySV
hZV44hy2LUExlNlWNUFSY7OynI+YZ1PfStWXbk04t3i05OnAyZSz80OKTeI/tvN8
rtH+j7zHOQ7MKsMoN7u8LsqLz7nxNTB7u7EBrRzxEa+kuQpUa6YTGvKGHRl+bWpl
QA1hBzsTVeUUn3TqQQsH4Yprt4LjDWisyWQnJgnGZm/4esDIIX5k//Sc5+wfUXan
gG6my/SisoZW/EG0GELHiDr7+NJDiCnecsZDpG90siwlUE7VrnB/onRXGHM6ah+a
pbkZeEkVs/pzWn6IFAw3ToBwtUf4Ni+OaZ4hemtimZn+wTCvY8OMIKv5EmBC/uJY
byQ989zQIVwzK4VUf0btOGuhWfcvEXw1DfScKk8NFeOgqdqi9el1LfbThR4iJvNa
IFir+h5bYguvP3y4yoplDyuAQRqevXWemudq5yXHgC3cOL7Ak92JkB5fA5JcjGR/
zT6AxKt6NvI5B6Su84lX7kaTXsmOmmyt6RsdevJWEjwahHPD4UxTTKlbzu0RBinm
T3Mm/4zMOklW0kr19QSirU8ypE3rI3C+JQXTfRh6adFg5GSNrcnh7lrkLHIUDSpr
UYV/rizFeC52yDveiY2dfwcbB8uUv24u5nUmS6OsZodBCKE2cgn45e40tYs1FhQK
vkWExqFHUJrwY2b3zAf4HIyRFZjJCp6VuPkssufmFIAPWUASmUClfkXc5wyAQur1
aAUceR5NlDSWYJVWwz7Ema4gt3ApGrrxgn9w2Juyt90nQUEYG/ty4+6eGWYyt4cM
x4pkZPdeVlWpWm5GIdUhJUemk0o1rs6Prx+uns3aLkeY6V4F7nv73+VfXaDzZAA1
GXHgV2vELY23QH4ep1a+x0tvy+yoJu6QF5tcfyOGDQEu1Y+c1pyqzMuoY0aW4VPw
aj/zFYUB2upAEHevC8HWpIqyzTojgGeX0xzBr/aMvG6Hv3Xdu6Bwu+Ei6dYh1Juj
flL5re4GY5caaPRNfIo7+T2K9NgpgPuPw2f099cPeu7KQGPtbaL0afsMUSz/+hnY
NL2kzWHS6yn3879kDYT6Zji33UdSQocWqpiPT8R9j4nTcRLN9OaL5TtFlhlVDB0Q
qmfnArJJlB3hCmFtYg8GIU5FSx/aQEFZaNwm+6ZF+rJOSYscrlbxQkJJp7eXnokd
mlhyY3U/RCA3gLz36idN5r7AfNlVtVvYBrfus1y+nAPF0XDGwT7rJMcKPJ7FFzp0
wLoZ+m58XzmJsU9QcZ+L5p5KVzDE2UK/4R1Ip3TcSFFfAtlrDpt4uPnJwQOKA5n+
aqLDCyAULujdR0s6LtudAecwhNHT3GLExFEBfWvLNViYXUZPbxkzht0ael2yb2/R
JXKFrucF+TR7vifsTBomR03Orr+JYbRgZ9zsGlKHQExEAhHOVOfM5cLvG/9LlVGs
riT6uoGXs9yhKi77jWCwOc6BMZurZIVEljDbB/D37nJGc35Qxt1Q30W+k/cKElSy
XJOM7JBHG/tzvFyM+KgQqOtUAQmx75wpO4bHPy4v30c+2TgkdjlPcG3qWnFsLWKO
xSAcdk2VF/Il7SJS6VtzHApMMipicQtrmz9v7W5TVjsZ9D08uEJNTQv6aLgFCVcw
T3+pg1dgRYV2KjTSi6WOaI69Zk8EYXQESGsbYjAXHyaZAG+3ofDWiCsSnCiCZfka
kzc5+RZX5f2P0n8CPNH2KyDHQJkDhU3i8xwr8PQL8o1D0+sxybIl3p8ak6T7ML2X
/WQ+GI3kJGNhquCsauPqma8cDaGGoH9xeEBps4cd7HTyduP/OJJsKsaQoW/WNlyj
DJPqN9lRnecMD9HVzF42VYFAbNl5X0jYpcYdoA6Ab2HmAteJar0qe4wXub7Jj5vF
jWfRlJgpqm66R4c7V4xQ7nKFbtuHiyUrNopKYg+9D+mPNEAf47wm8Gt8BjGoID10
okEg7/lVhILgO4KZHOEPDfu/+3t1UhNPqIhav8bXewE4XusTcCFfbFYeOuQpWOxa
D2+icpB47K1UHslF2chS4XGWB6nnOTZ4NhgGPLOkcL7+wgOKkRTnASefLnvHddCI
KgLgvoJD4kdh6CWiBtjIEPp9SjO0LpgP5BAS/B37LTxcTolzL3C8EsdWYMzIQVHA
KRxaEfzXm+tu6wAXS27RU7N1hltCAxml1FqRO9j9S8OaFN1/PIsPbyPzCEr7xnuC
L+P32lwbfJ8yy2gDnr8u449EIOkNEMAaAJY+6IYwAniRQ+z7TXDFVtRYnCH4T0dd
R12Su8eikHajMyeoLKLdauVrCaKPI7LNxSueyUvm/W9uHC4y5/NvdUrRWDl39m+z
wNYsUCVqxurJbSU+lPjOvXWQrnN3cKcJUorXy4sTwsR2Deqhp1/qWjN4ZJ2jk+UB
l3BL8M5Gh0klSwKSiDlCpH3bt3hdQg2Jzk26FgEku0+GS6u+wihqst8INxJDBV4c
L854IrtwjkLlU6lvdQN9YuwJrIVTNmV7YKIkc1JDTktLWcquKzmY6dmUEIkXKehc
CcG6riOBRXAPXwr4gt3YcNmlp12/+/m0edL3KKiqFNMJXLW1YXdVxgWJU41xJkN7
n8T9NzvXjAaLApJbkCou3ZaI5M8EH/FmpRBcI4tLDGCHZl329/wvxrxxROwdrjTU
rqeZId+bhjlLrKQVz1DTbT52C7pKgx8IJ4E7sZIiyO+z749iIPIe8VK23o+wIV6y
+0LICEVfatB12XAnMr9AmyVdrXRrzZPwkXGW9vZ1qWzyD7P0KeNOC1E0jNtRr5hq
S286bAiKuMfxlBcxYI6wq466pSwyWF4IS2hMp7qm1EYpmiopwbUcA7tX2CnpsOUg
maWEfXbXMvknHnK3AA2BwMsn7lnLokCCdaB65jnjJ4QdJcAncSvj4fwBmry+eOnA
krDIF7/92BCjtSEOTkdPtcFtYj5mC63nO8ZpQRkoKnOCRuyflB3kMkgytdmSqmIO
VDhBCbvZZ47HiaUSvnIDHRkXSM+nZiZdWS/BDtwxcvHyKSuXkTzvz8BcsT2J2HfJ
8wTyd/F5x7gu7K9+bZZfGXee9ctwhdjNMSLk4rzTnd/rvcxHmi2InK2RsppU8f2Z
Gb6Bdiin4j3ivoK6LGXB2XbuKM1IKbDZAYqxCTmUIgUi64NSsrHOzHSS6FY6dsxa
AyFzUPkpwojwgxTw15ytzEnupxf04Uhh8dRLDWl+I6BRoTGiPMHZsi2infi937dO
fDzPIlWUajSXHMIiwJvkxcflZvo5ZFdSabNOCyeNNAMVb653jnAJLkzvHDG6rKA2
R1N4YCXGbHJe95QtPzo0hZU/O9dIo6417sQUWJ4cNTLMfXW9UEOzmh0OMTnLXuhv
kJ4CZTxUlyar1dU+5h+ueOpOsB5/wZ7beBbUGMAKJIiK1ow3hB5hbc0vwa+aMida
BcLY7VmG1b/lcguPWdEH8NsWu+Ah9JfByOBP9NBPl12PvqrooO9pTX4dURCqUCzi
TznYgPCel0LFlDQmnz4FFkL8gGL1oKydaOVolXBQDal7yxZuSnbw4glZn26r4GMd
5RQeXQWJ7djcFAMD01KYHBHOSrZQ2ku9xDaDHni6uNqs3zDfi17c3tUDOz9L/E7d
cbYcCnBSiJoq1Pk3vt5hdNjJLhu+P4bNCHltg2Tvu3i5tIFnoXvbs0Y/AmV3qudE
6VMdwgRzTo2Yu1uHiIgZUGJ9tCui96ibuScndf6zKPkYDrFOVo+auitQMC8kAsWs
kUibqCgGbDptsNuA9W0TU1EfSO82neh9yrjDd6srcafih3AEbJPWcNhQnfLdaOVT
EGmT/z0SPQ/UZhl064HQsFZDWJuOl+jDSD5W5pRKa+dLbcLNj1LO41nCyCkIZVnI
XZGYUUAAuFLChRZQihSOQJx2nmszpT57lUJOmArm2dA3mTWw7Sd7WbQ3TeabV8OP
lVGAjvmyK467/Z+sKpZLc2jfAp3QzzthiNjJBTlwo/XVPAZ3FOBK4U5Suy1b79dg
xrDuxDhJqZpCdqQ8Mfl4wgeQKPtz+Vdul1vcZm51oWzGwxKsH87XpRncOMSgFyvh
HfZtoorXBDiwTdDkNGVISqMDxKsVJ/PFe1WCzBVJ/7o8PLayIcR/yg6c1RQu334F
3gX0YcCfEWZAQh2Cut7YhKtnJ0D23HpsPdcOqOi+5lzCKeI1BOgQSquka3swT736
UTvH8wuB+oEDlvuuXckWk4qqFPBuUZYCRnAfdQ0/Xdl6I8BHZCQsy0MScjG5kc5z
v347Jpzx7nXqwlV97OFpm8DVxqFkFDJSyUWqXJcTkDBI09J502RnyNZNxwP3PWdV
llbKgOSmJ9OTs0rVe9Ee7cpDkByoBJIJMbJtd7ax9h0NePQd+/y14AUIete4rAEn
NEuoWtE8IU5xQCR7ixScxJ7mdk9qAEMXM4cyi+AhLx+dtkQweniSz474pdi8Kybu
YVS5UT1Wa+LjJa46Jyrd7D446Usv+GR4p9ZpxVJ1zbffyS/uygdaUCDJ9i7UO2Rc
GkFZir40t0OFiWX1p+vp4NjJGvAOdb4k+zdSdu2Lh0VxiZzdGq18ZeM0t0AxaM4x
oicw8v97MXkka4KD7bZmW+Tw9PbuXq7p/kpbDdHGvjzu3f/49llb0+Hx+CD0amj/
UYGZYv/W+8cAV7IFyWTfX6HGzdzB6SDxBPlZKA9B8yjsH5WuCOEnu0p7kBmu2L4g
N2AynZjxpNbbInzBFKmPVUTVlDi47ChnkNiVl/HqdO3aX5Rds5OZ7/l4o2Rr3DVi
eaKCy4zfxTMGc6xcahmgLwq1RNWmG89xQAIgWKirmFjeh1MutOSgdelDE7Gc91Uh
3TGIc8sJL0GcMntENaVCJqSwvjagAQfyjQaOlJTrLX2c0GkZBKuWFfuUVrzb1XxW
6RqGnrm7jX5pSj/eBs0gSoGxNEZXMsXJEOwqWdMa/IJvm5E46Q+kFM79vgsyknYh
AMEH1+snTxxM+fZWogupbSquGbtPVBq1w/21U/U40m9zWBCjOqXvJmE2x7/41gBS
qIKnm1X/e3zMVqXsTCEWvR87xuWzfN/KPn0mS28ae95BdW846w5mkjX0mobsrt+0
+f9WKNjhZM/MSGe+YrC1hU59W0Mg3Ax+qrp7vNXKcDmYO6bAjynhf8BKwCqvs4cw
pFZK3JHg9efPvVJgu9ao9CVpENo8IvRFwqILjY3lyOlFAQOQpOCY8K5mQouYVDcb
oVTez6LHLBMs/MdcpBzJOGHoZvie2U7mfPvr/BCSUq0uc3h8EE/F4kYg0ehjmD9D
JGT5Hng12nil1pYHfWXOSuUbeNyD6EU2RVTM/EeNs89vpODalud0Tf6z111ogk1B
gAGvHfpxUvXr/qFos1kBlIGFAI1xueh+Ka+/ElUVzQWwNW7ICUmGs2y+Rd5l7FhB
dwQeQ1vt5PBggnObMmpVkS3PknSdrVHnZUuv7nh7KOnRE4eDEISBxe6stVB8gEJl
6p3IxDq744kUB0OdjBMwa8azxhoEYYk6EMEFZHncETV/oZBjfVzuQqAMzVmb6hi+
dBuixQywW8RnLJm2ZfNdEnMFiza+Qjf4kEo3aRSC4gT91MWu7lKt2eC5+TL8vfZQ
JNxmmcgtefLC0vC/SinKHQoB+hUlmIMciraQ2b4e+i63eqyodYoOKR7dlsgnQLGK
hKZjz//4DDkYE4797v0L8cNgVo3JFgh48crhaNRctuy9Wxh5r+T71FwjrR+wZTIS
PJUHwlhiafnomLt7I/J2JoyJ/AeFD8AbMklY1m9Le+af7PSMmwfyNCwyFLQiXvb3
SGWd5B0ua9ergyMnqqn1X9rrVwtpeYZgNaUykvQy1TTYYCZ9nkD2ovkRxMud0CFr
bSJvIvI5HXu08x4iaEcZu/YLwAtBO6vioIRc9CmsraJRdkQmCm85/WSf9dv6j34m
fuqn+nlgvZVoFTtbnqUHC6fcCnFdIpXwztLHkJIxjH4AsOoKf37557mlXcWMmC9s
vUnZOuMBDKkm/oMM23xT6se6SrFhh01MN/csT9WW7m1Ur3Zi2CZOGyJqGrB81aeD
91utZOfxxMDv+CCWA2kLa9t27/GS/m+b6N8P2Q9BKbSQuuGaHcZcmO0cMuuNgA9D
I2hiqjqIBUEWR0YdiUU3SahQtoIMnDw/xn+mgLg54PEsNBzdEQIqELBSqXKn25/S
hZKc6yN3j+0wGBSpqXkTkFWHezPnKqbb80kJhY5w6sjF7Tt50xN4A7M2NdjYSqxr
JnqxavJWBk/WBiiaw97cOPsWoox3r4xUYo2WuO6H3UCU7qa4X28CHQ9crLaaTH0s
7QWUOpWL4m6q0GjBsbQztsZ3UPUXSWYytlnpIeRKOjUheVi+VWMlEV55Yvar1rDk
iGtzie3cXb1IdW+xX/B81fxL0w1/OTyn8ZRm3O0C1+NPmP1gkbZ4FDWagM4enpMj
hHPiwT5NOaGaijs6EX2e85mCVUJCPVlOAjtc5JH4ylFzEJEBRUnxYCR4RSKqvP6U
SXqPkxsodnpMlUzFsaSE62NxvNTuOGyAnAr64xpIUt2k3y2yfShn1LUnsrsmGG7b
sEmODtwuMj1WHtBOdfMYOh8chgq7R8B/Bfv3JSApCM7o8FAQUOTNUoS+W9guSuDF
UdvCImzStCwHebG9EmRbGBWA4lBVbKEV2PHdjgR+286Sk6mv/dSbcap0dXJ90K2L
tydnf2W6yQOgpA+mFQC9iZJrWe73s7geBog3+xaNfmKJOZZkC4nii0MyJEXOMYbF
MFDT350HpBx+AFhUHz3pkGl5EGfPW2dy0aRsR6+nCYw65aIWE23jRLfjlB7s0J+O
CL49lt82nBRqftg4pFqUP2igxcJM645HZWHSztjAFFHO1gN6FgBrZuUzWgj2142D
+mILoA+/XosesN9hRf7T4duoKEg/Yp6rIMpRUN8K1mBLBBBHkUgJ0h/o1vy1wclu
8DUi2GMSMZ9n14f88AaWSJj9gMVhK+Fr/5j8Bnz2PNCOHqdaMQuKI331yHv0rvi2
LOZfgT50KLZdLNQGbHqbX7SMqUBT4OTOFEEbJm2jGY3fUA3hzoI4juIwVbCuQ6sT
iYp2zjJkAEYfVteuyNIrbcis4U7YlKaPRBoCl4wobLHnmlwVl0oBkY/Dce9IRG1q
rh/Va6JDpa73xRKho1M4XO+5m4t0rHjWu4tbAIgDSmctyGDJ5hexCQnVhBBOmWhc
yRMIN081igwsnI6NN5qIHlhOusvjXZOIdTXEGCtGAHFYgCLyYAti5RQP7Kqz0AzO
GoU+ubwL0TbKApY9oRgJbYYQC9jSR4fhDxLvA8ceWvpdYMp89l/v92MzV92cwwFK
pnP/y8m5Mjqg/VYw7vcAm5Uuxi9FccYNRetaXuf4XlvBRI2emMdGHJh+f5wj+1wu
qz+5nj8a2cCo2RkvrpYh4psMGeylx5zA2JxTb1jYOpOAKxg8Fj/pu6xLiPlVW88z
yiWxQzH+WrOUMQ9w/JG5tzIuSEzls2GEY5KW8d8u8LAgcfgqUNm5FzPDHV/GaYVJ
6YNU8TKDmycmWo1ojaH/4D6LF3NPqwpAsxemlNLkMOJNRzasKlVR8kRNdM7DuDNx
PPBvUVGdualtq8SNKACd2ojFVl7fSohmT/mD3qcY49AZV+ldmlbjHzg/engsBz17
xJkxwT4mj19Gf4ZP6MAxYpLwT8aL8vtkcUZeFU7G35MSf5HHFhFtZc3ieQASR/5n
s7/6ki76s3c3Hh2BT7H2YDY7Ewi85en/786+yMu+ps7XYYV2spGRWwkkbUrjcVKZ
KwRXctu/yvN0PdtO9DNmrRtsESJ+xvc78gcUgx23ZoTDz9lQ7eUyE++XJHRqSOSk
H5EebGeNBRl/7OZxbnrKiUSP8brYy4HGf/kqsW9ePFpyTlqMP0ATKbzmcOyqIi7e
rwIBEwJm6IldEBHemImzlNuRlGnbW77Dr3cJyuP15FF+d3GhVQpstYqDu2pVbvL0
0EYQZgmfAl7GsxQ2VKFckCHqA7QBsuL8gUklGaJH82Dvzygt/WRqziLJ3LS3Cq7T
dM5iCyiz7rDGFiNKH/Wg69DbyEMaAurKNkQrycAmppkHANr8JawL26kZ0WSl4EBm
fdIkCYtweHC4mMaG9X/ku76LCuENQDy0loSu5n9C35sqQuSFwNGtdgLACPKw3hI/
BvtcaWgfyF4nBVuZ1FCl1GaP5F1zH+slFOEmJAty1YEcfwEIeBMb64ZERgXSjiCO
UOnE8AFMGphu+QdQ+LHFIwb7pUQfLEyB17r5xQdOjWPvuvd6UEMQspxbMe8dIHOX
lJF2HP2vXCxbWCNSmLxi0yFJDOVE5iR/0keE/Sz8i9UMCvgCdHWY48rvPwEoj0GW
nk/qefECfvrs+EPbZyA7rchfykODtWqFuLpihKI8sdkW0wEH5c2H6cBEjeR4JUyX
YS+bJegPgx5DyBq4zSVc8WO6jwVMBgyTgtUcXuJ+uFkdsDtoyAL+s0rw26a2qngu
Ms4q3fbt7opKx8CkMpgqlfeQ3z4lpTsilzVMvi3M4iUv40SU7QOWHU+sOUvFnTmM
2MsS4j6g0oaHU41rF8wxcRWiOaLqgdyDPBeVjPvwySHlW1GeqCWxjib7eIDES5Rx
w4aYdr23HWdo5Wej/IKFrvJpG4ClF9u2Ee+GHG7MCk4LHLYFSFsUzeCZN03mfTtX
+VAd+W9rCwIftygWePo4Hya73mt9d8kzbQsEgxG5diHO6FtQWBSVe3LKGWP/c/3o
OzAOanVp+rbCHBw+zMxuJu4GcmT6QPugZ11VTcDF33PR2VBqEbatXDmwmCMRiGLA
2NbT0bMNdWkJTtMtd9jJ1HF3b7VqVTvRyScPcf5KH4OUh3ogrdhIkKgL3Us7UzFf
1JG2816EmdKoueXkLXsghs6XdLyC7SUrzkjhGA+IIyQmyyYxljMvIp4gaSlTfZUM
Zxwqf9TrUbaqz3PaIP47FihV5L7r3FIgpHQG8uFkQpkXGqVZCnU24I4AxUecZOAA
FRH4SxiW7QgiUN8bL7hUpVHHQmNFOcgHi22nRIQGj+kM/HILDjw3cOGOWoRpGpGv
Knnreg3GDdAjedtk0E2h9YYNNnsv74h+erH+efc3o69OgwjshgIglltU1GA5O10s
1DixFxzayJK/DvYiY72NkmG/Mi4MmteAjcJ1qO/xGXYOogRDQnxQdbVgC/orz4Yp
8nHLijFByE+FYOqjV1MEqnNun/Na/MH7Zczq/joHLrZiY04yDI7e+aMEUpN+AN5/
L65nlPcHl9VStBRrzOQSwkxK4Q9CuOOLsIvVU4N2tP/YCXu00XUVsVP7A38sHOia
lExeEAv78cPYX97Li3uhM3shJTPDYOzTUzC9LKtgck8n31bVwyzVhx1abFzlED+x
+uoieMMtb5TXI4La6BGXG86SRsz2BV5JuCj0pN3ngY6qs7YAlwD7CaO21K9hxlKf
aVMAXmcY+/73J0CluPw8oVB7Qwy0fhod25seI04/xImL3CXcHQGlnewp9SHCWyRB
vFjkqXXB5os6ipa9wVqU3zzqI9LFmvqI92xgxgV+Whz/8qVSGuEQRerqEKqu4xhK
hxSmWYEcpJQQWvIpQHB0BY0fcKdJvAvklXAAchoIFuTifu2u50jw1jpavGcjeOu3
nXhq7ZMxjF+5jY0XoS2TNY46zVdqZCABQ3me/J3iG/odgHqr/fLdmBiaaFr6R2JP
RbqCB/CPaX4itk1mNk8APPegViM6PF/71hPA3nTu/XpI6NgCg7WUWXPblHKqlCvN
Yz1NhLaYnaU15Uo1j7mvW/DKoYeNGWeQMcWhy7fqq8fWrvdhB0bo6oIik8VPfPc5
BtJs0dxUtJVqm8usWW4QlTh6LrIsXFn1oS/vXZQDLTNejZx+CzzzBWDtMZpsweQB
zdp/bS66cSxmEs8iwVgnQZHhtuAJRvMQ3BeeaUEkg3cOK8kuTmNO/JlwQ+ioI86W
WRRmhK3g/wZZO1gkFTUS0arvK1x0exNkVSKSYxrJ9wha3s8N8EWcfcVie2CamjVA
qC0y2hwDlQr5fbKWVqWER7cPtQxfhyBoOacI1niAYHkPSY6wOotQGP/p4C9We2ee
EvBTcxH9vMmkFsu0JmgdZdpr1wa/Cv7oK6jounFSdj1FZx1ocF9LnfhqUAEjBGQp
CW9U8WYHqW99rAe72Pgmsme8aRPP3Y3OO7tKLYlm3jj9fBvzHbYi3Q+7FhGpVHmy
l6L6lsIR0Y12gBXJEIJvpcdmwOOL80gyyHpbk7esv4M/wd+SynWMtmF/sn1Xk5y8
gmyfbYrZE4YUjBT5QK3vx7LQDA/GtkN3kfyCAj8GDemIbGLf79qeH2TLBs0B1W5D
FzdmIuBNQs9G0SXKD7I9UvlF/wK9Q4mSoe743OIqVhgey+IdfmQf389u+XpzS34r
uaTYPCIf9pqGv/+5cJOkz0rf+Drsdoip/HNzi3YoxBoKlOZJxhF7PcGEB1Cv+Oyd
CKEChSQN0ye0Up6Fle3FrvCwkE3ywKrJDDLguQSd2MsNzKls+XuFavBAhh6DAxdr
5p45N5f7nHSY0RJfWqb093pMbXhLq+v9D8xGvfcV3WUFWdoo/7SsyC0komhV3H9w
LIW3vJ2wTMX6MJfH0a71YMQSfCxH2QPZpTlesRCL2AxLeWOnQ82GqT17GLJ/mOWv
Ytv19b6RyiELR1BA9KPBly5vaqmn4rvZiRMM4wArMxs+kHq09y1qGvLX5zNmo64e
597EeLx9awZ1546S7AUr2jQddKv/aCIMzkuejzymrf8CFdzno15d7L8hhx9OVXYj
deCqmuDAewfwszzyXsNOtXp+l3JzhQEOjG2oDU8m5Nej0vmpb902IAb1P/Ac5NQn
kq0cRokK+N/G7G5kzXpRix0Ic7dlSapzlB+4gPsXrY1cu6P406CM4KJYUVFwlW6+
tgy+ZB+XURTvQL5zKX4lBs/zWwirlpMRU+KPaxMidEBUneUDaE3gMhtSPiJqAcru
jIreq6d9wLLjL6TMfTCkBJZuVvHBqkJhffXkz3GEb78TuEkCUAI72DHo9ax9mhgS
RjvdQTfs3btOhMSHDXghx5q1IR7BE1xESGZf9Pl0PHpo96Q9Xx3tXkP0Ba7Ekfnl
uKYeZdYQJB7CSEffuZcbVIHNDLpuLhixg2RzTkYX1+Kg5EcMhWuZvwGV20bvZS9l
D+05uimyJQSeHcq4szD2I6CUjdQ2YwkqbQK+54ITHKDl6cYwl70AnQmqFlDsvmmd
A4V47hSB2jG7zmWSxqhh2BJlH0SRWA29X/vxyOZtVA9y8JoN/bQXvsDN7dpI8w24
8G62IjwM1Dn78zRoHidZsMx5szJ9GtYtzlBdv9katD1HV0lzCLTik7IoUC4XrByt
Vq0U+ooipxQWUTIXurbX9HotbjBfqN7LiwNLkdtn2h50sgrwerWSntabgAM0hL/o
qDkFyrqEOcQOuUQmbeU9rdk4dWAwhYiLSoulV4YJ80aLs1viJLPT4t8ZE2zGPQRk
DFu6+XVkHAcEkYkh5ySkt33u70T7jP8sEi5yIA798/zlO1dGZY/YHDRIcbuK61F+
mTntjcb6/lNyMUSIrx3HAR+rIL39b4PIYuHgy+Sj82e5FGzwKBQExcWcD3FpUtVL
DDuS9EwhynUnLattNCiU+jNgJjemYw5i9f+TdcuI4MsZunWxkLLOheVoIF1+WjvV
/COrs2oR2+prgh87Q6KMrkRdJwKidSkFfTDEh9Tk7UCxe8MmSSyT3kKb69GOuSy9
VKnrWQyPCz+0qPLq1Lnf/JPAUkf8fjL/tRPpBx+Nfv7lx6OVs2Csyu+ZVatNC/zA
4ozGVT2JElbBq2OgmMRGU8IXsux+8MOHzy+x/pKncwrBZYMS/CERPf9YOuH94pWI
nb2Q+Ocbg9e2+nCzD/VYBAN0QfizPRVqIGN5gV2cWOgNz015ThfTny2aEBvP5B2v
Ipi1HVXsbArVNMnZWSH/SOxWshswzpSZQFpWIYIgkLvGDkw5CYnb69Z3n3YC+LDN
gWzol1goku4YgdIJmmd59zBHJ2nOXr/RrFdv1tuygHn5dVYusGaU82LxAslGhnQs
kB7kTdGUKUyQmdy9+jDQehjQURUZeKnNCohlMpRGxQvx9wEUyaI96awq4fwJzF+Y
S46B86RhDFWm4XFeeJE1kEsqCILrZVa+w3J/JAXr1f6gvntIdznf1xajduGlsCH0
hKirzyz3YQy5DX092SrDeLeo+YIHb1KZb6M/Cn/mKsdNjDQuZg9HoXRgiVedQTuo
3AqIeGPOC8XoMn84mdp1/eVYZWboeqOvstW5zDdy8mxZRLzMR0Xr5hjhMw9d6QVL
sbltrZ5twh2JBhUUOfYIJ47yuMeVAtASH8rochHGg5Fhfn/8OjIkJPyF+b6plujf
rXusqTsSjFWOLpnnXSp1KYrfA0vswTtQ6y87+C6PVxuoSn+Fo5mDzWeU7N9CLJDJ
WsXBptfKPtXX7zgR653jG6MPiNF8R5+R0lGk2U6SpxtOsM89et+GWzQTy+sPQoMr
jidVJsDRUpSRGDsqe3FYUgvKcELhLBO0VjyV6bRbODmfwfKDO8cSfAWseImcBDZA
34pIsFeHgDzvidNCEfp+ulT2yA/gVCNLpfbtXLPF4DVgmdjO2xRHSNtPtM1/teCw
Sb24jBzjpdvjtySrpf4zUi3pffhEQUrMTJtrPs2bjXs/aD1ojlFfaF2nuRQgpGpr
NVfpJ39bOoefwISVWG1F9RGA41oKm5WJXHoUm/uks8CV34lgOuvVaADbcBJGuJAN
hf6NVzA5nL6EJqIcUb8cPrZDOOnPgmiBv4HKIIknVvoEMf7d+RH1xGFEBr3ek9LO
jQH7hPzJs9s2/EYh4WQlOprabYwgvFD6m25GTg1TH5DRldK9Jto8BsZBdARDE+rC
PjB2zTfiUcbVHTIWohlg9T/hbCHFL/7BVKALxxB98sUgSKUgwiYYYZfmzoHQ+hf1
5iqipqdOQAwnn9cQWLRbEPDjN/+EwJAxsy0+tkOM4Npk2Tb/kjYcTVGm7Dq5ajbs
oYhAXsSpEbqL2SryWqj9IcvHRcalysxv5dKgCTbDGzcaezs10iGxzhajPQR6xvNt
nj9XtHEFweKANr3nxp6jnop5s7l5F+63G9fxmN6EBEEpPNO1i0JHgI8GEd6YGvcr
bhuXUV9SMin6PF7u71G/KB5Lr1y17V/oR86WxPPPF1Ig4OT5un/3Q+Tip1IqTVdF
g5GpNFSl3/SCdlSOoYl86vP8UaDwGHdfJ/c2TJXZ82UZIvTSDbP9n5UQRQ7sYSPz
YJy37OoICUsrG2QCTGsFjKB0l8SwYmlVYCdQnx5zV6enN005XBA+GgvlyzkmARBQ
xiU5rQYRJWjjOhP3jxwXtFZbh4oTrBjkXjulERH3Ynf4ooVNT08Tnvd81Lg4fjIu
34CYRiwxRs8N3wZB3niXryd/D2tO/oYZRHq4YhWidZWPtl/AMgnV3eaN3Xq6wkp7
ATqsd2XWrR45CmsVmLLWXg7anTXXIVLjx573nJBk4nf2jyYq1M4nYWUOzLWyYGXT
o22OOE07dYx/ID5xbx9wu2pKkfVVL3Xc4TPDmpQNN7df1Ld4ozLaPeVsEGiR2Gw9
vCP2QySpJCnsMNCYZ8XGX+mrA5249jOUWoBimCHhIhSvOWak2KDz/UKNqo/1b4MU
iymoflNlc73vhD7bmA2GWKV61S4bHEF9MInw6GrRocDVh/VWOXmi4shvHSb2PXGy
qC3U+dpUuOdOjx0UTaoTLmxbNAsqNNiBJr2+HuiQCRT8Cgm69lKSXM627uD/LfFy
xYwEdY4i/KDf+i9n5X9PC9lbpRpB8+rYbxfg8n/99w7GrRSoK5kip51O3cKjz/G1
STzb4SN50bV2+rMLHd1B484CW0zNmrhYJ0+UW7N2+wMd8t2VlpVUiD+QkGFxaylK
D0Kk64W2KXBrjWKxE69cRow3A6GstE53AH5TuQGW2Rfk4isgB4itJHXfv6cpUDl+
umNmCtWKSaXAx9Z1XIni4dH10WThcgcTybLugNGG2c2RCiZELiE/eew4ztibRaqm
YW9/jXLFz6DlBTVl0eAy8X4DKt6GUH7aaqC0q1cqFxRwndt2i5kom0VvxkfglkaQ
NGev3CNYEuSdXzH8klAFD8alqM5d9xGP0OZFnf+AllU0rgMOur01acO3SXTdWtGr
B2/DfREBzZ6YBgxcl0Dtiq0KSlkxND1tuO0ZBC6gAEBH/ZMyZa7lpIH0SRpy6lxK
FYS2Iz6a7CPerdhQ7PVcAtEbaBv/PHy9UUtxZLLNkeL+GViBonExTt9A9UzXd0N5
Ua93yGrNfNW6q4PTX+Ytc7VDBtdYWyJ9FfrCzJO1tBPXmdQ4OBvrVzqLeOQxpKs8
k7452kig8JXh4nI/Lp5I1vya7+hcJr3sOEnP0oWBxlYnRg/4jn15trqvaNb+DYht
CPQk59CYmUi7zfMDn2eZuQvxX5ZamYFmjxlIZQl1QwXaUJM2pRgpwDzEfKie6bdO
VIxSJ6Lu1cBQq3vyPIx2AkMufYhD+31l0tjmyxK7P7nxuyJyGQ9Oa2savY3q7h7X
ntM1Q4agW8T4Iz/iQIjmjYrkly2kE4ypA6Khc+SiUn8kucU86uuv8oh0oD7tLe6j
I1Jkq39QS5iT5O4QVsJBYmCc+kT6T/G+m3bFmE/07DjO0SWyJINOYHXoUEJBzLDz
XHcjWd+1gI46ICXJF8fftgM0lXUFVIY7kI7QMTdrhpuVsOwDIJhugto6DkU8z7n/
ExvkLkeqrFezy/s/taEM+igxOJ3/i1qjNjLR9Wo+e61ViWT00R+A6zDHHxwPSV31
g++EYVCvbr1EEZR8gMwMHk0uWjcWg/cgpa/gh5sT0W4g/BMZ7ap4NoTxLBO9DVlf
OLSaaKaBVHN39xhk75ekX/H/fLjmk7s++2Ecpo/nkJv+Z5wl43DHMQe+f08zAHaV
jyKcQhxVZ8hGmMvpJdwsHLkr8pcS0Vt7U2ADQKa8P6MGmN5UXcVBKiffMn+K6KTR
+bV4CF+2Cwpw0RyZf1Lt0R9+NgqgOkMD1cD0z32aj/+QPgndwnNt53wOS6F3JTu6
7DiVhzLJxWcJRAeniqFS6ntLJqlI2jmAukFxUNdJBfuNYF/UdqpYlJkeKd68dBUy
7LMQGsdNtXeyLoEBOaxPSMeXR0iQd+lbFyV8ww3Xg5ts90vJ3Wx5ccbYWnQDEsjM
99SvQuLjwZpx+iI04Dght8aFhAOErk+VDdhm36UdaLcQ9MEt0spp4gdf+YMry80c
mzdg20CGNdnREQY0IgmVf1o8tydOH9QyCMio7IEL7k6QD+RH04J8JFdTPWZuK34T
loDlpvE5KOqywRUL+WZbkSuVxbBdHZ9OlzH34ttt9zQymrSqUytTi/OgbHty/fMt
CBmov2lvkJfv3wA9avRjv243TNqUkafKL/jYFNMOIn2gwAoppVflcO1/2KiWXbSq
nfpJD6r0X7FdS1aHylo2JsaLa3uZSlwNHO8v6GCUzxvEXMIu7o4/6zRLR2XfslVN
xqfaz8jByA3wlaG/zgf1CM5/BbusfSNFRfGN+kaSLXUKALTqn1DMnXSfoO2m+pRQ
SeBNJ7Qx7wjrSWvh+0hz8wcTaafuj9f3qYAKc3jq7Nbb6iSBB069nhe7A7zVWgrk
7ZBDUqzuCM3oPYMR51MPc3iPSHayQHn/Lg85dl49yPhSJxIHUiqnW/joj9XkGekx
VbmKXt6DkeZTIiAuJy70QdfSN/r8U8zeQRM5P8eREzWg5A2RmILxaHQnNdql8dZg
xzslv4CYO+UlBmjqraEUGgUFTNnnGK9H9YyLbP9fkwl8y17S5HWh/uG7nYOf5E24
7qlvon/aYO2vSCRBr5CQQuJBV63XVSU2W4j/v0YSzUhNFM00CysMxHfMI69TIMyw
5KlPu2ihEk1KdbNegHDhJirY3pZLeb5Fza8OPB6wGiMV5WgrfFti2PixA+2QKadz
qBSttprcp4XSkP5byDoDyjFnFtofc51gprPtI8P0+h67hZ0z1WyA4r/8xiE2a/Ie
x4+4pvLq+sxbT/hHInVzwsVcnqjYhUajgIK0LCAuva15bGROsFaLzZ8faGGR5OrH
e+oEXrP59A3XUoWGp9myXsZLl1FrCLZtarE0GgIOcHCXWBAdyP6g3OpfjU/3SqmY
wYgVnBFwQM2kvxfhtryJE8ouKoG9wUVYT4z1/V+oG463Z9c5cJtAXa4UnmwcVvW9
/0RSZc/ndsxM/+BrAlug+Z+7vOpUiZuNx6PbDxWfVQ/BLpEodH3uRTZqydjB4O26
0+WaAS+ZyC57gwsqMBDdpQIWbU90Ub9xLcFBRKRhlFVZee588T8Qmw3yI2yhv6/2
22MEh2kIF/XPN9/oLDby16Dr8ZbR2X7Ia8dlnwaKhSaFuZgoyQQoF3FYWU+R1Viq
gihb2d6knzKTB6QE4Wg3GT1tpLywf8WnLdqbIPwykL4nu8+/77GpOJZzQ8luFrSw
MAohKLN8d1kexI7qt5Oo/t0SBDoESBS6qXqBTb6XA4Z8Anj4P7mlqVE1Wp8lwKd5
9/zwcs284a6ooW3xfLvaWJWvssE8wCv5tAVCV4ALvdHQG0iI/16nj2GrvVSP/G1b
hHHb2mEhKW74eMrOPFsxB9K7H3gh/+KH8eEqdxAj5aJMBGTC2d2phT5+haF67KH4
zhmmUvxaobcScLaUAXAVCKIaAO1AxKKMHLE+/gXtBtNMC7OWkza/bX6JF63c8OuP
Eou66+Ryr0cIs9JLqXop82XxnUg1inZ0FGVvuVk9snUtj/+qmXi5VwDzK0jxJ0KF
04gnBa0OdJNJygClJ36NQHYoVt5JFXd4j04pgo8gkxwOwj/ywKYz1WHG+rc4qBki
UwVKjbE60/+F2gm2OIOzH/FkVRVeAWE6vOl5itUlgBH6tRgjNkP5kZD+YLwPvrtR
+k+4xyMnEWKDAAHNGu/MI0pwimiNT6UpkSfxpWhawn2PUhKSRRSG3DEcAtTGkGFw
sYIKmDMwO9UWYM7lez/kw1bfM/ii6owe4rVBtyARWuChaU/5yH8FTHC2wDsC73w1
Sfpnc7ts/WRV4glEGf3JT1Aa+qp/+9rN0fY8bKYk4+CsgQLdmOgTvMjrlctLC1BN
+cSc7kt57I5WQlmvN6CkIiYsE1uviXGF9fAX923Z9Up3WpdIfENyLjq54vh+jv/c
6IOsSV6C/74u8ZB74zu3HrzOJEbCQE6gCeYJEs45xzVUkKZjKxqbRadfhAWZ383c
mzOz37si2KbOx9Q3SzR9LGd2oxb/y9rVSATB2BqFUTzRgg53bGwwA9cnu4URdEcX
dyFGlhKW1cljQ+28iQKFksPyOpbZfal3RVnYCutP10elkB9XE0TTwesHzD1/Gxya
IMdy/Ux9aqHAeU44GmZ4m46TrZFZDJJ3N4Q3oXniztCr5h/DGxU+HfSeaz9ANWzO
ttCHFSYRQbueXh0tux6wWuGqcVL4HW7LNe7LOp7a2z8d0KeiASlCRhQ9iWfirOEB
L1102mTG38oVHqYWaueNf46akyNkSt8qruaaRwUdsWqPOgnbUOLWq6eDI2xPftwl
AEv2+KNEqW52WfXXmycyIvYAuL7jTvTHI+aTIUJZJYWDyg+KcBaG8C8QcnzfcBJg
KCg1bIcs3BKLvnlEAgGm6t2n7u597Qt1KhQjUbU1h2OHdaElx61FESd/MhuZ0EqV
nt/3MacuIFPzcctm9cYsz0magWxwmScgAFyvzH9aAj4cJYrDqTZC7QbopEQ2I4px
AWdhHyt06GAwuMhwRaGYsam01kNEczY0rLxCKN6WN4nPgrHV0ErVcivJRt4nKxx6
WYLI/y36AJ/gupQ9CAWNw0qk7l8c+FjPem92WE0lr9xEeZxKI6UflhPwXRUw4wDV
ln4iE2/2KIwyalL3UUqAXYkmwfAlzbZ3EL4OrbXvUJEL2U1+kTnd6OCJY8har2TM
wL+mlYZh0jXHNjPsnD338A9XFWKoEA9NkRDasI3nLDHLtSo8nkWnn6U1l/To8s0p
GVT4tSjrJdewUwIw8bV4hVv1lQLSPZYaYfdNyebCgxqkWyKiQadHbQtwFLMyRrrt
2xCYZ1uirV1cGPQUu8HZdFeBhErE15DXnxRg+C7ZpsxSCSo1mqSZmB2aojb/qrxI
HEiAbDHnNqQ+mUtZjqGEJ+OOu425ITGoF81rbS4VPe9Ab1bEUOXb9QcPlcwaLa1Q
bw4aMobX1EayNKyPK28JmcZmxMf1HjTv0V2actTu+y8VczsNMAlcoruWusNpxdLI
c55vKiHC4IozVGRNvny3FAD8kp80MPv9NeyFIvp3DSk6Ps+Hx7P8r0LkI0DasEyy
AzW3xxL8H7ocOP+gHleLuf8zxf87MAZ+7XJmTaehnXF1popHa5s0LEGRb/eENwBw
/vjCPvUzIu83dtoIy+bXF5ZLpk/jJvtnVxzZ1WtCaZ5hF4nhkvSKuVKsb96Z2PiU
UzaYsNYyTHOAl0lS4QOJd/Iq2v1kHkT0g5vuD3fkVJGsdkis1mfFciqTxF601Qqr
Mabl7uQYfnlF8+J+iIi42VNXAVeVhn/mAbrA4MRASeTjr6PKKxVJroiSo3VE9QCE
A0O0O3ATfRMDpGeVOPv4GOKsLFJx7lBfi9Sa/GCeA2K9nbri4q8eyRyTprZoMc0Z
MSxQdsx/AFqjVuucOGMZtVgG0dkc2PJ6t8PRognVNJU1lBYfA7CyHvFImCgRq1GJ
JQ4wdxQKmjKZeUSEWVf0iQDZ1z10tez7SCaTHcJdrPZJVRftiVUkNrWyw94oYO45
7wgxkidekaHU2D2QLutrsRsxbcKbaOP0vvhXvA9bgpZDHbmc0/67HOfCF6kc35Ff
fWweBFBOSb71qsoAZfN+y4b629c4GzOXGB52LdtQg8U/6iQaCIkb0g1u3Y2ldvSs
zJ3+OoGFgWBlCbXxVwfyslODUi55SakTBG9Xia347GkBvud6heLzGh3jzuH7ivdI
yRDtgNqfz4t4tjtiUidGumDe4mrlUks2ao6RattNV/IL5zjJvnyqclH0hMiZDHYU
4e9jp6phMPqgT3if7AhdXlA8WUlinRVXAUfHrzWl5VMwOBJrhPSI+Q/xRkJ/PnKn
N1HE0HrC58bskz78diqtDxJ+Z/0k7ZKPvJQ6GPvpfHNGsAMV/5yTJnIlZsc1YCIP
WsaOrm0Y/U2ZUJywsn6DsxidWKgV2Jje6S5Fsk7pV/ZViLpMZ8ASrrG7bRAS+sL9
r1Ofg8yVt3y6ztUSD4hFJKtFnW08B3t0TT9btKHGXsWdhFC06OkzY1l8NmZmGcqG
sv8PO1X+tm0UnC1pjkWgYdM/Vd6IVQHhOhBQiA6ztnixRtyiKJVLu0bXtPxUDV+r
MBo1M6B3+nqkHFIiccXPnq5+yeCrZNnAabTV+Ssq/euuEdNlSdwgVqpC0+ZyrHRv
5sY7R0hIxQWoejjFWQIG4kNJkwN0vtHtfpeWgUc3uR470UlczhhbDU2n17rJ0njK
qStuLBIWM+am6vPhUJaZ7XoiYFLhVN5xh8gbuW+KJwsTSLkq8UbAbWHJvKYB8J1I
38MtSFj2Oym61dZ9W/ZapQbHt+jcBSJpUSGFD8z//Zf31UnP0GOPMKGwSpdekhwo
asf8IZoh8XJTYMcrENBwUFJ/iQF/AYLxlsGMg0ZFWA6pVvH29ePfKrEfguKgfWXz
9fCigEVwp27TINfURquwaoZQKXs1nT43oy3Bf1gaj7S9M7A6y9yOcFJcUKcwgmRg
P9j3xGKRGS4VGKei4Id8TpfkDADObFCVsytzlg3O0ocQotZAfnk672m9g9jnj4Ol
97Ubwij2RG39hrx8yfq+EtNPWqr1d8YMgY3b35aWtRdpJVesc1WmK2n6aWJXz6k2
W976/2PncPl7rp+NudycZVy9r0IecZN3HDeZOojsL0tfpERzrs7lf4I6rm+95rNc
nhIPk+YlMW/KNrundxYrUgLIPn8QycbHXZTUy3FZ7I0vWIX2cteBzX8OsmCKh/eD
eQp5LYdgp3Iz9tckBE+/mSwCR2chtWB3FzIJFkVtJbm4jOS1yVU+KgZYvOe9dzdd
by9mFs1UrMmh1+cz44cQlFeF7YLePMpYH1qIWZDeeK8TeLCsoIiisj2v5w9R9Ezh
gp0fefrdfSAjH0l961Nvk85rxSZc5LZ944mw+WsG9sYa8BKAvWI4HYH7v4IFNNPy
jOaULkKKMPGsOF4VEc3GQthANsS3JPKnO8qZuZfcxZfTClFEt7yWeXt8MxSusgVF
ZDKQy3rLFnyPGRlNLe/wqgnJrZbKnWjalMISi9YlJszf7CfeoKLA3+ufITQpSoAk
Q0DmGDfG+Y5jKmnwkMUg/pSuZ/1ukCu2wNCNoHc/uV8z/TjINoa89trKjiXdDdcE
ZzpzYVsA/WJ4dT5qe64QiRTltHylDLNHHpsJa0pjkqQYPXlD0iWGpIR1L7ZGs7OY
0XX/VYBu8O9mNj5eBo1ITWegK5xTIo+qAk1SZ4Px+MFEj4C51pD+yyaPiq2Adsm3
ouFMme78Z/ALlKdOoRakXCYgCGqH9zLpqORqKalIZkIZF2w1AMu2qmdWONIOg2il
cThOD4EnVnz6sjN1dz8USLHsqWYtgaGRcBiHdr5vhnec18cRDfrck4Wylge8mglU
sTywv/k2J0LsJfi92KDYUUt2q5GmrA9MAB8ywTX229j2r9WDchBksqY3kw7RqpoO
3hVm9ip9mOD+K+riFJKU+8p+7p7MTJLYUCrCziLcpqVoCZLbjg2vQ1BRutY2rSui
PFoMNj+glqaDKTH6/c09M/pJxXj3FzLQnHyeelCENddSSZeiNTizG+x1P2JUvuiB
g+DwGZKH/fIlK7QLM2qWmlaeAve220xLr7pBCHzpSAXzMQNM5SHQxzPUah7FzusW
3iso2sfBPdTeqPggxylf4znjF/2Ur2UJv4eSxlY9nrghu81M2ofU8O9cXHlTkwyz
w+NqnVRi8XOIFMN3p+STKsBE8cMs8G0wc4wYvMMjwMBMR7cq3SN8isNkWsBcgnST
8j3ywnix9sC5Vf3fhrFrGSQbEIVGS3ksPpXBUnm0CEcNcY3mN8zx0Rawxo0x5uGc
IrSOcjdJRb7rbNFW8Lx8ctUisg4RXBJyyGCKfCO+/Ja0C8K51m1qOz3jwz9xcAVZ
x8vinEtALPsgWENWHBYVyP2DbtxBH3mUmij4AHipXAzbNDP+uDF/isOCGoUvLsPe
Sr6nTJdYbNdxvBYQ4Ze3B/KKNkJJmDdUJr63BxJy4mb3fOSImYi0GYXGZjws+jDi
RS3YHjOGRnfKJCDdS6QNFiFna80B7GPqDCb59jbUXm/acJvhyjGxfgo+VszbePNE
FO9VlITb31KIkX1niKkT621+53KizSeOYplPkcyPoTrOys1gOErg9Ip7x6JbCU7L
cwF5bBP62W5d51RIAWNjUwyjAaR8jkFcByDkXJ5M0bsyJOfaTGjRN/qJJuQWtR3p
YnZY5h5JsTCWC8lDAwFeYhGvAQYnuwd4aCnWFlMfChIZketrjAOA9672WIHqsrt1
3ZeEKLpjY2U7Fc7sttC9YIXDQKUw1eyDTtiCyUKyKYM1DBT/uqYazNW/39AjoRlQ
65zpM54NyLo4sKtBuBP21zyXLPJPnql9IgF2CAUCiLHGwBk3OtjFiM1IbXgdpIX7
wL4gWExkRcrlBRO3+stPa+8t67iaqkwPTVbs8Qs/3114pqiG9BicYvRZATFQbA3J
Qc7oAzghsS84nd8R2vcDz/2wpqLf3LiyEFZZUbHFqj+YbO0ZfB4fM+0uDlj3dFU2
M1t1spysZTYBnv6TPtoP+P8JpWs+Prop3A+A/Sw0hQyjjPPdVd5N4kmeXuXKFRO3
3pEMsva4nNq1+OBNxzclhXZftNi6tYVKkFBVaHP/50yuAF1Qn5sR9pcI0FsVuGoc
oMQGbv80//JQ88aviaLTU2lijcFQnJTNgXUmKaKmTFdiT5rt7yZYzUCpDCnGMee3
zpK5lCpyzkL9p6PAOB0v1qgTqMtXzz9u2AxI0LMYUSMe1MCZ4rCQ6XSwrTGE9gxP
U1RKu3QZd/GXq/8nrQ2MqHwHBjpcnkU32CQDz5hU/Ytv3np7nii9NC1UUthAoGPi
0YqhbIv2lvF5RkQIo9BZqsVDWlwLOLZux5BqqD9+jU9ueVBLZx1XrcjgWLIANtyr
leiD02y+dNCKCghRXZj9LkRgWbGBEhrUUlgDcD5L8FbHa/gLJpzVk2muTumm8Yr9
qM4tu3TS0iwUNxoHcE2s4b+2kWMtSXn+WYArjAa90m98tTWn+jbzubZckiXP7744
/WSPjQ6HCYWX5oc1Tn/exoYIu4ykNZocfwuEWKPLnDkxq9JyDf19CGAIe2GooO2r
jiPWu6JaP+71+NvMZWLR+8e31BUvUFP/thSe4CyzJX/3vDrkdR6gIE7qnhpB5LrH
S8fkeyfdSe2jC250LjsFGRF0LMqAsBCPmgkYZQ2u+R9QXPGCmMszkThP9oEx5mZT
CWmSBlYpmPoGKNlXczMM3WUyltCqHkFDCfuToIZ7b9vIJ3ssQzlx5Pwtdx7MDkLD
rM9G5UKU7CHwtSYy8OQ2yqOAmPkpoTUExsfUv739fsTlcc2HdDnvXeGaBSKhReyB
5O8RXpcePjBLd6jcR53mCNR8KYu8ibmdzzvH2kwqFudnfiieuisGNpEUYe8I/Euc
gjWENt1hanylX08HL2ruWAbPvtAoo/xS6e6rhHornYMHrNt/0bxYpD6odOVZhFNe
0wi4nQDsGQIk6rQSc/5dhrF7AqlhcAg1ynYk+MFwEqISZTWSTZCTMUza/sf3UIGP
q8zrgy57bYHDOHE+kT5dgt57wUQUiToh/p/kUfs9kHIQOXnj0hJqvPiY39621wRf
B2vgAERln9APLeBvL6KvzLBQyZkXeSn8Y0p4WzzBiGwmySidKPleThBFsyfg0/eU
+byDyRlGACTrTC/TfafhKokrPHjmlwoPiKZM6f6dLAaAFbaiRlLG9kTeUlyRICQP
Fvrhl0D2ajHJKk44CfWpCuySjr7u//VAxLwmg0ittxHkVkZ1xyRBRx1nYWJ3ae/V
YGz32y+PzDi3RqKIVf1kveqhN2CaOUW61pRcWjZ4lT3K11rxlm0yMs4YOaPz92tD
NLt53qWs13+GGveBpz+7KXF1GlCfkmJMYOBDUmeQcpJ1PljmU7lNAJXaQm8xLXke
t2GTzT/KQZQouSn4BKkGqHd5YlVBZ4pNTv6qdiQLb+1VisndqVLhcUEZPhSVfZMR
GUrTULblLAfpTPBCGybNgKm4Oa713F3FIAuSS3IaDtw8AtGdkdT0o8nlCrDxDSbv
Q8uMhd9gU3xJx5TL+QdthgYoRR5uQTlV2izY9gz9e9z5XAepRVafuySCrwiid20d
sscP6VJhpSltzHLgDeyRpieCTxNJiG+947dPWDVj+espLHDo9DG5CbafmWNEg8Cu
6JKYT1Tmtj0rOe5xDGY35KA0J50u12a7EoM7v+6bfTaQoS/uSXSlMhOjvrzhe02l
DDShnJGVZzPkImJeD+evLrspB4RMWdZRLSRym5GqkXZ3XKvip1pMllvOEvOhzDfo
HvOvQss1iFCcnZvpl53wDMjK6b+KpXV9DI2buENAxE0yRFdR09cAZsYbOgLsgI/M
PXScj8QQkXmtb6wNCzL31SmI+auTJ0Dud5nRdfBV7jMAU2W4PMYLYPFw3QgFrvsz
D5aoI1g1/d6QvUvSp/0JxFAFQtrGUX0A6twWZFFZCIVFZSV5DEPwIx4qvvCa71Th
4pbV/pFUYBIbgHEB3a5U1VBHRGmrqQpNjBry0/dWZ7vqged9Bj5CYtwRwxQgljqM
CRqhPUc+Y1SfkS2ir2s+zY/q4mGDp/zxEfUs3GRDPn8S/YYcL5tSMV4dS+voHkh4
roaa/SzLfd0jmRAeT09TolP1iq2qTnnXmh7eqFvso99sMictrnzV2cUuNtQGosaD
1aNjjXj5Miig9+IkDMmRet+lkKruQaALucARJqbRXWknJpzkeF1woX74OCQ8V9bv
qEUxYEYJpcBmhiKbKHdWSUu4Q4hazpHT/yy7DB8eZO923+xQSnhx+NvWsV/GGUa6
Qs+qC2c24dFwnLr9XAIHulELC8o6HudEKxdVEWvI29L5difAYk8/wDX4e/xbUhDH
HF0jRoVqOeTnrCPaOp440FL2vF2QdCE64nr5VGaLZMahwV9yZFRdjTHIgVA5WZRW
OeY6hvI+TMngVWyP0pP2wYig25WHbigJZ7bpU5m7DGu+8fR3p3P3O3DY/UAD7mPs
o49uxlHO0Tux5zoMN5EHmTj9QYpteNsYA+KGrP4yw0t3vPdRg2e5m+z3sgF8zqM9
/M9cjNXLQn2kbWb5UJVZbLNW/ARV3qnkEwgjcsq2T0eGRHchcVJM30rEchvaa7oc
wYaQQYDKG7JXN0mR7N6a2Ss/cfPKFNUT4u2J4UZJ+tPUnyNAD/owauxtDOy5rszi
BVNJsI2H43k7VME/SV3GMarlEnoksGAzgVpAr2tWhxl8asL0qW0SdIUrM/O7P67N
Ge2LEJqgNTrdbQn3qpFs9PxGK8uGBaKps6vz8zRvIBEFtg51XWCcJsyh3Cb6oH+m
MTpxf2CAItA8m62ZXuNIRqXsXpTKqlL8NTfZ4FjNMspnX0nWjH+iQjZCy2Ntwno6
45qeLM4VHjloCLuMEsshkIW1yWb4S8JWULjeBvh39ZT478d7+dnNJl8J6fxDasQm
5g58dWVJHOUEV8s8b2gxAWdIJ51rg+tTAT9eJ/xLGILBtMG1fTG2JkkOoz1GO0i1
Tlkq+079KNFDrsjt2jlBLqD1mpYEVqBpRNDWHznEn4TAWKwJDW9pPFYNPphuvM8X
HN2HjG7T9UeT7fszuNn6CfuOfmERAtyTzZ12+vYBuCE0ZVtfhXBF4bO9lOsoKAnJ
t9uVGSQcbin4t5gLNjZY2b77+WwbbuJMzMXCT+nX2gJU+65oOggEiX2/yc+f0/J/
9iIwPMZqlMZt0UEZ6AnC2BcEwVqri8w6AFbouaEUgelKO9Eob5ojddKN2axEfO1a
LJhiR1jJNXhyZINFf8KK++5getv+TCSMu8iS7+WboYv7znYEDSWkYN7S2bYl9kpe
VobZu3b1sYiBCJx0TxIFG7tPmU6ivPb9B9EENVAg2m+duBotHg5Z7bu065yrTvUU
RWye++X5HDAO9x8oMIeT9mKZyiuvwVAIiPyWcEf6+EkkttVuhEPamMYiejOTXF9l
gVnpjgg8YlGn9q6Zg51pTl5Rwqd4y+9HkuNWrzDG0JmMMUzHuaXRc/QQhyqh/0bq
Ai8SnqOWyErZppHspyEuRFC/2m7aX6GoYI0XtRMqeaz5s01BASuQozDpAgRaVPYZ
ghCPMJKXtwLt/1sQId8FCJJJuPTHrhc4BPmtE8Di7hYypVV14DJqqBg4EMbF6HYK
NjRzdBOststGpxsVguoqz/Nv5Jc2Wl0wI/HvdIQ5+6mYbq7GxVcMNGqj1VpJtJx8
sy8LVZwhHht5i+iJsj6r9OVor8cVuHckb8NboSkvXATUqNwqMvqiMbO32Pyz1En0
c4Vdatp6+cY9VMeAMDwZUc4Q1uVvWGIRmWNHTltUvBE4BitOE3Lm0uyY/z/iv+A1
gi7MD0uCEKTeOTjqFt2DZjABU4A4UOIN61DyW13rX68snOXU8LwZMjmv0jOrwhYk
/DBneZkbooo0fQiFIzmjMMN4mNECKbCy9ebGIsNYaCzq8W3O5XKYmMXx48TjZY0c
/SZm23XDtW+vroMwRJkPn98JFcIba8eWAi4fe5d3IESqKJ1S8Ru6MOnI/xrKcxc3
Jtqn/HA/pX1V6vpDl2p6hSOeRr3veN1kINYTOlmAUiYtJ8KlTXcN8Gi2FO9Y+8yd
k8/EEA3At4VY4/GAbp/6B95o+9GlwN0pT0dbrtIY1ZF+RULxPa/9Q/RurGcJXtsg
f+g1jkMtUCUIYRm14qmN2YnT+pwgeSAahbSiE+9CvtR5/SL4wZg4tVNvh15QYvWb
FW+TSq6Ix5bdv0lgSPJFKgHRKDAwNlOieah6Sx5ziw+3uH+VP4/BuXyCsmYWf8pw
cCgPdiJiQgvE0XO1Z7t3+H+mU8F/lyKuH8lKe/wEbpFd/topwbWCBmT0lDar/GVO
8wLvQyy7xP+6w2itSeHJzrzYFdYAaj2fABo19CHfPEDfgeJFG1TlfROm+Vfaxhp3
LA6xU/lRkxC6Whaif/jc+SuHcCPm+igAZwN0A45Hk4LLLfBOAQJ3+yn2meGkcK0N
0qLiMEWfG6YS5HiE1bE96XvfBqU0WPwCYYvn0rArOK8G/JMW6vu+uezheJTa2Ktg
qyrZOQQAyqLn7mM0aCHO/i6W7fDoiM2AyjR2a4YB41qOr4WMSQN6FijNTl6th3h2
V3adf9my94e3vt8rW2HtLcKa3mykH0Se5InH3IoWpZlqk5T3kXxWfUYMTJklNxPL
uLVTlYp/XvJzVhTWo96JXrKeaQ9DA6PnEqRHQH/GkMPVWSbZDIht+Wgw4XmhLIuY
0TQ6XnFTo2XP5wnJohcUIq203/t/KAH7NgJFtSpbpeiqknz6nEN+Ye/7fuH5S6NY
3ofluo5uJXQsgiyW9GXQ8vTaUAVXslGS6qKf7aJtYzfajjOTughfzmjbG/0zIkrz
yn3rzbahFcYjaNV9v6MZC/p0HHK7CtEREUNxwf65uumna4DGOCwX29t/0J+ts6LS
VWmyWQUkVUp/jbRzff+4XZ5DIHN4O62/vU/dE+wH5WbCk3w5qijdSdmp/Iq2oBbU
acl5z4oTiYRjj9fUWf3ceGkcBawUM7KPD3VLcL445XIdhy5iSmrFZHGLQOTzg/YQ
5D00Bp8iEQP+6bAljVe9ddUCjQWmyekBlQGO/9mn3c3fnnJytDyr36xp1YNn/2+F
W7sGOJZlnGYW+qv5J+fH+r8x/xLOpdP46/x4Ccu0fDAzMGnzs13LMqqr7vYEKbwz
HORbXmAKfUzXBPSv94/OijKubsh456vNQOGPy5DJDfGkBYOsbSkJZDSyJgBLC8lX
ROmXfQSJMZRMjjXOiy/XDRE51pKQaAPrpnm8KAj7BdsNQ59Kn8w1XflWqIyQ7+5t
vL8+3TroJFoXtVVx5NjCAg9paUGykHXjubY+A1/NX2UC/RzQA1XNxwjTUt0UVoDT
Nj/sBTGpjbKU9AnCdViR7IFEst5fOsDqKwCxuk2UCmzop/zJ2ahw5Gk0q35xuZFn
DP4/e9250RU7oKK1mTzh13oUBtrjxh9n6j+rLZ05Q6pPnjion18dliOFSjwpomJ+
0UcgBpu2CiM/BBKWVndqC1tiQaAPtOWgTaEuGa7I2QROlZq9lzXT4CoiRImpyN2q
9eb2M3cegUwt5xrFsApnte+q/5jJGm1PCrZ3uswzAPFB22ayR5K5BxPk2wwU58an
NhJbLEUs8Y5/qqmuHtUp6pIC4EF4JUlUqWSmLUqQtgtVNPs58xFueto9ZZ0Oq9wd
XPn/DIdeR9Q9Y8lPrPMXOxR4E8Z5fYCuQkB59J/NaaDSfj5EB+WDbQHdQRbrUv7O
b2aqXr9g2OS0Jq0D9qByO3ag2bSKvGuRxr+ND20o+95yP/kaOxqsVJxZXoftpz3W
E/RbmNriLRVhJl4v0qHmjF3xIgGmul5+13VEIpqSvwMMdEGSVdEEoUBt+YGKSjGR
0/3a9EsB4sRHknTwGINsQ8SnJb6czyqPY1dLq7LNqKG2yZq5eK5BoDjhDMFK3ifs
mmwoYkAMjuVEA+QnMA6tG5mXoDn7Xdgyn3LsTRgwqLpyQ004fXozDr2K7ngwjsYO
xrvKTtXWjN7O/q/V8YVrbk5rXJmyIxMuDERuOdKJA9WLKVqhmCN73FfYwmb5LqEQ
Z3nHU3k8ciSBNMckjbqgXcZIaj3BViyOf9vLQMSkASHli0W3vuP2iSR3dd2Ls1RR
RbM21/VfDa3b+O5OiqwFgfqMXg0+t17bJTKitXiyu/lvtOxPCzR7/8L4y5MWGzHf
gCrzSjH1qhGPvknFReS3U4ewScepSVOQg1RmwXHgd3Ag0ZZ4vBSNj7Iz7S3MLbKR
XteFtbRETwUD9G9LaVmLg4YgVhYuU+hqmMEX6J1lmFVU8g3ajED66kYP2yK4meii
O8N32MQtSji31Z/cPGgNsbmuwgL7gbVp61XZhVFajddCtRoLLXncMFuG/JQBQTHo
u+Yo4c3D6ZQBGPUhvY7LAVFEX5O48xbRFBiWeIccSXjM5eZt/jZwpH67X1Hm0O1e
igWPd3qddIskEBK+09/AuL0HEdf+1LsBws9yNMPhck8RybOGt7IAT09Id0SteJ/B
TRsRDIvURJcnc4gXXqOH7uYkKPbVGShHjhyPuyxcPc9VImVDX0h7Qd/YYAyakD54
0CWZI8LCBAYO9ml+qbDEW1uH+E7qSQ81NeEDV99UOIu0l+ZufBq3OkaUsGmDIa2d
HtSIemxomWP/FfPkfAAHhvRLPGHbG4NIEfgbn16dTPK4ifsmUKzzra7r3PdMsYOa
YzoCpzl5zxt/B93EDHA+lA24svpexTodKZW1rrxAUZ3GgSbI69wVqHAARzPRei0D
WEYyIL+9BhMuqmGQR/bIXM9T+QhcKIQTUEBzYDW8JzR6rWX1Oh9dC0qcC8AIT/Gp
Kg4IA4hABe1YLTl4f1mNP0fgtDh4TC+rdKJtzE+dd9EWSIuZ75zox/aYW/Lo0NkP
rtYtNCDWK511gcIK8Nmm252VGTGb+2jiqFzSLXX1YT/d+ctzHP1nDNKFIBzDHNiL
5K/LIdGUztr8RxO9whkia0F8N9dqYvSCZwacvZHNefAVfXC4uwzlEtx+3OuvukuR
Ya+OhDIyHJde5gLV2oJU14Y88BSJMkO6rtE8PjjH4c32lm5C5enCgL52dutaI9P9
7lw3wOEuMNl86NjXeUjFInWwBHdQW35vg/YIsSouxgi7YR1pn6G3TlLcpgAdRgHI
39Wo+IfAZQcl0RFMzLBwW7rWLlYV+DXTGj85yDoAf05+32InffXVSaNKQ5Rght11
6HtWbL9ksrE4YLv0IyNuLTcBDTUac7ILZhH4mAG6ZkMYLHh7Ah7wQwBN5sq/Qr9p
IT7jXv/yMBX7eEaCPxX08MZ5tk7kwEWFfPg/tk2WEYtaI6KHdCycqTTe8fcqAscE
2ZqQjIja33GaegJ8onWnGN9tUrKAGt6x4odFQYJlSsPKgo/qMZuDFDmqv//D1AvU
ouCvu6xuMahhnKy6N1J/28G7gotq6PiiPo5TgrYTGzE6jmz2rLrQ1Rgacvrfa9tD
LUSg3JYKo0yWMb7Zd7tRhzeC8KWtDbQnrQvKS8GzV/s2WmzvJTYK4QiWk+cJRxlt
kxMqVqzNtV71P2G6XsFDXphp2ZEwdMVgEoFLnVkhLPl6DRcMCo5exsGSU6j3mNtM
Isz8pKJjQMDMMycpA3aVyQwFMX1HmWFY2qHRpnnyuLlQh1AfKUoTw7WodvSWy+xA
dizh0V+mHxrLWX5hm06+3uwqAbhXSrIDHvtk7bYZm5PjKhWISon2zxJ0JjvOTHDa
l9d24pUBSwGQnra4zcC2Chb1n6CqAuztCPkiCooWelmzoH37ZHZCrjV3j/nE1f73
MPlFALQlZdKLYj2FvRD5kuVQZs4yd27ibXTcToOyAlPr6cEvp1FrTPuhKVlXk7G4
cSPg9RKIUWS+uqcC+/EK6UyMZ9SerUa8YwEZPThaGI5byTWxT+Eh+s2iJzNDoMOV
McIZuId+Kn0oX7qFLVonkl0RuR2tM7O4PTO9Ys44FqtYtQo5gIc8gp+fgOYdW7dT
eduhYCLbeEwMZW0LeQj8ZBZeXwBoPHYvnydodKERLYoCeYNawDDEG9gxf05TlI5c
1zzeJhxu/2DbUpiLw7VgSt1U1EoyPIxUlgRUJQ4VEWjoGsoA5+qoeLXqoH3g1eJ3
3MoyNYw+5C0TD/S1F0pI7JCzt7b68DMrMfSw9DPskwVdl1I+DwdTFfQ7P1jUOMne
RyrVfb2kVuXXe2rLeerxfzkPnNFt7iD4DFI0JXa5/nIk2uGzy896b0ChLw9AwgSR
uRMTEW6Hk1DwsiUTWlLQl4k3lnm+8Uzn+6VvQsCGaIUEga9uNFCH3S1MekjFJt04
oEWLoP4E1w9pap3Qpq7fxf40iM0RF5N4lqTj5w+8Pp8w4Pre+uXnq0aptHBPXAz9
7aTmzaE5dQWKaBcX2QGIVaRJnS68ng5heKm6yakiwgZb4HTFhOvj62fIfT/G7IU9
yrupGBzOQfgeXEvdqaMNk8cQIQJUq9gD8oIpuTQHWjCb6+P4LX00XVRkCa3PVRgP
+/cgWLBdhM3QZXJntkB4jpN5jAOHuRO5jfHtGRfj8JmQqGqN7j5XAhZ+aVeZh5Pa
1WV8QFW8cUfRHuIp/A90YsQ8hAXcShPBv9/KE48WSkGGYcdzPtlS97e8pTI0rTw8
VmWwSEwNOJXDv0NyUUPh80s6+Yu/MQapRIxm1BnJ/VQcSgzqYWFV97Sx/sSIyeco
W3GB2ShIw2Nq6VGBtdhazfKjpTFwb3DbRrcjCnn+w0lYjMv3oxRAfL/wD7OOxwKM
pQKmfcSO7VCCTYOHOwBmKRc0lW5ZOM2oUSaxSKg2redBHTNnMs/hFSCIDylkzTEc
qLT+ik/8UXj4S0NCPfILw5sy7/ZEYJ4iuTnLImDRWBWbKYwf7eUYuwJHqNUakQUG
NC7tDVgQvg8HruShw6wC/FDtZJBsq4uoKM4qCCWB8FzXAGcd9zCoy6PDzYRTr6jA
eWWIMxaURA9Y+RFtnzEZdB3q/hsGrE2Wz9xe4XVFdlRtRyjxd25yMjcm7E00EKMb
kD0THTqbezZhp0G6HOj+Npzl2tP6/mh4pb7LoRSXLhrJiagHOSY0BRKR4XAyFt3F
yebefANMJ6Ki0i6QCQg7ZWCGqYeTyyEHajdVb+vjwNIqnBnc/1nM9G4bXo2+/fu1
TVbXcIu0U7NvgsHbM7L0YJ40EsT8/S2rXbq0QOmMzzDemKeCwRgHH63w1dT2/y+x
56qC9ucUOauetzlIrhuipTnD/voY/m5gWnJg5mMLEX314btamm8aRBALIjG4ONYJ
huLaXwjWiLa2Io5UWTEvQmdQj76v0rhq6FVN50b6PDFCANi2GT0H+aSagMmTimOB
iQS0qz/itE+dTP0ne4L/yeboAJMYqOw7DitJLfoNkjtMwshAhjCzgFkLGawby5LX
flNziqrCwl7gQumf6+RBYxPdxf4wXNDK4fEpMztMHsrXf5iPuRLYHTQtqhi51K//
ID/+9Mi2oT1yL1iapbbC4pZpZeJ0Ct8mVUbnbiWYcIkF1oRCJ1tmDmCzFOJLZHsl
p4Y4gm9gjeSeNI5KRvm30VyXAa0Sl22BcSKd8LPGV5zaV6gW8GAcDu0/M7B+Qa3w
mc4aQptQaDYWo6Di4FG9OhgJ9XSp7aipohYvVE1ewrYkhwL1FsXuFFJBJAaAaGM8
jLBDXAW+tGVlyBgsDMDkjxqVJlOTIIkZkHjw7k2SO7bYuxcnTopm4TxWKpjFAluY
OvrMgyWZDuPB/u606RSgjItIW67SzTVr7uxDPVXspH9Z3MpC50JZhv07lvsyKwHI
N+x1/RpH82YE0ESIFrH/3m40V596lUH/IW9KV0RYP1fJurrUe7HyZTiCL7s3iEbZ
3zmH7VN0JGncPPycQLGLw+yGT0+jpr/Cdw0ypmJAtvrUqx6D6f5nCe+pQh5BmiHK
u437j1GkrU6FRe0LKUOJ5B4/tpTcMsW5Z9CWU3Ii4J/Sp3uPhLOIHPRMKiUbq/Cd
oQEWlP485XyAfKPm4rwxY8x5RTDstHqcFx9QopUwipqcSPwq+5xueYtqXHJ5tpJw
znpZAlUb3JBR7cPKi43y41FPcbTxPOx7tQ0B6qdGA203ovM8MYFwL1ZW6diMh50A
LCsFnFTsWxl0kSi07kNcDPcisT360+bOMTPc1SMddc4KnLkQa8LGA//PoVfqn08A
A91k+H5/XUUMOtmGb6XTUsU4+gZQS1+rIhHGxvwL/jKXpHwOFNMlilnEuCwj3yyJ
Vxv+MQ4A00b7KEwFMytvMftpbPrb6rhiaBTOVEyjKUWxQShnKIYaGpGVaNuxQfTD
0NjbXkOxl2aDpaoRdPjKwMYgLt4Bw4WY8eajfuMIkj1eSPvbxBDytvqMvZxbFt5g
B7S2Gpi+xAMvn8HEWIfVWSwzQGGjj9+W7ab6U2PsTYmECpOIKwUgmVHk4JKQqOhH
CHUj3v07MpMXD0b+40yZED/lg3mWFH57W3Wvt8HOeUDf/Eg41CtJGmZuw4ghZn6d
i2zx0q2GMIvbrAK9minkq5feuH9ZMRfDaQnloc46LKEsPW1yTlDq/DOE8v4/TlTf
0gHDXjLVBV2jqgUPz/b3Q4E+gtfRwMD8EbCtc5Xok28VtaXWkQw/fVDY4WmKIgX1
0THaw588eGUy6OaYdwF1qy0W6U/jwJWCfswIn2h5NzP4dC+zcaggZ2Po4GBS7nqi
sp4xU6TY0IdfAdpVYR0EA0gseSrakMzSo1DAk5YosqrrnEZ7G+LgwRupAqc32MZO
gpGcHgKpnSPiZjy2IwqrEXvMQJNXZ58qcJX0y2fmFlrzHKf9eQjiQOHji8DRJ/E6
0I04EDUWu84lGAddf2M///0CU+p0w8V0EP9DBO01maN8ZNvURocsfmOEzF1ZMlEu
aXf64nowFDxMKEM/U3b6t6NZWPHmq1OaHQBxnkBc82ZJRrrzkTCTwKg6pIKljWPV
4QLEirO5Ayq4FZm8mIRngxU1+NLU0rEndtzPTCgkVQVyGzNJuAGj71XH3/Y4i3rM
Q+sNYt88lHdGJxCSHbjmA6mWPpwXgGnOAdmZR2MpPcYKuJ5U1fqAlS/l1ukAc7E/
svnkbrl9UoOqqtYmPiP7uTUwWxQR8Q7wXJJx4oKSA23BEddplRUkksDILxnNu1i6
tl1L4LAr36inft0zASCXo2D49RX/KH49K47FFRi40dimpFBsQEhlYt0wZ/vBeOFi
7/xjOoLfHRqVsizsN3nIIjJ9Q5AX1Yxsr7/8e2sUXFuDg69lgMNh4Mc1dA1pVQbV
CZU0AUtd4UfwR0taeC2Hlh4ZOk+rfEcoCfIwCSI5ZGAE/EOgaBH6lRAZcUV//uwB
D4Zpw07seEui6sjgkTPV25wc0INV4JOD1yGE6edhR/kCstIJ2w1EgHndRBY1Pc7e
fIIn6UQV47NxqN44gps2IBjuJ1FDQqgDPsKmsIo8nPPJ1bJbVSMaav9CfD8H3WhK
oiiaBcEKWgpvgugTnFGWdb18TrgXs5mGaeHIuq71IT0Pi8x3WJGhZXqX7iMbYXSz
lVjlo6FwbZ/JWwCA/i1oNXqYLNAjDpXNamltmsgNB6ZQe8w3rvqsF/8NQDhNueLR
PEhDDyRHCx27Jt4sO1nQIwZoo0aHI/1/nfZzYZMTHU6OCsjnLXAQAZODmXYfzW/i
0pD6PqZStAh6DDbsgUeJB66QJZlSWo6WiQ1ydVKRYcYNM7IcTrCvOwdThCHZjHwg
Hl09YHO0t+ptFMV/Ob7yFuQc+aao9hDlHk1Z87BOwuKrrhiuisOfLDyd6IUurp44
bh8gEIfDZcoR1rys7956WC/Gt3B7jZa5Jz6C23I1PZtjAVZboSBWFd2fVJSUdCjD
6TAG7YGPcYvGRzR5jQLrD5U1iyXBp4rLLN+V3ErGCVC8t/5C8CInFvQSwqHlV6xH
32sFaDo3qzQlK0DTNgLwj+yS5xoaL3bRy8RzSC7+6DDWEEjI702zYonqJlQX+lfb
MvVbRHZPEx6iHB5+o5JRPOE4s7wzXLfkDinRvWnSmHbVSW54r5vQMvLQaGTnOZnE
2PGtpW91Q07XrQUdLUjFdJE6w1h2zdkJWkhAxaC+p4JVRm5IJiPAwEJsOrL10W4Q
4K4NUSOn2+5v7mlxtU3HmpP5TvymoGfF7PKgcyvw8c+t2gEs+NSJxpO7eyY/E1k2
SjYLMELpSBvxDBrZOJoGvSJKIISkNWL4n8kf3NdzpGYySQ/DBQJHjum51L6x3MiN
mxHhZfvsNnwt1dvxsU/8CrVw65gBpqawGg0cN81BSKZa3+E7h98WAefB1LK727b3
4diOOJLqgD1mBb7YjXW5E+Veqhk9RwUDzB5Ax6jjCIzdg5mZE5WaL7llRlT7SDFl
8V1Uz3KPJyS7QVxlmS+BrAU6Pssy5K9c9erTPkKC6Xn/qAsHqHn+WIrk9ATgj2zb
GClooBiGTG8VdKDTbXeUzuvlmNSbPX+jhbjjCjwOMKMCpxgF4lZsxAzbLtliMCrY
SCZdLpUK0g9PHo0FsDpJdAUU2xWuph2dvMwk+Jq/DUb7RuFC0oduUgHHgDVPg7wE
ar/f18B1w/7XoU49RK4vhOXptCE0Sk1OigWymEYmnUGlBGFHa9O8IthaSG5V3CzK
uSZrOl2cIhBo0UBl44rnzn2jUQbgCXxlXuFmfJ2pToGWnoJXL4fsQBsdKp3euhs/
6CArG9BcDxY5u9NtLon6gkNLZupIMzsYGxR/L/NSUq72I4CcJQSWqVPef29rphVf
4eenu79ZH/vhKqnIeBYaI3HtwzDFqP19IICUUUK7ADg15o8HLXhpnL86LIpsGI6T
9OMRF40SSFltZ5qoJbDF2A94s2wlFKmNmwiqGB8mFzVZweFbPch9VydD6u6Kbvrg
sJupW+dioJazV/KvxyWUNsrZlr0Yqxxf6hZ92JVQiwCZGVP8ei/Y0j/1EEtoWbzQ
yAw60B8wiFiSyhUV7jdjYVGOtwFl8jnI/eeR7eqYUT2wfbgw/fVJ871LEs+WEIaK
zbZtN8ytwuPpE+anXFYklkBzbcGX+kft2VnIY6K3uj/2nxi40ssTLisCs1739RZ3
Jbqoe8kSsq8pR+9txUDNwpaQwNG3iul7eLmI7qJD7ggbxOzBJqGnojRwCeZH5gSV
T2IHLtHye4Lc4zeNs3MuWoMCAsZB3GQ0SwILBrhiZwuXNuIF6MGfVeN7Gfs7yaTp
LMDCq8TR9FYPgjDsTU4NiaLJYGIRFy8e3/dqgchBwJlC7C0rXZONyEDV5UNXmLpE
ah+MeB8fSE9DgzL8PfwaB6if06J0EzwpbGb3hkAp23HEcK4WslEPbozC01KdlTdg
emT5gccjG2l8+9/c73LFFHyMaGXWzETpuMns9Hf6TUjhOifez+Yl4lKJGrABASnh
4fb6hXHDKe5JYroWP/5Npg6o7+p9ZeBIAuaHRZCgt4sxev7Q/bXqDJWfYJ6f70A5
SnP5P/pcOGcBZu8V9ts4SkIu+iV6cPbMEg3gkKgncPWUHqJfypLFtlb1fnX+Pn4E
aSggWXt9SsMbTM2Yrg2c23Oqya4kmt2GXpc+s1qjRtyzgLKp8wscut40Gk9hQhm3
D/g3iXuMxnFKDbFSNFz5t6AjC6gd4LBQFIwr2EoREkKYlJ+CnJenULzrzD0pIr1M
NaDaskfdsgq++lq2CSbK4dPQ5KihxvmDHS1S/HW/jNdNor4Sn3PwH1mVi6Fs6TAL
A+Isegt25bjIe7Vo+N8tKIht5jyC1MWwlDz/7LoeFkz91nkZtWCcvmEaVEMevigl
hFPjWVeL0aNzlyU9OGOoCjNnqPkfslGCYalTpH3kfZxiWwLRNd0k03V4eb4MCgbu
si6PlYMgqLgJk3menVuPN+BJ8wXyblKcS5BBSjZHv+j1gug8mKiH21/DSnW1bbd+
tcGEVpxQmGBO8coDlAANtfaCVQXzKV7juCMBhnUtfLWEbk85oFI5gEaCKIgaqzjt
vqEGgU0MO0XM9sTl66XCUZMOQJmHBNfbejMeHvYg84rSrJhjp/bN5Xhm/Sxc2xaI
PToSkAKOhGo6VJGL3wLOrqXWIWLcKDbtUbEvod2VlXk4OnP+wasTHeGJFeQFJkyN
tFs0WFyTMr2QVoPzHYMIZS/FzVM0HlE7QyRJMFQFWwZhGM3izIhkQpeMSKxgrCyF
nOJE46NfdgxWacFdvYHf8e+BlHJtPPoZ40lhYAQRJUCHyj+//xtbZfab8dS6RMob
lz2Vo15R1UNAbu5ggzBbVbO/qh1bJGhmT+NrH0YEx+i5J/TZguOZSXELRSe9XxvY
jyI7ZXEfp8ZQ6zV/dSriTEKD5Wc/G+TVD4Gso01U40nJ3r6bAqpmyt3gJ+gP8Zow
XM+1hDo7YdBfbLAElX7J257qOaO1vzp76Qctvle6KqVu+yXWG8o2tsHGQdJqeC78
NQefi47PrglA2iJJK82oE/hAmAaSs8XsNVkisqLxTBk/DBNUY49bqyX+t1eak38Q
m3TY3j5zeaDqnfwnpP7B3yU2LMSrcr2mWYMP1ACTosbh+bIdZxsAUkmxTCdtBYWi
3q+DnkASBQsYG1O4+H/HkHDJQ3jRmdMxvtM8ViUlMfLCBkglztTAP1UU63tPyGWt
LWtJoxpOQKvKJopxb2bfnAFa2kzCsvZZPU71N9G5RSBewJX+zMad+VEKaKeFIl/j
h2NxP5xTG+G9v+YkzqufQOFqhDHQKM9H74ahbZXgNprdY+Ygp5zlTXClAo12iJfU
Y5zKJU83+Uh6ubHQMX+Qo/6jPejm0nmcFA1AEFEaK+k50RzkhuF4HImLdDLgZmpt
8wmZjygWRUZe0my3znC4FsPnTdlWbxvezGt43RQExINscNcyPlDCoxrrXosifQPm
38YmtBPATCMaf5wX4x75XXCMCB8Jfj0XZA9pgZGTqz5uS6pCYUCWYM4jock/Q75k
uMCGPe0GIG+p4QhtEBg1U623K7vvk9DRRzmvXE11LacNERT6Ugi+SO+yNlRt6OEJ
arP1153UGQqxIMr4fEyJ1vtmuCOBXZrq/Mqth/MFOc0dpcDMeUSwIXdsQD3483Oo
g4YISU/CN4Yl4scIXb0Nd9DZIiTAUfs8bxIogEWZ1qN41myFDShPz3QPM4/DLSkZ
N5glIwnCymVLqdfEvAe8HUyB08MY2VgrTlbdt6wAWx/NUcIZyzZE8kyWG4woRSGz
AYOnt7MyOS4IgTAaTDo34zy0Gj3s6EKBQwr6vvGnBVtIarXQYxFJoN7rQ8WqKaf/
wBTBzRAM7ffgY+fnSK3eVceYhv+++7Mzg3agNcCY79BWMSIq9b4x2TU5LaAG1ZiN
rTHuLJj/nlQWIsMRqjgcD5jT2s5KJXxuU9tyzvM74L6R4SQ22nnKexJmzaAvk+lG
2ZkWs/IZUtcL4IMO985EArtXlE4FaHBXUepxaZfv6cxVKaEWG6cFHbUArrnb34Hw
pWj9EyUyuY3zaExRuNuhcixJq67AxqoKR05k/lbr++V6wLsTi1aQIKJLl8PokWPi
Sb7DcfHhYBgMB+Zlkfr+wJt/JEN2OLiWtHwdu+5efAC6i9Y5tcjY+MG6CpYfpteJ
P9am/y6AOBJq3CWB411TYBUKfMOwsxCz8smi26Yb3mdloHlAx4emAYMIizcf8ACE
0JuyGltBre4GpQxsgkZ8nWMgNC6IP/2olFqmolZ6HJ+H4aOWsIvozeLsifg8NnLL
amvbq91/44KzlGyMzN2e205CbwWMDRpLCfAK3BHT4b003DGoZc8UgidHMuhhKxqG
vlNzDiXauOBiuVbAtmCxilom26/VnDt7iLHC3qBsn6YJlsAlt2TuqqUxtHo1CuKY
ncTFfY9AY2bUgsvhH2aantTm9KLebcGJ9O9+2UnIos882H/0xfOyG6gkWORmDNYQ
I6wq4ZrPP5BL8C9Ogkh6j5cu2hYsiCHn19hO3HZVnAW/+7UM8K01zgDf3kUmCakk
3lz89iC0U8QX3boAmrf8WaMJaStD6GbAjlI/f4+a1Y9Q9CbmwEqmzGGahFoMaQYQ
AczPEuRh5C+9uxTpw9PVMu1y4IvCazLvSLUBFEvLxR2p3u/BEkFKg7N5DyX2ILNu
N62AFFP9rgJXOflFLDp231NZ1CQXBcxJsRAl4SCiqgdbTLtDnbJIDr8domDYL9AW
Fx23YfDYYmF3cFzZhMKrD7iVeE1NGv8tTS8uCgFkknr2VCdKB27d7H7CLZ/UFrmc
8hOewGWVrkj2zuTkWPyxV5unhSd43KLfRsbdKYy9jc8l4JVHHSH/t5EV/aPJsrAF
MGLV+v+NkBgt7YcKZIjZ5P9RgIIai09AO6SzGuXeiLDySaEP07JwTZwHf7u1RW+R
0wIUW/dcRt62S+mfCxjSyQ1rdIaOG3c2MAS0DZl7PsgdKJ3HqX4eWtfVzWzOHNk4
yFd417KCIGo04HiNJbFjh5MPLOfFFtheo/CVpdEWWWIsUzFteog2qryVtGETvcv3
9vAF/daK5XbaFPXtBGDw4OBZTCxWDYUsEwZS96Sb1iHvtli9lm73+v+BB4Z1O00i
IOIbygrgAgmYtWqgqSwekLlr7rgPSw965i7E9EeAdaJCDt+mZus5Tg74xIgIDXUY
VQ3uJ/4hKdhb4Hub6XWDV4vTcgSEo7bwHYNOdBObqDCGRfgdN1KfosHCdi+k6Gwe
ZdI1tt1TDXX54BkSX6mO5RePy7aJ9dDdam+v50N/kOfeSTDmLwamcXxgfezwxC9e
HamaH8ZETk/l1gnMb0BR7AsraD29SMCY+4A0RZwXLeEEVN/sGYEmTg6GQd6j7KTY
ZU4yT03Z5SQUQptNQwzHFbfL8ZwWA+rotwl3YJYC9qOGnZFYWdMbb5n6shuPpRad
UuFSV4G1L5we8OgFazXiVFSzrvHMb6i5HJF+jFMID+OYazmvwH90BsyBcAdrj0e9
v7K2cdqploSJvzcjOHqoCdYTEHxcd5oroBJN6/9JQaYWqndYhOwR0EswxUC/5NlV
HWw0p7xDYcbapGPMNlIGkC7XOSrAcBs7iWDBS/+cIgIPY69I1M6WkczK72zMNGPm
w/r0xo+wOH5ELfFZAl544AoB9AjZrQNAJ7EGkYsVw6Awhqdb8MOVTIKSqDDqZ9tV
4R8mtiSzaekWyxhStSKQeOZsAD04GZ4Jq4QocsNl8Og/nmFs2DJwoQPfTdVcWuom
6XXXGHSSgNkfrJugLWL7mimQh1byAi0LE6x0phXCG8CHeTT96l/IX8OMrn8H26wg
xdAqUqqFYWImdbI5qlBis4GmdBvUXDFGPCvf17uDYEP8M00k56LF5bJbMKvD4Y7q
Nxf/K80Mc1UXahWY0ofcHcgEKbkAMX78X+dF1X7rKF7u1uU1++MKxmG7KmDx6W5K
KzxYPcCjV+c7TKZ0sqL28CCHB+AIQIlAe/TKolKe7b1AOMGrV2DbSIl5pLLFiAUl
QrJsAAchnLFQaIAmXQsHirVSo0dAWGdxbgHyJSX9pmSQCWXLqrog73R22aiyHP7H
VFFCCVuwJmjwEjD7dwIRE2pMNxTyJhvG64nTUHBNM7ovU4sGaVoA5Gi5qLPdxwKL
zpFa4qBStvzIAW5SW8zrb7USXM8Lsj8SONVFfd8eJcXmNlfKKAqcT5XY3SG6R1YK
pWaX6+cboas7cSGXLYvkBeaKIzi7qIy7o7B7rvJkHfkTvWM2UVLTmPzdyiqF7NyP
V8iJzmtU7yQDdeINe9ElpWEpB+eB/fW2G5UKSKkAHLnfqhQ9BsmNztcGdWxL5Cru
nrM5sWZL0ZARpicml9gkRHGtXONWhGBWo+4NFbrFiHF9+e8D8YbBBmSnAs0ucsBP
BLj2Xun7DI156eZFoUQ5xK9AepUW9G8J5ZRRNv9jxtkmxsZ28Od363XQ930M19PO
8VMyFvijFcO+d7BM6l3aABqP8Mkw/gHiNvoo1+ic5lChK8zOMPDCKpnRKqZmqmFv
29SOQ/KpQiX5HoT3Xg35Y82fILSIniz9SGmxade26G+Upyfb8PAjE7GK1opbHM1O
Mz1tXxjckTTwSS8sDaHR/ePuAGwGvlFy42b0aDm/NP6WHKCPRAd2L1FCntRFCsB1
bzF4Noxmks5Nhg7Z8eteEyOMWBXX7+2lL8o8w2x3pNA3FbeY0Xxf8GcJWA4Zh7ym
2XwQCzJteTTMcaXAS7jUdVkjRN0jdwBXrMSZpttGk1T0/pIzu66H9oX/86MFdFWG
2sZrKNDtyCm/M7IcIgURSwsW7OW6Lf+OY9if76wmTQwhE/2u26FhTQxnmYaNgul0
it+4kLV4ZLW1AKGzLT7SUkSx8cWMSx9TS0pDlZvL9+uqGDNyOK5Udf2tPTJtTsR7
7QY84dGwZ/7TqivjVjKTdvtqm2Ja+fBC4hjGgRAP01LYRKP6ix6VvnZ2dXH4lBL3
j0JO9TYDUOWqd8Lf5M4Qv6XmENJQSoMnz5cbRH33WVigA60xV+WB8zhCoBzupaY0
W0CGUesw19/zHBx86TS1egKfbV/Vk5jWTWnYezZvzXylDcWQ6sWiFM9HlHXTq2Rm
HuJ4D9xCo1I6PmQX16EvxgH3gEptCDKdmUS0bXu5pXZOusr6kUFLbsY6NsSxfaB5
2RSg9ByViv675xhhwV5SDTRy0sCwzj9e9/ufCkMJm24Iat1QJAPa6b01oHSzlqkg
PRr06JMVwyUHFVR4sVdJPx/FT2BecvgqqNGK6sO0M4iyEcj24GOryZcx4GENxe9z
HIQfSH8ls4oiMsy8mRQvXJrS+6Ki+KjJFUAEPXmSYpYKMN4udRocAyAwmSEBQNwU
Q7aF5V/M65HAzrTQt+PdMdKNqj+ED0Yw5qIXabg8UrUt17mwLcEzHnfNl/8quABz
mK+qOtKzOPHSE2dUWc+XROVpLU+TPFVT96RfRH7dwXasdKKqWQesuJDJ3Qq275TS
MErhsd8Atoniq8FBf2QxTexfrBHU9dy5BfifZTSEfSmiaJPIz6kkSlJOxNif+Vke
QGF6cGeAZljrhRM15gT6jN8ghUXNYdg3WsBXAGXXOLGjYWfzOqwpzo7jjM8H5ltS
88u2qqgYRmyJ05dnCfA7nZ/OUhVvKyVbB1hqwE7aunuvuenY2CVjpC2Tf1BwpmZR
5NPMVzJyMCqXYoPz11N1olNbq83f1iynzASyxtSkWGzAXpB0sNANj8QiZ04fzEhR
5xN384z2ceSjQeMHu/n/wS7Oxomkk5hgCu/hDO86XsX/+vQAazYH8Uaj6xKhe7yL
Ug8VK8/GhdiokMyuBc0DcXLA4/HhHJu5W8t+8dfRy5zwjc0gLXgJn0g4RPQvSAX7
XrcvNe9YAI1KUSmn5LxWmvJoWPFRYtv1364SXXrmAcZQEjU8eXmZ8inqiAVulkxR
0VioVMSLkeqm9Oo8n/RPKlr6FH/d1lOtChcRWKdAPxwboS1OGeQ121LpmKovXr8+
Gh0MI0oouTrq07gqH115kqzOw0pE198z3D03hGS6IXhre76Mqf4OmZz1xuCkPv9y
kEEc3GJ4J7bcVFdHFJv2iXilB9vDKnTpwDxE4h5T+WshqPjBZl8sdc9Ix38NDuIJ
m9t5ubEoSUV71FlquON+W7iPPqxuZi3I6pK6Oqjo2//7vsvipJSx4bc9VcpoeTel
G1srz/zGrNP8CKf0a0vQkv5Fuc+6/ll2qLf0HWui7U14tx1xHBHUMaVPc9eddmS3
upxi9KwvXf1Am0gTV+ucqBG6SegpZhjPOuZuyLgaF3RkExWExqyNnyxmdp4gMNDS
ZNc62JMkE6niUWhxrud75kx1bQSSK3AHiHd2sEIYPKcKr95DDUgqTe+wmw2GnDto
vI2pKxVg/r6Af+RUpZ0/ENQySkMcMwP2FDS/xFqF5oukeCfbooTEdwjcl18oPXrm
THEa9+Eg9StlFKEBGG8L/qFvV72/RI1nm5LIzhhaR41HiS8bzPvYZ/rrw+fQbn9K
T/j+NJIjbdlAhEOCcfCeyUzywMr1imZRQJ9uJedvQ83wygKY6enliorI9LPsz2So
5XhJfiN1NpJ5cUdZ/3hPfdO1/Ietw5Czerwxnet4qziHNj98Q8Hz2tMeIaEnObDR
ar6/dm0cyUGUj5K2GxLc/WwA/8eP5JNwnZxj01ciX5D528HRsAIQUruMwnIyH7r/
PldQvzOQsnLpx5TdC9+80NUt4Wd2spBECG95Hmx7da6pIL2jxJY/1OCDbHU+Glqx
8f5JWPzchLVPaT55sX70QhS7IfggN+7Q7iu9Qnp1KfWdwv7xLfnM1/rpvTG0Zn+n
W6e2y55cmBq6IN2wbHUVASgFtrJMUzdhIlShUw/XGy4gu+gaKuZhSqoJ8DITnqkB
V3faUswuUbxNNq6c0o4yOAcWDVOL2kEUd0U0RZJkFIa22Xe2SjjTDAcJnG/1Mb3Y
EHjfpow+95qwDPTc6Qr3XdJIoiM+Qd8+wwc4Z3qKdNUvahkPTSH7iEY8cMGF3tvP
TXjA1Dmiqx/e7xIw9OuhMpEnoGfrM5SkabvSgmexafvgxOnzeoSaPIIIrlbrFZug
hwjXGIPIF8qnIjkfu5NF4i0HDfbo4QmTGo+uEdYBp6h6Dutdrv1dhf6VpIkvsbqf
w8aGgwzY3kp2QlBR1WEGvL1eOZkQq9zYi60+5RC85xcBwkTdjt22I1gPxtUJ9rAu
+GxpZpYSjnz6lG/Vas32f3lHB5LUGeks14Xx3klaNlPoV7r9SF7axoQkDiehQqai
LCwH618oCbemmKXTb/OvNXQqfmyTHEysGGHqu/F8FCWwSyrLWdeYdVpkUWfK4rfA
0gTX1O3icI3DpQx5kOgideex2NvvnXAeOz97ks/cLjlOIogKZVi93x1kCGZOIcH3
J5bqswZDatj27gd/SChNwBDTJahoiy0G58YpU9kqLOUT3kglp/VDc0q30eiqDiHl
J3mqUpOKBV8ryFCmNC/o56vfAjPM4kMr/RyZwLvl5ZTVVl306gXtrK1mcjClAsgU
a01EZBMEJDC7+Eqmp3sir5CzE9/flUbcPD4Nk/Z3kQmSRFS5Qkxpb8VnL+L9z65l
Sjk2imfcWObeeJ0bsKcvT2GszFn9fI2B+Hqv3S+0A0gR5/i0mt9k6lGtRId20R2n
q628XL4uF9CbSPvj9qgfkJ3kZvigfFEcOd8dahLGXXvZFFhcmTBAaL//XONaRdSu
yW+pZ472A+UaoTf8r2RwE2c6RPFmC7Zn9qAjTJueHbnoYurBqDn2kYJ2DmV4lfNT
HqpxtilwbfvPmdXFuSxKTEWO3JBxiJ2ExSGnGkhZMQDZxNwE1HmmXf1jkxK++o/G
K07liufUmLORwJyybUzYVCw0MZyBjD01b9mQm0ILIshTCpRlrE2TP9jKDxNPa4Bi
e1HX46h2CMPaY6+EYmLkni35eYBqJ6t4cMi/URIb3hgRm3+D7CG2g+4NH/cWIrd6
H6ls40A37Q2RyV6RymyIhCsTqrx5zESf/d07lPrVZSRVKItWHjKs7NU6l1nH/KNf
fdfHBWMTG+2uSErLcVz/gIziqxFdhYmmqe2fRT8T3fKq8hvx4381P2rK3brPHpGV
vFPFwb6yD7i3TAeqNT27mlcxhJqJjshEQPtwdSTF8bQEpryth0vMVF3XbxhUIRUq
HPRjEQkdrXdpslHC4kIEOJV1t+uPjKqnTWtVP419WFgsNf4X8s6+bwBkoDeMP2K5
KhFdSnULT9vlfQRlx+FNm69aG4yJhm/uwVQP9vijyBXoLZuyTNXGWBMroo1PQRKr
DhgyKTzq6brVKp2FbhmWYwBQd4Vk+GxWoGWHIoRuVvPxABKujLwqMDMps9NOLduD
qHq07/2bIrf/Ng0KZsRteHO70rHf+asDwZ7llI0kN+f/dyqM2lFOL1iYgaveo9Uo
G1UuKidnitSzHisvTSkWjRxxakB0ulGoxahtnA2tTRtTrT1n9nEJFJhdLiKW4TpD
51RCUvL7ykg9e87Shp1cn7b5KH/y9Jb33l+5MZeShhQEQeDi2XhhoH8e2wxTDlNy
ZtW7VXPV/dlL9jkxWzNcNL5P/jPKWmXsinsirEzF+3ccDE7B9CwBS+Elv7nRpFOo
LjcFLxW9tjb+o83oo/xl5NPYVuJez0Q7bXO9+uE/8IZ8LD058DM3KKlZ0PyqrEGh
f3UEbgE2xUSFSDBP8L1CUbqUBp6hOqTbJmpxvbGP2oiuL2nTrkEKGpti3rGKfl93
P3kfRoy16wlVEOR08uEwvw2KA6UGJV0zy7UB+BgfenBlFXmoAQCYfLWlwZZyD4j5
NxvMlq6goM1M2NnaG0b3An7qptmItQmoC7C/5cmyQDh0Vvj9qCIk1oZk5VSfbcQQ
HR/jUcI6Ehx2K/J0jUEOZAP5M/dXDZE9DhvBqjIlVreiGsS/kRxn3PjEWThLfNYa
JPQMjCgFJpyu2red0aXlzUD+NjMZ7qbA2l5WQVppg07entzOARX3z4l3qaKcHvw7
qR6m0QNSg2TXyhErj9gsvdW2wK1GYxX38EfFe2fTWq0uoUUex/dbGV3T8KkK+68x
jHhCNRVO1ukk9jPbcBUXJ0s4O3OqiP0vUpoabqqRFT17UIHabEWD/SFnASL/Knh/
n2wPQlvbfW03UCbnJgLAztjc+SVInysOUhYGvvH099INt8zc1Ch5+A0z21odM8V+
/Di5SWN8hImR2yFCDhZoSqccjcM3dR7AwSXMzCxeWqoC6m+fbPuEmGGTq5gsUK7a
u2XH+x60mkxoXDXU7tCKql+xqdK6//vgzYOO7+cnfveWb3p8WnBpKUocgj7GLzO0
24YYU+t77mYUfzTkX81WI7L9IrZMKWDlT33iW4Cwd96TH6z/UKiYkicFN/5QJGxE
iZj6bJzfsMUKzThv+xdn/vQqq+G7FzbrLNCW/3GvJ0szKCJFzXqiyDFewyQAD176
7qOE2rv+OCpLeheApadtkwYNmSZPQWTDwN9fiipou2pHdEA0YvUVMDaybaLa4tZA
osLHP/VWaxyCC+Ko4yJZ1ZbZaHm4FOsRLIiB7YN+k1p+YG6e19DA5TriQe52muLT
t6vx0eTnSCE0pCQkXuF6F88rn7nxD7YrSwAFfG0WoFEbAkQRTAUpm9wnd1CAUPM6
Y5H4dbMisdBVx1Qr+6+IR5WwmCsJHhOVM7cBAJAxmrmYshUaErvdH3F7+T4dARzU
yBuPYHBzt6+KZrAgmT5kxbZYsDXTHgxRFau4+ESALDK34iqpzMNt6CZjnjpwXXEU
VyXxR3WxYklHYLGCP9G225Yz2l6Jaum1G0eR9+334/8ZPrEpHYWBWNrwNc93RR7u
kTSyeygc/1ZzlAs2ChY5xR5wkvKNd4HNzpOoh428Fb7ysxcRM9rd5uWONkr9H2tI
1wJ5mQtpGjUdpdueStGm7aVJB00rVumVfjlaQ0UKnyHBb31QXxZSSRaNOshHPrXo
rIBSE46HhGZMZNGdZaZAQDMds4bp3hA3geNlrxen7zI3kyiLzmOeOX5sZanl7qJ7
afNqiY1vjqbquZlcRqEbKxGRLNrmZTTC2HgClvpLnd5bG9gb+Q7qglZ6F2V5eiGm
SAZGfQ+/cOu6SGX6vdbhzA8U5Alp9hsmKQHulBEtTklPHszpTQ689qdUzd1QvK9E
dphBfSJgTIk279FVqMZ/T+UtK4mCuU7fQT5FfjMzmaoqiaoEKwjvEQbyADZZw206
pKCG5wXF0I92Krp0rkMD6rPJG7wuC3cU2Yq9uD30hlDcDKSd+sPV92URE2kSpFRS
BjtC6jLuF7rj5726p7S8wgE3y768rvn9CFqT0TLlLfy56pLWjiK3NePzxGpZi925
DUc/10c/h9zQNcvsFzNyEI7t00LOEgHcmB4iB9Xs1RUYQbmgRNm+MfREeYKwZlc7
eUhNGC0dLGH3ukGlFZdgYiaQMRFckJh5mME9prO321GJA0/WVtWfgh6TVG1NCkZB
OIBCdYOMlHTOXX2zSzoXq1w5aQZyseaJkuICOsyf5sONcVBJsomYgzOJ0Ov7Tj3e
s1v7hs8Zvr6oz9MgVEtqrHWEOZFeJhDPrDXo2ro+GcsI8kPPza1st632hAYQ9mdV
s8q1FJUJyjGKUfw4iXyidPZsmSYk1w2P+DoYjJysBkjC9Z6oNL/MFu/AZdlB63oc
ygpjUJBEp+LJeHHCDBFWRJjzU3P7/zI5NBurW5ytNVf9SDJEdAybH9GEb6pha60J
lpLfqFULyPEucj5Wvl8hYG5GzkDIzIccx6wR0uu2K8Lst9lyRUzkRLJcczsSB6fa
s4TnOPzR0eqiVU3Zo/8wE7j2goR7xGY7VIio2/PpGixKUFMMMctPFMOtfhk3R5mH
56xFCO7rM3C+neS/0gK+TNRcrY3joI4hwqBDGAG+pMXj5PHw9pPQKMn7pzTLAJN7
npRjdF/lElT7p/5fX94CIHN53GL40friR9NW/FdbJ2b6caQo6Pyao8N3OYLy32wo
5VriGWNl2flK+XTA7M9srabm8lyg091mAntufDqD7uX96Q/tFOB2tT1c2xlrayAA
SkDLQ1zb526a+khyMdKscH6PB2sAoylG35kUOWbelpjUR5uSkiYFkhUwWSoi7KLi
Y/xGO7xnJjUFHwh1hDWPzdVl6/6fpPRes2Fd83uhLNzeWjRTPBP79aDhxN33uE3I
lfdGLWR6DS/VWmDuC8Kp5n2HzhkmS45Kx3xJZhXXO5xtqEKgR5ZNAP24vbfnszXO
XQbWXR8Dc0VnDll0OexthQpmZ+Pf8t4br/H/AMMYwehm+JrhGRn6h9NRhVMKy6oT
wjPhJjNtsIiAF4rGKaSR2VQD5uJNTJEXuJkImp13oRIqaC9RHsgPLBRwCSm38SHT
OCOzqNqA9pZ8w4i7Sod+10l6dorym4QmttIGXXQ5bmN8RyMUG06WrAzDY8BqBus6
6zN+ZvMa6Bb7J2kCnvYT4LxGJhAp+XIMMn+HJw3QeRDSpm9w70s7yTFLbOxBeaPi
iO4b0IocdkNfSmVlIl3Vxk06epi+GM4a7qcR+6kJsFpxS3VgjaXqD8jomnHv+1gs
G96lRqnwyhiwBHB7tUSCQ+8FwIs9cMvFpFTd623pqxzh4u41+17QUNdlQEZOHhTi
odhwizXr5gIda6bkqlBUcrh8Hs2p1vUUvJrab2bAeYxYzykqvPc5hzTq6PPTmjmE
O7zEMY0wBOaOUIIyWSB1w3kpxSgEgbqbQBxwRdXihsrr8Xl/ysNzZzh/WoZyFxlE
HMTnZViRbauxynnpJF5C8zzA2W0bSGqWyszjkNx+82M8//KshjQURc2TcI23zH3h
ivW5ZyE+4yz8ZxYCD1wEVP3iN34vgakFQz1IrO/SMsdsoCBqqVCEGNwIeRCXYa3g
e3Npn2pl5I5uUb5WnqZe/qMgfGaO27REZdY7K/56I7r2bDi8RP99MC4lROf4/k46
uSlFpdAb09BrAv7cmIm3qTJiyb7ORZYYv/SzCJbCaQhQZ22onRkdSCt7QOK6jI91
kaHxcwfeC12sXTPfz1csuaVqfQpZj8cMX6LPNRDXl2d2Junzr5m+ftJzT+iwEaMQ
/vdITLxsENrPggUm9nt/nDATiJPqoE7zwYycefWQFl11bgs/RM1M9snOf4ZTyKOG
FJxP4W6OQxbw03WCOnaoqN3hYt7uMtNGTFKmHfKJ6k2XEUt9KVzRt2i3NnVwDq36
HW9VvfM+xJY52XSug4Qal15CI5P0TbdwM9pvm19nWhhNO78TsVgGlex7jOw9QqtK
scGmGyafjoK9zDPxCaH/gSxHVjnWJCTKE4Pwk87IuPA5do0PLAd/luX2+0RWI2v9
M9q9eOKziJde/2fcL9HJKUnZnQS3AHnCKoZroPcbIgG7xVPetP+Fl1GuKS002c7r
Z2JaEWKO1ljvYC760VVbzwHrdVtUtr05zt9+FfDnb4xAamFKnwxS4M6AV+b36ewl
qRHKNF4RGw4AYN9jdvTLqxoIXRxamFoiGkocjsCZYPtBwViO4mnMwOF8DZ15zn43
6w9loFopzjm5TzUo9YteQ8qWI3FXRqyiFCSZ9Cya3eWTrhYALFg6aq+jAJp+TE/y
QfLq/ePMX3MQhJaD8Ng1ZD1nKPd0gaIMXLoyVlRpbVxZU2ilQgZz/eI+E4KH7/bp
xL15JgRA+mHRHlavVxsL7bd6jWoVyOM54Bt3JyMFqYtJh3on1WRxngvryTlGqJZj
sAh1a3sw+ue8rycONZ5SzAk7MXA09EEgB12o2ipvKR8bFM35DDn5Y9oE1R504KqV
D68iof9auJ/ouhB07DnG5d4UwBwSX3CdkATTyHMXnD8SKrNwxqDYrKHN+yNwTXiO
ZHYOGP7L1woL6O4wpE+fgv92dxLSqDCO+1qcjpRusXqEg6X7BuZwn8na7lRLCkC3
9ZGY8d3NWHlWLpCzbaelA6hMUBgTj2ZIcSr7gE2ZIh+55Yn46ZSHJBu57AnGW8Ds
LyLd42fOkY+z81ptrIz251PYSa79IgV5xo6yBQvD8DgoQJQJJZDADJ5PT6s7xOtH
Ea88OfUjW9Opvzwau4xFQhC0N27WewWcs2FmAI/zSCQQ2r++TAyerY2hYwx9/uUL
6LINSXC/WZfW9IAC9QgKc0TarQBbjRK+NH295OerRT11rWPcXJOWRURHWT76Epl7
Z8Xow/oyvr5eF9VhjmOh9+0y1QBOJQRcBXVVgzziL+sUXeFthCFy51FGDk3Gj/mM
6KFlkcxnQ6+0707yZEJVjpqIMqSLsaUZZSGti5wj7LPja0lSwxZiBNYX7vm7ZF81
rA5JgPqIJlWbWZ7pgi+BmiWQ+dc6OLiqWsXKwO8IUlIKounMTtZ2DktkYCZzJgDB
E1ETayxrsQ3108dxvKyr1oKDzIzg5xgIsetv2Gh1H2lw7UCeM6SF7SeoMdNvik3G
EsCe+G9bEFv8F6Z769fuZJZeUI/SZcWYc6DHXq85oY1pi9BZwFT9eK98zbZUTQsu
10B+fy6hI6kDheGN1sZyZjNMi++KG6ASWuHEPm+gq2YT0iQSPZnOTJHukNfP3oIb
Ns5HIllsYXs+9j3DMALbauuqhAw0we0zUg6s7oZVx0ohq2FGS+/bLJqGQTOM4kdk
NNaR7Rq7E6eHaZKXOIFzyCAEAgEfFRm8Ez6GhCAvi/fG0XARxgsbCPr0cU0cweZD
8qgqE8qgU1v5xPFPnbz/EJvl+GizCBue+VxooARvoW1xFnjZGsDJYrkiKcbKg5NQ
JFxmKdKJA3TzNhv4kAHHCyEaRXoPIMaFZJnyou9sQhOIEKSRcGuE33YLQSAz/WXS
EnJa1lzCwWQseJX4L8SnX1r2qrPrSAbsR5IHYnbTv7WZ1XOacmYuYExOz9Z/b28d
w9Rpa1lso7YneITv1hr1zhcBfdENUH+Bg0s4fgHdVvZ7fU1zZCyhw7FZp8V4DVct
8uhYxIe/f8YYRvic1IDCcLtY8M8wUqTHFMndV0wdenP5jaNhhWzmfms1tv+98RY4
vlaqrDHC7anvmFx5qgpZ+kKmzQlyI53LS4JiTotDYxZd3iVlPIKMlXziupyoVoOX
2/4e/DKiyneOFu04PWKNHmiHm8KO1q5MhbUjMGjiBUbLKxOUdkZ93vcbNw9LwnPJ
pKicfIkBwINFgyigN1SDVScRDZadugW5WQ8ODs7g4+73x6m6XEAIypJdh+7dc4wy
9+fD45WuSmx6X+w4FqSOVddJ21hkBcgGfSEDgW9QGH+lDrtnA2KZv7dDyPGLJ3c8
Xa2hZlzztbzwfbJK85wWUYsVysMpIy4UYqHVufqm+izPZIk5k4ZVPw7/vycQJw+S
VVZbUboIrJK9ebDh7P4YAonXxIYDQiwmw1bPer0CT08zOXuHK4YXZ85diShO8YsD
TNgcMaSuBYJfZPVjqACsdI1lrh0Kuz/R3jBFdvs0D8m7Gnupce9dFKnWpRXG5i4z
5z0r+h1V8UqxRMIsI6mPIC/DWNjj+gNCWCTNQiyUsraNFVEzwiIjXXSOLKipovFg
AaGFC73QcOUkgduhtkpaFTEQllsPqm/LVECORU99r1qtofg86Aq4b4OehhObc9Ci
Nn7fIvE/0Oeg98GfDIN/KtZxkXrtli4pgNAMa5B1vjw5bY0Rlegk0ZBYTbztnCi3
+DwZzCYje4aYChtwxZ7FOTwMMpIeHZM+Csmr8hCs4RQyDSracTrm94bgFS/W+IV9
mgbmWXxlyvykMP4aPHBXyyBtqEYXOy8huf/18znkj1h4pUvq75Vdo34JZPjYe+zp
CpcmcFx6SPZ43o1Pwc8+Ios6kRcu9hhFyWp2nLluaoY/PxgP2l+YPidTV8/E/t5T
YGgyiieJtK+04GD19inozAlHuKSF5AMwkMi3rcrwHaoXHk8nwBtV6LLaqKMTa6dl
GPcJhIDyrlBbqMZfZMaq4sx+NBkng0pAjad4GNIioEIIOPDEPUM3+oIdVDpY3cE+
YC37K6ArMJtTBoscHeILIsfW2DlYGkeAgaiEQyRsusek3uhAsaqlw1Tqa4mEl2RB
KDkv1pKnj+DMw/UbBmaWCddmhq3EYHPyyD5HRB4Bijnsqm231KKm8r5xtlwdB+dB
5e/NKPKMobA1fwAcopunsHRYuATzmvE80r7Na2VuawFnAbBpOcgm775ZakTbgR1k
KR4Fn4lDuy8YMHztukHUKsjIU78nyLHky6RMtJWVeoZoVGmLxl9dgOgZS0/9iw0b
8OwjU2+Ud0zynXgD+hNlUHSZta86VYarNsrk4jHQqXPVDEf5Fx4ddNfJ1Q5Vnmwx
G26GWZC3BfLhuI7Mpl5DVV/AAr3g9jVVKnN2WBYEjTVbhZ45d59T4PSq4R2jYNw3
Co7tWQhMdHc+oLVOkJrftqxGkpMZdJQfFX5R4OJ09blwYCpkZ2mL2E+BTfw/kVlm
9HJPgD4y9syDUWihjJnLFCaBMqoiEgBwWC5ns5XyM89d9lSZEl60YDdbd3BfT2ZQ
N9y1h0qvu6fa+i+qDxM1IbHOsceZoA7Tj+3D4fJkDmoMNB5MMwnWfjJZn7Dtbo4l
q5peOFcy8UQL9kCGSd9rx0Pm2BO7M4PZWhqmXbTF7SSC96etYJ8PE+/Qmjfs9jz9
hHFUH0a4NEx7Ra0X3ereivAs6U95BxIbjiKsbQb7LNA53DAJ8l5QEW2a1qgJNpE6
XsQ4QsLJClxIaDTttw1+jKaLNBrdsgWFFJkOCfq+YIDVlAlQaTg+yA/5aU034iCE
i+bZVkF/WdkXD7wXcDLu79U1gieoLnN9FEzHqgxZIIUNSA766ZM5DhOQ6adceGlp
d+rW9uMAFaRX5QclfQet7jwqU+Z+IYwlm2v6/Sj3cky0C2mmmYohLblhw88btr2p
P3Chj+t1KzrlygxXXrlpqvFWX1monAnFHqfNVmCPRmR/0wEgD5lxTKitkIFkYOdK
UV5Yr8/yzgrGA5Q70zI3ARntstiCku6yP7hnXz/BO7a2E5DyLI/8jmDeE+b3AbPE
NtTdpVIZahiS/r9+aCF1DLGcvMz0zGqIjI6c/DcCoQkwxFw0d+IwCbP7UnIYMSvf
G+AuEZaxSD6i7/TNa1C1xAjjXTYllRnvnk9l4tn5kYuWPqZPRfNRDoDjxuWhnRz9
AzCS8oTTLEsK7fSe3lK7vq1zwm1MV03Pjdj749jDKd+lZ6TNiHirIFEifaFia83Q
cJ7so2QW+dj4asos1E/gy3YfFs8KFCuQ46p2MB0LxFud6FFTTLgSkFpw5cyXUnyq
vfSGt+6zKMwGGEVwO9Q7Zk4hs/3EzRE4lbwRdocK0Prat38MVXGMoFlsM34zSWL5
/CHMBam1k+C5jE+IEIVUz8ePazp10mcPqqgoR9O5UK0R3dPdFW1mzUUvwKX820qk
9RtL6dR+PohuywmRba/9CW5dUP2yVoH5ElhP2SIErq5KAIWhNr47AKirWwWww+dl
BYoGjNtNNlzs1HXoBij2QP7Us6EsholFrzUOSbBvFJwVPo9XcYfQLuBA5XLxKluh
vkp6aDE4SC9Km5CrrpGl6GtfRdtMutTHyMVByUD68AIg0vFBKclnBJa3r9aETrRx
OzNuVp3ecnRrCMjm9o2MFMtfyr98+mqGIrQugDf+z3eAG7kD3+05YonBLsytzjti
+5tmlKEP/G1ybJi6gACN49GnAhsKL+5yuOefoOIw9bqQI/NMtbtwdJN5WdgDeY6I
QcMhKIFZsrDvrHQ5VqWMr4DrbKsg9gtzFsf1m+jOY/IOtV+3/GY1viPNkOV0KmC/
tMAe9v/Ni9ynAo24sxAYhP+6D+1KlLnkCnmTNFg4qnh1rGyKJJDWpfWXvs42mBtJ
OYNWfkep3pQ1A3WnKxy/MHSU6b+kHeCGKnPkXeeJQtBfoNasqokPuUzMyHGllhaC
QxAJ0iiGWchQC0qg6bIiNKttCFZfc1suEt0c0tQV5LhSrdCvUzH7H9evNE/PGZhs
/jgE+bwiO6zzGvCqXEz/ttqM43wKfpnGQQbFLM/fb6vAdgWiPWmQi7El9L+L6RX2
5rbptJrhWVlleu50YR8D7UQqIDDwokbVlnWn/S2+xvW2e5Gcy9KLolBPChHOZBcV
HvUQOKRTvNI/JRlAoHnzgbymXO5qacMh++fzVATEximRV/Lxiv9S5rnpOHk2Sroj
QYzVc8oB+7mGYfGISfJQDPk9WtbQiIUvpcyN9WgtHm5y0/vVDDZnPcYnWXk4V0G5
5Kzz63UNF2iLYGec2SfvY/1bmBf11FmOaNquuA9pvpUtfIN+c0ALmuh2ypSc3fpC
ifBDPzySANWc7TkYwFwZ6Pgvpg44jecfhn66Cwdvo0gjnEu5VUc4a/vtHtZvRTub
XGUXfjH6gT4lrVAgdpW8v14z8qgjD+NIO7+zQkVF3RF0OB/RRhdLWcm8Y6mztRma
7ycrkwIOsTvMLlq+LsveuD/M7j0oM2G69U0kowwazX9IxPsNpZMUv0ktPkxKF+pM
yWMuHHOXT0PGfbx5IU/wUHF2apguAondbdMrMVc2YTLFBeatgvP812BtvRTgTc/j
TNPcWnShncW+cQk4ZERxqOO2nkBaA1q/gEpykbt+CvAZv8PuCZBOC2XQDekV/YCS
x/F6JIG9DTDqDNZrXZkM6+S7RqMrzVGCFQ4kdi4LDeCJDnayLpr9YbJ8qDkhYlHZ
UfRrIhC7nGWZsYBURf7dxWypL04tTTMbyz7C86sukTL1t3TtIGdyJr/5AbV9z8Jo
+Zo7COlMidA/AXPteweWcBssH6jbW5Xb1TZszg8bYzI6YJNLD/3l3U13dJv5oMU8
N3oJ51b8z1ILZVBMZjVIWe3SJWXFDp5c+dOxWo48mcf4z/r783ZKNipRqOwFFymz
BzZLL87Cse4KHAwqAl2iOb01NvDuI+3kVXMJMTO2Uc5JJM2O6JxuWKAbWfAG8NcC
RcsaSgCEuB/PgDW+BmjsaMTQRe62dMhvauzrgSvGzpq19PL6swPbcNPL7Sfmkzno
VgI4UP50HGLuGb4u386/7pH7sZG2M67+yF3ifD1XEwUhYm27I6/Uv/tX7EGUYine
KPkUctPtH3WpL2xZkHtDlkzwb6f5pdt1N8Qp9XaWbTPX/nqQZVKyIf2BAYm4u0IK
QwPSlYibdlhk+RXCJa0R0bzw3SkVmBYs4tBg3zpub9QyVU0xXFOLRk2iTyJdHlj5
hn/eHFnfvmrtseD3I0aoAQWu7qImP7n1PNwoZgFCWWsYVnxpGmyliKNKs0ahl9Jv
LIgzUgweLOxJUTi3OsCN3Qtho7tQDIIc+pq19y9V1cq+8XoFn59d62cRue7059R/
BZXwFtlEzGCrKJJPDAs6fxiJF6xGnnjfEKJBaO0Lg/GXAAHcrllavWBHQWrdsxu/
KHjfr91cB/Bc9vzrdE2iFP9WGpar8DCsMLI8MAYIbmlSn69KK+VGMk2BZBdW2Zh9
pw/B+H4oDDTi5qANoEHjnhUZQa308xNVeQpdv2K2ym1okWPX2PLJmXUBkV4eO+C7
32/YU+4wQAXTyZAzHk5cSVUD8y11lsLIYDv6fguVENc1WpKvqyL3kSLQlQW10CGd
Q5W9e9laiC+qjvILk9imyf1ToF2Fsu6EhjSojISdyh+8eVJCuFZXENuSeQekXsnk
7hnLqhiRBU4ngdxdJtJNhmYYpdRfNFRVDlyc3x3LmTvgKrKg4St3ujGo5HV9RCKa
eeYQY0pu8XQhlOTInc6gLbpzShmJgYG2XoDHZnWc5ynnU1BoYJ2M2hvy5vt/AqfK
W/dDCR3ZnDAH6wKJpi7LgEPYgC9rfy4plVDj20EpYyH7RsaZXPISkNxlp2vDcMjd
8sB1t1DUK1y0AHuTpH1c+2zE12rqRwrs+9o4KMSYIpFRn9YNhJis8vl1+W8Mul0V
BZ+aph/XtLWX3rKQm8hyOlZGNa0kyu68KIrSfLsrstUPMN4jWg1bwT4aW51SANtk
QP2BEkWZt9NdV9+DAK5fYDKTij45NYdG00WLpXScJAaxC1pn0WD9gwTtQ+sYZvzi
qOzCO57jewjkvKU/V80bIJROF2Q7Jz5IofVlvaZvKYJ5U/89oMrlcg72MW5UYUvb
6aeUWiHyO3F8QalA6UTkdiCv0SlT9/4l6qUb9P8pR/PURjVxVLio5Jg1QT4Yicgw
VZoDzSad3MfeN+AXeCM6p12bWHk9NrbI+/mIqDuttEo2UyL/Vx9iIatR7wmiNcnO
//HPpMSZ7KwhytD0tiqvY+oLnShOBKqGWhSOgxDg//RYnzHxRs1CON8mFurN0rd1
X6gj//vSTq0cwrMOgl/cwWBScwAClEzJcaaWLDwSPtvsYMyCyEQmuv2zUUucNYN4
lv9jqGUExQtbfqNoYb03oNe+gO1tZql5Lg+57Ubdb6aLAh4d+gqW/xvMnYvRuD8U
XLdcBKShVfimzvPk+R6ohumtZxXd0g/1QIIQ/bJvJsArR7FtOfagGmyv2SMmwWRz
ws9Da6vNVxHRsBLB5Rz8MR6i38ND0OtrvJhHcy2dfSe9RxFhxsNBw2fCURF+NVdW
tNQWlcK0zcb38kGedumqiA/NUhN5hm1GPQy0aHQVVBwdcLUKCJy/861lga71gah1
O85i+FlrM6QfZ/GZN18p7njfFfeAOf3HCKEtNFxtTlWKHF3EG1ZgpKsoqRAFxEK9
bA5aJsAmFIqSN35hvwcHMgTG7i4lmCQOJWV8CgkvF3T63+ZFvp9z9/HZma1bd89X
3i4FfICa7hycXGYfmybv45VNEvrdeeLKhHvtXRamG8knDMXvUIwxAn8xiN4WdmC2
9NaKdczhj1HD3TGV13+DB0qnoSCZKR98mYNtKNvTWzKuJgXpBL2LQ1IRN6/7rnkq
zuJD29feFT4POd7TUixs4LHLG6GhoZm+U5zCxFGTB15B1EXYptuMPxStkIwHPAcx
JSMzbJY63JsqSnuwoNr5PYBbN0FueVX8+GfSWhE1cQsqc1uh5C+DqUhq5qJmDYd2
1gIDdGEyEcWJjlomvVpgDUv9ZQvIIYQWE7mIE5HIGPY5Me/9bj7/0SY/D/rHD32f
0jsHA0hsmCBtnLmy5Btu0qzDjjLRsF7AbEjLYWYizHHckzlHBTFJGTtw26geHTZC
psq4lZgAYJXukBUw2l3QdZbD8bOskN0Mflv+8nMEH2uBJYoNuMY+nuh8qrlukzNI
UtudWL9HBWRYzUyJt3c4WY5IaEyn1Z7rR6Jinm0ikPcvVQysaLN5UQP6sAqv5p36
+LfnSqPsbkSVZqNTu1I60PhJXGt8FKnhTNQZeuUdO8e1+41EoTMqa68AGSjQjPlc
SNmv+ffuzBCxENPySwdD0J9K1IAdp196CEzQa2aaTUxu0kpTauOnJwVNyif87JiQ
+qhTrJZJn8iDBOO1J5wCQFH4gPldqlOIVE5AsfRf+tQCy7fYpAOaji84GuyS2+hs
DMtyjrpOk840t4BEu+Arhg3sL8/GKfiWRLdqvJAlc8WhxQjIEPDVK+dFk9HTa7uN
WYckcurlpK3kIp0I2kJc2NZpj8GJLk6IjqmCQiyxb7SEOh9KB4Xg5QFQE6LJTNbs
49yLgpJuZaC5Anh/UOzFuzXt31CWkRBFxruRon+9x9CroXz0wg3LpZ03RgclJCfk
caTMqDSxsa4cfM5rhLR8bDjdHjQtvgmuSNNHuowIdRqp8uIQrEcz4+/KxtfFSc+b
+t73EXlHQLJScHU1d/2FFcYXCHPTd7+X+Hlukj3E47qpomcBLom0Zy8wL9nFfCbR
rlGfyWeiEZQ/7MMlfMtUMYB8My/jhDxZb1mQV8yBzcJ631xAaBd9ZVP8HwrC0KR9
Wp2lbWddgVqCM4tebw61u8ZRBOjWZpvhEMgxAD4J0+iDDOVcEfRUNI7A9D9z1IkT
k36fMXoktwaolRhhl1AoPhMBY/CXoTmXS3Cly2ENpm0+PjmlfGyQPN9afWcQLTBT
lPUrV6s1YiS3eOE4c6xnT8XNi3pYQi2MP0k6R6W8BUKqHNrEFWIrEJb0dlALW1I8
8FLkGo8gzN9EoAOXrFItXDFFgtIqDqxf2KLadz8L/a88NsbtQztvp0VASDKwrpnV
SIHEOGvITHljUzPS6qx78QGE+RohjeaIeKbLaNXCgBFadRWTqjMJqwaNf7+ULStP
N37JyNxS8X1JaPS4DoON9eGwtGqVgn30/0N5Am+vMJPdFBUVdmbd2azrvcVgQW8U
Vt1AvA7nCoQgOl4odMRYj+Z844yY0RHuD8UEWSoofZ4t1RcxmaZHGlh834GLRK5o
SRHh1U0i3uDX//NEVOQ48/WCGEodoisXyUA3mQRGuTmDTCB8PytGXDLptlKFd5U7
+eLEeYaN92fciQYcjLWUBMHhWBkw4EYMjUle5qpItJsHJ/3JoeN97OHCnTXBzgYx
vNkPcT/Epek9lKafg/kDh1Cs9wTsacfMn7iE6PJ8El9bAB9fGpwpLdE5Bi2F39Vz
WfnK8QEnH5k/4mhTEbLudb4DyzN2774tYt5XCYgn+RJLm2nPL3ZH15sOih3Wdx7D
QVLTMS4qfYW5fLRGUz5mcE28lVhX6sHGX3ocoT0rKhLq6n2Ad+113Z03jQIxNHjW
GA7cQbI8TwgZFFd1W8r/PDGpC9AVfxwyXtk+6B1qfO88oxjHL/bKH4mHb8izV68V
W2HhAIfuk21ZE2csIQl8Us+NcjSab0ErtfgXMUPtBu69+4/BKxJZrptT4DnBJ6S9
d40hK7dbDyzfqwQpp5dEx0MwmN+KyzlQPE09EszEWscdL73AuCijDy7x4SAVTymb
j1+DBWlDacX6sSjsvzii0AT4BDIZbEHg+IKV4f9zUd9MicHrO5pKrZwA0w8mVEcN
7mYjAHASBAhZ4JIY6HQbelN68F2zM7yw0ntmpRxn+uXvvtKrEM3oL+d0K2ECiN+4
+NmSAMOkFYjK5wdlKZYpM4aRKqkPGyLHbB39NPwxJIczua7rq61tJebF7jNzK4sW
rhwYyZAvxNkJDLqUzDnOKFi4mY3VjpoPVeDj2zKeelpZ4OtbLYroSKB8PH3jvdxo
Z7uyjTygPTftLyBiEgcq8ORkrKUUNkKqSeFeqsiSqQUx3baT9Y9/BwV3AF+VmG/m
b0ECRMl/v+L4t29Aiza7RV1l1W48h1Lf07WTjzVhfpB4y0yjzWMzQ6/iEiuhCq8R
M5sjHAqbo24IIHcpGF4ckoUyXMyG2jPMRNpO9Wu0UJ1f5MwqrON+4ShQq68X8eEc
3ZVe8EIkz0atjiSs2ALIauKNQB+nWjwJHgVxA+oZb59cH2F36+DKpWDr0Qu1Ftob
/0gmaId9f+UbpriPeJmrPZSRmfSJRdW3Iz/6uQ1EZRTkVmp0DGOZ334k+/VkKBys
YCISJcrrFvNWiEKhkYv+96Ut5i9TWeHJK9JzTAXNJG31BSy49pUGwjw6QddVD9yn
o9W90UNDHC9RjP0jUIiTJPsTL1kPvPpJ4uYK+EzhtMK15R6n21oAvF8E8Jt1gb1M
h1CC+wmgpu1IrRtS59dEPhdLZpU/eE33l8eAgOY8C0ogogRQY6Za4351yJ194ONi
Gi+9wsrHkrSh7zjdBn8kjmyBEyJAElHgm9ugGFDEpzL7YrMz0Z472zzMEnO72S1G
160/XhMyO0/ihFpeMkQL9tjcbgGMsQnlchak8/l48uUj+qhf4gnSXtSWqDqIDK03
Wg8EBw1Vsd9S5U+6731W7+dpuZuGR/yWS7UUaZx1KMzxeJFO4juJcv5kKh8E84q7
sBpYSzKhC7PzCNAypwUJ/I/gwKwVINOSWGf8Awjc0FyMH0ALrUe3IGdVMiPIx2nr
BbZK7QtFj1lXF+BpQhpRirqiZPvA0i7xS8Zdd4Lmw2bbCc7rm3XwrNNLgBV89HsN
MLEIy2kwNy29on0kjjDEia6qePk6crpjqQ+XD1HozoWskO7Z1jkiBsanXSJ6WkvC
fTunq3edHNOo6D31GjS6amg0Z2Arygy9nYCoRbXxysJryGMFiNRZkZ9aJbaoTf3k
gEfZDME6096LzspzT+Aa2ies5exp6/AJRLzKp8BmrlTer3MK6TBDTOQep3eZAlMs
Llr1fPTc8cIt7gu9ucHcJiohe9ypI+GYcfCa0tUjN85bvewMN3L8A3jDP28bnVJO
iN49zH2N2bEr8RI0j7rnhtqqiGD/ihlSlkRQsZfhddXAjWzsnvviobHsBRbcINRu
AZ3qZh0ygc1Pb/2ceYwPe9fMF83teO4vMHhVUpljOOqr24cUCqgU+a/+q6j4gt56
6bcWkrzamW02AGZP5qYI33Gc6jzlSgW8jn3zRZki12MwhxIKDBuG+tNhQLxE/9pg
1LnNC7K9nNW/hYnF32Mc8Mn00Ga4wx89GEf2jQYzkq6Q+OZAx8AAJEORs0CRR5rv
GTXxNOoP28r0up8SFovu2HKrwWVmRKUcdL4dFTrC8C0VwbWhGrnog11T/WnLICah
/H0y9qosjhoLvUheSINpvxMJ6VxZioN28HYgqNmh8XwLSD7iKdPqvoVHvYj7qrAw
3+5CKfyqfOxtvTLygEKQ7LXi1wSMdNK/4fbaiQs9eCca4QC92skg32PzbGYoQDLe
jWVpH1aQLviogzAADvg5DkADBzmUVcoR0ZxIVR70oeZlVF5SE037gz0cu11q5vYS
nGEpOZIPpNTG1GSWHvMCPDKkXc5ikbC/V9siqWdPkrB7SZcSt1YumfAiXDlJTNlX
yETtcxP6dZxQLUF547KEXktwmyhDtHpLD5/FE8hx5Jeo8dGUEZ+j+TTYk0Y6WkFT
47ju/ozfhsbnWZ/P2iBJ2hS15FNVp/daSbCXPyK1Oiy7LGAHBIx70Vj8uFOfaSJF
jrfScOzzeLuMqIRzOCNtTTKTMQxAqGup9jntNTTHxgXZQnYyk+JoZ8J6o2HofoPL
NsHSNZ6se1wOtnO/w9RivPApkCJkwTxdISQuMYNoeRxmZb2tevL5m7mlG4ro47v1
21lBmyB08ZEl4uW0jDbFpuPkDg65PaoXLNvRAXPvG4ktZlEsLTPEosLiupdVSYOg
rlzpvCQJvYdVeYfuCZsqTjJsu6ytmIiJ2s14d1RB14jG0QCpBWic2OiOZH9c8eWW
vZRi4DkD6Wg9FLmYBfqehqMSVRLKxkycktQjLAGx/ACTyoVozwWryNUoJDRsEX0I
bmWx0R1w1wZ44/O+ed8onK9A1Sl6PxVujNxAWsC7fRAngWJPVK0JptNyjg4e7GnP
c1nLBu6ioiA2GrnYE10tuAu1qiL2Bqxp5fitLrn7daEYQQOvEOJ8JKXbf0Z1hhsI
n/+6OxkYYa7pJThBPui8rVo21Tc2IFeCX8004dx06WZ6KDR/fgHTrhkz7levPOMu
6RJmdFmyTgf3b4+BLYLaw/F1EdgaHRhWMqpU43G9i/FxDulP96bTYlTCXGGmeotn
PTO/OflufObAHG56S54tqXMWnYnL5LBKRt93ItuXlC1I3lbxZYTK6lO6E3Z2mT8P
kCbCV67CalkCBfgBPR/8CWhCNARfSGcBe2gkYIPR0SEM4VHODPaKwbbHsuosIFRs
oCoqVuPEjPrBEj5zcH70wWSJOfRCrZlaBatxAuLJqSgWHBzDQ/Oxy433v4+OGWHF
aJsparGFxSQSSoJ1U+xEk2tUunbL7153iBFDGMP48PKmaNpTEntpouqE612rcDFO
OR46RsOlVOZ3yNUJTXEsuNbgP1410iAjqeS7C45HZdcMpZ3pwTQfLpie5o8GKXIF
AP3FE1w8+1ExUzCfuI5Ku25JGXR7mgV9JFiDRwTGuuMyQ6Xa4IG3elNoGNDiYoTi
EGYxWqXqFfxs65jqYZ4YjOfWqdkkn8cUDOMYzO5N8tubAYWWGxZ4leAFn+Spzj8a
6W0/Dt+xWebRXrc9SwKbFwTNxdj0fjDwPwSg7h8VLLcoZdgw2/y41ZNxqOHhx5cS
vJTw0jBwMGQ9p4dE5sgnsa1gV4FkpQgAF1Aj17eIPDBAfZaZUTKpm8znHlHN7bc9
/RNAWl72+c+W2d72eVm8tQszOGDH7Q/iT0KEFTZsk8CjyTSEx7dHmBkC0NK99tUM
SeDw9eDNoB9Xf1Ols3k6Fj3bizlkR8mpbypGRHoNHd2Kw8onZRB7VUMJ/8QxpXiA
WIDBFCtV6y8CYNi6UZU2Np5YN4GgXbP5BGjYKQP9eO9IY9AzBP0saX44ZpAp9WMY
axGnRtks3c8RF1Lz+1+3dyjV7J09j+F7zoeFo7U3BB9iBSfwClY2YbiKjC0UEtFQ
Z+hrfz6QZyPXCNpu6CxtyCWTAZK0eO/rPdJTvF41S05EQDotzQoThwdoKEA47RA8
+ATLmg3tWHdn1R1PKKBGTafJUk9PKIi7PhiBdD37SWbLqvEv8qFgmA+YvGivAxT+
0JnS8onnP5RK/lPdS4DljJOA1VkuABXkD+sBWtvNh42hsRdi134RJbuLec4D6I/D
F78pZx9bRhx6xe5tBVmMObqKJ58V/00cRsdCdxaRd+B/oTmJ4UC4wkdUKAuNLPBn
b5Q6JymYZDcV/e7p/l5r+7jPzv4603qTYV34Mfp1WVDxYSOLqT8bIXp442uN6dFd
BrtAPJtfaPoxXRNBJ5F9jPbMiuVpMbK3hGlTMJDgoCUi3nS9lkFP4dxPupjQg/Pg
ZNJKovETqEWSI0hbNrjLT2hHEUdYZnCoK749smg+i3wfUFMWikUcJuNAhm4G7Eon
/YPfLIU7nRbjbEZhm7Bq8DeylOPZYSeXQjqWR5zmfIbc2hFm/DRCCZ0f0wHvJh/A
AfEZDnmlwJFgkS854lK4F2M6CLNeICgfgV6Su01cjwPJGqIef7mS4//P35bQ+Tck
+R4AW/xFraGBNQfPdDDALCjg/dSM4we03EpCKvgTg3rpiv2qnYWPVSK/AFGIvnlj
YXivCxwk9chx6kw+kXHFSX3vb6kKTYCchvNQvZcNlk628lVwWpaUcV1tXiKIuwRl
5irf6hYsd+nd9nMg6Y6c29f6iuKjL0TmG9A+w9YQi0T97E4zYUKen32LFE1dPTKu
wPOMeDmHbxqD2qhPzNse0r/uJxW+B3umvBjzYoIzOcwkqXNHOyB8DOexHzNiRTGV
YX1eqnAG7HOT2M7cJkdpcOcOA/iYitUl+R9SLZLKCq0NLW7a70lNGTbnm5ZK+6Mr
l0mHTnXdKp8y88en9Rr3GXPm/vKac0ZLIA35Ke0SQoUZW0jE2ZQygpdjdsh+Sjed
+8Ew3yDhF6y4M4vKhfSpt+1uXiTUvH+K78RQo2jB8K1Yz6ky1Mwx4ft+nTkSm4d+
+HPVfhrVPux3HF1FAh7VdywSBLPPt8WhJX0RMCeEbwHzo4vYlIZCklguOaevA6AW
zhH9ArpnIN7nzjM4zzUQlg83I3xVIjJVvuoTJYpNidnfB+AYinhqPNxBSWEROXCp
5vlHrJ2txLdaHr1ddfFi4CvNTCeGz5SaV4x8pLhFH2SYr0SAu0xwdODJZZlv58/f
xtq4uRDWnzvfVphscoIf8YHBAy3a6O36XbfzlStrTRw2407g0ldqighSUwLonIV6
DY8w2bC9N0GYG01xE4RsuTXhbN4iXjoAU6EVyRmPcAQrq87cte6uffs9pcOheG0k
Xdf4fbv7pA5GXOJDcbVCzAaY3ei7R5KHIEJH5FGHOUY5JPwdVJqhYpJYa7zeHf64
E8PdRrzjvGy/3S31i01sdStdUiaPSiTJBQ5eZS7HA+OZ56cW/VT3irDlua8b/T/L
R7tQzDG79Y37rNKA8AGZaI6xzjcgRq90Ki4CP2Riiceg5gSDyA07GdfULslCqQul
F1aWNSWfJHKvq75V6WBDl880AEJcEjPPbLv4oQPl4pOSqEosdFT+rLG/Ux2HVhcv
f6inYk/9Z/uRxv/ITR578vye64h8lnj87PmE+q/7laa9HKRRWrTRxqMxN2wBeAGK
zQMMqSSwFVZbegyjTucuc/n9r0DllB53fL21AisG57I82JYlvDKJ4zvb+eu+T6M8
UdRu27yyAhd3niDazd00T04r8GggAPiybQRrtEd5OF0BpZIuVsRD02u166HTM8NE
RGx5DJoix1iE3W2xCpgSfEpHxCeOZCmQutI2sV6WZNz3t+m4KvLQHnZc+G8SUO6c
AAlU/gtTrfCVWo2mmWcQZDVLBCGHUM2gibzBHYOMaIba8jxaDZ6OSuqvgbhSUJ8x
AQHXILDHAq+/WbugzQbPSnMFNTYHtwwN0WxhUfRyGvv8YUc7Cq+C+VCAqihrh1vW
4C6mnGI1WS0BSX0dRSJk83Unam3n5FQ6qlHFBOGm/d1+IroYCd69dpJU4fwXhxu1
swKhBz36R/kvixSOaYDRB6UaXJIg74rXQPc9PFHaBOSI905n4TZ+OWYxa5gjines
+IVKVQVdAaevUY3Mo9f4e3sg/fOedp0p6ExwUKBSJ2MBimLRpZx0yhg4TgSqdC8N
xydgKz18vf88OBxHSk90Vpc4BKQW38zSLOfFLVgStjUEtytvn/6xRVSgdIoYnV/5
TMtlgHViotIoAHg3J8j62rU0LCPBTMk514kX7OK/up9wNH1O8pcFr61sHbl0JGf4
vn3NWp4mZrGqsCQxMagq2DxWfCkq6kfEKJQK/ohNYUwtUnDgTIIStBTR5nhCsvTC
msaYz7SWMuIs5WtpES+OIpl0NvyyqdXsKJ9q283rKxGSvCMBZ1D1V1otXa/IecmF
kn1mJ2kaCyo22CQzhc14Mu1O5A991uG/RJmEmLZXsmkOUvlIZ/u91UOMndypOMcu
dgwKsDKRMl5Pjm0vv1AnOPnxhyMuK3a3zkHlUKa4ojfiEaUJ2J+7j08y3bwaLDXw
dlQSiFV3N86+souh/AKyx3e7YyOPROLJ1DqwT8+REron46YBQW7tjcjeS1ErQ4kE
ygchTLIZvS3V/7yXa15fBVQ3KGVtHFNDJhKVv6AGPEpClMoTvgbiX6Q2qX/mIMOM
G9hroNFSYwvYIsd6MnMVUadZoRBa+zz71tV1RuyYSHT4yg2e3uG9ssn+dAmab9XR
+mgM5pD8gQu5ce1M/S+1UBtcAjaCWGRuNpxbkZhnNkOH5jO877yTRJTpT0CZq3xt
GQkjfyRMh3BK3tABfHOw6sW7kUOl34lnqJ5jDGLK9GmJxWObwd96hu1BzubGK9/F
fgbC+745mKpL5oRW6+ThMsiOCmAuGYa9uMHy8InPKvNGIA3UAcVwkQTrw+hd44Wx
NycIjIMqb+1+WX81l6b/NrqJ2PiupIzCcmR2oCjy49Y7qyga1tRZ0Vpvk8kvo1lJ
SSdFqpTpBeQyMpuB/7Os2lMNPVb+LX1duUWNDg0Bu1WxSjU2wvzvmzeu/VWycoUm
cGPEykkjxQMPFf3Gi73O5GN1Sgaab4QlzwzrDNCUZzBemh+wAYxo2EyZz9dB07/O
l4Aadd3/GbMd+gzaZZva2YTDgwhPJj/6Phk0ffnwHs4VO1sdFrt0mPGFtzg+NxLJ
QiyUC6EOahLfczpXApC1bbwxj9aHvWzCR+VyRNx7Ku2vwCfdYREGx2T6O0E5En7d
9iRB4IduDfs0wj4aMtSs5M8z4vMa8ExI9MBtyoXTWJLWZtMPZVvSh89xDQiSA2rW
yZEPZFIJoBQ8AtzhAwznR+f9DeeZS+3VtIweGArU6ZuF1clPc91kXrdfLRwZPJP7
fvh1TtWGytlbAniHWT6YZkxpDzwLRU7RnrYLLt9aW1eoTeacjyY8j7c4xWZIEK5B
vrDrp/0SEcqBsxG3PygzdnCdmEyzQVGvyogLtqxitEYWmsVhbe7SdElvHU6mhL7i
9IP7jmPU8voeQYTsIhJUriErlLQDMfM5D2PhUcgSsk7UwYBQwzR0Zzu52NR02wJe
/Q1za3SO10Ovfg5P5IPTQt3Ak4IYWxvx/CZ0gSRA81PDKYRvPdJnr87gw1qzRW47
7RDqQpq3Y5iTfnfAtqG6Y2JBYt9lS5KizeIpaU6Q7+1l3GAROxWBr4lFWxPx6Iyv
NVirndCUhWWr4+x7eRcbIbK+GRFRPMke6pIfdPmU46UWkncYMrfa9291TFhVXBt+
sSbARA2j2xxsMzm+Dil3+AMEqd8ZPAZ2OatLh9uzZKNcwUq109rqfIkU8Gg8gHL2
gUwgmZlLYuSJGkOtFiYrEvfoOrf4RTLoHLPiXOpJbUSvcpKO/YngZ+F3uZFcMN75
kgBNnR4IJaBcp1jFaeuIPOHpKceG3blXClMcqjgqQ76hsNmOQd3yLSjOiSKRJz2p
s8JhOxAZJF6W+p8O0wugSnbkSgx7lnWg18XV7AzRU38phP2gjHxJs/6vtHKcyFRE
GowTddvCqyUf3/jGAKhBWOUgPRZiZbZ57aFIJdRes65ivHhJXdGHM9jDH6KfH4dz
i7f+8X9+UNOJ+00swej1nDPvaFaYfd7S/e6wl5r5h8ue92P0YdKAWEinq/6GXkY2
xSA9AyLPWb9pSZfyeJfDQX+15l6T8y7vdR3tEfSjlLKL06tMJpuxIU2+yqMZNOkk
l4gMbWiZXftykCqinGuE17mjRInepETHEQ9h3tcX95ZZbfpX4xhjKuPrguu59+CH
ekKIMMuyXsi1rjSwS+1+uvbZgLHS4RS7h7eDcWT/LCansoKer+i9AuPhtP37fWfv
SygqGAIqi9JV0IE/RuDpjw6E5gLu64P3OFUylGQYBx/mb+nea6/bCv/umExmH4Yx
si9xk+MqGjbXC+b0ZICzvxzBNBLJUkRlTvHJ6N8rWve83tTMmApvn46votDZqYQv
8W1hHvbB/3OHQd9ASufgiWM6+upu281ISRGHk8oM6BGiSqFq3FmrFwSiyF8mGH0C
C0ie0aLPa2DvaeaCrO0eCHwkJ4JwGFRMyyNPFhQddwm68YBF5sa48av+N6+EhTyr
5NEPpJCssaOxBbIvJjat/zVhnY2JztQ9ukJnBN06dwcx93zlyOKoNcYDQugne2Xe
GMA+vl2HVieqtSmsN19tPHtBG5oXxlHJQaeuIeyjdbRD/RargnJE4OKVIPLsTwX5
WC5PId+dyyEWhMdsPgBVCUfX4a21gvqdK1xAbyKc4kttv7RZaVnO2XHmr72drcSt
mPMGK3gA5p5EY3gz3SKLU7cGfrUbvShYs7g/QMNxoA8tUJfVuGnSbJNDHN0yYg8X
CWoes8md7NONFV3K35q+tKeuGnToMAi7PQ57UY7dLYNnWFJmjzJ8XrR65lkOKWrN
hmn38faeYsuBP5TPpgWHwX9Xt9bKt0z6xkmsJXWZ3STWXcsn6FjTd6sFZj6/fe/d
0kFYFwZLHd3Nj2JnbWgbvz48yw38m3D1GZ63UPFwe7UAcyobYruM/JA2WwvlUl+J
V0hqrueyuqWbVRfQx89u+vntldavCxYw9iYPVoMKJ/hpTAqHKVJy9Runef9JaoNr
phOUl9JH8EyulBBDruBaNmTRJ2JOziRH4Z54KRDmqepHJYIh1lZCtkFAq2LBKyTm
IfKGkHr4cNaEscX8OWTIhiF26hjQ5kvW9tDYx8dMSEtV3puKCWnZjyCPb9Wnu9Af
vHs3hHoaM8YXKripTmai08kyPtFPqPkwCn0Z++nPF877n4ERT5B+dg4yss+S+77k
fhOZ3QXvMuySKQ5EilOERter6I2qJEa+WkmOHFhZEXreN8/6qivD69ir4cRMUHEh
WhdpFUm5CPjWTyqlJBjFgA40AuRA72YDFoRC8L9SobfZvuotWwtZ/TjA/Tsr5YV1
3QVQyYAIHkpy6fN/iSNA82i38oL07UMM85ct7mkesXnOavlopJi6Zn+Z0IB+s+TT
+7m2ld/vDR1ymYzsT7qAwwtbeOlTYFOQi2iWT/RRZ4VMZh5dLOQLqohmUhq32DZ2
q14UyfJuB0EhkGcpy9YfS/3k3dAX0+byFmJkUtoLFLS+SWwXpOD3qzQRiCY+kLXM
ONvo7ppM0tzP0CQdwZ6NncY1m6eIqnHIePkDKsTP2H2Pzxb4/kuWZm5phKEuFHVU
y31X2qpN04SYPtyiWcXd/DrkVz/O6uyCmx9yeAnAwU5WEqzfgYHu0XiReQhH7Y6l
D5vhxGD8uXPgjR9Vfdyr3ZeGEGYuZ45YlYdzIjYwAp58yzv6M4Cif8t1cN1xQnhD
FSgVgVGv1CzVlTrDiISnhdoz+XCi+77+Dn0aN99w1RmZ2vBnjmkwEtGcyZTc899X
lD5VL33LRHngH/5MMsBn+pf/ahZtrYQfRtiMd8SnQNZIcYnJLn5BlOxY4oJ+jxGu
gppW7GdLqcBjKcN7vc3M0cNMoOo+pyu7XPS4Wog6ZGC0InleN2gwyQg0RP+imgVI
ar3MmNFpONMuRrQBVIR6dRuPlJy+CFKeiXmlf2kvLwD4/iZKVvXSP8Csg4gbJiM1
Zkc4Q5RtZGZSuxfo1TBw0ze3hcJvuJsTQcDaP8IWk2UkFnX3b/sUsiQdpagOx/eh
zeTleEjxQxin1V867WP1LsNkyj1erbKyYRa4ONg66UXzij81ram83pzGfMbJQNXM
F+Wbam9lm32wOSlm4X6kNpa808u92dgL8B8Y9qlgzSzdLo3mesuowcV8ZpozW3QW
kEyW709jOdOUAcidF3hsXraNY2pu7Z8ZkQWQLQFnRefPQvnqA7m2a36MH5mPwfVK
z43FPCPC2GZvJflQw4/MwoY9LOhcVtcdBUCU6IC2fG5bbZUqbcbDWc4L7yIGNn+Z
Z+y9vki9J+7nFHn2klFoAfZHVqBQY5vdlxOriN4Vj8Q3vOmBO9jvAa2540wjUaIv
x2T6GCqZUtC9dHyzAakAqzqe9l+ToxN9l5Wm8AnmBCnXnjeDQFOGw6HcDzIvyOrn
nosLPFq0+ZuQYn/ez6I6bkw/KMMHELZZBmGhLidLfPD69H4iCjJNk0YFuRmOqDjL
Zfsi9YjKbQo5Po7/UZNAq0DgFmRSBQWLgLTk0DGTVlXoNxGYNdzD0zoE8f8PMyll
LgTSfq9OvGgbJXpAadx5mO4SfyfyAfhPUvTR2gh/u1/n6RQUbYUeRFag2f34crF0
fIrBijiFiWeMEFQNlauJOPHJD1+RfakY91jETtu94Yryr+a94/ymb140JvxnTjNW
CLPz+9rhJbU8QO+MmPouvHhpCXGbglh3wuJr7Iho1itibrB7Y1m1XE14zWWac3JK
kBRGxB50lOIU6aDMGOyCD90tLS28/7sSth2L3VytdSiqtFRBRO0Xt6jXucjau8ad
sxfBJh6fdX5IRnwu0mcjlB5u1lbSXAm4c0nWwTtKYP1/UXNwOqaKJ2D8/wbQHk/C
wSfclye9666pHHt643E3ntj+q/RJYekTIB5epijFSMxyzPmz4kU5oHESY1x9Zgbd
aPSu2WD7JI2W0BWbG2baoUu9gUKWILsTiQlVIaJGRP9yWdckfOnvjCad2R8nvAy9
ZztXoEshAWcsGJ7QByf9JTKzQhLABH6k1Um1DQBrLaF733NiLEH4ECpqXXc7EEZA
ztgsIw07xgDMIIJmt9akLM+u9hmYlLrsUbPGSIGweS8ZJL/5voUIrh5JJ0S3L5dD
v7q9SVqcfZynOSm02sPDTFzMUGAcA0xQicz+4oIuEDfZt2IgfULBnhG4WVvyEYUf
sOMTiBxQJPJzJ8PStClsUqEl5cFh3dN3DYo8us8W5lxMRW6azExIgQUuI0XALBgI
CnmsrWGsFOEYaTSvscz7E3a1fOidPDy0IIiLqg/Ngza9hoxrza4uoEoQMx61X60D
k1A+rrw5I7uwtsLuidTgtJnh0Ee3i/7KFozjy8fyT+z8KkO2oZP3+hU3xcHuPayN
r+EmV4ZngWXbEyTu/eFbOkymcqKp2RaL4k4wG3NHIshpa/Qav4/A3zLcNOY5kZMl
8pVCYZ/0yBeo8f/AI9AiGHoTTxfzXjOIDVdujbWZBdpgnSbcAzjbE0/ZeauZwqI/
g2vrvChNUMdTMxPf1jIUM/ZkwM/2di84KlueZFGzGKp0AFyX6wBe4Y/D74oHHh+h
Kfpq0SAl7fyDK/2dr2hzFpszvrUTJF0NhDDPdRdgj824CBjZvW/ZRAWjXkcTNTqD
SjFEWD1l+eqVp3xGy6xbc+imf5KqEAl4QruI8iaGg4qea5c/BoAbFxchWYmZXaLK
6zX2lgeDtYjCLTryXxy/udeG+YzyLXqsTUpYmZhz3A8KrAw1wYhUJRwCJRLzZzaU
Ej8GtdrbvsaeEWXXyW9vvxdXZxNDOM1n5cSOij6jUbzcoUG1hfSA23u4LAjsrJOe
47vXc+jqYY3kRZfTNafX8M8QIAvFmjbm2KIB3AYNCiyJ1rkhEth+zd1TTiPqWrnz
uz9bro1wm2KAhSbdbBNC2VYXgSTjj/EmPICnIEtQfCgCLDKiz0mwZyqoP78NGAuB
XC6FYsSM2Pi5UgMmp3jhhL8atOoa2xXm12WYiQOw9kFaUzOsA/Ki8TXK5985KKm7
ZJp3iKMSYQqslj6KB2mpWa0N9JVGooqul3KvxIx1hIjuq/fRuZgE7l9g9R+24STg
OcIa3fl6vz1uJ9kRWBDHFYaIiUfdfcVv4LsoT5YXJ3K1BBKQCHUtRwFBhBjjXOwc
4+mx5hdQ8723LNCLWM5dK2FznJssfqYpaIgnJzf6HW58st6w+vkpWOghwxQKwUEn
hUuAGCiHRLui4qdghfRsiaDukCg9GwUwrPgKrvja4xQ50bGhTe0J7Oa8FYfdhKkn
OHWYkueru5VdC5+0D5zfoKYG8Yn8+9OM2YuS10ysdz2VzhNh353CE4gc23xcxV2M
8mOf9suC/mMzGwMHHk/ftqIxYKJFEs3dAipfqhdNDTrVOpVZi3l8iniupy++eICL
hlNcExz7uRExfzNmgvBvkLRWNFjdbL2KNlO1NglenDWw0dLSEcnXzYKxEOAAhJw/
+1L77NsTSmvCf0HSHCx0HOyEENjEGntFoxbuzPooP9o+xjC6jy6DqaKVq1b5s2Zq
jVVIrOqFLTyiF9nhGmgCjNqBlbcpbrc3s/Cr4pQ80FtNeeXRYLn8vWQBjUoA20WB
Og5p756SRHTutUOWNkQ9SuKSRXF7cAczyPKTSwt3a/2Xv5t8A3H5stWw/D5sc6wy
FYkFJxHTjZGF5VZPeCUPGwMfNT9FdeIMXQPkRYqEzHbzcwp/SmR329Q4zoCX+a/P
zLKkGhaffdpQDSSfLEifhN0/l5HH+LkqS9B8XTZPzUYSvBWseJivFY069bMjZxX7
z8mre+259V7ZK75MnrIJKnlDlGQyDDa67xgjssjl+c5U0644dwd6TmvLPzjAIIzY
lYib7Rs0M7/Ws9UQk2iOLx+vlhovXjfQKpWoz+/DoxlMV0pZPXStgtC/ONOqEiq6
TgZVaV9p56HaoYOyl39DP9J5AbL0UyJcelMGKvAeM4Cfsxsikjnkx318iWUhUR/r
JVM1R45lPy7r550F6L0NMfR63Zbgy5r85nT2lo1IdwhfniFzYchTh36z6n2SIcpj
/m1lK1DLf3ehq560FVkmwiO22teJoG6ZEFXYc/BG3jmpT1CTAe0SyO4ysAaR1roQ
/OidyOjLZCqjHPMNbWHtG84ShmM92RxuPIMFVwTSlmnHv04tJjf6He3oBVkIj/2I
p549ZkRLIs8Y87H+7xx76p8eADj8eyJMi2EgbzDPPLczI2oLt79GVmpBIp0JGiLb
AelfrRrgn5G3jKH8VL9a4kagZyfHUL9nAJH52m3DO8QrmpxpcrJgggu4RAmMJrNA
2nUQj2xQt1tDdzcodFNsvJ4uv6wZB4VyL4FGqROm3gllSOaGE7hnIMMlsLfxFBGm
gChMBQE3SN/ZFyvrIlDti6qGAMXEmF+harg2qAQC+mwbBDf5UJd52M22A1bEYvc6
mJ7LuIs2dfgTb/aCYxLELBzLV++BEXPpKIxSFrzf9vQtY89euexWstCRAnsGxLeg
9KXnLs6KH/SxtefeEkKpWJFDm47hJzG8/zgnLt3PU2d6T5zRyGUTNkc+MlTYaccr
gA4h0mHmRckLoux+KWIQ7aYCtaQ3qIrsYH5zCMBB0iw7Mi9i/OOjw+deftv8X1Gh
Y+eBSoDIjKxo2t9nXzuvTd81wE/3V3v906BF5ss7ZBRDf9AhWxamfNtk0OO95eal
X1FLWgJXgl1FqVBA/gAmVtOG9XemFT6I7UDDTD2KEYhaiiek+J/MS/YFhPoLd0js
9XmiuqSVk8dggij/MPrVboh5RVOcDWI8T3QdhTOP1BGIcZSIZ//xqQ7+qB8siga8
BbbYXKVVnG5DzRZGfPMNJwkmfrrn7nwG1L2feqO0uRE+u9QZuBomCd02aTUQh1lh
raw92pGFw5ZgzfZp9rCLsM7r7kZoaLLlde+5p0yxH6E1QH8koWoVv5tr78BnbzYi
xC1jAr3O5AeuE3hnvoRxtXJd6vaBSSOKI2c+f1FMLzhco0hHIhbiKE6Nr75JcIZx
PtOR71YqaQhGEJ1YvG7wYzy1Fv+GFYBbx/CpxidH1GAqJeez990k0mnRxm1lGZ1P
cwjVXER/f4zqIhZgbjVvoUByHVlH/KtipLp9l81Hw+qkI+VTnH2aTPyI4ATWuUXU
Hu1E3U0nK+BvUa1TcvhbsQUVKjMSAj7DF0e1I/zDaNGy5briZ5gnx+su5FJCZr9O
fOoPPApLwpwtmTkdrCdkXejpUxHkvRdFX3WVzx7DsD63T0a0tt+Ww1Q5EYLha92n
MKke/RuaVFcK4iLCRYPPAbUKIVpHUW5oPdpQrfKJ6Y52VRkv4xolEnEwyuAXGI9D
SEDYZr1hn8jbtqUU11hSDgMWmJCQzP8MMjbSqbOBHvm1ON1gpFBW/VAcDfb2SGcT
lzTawXhTC6DexQz7bGvA/XA4ue8uTdsCtlnBDIVnxjzRS2gu/x/beJS5UAyLCeS2
VMaBjJm5u8mpRHrak0rxdKUZLfW5fQu5O8WaD74R6NoFZMjjb2p0BzzxAZ6MqS9X
kxjpv+wqIdMDXQHcDT2lWplJVM35OOMr19XZ3okmFyynmpn1Mnefk/EsReM/hrR7
pyMYH1XT/9DW+LAGqeVq+kyPHm4xRDuCiuqsCaLdXn/C8CQkVaUudaAr5k59CkRH
1L1wtk1bl3WkLFlN3ftoR4gaZcY2yW1OCBt6JJ1AyqpHhyyPZbzb8KzYV3itvTaZ
GayOT7p7PWXbNgddCmJWw/PfQxqhGGkrwttCNWoK+hT9CKE+l1GscT4t2yuOBppY
gyMzLiJnZLsHOhMWbOMRMKcrezhhBHQ8BE4MuPBD8Q3zwKUugMoy/Grsn+ayYs2/
sAo2VrCIDtZobm9mf2NOUE2RklfVg2BYtMUiqYERvwEvfR8SOJmgUxRJYPp6d1Tw
ISw2SRl8hPF8ghkw00ECC9npzvrIfrmhaq6zZn5a6kYGaDr7NvRUQb8683+iDQY7
DPgruawo21AezBpLCidlC66XsHGBG0JBWf99Hie/OP6MovamVfY/uK8CTojvLZZ1
pwR4pjawibcFWRKPSXva9yCN39yEnLG+eMb0qcT2O8Zb6GZ1BoCpDXD1ObjXq8Ml
AC9bXzF1cQxx5ks0skbVmN9AtFx3buVlkwlOIj3m7Os07UVYV4qSRI0nXQiCGD3U
r7D6s2Xl0ccum8YA9e7i8PGB9Um/3Fe+j6sfGYD+hWN1iB0+JotcFp+v1dG4LmYR
iJShzMTMOpa+TQYrnbZuBQfTsKcI9chrfMYD6lBXYXBUnLRGNk3kRl8Z5uOw7M3N
2dSGJxcTE7ngyxylBfeVUhJy3FriJ3zUgNaGaQaelEIE73ROGBVGU08Zw6v1ANFY
94r6Ez2ccxDBZ60vHsDpk+enLwG+Gvi2DgzMlAHWESDg63PstF9Yab6S9b4HzUtc
dbsEh7Nwv968h7OrnSMsJg82enw/FP4nPBcndodNs87oxe5AGWMZQ/J2GJ6bJ3Ex
tbQ/2/rkm0W4p48MhoYBbZ3B4oWjrwcQmYIpmLwr3R2aq/A/CgYB5lL8cMUyIaXi
B99MkOMewDAJy6Q8998TaA71uoqrrtrXNuALuGh00fGzzHCe4mBHTM0hepvQF3Zd
wCEG1LokbBBoiCldsBQEOQl9rFFL/U69SAqccjtzI25P7U1daLF08uhLAOjWg2/h
kKyosS8zKGNsclg+cTv0VlOObTmk0pl2IeUrUYO/N9S7VJUgVE79EUubv7pxBOY+
9TjtQlIxFhp9qm2BwIPqAS7sCDDoXFFLTz/LaWdaUkvJ0KuZ5XGyee2djQrBcAs7
yOpgkxtwS6bztsK2eQj4wYyNno3ChyS32U+vLZOLhRIhNR6NauS2zUuFSCNp/Uhp
qRmfzPdFKYamRMd0ckCSh5KIilBE48Osb7XA3wN5UrVZYrJjMkwIqfuzb0PDk1B+
2woUg75i/iH2Tcnf6o8ZuFwljF7P+rknGLbTLCX26QsPkIX/iycXms64iLRM6T5Z
/083iq1q3+x9NGaIusl2DTDefAcGyFXY1rZglSAZgl8NzzSXUaP7oR8NQhk0vJ54
3DKsYy+fw06JXuU7vP+Mkhqw2Ye10wPDH0SaIlPy495CYOTVPrTVQ8Ora4lKQ2ya
G/7mPQZi7SkY5+efTEKn2uRvzjwFGf5oGOft6fgYDtqUFbz0A0yJlq1C4s5324sN
cPsx8Jz/RcezD/hlHOEWc5h5NL7/fu9FB4IYznvDJHM5GqybVxQhHynLkh87S5w8
71dEnzEIL8v8PsADt891WSHkYBKmCDQt2RUHz0eTfTD/adRkjZWaX5QHfbkLfcz0
diIUVxRszeKong2qxK1gbXu/iffa9RtD+zR1xX1pcuitrfyBlCLEcJRxX14PeX01
XmLuqRHcSmAuD/mVmVdwJ3cOtb7/5+MqGazhWfe8RXKpIqHQqyC2A1orQruLuLv1
Jmkb1qhVRQp28gVJ3He3IdhUHPUpT78x8z1S2svl15MCrmaQkwkinUHUiW5a978e
fL1hbm/ZKimPg99A5TMut9xO5tuorPdIongvOQ9Y8e8fQy8S36HMk5hrywwWO8ic
xIiVvjSOOHD6R9xTbM0wLciIVbb5QI+MTHEubZekHhG98hZD63R6EYDIF7YCH3wV
YAMVzGo21U8lYATkNF3CiAU3KYMnpDlVsna7JbhJjH1QLglxOQ4yRhP+nOXw4NmB
Q9c+4hCmA3FLCcu5E/orDDHE+JbppqhXajze9psooknwfJmJ6L9mxrJ0b7iIPj2W
qdjsfQeg7fnSavZ/GXTOeZSx3373BCDrIAolwty/y4fzDaKvdcWsb2s0t/wQMuhn
uS1wBrduTNw8S4N5NBY8+4fGwyapQq84AFcHRdxir/bWL7lce1079HCUUJsTP+1t
m0ug/q26cmGzZIBmrvgUgBae40xeyml/1Z5HC5NrAcSRDXI6y+0gYseVRUvZysol
CEsZEBtga4P/Rp+jD3yTs4G6kAjZ36M0RhXhUgRT28pjgTxYUTrtjVgvimCl1IRx
GAOkCH9SZPpZfke8hcTMbEPJ3RofHE5UhT1/wELAgXd/SLJIP5Uezcl4LUygz/Yi
+39ma1alYmQccxEJoVj3bcSCDN7INkmG8g4AdO7yLDd2qc3dsOCHwB1vT67fMm3h
VpaXaW6OJpVVr1V1BGGLnSZczHYUbT+9NnkoMKCb8uAU2Xp3P+U98pYubJyBPcTq
hQIIZLbZB+1Nz9oYWLft/hOPRQJJrBlsIR+nkOxRj6i1s0bcmFkI7yLUDcCmYv5M
dObaOXqodZxhLG+rti/3bp198ljUFco1eUQQYmHXa9Vndf5VR+1OKM4ztKH2l99b
Ft3W/re/THmYiks/es+RruC1vpKWFH/tmU2VVwCnrkUBc4b+OcSVyssAMDCbtM5Y
zqJ54gxNpmDxCqJEqPTgDS3YxYzZjqKfMqAXdriSKkxm7WXPZQr6BAX63zYdqJ1u
aNIxf4Hn+gz6CD0OQer3G9hTM9ggCEEmClx6vHrRi/EU3vNBXDZmwuqZogUQk0oX
6VoPzS+at2tSexRtLjWVCR6tAO2cEyE+nc6EYRYpVqxwI5yGI2XPq7r6rPDYWhCM
Tmppr1o0tpKAFVQgrzsk7shiToU/+KJYyL7eVF2oyHynt7eXnFyjz5wsEYQshY9B
5PtqW0GwDoJkf0rFGaMJpszIDezRkW4DNiXgS6lIrQfGrCB35CgLH9kJcyXzKVxs
ni/pA4EZgdssth/BtOIIyBp4adQIx+xMMDQGehvNreMpwvPiGNuy1V+edt3h3sj1
+fl05NYBbfLix1i7ZAhLAmZV1wyotxSJiDSuXmvlkdmKGj2Lekz/zKF0JwywXuGr
hHGuDc2z5clAgBYrmre6HKGbYh/bNrGXzohkvhsTgeazewFxXxzCTSKni5bLrk5z
UFJht6pMAfal1qlv947LbJ0fG5cnI+XQTnKftrIT3AGjo5nKxGxGqVcscIu5u94f
RbxMasW5uiIzlRgShZmv9fBrdQg639m64dSzb/9WsYBC70gEm98SKx7Sn4FkRydC
3FBjCkQOEg5g/n+ogb2bVfq4rx9lSjj240OZ7jhHUXz+rb3Q+eGeUBrqaOul+F3x
oQ1vaz3TSJ0EYrfEBuFGxKPIaXACTm/2805m+cMmmx9nd4T8r4TtjSjl4QSyS10R
vdkkZFK4GWAKsj2gL5b7QwfOzYon98vJpQg01PfszvsaqV0clkqtFvtaC6ba+NGd
bX8KJTNufkb5y79Q17lIUckBR3JEsqpfbwQGDp2Ot2QV9dHSvc3/oo5u13SBsucy
1isbIEoQChAMIkZtERoi12qyXEOOm7GMsdc7/4mkEGpA0XAVJVs/Cb0LzauJDHHM
wd50JdeoAjmrmMzGOrH4vPDGgJcL5KbiQq7nHGUcf06Cg9Ktx3dP74Yo/lF4VkKp
+yROkfj7+H5KA6V6+vKgvu1fk9zkzRKQ2baVOP8meQO4MNzGAqKdXTmFlHzxSNN1
RlXjAcTDEW8vZ0OdgMitocyPMe3zcue9lYFCHLx7FzZX1UAoCpkfRPwJrOldc0vC
xqzGtGe7LTQf60Y8k0bmHErylK6k1E+cfuvE9aDNEXiJ0SfR+VWSQYbRTY6QXjWt
+v85/l/eKXahqEHpeHTgPjdisIldhaRtDG8WjjP4qEjYCelxumLeuVK8HFBYwnee
ui+l/s3ym0fXnYytjk2oVrn6oKpVDKw6MxEluD3SEE9yZUYAqyNhurxRVQKJZK6+
Jrp/WSpGeBOGkcSOdjTkBZdIup3eSPRSkXSjy0SE4nRb/cG3rpNYeKBVjIOTGDwc
3GI4MFtN0GTtlPDzX+f4xkVAKuM9gd/7CMg8HeRhqd7eBn83AFPLao1R/AJTB2s1
q1XFUgqNpoVeCDJT2xGnoUppTBClSeUgdI/VGLRpU0pKYW880QnVjSGzJ/RBaxvI
V4v8JwD7qtQDhG84c2eGkn1GPUkEalFzVUbGameiHg42L8/vrQYndF6iwe9ln9KO
w/s7wYRJGCPS3vt7hAG51cyy8/Ik4fknYrGCZWJMpJzktSuiTVXinKo1GUjCV3K2
rgMXAdeZQhYiyO9THW29aUjyttOxtQHsARILj9L0UNRAHhZGEovjM8J5quIKWiE0
wQ9drRooTlUFAY/Cq6xkBimqEzN96myaIBAaNFq2WvsbxAnpQpEO8TVZ+WZEGXrk
AqDzAZcWwhX1XnjpXCTTORLS2AjJN3uI47Pfts7sX8Zf0qA0pR2N8GGAz7BERi/q
G9PIqVceXRK1ejJL8P7IH+MvStrze+K2R8COP7pHyL7OxWKXJAqlRYXdVk3B8gaL
ooh1i4EUCydMZIZ0v9TOOktMAC0HzuXqIbTsleyWH09LTiCsZ6NdNE73H7Kh9M/M
JSc5ElNiC5qUtucsg4tHdtxFFntJu7KaHcKu2e+Q29HbtfeRQW/46T8yPRF2IpfH
M/XMyRmcLubzP1q6UPXQ9CIk+gjdKPX7+zkle/9CJlfLg5PlWEq+GuCFWs3culO7
XrPhkTAL9yESGADKdikUYReymAwD/oaSi+suEZjRQSDV3XGEjJ9be8uwyOWJrbSS
GvdWp2IhBEjXwFYfF37vSz47y8xDw2s1fgRSFXUEy5QxrjxcO9/+A/wzWvOlH/HU
HrNS3kSaKHfy3V31bN6zZXSUn3XozTkd7x62fTTrQfz7vyRQlsNksEDl6JJiz/VT
kWG5gm3aRXgGDfBz1ENaDewYy5QfY/Yl+/h0ntN1qnU4X0sdpBM9DIgNxIP6OvpY
G9AqfAyvRRIgxmTifREPihBHb5ZHgWcCbnc13VwJgBZZdC7EanD+9j/AH5xrIqRr
zvpEsDJWUbOrdSDP6U5WnBDZhro2IOqSeoTDmYhsaAMyKmVAXC7/Mj0DuZwwKMb+
9x7AuToZKdiSs5gftGWHNocHq30RtScL/Fe5Vs3322BgBCxKXceCIjN3ussHuE0I
zuii5etEsLckNyTIBQVSxiAQyRkgEIZy8KuRimPS7ct+4dg/1kNHhIC6hWvpkg6h
qkKNAZ8En3HDxmD1VPeUYLV22rIYR5Zj9YETdWLgA8S2ZEIu/fvjBgRD3TPQW02p
lGRih4UsW5IDDOD/1nwMgQUX5KkcYt0nNfaWvDXBoCyKdg+50/C42ipOjdv2gxFW
bTOdRbiix175Y9KYw123AQ8j7o0ViSZ0WDMQ8DFR28tv9UB3uI8p+ft7Rd5qPIBW
gGBH9VgN1OquI+nI5ghmnGrNhwadHFLzWaj5QAO0oicuFH8xA4SSyzyaIC/3wV9f
/dIijRskQAdo9HPVJ5GPHRVdj6KPwF3MhPO8KwSSP7pyXPhz3aRZd1/7myRQce0a
PU93kHeAvdGshcTHJHdkmnbiR7A7Lx1rw2L3a65T9f5ZhZsio+hVfw6LUj+dxwyT
6kAxl6XQPZJ+WBtuXNXAWLB7vOK941q02Er8PGYj+XNLe6qsihZrXgfBSIxhvs5r
/xSbxgNoI7obezSlzojy8lVRfr7bv7fIEOvVOZO4FvMdf2smP9bu0CNz+wXLcjlG
NWVg3xeY5RnP1P37CYfiJmpthVuZFCF+J50OeSpYpOKtgfPI6pH9N8EMnVPp8VZ/
T6YtfBYvLksZXNdUUrqV+uHTC62baVrLL1w3r6TGpgLKZ87Ifz1g5i9HqjETiuRM
y9P4pGCHhOFejh26lY45WbQeM/+uWjBReXeu5+LsNluK6WJsH3eh133TxyQQL8qT
+JMxxKVCz2iOU3mHEC9qOiJ6ApS78UT2bWZcPt1EJJ6ivo90/slEYMpwLrIbPRtf
wp8uHHCsHOBaLcw9X/KKn9IYVbKqG0tYJP1TcZfd3p/aLobvXjEBvl4zWF7ZQINW
CHHc/CVb8Hv+DdNwBrb7jNwoLSVfYPnMu7Z4jvugN3vm1l5dh0Q694wV6oNqzB3D
r/qTfZIKBR7y8+o39OQTt3bUfATUSI1CNQ12eYOlOBKxg1Jq8wbKmafwPgb9dd/K
m5w1pgREEK6jkM04Ow7jjtIdx7ob8Dcyes85oHP7BzqBpnLT0rcJzmGob0MnECDa
CTPAtVcTn9+yUTswHiDEa1WAPWERsDV1KXKeLK3mKHiZ5MCvOYUJJADGNZVLsEUQ
evi6mOsG/sMW61VUXfNvSo/DEjHhcbOZanRG8VRWWiRYv4go0W/nQf/hlbn/eqZ5
RK+EIkgfaIImyYHe2oU1TsH3TcXdkCAlMfcNM3ul/YMD/P691G6IxeL4hoVHb+Mr
0kg6z0d/AWzCN5ILDPYNwu6RnbEw6neNViT4rrBu5X+5inBYURSsHXvw5oO3WYph
Eblw2l6VrFl5BBpQuorXHPEC4O0LPSEvmcv+XmHcIg7XPmD2i4e3E2ZaiKSvnEJ4
1BM07ikMJCRGe639kgQbBCQsWPKFfBMLLU7amQsAT1EKzsFUHNWdvJmXeQfhiDs0
/56e/C0ClupkDnHt0sVq61F5p+Xux9tI5u4VSh3CV58XybXvb92JHvET22Kev3o4
uH1bIoIFGlmPWyXOKX9i9T9lgm9IfYTiBZieEA71MZNjGXe/ubHtDVG3F0lrcxUg
ZqO2HLgZZgpAJKqE+XO9sS54vgU44zUnAyPBuwXwtupARkQnKki0Ay0G/ysJcLvQ
0YZkjkVCxYbbShOf5h9BNR1cdE18HsSVfoP3Z8rXqClDk098BI8GzLtyl8Bngtc2
G085MKWBWA357bUkYpGOkXhFMwZECWZbHEyvE7n6S2IX/fJE8fngzo0p4MT8NASh
NONLtT1riGF0RpmQ3v2b0tYm/h5KAZZQrg4ZbloovAehmmfLi5Sjj769GtGitLiY
mipiejeMF/Md+TkSZQ2WKdsd6sf8zd7nJieVCwh0ucGA20Vx3/r4Wywk0Y7SMMIU
kJDAHmCXOzcZXsSswjM/WoolXxGqeX5hNsVRfq+Wh5vZvqi14yLP7cxZyYrpI/XC
YFdfqN2j3caT7IhoDTUqnUbkaZZ3htCr9VcsrXsH3IG0WDSbHGZbUaZro0PEzu3g
/dtVsY4iDY5pBn1bU/3FGpGMYu732etbiU0TePc128jMBrJ8qRJWVOAnEXtMl5xS
eZup/LKFfPr0FaUSCm48Vn+5Wy7LhOOiEwDbHn+NnHfESUMdgbUP/O+m3hbpaDNw
72KYx4rUopwuisqRMJzIP1se5nlCTU96V9rYsHy5PMyUbhFAkFW2RstpFSiXLJ2U
RtDp0mCifBkq52cLq0zHngcazMVKHHe+MRWRPJKG23lSz0/vMG6RZ2HcOvsXeVot
8tqkur10GroTgIoHyjXZF7vxHoms7qS2sas3ndLafijaY6/8Lr7RvvxwnfZovStS
ITgne2dJZTFuWJomnev2/WsEIVzkKhBFxB14rtkJixx+MFx/qaXwOAmr0LAi5gNF
xA6+nv9cl8JJiHYngUg0xcqnJ6zLIxBfU1q6LPG41YCEz4LVkv9UyG/DErJtvCeM
MXkMtAuCurv538OdjjhETuBzcitGAouL9UFLQclt67sPQIplPzSNA9/gL0fAjJKz
7zi7MT1JiM7ChHQddogOpI2XHug5DGbnu31+caj+jspztR6f5U5HlbSoiGTvbybW
vzUocx1zoCI3Oh8ytieQRVF1JC9MzETC6HMLHXm2Qp2vuX3IZm2F56p0jrlwLq3t
LcYnKkWaTNy5Vd354A4iUTXlUePiS2OP4e8DQScdofyOAqyAakk9PtbLL6MRBXsY
41McwTWFZ18o6rfm5IpIOAN0BFUHHUTYqlv3c76kJim6QAY0AG/YAWpMnCGNzlbJ
0cYDI0NPOUOTTh9TJAsykhhGZdC4uMS8Q1ElcMCFNUa51Rj0REzZXHt4BlooBFfJ
eiPQFFJ+fxW770SFC2FBD4hJVAYuV/3pZIEG2gwmT7LHSdymVybC2dMqtbY3MO/H
xpQKzqxY8vU4InI65KniNmVd9jTAosEG8Lrcu3iWYkNQCJIZdtPvVdOBX57HsuAm
GcQRRL53a82bPUl+fTlX5gFfOExhMkZyh8oAMOGiETcAH1tPxh2WWhJPzRrj5xhs
Ha/zhZUJ/LJv6Fj5AuQKdDC0wNEN2pAS7mmh7ChgXezNJUUlTJuecwDUDVdVmETw
yFQ38hlliRJlZCn8YuuUKG+bl5VTw3xSDYOD20N4VfmxqeyAPyIzG3K3fKpP+n0T
2T+z0e9EIQ7k7R4IAlDPnaXEZDty4xvsc4spuhDasOa8zkenvLw8S01XqztU8dEO
TiDf8wTEZLyVKTVD6Nohtlzcijl7tS9akzH1Mf1a6EVsUBrzdhLGr9WJqiAtW+7O
d5dmtASsMNM4hjxecjMY38RtxrGNRzJx+kwLdIVa6HWH1GwPCs+Ly0pL+JaTAPmd
oejOhdiZhuCtXbK1SEx1tsSZGJThZKjSy/o/m5xXB80VH55UeY1qowcVFGiffmf5
CZsijoCoP8xXpL48E1HSSLeY9q4ir/V0w1ZB3bm6zY/108xEKS0Tgg/UUW010fPH
6IGTZPftgWwVTLRpbYsbIT3EP3AwsYzWUMw6xk+PVJ+uXNYSTkpDQ2Qg/TT0AjfA
/xGtzZqyyUwWurf+chKxVDM9ur7AN6nc9oDSHAx9hhy6cbbY+J5sjWjf6ho9Q8yI
aAYBI4RGht+NoT+JRHxnVy4kHQFAzjOhcAniBCmZSeIB8p1EoZ7EbnHCRRctYNES
RAp4OclFdRRP4np5tYfRN2LvHEW82AC6ZT0T6vtIcNE8Y4Tw6aAaZmwPSPm4pAGx
tDWodPdvjUkqlWI4l7SXL7XtaRv3kjVTasCNtSEzxGxF9rS3o5sBTRE6jqAsoXl3
a7mngRtrmey6mgd8SWP18mx4WGswmyebyiH6K2OOU3VayJfbXiIJWdY9UwgpObYj
czaiyEDn8wlvhv0JfOn/ab4Euv+dLVb8KxUnSQ2fUzlp0mAOg4/ZFcGtPWuOY8VS
ilYva6CorYp4BssawXXzOXAseVWrWKuGA0utcS9y0hG+TdTHvlwYF2CYCdxBZSq/
tgzvznqmF25b63IqUv3YjK1FqqCy6ysflR1pBYdXVQhneryHd9nvrskBn/meGkO+
FlKpn9gSWrk5UemB7qKyI8B149rhIVZaFEv6xPUBq5mxGneF70LU8wExM8MomwcK
ZiYdvAMRCneyhdUeQsqOjUtfrHUdSkzbqmQxPTjzypZWf2I2kHoXvn70TsmcFQe0
a0qWXdh8IJdBvqxo7WrEboHUjbeDnP6x7uowgsjJkgT8ruPuCyPBmOi2280iM6Ly
2NK1wg4l8b+A3VlmtrBZ49Okrq6iRoQk681qC068YZCQcFQaGas9denMy3V70lDG
+mdBJXMnN2Pi/8Nzu2pJ3BHgZ92TIKQi75awoa13fASJm1ZtvGyYHKep/tlR3Qr7
YIfQxNCwS6aPRNfTslBthpEYdNeJQeiBnNKykj3khN5pqVz1FfTq6PzN/sbTRupC
FvcT3MNYlwRrtCbkg94cGka8zSsdtCPPxyidetxA1bcnBv57mqiqF14/coyRPVGi
l5ZPCnneXmY78MwEsDAMF0RYfaFrAp4KCivHWcVhkueuaZ/gh5tp2m8K0ycSshrZ
GAdhuWpccAwklUHTO6OQrPpQsL5MbbSfwgOoDpcAtaiz6ciCm5BO9vSa4VJPnaSe
41sSP5mZSMMgyQwtjo0vgzjabf63xypB85ArMJC9Ei8kSELg4S8dAPC7A3/R7osR
YDLFLvvJtqqyxvo0bAaqlmZiaTcpck4+QtAtutsgprgNcCDnTIyKvgP0378cZCPE
lH6TrM9zjl2iIh9KjhUAXnViIpYrjrKLEvdT5JuOPZEggufDDUWTo4Qg4f/wUAfL
XpcBiF1+CrvEJ7MgNyGcV5x7bJxu8L/g3QBV4BTSQZ3yyjXBeYIBn/gJcJVmwzq9
xcS50gulZ6LcBHN9hGMBKmJ+xavAnuzq3U/YV3+6TPvqaXu+3Vohje7zv9AZ7d9k
H+5s8KYP1uf4O9sYJMsvgef3icggXLYKqji7kaXyxSC17x+yT/KYz4MYA6wW23UW
6D0wtJZeWI/73/qcDIw3Goe2bVidQ8XLQWiRuaiQfTNs0gWeALv9+vL0AznoSKoM
Oe+u9m6pbx8exol7jvGrUx4pCfQvhwxzYhVHxliKycvQPl4fsuh+ej3rZox27sLq
0tBW/N5tnvYjSl0AGbAq6+K3JmaE8OH+HDwtXdjXI/9d+dGVP4ngO94ePJKf5p72
xbfbmwldqlP2uhgen/9m7KVST75t1xf0mnPB/0zI4q5V5mJ4ZeaeMB6aGp8kxKrl
F8xO6ia79p1X3RhjigISwIVsOdA6ULThChngPLtyqa+YORvWDub4XCl6ONwLemsq
4pqim/e7CMRxxijGm5gEGnAyQ5rjpmaGEXSR/hcd3adaGKmMylED5o/vRG1M5e6g
EsBulkqxXkuY+H7h7fQmN2EtVw6GZEuV5GZ7VRRyeENozwHMKMIsjx7B8ipnOhkD
TXJcwKzfgd/oNDS/U3yPMe+5fftfUM2MDPVfyg0FnVJ1zF5qhJuMJsKFqx7xl5fZ
P2cuT+8HVawLECxA6kCKVnrrn3UNNEJT2wgElyDs3RuKd+mJURBryQHLIZATh/zL
kREDxjy2bpj4xKGhUcp5D9I/Wg7hGxp1NwQIATv3qxP1IVKOWT/y2Jm9pDp5Vp46
ynDEhDGjU1OgsVgWRyyKx87G16jPhBUlpbJ6crdBDZx7H1YTHKSFSks3kBPNR9QB
FBIfSlmxkv1tFP2UkPB3+44ebQWHR1YfI12gzWjA94hxuU9XI7jsc+R/ApfdjjBV
bfQH9gbnIiC0CNum8l1saqDztYIVgupkJ8dilQ7tZZAjxCxCF2/TABXtNJPEtSSQ
CtxxJROgHov+6wAiVv82RPkoV16uAL6tnOx2R9KhM6R20bQZVH/cHeCzkXEvksOp
VKPcv48E5NpAZfGP+L0pNmCsz0qS1sI6rELHQBZpy03/f9j58sYwFTMO+qJhHN7S
GqCPq7FGPx8maXRaHiRqYynzfqQoAubBZG4GfBrFEkB6SaQ5jWqaY+yuqYCWobtO
xcUxDM0CxclpkaAvK1nfVCZloU5N32Z/YM0jAr/XFJAwEIpaIANQAIT+NAUT0cyR
cgUGXOTJdDdvCFGr1p3xx0mh4QK69+WkhNvMJU06+T3MrXXOgEv8vty36xJ8Psvb
f8qQS9D0O9TWIa0yuyfPkJdr4ogrZ4vMUYHKaGnx/9SWxT4Q4XX19YQIdjOkHxvr
m8wwLu93QwKLA+TYhl8Zpk3QsJP2PH8SPOzrZdM34KlHAYdhzyrYlTiL2+QWE3HN
HxcDccj073m6KUtDK0MdCHiItB3kr2ZsWXCIFzfQV1Jxq4XRJeMaYbdNstvxSBQx
JsYcvsw2g/FVIKqzSq4pSDcpuSDzaoEnpZ9wzXC/Z7NRSoNOrf+zAypVEhFpARW9
3RyCwv5x41OM9bsrCe7QdcNLStNHXevc73tz2lui6Tl28DhvyGjOUrueCCwboD1f
98HS7bP0qfMzDPvA1RZYyoNWFMfC9a3hnA9I4/LBc5y/fy91bR1d6Q/+ijSBab2v
YeM4vFwP8fUCeU1NbeZo9dMxUSZFufoqwXavKwZmjrrXvlkyiP17EQBtkZ21iSYj
rYawJqbgSmGIcw+mSC/FqznsLELtMJT74Ofxaj/lDXLi6759iIjV8jZyrvS9+20v
smk+tn44n8WioSnobZS5Vlo93vzKCbPapGag1rLxELrTtF6ANoxPVvWBihHCzjfJ
axVWR9u0d+CrcpO47FC+v/szdz7qF3bk8xAiRBY6qQ9xutjSkeneg4RDQes4YY6V
9x66X1Y8P3fZPw540+NX9a/qRGRVzW5u8JCOdzU4GS0jITvE9ekKbPJuPzyu9WYQ
StTrY7BTZOk3unRY4DWzm/7KOji9DLgCMDGRqwYTVB4Fma3DG16384PiKDs72lRR
6ovty40wYoO6yWlCOhUlH7nSVc2bwyi/pgFinUGj4xH+g42mKZKullX2u9Lii7NO
0gCdYwTavIu/xHc2Ei2Sh/LOYPBnpx9LwNSmE7NLZW1FfF/lkmXmJ4WklBOR9MFz
hEc9IkVZDwJw+NUyB4HtjNu8gKpm1k/JzUHynDjojyA1fjjv/pIaFFylDlQ0Eim/
tpIdkNJxtHeh+BNw3L0PBAvEXcWsfR1A9g33VcCyKUyRtxL+v80S7cdySXJ8rjWs
7/Qu5NSYd6qjF3+o7ywzcaIYatLvQbuhspovtofjg+vrddkFrVPmLxY2KM+2n2WY
1lXobn+iRZBCwO5/XdXFzsVN+eUImanaR9ijPsoyw09+2ERTAsLaflAUYFtddotm
AGmrB+ZRA+y4+B4+R0swJsiSrw+7J4RY6ZucCl2U3TJS8G4lk0WNG5Dsipzdtoti
5CZi6Bl0+5YPaEJ7F1J8uYx4suafPEJJtX0jSBNlmUqQkk2PNzB/s2yeWxDiHQZs
REDFzATtTZ2KS7XmA52og3psgsQQNEKCp7Ezj806VF3IVPz7w1xOQCePlNLhMZ2l
DT/fdLrNORJS+eABJtzw3YKt+JOec9qXUm44tQ8OxUtyLH7FN0RM5xM9SZuRUQRd
t+3dGeHQw/zbv86azcoCizQvivEIGJaIHp94hrkE3Nx58PmPckck9xFpSsRuyFNf
FhG0ImSMwPZwr9f1jEam8womzkiN0wRnvEnx4E6q0JFMQdLGiuSK/3Wr/kqP3l5M
BWbI+Hgm0X3XytMIDQoJBizRrU55TRfkEK5h6auJUH4kIxAnm96HYlg5jNQrbHQ+
laEd4s9HIEOznHOmGhhDof26Aobus1/EffP+mxceSvnaZCNn9WxzrZVYGATBFztu
RtB00F8GBohjfYNMglo2VMQyAKyOeEHBIG+wAY3Li9NQ+NKQSFRmk9EFybGePmGL
c3YDkCMe5GALc9Rv7Dmp9pA0oNz/2sX5AB/BC2payq0eZ4QuepT/j5WGBAmXl23H
g9+uuMoCE69M/LRVvRR+HbM58n+KLxtCuC8Ts7N0IsPLZpefba312xyrkzYO5Bkd
LsH2UZiEelbJ+keAbyh8hIhD+Olqct5aXlrJPeWwq9pmBQsFvM5R2G0Z2G2OPOZt
BwFf0VPe/n5NLJdP7yypkQ0Hemrjb2RHohr4XMJWt/SwNxt5s8v5gnUrf98++kcb
0YBkvD85xzFMTtp5Qx5nMynT+iPAyWLNjHiWA2OwLVOgalXyhlW2aS4LnNFQnYr/
cBOJJlxAqPzOeE1Dmz0Go1xqD0E258tuNcpeuIwI7cf4mIxB062J595wB9sLdYRJ
br3cLhmXpsXUUuSJikA6rugfmRrzoPMkZXcmvAZMbkTdfHeeUZkkkSYCsGMn//+3
pM3vmZ3klUd5wBLNty8EPH2bAkXsJ5Khfa0iJuYq+tN/Or0IAGuo4Q7KkvmlIxiL
BTJwHLyF1dj45bkBR0mzqTRTinxvL8Qu+DCJ5t4LdGdz3cA2sSo644ms+cEwg58j
2hvJym0peKu9Br1xmo8a0+OWBPJ2EDiekFJqHK58DE/A3TkN/XA1meNTQzGyaZ5I
i1It0z6Cv97PGfc6Lab5jM2X+hkyhTqa8D67sI3B5SDtE/NyrzUVk9+Q7VRfziV5
QV+oPd9FxHTjw7wzajTOaAmjGyTP/scQE9FtwryRYRwBSGb5OhFoSfJyrLNJfqWG
SgxwB2zH8Njlm4UNGNFRla5No+n1aDJmTZd3KRIt8eaRD8VF9Ag5c2I24g/+Gf4V
oncm1uGTEmlXK1YEVtkwkALlMLzNHBFKVvECFH1CCEqcZaRQOWW4/tjuW1dImnEE
cLz7kXDMY9sPkYozErRjQQ39tgXuIjCGNSip9OGo8RJ4L0PA8XQb7qw555gMuiIk
+0cKNYfcae9Gz0qZyaAjQNLjsX70ZO+juqU5uN/g20LZMyN12mzQ37k8vi2Vk2VE
w9nKhj65f4tpQjNqn4UxgMsUC0yG7N7K10FPUEByMjIoQXubQ8xCSPe8hxaZxDFG
IT0RIh+TIAZ0OvKQpvuf2lQr9IIIbn+ln3WJrRgtYtrJvs2DUieu2ExWjw9UXQIl
Q1QTdIPyorcGhh1z1OkoQT0xstxm42AzBGnqDqsg4RJMuL+dxt3dM6Z3ht9jGKZ5
dIEoZPLkvUnzYMH6bBlqtplti1Ne+0PlQ6vk3D556/HVTkJWSeHgCWccTi8/ChFQ
WH4rjHD+nH7lqzziqDN1zmfsyM10lX1mH7Z0cFBofxQjhbRiWJ+dk+HZ2EUlmJE8
kYfKejLCiMfZRuY6Ej8m6ApRqoaFzoSDcNGmxK+DEVHMtAq4PMss8YfAemnS8eZh
KhiEp0QbPWoK9dNqcifj0RlOq66QEfTpgw3cYEkbU7h5MDd8/acc45/9bvWLKUeL
irSwQ9U50AdV224VeY0sIyeljO4qgtZhyRaCSHnKF8X4bWag9VuGIohtr5oHqnNR
Qb4YrDhWzAwU9lfNC31qKRhBC8UGwPGuigSqPVr+KdLJ08Ij2xV3VwFkK/KrSmMo
c02A7YOxKx/gQyPHUHmopAsPWvq6uE9BCHS8bhLNPPUQoVH/EPeVlEgOX1SNrvJ1
DKEa1wUDN4cau4z7Y5sOATqJpWKJmiBa5kvPpeci7qiHF2gIlHLXJV/bLn3tSzRT
2KTADS80mgdpPWxjxySCSZVapnF/JdiXL2zU4LU8xJ+Ux1d4+PZBVVj4tYdszwhO
8ev7PRq7Al8HTsJVb/TD0HtIR7QKlBX8AcKabb+7f9M8XtivG2fIseKXv7KoaZLj
B/bnXP6lFLGj7VhaIaYiXZH9UDaK70kOZDXtP8NK+OSaXF6gvURara5yMqlpuVwa
TJDeT6XdGd2xgJO/dsOSv4SULtUydWPe4DEHv/VoVjj16D7hjqMQRWTUTmtRZK5j
RsKGj8XkcrsG7OZ/0DjCtV/lvPVShondTdZAxSsXSvkk0IYTk9Zf0TFsjX3YjlQ4
FA5Z1Vn6s0PbsBQoI2+ruR32RTDLjkdobQc+W7J5ccZ0O7PPdeL/t7PUZUnKRYcg
O6Yc9nMw4gm6MUojGyzLkvnpA/p68W2Vmp1uyipTcb0cQgY8HmZyG6ZbedXalicO
lMSlpW6CL6RF52zicCC536YbYb5nZJrYjNtmRZTC2e05YBkZbxRpoh++v3ojIWMn
AyakitGIN4Fvjr1JHh8hAgLzjQIeCv9854KAzMHCze/Zz6tKS8zMxto+RgNYiX4R
8XswgdY2nmeVk/fqv6aG2W6S04EoeKCol6CDOdPBrY8QLpkJWSpmhEgwa7m7879q
2SRT0UJYN5UxDXzwLNF8hrpAKNvXHzO/jO4Lm4B+p/6SGQ8/ZOdus1m9kH7yDFG7
RMeSAmZitzcSsuwC2jY6PmLAEptX+2S8YWKaCtngV6ooT7WWzvnQ8U91+GjlGXsQ
7iPDNZHo+MZeGRIVsF7wgfp3CE8twct/jWWsASlsahIjLY4U9jz8teDLLwT9++OF
3NxyzjSniHcXa9jjwKhp1mbxlDRP1lI1aEu6JQw7E/ZKoojAbbksn9MXYoyrm1L2
UVoa6lsLF/ksf3Of7Xll5tQIQhyXqeHnunQAZ8I1hsnJELBKFKEK8ST/fIoNkxn1
7lNsg269i/iVgTLgJRow7EV46AMTSvvo+NFvmHY2GoFT95Gd0OHe9D+GrdUYOU0n
jgbvOJmeIo1AeGG0OlNAA1GVKF0N+P+zs9960OrWlQySfjgp0kZYCJNZq/2wd4Az
W4NH6pVU8SADqV2Z7lXy73Q/wILHyBoh8go9IqBq5qbGqLIFEK+zElxjBAeROcMT
u1R9bvxpk/w2VZdjQCH4U5s5B3L2hdlpegwWXKVgNpExjJYbLcXjjDS4HcX/irfp
HUmpeYdetf5+TuQysJG+DMPgqIXk/yB8VWxEljvi+bQaM3MVON3IpK/Gc57NZ4F+
RJ9L4QgLPBo9v3suzynRBtqr/a6cB/dJzulxFDu/BRQabC90hBg0kQYzirTUVQ1A
GBUThrw4tfUcAx9Dsk4puT8vzPa0rNCQnFfTckWcU7aKJZDvhSvsNyGCCj2dfLDW
D7+6HcmRW52boOkSM3uCglyyxtejqGErTF+lACcScFbPwDqevnc7oQsIvGb9igyb
F1z3Spfml3OaBcclpqdwSWSgUVI36nv7CvT/D33aCDWHS/xqzfOb4uGgPtrD65B1
yED7Cm2nev8ikjNFhIx5/7BiKtPr755NhPfW416TQoSJk8DEhpplNVJMSP1bbzf4
3rOhI0bFeLs4OSNLCKQfF4ethXfmBiszojYiYTTlKLYfZxCFf5pQnazTGn+2BITZ
ETb2shFj7ganijj9ggbVOEFpDeYexqZ9+5e8AdIXYYg/TGUZd3M/2oFIzAK9D2ZE
qkldA6K59hQ1V/a2eQXfVWL/0Xu2ykq2fM5i77KmKxpC0bdEsDBTDdX/KiMP7kpd
7f9DibCb8h5J8HJOZKdESa8Nxd5QllLlKL2dMIxVeBhOzhm/R4xSHE0EeCUe/29f
gEV3dw0+T49vRmraA+L02an/kzaXJkm5r8ixXokXJL1bLErsFTOrL/J+DZmc4HoO
RaJojF4vMJSMVoZMQ0F+ZLi01xTuHfPmXlPQ6ZgfPWIJdv2F0ZBTmwCwtGMVW4hP
s31bk3cPR6gXOhqJikPh+d2wjL4ZZEB4Yl9IObffyAveKck3kgRNHs6OZlyMoKjo
PQvTnjd9JRMZb6cGI+8KtR/kaoeaOMavE2znhNjq4jBja8CfQpwZ/Aprb44Mbyui
iNdTp3ahfvSzAIleitm42mHIOyXS1TIJg0uQyT0lIhn/mcySH+WJBFqON7HnZVro
yYp0MhwjzB2KPSxSeY+C7UkehzG0fn3IXEoLtT2ILb6ygTQgVU/eISN1P9FteQaH
Ev/9NMWjF0EqaGlomGwdywFWLX28RJRXV0XS1qibrlNh6pUh0Is3fZCtsRpAyjEZ
5jSm7I4612yTxPfNGvfmpb4tJ3qvxNbG2ACZLHiNXIRBVHl8GaPyhuX57G3j7Vyl
X1lcdsk200O1FOrpI5h7fpq+4mEg6Ct5fkZhsXa2LaVwyB5X9Dksugxfjoo867f4
6oluI3wqsSXXyGvznKI/0zn7USv/jg6ic5EjgqxmR210h++pWfNVaxtIwQ0P8ctk
RujrKZ7iKmFVCUS8HNLO6201ebbE+1Tc4ubV/rl2Igk2q+NnZd7oQnPe4N7iV5wa
T1JlyfvQRwTZXaSoGJ3Ft8CF7paJJvzi2l62l2y2xAKcvX31zSurE3B2v1tl7/Gs
k8CVFwmfoXeHCTccr321Faq+2rdzj+W7BkLVroR3D7UwGAFSss19JSE6D/DiX3t1
y09BV8gpISzXcAwge0VWzKmCH6P8iHGHanUo6FeesoOUx89Znx+cpspK/fS4R3zB
mm8MkisocvJ95xAJfwlUbP4JEFnZobrdLUjqdBejuPtT4Yav8t0xQbsaFe3fPyKl
qiSFCyX/QdnJ+sUlSpKgCw+7jWGT44XNnoN0SBMI3v4IS3M7cttHftbAJ44sis84
7yuelRxGtzN3XXpCZI2uTeqi6KsenAV/o3PjNTFlGfg/XdtRr+yaMPpiN/+d4zHl
XQ8SAs6AkaPgXkpf0BXYyGSO3/ALg2PgRugiE4HUO9vUGQzufW42WbwgC3xvx36f
EwCK2W5fbqGH02XOfwduNaT84UQvvAQ2MBaoorFi+tQjb6nMMSg15MhLOzve/FIb
M+ZwY6g1D/4EfbiDnAsZCRvFvZ8g6Xp2IrHTVW5gA3zZ1TdBtkCgpzntBnyxBkPJ
pxKBzCFGOZ6njuqDtDR7DEFM7SxmqSwYMAO6yj5WHm+qh5ffpMo6RU1rZ2eESrkn
pbX4wFrmhbd9DUAd0Lb+QGSTKkQL6M243dc763ERGjkJev5YD9PjazoYOC96WTrM
XrpcACE9AyhYsBI18Dtm+Fk7qToOW8TnEwdqxnPixt2shMpIbHm67LDrv7/HBNgV
99Aa9cL05j5QjGaRVx9ohN1hnTyK1s+v7T3ljAEduM1fBZh2QKv5a8ToUAxKPtQG
ewmzHJEBtKlfMJC6WYXKaP6/GcgR+nxcrNkhfP+j4PsthsLR2HYR/HtRljqqTA+7
s3wygtslAk1Y9DbqjaBVTzlu47RGMQ7qxOh/EtJfynloF/l/EjvwNpa41ciMHsyO
XLAYntVHs/eCc8CRnO1D0mFsUgA8PnSO/TRe6zrHtgrUloUwSRkJM1KEGl3p/Fvu
Bla4Lmrg29Fj7dcpZsnwf9cDnS/iKOEMfMIsHI7fX2Le1z7dw/n0wQeob2+0uAlQ
V/8UcvF0A4i63j/4t9WNCEeLehHF/xsjVUDrMR91Z6as8byIEtW8WexMZFLSSzRj
sQdw21mTBCUbPr0YrYwPzhpFLnwMVK0D7fMebqKXP2rb1MpnMzRSBDmQp0PW0dyx
P5ImJl7GGxHB3rCx12z0B6lR1tP0JeJfQknlS/4VB1yFud0BJhrMH8u8eS7x0SJM
veD0JBpu9ipsjvJN4b/p5NUV48pEC0n4abrglhZ/ZaodKA20KYdR1jfpaqLgg/vA
9btsoHlUaqAB306AdoTeJ2QIR22QrWkEDoXU+Ewq+xubyAA3Az4o2fsdnVbnDNmx
yT44b8Q3TPS6922ZJw/dueF+cbAMrnkdVqJ28stCPplASEbQ9KZkG0MbMEpb2xd+
I8BnrLBjf2rXPlDohF9evsrOzm+nZ0dQGewsX7BqobFsa838JkH6ZIXven/tbXAI
+180zHiFOUvLlYtS5KuAe79vN5JInADjZ8+/FXSVtt3BMfFjYob4qTiF+F4Izfck
mIHBbJlYfgETMhs7Q/9W2lr5fQrMQlG0lQczz0DZBybvKKyYHwn74rC9S/7z+uLf
pu9Rdx7drf915dgNoI2aKahqzk4LfdU+rDqmiS0wzNkfHyKhHnUMUmtOfQXWDrxB
vr1bSm1BZDrqJpf20Zm5o58/jvnBzTwGVnF6TkwU9Oqb8ClddGeYnOprYkKbMh+X
ynr/Pfn+Cy850nZTWRpEMecQxL6kOU0QrPTv8/FNuXaa9NezevzRXdLCEiUeIZ9L
0VXGZY3IcD0fvsAIQaZgZke7nCTggJVBuhgRaqyC+tFURQNfH4oo4FzlK3BDkB85
7cpxeI/bbEg0N4ZcMJqccUv4jxIDffqpREIQO6T9cOBtznh7yQZPtxRUSIa14A0J
u+htk/7VpD2q+sFaKyXRfTrG5EGAUcBgatlUDeEI1i/kgS/SnBz6YciNsYAqho7R
BZyxubqQymeFDyhjdsIMeXI0Z7AkxK//Sm2WxQ6llxydpX0owsXguQQdJH/YMtTR
HIhXbFJUhj6Oft9yRX/VOMsPjtM9x1cWK0X4XRpkuCbGtXWwUpc02odFOZ5nRmC9
TvSZHjQGIZS53sRPhPjFJjM9lS/2g7VHPwrydhBdco8jQ1ughkIFxq0OKJ8QvNby
Z65ZjQq1T5pvgWE+HQOmQbxH4kKSbGRgjo2dfoOIGfr0W1uXk9isMgExXnbP3kOf
zeNw8plp4XyEvROouhS7x8pkWF2opVm8FudCdXOpnQxprt4Mmr1SwugwmRqLGs0Z
gRC3+14rf9rDVfVvUHT4Nc5sNPaE/L1NSaP6ARxA12JcnciAOFbp+djnmDhr0j5z
WAPjXNIAg0MKxcX1SEKKZLPHcezN37dWM6TeacBMc8fwA9ssZZaJAr5fgFJMRiFE
kJSogcd8Wu2u8t3wP8Y3PaqOP4Uziq0pLW+2AWtkygrtfk29QugNVHpbWlOH1nwd
E/vC88qn0nPrDq0JYVJ/kG5rdY/tFYBCGISXOdy7eTwaIyql0CZQvGaYAz2sxOB4
hmhkr0RNyR7vXSHMvQIcyZTjBWzWvzHXEef+WZ30DiLUOm1wmIX0bFFgdPXoOuKX
mqZSWNxDtf1Ey1oOBKZJrhmUyP3xMM0IB/58NXr6oQG7QIgmQUdL4XqVkvVGSJ2V
K/sXvxAGLGm48wN3BljX4ac8d59ae4/5rDcc2SGJnlNR3Nz7gry77FaSJp/F/JQc
6882OemPfmjksjxpaNwyfH7olQThd1gHRRQWA/RepZf+T/6T4ie9xh++Vj3FgCzH
IO6EKk7LZuPROmKpeL1kdgUV7x09E8j5MBYTS/fZUVUvblbfI45h77etLQiEbtAY
sMcUXfwLC6uhAruqZc2FNLOCGlnKT6JDSTFVvZddZima9045hIJZGLPM78fbkVOc
zqn0N0nPqQGBKgrVwGf9iJOWRL1z4OTtM4ToQzrK+ELjd5rSnsnXa8pCiH7ixHgE
r7DTNHQLwsxDnrL3nKPTQFpAkRm0YSH130CTTXw0Lmw2j9sH9jve5LEFiF0hro0a
fmjgu6joDkvttp2IE9SuFMgJqit8RJZIe0vKpFZX6fL9TufOTERe4BorZsYKgERD
BbSdN1clKu5DT0ffHnQLrofg9hUd9AQ6mztcWct+kwdvShM9WwPpuJ9bQ97HI6Vd
OGwm1UbYjcyt/OxRD9E97mHcE/vBg14SvjE6cCXgN0RGwwI3B9fWuzvTgiwGiR9H
ApxMoWRGAmo2xHCD+Ri4SwsUncGdfAzygnIf3GR9nL4QzwfFqV2HLcFm10sReNwY
NsHxDYzCtU18YSuI/7a1OjKBz6IaLEeyXGPejmJdJSEEIMHXIjOlozkdGMGtfZym
IIX0raHuQFSDOn0QsnvNT2OXJMjBPh46hk/eCRBBzm6E1tccc66K8BtRIoETjTEx
PlwmqMHQJb8miejJ6lpxZBhPlcl0E00NGmc+TkQ8DUSjKL3oAUvoalDJIXzULYGW
vDVS9gM/cj6IZBLaztfCgqLMfG6MLtsWOh1uQkbNSvhHbtY03F9+4/do14pTDkoO
Rb0Dnp9F7AFPhTDvVZXzDgsY5K/R7dgwKZMhcBBKmWmcJHot3K3n8tlTf98ZIUfW
8WjupthYOTK8iWd/HkEH4rMNGH9IxWiER5IedlU6OSZJnJaHchZRmRuWUKLAz1cK
sKa9q4eyBV7am6aOx5DXozYI77ZZoVci1RpBNVrd/Ltxp1Y+Nxd8uaWh3PxYBC3j
sv3sFAK5qz/aOk5WGEI7DWUDkgtZs13aoS3lJf//oZ50rDx7RQ31JPZsxN1671Ik
KVeRZ/68VIxMdl/Bdc7R1F3uSSUWRW0ONjeDC/xoubo5epQ2SM4Xli7+02/KITCn
4os49GOQ8qAD0dJUBLFeHRAfI+kdBSHFLn76TA4bhaMF9U9Rbzkd6lqM29H+uvUQ
+Np+yvaCAhp4YjlfwBZE/6/73IOtIKfuxrHNa8bKFzWtinRQRbct9cFRgpYat1dP
O7hga+fc4Gs9ZexWfsUHJSVWR6JEvBp9Mm68Ff+56mP4k96GjO62c82MFfFqJEZh
7hYhwXj5KZzVr4w0//n7xD1Yybr31OTquO6RypZ0jR4h9Nu0miagZ0dcXmBuOvrM
pm39lcUBBpeCXnGKplYOMKaDBiXFrNZqi8+NAfrnqsWIGHX4lMDVUMOL0kURSIty
YWo1kI7Ik9qr+R8Ku8GwjuY+hG7axu0GH/eqeT7bu64cDivJN5Nb1030/COwI2MF
9d4iZEDN+JZWl3GGTsDlZJs7GokN4vyuo2YzHb8IQYPRpVS7fOe73ptWB2/cKRn7
56AhO31QI32wcgPL7OOf1oo8mbsbUnKjx7pcDw0a86Y5pPdYI35GycSE8D1xfJxi
HjuF3UO8j1/EKwStjFeyhamhga4ZirB/vRC6hjMGWmWQFhMlFv+RtJhwiAp7rxFH
WS2li0yWQIYZ5CvKLH+5TzixO/VDOAzYhpWmyxcicUQtd9Q8g0d7h/4BiXdjerM8
OLeUBj/zJGWfjQ5ZBqPctZlKnY1xO7RhOIkYtGN9nZMau9Gj4A+Re9QlAlrSl3WE
xmp2MhpjS4PungBDr4+mKz+7ZIyYuEeMTJ5ULnJuojrSZXw3qCjs7CI/lm13OW0i
F0CJ6g8NAYA7LfTs4hbnXk9z+mVEG1b299KfMqzeyN3lGknhzGlUHuu1zYWcagDm
14FStXhcKyr/7suQhfzS7gQSPH1YsxrDWy7DcCrpCGB6Z2K/XaaiMePnAbjNVoS4
VFreG/dF/L+P2BlSqwzo6ArIakK7+/Cz4wxh3022VhFKC9iAT0eo6GW+7tQ9bO0A
9RXMW5wAvZ8ird98Jc3oWcoIxNVsIFlxSFD0cWmw1EZ9OlVacCC1+KGpZNmNBQdl
EJ4so0uvZ9iSIkvzYea4z5XlHoTVVl5nuFZ84dbDlIWUpTLtXxsmJgfzaJl5ao/A
JaUaGg7+5yHiRpnsVyg0d00L3ZRUKHKM8CceFMzHiLX3OyoeDluLV+8BApAWPzdx
mHPeFYDlGMGTdE3grNc2HszB+PEs1lX9OcYQRVJwyc1szvbBF7cM0Mkn+mdy4A7V
HDFttRZDZifTqAof961hXUHSGAPxA1uG1WpAgvw5I0S4dlgfKziMHMtotrv33ZOy
Z7wpLryCR/Sfc0kH+iRrH89N3q0bDkraPLFGPg2rcknuUJARMmueTpDI24I9Przu
wGO2/3XconYjQSR5aC6DeibgLTboyefYp7JLZdelHmJ11dR9FuExuiRH4ZojbZS3
SCkiN9YsWAMcgwNp7d1PyVO2ZZ2/wpui62TNd85sr5zOKt2+OV0onC0VglHhhNp8
5boZMJKiXosch5e3IW6DuRslAQ68h+IAtLWBnQwqiNYjqM0SbsUMq5UIN6/0WY0x
DY/5B8zd15wEe/RTICktvQMHH61bSXI8YfAFK9maYuqNDOquSZpJgZ1w2zG4wCLt
O8p298qY0p/rcKATB9HgTE8lQCD5ll8YGlxij05TAJuU9n8tQbgNq1o28f/Fghu4
nQCaomTGFmqk7zPvzxuWc6vLD6d8PP3DtkmH+VsVRIQVfpq2bbkcLz29ry7r/dbU
Qp7datYIJrS2Mbz7Lbh+ZqH99eSU87mNT553qig1iXOVgN8T56M3UKRvyVM2Fsz5
cyj+kmEr2O9f0Ocxj+8meq6lBRK+mUuFtRvf6LimenJrgKXX4bStC0rzTdgPu3Ji
9RwIFWtSDPqzUwX0Xc6KzKcEjPV/hu1p61mHgkpXEyN4PBNkNB+4mgKfxFMnLHbW
nC01blyTOyNXYOX+Fuqmj9B6BS+AamvMTDIiVNZMAMLIgIlwCBSkP9uOrEIHE50Z
Zhp6byUn6X4JE8ZFDtI/G6GMCCiKVf+2y8Vi4d6fMjhfegDvvOOHgqnXAnxhPrVW
59fGiCaENnwtleUqFHDnNgD8oOtIXSCd1ANLoEK+VGeKNNYQxipcCDNuxkxmmRJ/
yiINmp+cESf0HHAy2z7+mxmC5AITUSHsj+tiHJA6xZZu0jJEVEs6usD8ln6T6QeM
Dk7hurLDpWSJonsMbOc+SH+N+iYpcNWGESOsmdo97gE2W0yLdeyLHjk0gq7I9jKR
HqPx3hXF7UBR3fkt9QLR1waZhqOyh4ORG6cUCMq7c66Tsh8I9jgzICEo0vt8PvfI
oglFhrFXhxbYFFQIRSvCGF/HD14fGjibX4EMK0UgeXGGUGxCJbxYFDNSSXqasECQ
r+ZobhX5BpaDDUbIwyJRYKrh/upC83Y5nxSCbbkYxlCp7aZPvsM8rPbFCU3Rsx5m
26pG3R+UyJLqt+SGko1L8dj/NqqTBXIjivOgF9nv1bZw356xYANvYWY1AUXZ6MpJ
JYWH2GxwHjgyTdZ5EJCswgvDBp3RudYwhsgx6hU35XzJDkRFQDPCV3C0Bqm2u+v8
m38HXKUBhdPNMd7GVUBInVhGS4R2n+8/MgftTkFQGdNVcecZ5vVF0q8Cu1qyFVeQ
63Av85JwW7cURvvKQieQGLma9F/yAYEHObrY+lu8Fatht1/MfxQ8XLlQwxIFLx+w
isuw6mkNVUAensqKt80sGmOJdn4+icAa6fXCsS6sUlUqlMLU8eiEhOxujZl8Bmc7
6cUdREhKr7JPGuY9q77Qz2GEHFQT4jxcWRRkwj30u1kJL89vn9kiXAa/s06WtATV
2ezD8eJiaIz1E5jeuZQBUc5uDfKi7c4F2CPtZWjRXiUQCqGNtFBSoLFTn/ogoZGy
PEUkYyj3njusHDgwnT5ZDLsu6X7KicXk+vYAyzuXbdJcljp2UsXiqF8Cem3cPgHy
5zOmu+zlJHYK9PeeVSnqJd0eAXYE42gnXGpDD6CTL/T1gytl7Y7I2twNzeUuDK2z
d5RhXcOGxjbhKMi4wECqvFfVzCtrpHhteRlKMVV/QcoqHnO2ZeFXT6IJasMpD20M
ujIbV3vn6Vq7j96wKa9ny1oXeMEKbYIXnYbNqvam3u+KyOayd3cIhcfTOv643rr1
3VEnNjNVQUVwuQB3JDBvHBXWc4RucyR0w5oKztPu9PcQyMf9FPOIUH6yOTxoNW9v
Q/lKif71yn/8aQ1cCc4vmSgxI7ODpyc7Jiow1QG0B3zlXuy/lGL6oXEI4CkY5zTt
7r2YngXkKGKROa1BbwjNdDq2PaD8CUaknvK3Fj/a6UNy13dJVVXAC/oi7iYQDJlr
Sn57piG3EbAMZDMprW+H7kG0b3iC7gQISQSe+rSCXOdkG+yO1+WAh50eonbSrYhA
jNC9CJEmw86IpdZGLeFh8im+t+McswTwuiFzKBXifMhhwnGOf2jHZMjuxR4WC558
nnOaY8nByKl4bzaoKrAAZXgYTfH0Itc9C0bjxEfqPCcPGEN1qbDSAy1wh9o6M+Wa
7bNQCcw9r/bm/m+RiBxrDqqclQ0AaTsrKgONHf6WWR8Cd++jt/ELqJ+1JIxyOzeY
vS90deqnDaq33B88+wVdrOOZCbBRtMOxLuapfMY42vi9m3PTtYHZtayoa0t1RnYo
miEk+LDDwlcNDhvM1IaltSo/QjSwnBaF/4FyDbI3/4F0ppJPKMpaqUxmCntOT/I7
YCHPtjFV/8y1kc779YD7mNeF1t7NBZ/k8CqxIAa0brWk3p4YBAc4pwSQLOd6cDNm
AVd3st0GWjFiMbQvlNV21ThBzRW00cWsqZfPAePGKz7nO6wVBYRb8PAEX9eeSbNN
/eHAOjxyKCViR+fnbFKqWTpbIglyJnGfqMTu/zqywI7DGGX/7hcMl6ceETuXMAwL
T8tkeg4gaKsWjSa0bLaSi+8UpVfXHNKZy5u6Sg29AvyjTRTeJAmBpP2WuC6VUSuj
mc2gf3QioUf9YjsfRkF/47hL5fLXlJKEtxvs8DvZOShRKU1DZ2CdQo2dFeZD8x0/
9oZoymzY/nnrRfHcQLmNqnaq/9uAjGATAPmNAEuMdFL92NhNYZng7vrOJVQKhuf+
he6w3Hrqrf+RXtseH1q1YQ59Yse9ITuLxg7kkcbGpXK5p/NPTM1qCF/iPTRZxdWr
AvYY/rnJInU9vWyV90Mt9Itfw0UHOIy+Kq69ylVzqlziTbH/HpNxECYqV9QkpxrJ
wl5ioVMnyy8P4w4kFAQ4+gVEOaz0GoLmqjY8M8s801xOwGa3fDXxN8fywy3sVnlD
23X80YEKv8dQvR9Okp+BDXHOLSTin7Bjo6E0kJ/6EF/IFcFbkhgQDYY67o02MT8k
oQMvDjE5MV0abm0IAyE365+mYd4TN5a+eqsUqlW1dAkadwrVwtXq+r6A183Wsehg
T1FS3I9gbYhJlePyTdTGrh0eVwBq+8VKc+N0Vq3Zr/mHY4N943SaEe1+oybK70gq
6lU7n3U9sQ+LK5ETPeuH0DfBTR0AzODAlMs6HLo08XVHshMC/jjZm+4SUSAt3bTt
sowtdsjrskLiLSmjJfFO2jH44kDKsOK3we9D6hW+Qu3Gd+hOOgUEAFSw+oJtUxFE
pmUzSkYFq+FyB6avhsOvBGLIoh7k8Je+4zio1DAMNYicj1n9iKvr+pvx0UUaRblw
PrOidXhdx+CBqFbQ48UmqVuBkNqUYfho3PUrYjlj7FFNaiFpsvK8HMVfCRuERskP
3EKZWOxqb5XoaYnlFJBFxklRyRrsQF5U2T4K+gPqN+K1hDKQNzozUTLM8l2tKgNv
e44nCQVva55OdgY60urmq7a9pEtVsuew6/Ny3GHI6eUyQaM9utRpgvXkactM40G7
FxtRXcZFCVwbfpT77naLxsgirbxMB3P9QnTDTqMA3+hUOyy3ihQaD7wbj2Rcx7Rv
Pa2X1NK+Y1BvBagpuWzXr5j0nojEeKHWHbTYTCLIQLYJ3T6rA5o1PCOWKThpwOrr
66AnimV8zZCDSrMoHbtVElv1mGFItY7AH2O937wP9mvi6/hAVaqcjv6F37YR0gMO
d9WtRbOlUEHDbXxQO21o5+M1DmXt2JYLr1JgmNr8B9JTac8PPs7yZ3tTBkU8A1Zk
SV2p/Xg1ZK/DcglN6JeSPb/NX1gypGi4MlN1WVu1u+Qhvi7/Nmqk2pnlVi7gHe7e
qNm0wY51zCs4u5FJ4CHqp8yAPOeTY/+tKjdoyXqwDMTGxMHYco7CUD0f695yJVkU
mEceDt5utXUrgq5bQFTkvwL1SpZ1AyQpOJzu4k19yRlXprek/0DgyFXKXVgry8LA
ttWvhXsz0WX2Otgjq0/7fTbVbM4i2+upRCeV0BE5ZGpTDoJWaFKkA8rmqDzwRDsL
Iqt3Shs2kts651+dwQW8UyfjIAroxGdgHsUsAMIJNqiocSX0ZCcIos8LZIxt934R
qSd/M3RmsGU39T/uamtoIDGTORC+hv51oVCycNMuO6qKP0gb0kqr2y0ZmO9TS+vB
tTL5S53kpbcRg2Bqe2adbPvG67fx2abKnjcabVi5XSzH4ge4ByczWgKaOH7qMtmD
N69d6Lm6DPtMHq7X89b3AShM0ldvZ+Zx+kxgCwdmcDhtL/bHZJFUshN6yv7eseOp
NVHB9XdqNTAODKgMQnn1ipQELh2X7uKicCZ0L/CyKAWtgcR0HMqB4z6LDb1lqitg
6kG3YEVlghRi1goW6zZ+K57/mQ03jaO5hK4o+T62WJf9JSDQOiSY0u+Shx51gJMi
VKctd2CFylw5cdgtj+sHXE81QJ15gSRN84dySlQ87ODdw/2gMC3q0YtHCV55sYch
YnVqvZdvwdfKxh/5x05cuU3JD/EDYazGWF77u6P6tY3RTjYOnY3XrxTq3oQvWrBm
d4w1zlV7CRCTyL49P4d12iuALgzm/sVEJK/kUWENPPn/IlPWFWvnmfJXR4Z8Wmz3
gy41LRp3fGWKyeg8lTRk/fWagcxGTaTEta6xtDDkJbnhqbOzjF+01FV9jpDBAf/D
ysoKzaEkycpq+nK02IXbzqqs8DDO9cbiC7QuoqWSLtx3CF2wxyZvTmTd068B3L9Y
6YKU64kBsd0lD9fBebvTWOxAxvsq5e30rN6NnV2yP4B9nZXS4W90de7bZL7kyNUb
m15PrOWcrRJxrdwndcQwgNmPF573YmOP3hk0HqjOErFM0aYMgim+GkmpGPZglOtb
lXYsvJggBFvKXWZEl8c2el8SLbXxcDqahMl3Spo0yLADzyg9uEa9Mvt1/rJdNTJw
yLgc2qUeybzqnubisu0fCO6WD0wAjyIOB+V1Eqb5lFn6tm7+zhWBYJYqMVibeegQ
8AqJSG3odGL3MW2lI6A2UbjEO2lVUlSBI7Y0AX0u0wtzdj7NXFfPksk+lkFCAffT
9mzVK3IV1Q1iXFhFm0vXf8bI0D0U8m6VKwX6V0zsGp550x/PRPZM14MT7JSCPmIt
4NdW08rXiepXU+DINzYko5FFWO8cK1dDh+O0nefOCcEqZtsCEmu+wt3FeFZzJvQ0
w+l6t3ZFSES028gtyoTPo4qtrLiTfwlLawlpVdDH8RVY/IRET43DrE3qEYJ04A5H
tv9Rn1RaB5kfDXUdAfMVIyE5sbJNXc/xjZEdAFlyFYa7yeBoFpX5J6ovPxQQAdE9
CymkG5MueDP9+gaWxBQWzMD9kPR3sKCU4oFxvPPouuQFRBYKCKSO0dA6w0jqzdUI
8ylqq78e6dso475kq2DyGQrbNq1nTFANBfK+ZwsL4w37nCIuW6OU6Lb8u1YSK/le
8oCWtq8qmH6X97lJ5QwiY45/98LNhv9zKFLyhxZXlp/7qzvXiZL/LufcbvL4+GP9
4Qb2qi4AunmYF+Isdldpm3K7UHaND7CDfoR6vYd4rFD36AKMGOPO6tyZGONlp5Ms
KVMUVCuRRNmE6Z2wpnQQSQ5/yFq6jKLRDwMaihLWcJucxvvRoMSjoOaMCvx3Z965
SneqFjLirX8WNPHJieq3BMi6xvuk7EeRpWP+YxKd3yC799sP2/jQLL80oELWYUoQ
40uozP3hPmZ5LtOYxd5aMG83vCY9J4nhoV+Vx9E899TpATMyVszCy3+1oWNDubf9
lD1xLK+9063x7ci4dsEo4dFSaQDC/PWOwjdLg2jPsoazmaLQ4fDdLxjbpMsdPvyI
l83fEF3Rbyz3Lz0Mxz/El5glXN+7XI2A0PpOGy2NEbin8acM4jEtLeXfFpGGTHZ2
vAGaj1xCSNzHoXXwMyGfWJq1raQBqULiQepZo1UCwP67PkhY8b05Mr3M4A52VcU1
dF/FdFc4axl37qrJ3IkamseqDagbs+DidtqOPEJl5TED0TVmQdzV4Zvwqfpgt1y0
QcE7EuduI77mP78C8IXq24uI1s0thBVh9RzaOU5OU43Goq4noRShdPwX/nVkCEjh
nRRHTdZQPF/3hce5J3/FJFwGEuwHFCspDWaRO12UM632YB+2NOAIOpnJOsEP/iuV
AE+DTxvBbUjevRs58DSN7TKH8k+9yvI3OFFXPXuTKLQ6DU+1pYJLx7iv36FJb74k
b9vSTnY0MJ6eaiLEO9WQyx3h8Oa/rc5HN8TVuMmOKxVkwNX8IujiYVwDSsawlJhN
lTYoC7z266wxok+Sn/j79/FESVhYA1mb/1N9lt9SoaCKCKVy/pC2I59lMdJgIkyi
puBIzcbCmSCf5FqGUwra7a+A/LhQl2RWmmm0+TZa6stMHPWicMAWmj1me0v/+ObA
Ga+aWrRJwZiT4uOUUm4wQ/2yDGZdiJLbmM+/3Isn0JVv/T9ZmEuyiUYS7osnz9Us
+DMDzUhS5yyZQtkqiZi1EMvYbgsPpfQzNod98t7mUV5Xe9kfYBReIX1z4bPOacmY
WjMsqDKPA9/zttKZMNOnW1oiF92lHTgzevf+QROYtGmdnDvL+TT2Dp69jisn6u25
gcb8hE8XWcwQ9iAHKZjVt+ZYmgAYfg0BnhzjTJMIgEQp5A3iBzEnQVlj8y7i1Nb9
1nSpY/KjIS3a8OtgceF0QTIkTxZNYEMFxfp80xA6Wiyg1GlYnLWjsE60uh0W9ANn
JQiWEeqd1DaD/Ypbma/OKy1mrRgoX9zbmuQP1kXgudg5mmkPNo3R6BzgwNOPIWTI
hwcqDhUQSH5ElGvIZgysGFsz4UqDOvOv+aMKBg9XTqiEckVIG63ySc29AErhciFC
kUgbLkLw+rLjF60QUwYrRbEYHfKkIZuytColxkUwEnPMSROgLWuvyR9xOaaJTxON
X7Gjrb7xJ/SEegUzaEfGUKzZlhjTVSqeqVQHKa/zkZjKjN/3N4VCh489FPmdK8ad
t/+RS6HSeaQCUj6IpfqyqDCI8mHDZN6qDQphI4BZkWKQXINDExCS0n6ms5mO5LGp
uL5pACQiBmBN7EU4JdyzwK+w9DWIfp8TdU6zoxzqIGE21qNJQn9W0F3D6XByjyO1
IyiD4AIz3htU+IpF3m4bpFqctJ8/3xY5RytDkH1c9hVb2iDrMNDLrvYDquYxk95A
YncQbD8lgpXIv3AwNJzfljCj8OVEw7XSxlm13FCHIv8kk3qjdr46GJZUJQSSsfNO
pVymcgzn8yWDkvxnv3b22vzX51pr8AD3PV6utm4qAVcjITvFjS14n0+vmoyzBZXv
edieaQY9sEJ2qFcgO3Okl2q9Jcgsvr+GHIKxDnglmBqE93ohGBd23lk2NjpClSNY
zp9O2xE04M19EkkFL46frF2Eg6xsRyE35sRpmgWo0ITaqAz4TGTsiSe4egGuy91w
euR4lxqtDxpVZHX7szrUWE5dcCyNhLSnE668jv1YM8XEHJphPz7Ju1pEHWKAv+Ve
VHwLjRIwr9CLE9AeV2GJ59oDa53nVFWmySMpujFVu+jX3ukHvGGAskFXAwuHcdN0
z3yh+1BECYM0vFxTKsjYX31B4kBMT5ueL8LjIyIgUhKpwIEMboeMkklmFh2LhL17
rtLy8YTKB6b5dZQ9VbqSfZ6yztVpre82O0kF/NSr8PZusQvmthTZNqIjv4BdQIbY
daO61p48kQRFOXMA/H5HAnrlnA8OkPo7VSF2tcCqDrSopmTdXmkFa+3WgnSVetn+
4HYH1lmgfD3iEIR1z2LnUL6a2V9X5IiXLFYTPkDZC1tuEzWcxCdLCLSR0SwYWOMz
bYEdXa4xuJc9h0xGdGdmPXWx2ncMLnWFRrAz09PNHOrjIcCgN5U9pw+resSAKCxR
FaYdRoWSvO2LfZbU5onrP19LuQMuyTr9qP1/tx3HD8SAsU3t2le8cW9X+BABqWIf
z/EPuQQBSIX2vC4VJzdV/8lSX1eWygb/q1Vm2tYRnUTCIfRz1U2IGjM18hGie3j9
UJ/9/6byXNd4D/Ku9cjRNPIefBU3ebg49Mke1p547krhyUjLMOIxHd2xSySmQmXb
t/eastxLaxNHZ8ZXY2MVpJf4JCtfYfLU7N3JA4xLcSCDoWgwz6vFLFFugYb77Hpm
OGgPKjv4yPggxLsItuyAmW6/wcXzlnC45qelZW2kmrb1CpAvFCEQ3vr3OlwfYlyw
n7bZnEUSV2aAdi8p5To4YFqUKfkaY+6gHnb26Dukx7zCbjmNii+sUWV7TDBrZ9NN
yan/xI0Tr0rB999S5i7TxGEunpRW6BDRe48tWVcwf1Tz+hZ6KPDWyKmWo4EgOpFM
9jH9FbKnYEO4FsQXDmOyc4NeOIBbkjeFpSWbcupOpAQ9549ppYsBnNMl+TPzq2tO
1zCqnjBh7vhmBmc4CL9rcbuqwZ1umBnNHUsWV2zXu4ID1dSQXiIUzeX7KpO9GzJd
k3djCb7BjxnMKTTuiEW2F25L9bdrTAq1TPk4XBc8zrBmVFRRisQNrc0FaNpfyKiN
vDpx6oj2GhMjJ1PbNUeXG1J+d1jD+WTaAS3+Cjv1iLSsrzNGzn84GnIIUo6sPtgM
pUR8f6flGgyQoG8YVBgWfLbo2Tuy2Kxblfl+97QlIfmInbQQxQ8DzHY92lcYpcCl
ILbzMnrJyA2e7H9Z4SM16fFRbsCTo7NFAeTnhaItTllh4RI04KROul3bLKFfkj8J
B9dwb0U0dqd2RQ+jFtQGxrTR4hXW9wyGFGekhc+GA7h1K9aWj/bsm3X+ZFT6xt6P
iCl736KY7hjlphs9ETw3Wfd1nU28NI8w7rdaCX2V4Bo3r+xpsJZuSZmfSKUczP/E
VDfwf5HCRDqCyNZR1ZeGwLsgelqK8C2aszONqDpM4Z/5AVbAty1kGeN9CKmh46nR
OzbCi+qtvM8mXgHBwZhaH5bmxUU75l33UImW1nfxd5/T85VRFaZ5ed+Ho/K1ia6Z
//7M6TjaREG4wR8VjCsMIpaW94SWnGxVuyYNjyMi1zWDduMUuoI3pTkTJRK00GMG
ikytwv+1aBvoN1MDseNQA8uNexF+XpZcWQuoLHY4QgcQqM0FQqUuKjy/0DzuHjfX
IKS8WJI+S4NGbB/PA4LNsq/FJrVBBHVslhqMUXTR+X0/7jYZ8yrmC+EfaJpzpGZS
eZWK4Uxl0IGA5AGpiBaNX6XSAVasDPxf6N7pTygrP2rdRwfAQdBRbwtisICG2dcq
Zqn19qxHiIxo0DOJfsRD03M14ydpxbLbdo8YP57X9c83FhDYV/8Livb4o3ZeFyxn
qjHmqJsQrr3JE6t0Ao2a1U4RfmmyamYmzHwyE11ojEfcH2VCXI1RwCNr8Ja/xE01
A8f6UQF/W7dSxh1Crq0vVSwj7Ls+42D2KyJ1jVaEFv0Qzn2KqIbDV2Wvy0DUV837
25P3cCQ+h2VhXr6+Gc1LQIDRScpJfiG42FY7dajxkq91BrTLrk/0JSLOB+ZrCR1H
0O/hIMrjlM6t2asXF8NnfHubIbK6lD7D8R1cbGq+azXPh8bWvzzdJrN2+x8O8InI
8q5X1SQD86fgGHgxBG1Y+RFydY8KO1h9Is+LJBvXAHkh+WGRyH+I7lRr+9LN/HnW
C4NKF//S63dVCK4m9WFyG4/RJ43WZLJpIRXVKArtSJKPEB0jh5eN3P1UagB2dzuj
mFbno3wW0pZQEhUlesIiBObhPc3eQhAAECYAKzcUvJtE5ZhmWkpx9j951ua3pxId
7QjNoxL15/yiZM77+QzcBvnb0ieY0EjujP4Bt5Ch/JsaPEzxw6d5ThBI8LAwwwEn
6mQA7i98aAzXoL7EOKbV/YQZdLroZ0d7eeXsAtK0CQRTjS17X9Kfjp0mBF4YS0x1
mNZQJTzxOdJZqaGzk4+obUy69wDF/9YiZAa01PAwQ+p6PSeJhYP3LHK670C9QXJU
VSKRMMmU+Cm5Be/qrKKZdixKPyZPRv8Lwxw/q3JFXuCJuX/S4XVSz1+UqTaoZCuV
60rLjpa9phgm9PoDTpnJKFZvLtI4hEClhQGsQLY38MxYmlLzezeLoagnwhkaxBIW
L6KTT8PihtOBcnLVJN+kvWbjLFbiE6NTzG0bLj9p4esXMfhm+cCM+4JaPwNDQnVH
OpklQpjm/9qswjzNzEg245YvpM09PeBe/e5Oj2F0sC5luNBTPbYD3S3fse2yXjOb
7YFPszxZtJjPTC5Iv2aKsJeNcETYvRF8VehKmmqc6eP67TF3e6DOaZEhuTiJtu9o
A2FeAT0Dgu1xY+Kev7WTucXkwKEI4Ric9s7Z1hy2xFiLogLzInWaYuOQ8IF9XSZu
30xcaVnbKKya9qM1ckSPGj/0pzedKxVFLN4dr571ezeicDGLe3B4KmFj1Z8BQSQh
kFxC8NQ1uecrQ4hnvT8babnLXZgib1oaN5leMSxzH9hK8GMZcI8SzUPlhv+tZ5FR
GtZ9WFaED2Ey9Cckw7cF024oi5QPYLh8DqSPPGhRp0zFqLU8yru+46P//XHNA0kH
Iffs2vWCoZ7pUfFJU6Yv2ZoeJk+FVi6Bl//h/jOPNFlOELjakJQ9Ync2tcFzJnxu
LUdLeamBO9qX2I+fsYktnnPMIW2EMyjzhPvmBJ3T57aior7RMusJD7BmmeqjB4a5
LpQrZ03sM+EIThbT1/Al1FZ1T+N8RVBKyD5HLXYu3csfKEiBnSYoD8QBqJswjj9D
X6u0W+yDaYS94klCMnP234666sw+t8+0rSQetEJkEpEc1jYSFwrMbWWzfDgaHImJ
sqpCvRlmY+q1KFq1F0iD3mG5DsHZprB5UA59AVyJ6JJYCHMsqe/r52l1Paqyd4sa
28mS1D/V4vmmIDOoi7JiIicwMk+HgNOE4vYk/3GGmpC62yuGjaHsDchiv4NFEOiZ
D3J1LH1yrIbawDIFgHEoIYVWDilrGvkttztpxQQE4uuWzuTaGzJ9f+a3xXEHd69h
aJGyk8sYCSiozHJ8YN9zGmxUBUkERBbMloywmhn7JLQQylUnxXU0gHH5CkF+yDbK
KGOQF30obzYzFcBOrZ7HapcUdbUpY+TjKS45Zexofw1aWV7ymDHdUmjZ/93eJmYZ
84gss8Qn2A0jGq+qtSstXDFKq9M9UZPxcz9KbJWrQAP+We3K27cjNhpPVROtshYv
zvuC6fDWyH8hSvzHImPUEKivgswCrO0WKXHUIUJtptjDewYMteyTsHxORxFEdVEd
8EL//bp/DqLkFH4Mo2zLaqm/OSkOVhO3iABNocOG9T3xGRpTmlyDp0G3Oo4EVQrH
l8Fxc/oRW4rtvfzQw3auioZlAXCI7fGUedoKvfN9XxYRu52f9hTf9gIXJ9jxHQ2B
nMLAueLs7xSP7W6/12qSjuq2lfJh5Zg68COZx6bW7bSw2aFeiHrFjlHixUeAlRrB
DwYpgHNmQNwV/7qNDJF1eiiBrEthi2+CAfgNKfL0xGv+oiac1DqGoDKqwpjTwvgr
m9AW/i5mZ0mGVOgIFmy4E8ENY+p9vY+CHunVCrhEctjJYV50irLp58U48VED6I9n
OXCjJ/RzpK3fRo64keZsAgbO31RcvLf6WZPWIiqK/z/Sc6WceZJf76dFV05DViMX
ndVz/uG+alYZgpAZ4uB6FACdgB6EBPseZpYmM2Qg6e8tK7rt94EyDCQemAYIJ9rK
W3wTqQIRZFRVu2jvNwmH+WjS3vw9aF+CdXMu6fxwUler9HaJY8QMhZzLyEf13iBO
18KOScvN2hv5z2xZCfsrqz/EcuD+lMcf7ntphNImtIVwyHoZxzcEd0+rZIMVjY4n
chGM7cdbDhv2rVitTQX2feKatdrYZaX1uMs1ipO+NubpqpaY56Fora6YQw1cHn6i
gFjQsx1Kc/R0hMrwP0D1D7AF79mLQJDU/M3XGExGsqwjDc8U4MHC8kokb9KMVtDf
ub+rixjjsjLBtPe6Yr8dcG202rQphbXIQFYswK0RM8DQU74gon8Yh6Ykkl6Cc1uj
EtGRaQkdGZI+tFAvV+L3rZN3bDgTpmlIC7abRvayQWRZ06F2xP+LaK6TFaBc5XgC
6U1fIMLpo4na0Rd5/hL0T8Qcynn2uI1q8gK+FkPHlSU3fPYnf1biQqDwkWd71w2v
77bPngcNkZWLxpLRXE4jwcqgLysLuA5cPfARMPPpwLLVY1uzdk7+NuSFGvr5N1Qy
aw+AlZNlmtdzBOIs7v3JEGoDaVSfEoBR5k6YMTMGy9o663FeeeHiChqDDWYPWFUj
tsl+pSF5xNx7KrvZYJY6HRN8c2ztxyCANZjuJhzgDmWpHIx3LHlQgoF5sjUky6uE
wP2wxVA1eRqv863/csxHDuhJ1tBzWfklFIAgmi4ub8hf1S2hmswYeexrRYdIMAPA
vu6MGHT7ECgj1110yKmOtZR0zE7ZElCP9MyyG3XDABJmM2OSlHre6VqCrCCsCwNc
j+wEVfOBZu1lkr+8ogolLcqx5hgmUe7BPrzcYWkdZXutFBG0eyNw2mWXo9NmXaSz
4brYU5h6SeOSdg7Hc7//y4qFF5qH/wIj+BhyEYXFdejCU1hEeR0JKsQFptSGK3NJ
Q7K5/5eWfENq/QXd6IzI0O5nmSv8ExqzG3cdjvldKlGRO93W69acNp6krJ0Dyp7V
JyqIulkRISc69x+KbPaOlEnc1FOtfRSVJZbDfBVRKitU+/0TgAMdiHn7zHHnnT62
eo3fRRnfvkr6JJdPLS5hnV/hCvPP38aKi9q67cL4eGC0BKxXID7r3ExwZTjbXR6J
6FyB1aOodnx4a798Glatu+dwrTCh58dxu21f4150MHpv94njeD81Jg/Qs7sRtBBI
pm2uT3T3Optci7QPTVjRFu51W87Bo+xovMxQueoKCQihQ84ImVSawfJJjC5TSB5P
DtAqiBsMaK0C+PEPw3J6yIpJPSjwW+BWiM2VtMSyvDDF4IsF2kD6fyBs4j/QVq9Z
gNnvSS3tiQSU6V8/QQH3I1ebu3JeXpfARXG4/yg6zcFjEPHFqi7rM0ZsFp+5OFMf
81iWiWNCHwosjNRwJwhZX1bUrujL+0xmhonAN1nobLTcC6vvXWIxflNoL5PYEZp3
neKtfn4mofmQIWcxJwkhBi6EUBjJdM+RROiZZHWl4O0a3jnmDBKHJU3Pk0TS6ya1
UJEF/IlpMk4er7372XId3uS53vGnpIOLrJfPVF8Fy2zq3hZd265sJLII7wi6L0+C
0VoMS7TCiXzE6BPhMNhbNN5dbtfWF+/qmHUgn+ejyQyAycNlVE+ZpNCIYvDR1gpV
u7F9vd6F23Docsfd3HL5bIurQC6FSI4/QZgvt8/bmQ9yoZwfnxE7MiRpI2SGQG8S
vqRHwAyZVI2PrZScl7HzouT5/59QeJZFlPEC96mNjDJViCilpB2Fcgrq4WGfAVJE
wpDrb3XJuIQWDxgJkgTpMRzec18o2WAP19uOLeKIyAyC2Hh+Ht4McosuuDG5sQp3
dj2LOnoqtg7IVRFppYYdrA1TINQKAIFCg8KDE95GEnwXAvMjwQSWKPy47Ha7H6cH
5pajatCl88l8hKpe35r6CgpqaC3FUSKkGGTCxV1EUPjYlLYkdduCFh3tPHLxHRHI
DCrw1sQ6cOmwFh/VSbfwTaJzqRGtGRAISZ5hOvDxeuuX6ShE6a7DaXtivsewDaFC
2BVE3KuV4zN8m8hZzkXPJA6Ouu0wrbC0uOGecxh4SvV3Jh0lj60kcXdT+Iot5xWn
9/rdREjWstECaUPG2c0zmk8LiNcEN0E0WVRv+SxjLs7Yk40Ux16mXN6QdR2fu5HD
ZhfaR7hmYLfibefQrFDotwLqugAnX4NAC+bGOOl+kCWUTWkAQjkDAFwMdGgB2l9F
RBqwXBIeSfYGRgBX2cv3G+M8vlriVNqIXUNoL9DJNB2p0giquZKGslRQ8/dMZHCR
j6A9iG8XqvaTIB1EzZdwm8GfyrRiSaNUKMczoKO5dez39UjNaLClNCF0BAS5FBJ0
VLR1sSPe0jHkFNPZwVX0r4PED/+wf6GOIjE4XmAwsL3h/wl+jCWzRgolr8jHG2H7
o4gAJKd0nCE/lJ1iisK1mCS/pTTO1PrMisMOQxQ0FG2Ri8f6Q67/1QT/NeXvCNuV
FN0s8VLh8OZZp2zTYiYFOmR6WPh3NXl4gziAxIcTb2YiXSD+6CAQXdw7TUIMRZzr
C/l6MQup/5GkEFxANBU0gOTEAu0HAf/AUdefcwTteqikv0vUMFVERxBgfVx5W8fs
Lxm1jc1jLVMfsOFPlM6MwVt5+TmZ0Db+WJFKpr/jWwQa43FVP9zhdZasAogh1hWn
sIpkdRMiN7ANoI1k9++ivLdF5M0o42g6FUpHpC6ajW4vB8m+C/ZaeXH9qS9DE96N
/FeRg3wQWHI9P3vlS7Iclj7Wr/2BrVDcxB04Edv6y/EcgP7Q/BAFs9s/weKUBsCF
D/uxXdyJLx+mJESwvw1NyWs6NKrV6xnlo79tnQhREaIIgHmMn7L6rnT6ZXX+yTOr
Sx2Yeppf3/S9qC2lvsTjGOvgy6hu421QDiP0JNQgrY4R6r/09o67g8f2t2SW7cO1
lCc1veSz4HJve4t+Dc3qhIdPN47ttBYixy4xVwzCgePAz28kahaDk0nDe0lQxEea
gs+m2RL4XFkY/5qaAGi5/Q9sZ74wvwI8tSlYsIlypCuhzNS6IxTkNDZ5IuzHF3bq
67hpyMvKmkpmQkhJCvmrPZTGMNG07ZQoMJ6Tjr97JqW+rQkABELotT/sk7cyVxRk
n0wlobpeaBBP19jFxZ9ObxgxBM37cs/cLOtunJDJ5nEmX5KdIn9tA5VcLLiXk2cZ
6YhI5+p9HIN7uxb3E8gI5OMnyG3CzB4HpNH+OzdfUTnPpeTFHmq7FnIl8E5MmpWt
EMG+bXQMf95WiBak9cU1Ze/8XfIm/oUYjcBk2DlsyHmx6Yvr0O8A7Jw3K42FYo7H
Es66IAZvuX+PKYl/DTKNmSimr73zDp4CpvWmOk6TdY8lzEV5RfM75wVI8ZpUdtBb
CBR+UaK1OiHZ2oQdoJjmsD+Fdu3tNRicVHd77fX/6geqcixsJTkr+IrVXdmwjRAH
i8Pze3WOk7aHbfzzz28HDNTMlVK7MRdI3hnclntHmFZjW3mKg+rtWqQFbKUpR6jo
EONIzRau8pDj67TbSvsDIpf1k4zTMjMIXenvbSSlxzJCDcG2jyOj+qPjAvBlMtXm
VYOI9Ea2QuICTNNrS/PDp7yhlwKnh3+dv1seOSrp42n/bYeaH25pftc6x37jDOY0
MKWqt5DQ9ci5OLkfARlXtpm+Zkm/DXD/IZQMXTAoJ1t3nCK9CZX5lCI/uU1zXzzH
pcGDXUdi6KESFutJ9ADjxFtHizWGTq7fjTeH+IA3fKoQxFst5bTZPGoywXpde9SZ
4KIkfIpqCdlH5cZ4UE7+rM/T1ABAZMs7FKplRIVkzryGkbTiiQjWELdL+jZibRaP
nH+5r+1VSBryo0WYeB0haWE8wbmG19srpnF7kXpXkVYX8LRE8dMpEfpRJ5f9b+tB
V/bMS8enW/FjMWBlvqYVQadAByWLeiwCrvrSOneu/QyRxPIspoqEwX9Geqq7TCJk
BLWBDj1gwjZ6/jAk0KVP5+YKPtGW3k+sjfU0m1sjTZG5p9MVXOS5VN+hdRl3z9oY
NKHoSReUcP6KlRehCez+VMPbQ8UUpzoxnAB4RP0gdZ9Tm3o5cbz7/y1LwUtqCqsw
nP70aWMlwruuPJATXd0pNpm2YhJ0M/aJ0kqMWstJUxeEv9Aj1Qot7+v61+Aqers4
/cffpM4EKSuPL9Bwjy4lLbVWhBDVX8k+icMXH2eHRW4git0PnIvJVmbaySacqITF
uqZqXpX1VUkIhX34Z0R6RlzhkwrqJX0CHXCKyC7dJt5rcAQxhxwfpA4/Qk+CccXU
f/UyYSYh6gcQvDg2O55CRoslwyHJX4bSa/Bo/7jRmMux/GAMLlfJiqdH8zDlKbuz
Cgou1DNOatHvWfa+56msx8T8f47QYBDKmV6vBtx3LhzYZNTSuqBshFSRyrG1vIj1
kpB6lsd0/zwISCp7ijzlFvdhcBHSLHzhRz0tfS3DQ/UD5v4byK/bYi1lfPzLCIun
Jb0gLdzuBLGqQ4PSuVtXhH242WiJDwkD0JUI+2VN4V1u1fIoKwoe1daSIiZ28+F1
8BqRwOrmbccEaE26m14NvyKtOSwYW22EoyhVqYaibhSbZncL2vyzBd87ubJMDIRY
G9DN5RX0oHBPWAMPNErnCce1U6t8Ktm28F5kDlDTs+qU/4JcBgzvZU+JwbjG/tfj
NlNykH85Kipt1tKaXeCdcRQYgJkFa2+CRtM1DvYOmf4dbCo04YKCzZrdNSTI9G6B
CkSII2emd9WwZoPJ2RS0MvLle6axB4eXFdOD9O5QLkB/CBCiyuhQHFHMgm4XhKYx
HZL7F7DaEc6fDhzJD0VtvqOfLAJMJoE5XjJf1BiWGcnUDv1xDvXTywRhrr2lXGui
44ZK0J+3ELTE4fuleA2h2suns3Wn2RemZiOJckcWkk1CmApLUR4TnZ227RTzv/dd
lRk5XIV6p4oxoduU+7mZ6aNA7jnhm8bxQxxRLTbXENEFlfH2lRCOhg7/AKQCGEr+
752irPHvsNpYZsXGNHM/oKKL0oF7n+ysluuTcMwSjH9Qf8Zv24KQobuMjFwB9neT
Xtmht9bIsG7moCD14lv5JGY3T6sZsDIhJ6+jGufD0DcTue6RAME7cFbkcjCvsD1/
7otaFfY0OXmNc4K+svB1lwvHgaiITafKPYNisBXhe48+IWiZsLyRDAvPpRRilYQe
LnBhAULxwMhxiUPdYwh7pB8YWldw2HJ4McQ1JzUA6M3DC0iECVg04ISY/xf7vEEP
nTR0AMC3hRC84NTqxe1PpCU4Hk+5XXutKiUr/Qv/0eydoXWc0kQ1VRyXmEPLGQHT
IGFWezRmMhFfshh+zEYCg8ptSkfLCCBW4DlVsP/pWZflFSv0anDMwE0Gsi62a7ui
Lfs0IoJe7MAmenw0VDf+6xUZgKLHaO0L+hSKUJxkIlEwUlfu4lqPPk8OxDo21UfJ
+ac8A8EPgEHXdITV6qr6uPlyE8JwfXxgislV/05i/graVu0TkFU48lC4g6lJixGv
80tDmbxNnTP29mFSMYjpLWYj4LXOSPmqaNQkIT62d5OsmlPvXuB8C7j2pwrVyBs7
nMCbAlfIj5whgDFmRpsuqwppfhQKC+g903hXRJiR9gW6Y1PS8s5/B6h4/Xe/s73I
/jiyES0WuLNGkmD0DYK9uPEH/u0AjNYcrhlvihKeatzK3tfp/9soZZ23qxfKqPiD
Wt2xuLJNagfDh29FvpaqvfKdjOnAMB7WuqOiPwJNLPByExVIU+z43OULZePRpTL+
akHBgENaI0VQpqzh9PcIPS7Kc6BgIXwk02f+pCBgsuak5gBx/kbS+/jnjSYhur69
7JEoX1hyQcGqhTVoWRhYxbaZbbjWOS4H45rmfrRhwr0dbIkWgPDM+M7IBTP0oDg6
pOuYQUSQg18Onx+zGsn8MVtSqz4y/FUHfOKOBdpw1uOjYWwr+LI/1sBEM0ky1ilD
nxG1YYZYZxnwTZ7A2et7gMbF6HpXlfTtdLEyQUCO0twyDSIIv3LXaZ6JagxHQARo
A1vnZVRz1zIyl2KraPTo9ODUU0SpOO8UuKs8JBqvgz7DOiAaAOQ/vHw7psUeQZzo
hFvoDrh6GLB3d9WFb6S+VOolHbtk/fjjLKTUMCdErJ57KS4iOVzvoLxa+uWrCZyT
omRLci9/1HrzlQd+7EyJBSaXvuqNARtpB5MPaBEAknbC/ZrJUQarKHk9pWGZQMPn
tExVjytM6kQJ/yGEBlVJLJ/0+0wo0/mGlG33gEjezx887gEc11qn1ss815R2jM9Q
Ecwv1FizkEnqkFVTbirLG123Ja0RW+RSWv/UoVlVDF1siCV69ZnqKM1CoHf/f2NQ
h4G7u5cUvOpSVLTjiChJbIgJgtxASVDk72oEuqEmTXPBtgAPZWgRIdwSz2leJn9R
yYUOYGjQIiEoFCmI46id3WVxDdUoGJSJSfI0QhHdX2hoCh7j+SS1kG8RUMfkyIBO
p2mxFNLoO6lky4f6PwTg6BihHqNq3D9HnDfGdrfGDKDg2nY/e+pY5NPih4lE91R6
XfgC1UaP9kuUztDEGSqAZrEgqOzKwIt2BufimCKO19QJ5/mpRc9DttwUvt54n8aP
fqijViS1rk+meYHFhUiqXnZzIX+1/Jn+2kKlRftkFzBHc8WWzZsl4klraQmM8i35
XlaViA12EMFdcJspyldVfvX94uhmBW+YVnbV74vMqVRsS1PN5PGfbVWJ82GDKd0k
TCNbn5frh8iDRUh13crn5YH4TVJA4cKOefnftIiEQ/99ROqi4sIPaVVsrz8621O6
W9OXSRRsF97EIM1ye+BkfAuVgZHvqIt32JYJQLrwId8PkJKy6OacZqGBRuY2lYZj
xd+OoPOmPLeFvb+Ph1/KmvjGRrFV5e9HOh4xvtzwZ9CJ+9FjoJiOpvwduS4vUwk4
FV1YX7y40jHYsX2MpWb3Bf1xsZovnhNGp5a45F8PBoBZWeV3dXaY0P/Z78gancrL
shGbnWBtwLVTPu5WmvRKzqLaa3kKFfFWPtKVM5RmrFFqh1GcBarAHQpjO1H5rq1r
/x+kWPdrPRBRTjcnQu3FnAQmTf92d+CEpjw9Jhts660cgoFjvH/0M4LI4Va8ReQv
Q6Wse9UB3BaKItBUpWuq0/++3VpedJF8ENX6xbeD7sIkkA+YqAQrYR7RBZCsuAtH
vlvocJUhpj4qDevbCzrHqBuRJSL3k1M8mSz+wXMQz0xXa48MarXccL2wpB8Ds8gd
Pu5GiNOMQo/bT8nPhaXSVJawkEIhKOgx9h2yjoyeU3yOgjjyhfSddzDer84b6NrM
h7QLXxgzLiLJAIHNtfnUh7CP61wn05s61CPtTDj8g64M0NZCDXe2Onb/5IzSBji6
JYmND6CqA0utBT6yyLcCOquhefmEmT+cE7LgFob1jtm+bdHIyws96QiaXP883727
lj1Ne4jU9T6HpGNihNYqpOV0i4SZDx1H25J6yQiMuUvB1TThF2422HvJK3u06kqL
pmtrm08WkiMA3iN5NmPJIETzQLZUneH5R5stC9O0e/rGeJvDvvpXeEWwYUZE9iDu
lGlgQe+mQiw9PEyPX99hXudbEPAL2XhyGBd+z4MBaN3WsSkkmVwkM77Qw9xIYOOa
0nLeR5n7ODvwHfW7Qxc800uD3wmV9SzproAXE9npukSQn+j9Jlbd9c8X7Tbc+38Z
uquzQfBfZUHosIZOXAiK4faF6wiJ6m995W5TZGiKMQxh2ND9+WtFFwkp1sY+JlHi
gzUsxjnpy36FMvyEoZexMg+UJNYuoA+6744nUUYN/SYaoMEq79FBRfOsLWW/ghxC
gAuk+QAjWcvWCnknQdDsQYHSiZOQYOffvEOOYCHc+T/cv32E+JK0S6H07a2krTzq
E+5IACkJjGxMvH2rj7Cf35wVrPXPvCAR2udESHcAd7hoOET+R1j4llCQoNHb1AQK
QTB/3D76K65OOeFESO7zoN/bw25QI7aeVvEUwvywA2KtlwEUDfiS5uLtsQNsXcYY
b9wbCtMdOCWJuHb3tRkn76RaD/JQXJjEPSZTYe1ob/chv+x4O8lRIJqt78h4BGsK
EONsqC5P5On713MsP4Wy/rrN87XheNAncE7KDqijlopT22JIiKpGL0PZrabbEy58
S4IN3gYaMeLd/wjoPDNXNuMfRisixRPduqsQH2XvuarxX31GUgOElLFM4D3CP/ll
kHGGlIBuInIEEWFQiOUbjOqn9AKtoU7pBbuCioxX1s2pyleXzYS33xqTTlJ4jXkn
N9eBW/G3ICXsx0LfINzaaDAqGLBCM1xVNJFKRdGRd7/ROyvX7oZxhjNseN2/4fRk
rRwyGN7bCdAPoNs+zKJ3X4sMhYVAiHmdw81Y5G7N2l1w5zpwtdaG70mSukjtlnk1
JoI/MKf3z0RA3xCRB6CNBGQUdV4XShzUHJITmMtelrSSCfeetRwrEV9ZCoWk3J1B
CKC2RAh1ijEAwhzcRTXEogcarKj0d+lL1QkPYLqRn6vg0u4zJjmHSQcnVx67dWuv
YI6sLu8lW3FPQ9v3V8MhcUzLNQVxvyZ2l2kTHXn1lh/jhTyf/WnldDL9x0i/yjC9
fxgdIMjWzmRy7MoOGJlM4Q5NUdfyS1+CNfrOMKR2M5BKOwsTMsHF0Kog6345xtzD
5LvRcHyYB5wBAj/EPekYL9zoV1ORD4iv4KQzBxFmk+Qmlycx+CoH68q+4oJvZZd9
Wl45RPd9lIkFQOvVRY2nUHGEcf6uaqeLng9Eb3S4x4BWPHUwek01NOy6nC2ayaSm
v4mZUgZFt8q8EjAHW+d7sTNkZL+XLYkvWNYFEkCWuGmW2GHHG1tUVMPmevosdO2m
boHPiHQsW5lJlXh6DCYpzOolbI2EaFmsxA9pLZVATVpFkpeb9P4YZSU1/RPp/Igj
aMvYl3B78S/QIimx/qd/0EqSMKYT+NowAdtnDfiEMOAvVVOzm7pJW9LBvt8/Bgup
LB60+cMiYIU7YHClNLnWKQZN6bg6q0rbEO14NSDdzlwr5Xnmv0IP719ssCgCFqYM
3nY79EyOlo/1MtLzEJpHOMDrcfPKv+FtZRr83/qA9c+n0nCgX2zNHM957eNGixXL
PXrssedZNZJvrDMu+MEDOABDrrs1hBeCqh9lNOic7JlWSrn4kq3o0xUcnqParh4O
yCx65B1WozizsUZZ2EE6OnDhgIX4hCgc2p9Dhw9vo0zKDlSXX6WAF52oMw9ukD/L
JvMKbn4yqskzo7bxIe95OeFp1vZ4GEL1MTVMmlP/ya9NbWO7+jpiHV3m8wu5R0fB
hkN81hFa9/gdY83kLXLwmNdwxaXtxwiLex2Fl7qs0WgBw+ubWrefVCsgaNF7j8qp
5gdCUPbu73p+rIfx9qDmNsUP6qdvDS2ccO5kisdtMct7P610k5Qe1W0W/gUbwgrX
V9uJTKGldf46nL5bR1mxaY48Ns0XbQOXmj2nnzk24ORtq5/B+yKmrudy1H3gOe0h
WGr0i1ZvyC36ZRk8Xm7Usti5O7pe+IJ7LsOxHJOi3egCl0hFzFTVOND6ckvEAGJO
/QMS8vUP8oO/OoGAulqH06OMJIPsrWf/bX18d5VCV6ZNmKJlotlZB9fu4A7jp95Q
UA3GUyjyeb4JLNppVR0p19QnlItqxJ5azZXVWqP6CjkxQc/PmJcVGHOBI7M+tSCW
firjoC3yMd6sbi2khczJD1izsrotT+wnl93tTnukVSLkm9hZEMS/TYnisrkmcyRH
+ttnotOeOr8meSDWE186C8vQG1kPZFvekjsiJKKz1hxqD6a7QZADTNJrMOqmvO5t
djfqJ0jflgX1PnK1fSKXr1iVvREdOlHinUn++VuffswK604onKpzlDjaAJD4s+XE
SJ1r0qYMYgjAaIcp5CXUqnOIKAHk2JsyQZE39D7PufBlgbDnuWjGMekPiM17Uoxd
k6WftMqU9SiuDMpHd4XXYDrLrXQl0+7uS4E2B0PNGGRK9MZFlHyJ9xLowK0L+cDZ
Y94yxxUlPmM97QEGF5wUvfQr8gN4ybkszrd7QW3UKhgXGdq6lGoYv/svQolqB45A
dUVEE9n6Au3DH6JZ5my/Xx+TieNbOwRDgnF+CvUdkyZG2CT/Uns7cUueGYJjVj7o
hVq3fJ5b2lSb5UfDLrt/syejvoB4ajunwaE745G1JaiHTeVAJyg3eMVnjx8Cmt8E
sRbUki4ctC5eCIYEOPAElOP6KYTMhJrRN4luXTDnCoSzVDHaXhhxi2ohSPaHEf2T
73NBehDTLZh9puCix9KNPPCIG+8GDuZAFjQ00siPp7AkxSYUy7h9zCrV/b3jtZmy
583CCZjAS7k+ldI/IQGlQ5plVjKkPKXd5NpHLMsEkGIiev4hr9xRq2RlZP06KkT4
r482dbFnzwGSyYVKeZE3c1eHIERP+to3wwOcHJsTU1+eq4szHNM33Oh7BV2oFTjr
VV3LjYx1ptjkQNr0KxqrllfneFm1fqWB6hmi3T/oxvPIbw/s2Z26vDRcaUO5p12Z
dh3s1L+Td6eXoV3QXfZDqu+Qb5JQ2HL6ZzRYtF9Zkf6V7ITiRKOG8xdHVzQGQYsb
5AH1KoGcy8WHA16hb0JxM3r/ktwx4mHMCZqgkfmfQLsiwP9ks3QTV+ppahz3A8kv
fUnBkRxTVdnUY8DgXtrjOwIJgyXobDHZsyuCrCGWFtk8EtxQ1h0LT760wcoN+hea
M2k/ewAX6i+gb3pBwLLNkeKGks+GBIFSLAunk7t2ciicw7sDBTdMaTxO7TcHF45m
zvz+GbeGXcqrCIldP9xZlxLvWOB4oG9Lrf2HGAJom6XZQTsNt9YENinPI5nzBkYq
T1bgwiDAHJOprhfM5b7ZucZHes0f+Il56aKTynUZGnCb9Huudy4jfJLxnfnlFTf/
yVtTtJIixUQPsDJQGco5dVWBvHFNdBfeYD4q0fe/x77woY6vQUVPeZ8YW+qKyE45
SvCzID3ClEvv8NrL1e+AN6Dy31jjZTXPSPPQBpqTs51xvSHyFNxYZUpNA57OX0Vp
+BQW+9E2k4OTK3X6PU/KTEukEWVYImQ/frfI4Wx2J4VsNZNzbiiAPLt67KnhPuap
lSmM8No9pFB5adXsopXuL5PIcNaPLc/IbkhDqPt+FCaJOsH/WhfHosQbMKeWj4ge
JTfCv0pcwKzmiGK62M3I8yhR24QtWD/9bN+alohODG+MIfrlB8U9Xls04tIlb5XF
BP7MYaZO8vRl7lGGMurbL13Y304nMlE4hQj8+VUHPzPmm82K9vfY4qfYdXfAgVa3
4TrFOuALjb5QEz7Raia2EJRNE2b5z2QgXI35B8d9z7WkqwTkKaQzf4sd7cFKEZks
tvcfJT2ZZwGVo5tfB8rfRtU5wQL+xWVRmWji45b/i6y3kYPTHh2n+XubjRcEe5FZ
+bUbB4lj+WqMWE6xrVay01zlbuZCa/NilxGKXKos4FgxkOHcnCNvshLuz/IANg6j
G0NL6R7teQ/y2MCwgc/EmtQLI5UuYWoLq0XS/MGn6DSnohNVnRXvwtba1DASL4Fd
fVce87vlanSuQQThg2QQH1onw6eXrBcervm2bgEYGm4v3pQyIv1I0+p1TtMeqg8B
X2tgjjwtxW0RabLgH1OIIEKATvfzpbVYFxInHvHCI25/LWbJR4D90yXvMBgAHuxt
aBdCD8LV7u2TunHRA/yQbdRweCRozN7jlh1A5UeiHddBHjXfqFQElSgg4Icf5K34
XwDaVQTEP20X3NpD5dGOhltFBBDoa+UREk/Wvkpfo3BtRQ28BDUjBuaBo6uzxEzl
YCgiP43zSrsZZdtm3rbedcRD0Gnqmw4HPHhosy79JCJUcb7vIcZXsP5o1L42SW5b
ayiAgmu3dlyPyDKE2Uv4LUNEjpcS+VPu7NPk55PMCfoKNigWqp6cb6++WWQsjERW
92k0cp8s5bHmNc2lBX2CHYJxRxREcxhM0ICb1zFTV/fsxrcep3S7s1nULZO9rlX5
3fzgtDvn2eNAoggwiIzXWTvXoydoHn0Dy77cOS55epNtNr71pl8RIjPXnlEo6SQV
B2e7xd/uN2KdAaWxCqvo15b3TpPM1RC7Avs3UW5Cs/C+euB9Vze1BDZ+dH97Fi/7
zOtEmXGBbJu86gjfaWut+oVvWflhBbpFOk40lOoc4TvrY7ybHStmRqDyxdinoQnl
5HgmfzX0aaulEcWy5MSsyPWO4715IafCknPjWsQ0Ps364YcLmMxBBsbPMbtE8OMM
UwRwJCZGTgynpYTrqX5jp7vbVBTdZ6+hRan/AUysqiTSshkOuQNGRLaeNwVISUAc
sdODtypwASqGAKb76KCvceRdruIQLc10xsMnjqPpUbhJ2+C7LghuQ9KWY1UCIvWW
4USpOuhU1FpxWoY8Umn3EHvDoMdM1XZttc0KpE4gJPqaFMjKSRo/zk7Q53NGrMP3
YbiJxQmR03sDP/VVwdIRQ0h01WSw4TCyKvECSnP9t/N62u0UetY/HxX3oY4pJ76o
R/Lel2x/+foEoasVrYqg2eHkPeP5UG1e6rSRi2YvIq+wzESvdpq9nC01OuB3TaXn
aodHCrTVNIBcqWgZLGtmMRAU/Lw+0d96ywTAzByhr/7K2sPagxT589MJcjVVZNuP
17XBAjH0iJk7FcgiO9yFqeGvMU0RGRu0/aYgJ4zVg2vj0MNdAltn7OVQAG+ZlwHc
LzYE09DhRu+zxg+ughnpnEo3GEDzu2dSnbCrR/NCYTE/fTL1h5e51KOoTBzxtatS
nHkuCwK2FDADGcCACKKwAow48LY7nkFGcujxz8wlE8OhJQE3xRbB9yg1yEvKjl3B
hY+r5PK4akSmqEvDg6+a2vWGJHCK16HIHG31gWbI8zrAnAMRLlaq4WsDJFzzMiJZ
yA9QUZoMDkgHnojJp1/v2/9F3cpPXzC4uv9ELFT+iXjJIzeYd0ChzQsqCNlvz1s+
qV8fA39KFmdojO9Zwk8yTgVZ/+ffuCq+BUc4M5jp6Byb3CGJZcvv25sNFo6PhL3b
z9BKsgiROcXq19r8nYdtkByCvUdQVgK+rujaT3YgvDdQhYYcYtNd5yuo8OIOnkMU
dlEoRtnMUYxN0yfq5BSGuQKICfVG3E+wTutpMmwhaJL1ey7Y/th3y37nWHPZJmIH
ImpxDalXNmGtmQ1EAUhYsKFv7p8COWYCvqlId0RpJDBCtriGISG6sHG2n2ymkg8h
1vMj6nQcX+h3FuuHe2JmcS1hi2SAbzQO7RCYbTEBEpLG6kjIC7jMSa7GGbY1rCVj
bmlV5S5pJTEsTENWaaqrQPJ3P+J/pz5WskxdLfEoSsbBGnz6k17cyk8sbfbW17R2
5zIPsIBB+WtHSzZU07JFw476AqFsmsyD/sW4ODLcTakgDveJuY1shxAx9cHKn3o/
L51JqDfoPINm7R3ypFef9XyEVO0dKQ0TZhJHbELyMW/60HM3YRn9A3iF6nWypVd7
5+3apSVreDX4UfWMh8ClM5iCvlZlEZX0fbBw974lIQhi6RdzMiWqztgcQUT0Ok2u
bhPOAKRNh4kaWq+i9YzqHiUeo5h70s24ts3GhIwC9USWTIvrRLMFQqXx4As+3ixY
pIdzaaMfJG2zlOC+QWBC9ucWXLam0A7mY3rd3z/F/wTrpMzpqQ4C0s1kpBtscyhG
FjsPQ9ZR/qbNgt7pOcHsMKLJTpuHgmsXTlZzaRvTO0P2VvbGxIXag5kj+pOfx32g
WnIR7HQcsi55UwNxTucfcomahFbxozSQRKmTSJFJy8HgBp41yn2TiiP4aL9podNY
W5eaJ51WA5qjWxbs7DJ+Zz2L2O7bHSAV27OAHSKK+tRfn/cQjpYp3wYb7BgHNFLl
goH60GMRxGX4s88cWFBm1KOjT4kefXcAtg2Oqy6SxICr7v15O/WLSmmVqdI7gRrx
dkVRf8BHNTx08zbi0PM4iI7wUeM2PM3YIV+TZ7U/OeIQEvuiBhPyUqbJ7pTdKAav
9xvhD2Fc3dfK0X1Qewi5p0Son9yNFyh2oS+zWmE/n0DcWT6h0L8Ex71x98pn/2Pp
YycOaakfPqFAass4j9fX08me9WwQyWhvVLLf2EEd749r6PL1FLLoXsXAXp0giS2M
bkH5zLeCK/7GCvE+2X838zvGvQXsRB6Ce/SnOspdRywyTnVDEttLdUcCBoXNvQFt
sgABZ496d5/bbIDDpXZjmFV4ZclGxzDDcuZ2ZWl/Ih1wVQbPM8cXXcxBupv4ont0
q+IUupmE2Foo2tSh9uuyOJxyHZYqqCdo1KiHue7oo62lwO19N3pUC1TtG9F0mBMT
PzcaeXWXZ2MA2pDiBWAAYl6wvPs6zZcOaADeEgjFfkyd6S/OyTm8lhOnu6Jjx7UX
c9Y8sAkXHIX6X2JWaJ3iXuvBi9YmEG6QyBgG2zheje9AejBOsqESOj5r3Sks+mG0
b/Z+5whx9flDQ/tyYHpIKMj6w82aKD7JcL4CstNXJcfsSj+HgWhWayp6ZzycPdzU
TMpeqcJUBxFjJ8lzfKULM0ZkNYJ8KiSYJcriOlxZtPLgmZ0xNUHZK46/0DGinzmx
oR/H6ujwSfHkzZPTP5woWGPcZ2iYs//pBHdonvIbEIPJMZQpnnoTi97XqIQ/fXNZ
BtjCkopghabtKyxrW4iw/45cDk/kInm6zNbMXuAKkctg+w5F4H55ZNmWfOEiZl/K
x3udorJiiccd8wfISPudxtglMcdK+SAZ95oP4ydoD991aXIJybPh9tZJqbveF9cE
yXd3TmVMHMIpq+jMqmGSRd6hYZfKyn6gXPZbQIfhyWBCsUXbgdWQnmOHUkNk854t
uAhxZvJnrQRh//6i1uq8XrdUfz+eSAl2kCQ2GO6BCoQctOzOA9aaGG0dI5LYa1F1
o+OViBYYRcENBvbQXa8DxbJEWs1LcQPuJNefObNNrf59jvmIDeYfNWlMwky+h7dd
6bDoN63vcfGM3kQi2AU10AtmcjQy2o7EmTMAWVuhMrE0pcNFFj0DmLBRsigNyQVL
jVW8KRXDp/BiKocW0eJeYwvXhneFOiDgX2ML+2dpzDckkS8Gqfksb3SVv74Ciq5S
N2sSOph7mZKJbmjONgtkLMXZw/zaeJrVyykFrXvdouEfvNPpKRUGUVHXGjpDobgn
2kxewlANSKn5hgeP3rREwsdG524LjMkUqADPpVJduFZ0MBN3wCla9xknuVmggU4E
R0xv/ZhF9sXfDGgnz/4wL5oP4iqmmFRth3bEq16bV1SlJEJDISFAi+tf3ASrU6kw
75EFfDz+fMzRApjfgMvQ9N5Jkie/9gy5YUx2LxnEn3cY97FkCQPrfP7NFAMMR1RI
pmE9FzAxa9MHLvE6ITfOrjVE0tHla7gWqBV+2A8P21MsJ13gK7qY1vnFodDu4iBg
6NIG6ONFW11QF6fRm2PeaVRqcLzovcM5v4omc/diuakbFKx0YcmeODxGk7CPwTH0
iAjWBlKwZJ+DKookt0fpYI9jo5av9GgFJ6y0TQhXKINCnympCC8xU6NcxUby/46C
lTSQc1Duem4WttEJgMnGP57dSDN9Q5BGnN4ELo+6mVFyW88eY2jRpbXYBdug4pbm
W/y/K/c+zerfBl+wRNWCrrNGK7I3tXt7ZTlkXPcJMnUbokk+CngSpF1IyTAc/wdq
gXUNlA3ekMv4T8OnVuut2rJ9/RB1kcka/zThILrwYBSCNEjt/OpRs57nv6W3gkbd
kCLmKX7rtYOrEQdUPbUyd3kL/AXO+A9IoV5T8/6dbmyMnCN6Wip/NN/XCpCI+fDw
qu0L8vMMI8kebfs9BEE9S70WGEW8Zascd6gGAPESPleX9afs2dleezDfhBqQR/WE
sAU6U+pLQTCqMuGeKAsL/uPltvtLXObZuJpv0Qj5jj6w4uuhPk8ML9fTnaxEEqNg
K68PswY6rFEq0Rk0ipWigmvTTUotaebD0vkSC1XfY8M7FvIEbPesjlnSxDiTpDwe
M59LKcMqYvjVD0/p/BpLfpOwRgy5B2xHzkmFXmqtlC03AEk5ChU/XsGIQ8FZLlLf
Md5y1sauza5QkaE2wmzVEfGiz4RA3yr9/Y40w29iBp1PCRDuGDsSRd/An1Z5d9eA
04tXDS30I1Vp3CgDs0/0ZE6dCJo3Vzi43LUSRDwo3F4zvADfunrzi/FkwmU3GAEA
qkwv1NzVAkPlgThABUn5vXecZrWzPWz5G2KaEoaytGcu8sROvfPnACjmiwLJ+3tH
0txMFhsbIvnGK/tCdOsqc1vrzss4E4CmgbZHosceBD9Fg5MhLSr5jSEcwCQzQ6cM
duXO7CQasF7Isgy3t9Epq3UuXAqcS7w/HaaUCG6nDtmGt4Wrmvn8HtwnDeVhd0VY
lnAD6yWUSJbt9RZzr116ZqEOMBhTpidhT2bxiZrsBSWQkBxIOF1TzLcza6z2Y9hs
4XcGd1DBMsQK7I9qsx1YAeifETL8Zbn7EMtna3vdYVMvBceLTFUenUvpeyNQyvIo
ndMq3aELafQkyLQfTM264vAwUDcQ3aqoAeDOXhjyaUD63moRb1RrDAVv8dUeaHg8
xTyxBwvXmSkMevTan+5WJeKGV39VrcM1ko1AlaVkWpKRIEtKI0Y0nocaQFFeRStL
3d+18S+jQIRrSW84yHOI8YVHWMEBUs4X8JX2ECg0FZwDkPIsCbJ2BCrM/otKQ8Ge
doZyELR+y4DrKZfndOAhdmDz/YcUd5vf6jjq6McIMVYITzGL6RNDi+SFzCCPjEmm
fAEo5Mhy5+G25GJnMnpNZ2qJoEFifmAMQ0QwfJ4Qxpj7xgJWQACeIgPGLCBErg/b
+mZ3U8if/1ByWVn9/HaawSgplaydcR2o8ZBnckaoINLQzEKLELFJfTYlZifzMtoJ
HbC/mZAovZLuAccS1fNtGglO3PIqsZ91Do2wxjvG4Drx0dTb+E6rNEfSiuo/GBgm
NOqlwJWJCUIlm0LYK1VRCUIChtxfnGsBTy4t9R20+43nz+s35fgWdhV6+t3kgq3I
4VP6emfPO0/Oj2rdBLdyPW1p1uQyKmM+5WGbWHT+giSfVuVnA+6L051GpC1oTwb0
MDWbt91kXHub404N1OOeCHwS2ucxUnK7HEchoUF6fKGSAMrFoBKJoYA4JkMF23sW
9MC/DkLTkYQfdDIWh+tblAm2tAzK/agsdKwp6/glTHiwM1HkIVepDVAgcTm91Klw
a4YyyP3LLmnm14Snaix8Dm34xonMeSbdLVeMsCpls8sPTkRmxAI1Q+ZW1Ll+YEGZ
dBbDRu9H0XjJ6btFFtzuTLh2daULxFmBe9CMqHOP/zkpeYmQcUBfXKW+QgNL6nd0
wVdrkhMlTd4xquSxRE0Qulv7OXTenT/d4gE4uWOexRpajdez2f9wehWYnw3lcxcu
4yBn+kX/rJWsHwWDtqNhvSUA5mh7rW30eHdO8JeBCA/vluQwhB+S2GJWMcDKxFa5
97f7zSGSO4ylTnDVTEtavfVicMrnOEbUeITYbYSBILnaJE+pGvfh+oQXWMmuez3C
wQ9AB15vKhVRjkyixmCmSkHH0dsCpXyQd6ajv1m0u20W7CeKMdVKmrpviGqVcwaV
/w9j1VtX2fCaJbdE0r3UEZObcIsQ+5cDt+faLAyCywXnt71fPSvlQvVpa8dRzAra
MXLYjR6Boy1ySmXnp4U+FOOuYP52z4XWCLmulehbDCMWUj87q68KWfJ4wk5uX2NV
HnDIhaTtWjDYmJTnTIHp5SDuFcVuOH//PpyjfPFfwFCMtTi+l9UsrKdrgoAz8CiJ
zgApjENSRth4kW0WRBoQwIeVmxWJdsidu2G4IxpBc5y9SVrMeCE3rAfBj96YB/TB
rA+NktkVXX+rZw4/2MT68j7vYSQ2Yj6zCT2ejkdR5AbC9rq5KZcidFMv8dVHs1Vz
ieVWIuEEXr+XrpnzE7P9JW3T+XDGjDF3dDUgzALKlaDVbtu+YpPDlmjAxlH9l9/+
tQx5skWgmqOFGq8askJ5dOfnANoS2XqO2QYVqEvXkf+i60/gQcUtVQMQuTAXP4qB
MmaD4FRd2bkUJhMoBGzNipRbuthrUUoMLCWFT17QMAGK74G6QyDWTkglK0fv+B1C
cEq87TRlGx2Cm2/cH6TeSIVg8T48bFETnR+6SKCrNbbcwnKSKecYKDc803mNbHZY
efJ2kSKQde4c0BMupFlJQede+etSsp9b4t8gxyFGEzHWJfFyyC3HM82361TrK+U7
kqTX6kRPOm4L/i1IUEP5vfVpOkvdvQocCfEgDgXaI9I87pKh0wBBcih5q9WjgnYo
9XEgmPgVnVUDv/4ixdrRt/CRj3mlNg0Gb+RT1RD1Yylq9FoghQ5zTkkRDNzZkNLT
58ij4qcuAGiyiL8k1ChxaTQgECxVlEVHG6iPCNuJ4UNTyKE4UPfI1kpgbUGInDUV
kh/WC5oFn+mAlsUsIFvjBuPg2xubB6rCQZ9CO7grdrAqr3H8xsT6fIeD3AkB0np7
QCVjy3liViBLR6G2DkkaciJ0AFP4DaSu52mfvR6/fclVZMblvyQOqNM0Lzi1X1te
WVvR/4BojUx+z4AILHYWZoHL+nVY0/4WK7mJnIjsl5ZaQOKp6pjtvwGi9NCqFTCl
vXF8vgBD1NFQSbSIsb9d2fZN9jDgNQ0JDMFUhutnStb+CjyQFyQqMlzz7WMVr6XZ
f2Q/CzbBiJioM9tw7m/C4/yc4sQthoBxnVggSqV0scwkg8Ijql4bYoJ+WAI1QQ+K
svMP0valJdfsESlwEaQEP4xijGOSy05rmXCRrvKW+NrtaFOmYnHfgtO/eUKruxs9
pnfQSxKGIxmgxlpb7/2tjtw4HggYHRBQmkeOHypypHxZZBdEaRB7tiP95payARux
UMywewi8p3vePrhcQ93AoJZrr6bm9S9vlOY20ce9bZZvbF4nu9mc08d5ghVUjfBZ
yXyor4OdJffLhD/4KR051+a4+UcsRGGvvIPCvHBcCUkwcGwrgU8kDbZVZRpoge4Y
5C2T8UjH7wd8nYJLKr4n2kUnV7rIJXncIZcCP4amWrQgMcy/tm3USo6AVB2rmP9P
KX2szwn1BadQE5scGC0XX9n4WCizcwB9+WS24pH0z3UXPOaadoyLUl2a2+tvWGUN
eSrudWBW+laB+Uypqt4FgO/bUo5xNn1/thZq/S26VFHYD8WUb1Ru/0FRQPkPDxu6
z4w81JMKUlkJMbvrAc6fQzJ5BMJgNn6KS5Z2KKopEBDY7Iter7obKRqB6YCOFjBq
/hUYgskHNUkfF6hK/KwmggR8N8WcwduH+XNziIrtZii8jLhvNhnUlNU44txCTp+d
RvExzzMt/JqVGUDVO62K97sI1pyLtfu3dY+yj5io1v36J2Jc3I1hsrsI1e19K+uE
yrH0PYy8ofKRbwJy0M6G5k/tUiWNZvcOKS//z1evC8YN997VCKDPyDn7mJQdmsfM
Nd9ZVRr41/R35gNCxkJMLu4QynJbuvEsMLIQuvW/3BhNgTqqVNXB4uDi3rmiR9An
56dqitjXODEGBgi6/HEl1jUx/J5NgU/+s4qhzoU1uAuBgHMe0x1BAkNECjccM0LJ
TnqYp6vAltF94VWgwTxlpxBU9nTeHxVcN4CD8fIA8YaR/2K9PIv5dCZJoWSY2CFp
77cNnfyN4HhzNtWrzm4jnG15BhpkGsQwsg/qTPqLUwPQ4VrFjGPuuv4B5QXleM/G
9GZ9khHXIDBXyufipP3bH/A9jJy8fzDCKhqMnVDWEPhSbquJbAK2qITAGAfedsdf
YVULXTQgi91QJYybl4OGHUTFeuAXVw4EazGK5UFnqKRAXH+Etj0XWBApkmYmnHlG
Gfm2JddMkQFW6UsgCexlOCyRpq+Eis8BQ1fnvjxgUOxrfCfyk/NisvyP+l6D9/GB
MNEkE6vN5Pj/kdTSHVm4WI2BW5LfbMZp3/T01QGaW/3mJLJ1Kx5Bp7zMiaSIwYbW
xrrGGnRPqIRyU688HMwwOyVwEfGMVjH0HoTEFK3ZiS/AtG5HTeTOBbMy94juOTFQ
K1rFyId3Pg/XKIFlHW/A/+Q+HL1qcbCG7t5fIBiO2RlaDvdsmggvdQGb+GDExGG2
hTUyjuCCnS2B9FXpN1/MAWZ0jSDsbJOxS9vf8naL6klfXxTfTGVjWLUGWWLI6Oxd
3cineCp8mVmLX9v30CQTfWu+JDkjQvi5eig7zbsdqq9PQu3NgfL2ByThynVCG7lj
FHgVUKfpuMber9/lzObyKwRPl45n6crawl8LoM6DUvZ5Q3a8bxXj0w5C0qaNID45
rBOV2kOPs5D4khdp1R45ae/dVOcvio9EBx74+EEhcqfadS8X/fQ6+HVDnhPe5j5a
0zmGNmXXpMX5fk6a1qYNp269CedxyrcfEvGHw0Ty6Z4WzpRgxgIL3XLVE57Zl7iV
wEzDKKdptDrTv8ITPueKh+uWxKeZgZpwMrZJ8CF6Jc7o7F22eVZ1ONT/y+mWjVyq
uAdYnlRIAe6rOmS6can7SfMaVXHVUthS8D/s0VMZ3/Ybtm/f3qyBeqikzqwE3lCc
NXiaWXE3OSKerQ3vadpjuxWkM2UemDc+TJH1AgG4qKOe5D4C0DTTrg2glh7p8qFd
af9wf6axkGXxS7rBEFi488mlyOL5AAznGr3ffLHCsqPe+7vo+qi8Tspu6Urpy3iK
3p2thWAh2kK0ExoR7SOWIwslLzGG1lxYZwNATLBONAuet3a78tCXcgkK7X9z+9zf
jd/tI++4Z5agUo8J/G97wbv6KXKVFoPN4NtM1Ujlu4pdVuBeFIj6OAgGcBceQOC6
SbS0hhAXWbNZ4SaqtImb3AZmRO8AnIbrB7cSswucahHrhBdeyXp7N7JuGp1zpXdb
8CvwJ3c66KlycOYQDhKUQXsfmph7l+PbOBllLIga0oo/JlIhdZDiXEjUoNTzMNww
5lwP7Ndt/l3GhqY1WX75C4UGoNiPF8qrc73XsAgjLwYASRIr0hi0aexlxiEDPENh
Il7YKL5aW+/PvAhWLx7LAbho0j19Qj7CHCJDPAo+ZJVI2RyTPVD/CQwsU9s8ROu5
wK3xYIPx4os7dnh/2Gr6zE+hU9s9+rrtZJwcxQaxRkaun/8bS3R7O3155Wsax9Yf
0Y2y2usDDEXlMq5CBTf+eeXU0v35qgJ7LtpdprVwwtCICeuKBwfMEKLW0gRfP4fQ
us5y8SrgWhrApig5KeB0zCi3/hY2zn0o5u4ybjxnKJGrSrh2Ags+hc9Dl2Uby1XZ
F0Lu0anfhI43RHeT6I1qHo5ABGiyBe72g4wNDi1ex5oELTJh8fPMA81s5jt7sn4+
PdogsY8MeZEZ6oP5zw46Z46RncyYkK6fcFHiZ71Kky73LTcHJXHQqWsIUwJ1qKuw
pRxFOJSPpslQPeTxAf7BYyeWgplCwNB32VhU3dyqzR2FAaF4lnOuAUn0QY2KcbrU
KSTDQloV/bN3xvZW1i1JdjqE0x52g+wmkgoxKzVIw9e8GJm8QDEhBkinFk9XDLqd
e1omnGV5moaUlphbFfzFuwm4CQzQBaZla3TOuxURMKrkD2xUjtz5GBHJ8ffAnAW/
2DRnl3GZV5v4MctzAxAeiNk6fo5WArsBlFNF4BDrHIqzY4O2E+udMM0nCCR08EEx
CUWlCiIBTTfmKF/c5PEP1HDEVRate3UhL1yhUdwTo4POm+hzOHqGNjADWHslVon6
uVsjVGo9QfCDxeP/+qlst6nCmcwEq0rBmF181nLEbsvko60ZTm/AmIwckOYeYhp/
y1Tnjd6O7ecuOqzPEmLu7ojIL+iQde2RbIZ/UY6cej/uNd1K00EYAd9HdH6Utf4W
lGf7MccGA9V3HdGFNB2no6igJElguZ9T+2xpwfVQdGi8a8NLwdmxU04aYsKEY9qI
1YbZHYZ8MM4l/Uj7FeesTJcS/RlepWQIbAOr0huW2DvdOjYPaLvQNSGKOtecSY98
ssyKl29A+s5f5KKOrnvtsbdS1gp6fZhmeYjJjGtnB5H6J+PY4izfkJqDaP3viHks
3f1jHaI8LgRgq23Kd7rvjwKgEM2j6SlRuDM/ol1Iu5m5gOqpfekWPATBa3jfFki8
PYSCP1oor967zBeahZt1gk+2gEJ/VeFvRrFsfh4Ah/McU6wSHFetoZ9MmSM8RuFa
nhSBvcuV5jkkOn4Y6J+30rg57iooEjfcAk+V237XtOS/Rz7zZTtm55jZ0HCERoru
riVrtp7IdGm5wfd0kMhfiPqljh5KTWz3KmRe/5r1afgcu6J5h6ZXgA+vQq6djPGk
Op2lZWZ0bnGJy1UtHsJxghmrDz/0zuWmd3u8CxxVx8j+ACGfomC5QbrsGaKbHKnt
BeX4obn5d2AxTgpuSm6pTo/Ihpa27GzIDRA7cpUXV5LFbiAsq0ZRZMxv9Bgw1Otd
1IAJQIPDZPbhQ4hmKxM1BYFmWBWbQjUDU+GdUJ5QKsI4t6chnxViLGq9hlmrdWQW
fJvt+Nuh6MSYK4+UJHq+Z4xxKOUfvo2B2QSdqEzadRJIaHNy+IOX1aaIFMD3UcSt
jP+GQa+G1HBsH0PGCzbz5GEjUK7pp5fha/iZ510h/fPcPmjGqN0LFK1fPILB2BTW
9uGvjAzUKpLNhqz5x4HJiedceZ38v81JN5gj+c5StXNxEHayocw4s6gZdAU9Mr/3
KZb8f1jdF2+ocrTNaBU+Wkj0W8ZMTZZ1L4xcTHzLV/m+cgD79t8auejX0JbWGvhO
GD5SxznySta2gnXwDZar+fFEtOcDgVj0C2G19crb4pqhS1pby3+4Pn3UTeCNLXfl
vr88sGmwQnAi0tTMZMQOs6aYHD0t/NjSy7DkHd+Prrwzpvn16Q9ir7csD+y+7Pn2
aMUwa8i7Af34JLro5+guGobjbSrmuuLUskWjeBTGt7OCtuHNiQ5cKYcXPj5jD0XR
1pZhTiGixBe1L1cdn3tCBYSVjJxt0gUSe9YXq6psIWORjoyjnl/SLBWdUUXlVKko
yLY21sqmQzRBG0HvtWZ4zPj79aLrcdsQqgBKZpfInAe3Lx6Rgoj8Io46tZnFWPaD
9dLWucNAgajinaTje5UcncPy16gJn3ASHQN+OoBBaM/X2a6vUqC+bsvbSSB1TXYj
4K/GlGaVyXqZtdf008SA2q4qOaAuhZI2Ty5b5oU5uZr71JrcJiSqnFpwZ73DyXxp
D/SqbgDMX7YKJxokNnD1CQ1g059z6dvLOkvNXRRAdIvbCW1wB6QLs+hQSioQc69u
ClWt1gpYotdr0T0WXp+CIOzgtNN/C6miuyDhI9U+HXlBZ59Uf0BHq0sy3OMMsizV
R6WW9NqJdukhm/+lLZa/jEgCKhg6h7iTc5MQFIU0PfgN/FOmsiPfFF/HFXtWoeLL
7+STcFdj2tOYk3bUlfqTSowNIw3hyUKP3oNXbmnIH1EuknCPpuD+Sq4JkClf5O4y
YI9H2sQuJ1tCQbiSRpclIwtqfDfepOToTTI+7NEEQUR9QX/IZ1pdPXOuK/ldOQpF
PAX707hGDdX8VxKnm/3RRfm/oICyXzmhAS9Umo5iIvQq0on67GHLa7V7kIUFe2vH
bHfZWdgJIou4ps/4COxZlI8JS5xSIck3pYxgY7j/nR54IZPpbcjVogKp6DpD8/AI
mzrbalPVKLvZqfRnlMqaV+bn9pAGdXL8uWnXPIzVS0aW6MUyGn99ta0wQfOwWc4c
9bbZ38NzDXO/8nD1wcgdETqnKerNUSpn7agI6LZdj5W6eIolbZMDg+mN3ghNtG7F
xLG9HL/j0LFCkfl/cn4F1akuYd0zf+K5hnHc3RmtaFNMWtl9mvsp9TT0QyBeZTOS
w9SReuCGPHg2hIYu5r7dTh2L+sVfO3KVeUunvj/tZX7LavJ2FbVleNxSAQ0u5LcS
OBsVbTJ7SVI4qUQj+WhK2ysd5BV87BbncBOC3lLVEVCmIOdTp6hcymRSw00QgmBU
oxESJ876/yO+eZkcC8neQkQsKn2MdZvLa8cyjiybyiSOpatfkHNyZAUmfC13qJ5p
JdLv0cjRWLPFedfHvmMTEl/0MFnu60FUe8ToXY+3BL4mw+lhz3F9Hip78pCmRFBh
UOOUQ8UXDxJkOkshg04GrdgwuBgye9ZlWmBvciKW4W9SH4+z+zgRlVfaBediaSyR
oC2G3edZt/k+58nV7dZZKpAd6Xa5gidsWoJL1MnJ21LEaZrbLQOVxbf09lY5rKF7
AzM7gFlkGlt7ZlQOPHfPyANPiemWhluG+NxVKTsU0GAlo8WG+eyJ7IjyLzzaa9N+
J9D9j9examh/rWd7LNA/JFupQMsH3qaGbAx+R7aNCeGrmm4bT9CrOiWrVA6Lhmzg
fDoOFDk5llF+bMCKCoOnEBBb9dm24OHr9+CR5do+4JWdhgDvFxk7oarqvqnw4oeg
MjHSg+GkUIYJZJf6HcTJBm6XnwATawiNKOZR0+gG7zyYyqO5nZonFiEBBcQl5rAL
RUAjopXBgLO7rR4ajTJJSZ++liSweEgwf+JbMU5lXgN8R1Lse6AjP+4bSl8SxKnp
V0e9SJanJ5NGGQNOnVGbzbTGr09iClZUk1zN/g12zsdTUZr1rj+Uq3v0naxBkSg9
enl/uvSpJMxB2eZOuFOpF7/Oqq/fImDyklnw4Flny+FYbjsVvFZBzWMIN/mkvt/J
2InfYRxkx4gQVBRDz7ZgUpkZrMlqHhTioLRUpkijHKaxkZ0PcymOa8HRODk6r/um
Yuppesl23fper+5zxgNVzSt8pptSTt/J9A4cz8ENHYnDKQ7kQ+ASEozOtil9JKqx
bZMZ1mS64y4UMdDXD+0Hr/QbqzE4wXpYu6IxEc17ag3xOojWdmd8gbUmZjZ32UUD
A2Coj1Kh8RnxtYvB0vjZxmVQWGlEFv+T5Dp3VNDIPAcVLCNPRPuZt4t4Q/DYm7Rx
C+5qcOhAiFsJ1j9p7lHJsjk8j1pKHwKR6dYVS2i7iXrhOqNRCjrWKtyAvXnsmXpG
PruX86vPY41pSeuSpv613wNE1j1K0uj3wV6a4hUeG5gNBm5cglF5g3CwanVw+0Xn
NBCnCSut93zqtZQsHn6ZYM2QpcxuP9e2eJ/FPBnELifpZw0rdkBATkKz4Nvehs31
jEzlnzAWAmCpUd7mAfVkblnjHDrtTNrPY4t4f/4mgo1s/V/KQxbyxP6uaYKh4UtB
GqZ44XX8HvHuLnCbFWqwPC1a3Qg5g63Y+bI/N7jaceFyYW6Va56YQcXmcLcnRek1
lPQNULMS9luBVWSyAnl7MZYMb6OPKMPOvkEijZirceT+XBooCPvhQQUJRIiWK2VC
uZRNuQvIrgUQ7xzqWW9wFlMiB0uxpNDfz39Ep7ruxsxcBZedUwq5GPwY9SrgLlTr
zigYUibgkkCkZbbia4/QAJ0oEV7uWhbb0S9StfVlLazxIL3Rba6CEhw/2w/DHMdc
v2Hg/GztqHOLq/OBe+dlKsp/RHKaKPubWuieRl1iQF1pKN2G2xmqWFjTmaWrKFYe
BQMhicEyH4FivUkfPnlvY3Pjk/8RgaLeTP22TShjvsMKTFnP9gfStulnAi447xKS
/WIqT+Aj0HehlmeS2DBj+kdVLmCumMLySIDwhbzA2CJ+DvhfXS331bzQpKiOt3tE
kAHAqQcAe4bKP/Uy2XDrwhrWk99XkF1VrzbTaRd2lLCfVbpjInYNJFpwWaKSvRUS
DEJdk2VAzsWuyuxC5iaEun5uaf6QlVIQ0eQ1/aiDahhFXWlfcAKimhjn6nG+AXo1
yBqAbDUjV/m+BMSNcQobIVcANtpYnkKBmufUil4hWSMOZkHWctYKSYM5RSzPGJ3N
uo1OB50wZD2yLhUTXXEdv6SIlTMQ8gckc/usZ83whHKSBPiIDlAVM4TxJZOgeMGB
c9Pzz/bxig5RCpyiVow4YoKVPYaFnUe6Zjr7JXsry7JTxjg2oPeSaJftldHesvL8
lsRk+8lyxBuwGQHC2phsPIXVVQ0s5hvKIwgyFQi/IWYhF7Ub3Yx5gmVhtbuwy/kc
Hi+Zl5B9nk3W+OUK8EJqECLNzLoniTCOIQ/u9SEuKiXg5BVynWhPJpWeTG3vBWbZ
4yJ72uAO0SVicpX+gRR76qmgt8pQH9AMjdor69f0PygPd21rQtUiwcyUTjMNTgg8
T0Wz6urnDC03zu/D+nyjF9yk+wE/1GmyvxKHHumLf1pKNcoZciBnjrfy4lNEx7E8
lnh9cQ3fMpSg/AJV7IO0eHJEHJZdiMhPb3Z1+maWVE75pKS2vzJ1pjcw8xijkXUB
CxJXi96Zs07w+EUB0ZccKSNVcZY0bWo9mUdwiUmiGFSOaUwMhA29AmjPtHDgipfQ
eULP+IuvXqg1Plhvo2+vqWHQXZiMf5VSniqG6glKb3jlxVG4L5WOdRZBb7aaClOH
gC+xwPLfG/A3ryXiPrEw1XxdRX5ZL+uSrcmU3pil+7h/epUU32WsTCDht5LRlYpt
xuuPqAe0OwHdS3zJec3H441oEHidPE7lUxyk9QyGGr51LZexu2XfcbNtVuwUpAbH
ClPOq2JFSvAyNT1IWNh4x6RVnm53q98yZW9f7pAXyI94/QS4VxNeeU+XKH4Ttopn
WwXQkl0nGzYbM4y0nRil+sMehEmW2TJMVZPDS64y5R1vXTA4XuHrc6liw92oGa1U
wXbQBIB46OXbZqtCT+WYiJdWmWWatHo9dYo3pys1sCQ70CAzcnSWNwl6KOJxLDRm
e3M3XU+fgh7mYt0B1UdlxUDxNyrrW8jLdMWRQED2wr55FJQJuhE2oHZw6DBAap8R
ouLeoymDem/iVEUIimwdCT4g+ZjXo9ezgRCwTcjMtw6c2MHyfMORihsU3LNzvn7z
MPiOJyUDTZG0pSLfwPne4xFtGVLTKwrGM8v8JHny4UOP8OWejTA7dp/JIdlTy/7Y
YYdjYZF8/vtEu8/Kj6P5Bpmevnwq0mlC9/6og2c4IAhSTtzEN5a3M03kNcC78rDx
aaA1eyAYkdtKQFU5DZCS/Rfv+HDhqEfFV2HnkvIaR+jN6/z84a1Ilj1Xxl92udSI
Fu2whAZ/jeG5Sx6Gh7ECjoNQbe8MCnt8c9l7vRxEBSNTp3uF87+AZ9hY4GPiBIx3
QqL37CdyOfhxPwu2u+amS8Kz0qsg+P1nz8qVp/EyNmO84QlmgvQUraO4yyt+YqJ8
fqnTnuS9gy0izf11yrnoMh/XS0b8VFgKOyUOGG1/qcrNANsrRjW61/jJDM0N8K2C
gESPsUgIdYs549ShKu0rgcUmLFf6br02FPsmwjTZLabd/L6EfQR9g6M9+QL9ND4Q
9G7+cwsYrQIZpKp1XDROajDckpEpjWwzw9VSEKCwe5Z+iNIrdOBNqmAelvost063
SUzoHFqtliGJXCI9cTDMIFru83gUw8yZZ//f3aN4/6RWGkUlym6m4QJJA+no4r/2
iCkx0glGUAn6A+4l9liBmtob6c8r20zMg7/ViN/FTnyKQxdcuczG66sEoBPHwBPF
41BYfxRT1VJ6apOwwp3sl1sZLB2bPodz/JrxEpP6MUsjqxSjS0bZjDwzQPSIhOP8
2jwg8bIiQswm+4ScuNdjQKeyyaV7emfEjjfJddzVvPIi8W4yRWimbWPrHaO+g8v4
FTmckebHJPKpojsmSPWQqKSXTrYeFWwY3cvSArtV5LuGqBvYVQ6LF7YsWuSX/sH0
U3jL6a3FH6V4jqpbnaP/Yj7loUcMOJiVoN7peAwwbT/MmJelwrzToMM5YntnQXa2
At24tvL2O7VZUUbyI/Ofvte7brYMwY2QwulqIa+iZqfNWarUTkatBZjiGCOyIFuH
UPCOdYq4/ognUb9boico3r6IKbms4tjQIS/Yjvu0JMvUgIEh4s6JklOhZIeK2/rb
sMuv/v4I9MRX7dZiAKzQqH+APb7c5Kg573/f4aQUK25M02mM0od8mhpsxyR/nrou
iogEXJCu7AER/QJ1YedA4Ztr/v8C+/CQtOcGhc8Y5b/3rFlcRAcpWyE34pXIJd22
LcWH/MXmWZXJd1JYpHTG2DdONMlgNTVDqshjUpB/v1F9UXI2LcpUrAxWDWMqo2b1
p7kqRIJeZpzudaLkoKZFQ2iKL+Mz8gE7TGTw5BqiyaJB0J1LmO3SzY40gi5sSbmO
HwyFjI1dqISqyV3ogzOu9vQiSxMA5QvqNwCdsmTpRbatA2nu6LOuXU9Vbb0OKwfS
sB7GB7V2uN5FGdXdCdK7fnvu3G7LrBwoeucd+2UgaXyZfEIHKVZXEdLfQgCM/zml
+LHYsoMKLGN613UHZBv3OJ4KqWDyWcKvtEzixh2q8JTIvEP8plVkQexIDBiH16BY
rL+NzHIrRVx+eDzoPK8Nxb6S3+mGGw35CFyT2EROGzD/qNdwGyCFiClYPYx9sXbj
Au9WTzkQTgcHYqeltjvFpMyVrMDUVU/cxXP9Z7AguSWr7wHxxlETKicwmxhH3D3q
E5Nlj7iUZUaTwjqAgYYLYcGLmC50z0bPsHQMujgabYncxPgdtZA76AfTpcYhf35+
7VEbESdzOv+M7v9GH/EevT4fToUSqdY5japlulHAEE2yWNbzUXym6IQjNnnrzXz4
dRhxJj3nTV5L2DI2B/xrawP4UA7SbV+L8qQspUj42+aFXJefdZxtVL63pIOo6Qfj
bfxftAbNro2pUVLjw1OYS9aKovK3NFKUHX1vKjeVIW7y1aGZn6xYQcU+dPRrNlGx
WUnPEkvM3x59Gk/EXI2V+opE8574rxYMXtWF+y5xWe26HYBmI00OyaAWfXmn0nC7
Jf5asGNX+U8CbbICbCWbUWj3Gd0zbZm4KcHPmrRsbZy0X/dH+cBOCCtQoRUC1uA2
Hscbu2AndJrzfRa0Ovg2I1oqD7ngL+b0sLt60gQZU+cxt7z0D7lF0mhlPg1FZ5DO
1Wfi9/ttbPFFuzLQ8qQOL9TVFqcR0/Nh4tUaw8EFNiyzq4gFZ5zQMmNXDnF4X8ML
IalkHyqyd+JWZQSHlx9Z+rrCmyidmK4i1qm07mi82X/SyDICbZ02uDbVX9PVsoPx
RF7hhkxGIFNi1f4BBRUaQk0Kzx8vv0+gbY00aTcjgREbpB/zeUc4r00zoYRAbV7J
FL0QcvGP7U/xQyV6hoIfGE/qoQcQiGR4qVsiT8I5FYbnBg7mmN+b4ygw3VhlNFFW
aYIjRmpRV7+Z2klLEsf9/rmwnHBDwPbX83PHbnPaXlQYCH4xeOhvLyvB3OKY/ZOu
GaVcJoxE1VkURGNMnHifhSQzU52spK/xDU25oFhi1Jy1HanybxhR9zLQtwD3lBjU
nj42O7hOQjt/i7tdLy8vDmWii3KjNuAMAL6cU4j/EEICxzcWLlVZp7FpiHdgl2+Z
Cg4GpBx/25PNv+1fX4Z/YAa9i7sQ9DVfRs/HbBYnolTDRWD527qYVMg5BABxjmRn
F75/Wker/rkTuoEveMVsMvmao2MOsyxbgC0ey/BAw41NCwE4+eLTqiBsbrxMe3Lx
EeyJVmk2/RS4ThkGydYVs8yMWZ/ES4+kch7uQwC5t8QMiMV5DJ6Q5THXjZFUCvZd
J9Qtv0Z+bz3lK4NKEk4DP40YSUr5G/qwn9JFJhC5+6bHYblHUiHiDkI8YDcJ/RYe
pRSbZ65AFlXZOStium8Z/khcHVkjFKRn99019JxOx7gOTSDmBM5UmfN0XQIaQ1cF
SvnPJgBCIDXeNG+D8KIu+oqBKMbS3FbFEzdN/9HQ7Tfyw35Jobl7FBeNQoqKKYiz
ybGjaQt+Q019AjGWXp0keWceyLuQz/BYhmNsehqp3nljGu/0rP2acV48ZSHZaP4V
pMhvqr8upHYZnhcxibKnTnk3rLXbqQV2hw+2xWqzpMghKJjcH/7tnFJaC5X1IE5P
t4LIKq1qfWmPHnnwHKeU0IXci6d+5OyecxSwhKyq7RnAfSgdxCjzQEs5fhQ4ysyv
0w50XLpA5tlpszKFR3lrT6NbXG2K/UADyhiQlwieOQSFLjcuyZxsueqJsCc33jIM
T5pCfS0E/0WKpbuAepFBg19gmxvN5ZV8cHEP+16i5VKHQsKLdsqo/V03wrJ30tNq
o8Ofv3BaIo80TWcqxtuY/UJ01YXZo2ZXy9Sn4SpW2mr5uMsUneSO8xZPt0FiwmWq
bIDL3s5aFYbqY4dRoZucIDKBDgXwP2b/2oUfhMz0SEJqSd8USt7QJ+5tCeibAMsY
D+K2HtnIB0GlO0jLJeN/MRFuQKP1NAOWxmhpMNfm74+/yZ5VDBj9UAGOjgdnCRnM
hNN0AJRU2mr4SfpvSUlrih+pIYtW3sC/T8nF5CdjfRylyvPietVzJl3DBjwvwF9A
EyH892YhVrjzCUBCiXHWfsrI0U+iEAvcb3QDWtPuf8EstFoeWC4eMM8A0cZoN+n8
NlYJtjlYCcNStYTrsS0AthNgGl13iReTvkB4D7bNqzc2S17cWRO1I+2XJKyZCiEK
qgBjX4Jdja5Ubiwk5HGXP7wq+sIJz7Xo0lnyGNIPYtmGRcFeSB1q1D4rP1uj9wg4
ug45lJmaBcu2Zc1LXP5Wy48L3L/SSUjn6WmPwYLZW5CNRV+fO7imcR2ivBOe3yCC
UpU6Qv3/SX4YVJ8mM2qjibEbQus8G3IsIObZtRqMjYt+KpudFg9aqEuqfLXnNT05
NWe9ELOD/5fxp4qww+KnxvP8e7YVtn1zTRLXSSnqTL+NrFoigw1LozptU1vB+1zg
5t4sPHMX6VTgTPMg2No6EhnmTGBSojEITEt+Lxu/MUTSe5ATPWUrPw3usKqY9ofO
qEYBAfZLM+BgJGKQiE+z+NeTWnYHqZ2kGokVG4ionS47wLyAkw5ABywmx6cTctTj
zChdLLRHWVbI4cXmi30Z62YzsSRt4ibjRgBjZ7oY+ZMxDDYf84SnT9qJ0l/lrwta
cPo9OQ1wtPwsgpdtdAUbfbw7pDkLxWLgM0z43hz718T/e2+GWBE0ZzMVtHDTIjcV
yHJE6TDLVHvVXuVxayigbTJR1W546z80WsnBWHenVPxtObH79H37JJdtCNW8yp3d
eG3jx7Z7mAxjGq6DdVja6zpXVVQBACCLIyoryAiOzuh5qj/OTS3d7h8UXSSJSNQ8
JX5mpVaoTxIdIv7kKemFob8qLf8mwZy2F/L9Ph7BE6sbRsOb5kSf3hDxwLAELPLS
o9EWNyZn6EbMZvihjNb9jKOVwB8ottHtqEMH2PjIoDlqhNyaLRGJIQKR1n/S7ED/
l7oeRqccssS7JRm64s2a/etSuaO/2w+RmFATIhPJQSrH0gknDh2Lp4KBNr310nl2
OQCzr4IcSvH2P3+R7Bwe+RhrFIo6BwB6p8KZOWXxMuGN5bwEAA0JmumRUTBD5znp
2awhR9P1MRrc2Re7hE5rY4orUW7IxzE4Djqr7Vm7d4yhC/L8oilSqeZ/ZGFcLpUg
JiZP+1Bq2YpJwi9sMcU6AFpDh6INqp8+8ADVvXhr/r5vgMDGJx6pIvd6uXZIUUXO
jI0hWYhkNeAoWn5vdHAmYX5GJCldJ6O0J+vZzg7qqQuDM+HMHep0Ifcw02VEzwxO
XM3cEkKy4lQzsmHU49+mhDX403a5wg1K1Hr9oGEYtjToEHBs8XKarkg02gLi4/VS
TKB7RWP8iWNrNU6MwCNn7LTSKUPIaCslOlJjYlhmSWG6UsV9T+VGrr3SG9yA7/Vo
Z/g5a2LqXfcAsUaMuIMFwy7kr8FDRQ4PKKbdB19glhMMHuP1g/zDVHJEyWOtnmxC
xD5ObcIYcDKeqh9JS48/ZAnxTol2SZob6UFNq3Hpmw3ZQc76UeNq1pNeeZupa3W/
cwauzPy2MIqmD8UFHKwmOVMUWvtpoknbSowDlP9rM60m0HVtaIRUZ0VtzewMeZFl
x2d8fR/VvrzRsN5hwjyqsmrcfBCQCKS2mPCxPwIwghVAYSljk06vNmSZ8dOxusMU
e6NNVDNkfceuX5oQMS3PghITxJ7+J8ROzBFxifx2FWCnRICydJzDtjY5UzRqS3Oh
ZdPTIkhWiE8J1XPkPh94c7WQXOOTzhHOK4WpfdQNS1kJk1ra5khd691+36rUEUMd
t69NReBLwwYsCvH9h2qgCoGPRZ6ENwnoYOfLo8+hrahjWbo0o46fp/o4PWSgNgVX
2oYZ00D5X8C6PU8etujoIx+UyW1b0AU5eAqmQeOsgA/8W4ehiCJiZONuhJ7t35IA
c7r46fW5xZDIHCkoZGs4SVdLKR+8tQiUBPCSdAo71PMTcmUXDB1/2nouewPVgEk7
knd4+PeggYi4KDTIum5E7VbR36B16+10rAt3C5C6IGwH2GSE3sFa1sgsb5yzIMU3
tAXYUCfKprO74oDE4T01K7CbCUJriv/dKuBmXc8KIfn9yXZr91I+IiU6aWs0WEtv
2N1sDZI5IxW0TzsSKGVOIjFsn1V5IW8u7kioYY75FoFCo5k/Djuq9wjo5qFeiXpE
OFmQLqNof/ujbYorokuDVk2lkBKLey2jwyErX8ak9L1/h3YWQqLINVZ1YhVqa+VU
7kRy5+Pq6mw4y+bWVUx1ljXKIkN1fnSwfYzHN3GPvfBhQNx3OsbC7R/DrgDqIQ3w
xtrGFzKcz5zhuD9OTEY6iO/UsiQG1Hggv1y9MlaG+9UqMOXSJ5DSijCw1I0VXR/o
8ARz6aeXgJ6HENdEu2CjuR3HXZ/EMF/0GP8tLhdhVD5LVrwxLav87ndLlutilBy6
GFw+WQaxBL26x3ewuINLVBGTk6FxRklkjAcfLuha6JhcV91zbDgYr/MY+OdmnPci
tEUYS6n6WNVJYV5B2XrW+SU2YA2VPNgxWmB0vOU4+k7i/cxEDTlUf0HT1jhtYuTV
RnY+h+Oh76crOjqIz0LuWgFvQhQdFUwJ8/PGELyaPsdPDuBG5HeqsridHwjGQ6u4
JxSlgv00uU8sYwV7rYWjhgIdvQoWXihwTQEbnWHQwxZmkk6M+SMJ1CwFQOuzj53A
8Xu9EnimdSHmLEfxSItsNPFXY4EhoM/0U9i7T7GFy/SpRgttvZ6T7li6VmbnNfoA
qqJWZcMpK+vmwM6SX1omFsmBHRL5Yb/5EstaRlrhfM9PvbJPheFp0uI4oMv8CqY0
PAPCRLYAX6bmYQ+Y5EBKQ36AC0rLo1uHlQaxyX/dc9xoEAgczh+vruikSy6mFpFU
Wno0goOXPiVk0cQw0u40kuGIz3H/nlHlCRXmsFDnL8Qhbxe4Lh9hiEV2KNb3vFMy
rnOiVZxcnOaaeB663Yjpj1EnxIMXFABvpdz2g4wezdhbv0rM4KbSvDJKAtWqkwqA
wWGAvJkDhp/72Qmh02P5SrDq6j/iIBVhY1BrVWBGTVLzB/iG1g5fTlkr/EkxuDIL
HpwoF6UHljot0BrGtC08RywqsG7agop1gtIV/pD58z9VEo0FEeRmiee1ynRvngu2
ALvEia4SpgTpoTqTvKs7N3jmvWl+K0u+65hRcMr1YhnnUHvw2XOaJWOhjMy/Kdqz
65dU8juvEfu1JRnNop9/jTqlfZUtfk0zRB6IstPVmVEuBQ0xRlfs9lpSCI/lEuWy
GrE/vxM7V/nVutNV5qS1nbbh83H/OU2pGAdTfEBCrmWetkg55zxV5ltGVyN44m3b
+ML2jRMoqcsXyEeGmSxugNIiZKeTlXAPHWAx2Fcm55Y/CD/vunclxtYO8flCV3lE
qMKt0iep9uYfjJrE1s3mwpe97zi8sV+WPubsq5mXIYOTnTReQ+tqCus0roAuJG7V
jzVDpEUK7/R1TY56JP3rp5EFChBm4v/G19zPA+eGiD5KJzxcaPKgVwkcrtgtlD5X
3EnBzNd6pdEA3TkktEZZV5hM+aVBJZ7O6nC0AzWJpu/I/5DuBfMFg8Qo+4kpoYgr
rV65jFUfFah9Ng51z/zmd3H0A0P/vSYBT6w/XWHSelHYSHe6vAZ60YfBAbkN2ETZ
fCGQ0vLOki5woL28mnUh5HmbgqcrjLkY3xCTajLt1s0ysLlUt+xmgwnz6ETCoK3I
qEizDlPKcIcwjNHJbDymbyAKVq6fSJjfQ1VeGZ72aGikXBTYkZqYAn9TEcOpZb7e
oJqCpuKqjXioxaDejIWLkDBCDbBY+IT86xxVvaE1uu4V1k8JySbyganuDi6i9RbJ
iK2AQXLJwD1kv9pS+2adR4iXh3svETwsFXxj3YBxlF2VfjuF0qVfnW9mIOmZmgQN
PIvTeTn5aGTJUdlnSYieTWl8GZOmAfE4n4z+o8A84gpFuwqt+6KfO1TnRCZlN2nz
Xu8I7C8KL+p3XGp7WXh6hxHgp5/pZyJ9S/7G8Dz3tNjvdsr9LR4ONfYH340reriW
9KICNKTGuxgO/4p006/u+0rJy++qpEfkMowlJnJmGNAavgwhMha8mVM6kSFYOIm8
xgRtMH9zpOtuSnTSoDVTr4HZOhW7mtG5ozrCyegRyWvH/QkxzivdI0bIB7Jgl/Cd
Mn+yC8XqKgcvqf+Q48tmMk40afdMarTrPKJrxbVjmweN8rmubRKejg66Az1CdO0U
5rJMWNhYwRlAar+Bjot++UCUOvnGyiYAQuhEYsfcETHlSNrkOqazxPfGvUY2A34Q
rjM3NnXAVl67pUF0OADtWZp4LGrozID0L3w84OxCxOdp7EUwEfpS+uwI3NR8fYCH
KjD8wwlR7qZbtpJoMVKPPuFxhLC0T+dchSVj3slpuL3+jCgC4QI1b4BGujHTx0vm
oBdb3zr12zUFOS5LxowkmPAZ6tmtIZ4JAnWcAZZqAeO06pG8s+0EE4izLfBoIE1s
w4KN1CXFp19NKaZeMN34vyAHEBl/JQiTojnJK4Qf31VtEOVFALSN/uC3dSTv4BE/
pbMLFmTbC+SIpNiULPmE+hfpqFXz44XajAyLP5+/sGj+L9FuBcwC1HqMTd70vor0
5h8S3rZY6RASsdOeRdOmcWXFQTdPboim9Rcog6QD/4OBnqJcfmtuSY/ugCmUzx90
QEltQoD6vfkn/xa+r6ptpYZ/HJ1mAzaJ3yezefDZX5E8Xgi0Fdf3TSnao1eSc6rq
BJR//awcb4cr/ywj2KAuLyijORu9zRgrc8cWwPca4Syl4uQiHc1W2UAunFr9bA8f
Apbo3sCe8Yg36Cc1jYcVK1SnrDR63RoqYJaNPQ6N2bIVYOpXa0CgoP+geeQ+3Ffe
qCAsczwjBkLUdeN/JSHZLTkQi490RrAOoloEk5W6DpQkKrvsqpbo16c2tDRYUc8c
Mj0MG3HYiDrmt3ZkPyrPKSUKGtamEjL2FDzIa4T4ab0PVTU6K/jA5lPDauhGFv4V
I4g2RODvQq6MUMhpM7pjRGDpe2Z+jHfbYthUgv0r9qUg6pKjR1SFKfKuhs3c17ub
xS7PJnv5jMuOt1wLhtIBuz0CpfceAD5FHdxkL/3nwN8CtECy5EVzM6Rm0W2/N+g5
udhSfDX/kZDWNIIwAQKh3DYSxX2AvUpF4qvHwL9+Gb3HYVQOd5Bw/j+HSC0CO57a
TLQ5fkT8RWjM1ii5+LMWO8l98iFIP/Plt2vKZaW2a0EGS9nuLqf88hKXI4aR9EdL
j9knH4HIwUK7oxbs6dfmcPaRiokyen4XMo/wbeGBjRLOp55+ixmasjbfdlmO3xNk
ZOWvQmdcvvEHPeg8ch0B7izOEaecyxLVlJucTpfAL7dPICswTOapWkKFQ2kvx2Xd
tRteMgugnEmopUI3guNGExWlcQpIljqGQr+M03IpxhnqHtJ0vjcXCJLInGUssSey
TeeLbohEfgmcLGCkb1x2sHwh+kGhZ058IfVTYqlpbRPHTd+YgXTS3+05tfMvCbc2
NKuYOZn5Nv9JxUUkQSOL8ZYlOwWxWmffGo7Hpsz7lEj/gPtMFe/yJapqtjvnLlQm
GTII4eKTv6E7vYviBtO8cLw1VBX6n9LSrRuIR+o1D7EqitO6B63XodG70rSYG+O9
RJV4DU2EJKXt21S0D2Cs/ukCtMc6NznN4GYJTppQaMaRw1nVcDt3AX+sYIf4uQXs
qW81XHZn7r1x5ZSkhYjoe01XmiSpu24G8XZxiOeKqrstAj/HgDxeuk7VulmGEWmx
9sCm3KvAZP7asFBWj3otdCJrDCaNLSgCbf3c5/6lj0HkNwOs/ASxd8/yeFbgNltm
yN2t748sK5B3fDJ8fTcCAMuWm51riu/AC6aPT4Fu4hSVI1HUPMrhTJkP+jF3JLd/
Lf0CXr2Ow1zFZTvO/6tRr/6rn9mEHzG0CWQlHr5YI/zysQnjVqXyDijpzxQ2THXE
wQorI5TsymwE1UF4Jf0TRGj2STRXrmhA6qMA3TE7QOj1IkpCOrZrIDcWtI66QilH
NIxRS2FvVlyv3+l64U0mZzbjx40GR1AxIev6ra7kBMePV3nPK52dFHll9fq4Uykl
nZPe9WF6iuXflm9QhtK3OYX5YBBl+CeSFduor0zMXTG3Kxx3S7/5RGkTT1GZbG/w
LUen7Qk79jVUovzsXzIe8TtxFA+viL8NnG8Z8xtyCnpMewRSzUqwsZvWAVxHQifa
K675geuyCQYICjKZ3eatu0qpUFjbgwUjHACkZ6zePUBtZ/uVqmgoq8wUvm3i4GHP
XMrtviFRvdObuSgoh8TCtwb9QFUPM4pQ7xNqX5vgT8DLSwiGRvnEP7OZO4fFCF1S
z5CNbX5SPyHqxt3wK6Z2+4WcBB5nALleFXDdagIWHL4Q82ktGUUFIzhLklCrsKpt
d2+ai3eT4NA1RLpEEqeOco3y2wwexLh/KK0PdHt4v7nMfYevuCOwpm8Wrtd31IeI
IWMOO2fWP2AcMVCWtO6ch5AdwX3j1FVMx0RSNDflTKAyP+6Fu3JelK6dp+q9mlHc
vZAfb/ca27wMInipHH4V+c+Lc6pzlgFFnxjFq+Nx4QQ32VhY/XWdeK06G0s0hcBf
Y7z2wpy+IftmBnztQxWuLWV3gH2K1AFF3UBSl/7CFnp0QXT8TOlJztdsFhcD/kmy
INroWYuw9wC5vYvr5ccgiboYdMcYAATU5/TX6fZsnFCySLUvywAWL1l2UNtF3FSK
JNI6VDCuAgqZD1cXU+FhWEVShgkG7zfeHlz5i5jac5/jQltKZAEBdqWcD9/5ET/w
PQKzm/y8AMHX3RxM+R6p3Uij4gfkTuxc+oRFH1F6kwcoMx5AnXh1IwWXVhqpu8tf
txPnSQnsJfaFQNJlPD4yO4PBIKudq0g9q1ygs/Rm6Ep4QXeyvnRVjt0AMtTJnnFa
47cOnonYBN6PxRwt3JyLFAKClRgH2XKULpzCmXVPUOTQrshMidp31ySkoyGN+VvR
GL+DW0PotUmCGZ3/EWAAnIQTWSQEWrslzbe41RmdIiP6/kDIPR1RuoPKdBVNQDVM
hdGH+82IIs7HaAQqgJftP72RHTk+x/TZUVk4aH8sUAsJB5Spj4xuuzDAVAeabyi6
6iEswMib5GIhKzOSjB8nekkBD3MqOs0HCvbH5kSGKPIpwqoh2x8Gk+G+TblM/JID
t7fZvR2Td8uEFduWO8n+vqTHCKqCA4ydOAkNua6AEqNogYx3eu7Tw3eGDSDa/ezp
9zCmfWPTe/ZPzZ4+Lc+/NegFY3TJqGZoEouyjpd9cwYNZH5L5wxw5uQV5uMFcXAy
gBWMcbe6ApdCBIn5dZqkuKUHmw13v0LpkmLcmOKyuGPXAnPKYTTedswHEeuBHGP8
Bi6KmwbnZQC82LZ0TBUl7zWhlgUkVM8hUT5N9TOkkZAAp0xtQopcCMQ7PGGalPyC
J3nNeDQ50HWQIptnl64hN3OEFeEU5iUZ3PgncAH2+wzrytSKFpqSlzssPtNlopYx
UBoD/N863PKioqFaR7mXIpAsu7MsRAxV99DRWmVdfpGYm0ZEIaxX/IXl1jtixzEZ
USzsggj80uWhLt+nQo7rlxEe2sUEsj2A+e3suqD/k/uxrGJvpADiMpN6xZ3ZZhz3
3Z6/wkbE4LsbzojotGfewzxP3BKuOR2cCT38NoscwphjKOoGEoABLFdyiJP/1FiH
/Xc+VaymViL/MZkDjsd4YUMuHNXFe5xtWGjbvpPtXJAIz395XaT/eLPu7wQgfqwE
4DACvKUKVunPthzCPwjhYo49xHp1qCckM7ro8f78VUwI/J8gnZAa488WI+QsKvu7
zw5aeOoCl7dpskmi3g/NW50g7Cv0Pm6CedlTuWvcBvkGg9YOcMSOqbpr/ttjIwtS
VfmFOs/cK/P4dZTSZ8ZCgB2gQ/uk+1eWK/XKFOY/0rUvfg3UxT0849z2tVgts79g
pTo0tEFGo0FAlrZAjUvw+CCBeCPih9r78Dkr2n/7AWLSVET7aa4J0efpaxvV5rBV
vLTVdtehhepsjtWoZls83+U6G1sUoNofCtFEE1Uk3Bdg0kB2CgbtbnFHFcMKhRUk
BjVoUpv+YTPAvPFTq9UnfXjRewMvkKwlVriobL/IimZnLsIZQndo+vT9BgoQY4rp
tHPdO2cU/nLRyvFq1dHX5kBeVzaZrGnEj8CfzP0Wtwp6WTzV697i8pZsa5Cs5Gfu
8FujQr8uQjieugBZYt0/krchesFg68uJv/GyydaVbGaPdFXrheQD7uJbQ9fWZS4r
/z3i7k34Nvk7KNuAjg2oLeJzLwcO0tVfp2OPW0iqjtIGxvcCPZWGsSmfVUW6q1DD
apUlFw8B1JTOKQAXJICHYTlaH9BeMimpGpHjsWYnE/vcuXvTwcVBgtw+RhHdX+Vl
rNXnNUPrOhXG6hmTWhClyAajUsFtOLI7MWgVDbApS60BdlMjie2gbzmc9kRPQrdr
rLFi9tS8xqlRerbJS15n4xzJaG2P8esZZevwX8I10N0rh/ny8rcU1U31GpLVDeL7
WWSo/pHmhHnomhQZ3KcZDGT/eZEsFtXSXnShfRI3ZSauXhTGYtfxZS1Zg4F5uuNI
RtpauVPZcVmnkfUU0I0ENP6ERJsFlhC8VAfPYLrKjZXjhH0EaZyTGtgzVyaEVkX7
JnWyfqHMILNugGjOvjx8qsLav4pwHxam+8VVB6JTFYEjU1ysmwQ58rQ1bEVXyVlB
BPUEKjMbESas3Z+Up7Yz0mEp8GMSSU2S/NFOKaZzXLbkZ06cPx97p1VCqASF6ckE
+wxcUTTZtW3rSWhHUKH7qMohFmI0VM7v5Rz90y6WV31YaPAoBK3pob2DKxKJ143y
XUBV+mokZdWcUzkrKx6DaoYizUZwIcQuKQa13EjWXV5e5ICBkg5+aZtQRWY8R79o
4iAbn0veAvEGoXw/f2+9rx4i+0lw4Owu7SJB/Uwcs4r658VVNd71tAPwRmuwSSE7
ePyDO4sNNR+2JTaA1K68jNZBrmAcOnQKyNkTONtA5zxeToOyOhH/Z9Zb6a4x0Mg8
8s4ZUKrupDdFdwFxK4/bxLfva81bND20znNhpGM/h2uNJSIiGL8IZ5rufdVdfFTD
AIPrQZlpwBbTH85r/LbWDouJY7slHDEkOsY6P3zg4rusAv5jzQX2w1Yby1zt02GR
b5YsPlC/GyPrF6Cb0ol00FZsFUB9lF+2yf92guXi0kTJ7DtH4ucg6yqk3EO1KzsB
/Db2GmTB6BXmyd2q1CO9apdJsCsjmAr10E5nvbj/L/cst1MuQHoFNz6F5eCNvRar
caFRV0LHM3ibbsTJ5Zbh8hhdogbYVezCybpaMo03HzqZgAiUxh2oYmMfYkFVBNTP
MVx2oouPaQJU9iKS2ia9S/1u1lM4KZ7J2jhUvfdJ6auNox1/ouUkFkB/EPQPPx4H
5HVxsHvuzivqnCS6VVbtw7oKdvulC0Qe3sStJGls0/4WsuvPIZEDZjrHY7dtlSw8
Y31LXu/35F3uSoieXjQ06ba0xf9xDnS2d695NfEpgEUObDQBGTu9HBliMwh0JapO
FiB356g/4sImsH2Nf15/C6PaNNT2zXfZqqYNrPnA+6oYt5Zvc9rOZQ8eTdUzupTQ
Qj5S7z8d6TV7Ah9j6YCLX0rZP3b6yLBHEz7+8B2RVe74dA44u0WTRaA3kdHMP2lM
vtlqntZZBtj5SbIBrftmVsfzALQnH5bEuJpxi9d6EWYnFqdjtHEQS/vT3m3wpYXN
Z0Yw62pGeadkg1OzaquRsc99YSowmb5gH2YrHEGq2cJT0MigZjIuCzjVt37xuwhG
+3/VAP7DpoW6fR1yqCtvgqUgPCB3Twn6Jp9D782n1zyAT+ZpCo2BCcgTp+uq0Qud
J0CZaywMnxQn51IlYrq/LmOfk8noeDbXkP3RutN0dHUY+uN1dvucpUXo4vxkeLLW
bQIHAKzIof30xvtt/yPX9l1Ilew8P1O0dospJUbfwNnYT8olnRmex+pyjQyPhFe4
/LFC2FdZ9x+cT3RjLwHkAiysQjNkD66BH3l9T+j+ozp4q2GAnrvf9mLIWpoVhR+W
m2RJqsjgqxU6FG9FOpZtZTvwtL0A7LHO8Si0j5UTKU1yV417JrcXpjSR+fGD1tYV
AQGhXtZDjVucZN0XLMLUKyBMHh7jZ8naoXyG8vi0ZPzD17NhANEPuoYHFJvOqokE
++TBp5J86GdKfBZa+OEPS5v2GXxtj78/87OMEKK08mXEJBL9xAV5y/UEQe28dgv3
dOPIG+pXAiiM7UQJoNjPdOrgN42gKBg2fDrzTIzQcBw4cnYjsTZ+S7Kez32rMT1Y
2yT0hC5uHPm+jC5JBidzinOg1opro0Pf+mndZdCluhMpoB9s/YeHMoQL2LadgT7O
FETCXXH5uA3AzXghxr593lYZn5RPJqdV8/fBAr05cQHt/gm3kutsQ/7tYcRnAQ9D
C2XUkHC3sk8h3mjlcfVLSbmuyEc+rrijOQhQGk2uaX7mPRgZJj1otB370dHtwrym
zt3ZTNggivPGiE47F4+WZl9k7PZV+sQnWyVmzzaHSnwU64SvXgSDMWesR9qu01fJ
46o1wj+0u/hrGnfrnSv56vJ75011pGjP1akVlH2Lz2RUAPG9klAyNE9yGO9fWuQ4
yFizqRH0TiV39VIzWZvw76Iask0QVE1ZbsTzjres3g+kC0Zl8/jXENQizcXIRHfL
0r2oqUWpniqzELCUk3OiRRAIIkKFAL4etnlU6VCtTmwxUq1bVWwycr9Asj4UCVkl
mecItjuxYbHUViapoqTa9UnDji+0KpQin5930z/oFLMV6Rp+s3fC+1DXvhQ63Yds
2uAwizJ1T3Fst20V+WMahaAOjyx36obEzjWwGOM7OkoeWZTBbrB9nQvF/IP3epCy
I6mwAew2DCQtgnadFcDBhGk+UAEI/pi5CnFlwF1aNLcrT7TPRVlFo19GNLScCXEK
QLtDo6atfxU7RhcSiSmS/gXAfz0+U0TT7pKfiNpgtbQkVLpHVESeiu2ckTLH3/AH
UngB/B6DrNrXmdLJK0s680SVRnLFCBaCktJkYeA9KQUPy0TEA2XUZQ5vvLVzbFht
/usITtFXUdzsuFxP55V9IcO7Moi/6XfKsQV8MlbyKnMR9oa7lAo32y1d34Is7CV2
cIFAbS5xRxul8jrRpglQK4G/hIY3gT3Rg+IrZBy7nTWUxfZfgRzTJRMJNz+1S3vd
pLgo/Y6Cdo0AuOPi2DMtqvIJWo2PMMDLET7u3qyeXhWM+F73OBENLBAm9V8VZq83
tutUKabzjTDd5YyIafL4OV2Cgt1A3OHK8xfRDwnF8GCe64bSwhNhAmwo7cY9H5gm
P8YQ0Je4xTdg916p5tQ3V85pyx4ziN/o4jxItAZWakBMW1ovo2/FUnmHE08FiYxD
suWayGKEwE96ADGqAF4eoBDWkfbT2iN8O+QDVQN54sFwYoWv+1wNL7cmkBnGlDhi
j4PyAZYXxhkZItCNIDAwEcS1fmoioBcR3gqH20KNZhqDGvtsDMsIQfgdNdXvZ3XD
LeLJEkCncSxO1jhrZt3oPkbhQZ4V2P9CZkGdCoC60Pol+xQ5r8cl5R8MxvfR/9wl
xt8I4tQjx2tMw+pzAYheMrEh4W+QAIESGR6LPbA/ljF/zShWZE22bX60G6nNX8z6
37db3F3aE5NXwJNaXUH0+LmzUVQvlZlcgNDsz5a1EQf9pIr0opgg9xDgHWyjNs3M
AmTiGnU8gYNCTc1hOvaJttqJT1hq6KzjmW+/GCiMoqNClh+g7WVfVAZrHBGEYUsy
ng/nPL1W656stc4DzP0KnrIZAPVAGAWxzqx+uxVvzVVuhMRzsfCnZmjbF7S0rmw5
pGlDnOOHdTT/4fJ92BPlZBVTTRf6KzS8p5jlfPzTSy4O8VehoCQ5eQHXMb/avyzS
uqJEy8a1ol3T4BqQPKdC/ftbZ0rOjKeyDV5HjO64xznZkZlSdtnXd5MAdCU3Ulj2
hTFMtJCJht/5ZXYhw/ewfY2FVtMC0+2kX6Hk4FOxoZHMgmnB7U39dwS7jvxgqNlS
Q0Kxl6uVFUaWrlqKw/ggvpPzSmgRkeO9bvQrJ9dhswNDAIG1Jp6DNPUdrEprg48t
lnuU7FkPY47D5opZoebTkOEcCKkVymfSLbqny6VBnVUrXD1SomShL6zZRtTM7ymr
DlamZ/4l0n/mdP5jMXB6fSv1sZLh9wCtjUO9VyMDLiO3EvDhBXfjdoGn6BiQLT7T
5BB2AKP0lTMszr8Q1rpUk0tyoTQ97+u3bXCLnZT6DffQdrv5UWYi2A2L92O2xSCa
m23rs1ua2bXVd9XOmdzIKHq27lCT2+t3KXsQRFEWvb9UdD1Lxu5Yan7ow0lLyUtj
YBSkLCBSWMq5rBY5E1yDBAfrG4KPY4L/KboxXvEtz90GrBdrYC9xdyYsuhQUUqge
7XHMdQ03kfeYC7/aH8CIYzCiDVQQd3F7wACA40aiZraW2ek29M/sMxomNGg0CkdI
UOfu6l/aW6IzJ9+t3v7Pyo/pkoG253zE5ISn0m04ZSU3oWSdLWqlnD+WBsANyC4z
Xo8bwj3iYYqxr8PcMkPi/FVT33oa1LTQRLJ1zJ5f/AG9kPxcN3b2maA/huFKm4Dh
BecANYyNuYgjeGnhts3CMAF+ctNhlr28Bf4OhrekDTI/xx/i6K2DC9dUlgR8G+gr
qVRGeTgYFc0hpQcvsvVy+BiYwldKX7Awepfbp0m3brwG4ZtUM0cEFG1i2+8d2Own
57z9XzgP0Sdbl8s2zEtgNo5jd4JmM4+APNPW0GGKH6OQaL0ikU+6ujdWEitAOBJX
NQXKAOQECai/FxMowkjhY3MlUMdITN+VBG2dFZVtQTwXc9DzPQDUM/4JrM6/4M1M
kzxi62tnVHgLPiHgDZRjezKFu36GF6YpTftefUJKxtvfIl3MPXTv7CP77LZGwdlb
y+HRKOnuiiKlZ8Q2hcZPmrXfm/sjYCWWg8ABMnim0hHekQiwb6AYxOwLoFNk3oPK
hpUCfEWBAD4++uvXznWTvklVUScVjj6dyxohSLj9CuEygXclf7yVh5YOjWU5KCoo
se7GKZyeouGafMiQ19AEpnNqu0jm9q72ZpCrVdllTtBqHXeSN6TKi+j/D1SZrAhC
ulGIleGjFP4KbfQCNhSsDH63J237A7CCraCwm6p9lDRGWWREHLfxe+/zRI+FSa7h
vq59PkC44Iylq9rTZboGqa1PcATH9plsz+kYVctB0AgXvXBemXVIQb4oeiL7kfI5
Hx9ygvXPt65z86LNkmuLogPtM3XlPVIxJv9gndNaFcZs0U7hacTeUJogvmyGr8uP
115qzvBsEKJg9XGMfmasvycjxiRbOpwvFsg41LHi5J9F2C4hZFuNUS+Eddy+VDeX
QM26K/xWNpXOElWg2j8YdCEpTnYhKPyUNumACNJbtvJkQ0JdgemczQZLJVSTGuQZ
cdkN1cKdrc9ii9BVcrRMshvDMTly9h+xMMr4ZfWzueIKrymgDkr0bobUk4sP2C5P
rPIdvyrobwH2/hASBuhCyN0zYqON7fBsHIzXCX1DjeoEm1v0C1QFQCu5jcxFKS8n
n6KdUPH01zrLBYifgz3DCzg52otb8J9MBEP2gGTaE99TMVLMOX6T/Fjz2IA/Ekzr
chhhdFWmcj/JXJdij6pyjrE72GNlupWsE1NWjme7JP1mm4GZ2smDohRQKlVmxhi7
XwtD4HdNj0aA4i16oiAjJ6BIEYfAglVFi/xIumdM25fItLBVQPwZIDzRnGAvbhXA
VgdVkgjspLYxhjukV7SBTIKp1USw459bFz6nctQbDvzjh2SkMGPaigH2vaLMbjVF
hAIvsgAgF8c3hfF0D9KWhuxKz+v7TkqC4GpKTrjwGBpqfDobmh4AJKONjqo4kdEh
GXnmIBMLay2Jdjy4EFSLWWk+oRKofBsYkUtDBIeBt97wrtjifpL7eMcKuZQDu/iq
8fa4e7/3q15oi9DdBUaiiQZugnc9ehKAEeg8KHMfPQyYGbfiZTPhzPWq6+Jtz1JY
JDkXUPJHm5qbqkrL4N/42/FKa64afNyNfMa8JfJr1JfQMtebGWdvGxHZUUVkHzGS
3w7ZQbwwgMaDz2QFjla7nQECTwh5hpfe+HIhuuYXOWVf8+pgA3Qx6o7RDN2cdNHk
DWOfLYu/DuLRR6dUcp1H4ea7S3B3OLVW6SC30lkYMztnrp1E27UbH0lDM+LqXbml
YfaxrdpjYnRR46ehl4ZMApHK0GBDyot1PYbdWaYIwrkWo0LJcTq80Zl+0tLzoj3t
Le1dg0+ozs1ZOwenVeO6T4Rckacv5Sch4hBEibQTNRNyf7NHAqsTEnT+ygWw3hcq
q9MSISStRjRYyZAOPooazEwdhYAVpnGKXyGnUViR+X/+4EPiDDXfKHfeOKeDCn4s
LN+cYFQligRDiI1TQP4bKN+lC4WAQm0Cm3yaDuPJ/4PkfBH7SKW0CruAsjQGkW+o
hx3YpzdF9rvTZ6c2MOhetc4llL4aAvJeGv0ok0vpOh35bEgLTlOKXIZgAAT6n8QW
Ab2/fKF6PaWitkvOZRmC5Y4oaLxkESts18mkqwcerKbiYae1xZpo4qAVDeXj69Li
XeNDarVu0KoFQPZgvQ8I/3Hvku2tttjPCg0wmWPOdZonkNQK2GJDqUNnXVDCXrfB
jXWWzb5/6NpPr7ZRkPMY4a7UoxCunh5TdBQO/9Eyh154XKOdNTRZe7YFIS6aQNWl
yvmHTrt1E++mAcyI8kDmcOD1eAvkzCsF43ONmxVgGlbO/w4P1YfbLJdDmvbfyjQX
nAdSdSfehOKexMsTue1XTGodzmLLdfmmhEILAlv4RcrXsoOky0BoMtbA45QytCQz
r87jX4PgRxjQ2xu6yz0NoYNgcXTC0laP0f9XzQYP/pOTd2m7i4PlyaXAEWd4wucK
dIZIyUsZyR7U5kLhfzZ3orQEMQNAY9CQbXnq7dOXBNzgiBm0C5a1s79JQefRfjnq
3QCeGqcUr2zdfw9e6bo8k2veh42ScAE+ISs2RoEyIKRVL21aNuN9MnlVOWCkonPs
srOxGrkpTssuO5h3Xu7itzD46ppRf9pk4nQMDBNeFhLHibCYTUwxhp69R6HI9wY7
K/qYoEhIkDTym/+porEvesE+25zyCHrFkqiN6m+jvZBAddBQpeTSlrMyWpdDiyIp
QZeKESNQrlMEhZmmreibYVtluDLEbnbLSFrWD3yCCpn3ptOFw4y/Jm6q7XtrtFE6
sIloKCGaWsmevUxpvDSJ2Pe16ChypDFDfKcidbX/IKiCe0HmDpv+V2IyZ71qvLiD
OAzaAgReSQP+Qs5oJbuwNiPsMNpyEtMlsLh6PXDiS8dbofFZXRFPyWk+ndJQyPw6
3IyOHa2ooLVywCKmkDsIJXMp3oP3v6CHvsiMktQVJHG87kovE6mLF/me3HmeNvBN
vBXEhhOL/bemk/kzTVd/D2HveiAiAnUw3s36C/JIlXrjY089xN9/AWuROsYcxWUv
pwhxfic3IwJH2S3PpxJrG61aUBpYzE/1Ut491KDtWooued+16kXzP0uvALq5e6WH
1HQAghm+HFTtA2vjcwcksE78X8YLazah0rGZTCXYYtSkd92PnWll+43xRjO2nAXE
hVTxoUgjb1kKeHKNDGBmb8YqyruCiIKjCA2Yi98VhbrmEGz8HnPjQczExRV4hJl/
UcFBQrcBuYuKbh3qOM1p98sXjj1IIHk1SJep3pkmQjoKpwsleemWJlLzMPeCEexw
/Fh3bZZjtg+d0hapE4PN6qDIleDYqIcek1BTC+hxieej8lq/L1Fu0YjZHmX7+YRG
eKztr8f1H80HhItd1KtUzIRsEgYfJRgrH8T60u6JZj2hScUpFCEQ5anAaFrFLwGI
M3QePsiQAIkA9GuoshTQK5ZMrJ9bWVREpL/RVU0QkXbi2J2BO9opnJWTJUTAMXZ5
ksUpC2E5fN4hQik/7s1Av7i2RP8yc9R2K88OyGU730Zv/nu+BUc+zLNjTRVsMDDC
EPiMR6qkmXLpn2IWNOoJlm6Iv4+S/tctCLn/DWLq4Cwshg6Nqf+TstsA/aCKWZ7o
UDAjqFFg+Yp1j1omGVG3irCYS00ew31ee3XaQU/BoXl3J5l9Qeu08Roh8D/kAUmV
v0UcVrelf1A8lCRwswDuSNftZcCk74RMYCAMk9v5OJj5YapYYR1xlw1J1R/m8fAv
szhHMT0U0dDsHgzGwjsvbjIHsxVAT8sJshucNOwBtk3C6mwgaxDDQy7DqiEJp5M3
lT+Xx3VA/947cMAhDLv088nKwhNbiIVzNIvoN0nkGeLoSqkljlJuBbkAW+o6f/XO
TXsThhEBcfaEjtEJA98MPej+M8Na6erWayAIyr6eloY2o0ojKApUki/2gJVSApoP
V6r61+mZqnCMJzu9TMBEci8jENbmKWP+t+eM4RpclbBVD8E3V22vG0d2RootzxWv
4WLnki08c0SyQ/pvmTUgiPp9HVcuWyZCPotRo3u3xKIxIuCEWZyGj88fscdmCF/q
kn2nq8bG5UJiYVkAolnSD6N/jJ9dAblnEWoVoVUvtYNAT4tzLNcP99S7vPVpWOgK
SYW6gIeJHLBWWB8WEVSiKhCuBagQF54yKH5KoNP/4AON2u5QJA/UvXCsfXjlkknJ
+5p9sWpPLvtYcsc0kZfzO4PEsiI7TW9Kdoh2hAz+6//3Q2H0lzOl2ELYsmia2TsB
MjyTB75GsDIengpl1n0REv9ixsYhkFFK+6sIBZIbPVGLpvxTvfEvVyOOfnxmydzN
dlRHRXGvp6hxG/dESpacdW3sTP3WgorBqhYpq55LRMQbDMo+jQKujg5qbt4EO1kk
z1CH0lLKQe17ly1z72x6qT1mZlLYsoB7l+RN6kz0bSI5Zmf3Q2cOZqnllN1thySJ
aN+CV30y1WMg9r/c2tpfL/a8cBY+DokScQevvKT8MMKvyfX742FLuRH2DJfsr/HL
05xVIHyxvy7g7Sk6JhGLJGb5yb0oC7m5k45qTdnukBkH0PgHixkTq3KS00U2/9YZ
K3jfsQxGRh9iJVqYWK1k6PMXcBA1aZJg4YCBvRzwzRK2YIZ/qDOrsFI3Zi0xf0bs
GcazlN1LX+/LKUc9GGMd++QLW+b5rsL4XzG8gpbtAxXVRTjOKkUyREVqhAJvWJg2
Dr57CUbSyvuGmvDjBUDPS8w5iJ6pjRxHnicjtzuOjLYJSeJ8iwO2GWqsiNRIiHRM
dt1jRz5tYfBGe8e3x3i3dg2oHWOM9U+w0TzYZyrogm/CFXtzR14q+mmWwVLDveaq
Z5VDTxXR/1Dsw29SwISPp/AVLk/6j1hvOhDmqMSaPC3tZAeNYU256tKcpIjc85Wn
2A6QNiUg4J96dQZQpWBIzSLW0tq8FVjdbI9lYW0X8ZWsy3mnrF6Y3HDlDgFaXMHg
TOFxIjLkIhzNqESisyDnrnB+aDAJ97cZ0t9PM5EyxVqWpMdt1CilCwmIyeMqt2lX
ebWj4CdPF+kjgl4fSYgWuocZkKPXQo8BdpBoK15QjQ5Md6yMTBCh52jllhTtwNbI
EERBXB6pJ8dPCG7q1WM4/n3JCH8S/yrCFpoWlfHEr8C7z/WgjSckJolhiAhRIO0A
41fxB4TIoSjoLzGDhWn0Cp0PfvVlVJIHWvBlHmhRjylwYR9O4weYJLF4/qmA6u0i
UMtULaqe7yLRI9nQDwAtnI7qgc9J75rva2sNAzQUhFKf5ucog3+MxkAx1nJPX3FV
mwrrsIMKAop0eByivr9GlqlQViVbZoPuh5Zb6ZK4gw4YU2HQ1dRlLm26sA4COpdf
tV6SPN+lJJGWKiSqRayqHfPuM9pkmfQPbm8tXc+GhKZJuJz3UVUX47i6s8ue02qg
5uorhWho5/6L+1SVAecIXAcwyNiZNmm9WwWIZxjUWbrm9nk2F5UZUMrYFF+jJh1i
4pU4Lrolbx5m6KNHr7oF8lVVNpA00t5qlQwCHVfGKYk1z40+WzblYFCuZKDNz41H
NCFD39xkCD51CbLENWeYbTM/Tbe+8Bh86y40/iQxbkSjtiTNei9/M3Z6CDMDeRqA
Nto0qJqWAaoR/Fv7gUUCmm/5wezcm3l41zVIkgWE1LWU1C20653im4yHdLGrPo1e
TAePjlaIY8o6OB0+noj1CztY/lO8ByipN5NApJa1q09zu8EAk/dC91lY9yDsJIb6
wxIyWx9j05DdhhuQrBg/JU08eKDybJWOuozwOqgUD2t0xaRsMYgZKdcc421wZo4Q
y9kJu9gJe+9dkiavixOIB+Dfg519WemEMYNY459isXB30roU3zM85DXXq0fl85lo
Y/89as7hlsA0Aoq/Ia8JNrQogr2rXR0FmTtTJnTflgM2NapZ+Pv4Pfr65rPhf252
+Xo7ejfyGth/FDJFPhTGBWCJ6YnygJ4lh8N4Ozeti7aoAN2boTX92GOz1tsl2YsX
/JJbDUoQ5J47rGOKs14MNF+YXLbZgqfnWb6SGzI8kvESI6sweKTQd1Y0UrXHniIW
8KuJBK1hAseqDalVrJxK/pm6wFFW/kn5sIu+1U9gD8JukcSTEqImsPW9Udpl7ahz
JwcZE6u25PqPIpiV2w8l4Zzl0tx0a/yj5fRZAsrcXuCc+D0W/rvbDn0KJwjt33cg
QhQIT+j2fBGoC9hoVbGDr5ae3Nl/MXLhSk41tqu9xMnq4F+OPFnGd2i1aCIByDMv
hVvTgadwen5MF2gz2Heb7ntGVnPkWAcbwOxcCYNhIJxMEbtHsk+PTSFKe4MCplnA
BUq7KFdUBj9gMO3NdxiZxcL9cdUtgP11foQduXbeqRaZdSqTeMaQ1oNCucUxA6J9
rUK3eSqltT9EwvdwGF2E7jPGp7TKCHlYCxhaLbRZJYX/3kBGqyNg5M6UPGvrQRr0
antpXnMf4NiLekcmRp27T6nz5Mn5kWKyWKfuNo5e3k+MxxHvKPVfLAaMyvAnBMnN
27yWPTWIWv1tfnIZ7aoir4FwfEyJUjRIU2PU/H/F6UhA5AKlzkSMmLTYya66urfp
bNJdUQH6GHbqhTGJE1QFj3egeI4RPjuzM5jj0qA6QSgZGmdGWo7CB0oOHapWexEz
wO9RjJvNhR2zHtvAXzfehfg+B5H4blFO7GckYt6teqQX8sM0sEdgRte33yUZ+h5d
vPVNNoxPUI6Bz7OZ2RDums3JSvAIFUcf9AsgFfLN7FLcixdiUiyz9f45GBmb3PRK
JMmoT/Nj9FhmRy7bIoPTDCf+GPyPbp4dHKBC7DvKfxH/wXXxckg4PCsRSUiKdFEq
7A0ic/mQuHtnYnILO/y7dXzdkw1GYLyiDRVVaCMigGatZadddEWuQBndE9l3viUg
RonKi8bBP6xyoTD4x5rthPE0OwAMFjCYRupinR2fwTeYBZsFYjDmvrnVaEhkveRd
c4Z8Nt10xkcupEdUNyZJsEmo/bwO3PsMa7Ileo+X1wlhRtJNZIUwh8X6gkRmOFVR
scqUmnq8rUfGSU0KMe/74zm7obwyIKSofWW3FjUki4Nz2CjTdkWIGLkTRADjx4aU
LuzALcKM3CVyZUDueo/8KaJXsMi9RJUa272ZXRqQ/EK033//fTeJtgTin2tBbxjv
9PEekUcnwCRE8s5/a/4cb/+AFkCO14xl871pmMPGyFWVt5Cq7p9m8NYPymKf6Cn6
5M84LIIhOIAR6jm6IfJCn+H1gUoCGq4tqsnEIlAY4/xI4wzJMXhSxKAUqdNn1fa9
390gXspxiMswwoUW8GtpsidahPm8zuFN2hsbGrGsCnFPCnpbZQrZ7ri1wJc8l7g7
wPi6uBGW45AVoDKx7o47TImOAQTjrK0ZzC5AvDOUPhdoJIYjOR7OIL9g2aw5RrYB
BUiGfLZ9argGxmJjs6/Tdi88Al2r25lwyurM1NKaei+ofG0LfSkEXU6Syhgehp/N
/5IFL6WGX+ntMbXUhDt8JkBxavlnFNI/sFgrDXf0214Nh6m17N2KNRIwJOvhKOU2
wmLjhTpwRrImZCkF4SapSJWiX+rbJ9yasaCrPG4J94pW2th3mvx8wxk7ozp6IBWr
6cz0gNr6LORUrwthPCk+7i891s46dBrZzktx8xou2WgG6DjcJUOGNv3GiMZ8G7V4
M7jt4EYK+QRvDIgKcEJ3jKQlPNqhHRwUGjM17vPDt1rd72GXlK0uTgq/n+PAphYR
6lXEnwyyme8suklC885gmXunCwXzh8McFkjDzaL51Yz3QjPIR3o1uNn0Ao5roHJY
Rarr1Dj54TvQU3A+WNzJnU651brEObC+F9dZr92M0FAJ6ohXDxneBZSbv7uLFyqs
wI6cdkYs+kz8RQ7ezCrdhoyns4B+ATxAKCfZSOpc8N7hJNUH6xvIgQhT2wXV08Ep
VnN+GbjijXJ3W9jXv1iXZgNcnYJcUU5Y0v23ReWRMd2FXHg2BJW5Ze23s3uTpKuQ
MEREI5zXsRsJ/OMhgvY5os1cHdSzeSzQb9RTQlV5L0EBD+/JVgBt3VByJoPsqAha
ubsrAxKI/GQ7jgpmxiz01LTyKYCswu9KjMaJy1IpuPygsluOcFPRnuIBF2nWw/Z1
sufWF/6BVTaE5hdf+d5pr3IeDI6M26KahHznNonb/SvK62Cxo/jlc/6lZrP8Vu3m
Xmd2dUGvvqE6AgRccfYdUL8HE1a0x7f5Kq0iIpXtTzPQGLseze4DOjCkvHgX4UOH
4odw2+S4om9sDOdVnOBUWYXPunoUMMkuycG5gHjKylgNgu+OdVaQGefBIb2Kr3MX
MyvmdaofxhYmNlierCi0H7NZAXxSc0yfoxms4b4m/tJTi6pG9XDGqTlYVKpYc5DR
23VCaxl77lv/DlNFY9LkUGdz8CzWPYYFD7lkROMPdFqm3MoI6QY5L+kvKec3RN2F
4x0iVLdgT+IpC2Ulhh5eH6bRcb0lI0VhR0rPctjKL1C6gaqimwjdkQfcg5ULPkks
3pX4p0x8B84OOVsRJWSpSrm/1yiFXlEzVpeJdtphQDOWMyml3km6XSyKbba6j4FK
DU1QVuFW0fX69vhPIyrSIEe2AjQ1kZNTICLNcsByGgnWtRihuNy2pbmfGQmyCzyI
tO9ZARcYqzAXSf0SlnhiSoN5wpovxc4YtmJ8iQZ57RlbEX8apk+auSvn33M48ehk
EUdXr0GVLSJvWxEkbGi3odOWCPmd/eind7BBjdmlzv+TwFJ2Xx954y/e8QiJV9sV
MG6jQuFR/9YjwUiErHrqkB5rrYn1+UFHQlt3w1aaPM6WptCeQPiTtJOJ+gO2an4M
6J5po88isufpwVMC5KWy4TzhRyHD3O8M9v+qLU7dGMhYw2DW6IzUEVEfr+8AehKA
zx2RMsbmd/Ft2hR0iggIf9k4F79bX+AFd+ZRqII6doI2j/sMcAzLDuSQhjb4JrWV
XeAJ9Sk1U8wvrXZPTfFYOllHCoB17k40p5NofxBIo2vngc1ReVCwLnhC2J7sQqVP
+420+AJeD2l7qCoMmJdz9X8ixechwx4vtOTZE8lIvz6xh0XGapPdOqJd/SwKGbdJ
PcFERYDlmW2TCJz/UKg4ZlWI7tm2TSembeoLMERXLm6tY0g/2G0krl5SIEpXs0AI
fhdM9Yn+0NwnFMQEwGivMM2iXIPVesmVkKLdx2duQ5yMZFlZnD4a8CnfHlSNbSWT
5TG+Qpmbg3q7fHre6fvomr3Lmhx6PLBVVHpEaUNnWt4Pj2C4QSvCmvR4mvAuHMgd
jiqH/EJJa7dif3OjUkS5tFCsUfY7EatJSpetyNQL9RGl8KDY7Y0gOHQ8Np2suFVx
5zSV86B3FFM2K9uBWnT1GdDWqhn9BCo06ON0WDQm7CBS+LJHV+Z50WrAoux+nv9l
FXcxp6rPhy6ZxsXUvdnFgYZt7Re2x+c6QT6a+FGdf893dFdHU4hrC00dTwPPTLNY
DyfDnXNyM3KFDHI1iweqtftopoRwApEeRI5HE7dG7GyxGpTor1np++Lyl0x1SlBz
mltfVX2++i6/l8QZT7Hw4zfwvOuA9k2nyDCntwY3vpnt+zok2Nm4pWDYvLaBGZRS
whOQiwSgc+LcNrk8QOTjWPloAg2shgPfhqOjgm7ideoL6mHJ1WThGqsdDFCulaIX
ZeQ8Xc8ybGcsgRt+dGWusa7m+Dk8eXw2TUABGEEjvdo6O0fWuvIBozGKLTQeMMqW
Wyq75VBsP5FMQWRO+0BFrKbBcLzIPIAboyX125X8yvQpjidPGfbxmbEYdUgyVtEI
8/eZPlFt4riaEopnEXZw3XcMna8HQZtF0q5jsnDbngVwD4EvaALUPjYyiWBZ8IOa
aeXFFMF2+hRrq25owZs9mL+//q5K1BI38aePDLGpPYKPlbLFZ9598eXylnX/KNU8
MN4DM2zxAKqfbO0BuYf7qHxuNe2HT0Khks72F9x72UhEK1iTN9DxC9/AvhLj6CLG
6ujCMfh8NcTf1+s8RxaPDO8dOHUF7pg7+tBK4nRWWZ+u2xjlM1uS9lkBsuhbjrHk
vsmqcxercRDHGX9SybcTtAiOHiDJsp6pRMamnPbEKVRXeE2zrAPkJqTlSaD3xzBu
1icK0bmwnKC3aUQUDDvocQ/1HEEUntK1B23h1hbguXSIJvgaoU9Ym2jQ7gwDBAgf
wJOqalq4NvpgF6c6g0UulmTp6r4rkzZLhiRiKKTk/WaIakPgyAgCRixYwktSmGkU
Y7rCV5gDKop1Z+4PsY/5hMOVjsbxqnkylw9dpI5N/WTtypn/A+5BF97APuMYgVu1
MuHJkHZWgpeVQ8oZxjamQW1W3Bvz1sHFxwAXvPQBPOwtxpf2ZUhQJxrfuWS8rGHD
5ODBX+F4QymJlwCNsO1Qtu3VJrrfx6Sbp/3G9BfX9qseAaR1Pi0Em3D7hgGl3bWf
Eia5Yc43m351Mu2q6san2SKLW/uxlHfQRJpkKuhQmaGLKkYzwJ/l0K8k4rFZ0vvF
L5FTRuSzylodjg8rrG/i3kRE/SIH0JfUO0kStb5GGs+vO9viXS9SbG89m46V7pMx
UtjoJV0EbtU7IIbTg9aD8e9V54/U55cqxwTFcxxGSXYIuN/hMSZPm/R0hP5W0YuH
qxQyRHyJpcndfQR/QNMH0DFXRmQ+1oTXPByJkMl3tP8USDuZ415HHFPJKQoUjLDe
SajC4Z2Cd8Nk/f/pkLLIbxH1aSpvt0I4FOgC0QJxoVSU1i7MFRkvwdrt0Qr6hEXX
fD7GdKF9kHmYYE2ra3G+chlYWI7LB2VZCg3KnPILmIyH96ivljEq0uIreZ0hdVuK
RLsJOqNz2/vl1HX1JxgS2KbHh330Oq+mRCvr27lu/m+jqiJpUd4rZXVXYdctv8Nv
yMvfuKcu3Ogt0wObXphtMsWGpLMJzFpBRo4EwSTrK8bTEHzBWEr98ZVdVZBZOKKu
8eJAHueGfHX35gaYbQIgTZ8u4N8Ym48Ah+skl9T/X1EScRvYMrkxsoU77TC3K5bu
r6bt4PSElfqeYFrZWgVwos5Rf9L/rYOpxmLsZXwCgVwFjDaYyiQAjvl8FXgilveT
oJoPDhrFS6VVBHifL2X91FfEWx2nuE+ALpWm6DOa1GFsJ7TkfAmmznYP4gdvUSz5
NLnTpkgNnuqMYRRB4V/D5XeAj1itSrN9Zdnmm1c4CHBSe60pTaBJMp+mghaVtD0J
hdxgbg6SH+zCrdtHgry9gh6jbyCYqzs6Ydj4F9/eG3iBMVc7i/q52cdzPyGGKKvU
cixx6Tnk0w+CNlIEeOYfUNShdjqId0V/lOf8AnWfoNvpC8PUau0XssQtKHbIp7la
eWDZrviZMwf+lchPaUPSgqT0uoTNBtoqkG2Xn3x9ZOgcCWpHM4wHWXEkuWgPwk/E
uZpS9D9GeqAa55Mr/L8eYtRtoDvW25w0iIAlqN/OGcwhHYj0XQsSpr7uK/zZQFYU
0V0oS/v9IVMJxfaKn3Tt5vw0z7rTZieuoUgQkKKV42QfdjvAZHaxI17WHPxXap9B
EC/UblCZ/nY2s468Xt6GxhekgQfqPgf7n1Pgil2fuJ6Ol+uDiO8lZHHgy3gZqBus
8Q7Jc53MBJkdvjRN84t+rG1rnm19PN+Hvk0AlLJ51UVOGut/EV83QbtCO1afIokV
ECl3v0ub8IWILL5yaNH6Xf+e6x0WTMPOUXzLo1zL7rPzlqRgEohl0kXWZy9ptBBi
ISX/inJt7Xxvqi7mASpebtQ8g3aqghIIZzs8uyMSxFdHWvE0ZmLTrWGbaA/SCBdg
6cpIG5k97jUz9Pp88VfeCUNKkge2A7quCaSWKNxczSRlMprrnebMozkcWpDuEEYA
/cpbdB4OlluREY+TIwigBL06VlyYiKokr1yCGDhN/1603MqS6MA+Pe9oknuGVubd
t98RAdIhsav417aPvrGjwRlaqMv0/vPAf0V8oX0562k0UZxPaCCww8p280v88izI
bfYCSF4dIYtXoLwzQ+nVgIjsQLiMpAnUJ7PWsj3Bu2ImQY+zE50+TzECH8au55Pm
+AXvABYHxeb4WQJpVioLmt7bXweRyC1Qpi2qosMKTUM2OadcymmW10wZ3oP2X6sp
R9Vjx7eM8j+djjeYmsUCxBjyIYK8kHWxBdMwk8oV3hfF3LgkpQU1rUjHBR8JZjOl
zS+wTy7vb4pRajwdc8tvYUOm7/vzP4g0NywryvjzhsODtkPpokT8BJCvuLKIIj6V
6MtMG+CfbuR6UXzS+cwjcIU7oGBj5sReLdyEz5d2lUm9uGOk6Bb0ypRDOEnVff+B
k+4Oi3yoJfzLEJjJsM7QZWJm8ylnhVncPRclnG/cWU4n2xbLm9K+S7CM1gwzbOpG
Y9G8lhlT/y9bL+E98pPvCfpK3Nb3qO3e36dCovwb1KiMZ37gvEMVFM66+xVMpihs
sd7CJ8ZoighdVosDQhRNgKgjYoO5CcRKcWvHsf6fzBoiDoR4j+uZBOBL/itoJVpS
+jGdEAjQnlAvI+kUisnkLfPu3wToHwo9yNvuGL37Y6EoD2H9xfeYfXswh2JYjk9I
54sLBMJnKv+izAuwd3kl+GyHIB6pal0rPruPthDUjKar177OTqsOC0hgq23QozWB
kevBrvVKRdGiEm5wG7e8lOcCv4h4eD9qTKAd4voGgHpSdF5qgGo6t1jjHoYYYQ23
0o9cm4oUHs4Fb6YRxQKbWrVVNHWL0Fab0NREwE1om2pr57Qu66oguIl/YhNhJi15
aicuglkkENNf0uiGSlu/plteMCOizMdmx7oCbkUe4Q6kjVD94aI6GpGLwU7PfE4n
vVqcs/Vufx1kdRDjmProTgTTu0CXfC9UAK0re/rB1OPFkzw2HL3HPA+Jo7wi2ORS
9uK11WQYhsONzTIF/04oZSQ6BtUfwuGgXm1iOnXd3Pu7MkOjWeUk2FtiGFVBrFim
JPbdYLCEJC7AUocbtlwCY40IzmigPeIC8toNFjE7pGpml3zMFpTKMakj/Tdc+Q3c
h5Y86II9kws7pLdqvWPYpSjhQznk5KN9uNjodJMxodlt2kmteidBy9YlKT6yO2eK
CZlgbXtBEkgeZ0EkQHPJE7+8/DTMQGye5leAGR1eb2fEtbUWVLuOiLIE04IXjOQN
6vI5cLYpVUCxhE4frUW7ucBrwKAwWAliytlAPPAWoVeeoYXLJa9rJkEFRUWtZGKL
Mo9RtzwqagrybjmtVggF23xwzFRbf6l5fgF0qLwvb8zWgZDQqQQ6XVJwtbI83mTg
P2Sa2j4ZCwilyn2zLt2toxK7wAcg3Qxc7iiZTLS77S2UnCSoMJDBVoeRtCOi/v8q
MfDPGJTiEQz995b48P+rUr3sIyTIUaqTKkeHmsrB67d59Lhx4e8+j058wdeIgFfs
cgoBmNBM5SwsAs7U3Wb1m5FhSO/SaP/t1/4PniSgMZ9azHrZ8Pbz9l4bti9QnHtc
MDoqrxrLKM014bjFwn+7LueRh+W+A2vaeE+Umb1TrcF1nbcRHcAvAI8Qfbt7KBgW
+DJ1QMWVFYx0tRXJOYlBWCDIPycfzBHacdXudCZLaTBFqfMGgeUVi/mjP2izMWyo
BcGK6x/uiFRNcIld7G3f+UW8ValTxIFW0Ifa6wOebZ1IAXuHDUQ4Ss9GMGJQNG0s
bTfvTAGGnwHqIbWSa34bvJE+b69DOogFX7iO8piwS2jm4se3aJouYc50Ss7P4LJ5
8lBlTjah8DF3NsYUL7zx21ii4I0Lgcd/Xj26lDU5SOmcISZ45ioZ9I4SVNw8rH1+
NyobiKk4x/uq21VW9HJtGkYCyVovaANahAUdDfW+M8BnFz+1314vaJ5dAJjPAsjc
5hZin+gU+DiTondbbzdDyhS2tfAQHAG14O+jOU3yQ32gQyWCqEA9gL5W9tczCijd
qhFGawYh8Jd71wzAVpDUaXGKI7yMfQVMK9BhbOzP47btS3vdc9HmjFQfJqb3mCK2
2F92aFsnbyj0NoO3nevba0MwN2cmOcw4L2+UVUKnKCMnOBJtXmiYWgvubOS+gipO
4ZfMg5nHA+uTNK0E4Dj3j5iib38eRTcPAy6d3WwCXLQuvtsaFC31AFbeC0KaSeuR
HLz2xI3dqLDVWLNKA+lfeYwsiFs3WIrbCDp5cxcg0WkHPbY7x4GsuBIVD09iv0yU
oDrB+bpdlS0e1f7BWv0vnNv5lveaiy41UmaZYiIp1rRg1RfVpLylyD7ULxcuCJuv
c1YZ0piK+2MTDCXJMvAvbfmQfxxWYYKXz3S7THI68A9j0CmLPVL+nhl1hcFDIEgA
/XoHPirnwTMiNg8JRgt+XD4N3OPxuxxzxFtY05lDXbopsXDFOsH2Z4SYN2ZDoRnB
SdhfTZG0cs81XhmVMXlMHS6CE/merbyD3lDi7BJW3SvFQwb6V2nLYStGlovFkgIt
pMDwQbd/UWy3AO0BLhwTEmxuqF3mWyhcGtIWW0u/OZP+An0y33VKq0z6u+dq+FRW
lyerbq1cYb2lO4IbiJ/k6coI0YXrRMBxrur9hYDCF/JpccW/+XaUR7g2z29BLDz0
cxJqpFU5XU7UL4jUIKWUoLvaYR7bCRDbOaeN40C1HjkQhbfCit+hHXDr20CLn4AA
hxXJ7xrsjNzUKifeNF1nW9a77lrTkkcjnc7XtkrPbzYJfR7jttuAM+jXASdX9KVr
olGLCPH180yJQ+1OSkREBys8AElhDjjsfe9EJ5pWJeMDJ4ST3LsCHsL+hdMRS83K
xRyj1lunub6GvcMzX6zKF9iSqhmO6WGpJXWzxjG2u/AiOsfLoLF60p2CCpjp0YTu
Md7xaQ4AQ1G0aCfSWGDpR/3v+KuAdjrGLu9NoAUVFpWEEL+YLjw/vjuWfBBQptYh
ku088fH7BV6LaSH0ITvj+6AeCZrXM6pz9sA+kRGF4tFggk/CJE7v7krb6tkOxCme
ejY83F6PJZNPh/EUlifMk/euUku8ToNGGW/7fKn/L6jeAvLak9KMKt+O+Xccw4uM
PK1Nb4Bja/ThDV6/nzkU9+Gt6jkMpQKsbzSo86XbNNHbeFo2yZYeEapKX5vxbCet
q4K9KMiWSGTZvxR4nyhuABzf/RxJuGoQw1DffRk0dsy7RO2sphwAxyfweU9/F/gM
2QDQU2KBgryv0M2RQsU8s5AO03cDHselvW5xULEdBmdBph55v6003H1m4gBqi2UK
C8QeSh1CUf+DoUGE1XmHLo2GbkoqU6I1xqEoH4/LIIIuS9dHT5sVYCml0QJJHLCF
pZeLf2AEH7eCvF65/3k78k8k79yEiIzKF59ge1Nb7fl+qXrwwiz2mLqNHFSzMAto
84cRx2KDl1RMXzgUKPkHiheXtG+HEhqVtXw/BaOc8269BrkOQjtPCd+gju1Q4Skf
h6tPCqINMqFOfQU+FmS4xEFgMevKXKxN3slmczoUOStVhxiy9xE53xjumgzzuu3M
Tw7Fk7e8fOpvJEBUFYf8b10HvmEhnf14hCtBe+M/ZnNQLopeTiCay846x/gVHL6e
i2pjEamJy8o/ulzgexRz4uZLKdnuGYmt44EAyN8n+iWpa0bmhzg2Omv15qX7NS5B
FOzVYTuqqRL/n2NE3kybZWBCqN34jNzaDqDWdJnffdeSmTOegX5Vw4YDglmP1CB2
O3kS9AeLOjwaRl06Qfr5EmVo7d7V+0C1If641V2gNfTWGoho8Exnc+WA3ZFG041s
/z04plh3cCEHZ3mvI4nJFyiqr6R6LEgGNi2ivZmGrbLySXmgM636/KzYhBDpqrtr
80kxd1JIsI2665LJguxbXWhSkG4XRMZ1fWWfUD1/s5j45NZllwPIrVgllNE+WEsy
MGUBKg3Hr6hFbbSn55cxlxA4bEcPkn9AWsFkbLm++3zk2lSHo1d3TbQsWaPPjJxh
0qNpli9wvG1WN7qd+oQqwJ/TrhwFiS7ViYNcgYLRWU0jxsvZGxbxkY4RAUyr/AbT
/Tg4weKICb6hVEb4yIbhoD6ytY9wdj5RPmk8vQjXsKqlOduJZIMuczxsZqHMF7UO
yv0LPDGaIgBK3uErvL6LRBwHBaz/gHXc6kBETrnnBzLfk+IAAjJI3t65/f0d0J3g
4CSbfN9PwRaTby7pRkDg2b7Mu3b3OHM4mv7cSOr/tWXZPV+lVtOiU4d0YaPfmi7k
cSh6AqJJB1L/fq4iPRr4Ac+pRjQBiNeUk7Y0iRQrCOBKlJOljm9S14s5cBUIGC/S
RqgKvZ9nA3NuIrVE983Yx9XjyDA+/ZzNLsqFCD9ofCHAXBMvRIIaEokczXGkBIu/
QC3lwI7AuzLAizXoYPb7jkYs6WlPyjNP+UaAvaKQcbPJOortuKh7gVUVRgf5UFyI
nUnmBYIwJtpmqrXM5RuPSF5u0ji3WaKvml4cTnKWUHJqWpLmP37URQ4YgwaVDKeO
kEf7m4/bT1Bz76mBSgRewptGjuNTghax1unr6NYm4DVDxTNpb9B1zi1P8gOfCEMr
VQnwz0A/jysX6zs1dcH4hk9KHt7DQ9VHVbfJl2m9dMKwwjH/I3tT+fmJs2lTNUEg
Rzk4fCnPdrDzBdhZQwwteO6SFxa38URrTX2aNYBob4rtlFKUdIprGu3H1QDr9fj+
PY87KNPk3W6dUVh8VYX/KfkwWGaeIgiYXyWIQ3Kh5hY0NZXW9F8NyDI9yupRJBlC
xP7U1Ah72NkozIlC2q7BmACeRLBZYRVSiZLnfSs/vgLbLLSJlFCKrPNwZPdTSHQA
JtAsCNIHyujohHOtGMP6ZoxH0P9oDJiALULrkNTTOPrvsEiW3EZzZwGY0HbQELOC
eUMguN+LAJIC8ZZh+/pp5yIVrf7gqz1wAFyRywE2ft9ouEXWUPzIdQ6dOwKQf57i
T2z/uBimm4rLgYF1O8Q39hVsHMUpKwj3mAdGuTfRg/4mpGITw+T+USGeBai1m2PE
eNFoPxl1oCXCNqQsAVSnwmo2c0IDzjCHokVa2+gUh45XHVc7ek3+LbfF+RvxoCmJ
aueleoxqLl5L9k620II61PZUZnt0rZIeYl1aSI2aawAkt6nGbbjdh6069S33nuHT
m4P66j+u7ky+bjrjOEigj4XbsHz5CjXw0b3cinXarIiTyGGHVdGMehuIr1hpmxZG
JZOOfHShOjPNNITlNa+LxDB7BMdM7BNgH9zUuOsuXgcduOy1pjy8SqvfEShYa8/Y
rSEQTAyVeJAYr+ib8uMoxFp1rJ9ytcg+OSyQOrCAwv79+MwJLNcBFdTbyXqYanYX
zEWQ3g/oeb0ywt9v57CPM6jp9NNvq+qXjDgg6GMBT81O8z33RPhEcOyLGByuopIU
qEBUNbHjxK9tUkW2weaavdforWTLZrMVqcbToACHwIzQCkSHJX4vuNlK+Y6SkHp2
oRXYaQFcA6Ezvg3nKnf6uP6Qn8eDyoKlipRgVhkmtUUtyFUmcJm24AUweld13Xba
S3X0lLSTqBZGS2Cc9Bu+rCkqO0uMLTgY/MX41UNS9ZE9xtgIG0Ixjpa87RHIdb++
ogIVeQRQN2df/eaxAELmY1Fug4gM/e9xK09bCbkiMRyHKk4ovhpZneEaoduAkdaU
N3PPEHdJioH9jRML27rQuK9sETEaah6qTyAIrw1VDN5AqoPdxKD2CNiTjnlBWsVb
6Ar9b2bcnTBGgcSdiAq9uwJ59muVwqD7Eyge0TMQXNtrVMxiIdbSZthi0Kzjo8ie
coF+MtdSoiv20I6o8j8b4i3OWB+Fa8N9Hma6grBSyEuxDPEzXUBd4szcbJXnjGIk
7CPW0q/yBRAuwdZ+1AS9mgq6klMzMsxK8MpWI1N2hO64twGMH18qNaPh2SUaCQcy
ZesziYFzrNuZjvmWfOVRnl6Aio69ma13JwkMExxrMZz2r00V2OEj4RcPAEVcArt4
Ed7eeJvC1/2n1acC58jY6uRrbUQciXrLLTZpXoguleERS7cBUya2HMXUIKsPOsbx
vZaV3ZzCsNrY6FwX4Id1SazM6a8s+f9jpHYEz6qHdQETfH7BhKoAqKEM5IFzKNvW
Y+CW02bEJkH5TCBZY/ILhALzrWmkywX7J7IPEHLuOl5OMAn63uks5HoxRAcP5Ytx
v3W0TkvG8aaSFgedeHPVOqGNEFTH2df2uacGVkZJfpKobB2wUo2dpL3mo+dN8yOc
LdqZ680zTuVXf7+s2B9j7/Trx6TfnsmPpBDmiYVTQootLnVvKe0YTS4oOAJa50fc
FwTRGHJ0jQpZcDBjEAKoOPz0ff3ivZmJQ341p5Z2tZkpGtehDRK6l6kt9pA+QjWq
AwQKamTJI2DLqM6fgH7FEHO3zky/bbbg6QYL2lJdqaDTC3p8I+r+4kGVC1TUaJvW
FAxQhGCImHUYSsZoL0mAf6x3wQ92HuNAVzUyElaIo06STgSD6YXD6C8hRbVYaEyA
wTshY6xJLHrvhKeG9qiQE/fPni6mtrzNw8PgtQAOqWCdMrAkb13FXqM8cv11b0u9
6hAFPPwgbS04x8+veReziux5Uk+QULShGS66ENMMGVRZKBANf2jhKAwO64cEx1zL
Tmk/HtemfQvMiRrP3sgrEF22ajz/JF2gUg7znDlk/zAFzJ2EvORjkswiEOpM90OG
Xfmkoj8eNzwYGWBhly1XgncNRchDC1lvZfMQxSlsl1iYQh9APALjQqdElLSd4LF3
lJyeb/LiKtxwBqQhfgJziRUjPENSs0irgVj1hKtPQw5UtjhvPXQtt0fdWstoJ7bo
4I9GCEjK9ITrAX2o8vf7mQmTsyOgrlMu+1x6hTOUvsSPNtNCTVsJv1OghGlcicr0
K3KrRqwEqtggl+Bojtzv6xyUOFHpAF089QiKlo/KqUKlnoFevWfm2G5TKxsAKouk
7F+ImnPVQsYo3l52w2K2mzWBM01uRfpv7tR1s0Tr47WZV+uDNTxA3Z6JHdUAAKbJ
EeVqBQrnmtWrGLIN0U8uZKxWYZpdPxsmF+34cYeemx9yDqEHWt6VbQQNxC3YiGuT
TTUuwn0WlFqjwLew8B98aTTJjE/c3Or1uaGJ2lLh8gt9fSEjMyuPTMLXSRmArH3+
EIu0TfxoWYH5ixKBtQ45L7NZCLL/XU6KXOlTcyHFomPgRyN9+2lMLDXf7LwPjy5V
1+0QLj8m/uago+93aXnAwSOM/EQAvgorYpDM7BFMjgOJ4b+DitFxNEFbwpKYYLi4
8V2iLZr3OLyRcD3jnm7XhYD6YK5cl97iSNRNAD0KPGnG3AOOVH9JyKUCb10nTrls
7PXoETavRN1WLc/ZJDE+f9K+LPtkBZNzEqOkEEGl64khyix4Afh9KSsdvrNTM5kL
RvoZXqUE8iw3Z42nqPK6jjtsOJBA/P6F2l3ZynJ5llyClLFwgVHUqgkqCJ/6gnWW
Z0K0d2TH3up3UBBBoXyR9JZIyqHKKVvrD1tksuDGmDVcPMUCdtvsdr/xw8Q8t7kA
VcwPjG7ullT5e45r0HPxfSB2HCv9M0sgvr0zIwJDntM8nFDaIUzAflofRKqtZdpo
+dPxn56C9CjbkGOJoBVYLv59Oy8HrJ+DFHPpRuv5QnabYHPkL2M45+R7larUKjdL
gPwuqSZ8eClagtR78VsjlW3465lLE4woeJXKuaTT6g0CxhbX1p0xCSwJ+vZK8AMP
x8G5CBc6SuiG6mttEN6DX+fE4f29Nm+jvxdoweYkeelqHeRmnQGwgPN1CRRJKUir
o3yHsdb4YieMrtWuYu8TtAfmK73iCCrgh3p6GFDYtx6rZfuM66IldZieRINUFmXi
nE0zvWs/FZC8MQw7TjrXt3MWBX6Um8tzxukAvwTKymv6BepYSYWP09cR0tcFXTjl
f8sT7aiuqddUiMsv6cAGtq/aBQYWaieRhUW18U7X3xGFzQmbZOtVYOeZnWYB6P0Z
PySvK+nJt+TpbMVZW+E90X758TEhfEuwT4Eo1M1CbvSnNNYVaZtHNtxiIW0fmCf2
FawOgbl+7vVI88z90khkZy+gpO0YZJ/VFQ/CZeZd5UxtHuMxyd9A9GZX9zqrBLMZ
ZbuKOlcVzahaGZ/k+dvOzS08iQm8HJ3oaZiw1MWzwYxuzvVds3PcOIn9zjVtSxTu
rYoV4Rgezvls5QH5Y08oYXkuOPH7n6EZfGwdztz908GIHWsLTcwuL+U5gR3ZHI/w
Y9o2ydEQwCcSpcFm9LRyGSDKJgqRqSndCpnGUyBgtoLcvAB/zxi2x1rkeui9fjkm
n4kDJb5oxtBkTmxfgTpaes6AbZZ1hqJJzl8ozpd+uFWwuQKPcCQns17p2YZPQNAr
U2aBhoQ0joV9HgEutneg0i1sZUiFPbmDRAmb4J40CH/kSzN9+JqiqKkjjGhTEmi+
3aniL/mqhFOig5W/JMgV9dzUx1osqdSu40JOSUDbQVPtVwxTe39A7JO9F++FKWR9
ufZ6i0j83lc85Ao47c5sj0SniONB4HTrvTUKMYklZB69AI5XeTqeAMVGCNgeBNx9
cCDQXINH6Es3WO6QMjtHblK8tVpQBoa4MAAlEqFmWpJPoKK1WSwzgjD8Oa+n13pW
PUWPUmuPL2/1MkLk78ob3yya7QyoWO+hETcB3SSj/Thfq2i3kIG4wCrKSIodNRol
4yY4CdRnV4ZVfFyfebkoAxbeeQQfq3NtHs+noocqbQ+HzfumUSZvPHMSO2xqvSo7
DoGBMW+KOLwIYNu8dNWvr01b8/Ol3p6iKfak9M+mprRruab3U/+YKVEKWzdmWMa8
8lbaq10q9TSteyPxUe7d/jGAiHgLPebiW1682dugyRJBwn2CeHfUDROpJtkhSMRk
E3VSomYhLAF1/H/4sbPkyaJ8DSFk6RN6ChUZCfHfRwZeVNlCBpkoHsdf18hcWHEl
hE1ZT+rzLnDGCKWzJREAbOluro38aIhipMfNyOWY21DiW6CExPSit8qYV+fKWdKm
VL+3KFG3DHjvrNBMEAJ1sfiT3uSeuvQxtRY7iKFpY28m/sPTK4BSXGzhkgYlttna
OzmOXdsr5rTVz6iUQudxDCp4qn7ne0Uw31VHWID4srmEOM4sKdqgEWPXlTBMvI3Y
ik3aLros1p2wCNi7eBTEV1KnY1zdG/hfob/005vy0Fe3FMOrNr8EiRqMDuasdVX1
aUzlBWWGe9g0r+v/cXUU+4L4t+VhRownDypl7zsz2s2AeDP7Qm9IIA4NLnuxPDpo
SiamsnhyJ2YxRf2fnZXjlAlYBO8YJ39trXOmDaFTfu81ZtObqmbOj+2J9ARcN9VY
xDWxd9vETyG7Yj+jlDS/T7lHkbXcHq48UR6SR6ADUjjI/Vq8za17pII8+U+JiLtt
wOaJWsbSXiSzTZH8+G+S+1awH4yoLEZu/tHTVuHNh4ZfGkov4d9pc2qhtVRYCfit
G4PAC12RoluBbRQP8VOCiCBBWOplRyXczSFxFeZKmvY27rlkLD+WrL7CE9TV5+z/
aARvcO9adWLngkMlzlRnrPMZO2gFtMLefTNUD0e+0tkkYaSYRmq7nB00KKoJ+vqA
365u1WokIw8po/J5KQKhYpqIiTBmHLoUyf+mAw5bbwu/mtiLeqMcH62BQchDCzMi
Avw/KkYjnzc9lLZRJNyazn7nbT+/sx8/E4zIBR0Is7ghHB4wAb80m1YSH06EWJFq
C0ZVnK9OvDwrIy9ml5WpqYhFdCwGZBTImDgp5R99ZnSedlMJIQfEYOa2DvuCYCtJ
/N9yR6E44fNjIlsDTkw2WQMMraQSFSZWG66boPklBhRLmz10LPZVGnX2IAPUKXwZ
IeUvGAyNtcIkqUbBbpSsZRcUKdqkO9debeEjN7LwC2NYqLAtVcwQAYWoAN5p8N/L
oqCAcyMDVXXJ8+K9cI7qqNy0TZuiz5jh99sDuPbmS5liyj6OyivtiO79TnGwypOW
rK3hgVlwhcjkSYWjyzelF3IWrxxKjXjjICz6q5lUfdrWvA3rlaFNrrjED6e0SXtS
h9OIpKP72vpci+dbwuT83rBIQnsgJSzETL6TEJnA6bo2E/krvTcZUxJcybfiSkHO
0NYTURNHJFkK+JvMsyuwcx7/kFJg8jeg0uOUhFxfEZfHcO5lV8II8so+S5fgoXoN
gaek9ueXAPsOGdPS+kWoDsqTnQeLowVFlx0USqKFaQkO5oYg3emUDYkEHDVgipTx
kmN8HQm424LyAFkX+b/AQoZmkn5935R5TobBvvUVD87NaxIciSDd/qlUr5eZoCLQ
h5MzDkGYWNnqEZzIwP7qA+ULOtDUYbyiBy/5SdGe1fL6BLO1BKYFvX1pUk0+19lH
SvL83A3piwzCfYxI+WVDs162vENxGLgUv50jXMel1jgMmhdqoU9FBRl2mHTb/rBd
nI2TwAEbMKS9QgX2AA+Uzs+wyD0ovITLfqy/Hx3rPXFayNCUgBVqrQ9iT0SY5ybk
4GVqbb2biruWcdDlS6LqdmrlzGKAVoVSk5sllwxMaoz2VxwOpzXJS6k8UJRR77NW
0jQq6M00Zo9eLflt9CTITaiL/39Ui4p04yK5BSqGXQQz5Dn4rAXBUXGqMC5EA/zG
qB7QLkgZA46mIpJyOtOYs+RlvGqt1/ADiVM3BNRJd6bofuE/p3MDCDxoAhAeyl2T
q/wYc9bSRsdSR13bozm/0q0zsFGRCkbaZXSxj93T3JbJLgwS9xjmOTS2iC60tebn
k7Hws8CIj5GrLlMvBHaTBdjL9xoCmPtjLZpNR31wPOydxIxM8eBHB3NQEYiFbwi8
oXXCR7JU1+GEs0UMvA20X5l3HBKljGqwgKEUrUf3LCTYpEBdolZx0NkPmiADu+Hd
fn132D9BQzlSU5Ke16k1eO5x9I+xd3s3aEfpKCy8JeEhy2AcqfVpvzMtQNHsJBC2
O4InHmrfn9WoHpDE58PCDxhZB3fJbDtM7gDF7Gl6IjsKw3gXHVU9PFc4vjvG1Vzl
6GDKnM6k7obudo3+U9JklDcFeHbBZ9vgtTt70cJk6CmIGfe34Wl0W9vANlKmoc9E
puox5GnAj5p9PHpKZvaKE2kX26V5uiUYhWZxLf/QKWj24d9Q/rqOoD5Ppn97qYfj
t292ZXZGiBl9ybsqDaKupr0YZqbULz/q48l3jhZ65iUIWZoehNoQOCLGXinFjRWu
Z92PMrpZsv3F0HKQPLTclPSVWQeiymq2/fv7fCin2dRe/Omlw68qPmaKfgfPcsaM
jJMzecDrUlE7qiopZn0VyGm7jO4WtUG9ju91GbcIZAPQxwfptqRqt0zvsVGzwx3f
eQEXMdMY0PDRgTpMSFKoyV1RQFfeAYjXKl3XDIDimHHD25tDn814YHVxruJlBgbB
abNvv1bfoMDciOj98tVodvL4Axab3BQNMKimXoMkPJsCfb+M6J7j1dREsFrIDgjL
a7q1qSYrB2M2yOjJ/aSxRztxOIbHDqHzVTP6IhgXJRheHpHtxQaShTffUSqPnnF7
SB5xxjUD9qK9oTSVihPrYVgb7hwg6YvAXsKxuu40zuOCHp3144QTxGcswWltQ/7Q
Hq5a1ndcfmny0r0c4nUMX3cr8Ut4RsJFxup6sJerY2r2IjZ28SKWiBVzMj7v0jyY
e3m6ytTtQGB/tyK+SzJ6TqbjkWknbiTh0VzK0Xma3e3Z2pKj4abGmrP+aY612Or8
QrFu864fvNtgV8uHa0ZC3M3KgqrdnYDmBSZbZCJIF/hSB2aHJtwVeIJPso8MdT63
TNZvj9skgbJ6d1qZo5CZiqgjNt4cbFzVSBzwhn6DN78YQbNNS2xSUgnLq8FcAiuU
E/vVaHtpwLl/vLVMmtYKfqOSjgbRiwnT3BseJJjs9ljF1JG01kJiekMHOFDoWg4N
5gGpZ681bB50QSacff82+r1UYhvWBmo2xs7ehs2Xy7pFWIPv7UZY+w4GFFDwg8L0
bEiJg5J9ek8dohFlbDdKh2gC9Pn0+ffxjvTCmK4tlFk+cbJNW4jlJqBJ1xczm/Og
+8rHfQ9SCPp4GkBjfll+Gw55IDqsUQLI1zMPKLyqfxGlAGs4Vh/8XM48TEMWc5WW
4mEVnCCFbNh4pXq6Tt1vPPyJWlwsKA1UJzD5JqW5yTU5SDE1WtF6oCXOpVdMg4Xh
wAnkNQNA2TgdMP3eAVLBIwGAGz838qxCeH9Qih/QisTxJ323UXT5NJPUgualNwz5
YSZYFL47JRV/YYODSNGjRfxx1O9CkVx+q54k4ryev002cMOJNUX1bwfogUz8HyIB
Qoryfs88GR02PT3KMt39JC/7jaGUPO/OwaGvSZV/NoUZaC9XYtm8X39Nsr7bX3Dw
Y4BP0HXdDifnMYncfQhRRp1BxEfRWV6+9iuxg2jxi2g2v5ZAWuWK+wGa1kN/LKm5
tiXLiSqOQUugd37H7PY004P3u3EILDlI5oMrPyxm4Co03BROfZo90Vu6RVtwlbY3
1pn2MXRfllxw7FJ/taH0CH6hjXkK5EShEo1Ue+MnxbO5ey0/QNJzsHC/r7AeuavF
QJYX4I/o8iFZyjtM97TjEKi04KR6y/5wxDp9+kqsctXvY4D1eZ2G7zdepbCzQb6v
7hB13TCbr/wis0y+m/O+x0nzIe72NFqvxpPsOTmMfwjCVDmebWd1h7rSGfNqQpWL
FPd9a3Tg1I8XpqeiajeJIULOHRD+BurCiC0J8eJE8iP3na4opZ3V3augApWzKAPX
Mn5ZX3GYvpwJXW6bfpvBCZkLDzHbNL5B6ahanBFnj617QGSdty+ZWW16mWGDHZrI
gqag27hx43lPVwl0bW4ygd0OTm8Jjk6Q+7lsyazeLE6Rc33ZlJscIEXI01mzTCX9
DYVELOdUW4fgEjzLpUffz7ppQNI/S6gjms8Dxa9tLVIm9ppd33u7VfLCFpcInOU2
R6hyayCPuhkaFYEtNSvJk2lZ2IEhkVBlmOX7I8GA1ZfxR0/ACd7euWQG/+ob5OJo
8Jt4GIGpwHnX0b7i4XOIR8pMTE42M+UlzDBuCgP9wNWji6qcfLbywruP0Jn7PrjU
4CT99gCat1EhQBISXCWLvEkoU67VuikwO5opseKlrJN/fBpcr05IVKGWvfuslIP0
eOMMEVwCd8QAtgiD0W9hoiv9dKASJqLiI7N6G0fZ1iFWlCKyp7IUhgbZ6dxlSt26
ZAsXCI190r59DBnXdqT07ncQrGs8M4lzSRpVJXZwQAfU6PQbMzkhzcnFa30NKxFX
TVXISb+km4hdgyOvfRC91MdPaP/SYAnJ2Sv66NIm2+Fm78+2bObby65Q104aC9P/
zWLvI+6FDspODpMjYc3MwAdDNP09/SDlXVJHoqbg1KOyLm3V+43sJvEh19jI1Oz2
ceqiguzXERfx26JBvz085HZkb8AZ0hoGjMUEIbMSevZQx91zPlNQSC/a4JPQivp/
PoXKXxjFlMZpin8ybWLuIHnYomJ86+l+IIDzyAutqiohHuHyf2kSQ4z49oAYvMWA
aMpIKyCPMktl1Ld/rkk/HWel/OIfoRoNeLdlhWrLJLybewNUi8N0jYe47zbKS/v1
H5/JJ+5VdSigBEJHAiOqUsmlKo60uV0Ht6ZevXhPqru8QgSadCT3RxMTBLGAhxeA
KYyXBRjlMtYGBOGVbw0OIr6WUHOXbko46UDEu8qk3P0OeDfk7i4FPCKzqYJ+owMH
a24qwzhNVFwJA65IKhDZFUCT57xhH0GD6x51FsuThBbBuPyyfJpE6TfUjNRx5RJ+
TuWydL06+ShH1CMmzn7OCApfEgjSk1QJbV4DOdpTsUWAQj1/545qcmmvVHxXAuNI
bm/bqDRKij7iZiERUAe8DMrA83O0r0yUi4ILy73Am5jm11vsbQagYRWJVUlpZ5M3
W4AD3hZWUWEYcIvxE+O3fIiO1f/j2h5pGVqnE+//2APjwp9rFpVtu/MhVt2FgR5t
KeWrdxe0zaTw/ZajfVNO369ETX0Tjk7aFwyeXMSoA7+ZcUFmAtisnhc5JOyibkCZ
gdvZ6y9EInmanfJxNN23k1QXrcH2kVpQ9p4wvJ0+Si5EmFeb2d9c5dPhR4u1yhiw
UdYLRUtN1OLulVvFYLoFfz5/Ea16ZggKA5G65LQzfUvTD/GA33RdD9xAy5LO3h+H
wcBtpqUDzcPC5D15ZTqbPnGK7Uc3u51MFT7G3qN6TSOkGI6cMLNIjgmVa8YrSPQP
sRg7mBPaCTYqHbUtsGZ3b3ZvKRS/8zqP6ZXSecSXLJjrxU2EqgbxNexcOFITy/Eo
CS2Kgyln818ElIOA941hawUbmpOA4lRO2TaxOGkC31Y27GJVyjJw1rT1ECq/r5ty
kaugYM+zy6h3ALPp5lEKOXzmHOs9gz6maUvP3hkt3LThrpn/i0bZHzQZ3oAWYhtL
go+kakfV5fxKqaZbavz2/DV/Xo6JJT1pP8/0K5/Wf/NIaL3yVRbg00EQLyJCvxXF
jOiHc0Fh9VIrMflali4NxrU/kU9n6delQRH8ZmdzlZrUKVC6vPKWIrub3ty4Jit/
hX2I/kgX3AT1GrK0VdUor5vlVuyFT1oOqs7mi+JZ7Udus3SbKRaF8mTFHs1EJHA5
+LXXtFJk4kwEjz4q5cCq3F0qoOkWB6ixtUokIynWRPhd52ZroJZbkcsU6cqeSaMf
GujvlM6M05KwG0+XbeJb7cxmS7jAcBVeNZpTofK3/c2NRrHU3d5487tQdhImwHA0
lsWgodSF13/joUxsS1EXHqJftC06cE3Ca6DBmjp58HZV11rvgSjmAwD5yGFMCk06
GVAS+m3VVEO102yiB+G9V3h9fnC5XbaGQC5p5ymBo14f+aKdjslQ/bEiYwrftTUg
bsjYCmvaYQPEMfSSK6LLyL8aOj3pGv4LpSlG2Owl3iKbzgOlo0e4gcKZa6iiVPGn
HKq16Ra/Ku3bP1tSb6qTASuYs/Okow1thvVAgzklof0rgDct8IQ4rGW0PuEtohgR
cWiC5sd0Md0QS9teYXPMvgp9En/QqAnkIHw5kkLAHz2oeaEqm5UVxmLvm0wZdr3v
8VwP9Y+lE531N8PicYBt3Gyqs2uxrcrTiFX7I7CO1YLjzUlWG3/YsM//N1lvpLLc
TxgOjINIq2UslFqvbk28kYaL77f7N3qT+osmAwmXU0XcIp0PXJpHTqYgVVruS+Tq
Ci1+K3j0r3bXbT2L2iBt5oLZG57r6dQQKk1eeEza6MpPOYRKg3j3jwRcQctoadwe
rlYKdGCJFwCKNjG3L3HfqHzcYsf8VUqBd73yqtN/7XP8aJeQKAOQFZw4VMlk9xmZ
MILmewqLvRnQ28c5UO/PTSU9eFFsIMeTnWQd4W5g0JEq12qOf9WmVC55avZ7XGPN
M/Ct2702GYg2UVsARJiWpvLFPnHg+Vgc1T9abPWCVG/D5yItSphlY6WqNkhnTLL7
iooLvAKVekrfq57nUp8gJGZN+Ybtkt1zIP9DLRCqqR2gKHpk841nPFboBumbkKht
xGPDGDHIZRDyIEZrM4bOOa9KQHn4e8+9z1yruQyEdaSp+yZCPmNqOsvTzQKb0zJf
bKiZKK/EqdCpLJtXGIhzLBXql3CBVlnq1ctSRfxhZKeV5Of7BQETdRNSJPg8oKQq
f3d/Kf08MQ6cgUb85QrocUOMMmzZxxJE2iE1/YKC3OMXQyCoU+MTONN28Z8OSNW0
iv0ZQ34oCjBThZS7Dar9B60/J0S0VUtUr1RqPrkbCBuDLH5cGMvP/UmEtHqef5lL
G+zKMkwnwymmj4cJ5mxE2ZzoASOwS/yYd21dxOg6FTGYs0q9mbVqkAPIBALDb7Cg
DbAQcs8sUbZYb+sKQ2Iif6cGiyRfcfGQs5dCyKTyzF2+kom6MsWB+f9HVOoTvbzh
wEU7Mb7kmPOTOKJi9wTDkTvj72HG4eZC0XD5weJh1+q22qiFEOD1LTBFWVB6Q/mN
9t8KAcWmLB3sxGcaZ971cTrd4tDpJWbisGBKsn3y+ycXUtXxuXR5xmP5Un4WHNUl
h1ktGLeXwQ+6E65yAeq6MoLVQu2ZfDqPse0pX3RVpHSkK6enTygCIRtK414pzSzn
BfQmrqwmqUWCqaTXwAl26q+keZhuYa5zF7sdnDdvl9r+SIhye9CfjDdAUXdAYFXI
44q3Tn6sq/MlSeTCmWGwgb1+JW1SM7yF6T4Gtka2HJKnMiRCpb4BhBt72kpoNWuJ
A5ZeKXxHy56mHP7xtA+ucHRa9msnoeBJv6saY5qvk+TR/0zG4PDymF+kD31xTW+k
iEqgxfXZOM1TUCIQk2ppjiyfM/ai+Qn5AHMB8Vm2nhmTLww6duUYEuVrTYhBnvKj
/0KUQygTXqngP/9GzFfdrI+X5sj0xlcVTixLqpH2/iDwt1PDxRIuFTu3BbisS83o
dUT6aX+22G0oj9CGtCG3sp56OLYjxQSeywTZwj88dXvtuSjeLIeVPSbi9DtuRyLb
O86aynhZYImOUxk0mJ7BNpZ7a8m2EHMzeGJvtpl1xFq338nigeaJPzNxejoGFRLi
tNsta6NGrNipnLR/swKAriRdfaKtJJx1oGKJlqwzuHugl5GQaHgNutMOPm9kORIy
tVFPtdeHEkm63O3wITONdrIhZhmRWabn6xlqfr5bCzW3SJ0xwgqSXS3l7WMXRoHx
RYas9pI6ZdTyvm+mS04HNVinjnCNTDoMOWiQkH32riRvOnNhi6vV6nmtTUb4ebr/
4e+3MCsoubbYvs5ZvOMAQ7Y5vm3lGkQnY4AgbpCbNX7ZVR1PxyY+6/6B87LixQXs
S+z7gFPYTZdnkVjRDFXJE/fY3pyQj0XR/vr1EEguUJjqbjP6y0cvVUM4TA4WCwn8
KUdscN3uTHJIwDJbnuI8wKSdlHHsAg+gUC0BjlXlpTgPP3xxuAUxjmefYiuFjnv9
ZPhinR0cuM9v1S391rN9+qjE+ivBDkIPbEzWG5h8rCwUTd9Ku1UrKp9dwuH0TsPo
bWY0sEBysKbcTaeS4wHhcj5BvJZhTvtbx8T2RiqNpAX+tajHF9A3PcEsnxy1MwNU
1+mGVPygyi1Hd77EfMfxo09Pp2hlmalGWOqnd+RB70D64AF0yErbdZT3RA6b2Jje
cACIEprS7NBfCB3PJMJJTXNxcLq/6tOa+aJ6fASWdWVPdgaDpBJb21bGrbaS8AWo
wH84IKlyPFcJGDHLCegjIMKG7UZFdHNljYToRbqL2N1QpcvaMDeD0SLMgnV6Wypw
WJLaTLX8ZncFJniudj9qtxM1KAg7ukm6Wz9rt5XFLO9+ImF246Oj/UvfuSTV0StK
oUbKCu6ahhPjxJZfP737HwrgggwiN0vwpsAyTvjFZRQRR7ExdMbhBwwuKjsMuALw
xMVp6kA/CHeLTP6siNRUu6rIR7gVAxFAxM202cevgimvlGMVpLJ0cIaBPY/VlXhU
wv6oOtAvId1shXKPeqpBZ1erpdkmMMPk/W3G6sszYV+jciPeUMeiIct/wz0JL9K8
W4l3Yasux7Mjt5a2Bfj0ShpQiVLOf68kBRHZ15860jPA2icjM50YytAQ5VEKDBK+
FaTWXg2083hll6gAmMSQ/P82CMrwTCgfRv1l8NSwbwD9IHfcaIiS3Q+NxQMQhfkY
GdjUZ7QrZ2/ZwY861XORCpaqnb9p6mPwqrbWRpwOcWOG0TAq/Teovf83Z06SQtry
sG1YPaoWbPbOULQsZiUw97xpAeB8AUWCbfU3kcUg4gv2D6f2FxDQR5ScQh62rqG4
g32WQmZ0k7rQnr1K5oCg0btHKr/qeB+sKisnfKgoPScXOtxzsItH1FKa2kA+nC37
RxyaSdkEb2qWXko57OyOdimzM6WbKnZTQjaL8/iq9vcKGB9YSGJCzOgHgdbWbY2x
+eRPv2p8nSEupfwm42kFcUf/MIm5OcsAtuf+Xofo6DBb5npYW5e5mIsXkvshgVh9
ltfZbtz/s1lSK+nfOoedLmyxGb2z/8K82xpO7s+LrNx8EzTKrh5EvL9Y6HmJuRvq
s0nt/Q0gEihwUO/QPHGiO+UrBs+OfGZxcRRLgG0mYj6kK2wT4JtByhsvyBBtoJ/C
hoZMqXVNkOIrK6hbWPAj2nZvGrJEo49WOcYU+u5NEsnJQrKOp/gKrK357GMWG68Z
6PmLZg9dh6fqGVG6SxRhrlncDgpLDtp6fHlujUq2/6ckozxfuLHLoqOIigrSiCJr
ouM+hSssLTTW+0TlHHzELovYbNL0MhKeF01ANUZ8QhgjHjrZjt4IbbYe69Hy9GWu
cA3lsN7UPIP8EYvmFpr47DEl24Qja5zhjXkEnIN7jdo9E/N35+PTcri4GH3ih6i4
rwzXQ+n6mGEiEvzdEXKvaFGLYfFgN/dH8pEPNRpHNJe56MV9QX6yb9Q1uG82oZAc
612Y+YdjMFjle8Y13L2a57Pl4M/WQCbxh6GmOgcV510FAMkGJrp4mzcqwAW4a74Y
fvu1s74W/xs47HlDPoBxoIqvSbsTUdOihZif0b3F5NXFfnKacHW4n7+4JB78HOcl
p4enOZBaFwm26BWqKYpgTP+PHR4KEm2jrSMgIgAadN7I2cV3RFYqT+6HKyT6B00Q
jgD9H8cQwsTZgEYIYGBv7MvUFv57XrhtqDInEAqa2ZlnmJ867gkhlMuyYRkS4+pe
bFwan6hQwjc8ZI5TcoLjcCIlAllrWLeroQkj/R4XQPH/j0PnC3Y8/HR5drmX/+lz
ziViqjumNuQgNIJWsLu6t5Z+wVUF7AW2vYmdXhByOXv1+krEZkppjvpiCvKWxZC6
6aJIM7tVOPbjSRzFsHKyq0HBp3O43PT7tGulRQq1FVKR5dw5BFw47WT1mw5Z1PcU
xpto8Q6kB3U7w/bFrDokyGxqsRypywNruKEdgoQsLEqGxWMjjIjK8akkUk/d5HuV
2GJjfePKd29bf0sKdMa5AukFCU7bOq7EBxyCx2sFGyx4Y67vLiiL+dmKadVTiTqH
kQbUboMsJw4/i4RD/DKzrLTee25gTkPxYodsLP3a+eV3lnX3LQ2mQS2C2o8fqAEP
xSIdVSInKHNWtA1tuks1zpDY3sA9k1NmTCEDSgnI++0Z4oi6YEu84V4vUNePAUub
Xvi7bw8v/8Octg19nLFiWJGjpotDGujD48+smmcmi7t6fZ+6W5ZupthV0+dcstCw
UPFDEFxi2RnMzylld4Sujue2pRdc2Yg4wdZ6jDhTPTX/iwq2824g3VCQnJPsZwAl
Q8Ny7ElDkt6rxIZMVLxrjokZLWYA/f2AyC8zVbUWQTz+Y+CAATv4ld6fm3M3r7xA
d4dp9VK4MX6db0x1KAR1LLU+4K832OW5MC/galAxI+t/+PKplxti81uCdqygrMKz
594V90/gBpXPO0+3r4HSQUiFlqi56wj+MzqxKnjM7eqws89R4DZYgf5c8LHqHZTE
pqWcJHnfVl08wCHXS/nv+PEDdHnmxMHe4kZ2jUdTl8a7viorTmHtWv4Ojc3hp63z
wPCa4Q5v4jMvcZ9yVof3evvVKyoZKxCZKzGd1AP+prkXQ7EThyWDB+PjQq0ZOF3f
6H7oHDW6mSeDnfM23nOWBPwSeqU5AXSfe8jJixnOKjCknOThrohCwk8wzqdGL+LY
9xXXhDde63RncN6vDTZHiKxSXPQknXvWUcdkkx1UMWbfZqRvVlFZ6UPkXTvcLm7j
7Qp20tm3Ceu2j7DZryA2hXV2AKWZTJX38JRqqycX1tKiase9jD8m225IsUv60t/N
NONKvEcO1OS65aiOg966+f6BG93aoc1Yw/L7HyskytOcI3e1EsyHoWaWfl3KNG04
3dQiLVovTE1tKLkbNfuZrlXMqGdAarQEiIkxKTNW26Fw3+DUEEjinOvizdrf0+pc
P+MsH5wfhfqbz5RvJO+8Ok6n0T9GIW3uJTyDevZKmxLS6IbLj6xUv0wdlQfxxS+3
D83b+4taiLm8aoGZXQYWSkiW4oOjFSEreVCLjK8iynKF+mKVMNX/2hO1IqzxA/+v
GcAbkebmLfyawfoTCGm2B9FqEdSyQYnIy2NjJRkbGojhwB0N6efQHthuicpqmCzL
9lvS6+dDa31iqNRdgkZWaYoSPBGfyd1z6IIThks3ox4dLEU/LrV59O4uSa4nk6B1
Xi79fgcH2sW/aqW9z5SRJCLFL6hqt2v3od/rfjKZLO2pJQz6fFDXI763ZvaMO7du
FiQlRUzYLqSn4U/tJJPcBQJ4mGj5A5mE425tIr+QSVKJIGYSGAHL20z6yU/FSijf
FjEhME6k5chTPCHQoH6IZUX7Hc1rwkUQRCELBKAVHUYjT+B9dxrtGslxkkY/Nxdy
gJGzE2CEDR8tUSN7nytnJfN+6xQ5dkptt8idWfgpHYU5khaEejDBaJBuTMalUH98
rj7Lqhok+Wr5BM3kRfWy2ZskNjwD+gIS6fs9wML8/yfjvHIYGHuDa2T2aepLxv5U
O3oNV/J8JhxGTGa8H4YcVbFss/CS3BSxifznA3vRu/AmKlMKdlBQ6CMy2iWFkINF
Ytnl7nUbx6WRhNfncqW/OXvbg5b2yH3N24f5v8WzNTYn6axOHLtU4ksLqMlMu+IJ
rmzRC4imBv4rK5oF7K9O9AB4pG6PdkFquBbTu6D3Fj17upYypu01zYdAWDBqE9yd
Z9Y5LrNrFqiWU01Hv/rjaXbTdpkbFMLf0lpezNPzC/bpfhYpn3Lt93UCjHIRHj3w
mgfAS4BnserA4dNCqkZe8K/OvEI40oOMA6rfoy/CgipeLGTSCgAhP4/TDrbAbdnO
c11uaJVQu2Cbt/jjnGMSL/HkOSUNeN0I7nY6925XpGSWb+Fe1YxnD1Umot8/JaR5
3xJO64aX7bxTZCgEZYH7+aA0PYZNmKgxMs8iVGw1LcXEt2fT5EGjS1m2PBw/ema4
KJdLPve58BLw4C4YWIFg4zi6VZx2/5UzcCr0IUlRJAkF6K+dsuH80XBtiCNRZ4Kr
JnvmYOBkAxCnmYA1Y1e/oQcTjDsXWnsDycnRMjreNHEkfv0Q13piY0+Mbi+iaEsB
cUAN0Y00kxoPgZZxGv4q2RatWniQ53dJURXOkPc6cLVnYtnFfoJnt5IKCV3GWDOo
CuGtFD4BMLR/JE2ksSYEiE6F37e+6aTUhhifUWOaoZwRXbruiban8IoKYy/LcSmd
e/TI6WBOe1luY2mlqNDPgiOuQM58IFcrE1DCx2ds4nr6eU6+syQ+kpu32hTOHVmp
w5Oz+xrfgebr2tyBUP1L3IKp2m2WTfZrojDalmq7mEQLlhm/EAPDAdADclaExllx
1FvLj4dBt7zCHDKY+lLuUA3mGZodls8hW3OL1mnEDGnFvRQ1+ZuWNZVxZ1lihRD6
pZYH+1Q3v+l75FqyCxqtLCTYSb5JbKNoPp58s4ibKBzRYcr3x+8PVJiD1TxJNZEY
t2xV0y1WG7SzzI2/2EJ8HoAhjx6LDU+0LT9cNxoahQQvnQ6JFf6mcmiFjdRcKAtD
H3FwHWsPqiUgBxlvh9G6XqKWlmm+VFYQitvfEhpfVnANvqE9ofaoDqEc/ughyj5H
QeUGBtbcvss6NlZv1eUyvRAr5/sdHt+QmT1fla9UC6QM9n181q8a1csMYUa+H59X
iTnz0sJ31ltBs8nUJEPE4wnqOoAWQGlj/NaJsbH9ucM/QCjKsyryIauHMY2kK3ln
m/k/8Jkr7ayCHPHuomNDbFOIbgoGWl1Oyo4x95TITiz3C7IuTD0ecJBZSSYhNu9a
SAziHrV/9K9dAZkyCs3ZqzRLJ4dCSFKVRJa9+7r5hHktdZQ7aq1Os9vKXQiatMtV
IvHs0xmOWUtYBwQ2isWxl1+9WHvC4y6GRtsvdqZ4X4J/rQOZsjKVolw1G4alU37I
XlBvWRGsMUkce6qWGcfKE5auk1t9Af4/Y4dUuPCEacJvu4aRmMhtvV7xz38LlbWf
snjc4Bs9Ibq0RBOznzDnL6Gpb9ajmwyrgsfTE3RH0F204ddJxar4ldpMDYo80F+i
4pswl1uo/Gi3vkZlL9IAs0SPhAjKOHZxXTGn7cIlmi1PRBU43aSPICpYkwCQPuDx
dZnkwMqYL7vQkfBlPCXEqYBxpSecqNWv9zWyl5ZTiH+8smBXkEo3IbGsOR7Gi+Cr
gL8mJOrr4EPFmDeqzL/fvqITjULeng36wo4sDEmDI1HNSUF9HGuxez7uVb2YAarw
6PShwpMwvTazQt1jtASIzY5s+SKlsIulOunXYUNTLPxkthWydkdQp02aA4zXZQrB
Pg1HjuSKXeGuDhNbUbnzrDVN/WqzlwYSzibj9QCoLikBCpvP9Mn+lp4A6pk1BioB
HZT/Sx3QQ9yVRe4q6qzfkmIlIUl679df8HyBzAqQd5mrp7Hus7gQWmQZPIh7vyP/
mL7cpwVLKB5Ngd8wSQOGZ+d/f6WhNZcWK9akP8gqGIeJ0655vZ6PTsbwC3MXAvkx
dOdcJdVfj/C2+RcXXPRD+HxlwLbuGxKO9ZZgTGSpyvLKNWucCAFU/D6DZvKtHvTg
niIpvopqoxtOa9+aWmKssuwXRhfuH76uzbLndWkyp6r6No4DE3+KbwdnThJKc5U/
HePf01EOc002jPsYv+gMVQR34yPqFkw6IzllFb34MoYWWEegjCO8Tkf2KMGxyeEC
MmRtpSa3UwDlUlIqpXOOiCsbMa4ftKouTUcleZCDDhXjl0yfQWS779MjAVJiy5AS
NCeZZEkfR7RgumWjGc4eI64TvQXa/lLd16Iy2iQ5VL0NyK1YybIOc+km1EDFT5yr
2YnjOrx0HCdZjX36MuMPUzc3AOeMjHg9wNmdg/wJsjRanZgZ4gJr3doPOIrT1In6
6ARjGByr8VI0I/Azp8mIQhryc7Vn1ZDDGhnzI/M370cpklRXT9CeRy8LCrdWl3LU
YECRvhBzVafjwxDWYNo5C0J1T7D9ZTDu9oYaEU5VQrLR87WV1rCv29AH4J40Ybk/
nqajYNRwh4d9t4YuQdZyiVkkOt64JOM2GnF5q68QX7ypHqAOCZAXTyinOQ63yAmy
Q31RX6FDTUfBY8Bv72eYV7oZqxdKUK0otBnjD8YXjbx5Y5HXnY3wl4+hM6B5x+2i
zf5444TF4TQLwZ74C9oIgxaN8nKaC9lo0TaNUO5S18jn1B7pubp3bf2Kkn3uy1iD
+8xSeKmbfAbixkIM0/3Tmkw1zHlIet1pC9bZZ8iKjarcwiGJ/D3p3MgXSvv6SAbj
CyTpH90Jzt7S89aRFNPmRmyLdC4/s0A5Dd2lvQMd5XOpBqhHXSkS35WBNztfjOfD
uP7HJX+pPs3Kx3Lr6Ad3IuW+UiGK2/AuhX3f5mrIaFXZ2IEfsBPzwxBVrwe6mytL
m0SDyvaG+qKSVbM5Zi0OJrHcbgipE4NiZh1jZffcbrb3qXjOa1J/pY8gEVZ29fPw
+efIQMdgEeuJtJSlcbx5rQwgCV18ugAy3Afghhfs2mc3sHKLvSaiOJ0J6jfFoujR
dcbtrLjGKOMQL33hRnI2sm7qVssYQw1T77AfxpUJ99JjMjio+BR6Xi5pZlZLbmjh
ff8xnM2Jpn1r5SGlkZvfcPzfYfuyjVnrxS9Os8P53J9+2ydwZKDdS3m6Fw2nTXsI
I4lpbkAAhb4EXSO26FVTt1B8n4H56z9RIIZKoc1LYFCcC4kHGTOsOyW8FStqVFY0
A+2vlr5ZjAuatyiDADAezfP3NjsJAeTpXnwF+/oo4c2TpjdHtmajuT+B73upPPO1
sou5Wsr+AIL259tJosucioce3OLytGGXs4FiasWHOczIW7My0bU+alTlrjmxZy2A
L+tTonBrqWs5fMpJuvea03eJcRzYQOVA/jta4m208k3ReSulck0ABzbHQKuWooud
dPl/JwznA740+FGWCtkLd7Z658WBbMbs6dI9ITVWvDizfPxQSUQw8hl3u+HUQwot
QyAhvdC7rABXyBDBQFWFXktiZ3c0TaJ8gvi2zQo95P2mzdsrUEU7OVmBzbD71I8C
9ktuS+n7lP1G/ZW8U/QILoThnGhHSgj1RE7kL73+hRCrlhH0420zxlt8x/ZZexyp
tI1srpVFhIyo3YltfLvrYu0JLUr5aExBo3ZaJrIdLA8UnfXc0iCo+Tlpbp9rd1Pl
Onnysx80Q0a3oibahgbV0knEQzl0gRfFssEjcY+L8iaQKi3uGEh55XhEE0KezFqA
/PJmiPwi1cR+7XUiyZRm4718WE/64KoxOji/5F7kC1Q23t1ycfDuUgdXvZ1srEYk
c261h3hHg3mqccE2oUKSpxEO4pVDf3NCYJ6NpUsNQx1psjAiDmPlIj9r3oL3PydF
LD1tJxx+elavyDQZV/WOGJwkS2iPhvV3+jiB66YsGuxVepmwl4pmLUa70ZURzHGn
iPoHlIX/ZNN/2vpmFDzOPP7VKy+eOgneV9YxG59k+tN74OKBWdCsIz9yLNo0bVqC
BKU2Z+zCSGX9yERZ3N2v5D2HbEqDUqhvJYIQnKHaze49+MqRzJLLpOXThsAYyoGh
2yVvDDENatwxjfomPbc/PnO1ekraiH+NJR2AKv7E26nepx5d8OLp+hC5sM4BS/Xt
kqkxd1jazJv012gZYQciQJagte9ajbHbdDf3xw4rw0KBvlB8Q7HahhcT/quOlQ3W
jAWWwA+1N9m4yEu5V1FFS0a2aGF5zUtx9PNsaYXPGHjWaceDDh+g2n3YqPnm7TEB
Y1IQN2A4rOznDwVzBIi+uZ5lRp+MVcGo6kv3A8Zvi6kotZs+DbBqOkw4wcCHV5OM
IRxkwNz6kCO9dspKpY0HeadwXJ/gXbYxXEdiGoCIyybM4JUW3k4T1Meiud1SVwsq
C137DVq9d5qHkCM2l5Avqad38NDiXHf6VVkh9bjWu0Jzv0eJ2NZR08jwoRoIWlmI
1fHECHPZXvzcf962X9aa2Jc0hFbjyE2JLA3eW4G+qyvbRfwGGIA2zjFTiM7hGkG0
V+xverm6QX7yfvkHtfwl0iBk38zQJjjQs5efBiCovrv1gh6oIWZgU8fvzzcxw1aq
VyPmnrohvjSsVpRhqQIf2Zt5uZJp9KUnr7cGYffUy/6XP6vTCpwwF+bVIEw0uoBs
TdZySXU1A/c+aoVduaYjSDSMrMD7V7A74T/A8MeuVZSGkWvNJw/iUznBgPP09o0j
j3dTdvw06H7x4s8KsPVVk4Dhsp/sBxtFeay+Lx6N5mzWxTw4d7Qn52hX824RRR/L
izm/8bkDqyzn3WnN2HnZW0hXXR/qXzWxqWcjCKoheRbCfUnxLmDAb0tVLMvDr+H4
obwN75awotN7aL/jOvw9mbG/RQ1CF0QDgs6kvpff0UD1McMfyLpjpNf6QXzumtxJ
ib/+cgTmPGwWDT4E0judLoSvIv8LFQSYNK8nLVj6g0Zx/6GDcN+Ruz58UsoH4WB3
YmFnh3ZKqwwBjPVx5qBhzxVEHXOF4v3A3+aT8O4YR1lsdj3TjclbQ8dltMUl3PvD
J8iATCLwYLbTp8i2vADQQuIvknpR+WVvKcw0mrmVER5oY6piJsHTtQy+PZ0FDLda
17zWHlEvqCZKbzw2rkqIfrOYpJ9aYvgP5TSBrmWj71wJ74/6yaHvyVTkVEANf7aK
RPupMKGbGoSnnQ1grUjSIj2KEhEjHaJTmTeH7MCCAdaWn6H3+uaymhbPOgjT49bJ
ov6YMj4feWRf4/d/eYRjIL4tK3upuk3S6goWefImgpzW1IkrZ9yyvP9kLBmJtwuN
jSHbWrFmubPsDO/WFuyb0uW2mtmMYABIkKaYZggmXD/eCOKclmeGvBMMUerwtniy
Pc8ZFYcx3CgfwuPb07zsG/i79HFdd1ukk5z8Yv0ehYEBiIpum33wypBDv3gbu2Ww
qRksdClTeppsA8k7w2H8bMQ9ze79hMGsTz4m5D/u1WdQagPZIXN4b1wNZ1w9xd5p
Ek/qTrwhxkLSgJE6wHSr0+bbGpTyDhneRF8RLHBwQ7Sdn3vXF09DK1gCvZ1Ad/BD
g9J790v8QyvSOKjAytzddWsCVFowAiRd5e+CztZycS9ceHoGFdMOiFRTAE9jPPNQ
JTI6JeWwdIF63fBChAD3f/C3G/vIURKCAptdFutKaFdKje/K6NjjzTNn9A8SYtSB
XbsCX5xn0eZvM3TFaKb7CLxGWGQ41F1iLLL6jYNcagbyo3ivT6bIKqjsBJqnH3HW
UTklx4FO/Z7TS/m7t+2mQ0mG+MQeTrn9UJ8PqAk6EWFSI2yucrRxKKtJL0Dcd+XV
1dgzwYQXcGmNDq8KQ+FAF9xaQfXQkX8jJffbTw3fu2Y3Oy1z0Ebmil+/VsB1xMLT
IYjOejoMttVt5ZcOUobf/dsyHb6i18p4C1cAZaMQxrn20DOU3Z9l+qzu0qcFr/2E
zD3a0VcwE7iMwe5NYesI2h/YTVGOS4xrzdbY1NU3UH+q4WL3BmK25n2LlO594xWR
W1ZpDoSWlG0OUAMs8W9jz13+F7z2AMhXJx2DDwD0/KfMPyFpTvJFghGQKRGAenBQ
EXAWIJu/rMKJISo5NE/rVrjgjfGmRH/tcT+pwx8GHunR6VVCdZrDHFeT8XjSFh3m
W+kUP+1zzvJAgSnEktk1qQLCzF6rapB1sC0+W0pNgxiZkKjr75eNkzy3cpqTR8tq
hEd1B0v035wBycswMqtsGcsC+4gb7ikgrZTFsQ6lO8e9NLGq96gOyO+r2UWqFf0i
RQ9oSVOqqdeLTK7IYPdVStYaax10F1SNJDGFoMzBlHepgO2cUtxeYDT53j+TXGFc
LqoRNwow2DewhPN/B3QaqhdvEumVoRX0SzO35HBdMogvD1x95Ra876rRm7ZxVvXC
C4Wi8RpbFmw/uEeKygllYYuzBsKDwzOq1c/Q9HjzVPi479DVITKdXOqkKirNnokC
CdNCvsfsrDJvXQyigP+ocTW0mPuzhfcztJKKkQ7s8IKwxCRCddtqER5qnJerh7WG
XIzMqwF8pYaqmtgAyuz1JLLp5s/rCWLujlmUctbMnTpBU0eKrf9zUSU7iCVWNp78
eaVlUTo3UKKMaOat3Lj/ZcZ6clTlfq4LJix7IxPUO8uCAQGaajT0IG3z0N5inBMU
2Wm7f4lRrkxwVkxC/tBHxhOeTZnAi/4siFW9r8hOZK29BQ86kcSVQof1anBz9gM4
Jdfx+cz5nriKeJRwrpCRt+ixGLgUUEEQgzLG9pHG5mZmRcqjL1tQkV72AbhdoOhr
msbM8vzTK0BMnSTmTCSDkpuahYljK6SX0EPkfChhHuZ6vN61jEFJ0XusDbp/ZmO7
PIb3U+9pNfrBG/fdEgJjadrOBG/0+X3bcO3/mexC0/RFyI52t7JP7dYbD4wuALn3
iUDBU79INLDmwWlxR28dxp0lMc407Fq6z/rbq+yIpNMK/Mc1qhQXQtsxtnolXD9p
bP3mzDmDpylCFwstpzPpEc1SPsW3yS7xuvp2rwD3hVLjqU2K6+/tJ8uHEMnl9Gad
Yi/uYmy7301S1viaPzXCqULA678VZ2kscNyuTADEgyw8+Vct+wwCFLNv5b8c0zYu
fL4uTwJMXF6j2uQ1ZK/OYAj/s7/FW/3pr/7XgKdWdQCUQoSfuDn12i404GzZa32v
d6xFgPG7i6X+dxNlE2lUU8WIF/ra7idX91OCBgCr3bJkPbIsi9xNX401I40wYfiP
hiYuhzBjIBrwAN68xbotm0LZfKhfvebHPV9Yhlj4HTJUkgCW9NS7XzRRTzXhiemv
kiq1etQtjrykSh3tr5DOwC2ZPu7oRFDH1DQg/aNLD28DYdei6rHnQGf9XUKxC6Mw
EilGsoc7yg2ooWfKwuoci4m7EA37Bz96MLPvSmS5pxcZkGWlrvs7yYcjyXMyqNRk
bVQUyzZTqVz4esYfqa8RTMRuD6Bij3XAj8J/XtxR3KfcSoKYab+HoAUSs5YMz7xr
kYvxWfCeesVVpbGoHPB3ejs6mqbdp1+KSiNZvpLYDAn7iocReY5Jg0WNQDFYMdb5
+ArOjOXiz1GoQEsaHBrY3Xi5KF/UvgS4k40Cx8yf/ADGi9pOk3p/xNzHzeHCYDYq
mnm10DlKnYJR6tG7ZN2CL2quIUSkSu4Pwjc4I19e6oHN/aociX2VuuZkLuG0D9J3
G4d5pE7KDkVSkVD6E2UvNvqGdoa/So4o5B57fci+JgwQ+HxhH4p0Um56H+4ow3iq
7em13qTETJKrzUzEoQS+xNCvWJ0Rb5nawEO+wO6070xbGNqhUPPlxT+xfXIviiY+
3xK8Wj1vBB0UpvWAGV612ZlMudVY38pcxOtMDfC19kaVnCG1wTOhnUVBYhRsmRyc
jNnU68jbHM+B5nBcp48gGImBeJwsFKLTued4M2YQHBLH2qr4eqEknp0G+WQu1Nf2
qoG5cH2QszMi3I7plTdMKcwulKG3K7UK+U2ncviXF3X6OV+RIsCABDYBdrww01r2
vHU9E/0yimveHvELTkD246isSclYFKPF4RZik/67HwxuwFqtWrixdXnweBW0fgP7
ynBvgM6MJzyoxE16hkYrhwcJIxUpOZiX7xAhG1cfNX2qb1riU8FfBwkuSwuqmhVj
WbSFtQSU3Icre+qPwFTuwLywS4WR+JY4U1I8IpqTkkMQYaqmOVoHRqdcImAW0L0I
CQlFzD+aQjG4DKGkR5SeK9iolycLQAGgFSlx06Dhnnqx8RJ8pKubopR1u/V1KZdC
7wC4RxiGLk6K/YWTjfhfHWjMdgPrWp0PKJjKdlMNrz3gCvPsYOzbhlNoAfmiJCST
gNKJbwRXESk+nPS3FHXcFXNrBoQ1vexDAmPL4cza/UpY/7YHz/Egtk9Ig/rm0IZD
GDIo1OSr+cwJw3UCJi/O5uoXE8UDCAlPM3Lr02gnXnD9KwlQHEz0zG9EALtLqBFu
FGARls9ftPei64ATdG4zVFUDJXycOB2j/PjYP0mFlWiUa33pVR33H8zIc0Psr/0e
TJY4PXug7BxbJNvCAnWgPAXWf0SYiNmgagbbGynVSjYxLO/Y9CEgy6kjdL0kz8Vi
AAf5VDdO0GO8ENXNjqzMux60qU18n9wBiEasvWjRba1NDq9SiqDQYK9zG2be/EYf
EDVpPgF6ansA3c5dhpOFUokjBQbr7CuAK9VGWqtYExUhpRdUcTnlf7FWBH3jGNvI
CX0HFp+zhr7hCFsXHS2AU7gFDZV+wCLK2Jvaa2RWY5j8wld49o0pREj5L4MLwFaC
Nl5vFpu9bkJ6dVeHupifIOkiYA0EZ6ep9FUvI6VYhm/OSbu9DyhUSPxlgklBSzm4
eIuA1gk/OrWW9W6IWppfNp8H5fb/pOTVQ7ZgBHpI1fSc6vUjIRvxf7MhsXj29Rpy
3y+3PHecv8Gz9p5r1I39ZPwDoHzixCjcT2+Tgxor1Ywz0cZNvCUZ6dunmH0zfxT4
PPzMBmNRsu9Nh1JjblRVEv0448mvX0eIeR6s99gxeyoXdXYkeGz5x5lQc7zmBMlt
QTXK6r7Dx5X7/srTIfYeFSjs1C9lVKBY/meG1loP7YudCL6/7UnQZbPgMViZfMkU
5ME98Ap90I3Z18S9SNuMV0+GwJJfApvbipYNxlvFsZB+PJ7EbpHci2u/hEo7/nFz
TJpPpt5hG4qT4fu1wCzSwA3D9mbRZql0qxlySNlgc9OZV+3HAYEo65R9YsZiYrqm
af/ZB3vbWLwusdpx14fgKJMmbBV1sf2o5J1IHTj2ohYw1w6x2nm5nxrP8kphCy8p
kXLJlyO2vQSRmRbXs9uuwYCUqY9XCsJ+6zTWhBeP/fkatBlicQjIkuYerzKjusIN
2RSuL4qkzBJubMX8notrsuCG/xjwGv9mwMcNH0t1o/ZxuqISE0BEEU2x+yqEjIjz
JZr/mnppbM+HvMF1QG6FyN5TfTGndABqzcYX0bC2aoSnotDJ7CRoSayn6JLpG+d8
3TP7k/wNxIVwPii1HfqbmjGze3OcJK1nWN1PT3ykF4K78LhSVILJkeptpaJ5kya4
ObByKLPx6f1AfFrHgaP25+aYM35XYMYC1RsLH1RFgUYk0KDEK2qvtzXMeamK817F
Z+3lIWB3v1jhkp34ZKqHEUGZdMJsXwIlJPCbuPDHo+hvW9V5tl9VS59fJmpPiAO+
6dGl1KkrkaEhYpAG8+oBM3/0dzoZTdctDaY2LRrtmlpD1xKOX3/uLTUFoZn0kUw4
pEMu70msfvCkdjk6zvaaQvvhmwnoTpZDQ1W75spMsotIKreJZFYRUYlE90uRJ6yg
9Pj1yyzpI1F9ju8P2mw+uBxF+LJWE02KhoDJ1YZhmZDKZJ6MVWUcSTvtRzakP7AU
VerBL1gYIxxznvzJJaLjXaltm04qsyyzpfzvgG2jD2D6hDUAoA8qQ77Bj6unbFmI
1JrwZ09Eoxsk30XRQsJvtMCrA9+eIW8nExQo9fgh9KHFi83N1toDpJPuO2iBKBSF
LvPFod/M/itJFyzPfOZxQLKmfBhJE0fqHUOVIqqotxncA6qyxC8G66ROea/ey8AY
kBTFgVR/0bxcetNhw8IpGuchi6aDSP0JKnaqRDf1zuj99Qtw+w9kJ38g7P9mU6K5
EtifHxPPg2WWLcEBZH1QUqSs5Xa8Uk86s5Gjpm401z48A2QeXp86lpvibHrHdSNB
l8ClryfWieCZlpVJV7DW3EkghINx9GSQc/xcLTH6b3BAYJNRt6DnJWbIYkE/428J
mRBOkae3jX/xXyCqV3pKZ9lzI1Fqos5Rtf/1MgdzRS6P2ouWfCVR5gWZU4AbgUnL
pMPE5u7I7hNwNs+bp2DKOKahaxoho5rVrKjleSbm/c2RdPW1jXgHNOZjqlpzqyNg
SlFgXhHsUsGTRavndPoMLd31F169z4/7eoUWzgjmOSIVWXYytKidno22b+kLJPIa
+pgPrtwX1R/a9I6DWCJ0MtkT2G6KdT/5gsgQp7VzsbTY/LXMC3NiBjQ4RwDDf73P
ItAaLcnUbdY6JUAlZ7/6XRXsNjxhEDwk7uAX2bMWYZgSBpbxfhkuhYVq9oBr7Z8P
ySUsWlp52N+POrLyYFlLWCs4YVqq5HmkGrhtYn6EyzvuqlPG+5bByU9MY2ea+iKY
Jzne/U0aRcdRwGAhceCkoC315ImIMXIEdoLj/UTBw+3sd30Tv4A8bT7IW2POq8g3
DrKzfCM/2IB/Zwqj7u1lM7rfYIrf0rtZMcLzcbzlcDw5pY94XOmm4Jof/CV/LbAu
+m30zEPRVMjFlSPqIMT4k6eyxuiMliN3BXeQmBiDjB7/37ACy9yqdzs9cjPbMQaX
fuQAerZDFnTK7eDRlWTvuDY3cn5wHs311ZUHgw5ZH0/PhR4vskTd+Ihufj3IL2sr
ky/SYSPMQyoZ9JQMUj6M0iq/7WF2VR8uB4xHe+7J20ncBG3//5GRBTTwWRqh5QQg
oDfoOuK2lRm+FPOX5NYeeFDusaKpNYVJuZuICtLb11qncS6ak8zlPoBo3JlKGixe
75E4AcDBk9jAXCUtb3wMmirfYRUF+2F+ZISSSxcw4wtTzJQBgNVVSp6yD2CQzFvN
RrtueliyUftR3B0uUo7wpodmTSMS2Tdllplt+ijWUuCJxZJVG8Dkgl1jwbiJEYO9
uemLaYatfiR+RqQksqZHYvb2UBtQ1qG1YcBiy4Rxwh83uhomkGrTdw/1xi2COVTN
o82osteoG+62zRbIINJcfAinLuNqB+pXrbzF2T5cc1HFCS4C+vr4AUxpLkQMCfY4
uyQocm1g1MAPlvbkpClnIrVrladMT9j5+1bNFRPl1qs1yyVI+mDlE1W1sgYXe4jB
r3BMc9+w+N7S7ddQSoLXXWQnaP8YPqbG+e65gdRKGcXYPC0OegUSfakOKtc4R3+h
cMX/LahlD/Le9WYwGrttr5GbsXENKOxqAEdZK4cNhyaC+ZJfbJxB8iqooOVWdyo0
slHdzhY38Wse1mD5saGWtRlRqF6ke6uyPiNIuonLfd9MyHq/OOoHY0S+GtA5/53G
18uETmDxgSh0Ij8z+Jl/B0yWZz7C9tz+ce6hUS27AmGfXLR5ccI4bOAxMffw4Uv9
V/0UglBGsUqP4aoZiBZp3VyZcBsr3qjeJocHqq1LVCajMHxLUHCitPe+G2a7h3ET
kvpgCsiXe4vaywa2I90lpUJUMYwSo1I2qqS9mdmj+PoyMLZ6+qNVtZzCm6YcbGtX
M2SWqkwOA1w/e44HwdDTk0b+uhiqDj618T4MXaZBHVlrNVYyIKhWvfSHSAE89K/Q
gVyICk3eeDKUTCMKIxI7WhtvRKfLmuuiLZnpBfsXdjm11cxgGWFAVWx49echTk+7
43MgQhbupzZirH1LRRM/RPTnzDLBW5lOdAVjK4BPXk7zE9j+qfD0bC6/4QhT5W4s
Iq7d1U6ZU7i9b33C4GwY8WiihZxDwoZik0X2kK21+/ulKbrYrsESnobui1r/wTpC
EYKIWDu08bbVic1/jkyP0OXHgRMYLXboMNkOJf1gvmCOwYSZp6+/1M081SBW2n+P
Z7k0toRWyRCu4qyhYQJZNlqAE6uXluMzFWCWcU6ee4iA0znTgvIzbAMkwh+d/Wlo
u64MiBh16C3jr41fE/vVZRuoMfkIS7w5uYEKxM/21vVGFpCmjpDi+GJTQj/S8/XH
2MRO15JYKCPRL9LLtuy/d9zG5NsgzupkLCMDwcrPhVGVpty9MdhjH8cwnynSFyMi
OgFbtPFIh5AgibA3RKu7M5zlHZoplVX+40J5xKZyVvOwLf3vwv+9YpDKzw36n9SU
1gFL77XCn7Oi6K38hN15jy7DTjFgsrbPuJb7hUZYmQV2XjIvDOdXvsWEHcYf6/FR
TaG6j4gNDb0tsy8rMf0fuOJBwauE6SZ0paSrrVxWI3fvnLpo6lJZgHCdgC5L+4SW
LwtW1zKY2yuanuRJD3VXSTGadNozA8uryXVCh6j0IAtteeSFKyHf39SERHoMMzE/
qe8W+cFKI4/4NB9gCJDJ/9avufPMh0srygt9bVkUiSXERu62rSs1FiHw9rky9BST
KfAgchkKe4is97dEBxyOmYzDFWS5eKrdDvCp9QLnJ9+QT3t/CMdB6Uj/kERF4IGB
vnVDEEQCk6n6ScI9WghArIdl2UIky8+hQfgjll6kWniHWanA4uwd7UbVRMCJLxeG
7N0BsZSEslsQEf+SnNsnPWQUQyyI8C5ncs105cIgjBYZTIywjn0b+B0kH63TuXhT
n6p7LBOEKaLZrxRdNMRIo3JLFC0E5SyhYcW6Lg8wZfzHN3EGciiS/XkjMhEpwTW3
+0Cnpv8gJyNrvBnRPbcQtrtSwFWE78vAwNg54ofRvAonQaO006n0j5uI9kemlk5J
W5iJi7Su1UF+DCnPZD3ekcCTGQ/waxzIrgpd1XJp8FZ3k/GUxPFFvGnzc0EnUE3p
zgZC/RIeib43Qx25DID0JOPifGakVwH3O7RSHRnXM2xSIjRvfyXOvMnlqAKoWTSH
fBCt6LB9kNq+YGw2DdPAflSClPEgzKTW1LSnYB0rVmLD+6NHEV6yrNqx46c0Xqg+
M6zEv2hziErrqCbP3mrlYhgcrGyJ9QeYrIzP3kTou2cwopiZswxkzg8JUO4J5bmV
QdDSlt+qCwdGgoyabSayWNcXAlImbBjE+NxeMSfExQtQELyTJ1lwZMRsEe6su8WZ
ahahKDFabe6/PfomJEVYs+AXHGPtq4Pkk0XaBpoAxyaOPcEGMYnCCAMYbNjGW5+u
ISMKEUeKXlI7169YBUgG6Uj3Ptn9FpDDVtSkrq839qmcINiDnFUxFdoSNmhX/Rkr
a3yKtml5TMU/oenRbKOVdLugZlGu/bnYXb8zIaW/ayV58s7Ps9yCItMuak19b0N5
71WUEo130vgeMxaZvMRMQffFK95xqsQ0gHy9QNkqsyXdzYIK47zq5RojPzvt71mP
kke6ThQXDXt1/uWflhH+6y3mDlPPU8zdUtQGCVKT6cBOrDuLPr+TmuFSDgdIcXez
5lyrGY61deM/tTmv/9tsjqKpOu0MoxGHnaYbjRtSG0JJ4MZZ+FNcQG7oxbI2LKi3
1YlbnGHBblrX4/sAMIOdYBCfOvdFqv/MSlRD9zTchRSxT6N4Z1L50DS1EuFzIGwk
n14PEUT56xU8OM13EK2XlITpXNZerG4djRdziJv4eoRKj4lbZ4lT2h44AHI7NosA
4WExUrKCAY0IuqDP8HyQeIX4oGX0o1uZsCaOuZajN+Wz97E8vhf6BuB5CYSX9fDi
hEWX0+QbEibto65zQNI8+n54LGMZWRpzkUm0Be7gmUpfml0fYbOucsrNlMmcXGYF
YJI69ZRlq7WVdceU1SXErb/6mCfJQN6GMyoQyHYAinoklDg7NatwOGpQzubBeb58
WRokJop0pZUVpqbHU0oUu037zq3fvmm/H66+i9xSQScJ1olPK08/uQ3AoQLCFA2T
tXSOxZOlt65KtJsI67xCxcKSD8bC/NbdJEkPQkQjsETkcU242PsDHOTH4rkpx9OB
03EvVayjeV4AfqAPL59iw76jVlZ2EubdynYZsmTAD7F1h/01UyagCwFwHCRu3mXE
ItPpKFipesfx9uozO0ddeljOHFYDZKgPOtVmTvsYrpy74aS0kn58eWhxVJkyHiXq
yR5xrfrr/7fwLdJIuw9F6/PlbfgmUaOLDn9jMkY+8q+45x/1Q1rY5vw3EjWLnCkn
aF1S8zRnA2B2ULFLZgMM2dDWtdlr5dirMbNTLwGMomAQwxlwEK4IsavDr66Bguq0
KT1wSr6yqQwSGne2uUpFWPoS6sIABLgtXnNdJXOy56iDhz6zYrBnvxsrgvbERwk4
y/uf4VAYS3yeYsJeL6W1RxdCOrPIMrN21YzK59upcFt6uGTLNoMMwaqHClz7BfrN
e2WnK/UWSHn94Ao3YXzpK5CQAmLMcWCjLOeNvZG2N/Gx/2B6mDA1p3Hcy2YLnhEa
668ZPAbaIyTBjdNz4iC/tEb/pQZb0N422ciKNl8Jkj7okL0W6xfnEarsBotZl47X
gZy+RYG2n/gH60mCHNiFneanuzqcx9bO+dRHErEZ6s/J+eJ/I8qD1w4PSzDgU+0q
8CbecgZai9nSgqe9naWhAFX4NfIKPSy/tZXalbj5xSW7+y/tpl5r7j8uV1x3zm83
Zq8cEuGXo0wRknArtxxgjJWYkVpmfobN4z+lFcMq+lzb2wzrnon5TssV6FxrSx4t
wu4FQhhUcWOpJ7hS8se0KsQ3Aw/6eZoi3rLjzyzYNFYT8JnTtzpMs+Z5eAYopct1
Y6BdAvUErUhKYvyVTzsPRjvjX7kR50JZUJI9z+/BXS3rdcOrtFEVdNCo+NnddcUB
4r/r81qe57L5KlA5jekHPE2laANpF51kVgMViCzyocZo8zeUV0SpNtU/C0pWKVcc
FUJM/KuOrikDckpIcBfRjamKVbUPw4OcHLCa9sf74q0UBiqfm0iDYs8UItWL5bD3
EEfNIG3O5JzW4NU7YdVbJ/GI54XOnttKv8qn/JX8bD4dyVYMeCjHIMsbhvPiiB95
bVr5Ua3P75D5rouqliEzWoX9GOD076RN6s/eAQIYH5AiWkyIaLI/MMj1IAMeiOfy
ffBB9oy2nEJWz3h3Z8WJ7mqm1qxzwA6Zz4Yqa0S8IbCTHdPwp5tHOHXItgyK64GF
kV/JwR57M0TWANoE/AC7uMn1Mcj4UYsQ4XznKTOvKEjeMrUDzJPjDhP/BnFU+bpM
AcFVLDt8M0Ew7qmPJWNqHUXqzvq4DtcoqEzV3SK6Q5OAUuPcA8mBuTd3xnNaPbmL
YY1g4iOgIQGsGsJncMAwF+VKzWEZZd8J53MoZ8vvml8S/7+V/UDf0ZCgk/NnIo+5
ilzGcuNfs01FIkfcRD4VnyPS2HnX55eqqxd1yWMjY6jWv+CcQSyf7G5xzBdwwCHw
oQk0L69qV2zpF02KN/fcE5OvPjkpU5kKghWIL8P9wr4SKlWO4oJ1sR9T11LKEtsw
W1oV1xBKxG+LZvnry2+35nCbnDJvXdm6oJLM9bHmFkq+fVaDLkoiPyq/O5JVyJh6
9TV6pvVk6gZHi2C5Xia+sJmbGEEtTUU25dBxF97jCL9DP6dyEJUBDjiWPzPxx/Bt
PWSVpX3tuU6pKqLFoWDUj2eXBK1jTq3htUviIt1D1F9edAtvhX4e+4ba7W8rwVmL
fgGea1dsEZwht+iVe1Vr86zY3J3UFBN+qDHvEg66zZ/jM4e4z/oCsWqOF0yY6aUv
vyrp7YNutcyVygpsTSJKKgm1UvmQvqjy8K8fQzfdOZwbca2uujJhEBgbiIGC3dJ4
vYF/vmRdmFJ2AJe4lQP6UpqjmvYvV1q/3QdhKhYJefUpMMrDjIdRwfvLQ/oheCBF
XOaBsazufTVYIIcxk1iMAg7LfS5yvLxR2+t8L4krohNOFkeKszwf4xSDE5wZBOrB
dIx9iQ5KcweZuWkATaUKK0neqVuF8ZQmdJC+6U7yURZMk7BWYhxsWJLYbVjX8VgC
xQQuIRSAnyaimmmU1VpbapWT19XG/zo5Hpp+Tr8r2fbLYq3GnDs8Thfc7uMnUoUw
pciV6rhUFTGGYg3YgIqtpAFByWTwdGZfzHzim+6VV3LViFqMh2cXnZahdH9UMy+J
YT2kRmwcb3ARXdwb5BG0mf3I/SHPhhEUnhPca6eSggSO3yJFvs5KE6bMKiXYodHj
JW+gmnpScMbESSBLVQZq2sef4ZF7t5kw5KbbYmsAiCIRNiAmCjXjCfGuKR0OOMxQ
Xcg/LsIAOlIYwpFYB0Mti05neA5L2cYhhKhT+b7BDgi04/tOHYY6//ubnQmHUIBi
DwM5OVl7JLH4QP5T6gVq1kD1tcjzmeUm7iQopzzxeKOAts3/2kl/Crnwxk/6X3Tg
mQvJQUzT2Qu/EQ+OEW6ZFNDyqHRi+hYfaIxm/5iKgu6/oy6O7x0KSZ5Ue4ZCLeTc
CQZQWOmMCEaOBRWDm12zG2hrCYsmLTl55xiqZ7YBbhhOQy5LsgcEH4owdnFWFOlx
ld0H6EAQvLdzbn1oHUuIOK5hVnzRFrq9bvcJfqwqVHKmB2Z93qBIOCfsKMggL8NI
lZKc5GqmREVY51SeRYDdmbnIxlYQxja8R0ZUc1I2G6F2367nOraSxSGacz0GxO63
wGKeFiVrj2j42UEaaEpOvrwz++9MdM1GMaVtgkxexA8OSbDpKoleLIGiY5d+aTwa
hQJhdkEE3jv7fwOi2noF8h33PItSgI2ZJdBc9PQk3LGuPya585iIcH+/f70VQYEx
0vqSlyQmIhNdQ1nb06CJnWaii/bDaTTmr4XfxSR4UO0PhQumFXLVdKAPvXLEgGLi
msZQWlXjP8qv+CAXClhuTQQnsq9TPzvO1jboY7xRC5UNgDVgA0WMRU/ifoCC1YFc
5r+SASC1kwoxRTXh/AMEJ3dbkFv6gcR6Jki05Ku3oUNmIU4dM9FSKcCkbDiD4N/U
ETvwSV0HCXV8Cou0Fy4xASxX0LGfAT2CyL5loCV9g0ZkmVTbgOMGiayAhN1DklCI
ebH0XHPnUWNSYGt36Ao+ITSk9MhyUoe5rICA0DLrrbrAx/Y6T+VxKP1uN7fSXr3B
QXRKQP2b6nHlAdVrBxFiokqt/CbovQhnu65NGr/94pgyK/F/54/lU+CB1UCsX8NF
I9o9KOuF+HqxwaOsBll+So7YDNAugMt9nQHqzyenkG764jGG4hcqQSeaHYS42Qg/
bpI2kbDxtYm8bpqbu1ZTowRLT8Xp6g66ITksb1IBfjfIbUVpCehg2ptot8CLb19V
jBW4t9EDgfbrEajEIQiPPfArQMiT94UXqcB/vu9pLCNwFgQ4NPklTMzO83+UIP+i
xA2fBkMzPcSmU2yU5rbaZx0LF9vjYGp3q2OlMPO1PolO82Wwj3ddKo/alvVGq5gW
ES8yzhBNd8sz66UV3003eYG6gu3OFiENf0pBOIJnskJY+O1k4QcRUygHvSWqbhRQ
dybr+13JsiILcdOE6PPyar9pP/VxQdoK4Nhux02sGrbMD5yjUoZA+j4mJe6DCb9j
h/LxVUNvRlTn3AXHJbNffl+MS4XdZ3yX9WQ5QN8//2gMpfRwVfzeLOH4jOFtZReL
umjlwAtqXwIXmQ6ZqZ86zloaJvHd7mte4sF2qAWKfI0skiT9mG50L3Pu2kN2gKhv
hReIgRixx1/6zWZ0KuL+9OMBhqwjAKuWVXE3ug4VXxErixlOhDJUL2WCBwuwW5gX
MJDmnHyEaZJnGNZGpvDMBk4SNjeq5C3Z+Gyi3YAYz8FYPICGmQWvEIka9WiJwxe2
18Ac5LM4yvMeYB6Q7hk0xrG2ucZdXq3HqfIFg9sJYgqcKJDA/xeE6P6vRVWuWauR
R8JBvx0/vniTNotSXsxdYE8IZe48JCv3G8lHjed0FLO7mk4UR5Oafj1vODml9yUd
rJYCgy6VkxnumW/XsGujnMCOwNj31qMaI/T+xqUldEY3DrfvxFWzsODpZRyqebSq
rIE9ukvar790qy9mRHKItXJkckhIgJZyq/rNm48Eyku0sgG7pUP2/hHPgTJAUDei
YVheXuqXC7czR2H16br5g0+nxAu9W3HlBnra9a74St4Z3ffdPV3maikU7uOkqeAV
lit4NuBgZV1Mxh8XZ3fLf+NpYhzvpndyDTlY4wWsECETo82FBAIE8xEvYSxcvjNi
MQ9ImPvsTBCfNSOWwVQqvLO0KozmikTmwId0z9wX781FmyjUtDG+C1TKvr72hYW2
WZarVX2wMoNfOm9boR1FEc7jPntfDP6zBz5H4hzB4R/geHHnlOuO9FksrFJjygFR
b5Ynh5cdekBD/yk9tJ/cZqKVhlEV4d4MfVmdVVPsAEx3dpPefuKxV5ISuJXEd9lW
pJB8GiBwUSD2A5erHRKW26UL5a4rxn25xeripnM51lRqXP2Zk7Mik9bcxiMkCFSD
EmlRRwctO2wHTz1i0Dv/kUNeGYGsOkPuJY87o+8Bqw0P4gSTiThmbbbwCcxoxUXL
IV/ReqehMyXKoGrUibJOA6Y6xpOkLanWuQsrzzsCZQR/bg3I3ilKpqZiWIpWWDMq
1CyKaHDh2difIUbOJhNt3b+ierY6FzSFpu76Vtjlfj13v3c4agTFbbxSubleBaSI
TFKxjuUlfXFfbqj3jGktIF6osWiHJ8Axe8/jZQy5yx9Jdrt3ozXmFANi56JVS56+
Rcg51Z5966fUcNnCxl2+dQ0NPWogsY+S1aIg2hPAG/7tqrFYeFnucVRBsV4iLOgD
+Eixnn7Vq3g8ZjyXHBlg9sQpYLZDM1UvBbXVF6rXD21t5HEgzkp/Air+x+SQerpl
zm1cQB9RHHJKf3ylIGD7Sj9KqVnhS/kC7XEPMwCuWUp6OtYKc1cOamflIPmPJq+N
EdwygCixSKqPeSnfnqpd3YJM823QTMYJOv0oHHBWonL8wheCHaXfTxNMUyOsCYpi
ZgiqOfRJjEQkv29rrhX/O7Jubf08kx/P9sJuw58fB3MCCUx5mTp16Ar+Mr/eFO7K
lCBZy3GCA8nW/8igimvHXGzYDn4SkmMqjR36yi7TFKoR6L+81d0Jw/OoHvZnz5D/
42IEM1BjkfP3I8Is0cScKx7Z8t7y81NJ4dT8+ds4P/Jhjk8MoO8qTHN5C/uCXcAu
2OsO/ibl/XXjdamCN3cJ70ix90b+IdMx18m2gvaBDXnppFbIMfMMFSAdkH1tmzfY
J1X41VBT+u+SrJRkSiwFPI57PYvP94WcEacjHP6zmnMiIqrvEnkTk8xEFltDZ/pD
atPgfXgEOJbgbS9t/CtbFEJ2uoRCeBUHKFqZRtEul2LK3rpWARDT9v63PvYOYgvA
vzDLwHwJv3RRvXLh0UvQD/9g9riZwYv7IgqNbBNYFL8ln52k9kv0WXj88yc+RoXl
2tHPqTYAAt+yEtYyrM23JMsjvjboV4jbDm+dhVWJ5JlM2qZD4OsEz5+QpWihX4/W
mRdP4/FpGFHq2mQHwJW9l4tFu9ujiGiEGaTfFiEd2VIUmAWwh/BcAWqufWC3tGrY
KFCoO0rUm3ROyF0KVfpiXqAwTwXMrA/Ii8dPscS+NfBITg48m8/Vw6hBdyNxinXU
0qymtRpWQbJYr7ek08fS7mRlyaqyx/OGelJj6fOciQie6Lv9GJ82DItwRNpYBaoo
nYO6mZeTkWZSLAToRwHP2A06zsGSb1whKgEniUfrIMvYDr0K3PxzbpufWPKqiXDc
WTQMcusG7LWiCHnntA8vyAMc0F5AQRXkakAXNEY2s7IKHsUm6SzjTHCTrunZ3GHX
KJAvlk0Q3H3vTCpGJ8E7gZedAWA87rTJCGe12nCDFJ9pHo/SSaZgB71KFJhBCzd6
l3GOcnAmuOfBYCXVHciasQD9lt2PVXt3ILk0/AzqaoT+SuOEGVRMq0c+k/t3aAEU
OHDUF3F3/3n6PQmvyh2le6N6LUXhhhzE2W4mNVfoGo26wQagVGV7ZhY3XGVXdrf3
lv/vN4lBr9nZ6nXUXgTmS7Iz0n+eQTbrstXmP7TII+XRM84Chgx/YKJ5n5kNEJO3
a7Pf5U2ZIXs1ypvHVCSZkzRRxHUmlvhc1K0KPrrI4t8bwIQ41xI96IkzKvN/anoE
c3Lw17EQL/1ohus+sb79hNdutU9pvbhqBIyN1hnCPpxNLJukGoV0FybalKXW6Bop
YHgUYKzZSVB0OajzUmhi71GeTZ1xbuKMCvI4/HTdTStiXJz4tAu8c3Jjl3D3kdN5
eeXdcfbzIZE5X21noSe7bQDFFVT11oEHsdSAikR61ltZk95ILifRJMd6V8eQkehW
N6mwQw3lIN0s544KDu+N24Qrpl7VOSX+Tk6G6dCIVx+RMo5GrY28LcDds4vKoM1U
etISZ45PVfBhvyRet6d5CXUCKxO1wDTBiiHwj9YCxt5rVXdACVuurZkMIkNy3lOb
rJFPstNnv2jFA3pqGJKmVI5ZbCoIAVTkBTnqWh4KVhrYWhGUbqejhBCDued+idC+
kthVYaqZnuGNxJ22WbpP9Romk67jOmZ505I4d0K2ICD+GaGwXyL6/VynTNW1HpZg
Wv2IiMC3gsXH3YcTnzrEPBcmF1H4TbgO84XnOcoysfchWU1+b1zze4QgMYVtkhHB
NCVpuEKcCeEd3hYMDCWLjf5w1ihokcW3xMjoTwUL5uoYKaUtirbiicAHt3sRBFRU
AaVayP3tU8bABBsRMHo26PC+AGTol3SReUFrfJZd6r75EcEau2SydTHI762SeS3n
qgEx9PdcmS+Ou6Lby3Nmf0Us6mvSVZabDO4np3lX/8qIDlBgA7ST6Dz1XUWq6F4B
39bOWk0EBVc5D1eR2YK4MjGN7EzdxYdaLoXcwPh+EQbmnF4Gbys0aksuU43BTORw
tk5p5QHwhTC9/2JpNvX1NVil4Ug/SsYhheeypKd/fPgJ5R4w1EUq55NSYaU4r8OK
54U9zXUN1bdrJf+CQIwupEQ5hEOM4KLxi5iSPXxBBQ1jaXw9xG8pf83+GXB8I7U/
4bEdT1i+GHCMDC1kSQ3CtkPEViuNGYq85xw4g6A21zCLFVOyTkUMGgwVXaq1G485
nIUd3IQGnoT6mNSzsk/NcXf1vBz9Amb2UY04dW80a2y2xNYtE8G/3Nq4JhSg3ulR
709v/2w4cVtYAccLiaFzV42878ec3Aizq/tTyN+1QgkFkdkmSvSEFHkFRB1nNXH3
AC97+dCGTbqs6n6LayMOiqo8gr/D2RkkqwwO13Hwz4hNysqtREqNfmwnc930Mfqi
cnoDTj2EkXg4iH+aMLd/cs/G9y1xgu870NpN0UIVTvZxLVxNy/8cB5Msu+M3P3oC
jcgzlNv3q/5uWAhaxxRMbfX6b1+L5eobFdXDrTo5V4jgPHMkXqGEEY7XUSxltYml
xi1WTJs9KZUKLxVywHzmFOgTd5C5BhTk7R5/Ozp505x/h7dtuxRcZsC1HI4J/mWO
NvildlBiDYIk0EsBYupahBJPx4YulJFVYTJpZad2VrCezzs1yuw0CyoABSCIY2At
7cB/r5UrQ/wF5ljvifdkVFTNvqpaelCRcl4WMlLXb8LoYHAL50UOcD+WSCAZJuz5
MhcOZSnn33ik5TyqSOjh6JRg6AJno6BshJ63tuz3wWojSoPFJwMxl+HG7id90T3r
qBzne/jfUaLn3wVWdgaqrYRbhHY+My3jZn+U/37/fPBZUIkTvZfAQziDdpqN9TSu
htSFVozveL7Q3tAi8k+IhKKs8zRhmtS7h6EEDfIaQA4AaGiBMlGfPU+dGhgLZ9ku
1VkwseX14P1IXNpilz9qKVNIMu0nMtvZeBE3VF0x+RBl8nxfJa5bVvP3GX4pKCnM
YqSTSUNBhw6K33iwnc5EVrCrPsUFNCJ/sfZR1D0r1ZznbpaXdMIDWGXPAm/mEFxb
H+LBWXFHxSxx9+QLuY0Y5h4z72ErZj2HpMS+W8UwQ0g7E2SbsjnVLYFsEVMIRbt8
aRZNufdb2LcZGWaQ0INItxCd6wp3swWfEsE5lznejxY9+57oe0HZjdbVp3AiUvg4
eAbi6Z48hn2fdsF0cUKa7+ZzV7YFfKLSa/1jBSg/TNfORSxjtwn5PCvawlGZm0J7
fCdLSlhMJbCz5r6MWVJBTya2yZqkcxAilp7O5frcUR7m25JHAasnTbbO+zZrMaOQ
WChhjeldFeeKHxNpCOiqi4OOD1gbk8DJQTkg4yhKwXgVzaZdd5Azf/7X8s3uQ+tE
DB30rdX/nzZ75GGWK25aZskVBtCZgT1uG79GvpDPiIrALIc/V9U0yHKMntUNP90C
UYNQFwk5Q1dLAvUJWg6z/knkdchJbmeG/o0YspDkzJxh0CZYEBKgE+mth/pQcELT
w0nYlKMf//S/hsBjErDi1jKN/ZjTj2Li8sJEQaVnjDU46OqqgUf7kd0vVAKhFojp
Sx92n7mLo+ZzYctlIdYV/DF1O5BOPR+vGs2+1/FPn229l6MQpp/3APsNNF1e5Ji5
S3Ck2qCXvzwMeuQkb5ECc8ZYfwIh+Jh8enTF4IzhkwDSVR+qL62LQsC/AkblxtZT
NSCVANXxFqweanBrblrZQ8yeGPyYXSBg/ubVqIrf+A6gTtD/MtnajfMbDf59PfOI
XmOsJ60PapKQgcZBvMB1Wf35cf1eScsuJzHmTNHWud0KlyYV/lJoKeU/Og37D3pW
x35T8njBr2NY8mbwrS48GXnQMtO/u+qYwt90n/Yp2y0tRgbYPZY3Bwg28Igd5zRt
DpU3mX4QyT0/bxgy9cW2bDj/C4yhnEQ82K/XAcEQsLvyV8udT3IQlYSsIRgXg6ki
6zQ4L/Zt6WnnaEEApoyJZ2IxjuWShFpkTETb4DJmCQeiS9Eg6UI4wGoIGzGxepls
hA1swtsYgxJHVf485Dp3DfPcgCEZ8DFXMH67HlP1NvHTYgPXaUHRDGcMEWrkt28J
pbFzvJtakn9LzT85xMqRfDmng9y+T6QTu2o+IPYlNCMIOTjfjpanl2heykj5gPlE
+IG43iKkFHxd1xYBJWqbxiX3FAkSruVszmfot7vjVZH7G506hL9vhxaBtkCo3gN5
KaMRUnqCqzuBAD1xFsVoq4SjuuRq5+u/w9SmGnl0F7cTaDYE+LjuOSTC24DFQed2
uftHW/38zCAJPs1Prq15LthBXrmh0+o9H/ysMv/IwDRLt1Tqvqd9tl2r/0sNzXJB
KEbSI9MBz1hTaHH1uxoiU98dqynyOEwqWO/JLMDij6kt/4tr5hz4d6mJ9gEScrH/
NUNzmjeQt8wYJU3kJ/qZWEbZbN0wvByBwOKVrkQtJng+H9jMW3moDiQydEtTTSzS
65QQU+xnwooRb6bTWLlapVAIITT3/TJfnokhm6AxiHBfX33wu87BehOJZsG4is1k
1/GvlAM/t4Gxe4AvMla/Mx6AvpUYdghU0J1uPaMcC2rh+Hxh+QrQYVsGad21RhFq
kdXJ4eJQewp4UBlVwwRtUM+zvKp0Zj9Z94IM7y1iY3RWIQElGj1iH6mEkbVucYVA
YMXuqc4jYoz5owIJudhwpKOeHzCHdXFmaj8HH6DUnfjTei3jpsvryUsrXzrqRmsx
TAvvre7nVUlRu7G1voaLdBZ1C482ci8O1qgO3UWSejXK1u1tc6Us9TXTy8uHwaHw
yRRiD49nbMKYf8HZX+5j5c7W+tl+yxN9U+AYSzNsggTNQeP+4rV3ubwBXqCtJir4
m3mRtrwpJD0ivAcMQ1SG+6QpdD9QFbZwWg+J6Gcd686tAIIhpnqluUqzJbHWegfH
DMesL8+ym3+pckBtTnQsSuXuKvbsKtOkah1UyuPxVvbnq5kKsRgSo8db4XRM1Z6j
Urkyzd7O9pBRp1fooMX8DpvDACjxQAxR4o/hLRcNqwqlZDNavFd7XapoxUMOSz0R
TUKF1y/V1fw5G6jWsrxYIfloMYD97ePXb5KCD28GpDn+NzDPqxUClJrNATmgf0Bv
4HOMGDsCKyn0t9M6dL2uRSKyZsr8e8Vq0jiqOIAZqhsSxwCzuBseB2whv2zLuPtn
RrGt/+cpYnuts+8GN5kasZwTaB6aB+9blOyMaNKhERVwG8gn0JnbQu6oIvguTAOj
E6oJVoy5CXHIZS7sxM4NbVS8Mpg3IQ2TAxLxMxkLChHaQ7PmFPo6wfOTY9BdsxA3
LDBNZrQTNdCR0fx/HZAFMJ9aZRiaLuj+LzgLedG78cZUcKrPsHysBYGe6bdr5V5f
AIEri9sLrgRrlayzmECgUHH4A5VyP8UF91qn8+WvmvM3jK50CtCrKJoucT4tSZrX
NSHRU0qrdRXmnXefxJSxup3FvJNKrjehtNi3VmsnaqJxxvUjJt3E/B90Daniz/Bt
2kEjOGEOEbIJS9G8nEokXA7sF4cBIQAvU6ZKLsOD/ugie2Fcb4mi0+FGYbFns0bH
gR7Z1rcG7hI0fb78FPEQx7vUre4Ae8ICYctxz+jcGgOQ3jMYIo6AeA+m+i9h0Ace
enMZJfx6/v8mA+z4SXPg+0GzIHwSnNOiTKaAoRb9vIeNfWvNmwWDxwbU0e2Hnf0F
zorU0PmzAaN96faGzw8hup03XFvv+EvUJXOscpeI1wan9Zn6NflJvJFqu867WLkS
eOGp1o9sLcX/suPzHikfaABH6gkSMOEDo2sEF750riwcRmQpcWPcnxm2UYYBdF8S
v5xHqkJ9OiXqji61YFivAZ5V4YqHCSsrPI0+Gu53Wjhwe7kvPFnKJ0vcngZvr85F
vorrqPSSZOR7ZwiffXBN/JoXszi8e9YCpNkDWhY/oWc+U4Mocnh08y/+zQVTvQzu
7zaQcDZlcZuOPiCvpTjYC1gmsdXGVig09RiddrVU64nf+Q4opjEpzd0Y3O3afSTf
FBvafLFcjnVVO1LXQ5RHTtS4FSf8olHxnZA90JHOllPsaidxJLXbdX/w1Yr5A6sI
N2VWLce7JMOV2b65/CP0A/XOCv8NE9zt/8VVcKEjDZFYWEcE0ryQ9FSTftMogVOL
M7WIGK2HMRVv+owGA1PJMS8HdIfrEuXboRnoejas/cCyA2T7OnHvSbKyktsHRD8t
9DAYGPSZ0AmE6BzCvtYnSkuvK0AlJMGWb3nK/42rO+TBlk2PP6f8yOHRYnAAyTj8
pI+rwmKvY+2nO6+2KSo7nMb/P39feTAfXzTkKv8xtp4gUclS6jZYRgM9qxFb2O2m
/bOXJTX9BfVFxrh71LvLC9XtCSMu7KpUfxpq7UyWcqbnejnqG3dFxUW2przuLsyj
W8uStrteTgXMWXsb6fM1DvXTnK24x90sD2IRIYJ2dWiRP1cgprbhMcGxd0GWIzz7
x4uE5wGouj2mTwv7cuSj7Oy7mx2d2yw6ybGmM760mLVDr/hfEoXHY9AmEzSE+bW5
OHOkXj6NBuvt33/SzVS9FwfK1PIry9hLYURaFciKBRV/+YHyqCFvd4VCm0wN6InK
6kcd72LFXI5qOY0v4bLUJc/i7c4eGd+LgselJDj4clboMWCYaG3eBJ8sLX2TXf9U
vvT/vaMyW5QwYkqttATGYvoJFjB429jYEFKuWCP4cC1QUrkdzHUPeESHL5BVh/i7
qEpXZv5JptwZjVtTARzmR7pG96S7WKVv6V77yIfck1FlVOZWnyTGd/GLNdXZUhH3
uQ8pdElLC32mnCWNRdxMZjVodVGvIXnRqfTiKpa1ssgkIputxM6wjLCjnTw9M2uy
Ywup2dsCHLyf2UIJw/+Gdc6h9ncLPBcWnEU4twB3VtZbvsVC3JCI18eMBAQQ9hDL
+aQ/A4wVzQ0HJ4x24DgHP5XXgyRvkwpF8meybWZQlH7FPj4sIYRAh03Guq6sqrYh
ltmvZ9G6fn7ju/5te5E1w76/0d+sttnXX45oW4c/va0guZuVWMzQVoUJ/lG/qEKT
bfcvCh9NEqkCmGTzD3WoXiDm7QbiwQVdg++ewchCGHkxzIwJc3MW5k42xvK7Pao+
D+/XlDLq3GQmtZFNELlKNAaFB/qQT+sFD+PKa3IiaTadfNOfQUy1TCVmI4tsYhjl
JifpJmWj3J8InFM8tx+5amrUupnCJRbc8OFaeJvilYoVyL1VQAdokmfs8NkSgDTT
ElvATjjvoPUtQx0Nmas1LjzW7aQdr/Luz7Y/n44R/n2Y9tXz98fuCNtw7DMNZ9Sm
MBP1Q2DzRl2CDjSGXWwy/cshHVVwWG9EO3tIruXuOGkA2eCIWlxbgWFtZfnfFILf
lgmlDL9OxTFTmhH3GHZQ3EWHnawR6bMxYFjcNmaL0my/qgSq4hYhkdYk+egdO9O7
pywrA4aFPCEgCKeDC4OWUiFhbiBy9UhrJXQtKz4yqlYyQwbp5tXb9qhUa13z3581
my3Ps8zvsT/523Eh+0FanYbWEZiPTcs5KOVirR9g6bBLds9+kC08SL8fsdKbIahx
emo3q+jN/XpeCDjvihrcmBmL2DvI4bPURN+79OQ4G1okbAdXzWQpPU6Tnb7bV3FH
Cnm30ww2PFeHY3SS7/C72WMz9leEHcwMoP0l58jBSX4w6PNPPRCtz1lCx17niYM5
VkqNmcIsbHI1TiE/imsZzCh9an8UQJ6ZVm48vaS6y5aYRqvRY1doaPTLLuOvsF4M
/6B7orBvnEKGOmSKpmwCvDCVi9r9kXAOmVs3c7Tw1mZdyMQnJKCukKQ++VCqFfra
p5CFKZFWBVbKnpyA2AnF3+gUgL3qgVHodrmKnTPstYXYjzzX16mIdPbklLBD2T6w
keVFQwwpD4fwdJ63bWHRe0Uz5iERi0C5uMhPuGYNWSGLYK//bb7lZEbsZwX/asuy
XQQGcySKzz4WRJKRYZ/UUppSBXpbY9bhHLVDYWIGOkK2/abm1yx7DJG2oDlrsfzp
bCBa+tPxMfAZyy7SwrGI4JghU3/3SqqrMluehEIeuhkwq2VcYbgFBUD13llHdJIM
y8OJnCrqS0kC9V0J93u0wFSDDXu9RbnGqbBMhKcUeNkx/aQzNCXe+yIs49VIpL/O
x8j8/6dWUcPmyDsIUcAmhRuMCM+uSOgMgPeqU4gpnZKlEsxmxhga5sggK0m9hZV5
nRxTYi8c0yM7r0NYr3iyHh0XiKxFxEUs/1qzZvI1fmDYoh8nR0BIH5umX7+aWx/h
9ylynmGcvv3Xb4TDcdwA+ZgXowVAmh/U+9ofeFT7p5tHS4Ba6IMM6ooLpBHhsFj5
0pjdRUVOVkeNyavUlsHLWJKLDAH954pIxf6lWd8UsuaUwIMOp7SrhwMMc5b5TTcx
Q+KedYvl3fvYXGdWZ6gp0+JdCNY1/pzqAJGbcan1M/yav1g/lyyH3W4KGEN6/wRm
nN8SJ5xa5eXs37MFNZiKKBRSSH/pLoYZ5XfePBQbhvPJNm8e5qoyrUOOgt0sU4Sx
3WGiWr4VLUEYqdUlc/rE/DALNFq9/Wboi6aJcE662qEG5rJLvDpwt4L650Opafkd
Nd/QQDV+4ZfG2s7SDsRkjIZImtLpH5K/NURRleW9Gc7rMgMEMERzN2AIABegbXqL
uT34cHU9HOMWDQrVnASzcH0ICH1x/A+WEydc/XhDe8Cug4UqlfyBKhQdXj0s2+Rr
0gZwW9DKjKAJrTPlX3P3Y3aeIDEdwH2ivCqY1y7vaLerMnotlYLWmLBGuk+nN5qs
bMvwDTmwAimnD0TdduMmeJdLytCBQQdFAaugGHGwktIIFLqmzXtWplnqg6Mx2kHT
flbvnCq47MoSpqfRePFBPSeQQgtqpHkjZf3K6uzs9pUglVwh9Cji1MZZxJDELdew
zT6zLm2QN10qB54pffQhPFENOO7qSKolt5pwq32zBihiDm+e9ncmBrdZQcYjUpiF
bqV8UVZ53p72SRAJ70fErVxh8TUyccWaMlT65imZkLL+2SHkHbWKniXIzphOiuuH
IclNaJ+7O104S+qwj8jyINGvr/1nH8j72yNmag8L8mt79+k5/9Qc4Vo0RlBnDTy7
3F+bggZEokimNPtbRiBlbfSxARjFvQvoxtij4GmzmOaF/XN5pRPlZ8tvoDrIgseP
PDdqRRpaN/R/58HlHsvphwW4Rg2gYfPswGsTKRTDGm4nCFEYWemFJ63rCCrzH5Nr
Im5VRDdxfD+PiB+YZ9W9mfLYqMVK0QJTlFN4+plUwp0ny27qNBFEccyMAEHmoIqr
n1fdsvcEh4ZY8c4MAoAlSPimnFMW9QbIQ6dAfRJig0kPvg3NBAsmI/KpXGo4tjPI
su2AypefrMVL2F14k2B0JhEf7YPW4xQ/pBFXw3a0Hzn5p8DgwiF9ThYG5F3DZUw7
gTqnFbE2PzcUPuhKzbhZfPpJd35bSpjmxmmG7HzQRU4moSexM49W/aZXr3iJR8WN
f//jA8eKYcHcqfQa5EPaUsUEC6vqqoDmfI00P6bovOBwyVYJrZ/Iv/qMnzg+czlz
lF8Yb7ZVcP/Xpo4gQ4fUp+Z4xi6wy6aF7blOTCYCIqO84KGYVW9oX4LPsFo3chwH
wpr3uCuWg3mXqGzcRlir56v127RM/VR3h6JwNn2LUbhc1p7gjEiBHH24skyBYQ4Z
jTsciqIYokgTXUJrUB5N+lqVZobqik9EXQnX0Y5cxOqMMuh8eMBc4eI94nw81P9v
G+FbknDT+VhdAr4kT5G+6bt7ABeBDhBwy0W/CK59U6JJyOktzQF9b3wCl8gKnrVC
T9fgkJMyFHemgJfkNm+PDbV+BF9ih4IwjkkfhrP3DC0M4tbAfVf8x0IXpgQtDb5B
15zQ0xFZkvPWhY2Nc4H4oNbyCOa1Q7Z6M8kAjhZFkkqOIJfZ2DqLYo3tTxO1mVK2
tqqWN/ksHyGunjdbcB42p+HkxsnBNZUnYPW8Jyis0x95aevkz28beGiEfL7ERP82
WM+Y2JKwEAP4KI0AgUvPKZxGL7r7QJ02EZ4qD3a/Bdqf9GztJTOW32WmTbXDzqk9
d5gMhpZ10m8sXYdE+6cY3BL6qBMBuiQeqoOLK37CDQe9HBgtC0RKBZKU+z/tMLud
aLc7UtnehF8VS+YSWc0SswB5CUSYp94/BcDdqiLoIkrfejRNKJOGpHYOuGGIqyZL
BpOx8ZDBQA23MGBoSRptLAjcuDK3FSICgEodONwt2agCMA28tTPxre7f2AMTNlWS
JJwQ5X2RpieyrzIGPoIjDI24lK7DHW33owR6eomjVwen3n1MOtM2mXirHG9khZSz
wKR7RKbYTaezqtRtvpmHAz3Ra3ERGOfDtTidNFLZROXO/6hLRYphzKQk1pMYnOCn
GITi35BOP0XnsJ/9/lbpAgmHf+cijckc7HIUazKtyznWmsB1RwTSOCA6MEI1nfj6
9bf6V874FpsF7lrup2ry4gW6R9ZZZRycL7zZ4ilYhREn1mgzFBq1MiApv61KKvpX
NppLzpOrMTS7sebUVqyLs5mGTDNbnwl1S1JXHTBe8JZV0tQllnybmahDuYo/H3WX
aF6T0TNg4GxynUJogDAU833tLgv43W+b1iuyXbA8XvGMGcKOSrOJadaAMZFiuwY+
x3kZoajRz/PVEX8kaRDP0xZML2B7Z/bdwJFuuTu4osOse/7Z2bOpl99NMXd0608J
Ttscq/0sCa12O18QoaityugX6VM6u9k3SEw6RGaVKUeWNCm/2zvE0rm2AgI6enKp
jm/a2V900t/KR8Dc5Lr6MZiixPLds+Fcw5Dcb5oNTC5EvMS8qVn2ePxQKXEFIX6Q
h8K+WN0kwIrMKE1u+piM5XbZFAf8cRIIZgKPHM3GBiCklkpE0l81QABlFND7kzNH
pfvbtj6ushJR0C3cSky47ClHzrXPWJ1HRM9EviscrpXMfC0AlVH38iegi6FSVBXh
NXDHuAWuJ1wYoGpZdyvxR6306cD0f8e68kmVEi+vRwWSGXaqPe4AUy0lUtfa+cj7
ygl/91Ftf+Sg4YNtyvBt8aZ2+n4pwDsFQSE53icsY71G/bUvtZ+SiditVsdTfxX3
bWgGHnMd6JKgMR36q27IajJ0AEvF2o8jnonuptmDDqsuapcrvPv+rbgjBVixeN+r
HXFLUllg0H+rAUPU4nMHDGIeodlT19X9LiXT+exQS03o4CSB3Vf2/9f34tTYiE9B
drxKo9x5yGoOfJ6wEESdEyZ0ULeajcaijv+gQGb9AGmh9EJ6hhC93puG5jTvfTE3
ePPgXxhi7GJtbDppqs5X3VrIR78vpD/+QuE17qLBduTFlUe/KNk/sw5le8RKoMvr
XlQls40Q6Hiwg9jS2tA0gf9DxrID+xxD4jwRFSrSMF/Ve23yl/pT/tiGfDbQHcFd
JwDtRt8oXf0BMY3QK7AjLz2kyw3v9A3MWkj5f18PAvfMCWXYXdDUCdQalco+vaRs
adukWPryrrl1p8DP1wOIbrWX1is7W1Z7IWzNhxjJioXF1KY2/p6cKhtzzvuyMZsp
r4b4+owV4ggULIBBfVilPqEnyf11rbrLiNZ8VJhgfvBAK4wrxFAZs4apd5eisK+E
xSZsEVH03jhcMrxPqgFe7OkGqUb4Sb/wKG/aBcblvVDlBBJs49GkFaMwjk/WbzHt
6PffG/VvuFOq8yCa77BxsCN6ZsDvBKnrqgznUuquwhYQdm1i9gQcbw08zq6LlG82
ssBV4R8ayU2brZlNgcapaINqFzypQPdc3BBTOwFPr6c9IDl/HrBAiWUxYiXupFYI
fRImtKDCn8CEVqw7q5mCJtBF7TRsa4cPy65cCr++oQDbQuV+sVYzMtE0D7vZXp/Y
qxvPosdkeBcFNahP9YL/xbvud8E0PTPDPA7MVp4YToZ/UG7aXJEgSAKYmkfN4KOR
wVrUbbOaL+U1gkX1t8EZNN8X3PJ5ZVA3I+uIYkVlik2nEhE+pgTt+m9ULhbuwrqp
+H/R+jeR6k2HvqcEI74cBDgjlx/KjN4ncus6mFAx3BaT/9w1uc7kG8gV2DD8VX/7
mcJAPvezy7dhy/jI5f8DqNy/d29i6PZTidL3kdMpx3vNmb5Mi0eN0y3oTc5CJAee
3XYFQGbOCJczfxqND0SVwAoIX3u12wByR1nj3CU9tBGKl5C7ZZm6Wx6oK4gYs8KD
J7fCZ7U+VFhIz3ra4s2d2Hx3rkHjPz6Qg0Ox4Wc+HFicVPLql6U+/3nIkYk6ulZ0
sgvViRLvbtbcvEgaVBQGWJuizBJZYznxmdrRGoGzIGOqXHhJq02TGa5zAhPRQFWN
lV1UuZBhfWOiUlFzwlqhZymNdPH1pO2jK5a9wOH2Ju6FbEnY/aDqMn9Sag+LS7Za
175udBhq/2aoan41C8dFtg36lU+msBI4Fh/2vmIi3+JWZsQqqgDRktZR9K9G3GEC
5P+oJfUCl4Zr1c4X1/V9AydYK6sTfX8cz2meJslCZQtFFJfKupzfiHcrqMCnE4BX
JoEk7iskQ0uZICTVOhsfjuJbr2TevumRCEqBhOCiZlZzR1zA3LBLNihsGaPyTT21
R48EbDXIb/j4VYkImgnjisDlN0kDuL7mO637aVI8ao8tm1q+/QjuayGUKL12XKHt
kUwi7lhb4WiFeV1GZqxRxpRBA1OYQuKfbHvmYSzmxtFfih1Rb6HV5FBkXOAt930K
dplm3EdQ8vPRayoL5kqrgKcV+WCrZD6ecc2mE8TmrFZd04dj/N8IG54sLVbrbDf0
Cen1TXUqKli+2alpqf+qF0eMOvvvOrP6IZwEXFExjR/E8Yi7bamjn1slKZFCFNEg
Hb19938qXh2Fw3G/kXOj6GhdzIdSSoNu98AB2TSkKNwORTCdwjO1mDOFICCVihMB
+wmbQds0YbRzrdbslrJSGVUU5H0zaJkRBJ7DXegI9bl0gk+puiB+yVDxPnMGg7VO
PleKxn5MauTXkItC/YFtOprfgc3M+hLemzNfbRbalja1Z28iYOm3+hnJcbhsmwz8
Y7dDhy1Dwz3v25MSzrcfNOcZjtNWqWZkFnppRLwROfnbynigKSWTwnprjqqUvGk+
YEcr+WIqHQORL37cCrxs3TW3Ty/w0q4a2PprYczedObmhHBbTlxVxWUEcJjLs1en
hwTutL1BQhkrGg5eAVA5jWx5RzbC89xM0N6iXT6mvDuT+a3BUhft0Xh1F2SjAoQt
XSUI6mps3NqWbhNwM5Xnpd1VuiprcQHwwNC1b/12rzbf9LFAePTopZ968UUr0G9g
g88Wk+Z+cUnNZVW3lKu0jY43pOcgMJQq2hA+jm0biLJ2odPjy3rWqzNgzopFbL+h
vy1utRlTuSMH3PQoc1xTT4HfMUU5RpUQHXlfxh2hQLy7V+x9WSZmYYCZVnA8jNWR
d5PZdm6hSQi1QRFJzbEn8CZaAuNxLUNfaxx0G/LCxgsO0/6x/dVDiwxIchpMVIRy
v0CVL7SXWS7YA982n1OLg4cz/eWPvAhJLsuK3hF093HPAxIifO3vgnGw33FtgMkM
TCzoMdf6dUH3SydOF83kwX8KHJ9n721cu7GdBrc+vpooiUFl3K7+EnUNnlwdnHR7
dR5pgWfPMXMfnLOXnYmidS/+jJEilJEZ9+c7NHJwl9PB4GUXkxD5nvhMZ+tmVB/N
ZUS+hVYP66R9L0Z/8EEUGQitSphtYSDaGsxzxf1+Cqbp2dXf+q03yzn92IZy4beZ
u5AcDfMhWS/Ewe5DToLMhHKa/Hzqd0OKjYpOz/b+M5OutJf6lIw/9c/tJxcvJWlU
nY/ddNV3leVhmAk2QMBz0Ns578bWxfj/IeMDz8JwDrxNEVAsLa4b88Rqgub945vN
DAiUpWgGGdU9giCzUflYUpKBWTdaoQlYju8lNpF6ODVOu3vYEFWF7QA4PSgUOT3y
8sU0RChhc7EyIGwGxJlCpK9wSi+zaeR4l0oqqunRQdi+ecVIzCgaPcMMOiiPHJCg
6fwJw57ItH7XHOwxXZ4aNWmg/eBMl2Fpt2+SuChxdkeCQox58bkw8NM49IxOci6c
NUnu00gxmAGQCR/iMr/4xtQHkci8ZWRi2tKrxj6Lhd4XTbc5voo8cH5gq8QrJbOY
sQIJemPBJBFl/+/XCJ+3gZFir7ss/VRQJVzh0trpBkS2zNSVuGlwHzGM43D2GO+X
WF3+EOi5AJeYls6frws+ZpLr6mrx4lFkduZHbClO9kEj6H3guao1PqVjp7oInuGS
E0dyFb6vCJTMcCeKn/ED3q1lCTNKqX1xdS9huk5u3DoC8Z2M2AaMP+tJ6v13V4ro
16CdN6oDnTZA7YrKqKZ2miMigWQPj0+4BZGfKuh3aZqPdfVAIsF8pRizqf3ZsReL
HtUi0HNOfRX3m43rPgKkzTYBElrfa1ugqHrNtUmzUqQ/JXCoigRbWIqlKUbpnio9
ga89gDZFSPxPLdgyNLS5V6TgmbSgezNOvmcIM+ApPDELEQXhJxUciLRor/0GFeYu
bnT9VA+m41qq3BnJ1v9moqNP0hBe/kWlJ7S5de5GS7IFqpbzXntcpxouWzgRhOO7
37gVgWmkSZw25g3f3Uz6KqwyyRjY4U60+DcS7LNRixZGjGywjnWhi0zYJG398V35
6BA8cxw1UM85hC/Oib8b8bn5SltX2VXIoESRrs/26840TIrDKtXoz0BJWjV3fT66
RDf3UIwl6d1m8Enkh4SofYPx/7DgjLeawbuPYfdQ3zZoPKxCglU5dDwYHalKz1vG
8jD7DYvxcQ/ZRk/n22agMEpFQo47jeCET75TT3702ZJdu+2iiq3BYtw6yQ3Cj+cp
hBl4/ph6ioaH8Son5IHtHMO9S2xRtLns3h1RUFIvdILU0sSbEvR+K58qf92atPh8
Z8h0kQc1QEhQld+0PLApFQI7ZhLtwZaJKs4f6JeO4Z6ilWOH97xOctFLcjHqvmYA
pZ2F0M9i73r0l5QC2ZxT9whGRghHeOvvLYx/q5WM0XnMpR1yuAoZKlngGg0BofZM
vVXQrzhqJShtfuJsjb0oUjj/KXeiR+h7Y5vMmkcwCG2wNH5Ro1h9UfkNXqzAL66U
QWyEOIBG+M5KNKJ7euxqfK7Xzi2YLHmyHotoKJ9szHiwnZvz3lasmlHqFyOWFqT8
0vPv6pT3JzFRpDNYmL0W4yYej4YfC05e/sjeBN4gUnUJMTjk6nzIy+pEDKTH6cBK
GERbfU4hASdJa/GokdmDnihnxOgrMQ4wpAEPO62B5hHfVpf0OE1u2ITqeRDghWvW
Ook6lQop7TY+EqOrPkwLAGWl6O0PLsWILvvUzA4ygM4uhTY28tHA5i3b0EDD+XoA
Hc7ITbCExTGnhPjZaJkequd/qojk80A29vI85Pvvt5ZfxRLZZI9+9H3EZAHMPUJx
qD701eZIMWG8Sh4uTRzg2duOm/G30Cvoz96WFN7cvJ66f2N5JunNpKyCvqcSwZHa
Ny4wvTlGVQWFbQ14J/E/JQF5K4hBX97nV15UaUUH27KITo7noaPsK6xPlnX+rbSk
0MiSMi+Wgb43VdbHC0HLYfAKA+SeL3NKURWinQkPXIYgltElLI4yUVKdgY9z4MEy
Ds7oFA1oF6KdUgJypIqEPCshQwea88Fa9yD6dZr505vGvAiKjZQ0tG4OOXEBiHZg
PTTzcNrpo6n59hzb7NxoxA/WnAAErcofOpCYl/v2VSJPYbe1MciDFfT/ZkhNW3jl
/JVn6Gsc0tNV2Z7Uh0AHLyZF/EBSP//cjjauLQiZ3Ae01/urPX1Ydz/GEKhnJQJG
1BXr8ALVv7sLtS1U1tanxcdxIE5l7tJ60MUsRD7wkwaGGqBE1MLrJ1gk3eFxeRrU
MXG5G/xZl8PHiqS1yEF2wxpUW08w81zIC3KqnlMKRnGitUjUAUm1WKpxnPexvgqL
NhHTZtAIEsRME5mRVhsIRTvNPX+7hbkwMN0kJnoSctMfM4k5ivvNH1kVLQLCvFgv
EDY349xXF/IrS4ARozYqvcwiP+7xZJ8N5dYXyk3T4C/CYerQvecHHcqMjUVnQYYR
4KBdv10giGOVmoUpft+OjFFL+NoRuJEPGZiKGMPDleisaNY0e6++ApbWIBfp0qOW
J6XGRTFl6PQWkH5EV3aRu9kq5tQv8YYaM/yh4sSWAuy7GxVaiPkFIUxlwrbf42mp
DCgkHnMHORxmt5d/RrtHoJjTWhd4PI2x4+hV5pbjug+uxgzQjKxFdGhTKfSEtObj
bCsNht7sXi5yUzAWeaaW5jV0FDDNl4yIvNejqiHPUg1AcRbKc2tflI1xl9fhuHok
VumGw9fHcQut1cSEawZckXPqBmHcO5s8tEAj4PmHzN+n7VLXKLd/eaflb7sX3zjH
CSPJFjtrmqKOU3WmwQcodEtXSQOa3Zngc+CV8OlqAN+79S2fPyvQVAGLDApDdGLq
GAtV74wh5+qTq/SwI+va899GTrFgzlEc+bC3GZHxAfEHzmCTZHv1UtpsnQeQUgXR
YHqq1l/DW+zd53k5Pf+E4Iex9Tkt1w+qdbIx0jwRha3gJuJao1uSJ/KPPODX+2c1
oKXp+OYPvuP7wp+A4rfNKA4yRQLB8h1P4Ua29eODXXVETP/hCE7jIl+ZtSknVNSS
aqtl4z2fmZH7vyeXUmlywFbFaWTj140A8qvL+R84/8wWAasaLK8Y39Fa9nJ9XJr7
oYOUKmkfz9Lku38KOb62K+8sdr2U4Tm/5HMJRS1pFvWLYvMf9zfiwt7ykxWdxjgi
QFliyc9lC2DaVjqcQSxfMKfAoVLNhgdIUYe2zxcYJKupzXz0ZmcGbi+Z8wXVTAC5
54SYv+cbyrONfSZFCFdPNkFx8Q7J/awi2wDJCySiCCY0ie5Xyol7Kx4JHWtQEFQm
zfmE7Smy0cFBVI8qPbNY2IfC5rOvrcm39ov0WE1X5cQkytZTuwLqS1r6Vif98O4J
oGZCLKBhy8bmP6BBfIbjsLT/6TkCCH6r4aJkBm7UEbqxIEWY1xtNkq8KP37djHwk
zdWfJHOGbdGqdmwbOhyBilucDNhE3hdOGC6X2oBabDqeyc3tEjMiMo2AJn0sWcHv
ks303RogiLgbABw90Yo/gC2qszqJCNReUZVvaOnjngqNDvGk9wubXiaCwOXFFBFK
UaB7Ftd3pfKZE6JhFs/fnD+tDDCHz6qjNaZQWOKlrSzGkUW3bgdy2U5AQ57QhbgE
kRBIa/l5WgMXkAQuoFSmnI6UrLyedN2oNauHyCgWko+/cgat7iu0fbiQVu7+Ah95
gtz+f9CrPf6tdU0F2zdbJG8rLnS2ohVdYsuQVpCuona5JBNo/OuAGtsv+xy32JyS
Sc2VdCFWFnjPS2r2UzSrXCRl5FlUByXqYQzKGJnfsiaSYoy4d2SXC5qc99ZnmWIB
oWtK/SolzZC7xE0iK83BbyVV0A6mn0cRPuAqOd9NCch4ojz+CI/Ka6CmyHusijIQ
nrLTWYSwmFiUjvyq9avtDWTYXxnRLGNsWlCvTTEfKNZ/p9r2uatZ68u7rLh9DtLy
iu1KVshP+hNExGsLMFG01kLVlOISJ6BbYTj9akQ74gfacycG6KJLEieZghtGUX3T
mKgTt0tag+QRW+IpyDMnwr8xRHUDGCypZSidgiqzgu2gtA1Dwot3nSJ9f3siPfdt
SUVFbdZUQe8nNPyWcia6VdYOCsLAWa+6endaB98/xyti1z+3by0CFjPQBel5y83/
9Ktdmo274BPqQmPoEVWqtsK31LSG+5oXMVuXI5A/9D100sqsBMIcaZi+LTa9lRmN
B/9fJqbuklzbvJSE1afEa1G0tmGQDPldP3IlxhY7+H2Q8+s8uxvsdNQDJYJgWhYC
l3VBeTb6U1mf6JP3w4FwDXLDtX86luBCo4UTF5i8QqYTwFk8TR7aWQG3xj2x9CIJ
u6KoBh8KNEi97IiyRKrqfBDtOdgXXeRKRdsoUMRnHU2EhZlBVxDeF8P556jx6JLT
TTAvgJwX8iN2a4Z9tZ+15UztfpPYV/0ay7q8NNg7NArIKAIuFWMJk4yxlTj21rwf
g6YTNq5bTS7B1AcQwxCY6L8WymGsgfYwFPNrljYBi0En/AtxPrZ3Lqn/cC/8Qpgi
AdpjCZgaX/EOpUqHeBK2aKx7t5UXDgYMxm8QwyNA7vu7nPqsGjpWl1S34vU2Tvk7
qiFLMy95n7xJKyb0JJsw8PZ1gwlDpc0WOsTzT+KUY/+Fb28u5dL+5lIFzM14Opdl
1nRbki7cSM07Wl1fcM1L9r/ep/f5hP3Pp7Ml2evfTiJ2vmvwBh0o76OByTSVzkhV
h801PjcRn/tcY0HcEm3SXQu9fO4hvdMx5emv8yytb3Wwz70myZask5PXuZ9dslbt
ABQPoNh65Mam/wMXZfjACpDk41/eXvAC8L7db2ctfhIz6Nj4QUWrjdal4QZfMnZZ
GrulifByNeHmJLwPoi/kdt84X65Hjt7bTG08SUwX6+sRHB+4WpLJcnrXgdG/dQPI
Pjk9DiCwGxDOpG2BrWNF7eqE+Xpdninf/nGZMW22lKXxxT/Op+6hefo/M5QQiKx6
KmmsdPiHSvWNy7Qwzi6O0SdxPLxh2y/TJBStr1i0y1x5D2/uIVP5LXJt9bGPw+wx
9FF9P1ccrfERhYKk53lnmrI9tfe8AhhPZZhVTfOHqLlq83w6bK96EXN9UgNWkf7T
4Ozj1c4kZjiKQie6z4/RwIlmetYK3Rlf1VKWFqrUTwTuumQl+J+vYn32VFRqXvQ/
nI6WpNT1kS5FI13kpniEknVgO/00Gxa5GaJxieAhR10i7Qg03oWND72qZfFLU7j+
uud9ErVN5oR4StDHgwM+ZV+du0isjLrJ5TSPRXfUmgYLert+Ol9pkyi6lMKPHKcl
jgORejt/LqKBGwNtMGcCrGxSi5sv9gRJ5ft2OAyg/hGhPTlldES/zfslMY7/1L29
0/NQFACjIALzIUdtkQ/yFdwEU2ca5h60TLcXxqI35JP5ZACZMK7eqmAegRXM6k2V
e+QJRw6W5DKvucucJZa8mozYSnq0ElnFYKZ/aKGd+Ar3HJxJFzknq14O2/LrbHj6
ZbapgnUC/h3EISL718Ct0PkXa9UO5sayML4TZ2lD2vOoAtP3QTyOgeXLNWi6lZlb
qclsB7Hcd1F56Xfacb2siFhZ9pez3JD/nHKOHZvsxhCnHd/BlQwTDs3bBIHHw9dx
vLHi84zKVyafpUbvp1gDTga768cI+7fyR0plii2KdO4NlejI15MkCffByD/T0BmS
/Oh+edaxjT43tXoAm6QQ/T35ViTjvQHEE/bwAJ24AxqTcYt0dRpVrjQuJzVedQJW
/dw651amMnsDfuz5l8FjUbCpYT9sdHnx2bPCl0s1pyIuI2WtC4fmHMXsPU5DhCF3
M7kK801Z8ck1vxM/Uds43Sk12P8WXZyKWnV89aicIB7D900Nk0RItjPzxZo8afw7
IM5dMLClGu1BLy8kOgChdL26+Z/WmhkQvr871Ste0/Skwd7RfhkgpL48qsWZ7kpF
Qzz864pZD1UjUQC4XCBcw0x8zZRijtJSMbMGE/hMpstAJcT7Ayd7eEfuttTm+I7C
9rBRsCI2bDQagvXSpUmC90wY2M+VQgt4Xd8xsyLr+qCnC/d6vm/AipbWaxWnNc+p
hMTOxYFeUMfxz7rAbFkoEB9RnxZGKd/de/6t9epBlGYmv7mauSgdoy+ch22JnmW+
xp7tPkG/tB4BIIM+umktrDfA1zQ0a1mT4ei503lUf6clh3LNDXYzMLN7dNMzmVxM
+SRwDSNKUgHZO5cDsdBvRvGsO0Oiwkj0YqXnYxjVm4Cy52bRetlEqM8G9nsmlZqD
WKnR7c4wFI7C7DHLtdB5NjLoXMCWXoJbeJeJTp8nYL3LphyShaRgwfmL9+ZMFDbA
0GII2yyr9hIgZvcneuZT/j6mHaNOTGKugmGqkrB59Xq5psOQpkfry3cYYeYbhEzb
i4Z6sZqC69iAReGiGJ/MF0yq4zhN1IoirWt1vPAZVxVyLoztQtunoLjK8EwUxJSQ
fz38z06kqPFyxxkhQFdCWmbCVUk7SSjjU6+XZza1XOeCRfqhuJ2quzYyj5fDUqXA
gBgcH2sAUnc0RnNxAsmGf9lR0GmKT1IeTDGFXEFQ7B3uklH/NLiIzfbYwlJpVimk
ItGy1rnsZPVnXLQDGg57xOC4FaUyJ+oHLKdtCSx3dxmwrJ6oqVRanBcoB/BQ25tQ
FBCEhYhVnnzOIS6w+s26y0tMOHncPMQt/aiGpgdQfE92ma6L666OxXuDDphA1kGa
toCbXrkCH7G9bj/PwhJPfHklHsWw5NfUx7id3/uXsNtlsHynhtJ8/0ZHWVWGKSj8
YejAHrP1tfyL8b4DngrBTblBBbG5MaEJ0wA7cJ3h9eSL3bi2msUvOSxAx+ZyQUbJ
8FxgSjp25BvNWpA9//H1jk3uctd/VxQ+0PCpme6aWqpzaOaiMnmN9qF50Nv+bvaX
jfPjvEz7bnnLYlPhmNRBApb5yb9GGfuVpeVXgCdpgo20naTmlTrcEmBM7k4HjSau
ne+O2SDlofKktmMOvhFt7ZyENbs43HvuhMhv5zEFewoCMzq2SIeo2re2NHGqVw4P
Cr3yHTU7yo6cFqgvDOp5etoyZws1lrslaA+4X3cehAyJJM3tAuvvB/t+eXjqXR/T
38lGeMalXx3rznzG2rSDpM8JUCFMlwOxgaGl+lrZgWHoGf69DIKywi2ajqPfMSsu
JFXgcto0bffag9L+u88+Hg00c6o8bVkKLW7q/000xk8oLR/om7zRjyEFKbS6Jc8C
cSabPAaT+zYEzLgTWQExBZjuDH7k+3rF9gW5rAPWz+gpe8G4mcoa6Ep5Bu+5irHG
vos5XgjWT/AoK+mOWBcval4W+8dmBKkX6oXUnDwo+YuJJyl0TPUFX7S3M5ZTMrBf
3Zsmjyxp3crqm4rwM9XlmYgsB00/AiwWpjcKdY3YIZb2ZkGxIcuZv0SVJqomLovE
d7HN1uMy//FvECoXKCES2axYYEmkShag5gJGQ+ocLe5bR9Pt4bgoy0/lvghgxCqK
J5EKCTcJjtsX7nC/V69IGDfGeWHFsJ3dJeGzZWONg47iwm2foLGKZIe54g67Wabo
MnkJ4GTmzj72RskbGkvmNYmZqeTdwpngf2+Jer2/zwddIYVd5p8rYAhlULeIxm27
ZDMIMUZ/ZYFK2oMoLTpkqjc3OY12rb9bEBVXRIs+QJgFslSXamKHDyYjhL06eiNf
OBPx4OtORQFdaiYuhHU4Lu0qou73z7jW74u5AgZpcols7cT6a9MMKLGOQqHUKhvl
TbwJO5JXWPRnPNyWCljQW2AJTezBogl1cgzTK58sFlN4jfs0F1TTVVYmreEctsZL
5TsGZNsbiO5Ff7rip0JKE7R0onmOf47rnvQVqQmO0mEBVPhjV5Oi2mTA+BRuBfHe
8d0c2Kf3LxPT5UIbLXJq8sey2LJUeaGVVyFZ9GOUSLQ5tVMqvOKGdHcRYVy9B7kh
qimcNPqDVlDyIfbov+qhrm5f95B4qTPMJWXf76cI8apKRgQrC3G2JnnFKMEY+Iez
uGXdDqdHAnLR3eY9qxrg9u32zhk17hstDmH+HgkjZEo7jWnVKkv1QEgqObTXuaAI
7tNKuF4+AdynnYOpF77+prQLIIWBxvKrbimHFXCFUSE/4qppGa1lwPbrDTcCZEOU
XhoWXY4stJoEJuCqnNovxDL+sZXg7/XwQyVmC6mBMXYkkjnwbqXXdZfXCbkla7Vb
Vlj8F1WH6LYW/SaRvcAvI99nJax3Fm3TvEK4qePCYE5T49+0JR4uFq/dCfPZetrJ
IC2wvpQ0zGYWKO9cbeabbnMWXyBGFqLXNnTJ675GicvbidKMcUVgSnZKcfWxXcjJ
CVbQajWlcUTnpErjbYshZVz83DU0XE1aSvXG9SzljdUpd+12mjNk40ZdpHqF4eB0
oImOnFTWYg17CpIKiTHwCQBlK+eC/Fzcj+wvzyjIclU5QPmpddnefiyWeJZYbY5P
fPJQgbnTxeMt0mIyAD9HBJM2xrp9V7DoRICd6ANtG1R+tHhr5abTSgblGC6S05zr
jxynxSK+PU5uoB43gnCAe4kZRwRZNvnVFm54xheCCEGWyRjzNLiLBKxQ9hsSFlhc
2knN4Z4+7p68T4ZLMzvkEAyM+W0Ump7TA51CCWfNvXluOrVD0j/E9zBqgaFEZscV
DBWtJrorlV9baQumhGQLIWtqUJExBZ0bY0uLVc3QPEEnVLgiD7unB9J8oLYD7X6Y
oOlTLvkHxch/fJw/SpjK7wkAtw7XqC2dhJ9he5wUmBM38I/Aik36hCWBI/iVrJ7f
M8JQarPD6FBSnHW/iaxa4fP9VdW89ItdGiEJ8LH9r266VLk1BPqwIndYUpEaPqkB
kEDZxmMCes1yKdKDU9J/9SscvV7uvi8GfN9bRaIy47vaJoLV0ienckR9MFO6aegv
t7diSygRzJykPDL5Evxrw3upq6CgPrd7YegxRACiDCswPQSKTnspoz02ggq1/jJ5
/KlK2O5S3CVxPFv18gAF2kwEqsiDr5eOgUpMpKeXK1ejAOuB1CTk9L1284t6uy67
5NYCPRM2UcZGNQAeKR9+ZSgQJEqJxJxCj3f0UtjTYXQTrnL7GSVZF906KFq0QZyh
oCg5uqjDQiTm5ZWteb1fN812/KnStQ43EB+iVe+K/G2SMY7/GV3nYaO2cgyWCK1x
SjuSgkPTaKffynbc+NBrndNv2x0HGdLI4RWtjE87KY1eZCH81/0LkpftxNv2WijF
A0YtRH7DHbphw7YVDZ1+/bGYMso0pTUzHA9FcYFbgUqRXdN4TtuTiJ6MOPHGkbr/
GmjG97dO5cusY642H6yM9a8F5rqE/702o1KdCNTGdaHkvWjVvrAC128/cpodvBoT
P/FJSCq3ZUi0iwOsnSgGx8vqqRWpVTB4Qn5uZu6jD+eg2Haq30PqZCsB8vvm5GC1
fFGyO4SewFUvrBakcGVDXLeQZgmhv13wzj0ooOst69tiWUp4OYIKHXvJs3I9nf4u
RKCcu4OqWGzXii8yhAzKgv77DvjynZWfZJ9nOsOYFZHC666ueoCI4Au4nO31EbqG
Iuq7QVzHYFaKoEQEXFs9M9C/0tZbRcu0j0gawIqEyweI925aQf7P8Po8eFsJNFyK
OochsnWKrwXSkYKigwUkoIs07aB99bP9oPQXH666J6RtnNx8X6w2UuMpGWnk+BZZ
JSB+886U2BvvKfbq+8IksS0n0xRcPIiIRrVjlfEyXrO4qQvaWJWFzNeD2nLrdW1F
4HzAwi3oWNNAn26KS5t7ZPfzNyAoOQ55BnDRyL+gKlaXnWCvMJ/IaVV8wY2sqIAd
/jB8MlUrHB/CSt+81Su6wfhsv8ERFVfz32Sji2qtD7XTcUzgOcdszJezjate/4pw
vb0jPTUifzxlvcZOjuEA0eWyheWuvXNQCpFsaFDa6ce9/zptLjvNg3FBW6UkKeiV
jhaoVporCc/7hd3kMJuK8r+TAl/LaAC81zerUBdtFh+nman808ofcU7MDnoJRGYy
N56h8xOkE1fChD3XlfvK8TaVVkuI6nQljnnKm9IwOWkmnXxF1rq1kJ983I+Dpf+/
CWF1eBIg2UkEBlPPTzF/lyy3kVZsTFvcNQzCvvVB1C5C5uQhmtQrzR2yAUQB3Y8I
YuxC8imYYPUtAYnjjiDezn863YorOmx/EDohDkstuXmQO2y3o7eKJ0BBnStW4/dX
KRK/Xx4AJFslJokib2y2MNt0GuRW5WMmSZpKEPzIdXL/faW1uctB4rGQWdDID3h5
u1lnL/D0qvf13nxgRnTTbJlmwhxxo6ozHt7uVV6wOPR5awcFZf21Khv0nuUKXYBq
MmGYo0+SPpMXJq7zATQTPjO7PNNbdCtkfHLGocIvRleBk/f6CMzGYhDQn+HGf/JQ
etjA7Xe+UPyvziiU1b/yQ2tkO9Jvk1ydn0nPH1Ej1HiiCJ7+ld9BHc61eog6SCon
+Iy4mO8zh7EUGFl+GUljMtU0+yYGfVfagjVJJZLAB5b8OHXht//iZ4aKBHcq68C/
dQYnX8bH0X5LjeIzeWoZMe6SB0YyLt7zWrvA35I152H0wtv9XPf5IYbcmlR8SKwg
DgpRCvooHefjZYP5jfjYQfNtz1GNt9gvp22lMAzMTdorFalFZlt6zjESBDtC6cMy
MApe3/ThER1ybp9pJcfEzo73f/W6FrbMwWhNSBq88vO+D9t5OHWM/BC7dDXN+V81
TMEQ53mF72O1RIAt7PrKBVuQFD57TGuBGDPTaLDbbQN3TGWlD8xOARTYuCx1ootn
mz2MSMx33sPQHX31lvKBVDb/+lcRiD5qQoN8INF8w0J3Tp3Ua058whyLHN/qzwDZ
ON2BfZVbTnqTMcdBajiRmxGDXNxTb/MU7CUsDLCn1GPpPQ9QzMLaDitFHvYyGYAE
jM41PH2IaXkOfwdoAKuDDoV113+twc+SKDl7HtK1Ey94ESHEMLgu0hdAQJXX2knv
hJX0IJmoE02XUqU9SaWQWgU5Sueo2hDENF8u9TTbZ0hErDx0SwmhyYuJQvJ+XKqk
ZRJzxbed7Jb3C+RB4R9hGNJnXUd7UzeuvtaqGiiNeSdY4MAhXtcKATFZrRbUFMWk
Nu9WKSAEFYrdq9+aqRy/SkUAnlydB43rLHc4hZk2nz1wpTv1kx+HiE4M7VOD5NX0
qkZay/15GrDzK9T7KnhqOks/C5BGV6roIQJCtiyHvgORlUje/qoMEepYFhFFN5nt
fpzAeQabijNTAjwkwVymI+Tqs2b2t3Khqgz4tSbaf2sE8iEGbtfb8xLRmeNvnOl/
2Ke2JmVtIuRvIkWexBDIC+SY9BrvXlC7QBsXNPlQ+U68VGBsOjSgMgxKFWkyZLM+
XYIUsDmU2jRvj/+5JvpjNcpbJeUVSljOEjr4f7EW9qkHRLFypTDYpeDOXqOvgOAo
c8FwCiwoXkLtMSajJHwQCqrv3O4XKc7LtO+kiWkH3PQ+lcwXNc2DeUoWnSp05sb/
gzBTQK0nymCABQ676SLL1k/bMkvYDzGE6swox5jiyFxgfzBhIEsjcEM4G4UsDmud
vhx/w2UycjkqprEoHNTMxdeDhzt0+Gvae/anGDayiQ370U5711Y7jjH099nGZWkv
MyCzIrCcb5dGMtLwmrb5uaBSW/PcUFKV4Q5Znpmk3TxLEvelLCJJZ8KY6x5mxNN4
DBNKu4fKKS4hZWlkXR79TyQ2MTKJioGTNNaIQ1SNXLD4he5rTBS8QDPXripOlvzg
s1D6d8udMehsYJevUXMSkz4NAHYdhtADhPdltUiuASYMN66mfoRg9TfMan+TVHb7
+fWbop5FAm1MsZ4WOn1LWkpeU1gyGMYwnQ+AiiPX9RPyMYlXQLGhANZndKw+9IQC
fPb1EYv5GuWbjeiPaQIoSKc7RLVx2cgmlUBU5EVZBNL77sYFUtuRIqQww/vJSvll
PwSZd/jmLf08NulWpDtChs3lEocarqhgS2X8RVOr8/kF5Fu/e2N8Zdkouo+EphPh
qZO6zTJ+8Mw15avwRM4gYY9PccBp7PUJCelkW+6XSjwIHPP/UcELuglkyYZLSfR6
gPup5vUrj/VUyX04lYtTljg7WL7rXtK84WKtEqWeMD0yL17RShLx1fpS5kDT5RCz
LVoE21l81aRSM0Q3gnxkQmL19SKP9XqIBqunDhwtIw3aa7NcZpLddYo10F/9zr9T
Pk4O+ueQJOFzXl8aN0AIM1w7uGfRPU9wl/Nlze+jNvHq2BNms927hXiLcXA5wYtx
fo9x3TU+wIdgIRq50L1UT80LCDMSu7HA7PbpxPlfK0NeJ2I3ZEeikQSGWNsQVAr2
M7x2ThhknsAqi8gmAT7rTK6+OXYIIRCtNvoYdpyhagGKRBURSF/x48peQj85xUGx
zMIYcTtHBN/FttuqnbF5pa4JrK0XfrtUHp06DizCNgUCVAMDBYpcMUwE3mKoswmZ
8uZ3t3uS+ncfJPWpWoqSfOVkXV+iog/TsvegHzYwuA17C8GUCXCoJJguhD4NkCkW
gFOy5nX7L4kTWa8TToYbCszrIPk1XC+w6x/ptgcHsGCU+FOgwsjAGN8DljBELzl+
k0nTby7rCs39KtXgs6v7ZF4dJSBdz/HULcapDLHnE2N4uii7kVmmfa7hZXc7Gg6u
L42a+gB8yzi/9HtR7cP08V/YdMNsZN5rMdeiyDcTIfc6hNrb0KN6rFpLoNVixo+J
5olUIoAVuc+2TAq4gZGslETHA/GWLZCYWgwHN1+SjllhqUg9g4PvI6QeeBlv/YF0
Bedw+SfuVGXuqLTRGevsAXc7ZmhP0iI4KM6kSftcYBS9KfeG5IBrzIa85a7d3XML
8qUJkvQKn1bo4gt0TrMRR7dRCxDP2XobtR6w/RDop8JZVFsHGQ48/FhHfSJCG6to
AFG6TUQoFnvVfaeDTYaDKD4RxmaT0DL8hnrdIvMm3lvrBSsZel1B1fBNgeXeGTKK
eiA4cA5Y5ms3fU6+/xblKoTEi0EFeIqgK6/Vnu5Dfrp/Lp9dSNjJFrtn7E2taEZX
8ZlnrQHYMEoJWCOQ7+fZfJIj/PCO8MebIglWUglkcnLa7YvP3ID49ZRUTao6A4nb
J3/uox7lG9461w9gnsa4DDWcbh2CpzgXizbxHq/QjkFkn2CvUimEpBAvwFmi2nqp
0q40b3tQJydWNDAE6raMtfjKY3uEL1A5F8IBdYB1EcEP1d9+PosPR/nIfBQmq8PP
9Y742ScX10MVr2ikHAxk6VEIQx83VpsO6FWKCAticQlBNgGh0bgo2tgAOsUfjsv0
R9Irs5PbNqSTvXWbiWVJ5gkCFBmM25KKaU0ir7/BLW0bNg7Xj9OEH7I6SADRPSKx
qwdabDhv3/y8TzWmc6T41rMNZyX2fDcQFjUBfyuI3td6pvxqUHgj2cUHHCgmkwI3
E1qyjW8JRq4Lrfj3QqMKx80iMlujeKRlaWf13oEVNt36tm4w7ROkHPvC5sW7EdzL
DWEDmDlUmS+rfakmEPJpt7K002x3wZqvawNEIYvcIWtwKBwhh818x8hfwXAOTO5G
H3JrXf+3tJiMoY3fayrYZ3Znu7fAmVN5lkTtKweE3Epsvi1mbdoDQVcIPT2HcGwW
7nBu3g5X2jz6fkblfCM5fN3uLKeyjohuG0QNszKDSeI2H9M9a3Mbsu4HEUPDMCL8
q5nzeTI7JWXKOcW8iRdyRB6I0VXrcQRd43GK7YEgNNAeE2zd7Ve2wuODvvfc8UCE
WbarjVbMnbqEZ22F8+6QqOw5th9mOzKq6UkVFs3jWl9z1c4BYFfGxIHOtU8TjSgH
rkycZ7cxyfJSU5M++i8yeNvYepVTp13k1pF/FxzDizZwTWwMxbTHZ+DQVya/KT3u
pH37Y9XIB6qHyugup1SceS9lxPUjWYqYaFlJyH9MMBvHgeswPgvCYDYi5MmFprCu
ol+fUnQUWUlRd2FDRYGAPRyCQHfQbdLcbbO5Ea3411E1LWpj51mdlMN6S/+urjJb
7XbRFa7UQ77Mbay/pyWA8Gj4F5zzKgfpzawacEjQxi+zb9D3hDrUPIPUXk6vy9JX
UYCEmDZkarf2WF4Y4ga1W1CE728d95WbocovDi4tTuVU4PvCjLhzqJDvOYUjhTUR
W1APhGLxG8ZaqD3rlT49T3pHbg3eLsOL0hJjCnjfeHm4f1L0AKO+k6FXrJO0OY2g
ZSa9oDb5kNy0b5X+hjIGD01KtDVSV/C4ekZMHZMEZZlnxl05MU9yWqHMhcd25ZCY
jLcMqQLXLb9s3xL/VAUnnu48BahCZzCpHRMcruBQZ4lUlE+3U/D9+CAu8L6ggbfm
BZPnFANhwtRs+wqrzNzOv2iI3h/MWZ1Yyutnz6cME75wNWzvr1eZi/5UU4Dz8l/x
lx+Etup/hV9OMtb5KR8s1qMjQnk/ZZ6KmTmDgnY/ZAQ/Gxb7gUx5nw3MnArcwCls
xJsD4+3B2TlTN0h+4HiBc7A4GYYQ48IsNQgFB7/eKxvvlPhtVpXAJ2FSbrOVfe1Z
14eJ9QN0HWk5kjgMXpWm18zvKrJXuhj9Skt9qfbkrsT6dz+aA7WPoJUVsgNfwgcy
0rSt+icLyYL5NLIYGr919I1UfOd7eaLVGHweKrTKlcZ831/+Hc/2O4xQnn7rI2RJ
XyLU4nOY2P+/E31gmY1YqDjeQSpzBhue+cZuToql2UBN13gyvjSFMA+14JEUS5Wb
7ImRZf3m0LZE+lPgpjE35ciHZJvHCubEDDqArndf9EhsrIGG47XVRVw9Gv8CwbRS
NSrxylKqHs+3uiovWgL7YX8CW9qu7x12Re3C6oHiRF0ZOgSJTFXycTGv8aY7MXHL
UjEKPWHmE4oJoUqJK7kmO0KRhpNzI/q2SG8EMDdMELYBvyOWquUcojQXgMERhpWx
H3WSMzp+7HSXCBZIbUjYSyc2eA07tXx4Rh+Zhf1tYDTosAIwd4pHAkMtDuceXnTf
KB6NX9la8+ZEla+td+/E9MdFeIBn4b0+axW+pp79KCuMG9gVY04hr+gRWsnzydEC
PJzrHIlmrs5mVM+LX4zIMQInLAnw9gV4Gz3lJGZhMM4HT7rPWGwjK/oBrfBwwbMN
KKXm692rvY/xSgA5DxKzGme8uRTGJTTaa+e/ldoYluYMjPTaSINXtevJL4Yn/9x3
zgJ+u//4jcT3jaydaaT9eRVce/mq+QvH1ceabhE/2dfgzoUX2uV6nqbJokK59XKp
RmaVgDOudkQye7Cr0rLt3nmdi6QvHxdJAnXWJM7GQZzX6dQqJJAs1fFzfgai8z64
Aa/vNu3XT0cn1OMG23Wga277iiif0mjE2j/SdGE8MYnai5p99CYFGGSd0UVrVm/6
Xv1u74fali3MvCbOslkrUhY7KUBFkRNCbukUwdFRp/l96n95BiCce1rQ4sU/cZ4E
n9HUF4CvhSowUxuUsW03f32n9fFGgRx60vdqKlg0zb2WiWoH/S/2LczMQnk8/7v7
b4TPOC94ZJKtGa9xLebJOzl7cxsVAjtybmfHC/xfePlNRmg8WzHogdgwFlqOsVY9
PPk1N0LGnwauxjV4zE+8DOibwECVJLPElMkeL1RQugnEEbKZn7Hhjn/S+KJDVmk2
ZvRqAHUEgYlZoiP6sYUtHz/gl4fIsayxByeGgwM0GHJ5GXDXdq2R7sNTbl/x5gZn
p1dAz9IRUMAld51jrbZgDovS9iJPsbvJYtbJboDP3bJ61g71ePAP4wEhzjaMWw0A
nvXLmW/RdPlytZysyLRt0ZBMAPKxtHjd8f6NX3/cmobLU3pIg8b2uhEvuNvA2H2X
kuX3IyJcU7PnSMk1My58DSaMNpDCuMixy1o0mSCc4u9EOm2H6y8xYJs0i4kTNxRP
p7U5cgDp4jyN1dqeabvdP7V9d6lXVZZfQqH3SO6ANc2iUZXiR1rtiUfBakF2hhIV
stK0dsjiML6UcFZPpQBSQNI4KX3FaSRr7ihA30GbJkTJv59kjo8M9DtaOVBHnZoK
GgYXGTz881aLZOXAWk74mFH9rVq1wbxA1nRVzxr+vWzWaaLFFsGBDWllL90P/cxI
Uzk9geCDS5q7V6JlfsR1r1ZgHySZuJk1ngm4olAaIpP/LcgpgePV7eh+rvVg31JK
gPL20FrXtnU/dyk/XiNQyhWWaF4bkPIg6SPohEwcq/qGSS2ZbXbpBBQ3uanTuCsn
Y/7yYqShgKgL3FK7R2i7mq5p7qILKGTjS+q1Oh+VTnqyCVif7iq3+Xd/N6wxTRae
ub5whIIuPjNdGeehIJeZ2b4Gg+hWoErvkSwCI6gNBz0FL7ztqPgy+41T4nz1JtHO
wZK2qBjkpJu3qzqEB7L0kWIRQI3XhmrRDnty1GGgBMQlDw8WeWlpAKNDEqdvr0BK
8djGrKUG5rMKbfXciJh1KjVeF0MnMLMH7xqUd4n/bqYXe+2xi5NGW9v11IYmdcLw
KMco3oY2pCvXtTo8elOakIBMkth5rN1r5tbDIFKSdffVGnpQxx9z7sRyAJwSDhVn
d6qVXgcAiawDedqdhuyce53/kvNcS9Ra81ywUXynFviJMCQ2SQPnYOrEAqyx5VaF
VFbDn0elPdsOzHnSdaU5Ek9j0Z+J05hF5AefV8IX5QBWQPZBO6jWji5odhS5iPBo
MEmVXRn/EuCTW+hfPxACz+TjrVfuv3Xx1KRETnxW7EJkqRZk2pzAqhObqe5OAJ7r
sy8TqpHkzUF3r93/JGo3qi7z4nB4dV9ML8MpOkj5o5Qjrk8bbiIppJq07S+2CvjK
fijBVqqgQpZjXV1FU9SaJlUI/PaHcntYsaqDZ8R5VFY1eB+U3i6UlohpOPI2U+HL
LJGeScXGZaPAQO7WbqcZbt0DS9OiFCp0oAAIvabZVMU4S9yGS/Mm+YIqQpvtd2uG
J1C6FPHoQalo6eUH+vE29mYyMNTXizaG0P7iq0Pdsbp/Fxr7lWf6cENrlqgT6Yd+
hCq8cBvilhrpS+zaxgw8ku8qKyaQCB7CZ8BTKlwa1wUHICFN/Unj3bXL/f9aYbLO
xLsB3DPDCIdUe3rRdOSrBUuZS1FYJgkDez8JfhOX/l1JaGWVoxiKWTvIsD9QVN8E
FH9lrFVUthUXNDlttN9kKrBJxFHxFFKP0hN9QvUmJmRSLxf8sPT1mvkZvPbjoS1m
yZWJzqcTKcg6Q8wTnrxZd53uNBdoQnGby/q3uHidpjhcFV3S3osLdV4du7xJi9qS
z/kpWQXgSq4TfJYgQ6wuBTf+cqGviIngTD+UDCPft80mHbI3irbjcJISAv56ytpt
mTu9tz5ufRi/EvmzQ3RvVuqa75zDDjxqYlS4WaRe/0kwVPpddaIsaBTyxW2oxfPm
m6mGdPcjYXJnQr57zsEeSWkJVW81QBf4fGwoftA4jEHIINcmVAAYwHC9xPakaTGx
iLM+qQ7im/v24d1B7BxEAamhPdTtijWqfoPjdH2bMKt6wgi313aZARrB4dXsqdTt
N2/zekTEPRxqbj8pVk3rHRTqAif863+ca0FHdKPm3+DqWOw+Jaz63yHOUhhI5fzB
YGciAiiVXjUyzMQlqzgNRR7Y3KxBwEwYyZUtDL+n2cheXzWrcxCdmk2p1JEhYmQa
k/ErLNxuHdf7lOd2LO9/xYeW0LNGYt7CRQltyN09WyKRInNjCml5FGOxRsxPoplx
LiroH1cT4Q7IcNXmBRviwY25uWGqwVaJ0xzB72xuVhhtXG8j2gMi4mDcibGwYkAF
QX9hosuMT62/u6CQsA+NCiht2P8FTKRoETZa3lFvcWfPQCx1w5E+VHLkEi0l65Sh
PwMV8AG8XJkMTVJ12vjpCghPiU1nSpop9CW7Iop8mtc+s+HRutofjKcAIc8MjmjS
tQqUaPGWDXgUdBcUp8yCTIKmQydblxzo66dXxzvidY8vsiYPZdTetjQ0L9Jo5Vhl
ez34O9NK9uS1NAOJuEJyem3GelsRGwH5rrywC3xi1aaV6c4kYZ7uYkmu4yT6NWxF
4QisAl/KaSaTjKY0qRqSt1Bmp+pQoXnWB8AW4SD6CVpO+Aq+rSLkDE4H4kyCVPqX
51J3NEX1h0SwFGE27a3d0v9PAVuRZPX5BZYaiL6CmhqGmeuwWUZDIKvOcebomnVp
zygRI7aWB96TXeVepGotkuEAIoqh/MyfetVyJC+28suy/g2pF7a/W0FxTwRryEfY
6wFQkFSb8/RziDB0EuX/2om6YtmrwoOCQX1m69zGGasS3vFdreK6rXl4QPf+8mwn
PaldEAK1CcE5sxwG8UKFk/0KP4g5uJGDShnYFgk7R5JFiWKPQF7xD+JSBUirOZyW
kOTCSxL9u48ihvNIEAFxigsYnZSkhbgH+zS4vRNO1S6R+eMMYrXwF6VeJb6G6EcJ
rQCXrsm1VJZZk1zyj1WNLcWea0I2jrhrbJtdpRALsuHj5/kCKhA5A00QycAWOOLA
Oj4Cgbl6pTwVZN4bvQI4aMVKjcMz2VYWF0rUjQFODQ0jIUMgPExHlgCQmHwoPh6n
5S6bIrAkdzvhSwiKy003mTKhahtupfqPnhW9yOTCI7luyuq77S485npEiC08L7l7
27vEl2OfdG93xs/E2/tOhjFpSvz7AbMO8NBgb9Kt10w7B0BDH3R6k5wRgRtW+qTc
T4HgUHDMhmcL5Kcahsso+SCBBl4xyXw5li07dcct0D70Qc7J40Q7ysvUAkRRfy9R
Gz7ncxyCwYaKUWTssbGCwByiU9dQYMDVrsdbBbtmrdT54ueyHkFWjU3FtHqUkqLf
dD2LLr6i/rK2O0QzrcNMFlwHyvAN1xnuB+Og53/h/r556QcVps2YU4Fcwa0FOInN
/8Mp0EGaipc3ebVmfegPsKYeHhRVkYsLAAEEsgzvteCQnmWrLPhTmawDeihrxmxL
/R4Ktl21kkGlAWfqXvSggv+Ee/QmwhX+xJyED37DtZ46eTsr/mznnQMaJ8HeNRKM
XN/LQSrbuQQCE1QyajJ1slTFZ7Fno7gbpr2bkk3DazkIR+FmrqYGOySsJ2reQWnW
hCWuJE/IQN+VS56CzWKyi7x+jT/0DI6E2WATabjtCMHotnXM3HplstX0qMHT//1b
l+H/TyZrO5O0gQo2pjTjxL5McsxbhkULek8c3E+ish7ypWJOO5WiB4MQvNSYVrT9
hNdQVOXkMB9WTbxw8ImfKLKG3OJviIaQheBk8WAXXZmmX/uQEqEgvwyuia/5XB+n
AmO/agDNCevpCUF5d9uKi18xB7XRMYMI9QoH3eM6FAcptwJQqCyWL34XExbp+hhQ
t5aKRyG8ncQqDfj6M6hHNYuIDzFmD4lP98hkT89N1ojecK0BSq8gODBg2a4P+QCw
a2OorDhz1cs3/9QXCJmK+xWuGVW6qFE0QtTU8jkRlJLVDYGKcFydD4U4i8GjrR2P
olxeNmXSkbETGvsQ1pNJ5YXHgYSHe9fk3vURwV/v4LY6p+4ekBFJrJZmqK6eODXu
Am0rj8t0B4/3iAxvh7jDcpewvJtlimS6223KljpRJmWkDeZMCz9Achh07oTGq4gd
OHicKXOiiH1tgWEpoM7XmrA9wCQHVdTktXZTsOqHlKOlG6S4Kqaw38fcuEHdfqr5
nr67GrqDWwoRi+IqQPfdXi/m4RwE1e7wpEucP9aBBmNSj8F+asFjaRrVT12DyxjY
nIu9Fq5cmYFvfHPDXl/KWZnKzoDRvC74Eulac4fzM1ZNxW3TXZQ8Rp/DLkr3Rm/p
8tNwT86pvpX865ruEFyxeQOecMmPgU4XlWiEYRHiaEdc5nEn1wfRW1bHJpWdJzYW
mv04uCbsKLzG8AR5VaBPmQumPFMlvwVifLHonW8ARW36DiybrkRsbvajMULUFwLL
HEjBjVEBTY/gBPYMJDbbtngE+48WjQZ2QEYaavXl1oCf3TeHrDMjgicdD1/4ZBcQ
wJOZ/sZczxryQq7+Wdc9NElP0xI68YYxFhgvzycXv+xHQweB10bCbsIP5LXN9Edk
cfVcabfhsDVQgsmtVmV8pYukCIQqSfAMOyIALasHz2kbqiUCFZ+nx3LLy0hm6dDd
/BzMCn6UAXDNoW86HfFpArfYgX6POfs0gl9BqoRRWE2Vf/Fx8P4naV2sruW9sUIa
y9nPNvZwQGAwOp43J/MrL2cJ6M5UhCZqIg/6flm4XfQy3CNphf/2jayVmGHE/1kH
QW86bgh5gWaOy5g7IJm7CYzAwLtaeUJh9YsjZJ/ifOOC3o89i4v5j+ClnFmjW4mU
Iolna5wRXXJfps7ymyVB6uemKKse7/wmzOc+HLua7/cHjJoFH+by98JI25HSQQJr
qlPknDunE2hRP/bS+8+9hDa/cs6S/OVjeF9jWFvnuQCUQh8eb0atanA8fXMP77vz
1lDPX2k1V0PBCof70dBc7KPTDroKDf79vSebfoSqsu4YVjQYtrePQ0/p4sidbyWd
P4CEfqE7Tlh2bWc6JTRzudU/6SIqI9dzj9FpXevNmUgWF4K89DhCSBc0DKyAm0QL
mJFJMchNbp99qKH1dgk9xR/y7VsGPl6DpwqdnYDUFDlV/BMVQTtyHP1RQgFUC1Ge
RoxwUQOT2dPOmgxrl+8e+FmKnNxs7P5xDA+bEGt6hP5NYsCqyxSqUpfvsb2s3p1M
YIO4KgJf7eKNYPrxF65U6Fg1EXZgPfDIuzMhSLiZbjQtEpVRlIEBUUn2w2dQKRh5
1089UOlDXgH0DYPRsiQXH5gm2BCIDQ+Ddg6qL35Vw4lXljVYOwmy4/8uyNi82DRw
NENrhYK53h6dNms4BwtKuil3m+M/mII+pBdn8Rg+cVYVQ7HQncdZ2v8C4HJazmz2
by1YVY0PVa6rfUPSLtq85s++wNE3ByvWIBGshGca8fUNHR2ADcUuS2wUSDjaZJMX
ywryY80AZgDAHs7fI87es6QdeWiZnj6/Ah3w4lxYv708oLBa4SzgoxagkVOeWYPO
5x2CXHHLdxOTeZLOM/oMfp+Kz4jgswkuhwQWmNHefBi9e1oE8I7Qa0fch1Te99KS
dRH8heOg3rv96kb35zUAfXzm45z9Ue05hRPjFNIb1WVxT7gYrk+8XrPJrew0Ef+N
m9guQgUjVUeIG5ZsEIA1+qz+92K4dFMQ7yL6ve77Cv/Dg8El3z83S3gFpsObG9d+
BHfJNv6WgcWQKhM3IlEqfbY53caBCqtfGLdPfQNFhOQLS8MGLcZXs7SK0/iixVm9
DK6LgQsJF41kjTSdKIQLXdJHUNF6fTYi+gYJalrmVfWDm7HykpzF3N6MazjQo+lh
46ZtAgdvGowZUqCbg0Z5GckU8/3gTbfWnxVr/Dc1Sr3IKXhBYEJW4mQIe5yLrjIx
6chQmMqbfArVSqiCtGPO+HL/ZTQx688VtpdPlaWN6Gp1snpnFMBVHmtsgyt2/8FQ
gAZ9vwFnDeLYStgprrPf8giT35DxUMXuVtM5cN8TlMW5+/smJPE7t2xCSQk6TlIW
k3CNjo2FgnLA/Zy8PiycLAOky94qMCr4VKu5GYy2wAWzYqNtconReYTDveAqlvx1
thK3ijdc+tAwxQBqyyWr5zJtpA5KDiUoEq1aCQVmGUstu4wu4s6+cmCEUGM/x2kc
GbCetkvBSC/f/v1pKQ1QZJz4aJLGtC066Ejab2MUWxUMxNvekGj2UuQ6QXg230fl
6LkYFWny4jGPrrAxJ4UYenQaA6ZsyxeDt2zEs9XUt++Xc356vJka1pKMc7zcIpMm
VDpVfnQjgspYKMEqfyEWDiEScLeP7UzD5PiIbU5AmVvFIWyjIKHExq+Hag00ZgfX
WELMzfiJJF9klNlOrlt1kbk67+VEn27MYJFsUScVCJuAYSbFKKSgzSTh581An3mc
kJg9b4reVSytxEaLDiUdArEyGcPlLQwvdIcvbq5zXve19N/IWjxedbHVyGQiCgto
AgSHoC+zbDiRnROefLcNqdowfjTd7CnQnoEFWN1tczyM65u3CWTt1CZnUVFBkNEa
NAn4HwA2H9qUazU0xdN7uiF48rGZGPMNZ2NhA72GVgaI1md/9PwHYwAJe9yL3zrT
ZUbFBrA3GdSnHXufDCy3mVj3OwawFCne8wPLw0ZpJptT5nnwBcKPqWxC7wpu0qN0
gyluYQ3gr5+m3x25oR/AEJpXqRImoADXTX5+rVbXBo6nbOaWHTjdKH78Qnls9yMi
yWQi7RY4gMbxpioR7OgWkx3g30nKCj0IaI/sMEshmhaQKSZp3+z/nX92pv75O2zn
neORn18FBJnOn+mudEpKlHnY89aNJFENxvQuMLjUok9lHc3fPe8R/G+aJbrzo80R
vFvkDaSHrpvrgqMa+9nfAiJ8mHlfAfCIPeSDXDaZ0LllSb4ntbZJY/z3kXVKDNyi
JD28OI+iM2K0nIXF+WM1VuDfEKnC4/hTNhTHWwpMaOUTMujYQT0LIHs+/U5qjhuW
XVyFFMUTOPNftcf1iV0188w/ukFVHwFSeL4UXDAxsk/Fps2FL4xaScI8COrxGKxy
O0rIDZneMuAdHzRK6dfNmDRVNO0q+FL4UOFSBBO1SCuNFtEfbBeHk3tHZx6KyMhi
gBv02ED2S4Dv76sgT99Z1X8woJx8pF8YsFtLbmhWhyW0X8cXWW1KKV37u2CYHFNT
A6irv355jQSConyvS0LxXLYJp7dJ/X7E057E+1AubaRoGRbYKvretI2efYzH7DJU
HB+qR3Z1M+3ej0QaM3D9ON+ek5q8DUeg63Rqqh86UsE+o4Wc1jdin9Y46ncdVf7u
gGqVUj/kiSxsyGk2gDL+UIIbrV4szJ0NymbzDm1CYSKMxqgpPwnuk1hMhSWbXI9d
P/NIVlITzvK/zyGgM0M/h41Q6g8W50hJk7F55QcDucF+7YRRruu/X0KvX6+SKLF7
Z8+XLmkVBauf0W8FUgu0/X43nq2QFqc8ODFf4o1v6LNaqzYwxz3cXf5GS1WTzzhx
9ZQWjX0bB3fvMh2ecrnrXbeHAiXxpC0XEO+36gm9zSnI5EwoODvxm1BFP/PK4rer
I2O5h+SQK76f0XdKs3TJK6/AKU4AA6rU6V0JMeOlOyjqa3Ck7guxINbZ+N99+DF/
hdAZkFVJ0KUdLbBb6wSwURyjzKp84+F9Jo+Y3AtX3m3Vy7DaPwtnY2xzfFBRl/0N
wlGnjHu8VUOIZGKuS7ykhs7fEgDI3IhEWtrpqqhwKdUeEsi0MfIG9bKx8xH5j9ei
uCQ61sxBeL+nVKdWcg7Yer30zVXopkXX8t6dmXRaJ7cqPaKrHWmn8xZ6BwC6h/jv
vxM/+hB0K6jNyOft7QSLQRCKE9azodBTlcjOLJu6lM/vGY5FsVI5DlXAbzRplsou
mv5SZeU0j6/NHYdTgRKltyxHxmZJjf5PcGYfr/eHCSW/RQs+k50rbknzYvSw9hae
yRIeRzX8e5tlRgi64diZgnRrKrCAWE8O3Ilw0d1kSTywT8nlwlRqwcP3kyPnXGXZ
sw5p45GIRv+7bX/1ABFFrxiIYC3wjr1PNtPh1/shix6lcc8C2NX/quJKr6t+3fyJ
M/zMw6P+SvTnhPYWQ1QFUo0PA4EA6Wp00zYEyn3jl7BOLnCM/0x1ZWR1oDLdT6Dp
w7Lme7W611Ed/1n9ofI65l1I4/epN3opD2Afo1TpJxZPM6JumYQ8fCihI9GpvOs9
VliqQTQiknTnyLkMwQVuKXl2iz9GmjBcJiw264vdjgZXvR0iz3RtCun1CVQDw1zs
k39TAeA0hfHOXGGvxtOCeqRTyUV8t160Drdf87BMXuyaO6wrpQmMUH4KXAVfjElp
y90qatvo0AdnVxYekUTiNl6U+i+qcZNfB/VaWmkpucidfCZTf03aCh92534aDhWs
TPOfTxdsGXOjYe5MkNxTy4ANQEpuRU4q+8hYd8h68muAcB9cynbEdetNCMT+FNkz
fJumMXJl6K6T07fqJ/UtjfDtCcXXdB9Je6OPsjhLNH7mGGHqqYq1+K50vnVitoz+
mDEgrExvNRt2qnFg5wpkEH3dYrH6ML0Ct0udMy7IYidGxZgiJmA9vmGpZ76N6gOI
YN0/nmNsdGN8goDTk56dMUIoFZWhZkuRb4wrUwEmurJJGoNI/9UKNHnBH0SMl3jp
xO8fQsS00p1vFMdJ400m9dRCmFZ7ooAC5Ay6tLZnfQMnhHb04vmJmiAvaxSSU0PO
AboFo6FkDP4ziMDNYsinMmrRF+7zj6wiwNs9w9HuHUQRiGJTWh9qfXc3z05qisrS
DpOC93hnvZqnRGWT4ISIT3tg7O6XnOOrRE57xWOvBfdTFus40YrZlJNgjgwKQ/W7
l4mg59ULkmC7oLLKQCgnH9oauQ87z7yUNA8kPdURB1CMbqq9CY+/z70Uz+f2ejf7
0XvWyRGjjnM+Pn1DGz+XFHw6y/CnLN8ZjzeB63cQKcS0w6OXG2oKRpy7zbIY2z7G
rBLZyOT3fzpOYl7/odK7lIaUc3dGcMZJVx/4ii3KoX7Sf1u52/mBwnYeF9cImsHA
MIMAPIrHgIsuqoH9h744+acGBGcwBEgvkf+n8rnM51KtMixU265YqTQpWgjrFuJx
7IeUTn2liPeppbol0zrrxmOCB1TRDNDWynJAnw7ycilObcOndWqj/invBIo4ixj3
8Y70FEQOokZykegA48+FtOFgG/BppLAY+zsNU7SuWg3Ioq0nrKMoY0PUlsoX8WiY
RSCJ0pO+wPSdMkGc3l0zYGab61vM3TaynT6MZDRtDlpznqlUkmbdSQIieJ0Y67c9
HF+HPPDd5OYZydFEXMywkYde2AnI+dUKLZ6w+eZNOrvKp/dxMbEKs3l45zMhU1Dd
X1QqwmRieWUDdV1JNFbEMa5RoFwUg+jLLtJhE6UKFm93qb7ymyL07+0y4zy4iRGE
97JqpHwMbCD3bzZfqxyuJ7KpMHcgg4fQm9wKI7ddUjeMWZbs9EQaFTY8HNR1IHXm
vnBgYDSr+0BdR3lzZ7qCPf7vaxColY6mtX3qmzAEzbDMtqKN8+6vHQbgA7sciJPP
N2Cs/YzkG5odOhTWihFMnt/wneC9rO6z7sklL1/7gExuYgEUGoc3X3k7sXSYgp2p
jca88N7fMGM9z5pjIz9g68NoA62gTWNhSVaxx1nmYkb/v80dAhGY9onh3AIeUJha
lFn5ykdd3G/C48lXoFltbiOeAZrsWkxHXPGqHfsz1dMYcSYoy0u/AOXMwSxkA1K6
fEnEKly/GQIG6wdzuufdK7LafR0fWdG9TvnhBhcjqT2alAKQJUT82qPPe37taxhM
kXA7b8SznxBacRZFxjgwi/Z7zT4GQ3FLTZhhYyZofNgZhN7zvRrCiHKRGYHEA2sD
BKAab1M+PMecAsSnrVSLKVWwBqeQGpa396J7imzRZkzVRE0olXYMO7Z8ke6bbPiF
/LsLL0+H6ZzE7aboorPtQDenR1gsKgcgHIDOrzwN53PD+sG6gSeBKbcMHQaHA0e8
KIp++wInx/DDMuzPd9ma/DlvZVgiEsoIPLDtVTG1CBMosbhh5q2KtaOLYivRUUg/
fap6d70IkmNiWZZxydeaGVHUsjTcV76u72254j4TLkSO/KyJNX36qJ1vWpPUWSBu
I7Ycun2m5d/KKu6BrkfUTq8JTfVtOdwpzVgQeyPJL9V5k91bQ+diP/JJHy2Iakn+
6244EdMbKdjbYCNNPkNEu06AI6Dm+BvE2ETy9V34thdp6YFXOt2ejHCHZGcV96Mx
0rKeZeNbSLUlfkJvR9m4TPRTz5mlopt+4ciRH7faqnkJxuRmPzoIiY029753kWBN
nOcrxx2737kb0RO2eWBqwmfPv3NPawhGNDS1UczFt4WEhhzz9kCjX8pHgixzh9uO
i1lSwtnEx6dgl0H1r/moEC1hBGlsLPV/I1nyeFQHtj0bJ0eyguHRpskwRwQqTRqw
0s2DVmLGsjePR8XmrM2fJMQd3+LwDVk8TaNjXPGy5TBuWfF81OJ4+P5OdgdPZxVO
X8xwt7a+egS7VOYf1vpOG7SB9t+r4veygdZduuOhglH/leRrKPZnc9+/6sHwklFJ
tZjTtWyMZB2Uhvr47ARRO98pwiMZ5weXQN5wKbVWnDrM6YgRbhsWUwOGdhUblmT7
xOR8ZprAr61xhsTe872MYDe0g6ZUX+jaZMG8uHKAmDoRCUhTHfUNkgKm4/7f1NPD
vfGzPDp7nylIFrmZxj4uuMP8qIUrAjJ50wy+LZxN+7eN7OzVy13WWj0qVn07v01K
Nl8tKaq+tVJgbB4+NSFLs5ggAsnCg/lgXYvlkf+0aWEYch3ulUfZd12/7ezo6fK/
tP0NKgtea7LEykZNdo8aB4HP9ddSBSMh9NhJ0ZQOQWvmKNZ3skKmiLaDIdFB8dNc
FBN3A9k1wkZdVgMLvB3xO8aUUIn6vJNGMhJvpyfzbKWwnSRroYhWAhjnpA/mupnX
XGtGKM6a9gji+8uU3RxZP8u5uUP9JR0qexgfX6XfPwKzJvdMcYXKUucNFueEJg9s
o+5PPF3m0Tvvauqne9DqEduT8FqhEDTiFxNtRJeWRAanYRPWOV1Cx8UAjEv5YOnP
F3Vl9iy8t3t2tYmfWuW84CRep7WrUpPSblpZGM7+a6Dkat1HGCx7grbwqfFr8k5r
pb0FmOFmZlvpBM5jIt5lHGzrFLlrxlq058vXbMSHP+dysW/BQgvxhngtj81LIHDS
YcHXQ02pOSCeOyQsIwxcGgoRN9OoUGwNGSf8d1o3pWKybkRf7fseGu7ebkwHSJ+c
dDmS7x8Fn5kuFemVaW3mhCUBv8uxKgNKwg/BSXRP8RVHoavbcD4izTgOlimZJwU6
hRSh/r8gNK9vvof+VA1MYCy2ntMbDw4fqmRdR0IMjOZyl6zWQGTyDeQl+gjLSfXn
LOVJJ9aKEpci2ten3AzrUzzOizEka1iJO4mWBIpf1hKytJxD9zjCe1d6ZgebjkNZ
U5IJyaL/jeuIxU4OO0CZHK5XEG7TazTGru5dECYgURtGE2+DRRK4asz//gcCvumw
DnRYbuiz3KrsKlQEYX0TyK2KmBnh+bTznNWSvEZ9ZwLPCX1hnknDj9I5xMfDOrlF
huBYcq9CTgWrUCc3WpLrSV0pgydhaPsbWgfDevcKoAYnD4v8XcQKgKOh4OSwe4C1
hypiCtgAi+6NG2v1C1HpCHG8NDxX9dCL0pZA7/R9dWB0NjxnjBVEgePXRs+KlnNC
x/9sb+C3DdNo9no/p9EM0A5+OFCZ1syDWBIORu4ERgQV1+MN8OdbJzdRfUlzWL6s
6ULrZ68uOQVuY+h28rJoMpAmeqSlQocKOVEU6P6JN+LC5uvMh3y5dr5Fb6Ln3kOm
BxOLmBRJuYifC1Zs1ziB/49e+UcEkkv+VsEo4FEAqs8rkTm1U6iIjOFMy3HzHc+o
jIsU+wVkbAZ2Iqli4Dg3MF8VauPd7ykiWT3ceARc5ZEeDzNUrL5Pp432nyBH0YEl
2NjWvOV/ygww+X/NtcvsKUuQsyPYd7rMdH3xYgURz5CbOdsKQS3j5LJmMEtTC4yv
ChNskrtZ1f0oGGDCaYNgGTn61iV9onP1QzO/EGSC0efv2aKsBHrPtCZ+AHB3MTNw
HoRX7dup/LCg2823lj1Md3U45H1C6Et9O/AD97zQCwxZXVtW9HEoxqvVd0f9EwcG
ExeeDwJebLsomX5Eq/fWjv+dS3P3DKI0/hsgeYIj/ourONH6WL6+yiGLAuTS5LHf
wS55pMsWscnlWI14CkBSp71XP38VOwhyzSwVgQMDi+sT3iDzPIo6FGeQpdgNYzFO
dSl4vh3GlgHS3/uB4PHkQK16akNv17AOE81GUwN7xtG0vuKcQZaSUpK1owiyiaZN
l8guidw0k+ZzykT8P2xGU3qd9eeti01qxg2fTaeOhYCxlVWneyXVCcEeWZKo0Kzy
L8ke+a2yGWTec9gLj1RntPIX0KGr/zBs3ifGXtgXTc2y52r3QfvEulIJDFvQZ/or
BWINfBNK23TMwaJVQH3ibHPyKa3OjcP+lsy5/MUxnEu8X0O36iEqecbdHSN0rSsa
/NhDzcxO2ymO73qnYo1pJtySy9sQStzQ8N9AYuc6YJIuULmBf5Iscrq2AAk/iRjW
GDObHmOutRJFNCikc3GfwypU7y4BO0GNf+bfDWL8+h3f0TG7D+F+v/acZtn1sYu7
gGEC85/zZTnDUupWoNCmnBiPDfJrRKpNK5J9uDmoeQFqUN3fkvwBR46bTKpMXd5C
le7IPpPwtJd6Q4LKH+Irnv5pNxOJIMWVovmzciFfr/WZgBgPXXQsObQ2bR/yqyDc
3+6pim1DFM+wSn9CHRaptBfn9blp/CFeSXorWkQ9FDrmeUnA4zbVqgj3g9h5FvBO
uOqrRaAsW8rV/AjJwm/vjoMWd4/aN+CxXXAoFIhtVTDr8pXoNeNt5IcxvYTBL/0s
mYYX7wH28E1j+7RKchPUuaRC8ctmxvbC+hnGOfkwvvkTscw4rv2FmFXpXQ1wX9TC
Xz8m5IMag/98mxTvwS9rMjXHlH0OdRGvEwV9gkgbX+xmUg8WbYRakZO08hcR3xmx
qo3bgrSr6wgZoxeBqQcLyRsnbJWZ/uU8AEZUvXnprqsmOnokzWIBZIxqLrqleU8Y
GOWuVgvmvsYJN8+wLzAxeNYRf3v+YNYNpPXmpBlvjLMMzm5p31Sy541LWNk8dwKn
1ROB70aWgYDSyS5eG55rwcCRMC8ol+MA47P7nghmI98QP1pW4FC96Z6lOwD30UOP
M+FEPKzHM/wLfBQuwyjJIxz9TB3CJh4wSUz9FcX+EQaR8zD+LPKeQ0EDNFBvqupE
t78QrqO1A/nWGhivU0MiFmvlgby1geXGl1AbctwWpI0J7D0XIiwfF3gRe58InjDC
Jq/bMIAIbDCTey0MqVt10KDNyViez+HGnl5PP3oKgADDX6En/M40eUrTq2XMGgc8
+bRr6PcJYDHEyVrTup9Pi36Kzvi1BZbQqsUHjm7P35pneRdjO8aDBKWPLnxWoiKb
FP7Yz2a1nry/yguYGk2ghDWPenDMIKC5STaWyajafRsJt5lzlZULmHKBX2+1PxcM
yokGlk4V4rTA+uwnw+UfZ/hmo0hq5YaZ+hDyLLq5fwV8gxh/DiFEJCcR1ksKj4yL
0B79Z9rqP9D3nq85Bx/jl4TaU5uiVVugOqRyXtAsAnuEzcrGLSVS7SA7ENOrNoe5
oOzngQUCp7A4X+2vA5QH5nsKgxXmP/KTDtSji3ORhbqMHIfa/RN8Efa98oTfzr59
+aLQwCdwrBBddZV/knMkONPoZNImoekTCbgy1DAr83RnYqcdp3ocT0A/7ohjH0uD
/HSNNkikNerq7NV/ljkP00XrTbk2fNwzFht2noQZUrTtJ2D9T6MSzK0wZbCdv+KY
+xTf/XmUM3NpwE26azbML6i9+UsHnqPiy1brlVQ5iK/EaD35DizU3UobxHM3T9HN
1/2oS+OmlIVA24PDFnCXc+PGOnXqwnfJruX5F4PIAk6h7XGTimd20SLxzc4wxrAH
6FMpIcijNJBETlZAXY/1wtCmHXqnFXtEWq47HcQpEPMMaRuAzX/RQ8uZSe6DcAYW
GTviJF9BiLytzjHA6PgaoTLySaZjytqD8h+PAWvatjiGjYrnXy0l/t/2yFXJokB6
x+NwexnW5ttwC874gQnrDiI3ep+WfS4Bwbw1trx4d7AkR17mdfe9XIRN8SLNbsKH
QQ5OEG+dC+tDcpce9yASkHu1YSxAPhIc6AWqkRSPx4xjmfjMZRXKmgWoE/DuQ4/J
QIoRun6MXbdyhNb7OooS72pagxipSDh0eYCCxZp3lpaHr6i7GtHRR7JmXTLqPWQP
cvsupDLeyK4dAUOHerdKJtwp2+/x7XoG6bRxIucdTk9nt60NRqLdy+Y7E/p+lKvZ
GJBCc4lyeJIitZ6dDmHUE8Fp5I0ZLt54nL5SPEOsG50wODfabv5uv8MCSPNCfQ7H
5GnQbSaJjbwqhjXTTR3DSXqsNPyt+pyYPvoLx2mchVpeoIWe5Lq12b4oEBF7uxMz
thPuwQ1M/twp+ADc28OoezLsGjQG/Eakgfb3LND05pqOa7/hz6VNxi1X6N9fMcuO
5jpWnnm1J5wQOcw7ruusN/Ve1OxmXKywIEFewbAp7gT2gpA0GHyeYfAMpJ04Tm6y
WP4dm+zEFDkxP0cWjpPGMxH7VrUu8Uf0JGUhnGknUas2d6cYKYLtvdZyqr8t/c+m
I8+2j5+X4yU7DYxMprmxpwtdtLYVRQ4OH+6RPqMPaW9wPa2/pX3Am7/mtIe9XQXT
n8p75AY5HzSiNEQkJRGfYsUyEdrz2s/Fv9TQs5hubMNtY3oyQgYL+l2Wb0D6Q6/O
nbWRaRPs1JN6uKf36XXdja5bc2QaM4I3xkQ3ZzjX5TowrmFnTLvNqPhlcdI/bMAZ
3retSxMgSlSa3KnaUAPhEuvlnfmTIv2UA9elyh2zyRBa9i1Pe+0plCvHyGaHweg3
0qJ1kPn9CNCwoDrA9+5zbBxo91nj86tqkztOVfkfKyqFLMjnT0iP37p42UCtgbkA
WmWE9b+aACC6piFOxVVP2Jx7JdgTefTvoCzQFrKgWJAhuXsPtULj2uHc+VOzwLss
j/ZgGgnognLTbnRyBIxZ7qNP5tA0I936tOM3U46PxK+b8Mcc+lziVOWeD5CapB8e
aU7knG4/i02p1IWl72kl4PaNiX6CExEe2s/ggBphDdD+vblwUJ6AfaxvqZ3Pjhdm
EyLTVNdEIJw6q8DDVyi3IYcQbR/KNdRD8/+sNLBRqL3aAvOSryuFGAb5m46c2Fr7
iy9+1laBEdhpVybLqQEmIY+MKA1aQ+e4hSLmarGsTbinLGYmEpx5oK2dNhUWM8Ag
aKkZJcdI1mcFmB+Fpp3cKlj64JYxKCPTWwPf4tQpZO+ZY5lnwBAHSjgO4lLKbDE5
8TnZMrzegS8JEPVOyQgqKJJG9XYVaLVQl4+CrDnYLYIbiKIbqsEohuCha0XPyydt
dCSI9mHIX10HJ730B5X0QSyT83Uu4n8gQW/4nvXF2JpU6WFy3yZSgAEIkAURLu/9
k9LJ+XW6HKSZRkwxwXdIPfQLynMAFyLg0G9SPYV1LEOqMqbYseIuEt03FvfTRAZY
VXnpUbcq5Z4363WxwmbvbJLf0S6SPCoFahS+tZ39MYffyJke7lZ90CvySvpy5D0I
rY5qOYDZvyOcmJNzwqwWXoPhLptfSBOczsHms+nkRqqL+1VDbjO+qkXDbZShsJA4
fPDdmo4CxVXwkELl0JWAO0RsUr/nFbDF7d58sVMaL3EfjOapxXyvyMkD/BTH5bHD
K3POiSymRKVMx7UnzRyHhAjh3oqcnDRzjsdOdnIiRwSzP+E4U2XtA1kDKo3ALYfn
Rvg5WkA4G0to7JeI1JVJZlgWXAxKsmBmJRuV79aJure19VeKT0o5Ky/1n2N23fES
xsMDSO6qiNIPYSDpu1zWk4fwfaubADArPuqfc3w1EBmDPKwAwhYLCREgSeescbop
kDZ5SKT8iFc0gJHOYROlrGOYZ9Ecjz+eRAxalWITyBYWp/RM5UBnewZChFsNUoeN
SpdsuF6GReI12HnrKoZ7yVLlZIoh3l1bnc2dg7j+QPaxMZvQsEd5bw3YCFH6gFZS
CUOpV0WGqZz4e18al5VJQw7XyDZdnfgXOyOR9Pyb4O+M1lBw8zU7pdddKmRKc2xX
Dclz68AJGq3SM7Z5l8edRFk4EDYiqKBC4ViIvs/a6ZVuZ9FvFyFgyrZvF0fGyZ17
X0OcO4UbsTGAS2V+ZkWc+7CYATUpQBt5rgbqFQpoYLYP10Wg/v0nW6UPdS8TjsWg
zYgBA+xBGBycNZEghJDJufQXJjYjcoeSyez2ww9X8U+ztXsO0oC0W5FwwtAcHwbT
43A8u63WahlcXNFlJMn2wifB+LJNxZb7t+bhLbtiuLyiZIPh54rpf/j0j5q1R4gc
4T4GjKGhN9vDJJpLvsVx3XVrkyuI7V8CkH5hJAPNL1kKC0+7M8WFBpET9EjmZS4o
L4CTYaFF4Ykh6zq5Lc9mM/1inz48J3XvXuxgnVgZ8UVsuvsp08H0TfZUgLzdx494
CPlgFIFYDpzcIHCXgeAdJ8A5DfvQw0yqfiOc1ffLzRtYwi0FYEwBVIqbhdFI9Sr6
jQVBZb65+f7unnFykvkv7L7giRbw75DIbrAbe9bl9fnUzNmmKcknSm2ePZIoZKlH
Uwh/+zLUeajEasu1kwS49+jtvWRHyKK6FOdFM+bUbgfv72csVhtZgIJFw8snwzMq
vqUFVAlcJ6TmqyLo5QFm4cekozinLo1zzbitXcE0xRm0pnMWKuW0gwtkUl477xYT
F8IxZanDasfGrpRwEXw9zMKp/ntHSaIMTUbLV4PJn/XyLQmSS0iX9pVIMgNuK4p+
MDqC6jkrTfKGxQh9mXlAtlDx0NFPeMHsjzcVVNzQOOyA2T8SX92lvg8Zh+YnFDDn
dkAnpRzu6akMqO78zT59LEItJnoKbvTwrY+DAUAmOW2nr7pUDnc5AtocuT8vCftf
eNlPxYbKb6lHyiRwJ0z6k9YQNSR8Vk+fhtwJHorMN6x7DpZujbquGb5uk92+xdRH
3HnbNrxJrjNfXmGse/ykSZms/xRmJBY0Jjnon7j4uGt9f+xW7FPPbUD8wzaLHkWe
DwLfT8JkZg9T3m4C6sPa69SlMPatgRMunNPuL6AbNN2VjFw8Ltd65EzqR1xiJZYc
4H6soeo6FFxbTDlMw1F9i/j6H/ImMecP719fYOVGNgGn4/TaNMwS54v+IhrUMV1g
hpM162nxebyOkNQmCuZTKEcTmLov+DFoxo2Kwu3UmoXZAXF8TqH5vdX95XfeK9+Y
8Cv72eGi3d8PuKxgwblLifOjLuwFjMO8lXLGU+8SMsPpCvPgsRvsCjHZxFO6eSl3
11ieHJ+3FShh5LY+ogEfKShEa4lxZDurwR5WCqpMgBOoeZlGrgZ0aZ5egRPiDZGo
GGEh3IR79UE9jddLf8trD1nVx9wCKz4/4fv4OhZRsk6vy+W6HVCGT5HAm6eYNqtY
Npvf3LyKCRTy+Ruq6vU3pWUbe9ij1/q0uSwdNZP1Xo56LyhJx7+lR+psTEJgDTvJ
MHSimjKPHW4od8TnOVkuSWt5BAp599IWbTkENz8cykcyYVQKZuYDjSpTCw9VsGbn
QeH/4+wzlrnxGgu2FeRKhIB32brwjKYwox29FuvwMC3YTSCkKgsMLEC/vaX5l3UA
/O/NwdJJxQ9K8esHPgIA31berFniKqUB6EdT7DjDCbUQIIPbcH89oh8iIfD1eH9R
lykQlLoaawugZrcBWDijP5oTIcR66bDnvyXBArMk32WfWCJZAaKJjRchtFtFy6AS
zRxbUR1u75l9RztQAH/GVlHYgYt7oZe3WjokVCJ2fSVH7qAiMokQpbCdxnFTvycG
ceGPHudyFUKAFhfm68BQYqB2uTxxD1Rpul4dsanCxLJZSu2So7ezkmJGIvXHiVg/
IOKxSbDl9F6NgrNcRlFxC9l61xtqUcc0YDhDcKuNOSwUytjgAiiXiYKSG2gnd7Km
ffVEXszK/hagMtVtcdd7YIbQHywb4PqFgXdsge5xcSOecQ3GZVR/jHWaWGPk1u3A
CY1jcmhYVs6w0Rn3XajTY+UxOaDuZYNnY6jfBg4YCo6b/jsxHGOzzcLkevG0FFuV
ym1TDY8MiQgKX2+NlCbwo0bFcQQoHENy8vGWLzVxRL5GML4PhNlGNBt5XvUeRLBT
r0qG4RppKze3BlrHI1zpmuE36ZgKUAeLiBgufuNgUSDxXdUrjrLtcbdh5zzaA3Oh
iHCtON5Rd6M2MFy0JM9Y1obTtiofaPze8trfE+BltpQT2xui9+rUQHCq8PjCBO2a
YD8ZXbOwmZSJltYq960EaI0Df/HCmGkVyzzxXcyXMB7thXCeih1Z6rhxXZeQ4sqi
DYsLUPbuvQcPJcdvOcBrtZC2DO1r1MJxwmjpFYeTZ5ANI3fDQDtWC+VNpwJtcJIH
Ur1dIthYolk9l8RlvGDM6LNdodcfEH8vK8+Fsofk6CWfGwDf9g/fw+VyTMOvS/7c
XwdkBF3zZ7imk5FbPXI7WZF0BMH5sMJEI+4ml2MhDW/gb+jpBumSt9K8uxtpwmQm
kBklRf6J9hLRKwIq9QzvcCkftYY35ICUKx3ZrEkAcPtuAvlqlQXLouT27Vmqwymw
EoKFD+BK2rH6hGh59fro/j0ipoPAAzo56iZBGQQXDPvw1s8imQIFNEg2R9AiWDUn
G9s+uj3cSOFYyBynytmIeOg7dhS5SOKpbnm1YPajzbIFV8CbEcMyHpfw+RSeHdPO
kc9nIzXxc7Vfmzv28A2BNhiputKRph8eN/J+grB1LhMeXsuWN0GfWfvzfSQaWqou
F38mdlqHVPs3bXt5Rtsz078qhNAhqbK29H9LISCSyCTziQg5IOpFltH7o2mh4iQy
SF0ZqF1gxYSKgOeJJGhKAG6zZ7ngxCLlsgkxMyw+A4In/ksRRcVzAzK3GaPPeMi7
DRgnROuNRmEtA3EEvSZXCg9HXWRsE3q7jEvfujbUPTwLSMy7WKXtK1esdPUzFf04
+4bgaFxUljV9hC7emjRa/g/qRNtaPlpNFuojlPRoL99SvtPCISODCrfeM8r4Q/B/
/gHhzVfCoXVU/dljYVGXtZ/LabuiBW1lEYyMzyYfI3ebD8JlxIUQLyR/bq005eUQ
xofFqAVKve5gX6RJS9Ep0kCoe/imtYcUdPwSrdonpNpX77d/rdLVuGtENzdr6sG6
Flaq95nYeybBj77LjeKy144GuxFbFFmAjo5G7U7gdQTWYtVoPO9ENyPzrJHu/88b
X3EcJ8upJ33s5eXOZwoB0MzGFqRfh/QImwNx69znntPifUjfDCCxbirjQjqLGijo
gD4HpWOiVxzt4Coxyc0h4Phq+8DwjLpUhQrxquwDT1ZSi2GUP89V+0V/i/oLE3Tz
B08JR1Rsbz9hKQQf7FFmg5qOk5ZVSCTlJHHbTn50vK9DkFn+jj0SWEr6QAJ4h6Zg
GHGhv3b4NaZRePyLDHugrynjeIULle/ngeSDa16XTqZqKtZiQ6wuj8zuL3rSQBxD
L9958ATVeVi+kRNdEKFkHy9Hz4VsvMV0Eu2rdGTKQxzpEtwUPq/inn4F3qajX8j6
xlFbntu0NI+X34xInJn1SwTXb3EeE1py8KCiUxqhdYgZ2CdOgUIU/xzqmKEzHKPo
FFXbqmxcG2RLbkdQ2NmAhEZSu3ppkmDebU4LH31FAq9pDdtot2iyOk7OZTGD/pjx
V+OQMKtVntgz3SbAtUFeyUp2npQ6Nmn492ffTsXAqwsukGzVQrcrdWoKu4yG+U4J
e7MV5Yx2To7iCnNfM8Dw1TnDxICgOZkEn9xHa6yN5xtZ0nEf8Owh1AM3q99DrVoO
QGqSvhXs0rNnwRxkyj6QDYmF73ts8HKOu4Ad14OwHtHb2gKzdw+dgoXaEnEy7VWE
MN+amY3mQ+DZBRvKvf6CuBhHaME7Ksdy/l512p+Gv6P0ng2rpa7HTtE0qyU1XA6E
iqCDfFMY/pmJS5ATDNNgSgPBPujrFRgt5hhsjdPR62ODSGHhUk7VXX+hFsncahXu
jh6JNI0cKc8G3a/pQFlXMmKi8/zC/H5mO2o2OUrxJ1bYRgpc83X8QPekJtziTQ40
DZZpsRprZCtOjOp10+bJ9qruOggv/E2ym4IR2TXGdOCO5u49t6g1UdEdQWVV6W31
DesEbw4IjW5iAaoSwUsZ4/XGE0+ZSzVe+rneWMXa7nOWSFvA7z4NEsy8tR2ywWNr
YFd+NQoD+XzWC4BrfePrq5UZI+/cik1+IyPMm60L4d9W5Cza/Q5jBcn6rwEDd4nw
T8sAPyn50zCQtd0GcLZbLGq9UmElHHDnSvBKYC5m1T8q9pMbvBeItZF0GO6jfXkJ
u/heVPcIYSa2I8Rnb4QpIjtvH9YCj5nxbl/TWwGXnHD/zcWWM+MiFoPTHWLHP9st
jHZtH+5+gKVjNcAoHF+U/dbrchquCEhdKhgIJiI6vsJE80WtxwZSPi66Gt3YUgJ3
0hghMd5ILj7W6djT2XWy0A+qS1K6+eNTzhaP8IkhRtBI3/ur8N8x5sZaQ8VhN7Ic
dNTFm8K8EvW2xlD91LcjjEEMZn+oIdB4kUIDBdlktk8bRZ8BNCbCCctskceq9T5E
5SHfp3lDS8MpfwYoyEKJInQ78ljgNOp34FL12ItlJfAYmJ6NeqNzA+I++1iLWWKS
fuWnM1qJxM8xx3Lnz8qSlt6VLzQ6JpUIYsEEfZ11OQ+q0gkXN8TP2pWDP9R4sDlq
1BxgCMghvO3WqpS+A4aZy7D3ZK6wlMZ4sj/Ixa4e0cHIYVMEZhbskAGL/nqzMvRo
OUZ0DldMNWK+AMfJqraZ+6UTLOz7sGWXmJJkGlDMVoPbvdVnOMWVGv1CDTsu4+TZ
0uUR7SIZbbwRABu/7eaGwoqe+s5k+P17qkWqyMDHxib/xaKV0ejm7okrGkNuhmhF
0uuH1+wsFsO+XchbAb+auQ4zkGOif2+Zux8IUW4C7fq5c805R+RGW477pi1sf3Ne
4S0QqdUgeKZ6WKAkoOMeSCsdBasmSDFX5shMmCPyvXZv9d5fljDdaPLPHZOzyNct
aD9KFkurh7QTjoC5/Agbb5GFHyjgXmZwV8cVAlD6nfQ0lHJ51jONKs9dLRmVAWTQ
syKP49eMKDqVKyStMrPCMLv7McxA9xMEcrQDL+3jn6ulpioq9INSjZiEcJ7VdeX7
FLTu+GxSgy02MV2J5luc53ja3zCjON+hLUYvYKyhUwzfM2ujpQbCxrG5rARzMFf9
YD9PLU93fLmenyA7KKTDv8v3bogqmZw1eJ0DgleUnglZ8ltr6mwslH7XYdIQ3FZj
TtnXnA44D9W37lQGK2W/m7VxJ5nknmzDSrkSFAVy3IVGpqLu/Fag2bPe8tOpR0Kt
vanRpLAqiENnCpQKJbTzVKKhu9Nd/oI4+GfLjxx1b/2cC65My9niJcUgjB+0rfrU
OGMetFdLFjgJ6OXfLCQYrdGJqR8ZjcdIvIH965JTtoaFuQ1lY8RSXgtuHhLNLEut
qLzktVppPUjwxlgrkoKHF2pjhYKhvtoMK+kv+1WbjAyodRVEvjpCg8erj87kDZJO
VcBFayXgvD64dPMYpAdc09iUekslbPfqyD9JYPcG+pJrM+e+l2HlvNru5BuYJmdy
2/4oewaat88hfC/p6eF3x7MLcQkxNJO46+qDsr3REnP9UfGJaRim98TqlZ+utnqJ
R1Y0WiZHCqpOB455TOuLrbWX+HMZrwvXdh5Z1rby4zGn6RpKx7UOzV0WANhignyM
beyJRQiwGqj4FmtMRiwPeld7vQ0TBIC0LYZQpU7TpYCyCWxfb8Njy/XUFkF+zmFv
x7yA5D93hAjE1O3CkGlFgOWRLdWKqefT9YtDpHAxitaBxn/oaPGMhqvJluLzdeVO
V5YvRT/aVpyaTfU5Miyt4Rqbtn1qP7vuvFWpuwZZkdMTvo3wzyUIq6SKmPGWf74n
7zN1xe+Lr1O0OcjXP7xSuyeBK2Vkpt7ytyEoYpsvY6p4LvCQNq0zgn3+fPfkb+MK
6gJB9zE2pitxU/Ut4uQvdTBZ9TGgu7SKYYSvPhibvwiQVtb9Xr36mHDFXz1Cdsvm
dU1Sh3bSHMrk2pYgUbNhvMkIidGEdMoqc467ZCoLNx1vvH+J+Ri0RWH+Q6+Dopkh
aTr25KShVyIxo+bAgaMuAqThSV0y8i6OOy3B8rBTKM8mwHGt04bQTUjor8M1wSTa
CCdgrAlXV1r6JZ62wblYxaCpWcS3/0KiB97+5F/zuMz4roLWsbXUReY0g39kzP27
mXoZn1j4EaZyG4UBokYrtPfnEa677cIPX78JQt0iTxtmclWY7PGy5gZ+AdZ3cQvR
qMXNxVsXRBfD6FPsc/1myxmfVROhb6bJPKgc80FApbJfwEEBVgKJVkp+eR68lgX2
DCiBeEPVutOka80NBEORB2fFZr3fI3mpbRvxc5uXWeajz+/v5nOAMuL0WWAyKgef
U+nVinVpQzLkqJcJM4GsL+Dn7mDx+fmNzX4pX+HaJfce/IV2+hJlCQbnhsiGVrJn
eiGNrlobY/eT6wLSxCQhtlJ+1Yya3DrZdwhDfPPiCGBqZ45SIWwkMNHur18lV1br
l0QmvlddHR4dRoAWXCPHO5bqLs7N7F3zePnwmmLSXM6S+jn1Kbb6ZiBAhtSM15/1
XmCTzzooxorq8D7bSmJYwZ7JkIkyoGQCN8PLyncuJO1B2t7B7QnA5ESJKo3ONGVl
iSTmNeQ3/D6EsLz4UEazpW5+RAR9IGQSiz5xZ3fJ2fVqNwEch6LwKT5YKNZsccK0
Nh8PKZhzrUHhvi22bcg6QDr1/WKpSKrKaEjlfS0gVu1WK6XlC2geLAff2zaCwgqv
qmjgDwx0Ok5rFSMC0peRgp0YjllpLLYQIEpX4rmR+7khl378E5lBENrGGYBf3dAx
uEFOpM85t9fmoPThrqdXCRCF3RyAZ4YWOxfZqjmVLaBkAuqBpZdcHAfX1ku6BW8J
r/5OwxR/iMePsRXs20M48U8+Qhpl7GM+j9wplinq1yXRQIoRSqqdPBMdUpKRVU9T
S8UwttAOhS29wGUvEWFaogMQ0skzaw9yz/hlz+IEWWYk/nLTb4LGiW6onKTio1Q/
Yqb+k5SyoXiSk50rvENT7ugZ0AFanhRubo5a1pETq5kNIm7nvwJcyZBW4eeca8W5
GgfgRhqWkK1FUqJjYlnbWUShkxW/XB8wRk1ddP1rR2AthIR94TDqayJdd6LfrH5U
NiPnvp5BBRNj1F9DehS+6+oOz5sgTkDNwzqD+2BW0Ps/Ew23q9hMEEiSy70iRWtB
E7basbIPck47ZtyxDjLDD+FtVMAmbHw6cZUtqDVGxc03IkI2iGWM/HJkmDeHz+y0
U6GeVsfohjEAAY3AnNRiZK7qaf74y2+uISGyjWv+sDfoHyCf4dmV7zcVATWHKQ8T
V79Us6ITGBJQrYrMbUCtb0qqP+TsAwWPtrtw77g1u+tCtyuFhgCAtYV3UsM+a5Pi
RhmW6JuYVM0o0GZN9GgSkGvGwyKr/GstuygPFPCTNN0bycAkPGdI8NWL8ZGzwLNP
LUfdmEZtOvSTB8mqvEQvQIV1255x7hR6pb8M0BwnnmTaVeOiHN8Dl5+65UONsicl
AAhoZl863iUj0T/Dde92comqZbUslBjPv8PQusQafX9Dg7xrjHOlVmQ1ppAtN5l5
bJ3PBySwhZObx6K8yF6BraaQcL+5JFIY9UroFmDirwU4LmrTRMHmen/DCNnY8LR3
A+SHHf6mMHN2KVgbL8NcYUHgF6l6Uo6gBtZGw3uUzvk3eMcuEzksaRR6pxTeg/zn
puqFQkjD6X8vfKtYAKXEdC75HyZdl1F7UAFv1Nni2kxfdAvuXjAccJe9SdjIbXDg
OzEU/Jrtb2xYses9GjOWZTJQjkGFcXeUi2fqnj8kal6W6E5i65q9GMCSRBRZbwfo
lmjbz96Pfu4L5UodNrF9xHcY2lsbsseypkWVyIMFeJNfVdC/jrb7OAEa1oaOMEyH
qxkfYFRP9fMDWHJH34N+nUotKFMExmjPAdc/0Ni21Wx/bSFtBqvW5eePWapYr0I3
LJlQ6hY1myredLVdW6FAJ8IFfICyakX0WoXhLxJcb5ojX9EvMImQoE3PGJagixrV
cRraqLvJoCJ1wRYU8hhvd8C47rYmHqvPXdivQg5BsspH0gN8DwTKFLA1WwZJiaTH
mfXul5EoHPK70WCsWSY9XonA+9+AnG4CN7RO3ZmyP32j9e3vgvVh6Ic+OyZrBoQh
3DfzW1u/4rb1n/2Ka8xPs6Y5wk8nyfnxG5IQuGvi7zlV4IZmfPs6wSzuIsM+K/g6
KDiua0cGYy2MXtsGOfFrEfM3tEyAzbkE7y5+d6lQ4mz40TXg52G9L2hMhVYcmVAN
NO6w6GQJFwS7z7Dn7Y0bp4azpYhD+3d9q7OW9sHdJuhHTxMtjolTdmcRC7CbQ7K3
aOTnBOmp6DHcZA14ipB2Fp/K+NM1sh+ztZprsDcOYsdnwh55Yp95S7WP+8+hIdmc
D2fhJ2w5d+2MNSTCyQcLQUrxcL5MKb9uaKuqPAd6x+F53bCqmxdGC+IabSQ1khJs
pIQLGKZgidcsidJ+GBlkX77Zw9GSAGSTV4HmpKjrKlVXNs+2usbiJetwcXxYoLUF
ZH8DPH2jR8mCrSQCP0kwXGswjaOM1YdZvCNChxnX0U6nu1ww57A6u5Du5Qha37ov
7amKmJBZyb4mTLM7JCJPrRVZ212URsnN+RioHmSehq6+72RA86SE258ycvRrZQcA
eJ37Q0jNGD+QOq6+FK+5+2Uu2jkPzM7ZRGE7vJWPivmzSjOslauQeBPJ6/avpdqG
OC/lTFbKKZY3YqMU+3zBWdlZAXJFVb0jQx5R2Vs/RpjQJdAs99nGwt2avRVmWbT+
GRNb1kIefgqUdprEDf8yA7D6IB5C/1cHX61o0v4NbmdbK9wD2KulX2jViR/ADnCs
XMwEGK1H6TRkmG2H2KTbmx9mD54UVdRQj2ykkVcFkPJJFt0cbLVm5BujOwmP/ynl
22R8c9F2vb+wCFhGiNwzRQVbE1ei3hf0yyklcvGkRybAycoLOZqjhO4BIoxPcQtZ
R2sCVJNloe9kB+4lv4tmtcUdjfmpdaVvmd3KeUm6t9qa2IzCI44Fur2KjdAcK306
tupYlQ6agqPbL6kGClbexNSytfXZ6u+CMxZGnyqA1gYcvC8g4Lcpg9tqJBI1BGPq
Bb5jLi+t2yMSJQ9yKVh6RBS81ao1RFr7YZ9NlpX1RSkZpExSIUoDWEz4pd5joMGL
0GeX78dBdg5KkHJeUSXZ1w6wdoUcx3TdC/Y1wk3g8dqz9HSKazvHJAc2+XPovjxo
9OOjbUrJx2INzeeG8JK0Pf7JUVvADMiiuSqPL7zYKXCyA7kiLACTZybOnpfMWhic
nDc0A4hI0pRNBHaDV3nIdaAh/D0sWRgi6JpA2WMmR0mgQ69qOn6h8q7Tv/AFBjXp
tcatUhhIuTAHrwOR1yYwSwvW+WI68fCkA6/hliM3D9/qNUXMkR8RupZC5PNxD2eG
PdLdnrv6M2trvr1ilvhcqBr7pCUcq48M+oJ05eS/bzLhJ6VHAyWSZhdIXE4ohye2
BX3az/mUoXwi861aJrefcMvUdZLiDpk124TPpq7kjKa/q74OEgFPzAza9EDArb77
EGlA8B59LnkUs4yZfbBefL0d8QsxlE+en6Jbjr1JDC9gZROz1v3xepZF52fSqRzI
+8PiROWtGfz9dEQRnthX++xc9sXbmp+ODBUx4oglzmGPGPqDvt8M0TaR17hrrBVy
ZBBe3nqFyd/XVoNFSEL+PuG2uwBpnd4vvQXPeHl+4q2kNxPa+nqcNhIbGxeknuoj
VHtfZq02UhkI4rl+/Lj97cz6lcPzkUYAVnaArLve2xAqOeJSfFHMkJnbKMEqBcrR
22+MiE0bqnsxv1rov1+xDVTLeD6OC6hwWbT4VN4JLjgcMyg40r6dNgKbduyA2IPH
VCmcYC/tYuWzgfLTLuToqeXrOVR6hHrTrGTWwS8kE/dyiRluXtOoOpA5IwTQxLpZ
Xyabuud1mjfBwfCsNAgXTjM/1uccAZ/G/kggwz0Gzo4mwODMiC6bsTcUKMAwueNr
2m2z1zaO20hq9ZzgqDd/YRbBIYD3Jgp++IvfcN98FaEgaFHIAUSAz54nCcOjer2Z
FjPIwRRRiKmmwdn3Fdu4PMGyZG5alkLKEp0YY9AkAVL9l9NVd5JNQlMg8kEkSPYR
TgCx1nJwfPM8NI7mMG7AGiE92fUbVsZ9FImUouH7ipJj2b0/eTmRSk83c4b7BGkO
HaaM8w8eHCoH4K5UeMWARS0KyL5+LcRjtwZyt8t1Sb9iGuOLJMarawTbbizB8JG0
SYIeZKAYExoISX3Q337pGHbXVvCv6pJtyyqf2yZ7QGBQD9+5tlZaK/bc9q8yodpN
9JQC9x1mf1TEJikImWYYO6c9HlU1ZkRFD3S2WyzABEYMsQxnNYhTIIKn4sXr2pca
CpmKB7W/DIWyPAF1tyecmzlY2h+5dNh0Y61zknkmrs+bokTCeQzR0KqqVWO4k/C5
DTNjgczsZg4msQw1l/RD2bbk8vLXh1S00zM6nqFZJuoe1a74M0KvG1HTThshbu1E
slIwm/jGW05Hu5x1V4whyTUiZpGYW8sdWO9wcpqiK72XUxIcaATX/4GMJes81hV7
ORBIx4tei1VZkU0tm9PojUrCpHMW/8t1J7DFeF6cK74Zpjtmc6wCE6sDL8HZpFfY
rhK0z6vNZ1BqoXbVvZS+9qWNVSXZ/wsrkHH20DgswvCwSeyzkB1GHgejFn1254Xl
zUn1w545ukQ8QGbwpJc6+Ahpn4M6RgGpwKfqNbXYHCkt+xnuL3YHOPgTLDsRUBT3
/eZpTl6TZekqRAq5JBq6iajOsywhbZrDudsqi372vUv1WG+PHtVpQIFi2THogaOn
JL/Nhmy0SDCX2+BAwNz51zWC30nPzFgC617UOUvET+ohqS7hPVMznCx2QbezT1s2
CThe/FzkTVk/cv2D4UvOW5iFXjPS89dpza/q5kjsTijMzaxIgL71UFqB5c/mVdFG
EvZWmRkOjXo/m8Ki9UTjefC+sybYSLjRqE8oor13VpWRlZ3/7S/YGmx3R0Kk5PCL
r0Ycp9z/Cqfbtu7/JURFUjd09JpWOZOlXZK0vFiP51wQEPHWzLOofXyW7iUdACNz
gL4S45Fu3z4mSv8y8aqkT8+ZuUgDD0ptuxIMwhZDn4sM49SRZdvriNzvUDnwHO9L
MPt1GdQ7owyeIIcY6sB2gJ97H8tcUfuOBbc/8bRUe8Q8tN0Hkb84M17rNtCUdgHE
n+eFYYbuJkfPN3Qmn32hfnfyu8csMOXM5G0Bwy3bHJlJzFIRFVDVGfCWQc/XRJYI
+xR+UmgLRBxAM3z7R9gislj+7EbGQPzx7b7HCF0/pYvB40aU7uU86U15DH+swS0s
vCSmNaufN4BSMU4Ub299WuWkRFOoRwRt9iwDyumSycDFjAOMFPvCTrSWZiWEkOOi
PD4bAwAtD4u/2CD1c0cDAt6ahdYJIzEdQtCJgTRCvAQLL10t3glE6+G7n2XsdWOW
ExdlotrOARBYHIcSFYl8YqUzzgpHrbntT8Scv9a1J9SpPPmdtNvFL5HMA9yFw+9G
98T/9QMOBXrvf8+2WTo3TSdCwo1aDy6o318J7r2pj1CPHfmLqbPKbQUfwSgenlm1
pNb4x7Pi8TOY4QFyxTKlJLg0TyQrTPjrkEnd67gO0fFJHaltoUUPENbK1qY5mZMw
6hIBTj/I1KNkgcXpONM02Bs2gwaQxRoLki0qPfTPyG8J4jQSsqKPdCYWcvaFl0Q+
5BwN2M0WgUCdXHmDNLTfzT7LoEvVAvyMWECUXQ5xaU/e0r+5clmD8aY5ArZr8vZj
PH1hgoeOC9SeP5Nliy0/srQMespKAfQXdPrdyNX3g4QLJe9y87g8Mtao3pvBEqcI
q5mlpeIrKUrfGrw3nbC419qggOslTrWDcle8Us9w1IKEg/lls01z6W9uESIHCgE/
M6U1l5WLS1cf0xxwRZC4mjKgSeg3RdpoMi8rg7npFNKe/3V9lCvbKmlGCqQxNn1Y
/BwQzQZW6uDhLEFc+JAaHp/JQQlnzdasRlTD+UGvflMSmNgePvQJABbdbxFwjk3i
902rU4aK1FxANCHw3T2Hb4ZrYG3pDqFjM2Wysi3XFXaANMznu7z/GSUwr0gbMkyp
Spv2gKA3fMQhwLJh1/+tK/Y6uNhFqbpCrFSdZO1/vDEfNoMOc/zl1T/BrppCopP/
OQ2lXN+yMvl/rkhqJZvjLb5W3bLcyMos58vUzFenletxITZ6FWvHNdezhBTms2jc
YPviHyFwM0n7n5iQYzhxq5ue1FT4j3rzEYDRaGG1JQF3Q90aozzLbta1jBX7rPkk
cxqDxi4P2BRNpQBC4ILVpC1pGYMjmMDGvZkCLv9DfSJqxYce1nYQDIws0xqflruZ
tLIzYiUuqIQAuMLpu4Am6/naMatM6WO4rI1adNYEi9b60fpBAVZd/FGL5TvVIcwE
gp/ZuYVIgkYk+W2pggpopunmr0saaO/xkIogjsk943GvghQl7Qk1hXqECqXaQ9vH
ltJFvxMVZ3w3cAB1c16U5B71U33OdJYnDHjMOClJGRGIE9IxjzbN0ZmJD+ZZ1P1j
MycR16WtOShkKTcMLWo0PT30NVDN1ZNMarkUMtmWq1X73xXkcurONZIPxxYfoHaP
57trrwecAokPstJ2CDDYInvtFdyf2DLO9RF1cRmKTsfHLOg0V4ci1AA3m0Qxga0N
HuFNa5d5Nu+pP5oqyfKfaMe/HUjmoqsr4Upgv8ewflK26JPltQ6Ra60zgCkoxGRx
K4phwPX1TAS2aER22sKUImliH7J44iRAiLhoIm964PBodd5OFwU6EhuaRjEEvZz/
fWZrk86KGyOklGg5NesrWKYggt2DSHvxmccHha9RsRMWbxDWNUvLcbzn5R2T2drP
xne635/ixqekROKQ+gbIp3cyw/lurKRA/yTjt77JdeQbZ932+AmnRh4qwcJ3SFVS
jCpZeRd9OBaXaxE1iiUswiP4oMyYtLwlyr62sg70iWIbKEn9VleIi+yPB8+02MyW
JRJ6KLZlkyQgct2q0chpph5w5IJU3CU8cyj+Ud96FhWR/FEghRmX13j5Ovju7kIy
bkUEO+DfHzMkk8CjDw7uubCS5DR6UsG+XMFZcDRmKGXX9McuoqmvENFlJAVfDc89
rrC5DT9hYTmkfvC8C5jRUJ6gcFMoJ8rd12AofpZNVlu6HftkoAa19mNRiM/VJxDc
BF2SaeFmxFYO8y8dS9Da6bRLHGYG0HG3ROc63pd7ePuiEvhynNWFB2LTCfapqNDd
HPfvyj+IkwStRZAESLb+Obe5Ws4u3fnHG7NKS2hXzHOCOAooFO6fWdPts8FcS4Tx
ulzmBw1hoNU8Vb7b54TUMnTcNZuwTSdrnPR+YHcbAo1k+MawlbgpMFIczEoLyGqU
xmWZ0hUs0zMb3QhnQOKrhMbW1I83buRhyZkchvo/JiOi2DxKQNZWOwUh87bjHERt
sgr9Y3Hdv5bFRyEWjw/stQY1WzzqLhIhaw+8YZv4T/oy4zqNiMduBFdTjLW1Psjd
wVThtfIJIiFG+SGbfx19sqnrqEDztRIzt75/TwMdaylRPVyQ4wkcypSIXggfU+v9
vZ5HtPDCTjNJqShJyBaG+u/yaVuZqHTgG7ov5femU29JtHFbHbrSmG0vMMLvLm05
9E4FZLeANc0ucdOnggaewhzGReqy52B/W3mGLJ/y5HgnJxrSxeELbgJd36u/bu4B
hU2PKJUxphR3m1jrL1K3647uCfN+C6u1/Ew9XnTwPCJ0JyqKOTlGWRlaA5eNxT5S
7jFiZUAsa0H7LWEar3da7gld0VyZbllQ25sedLhRmBQ7Dzzcfy9fZICuufUuNs2o
ZkrYr2tzKjAbVdjLid6d54DYUi4wHgx4TRNj89zXgxSeYjCCL7jEs5c+wYdqNVAu
rwKuP16b2Lh1d++XjQEZkW3osFuuV2tMRM/yHVWIatu265Oc0Wkg5hPGlA3yZjRR
Pn2BnL/iRizrAUvp3XnUfzOPUsoUi45qKoSUi99gt+FJazMBgCGS4BbY0lSkxOO0
FFOmAj/TBH0kV7TFmMj/ri/VQhOL3Uqjov5jPA9DCN+TFgvq3iVAD+aB89Pu2I1N
1ls9QO4uLMGBhYtsEjxKNi20Z5Zm6WrnMlE8NGvBo7dlAMRdLiFmaKWcQUZzZBKD
u5ZryCy8ScxMm0AN4RLeatVnBVrJ0pkn0YqAUmXHYpsTWQ+pahYr6xAr1xx5YLxG
WAtayAMB+dbDexn7WughFiOvMjnhv7Pw2n555J1m6H9wZrioxbIZFzkzhvTcdkh8
vfaMYWMckgVbpGM0PEjIfr59JiiHBs5QDSWylNfoA6a+UiwY5TcdZFf0v5a/GYdz
yG7JBKehBWMmouJpL4mvxpQz6AX+yAKSN9E9RjdG/IfgndwvR7V1NG6mgR1LQOXe
hITlgYBd4qdF9I7/+jAQq5xWTG6fP/tcnGADE5TMrSm5+/mPdRZJSfxT7DN9FWlo
3BV4Zn8gNG2wLLy4JO9o9iWVKpU3ihDevyWoXR8S54FEP5tHlbX9pOG9GzNhjDT8
nDweJ/7uBVZf7bx7fJDv9V7s+hwHZ4IIkO+2xdhxjvPUMm99caDRT8d18JdxOzP3
hcmvWzgIENksHJH6BMh5h/t/0iD/rYMs4JQSLDOXIVCnW7TKH5tBIxrN9EisapKt
Tib/NNl4siHFS52iVemTmYwjh/gZPhxvrovdkxDDqjASznJCzMgBalQjs/P208no
k4BlY1JIgH7yboU0qtxnNo0ukLD4fWDXZqfQDG/4i8n+q5onc8dMShK/4KFkvi9n
9QJlqIrEV7fstCXi1NeAhpY9t/m1d5V4XfiFnitNSaFEleP2ybQ+tDWToKoXm/Jr
Fo7lNNltsrd6oWc+mKALWkfyexpDZTRjXpUjFiUX+2ruv4wWyj0xLoaAJN4KBr7x
GGXahcObInu4J7xZvQgvG+pk7ICnCB7cU1e1JPT9WTO5oME3iYtL9JF2ykeWEwXT
GmPPyfEeiK2XAOW+8Y1EW7Jske1s5sjy87nxd3on3mublZrIIbq0IRH5hzJVbp4d
71A6hNpFRbWlLExRCwvxmEAXDsaeGxU4/Yh6qm77J/K5Zzep4ZF8XN0AcDraWqBZ
TyZ/GUys/6+km8jC7OthAVg+/ZM+qvRDZE+yHw1Ru1/2bGM1Yc4LS5mYyZXuLcWa
um/5/UvMC7RtwktSh5GEV3Xi7IHEwuaZM2Zmhnts8A/Wf23oyWxYXkLpA/HfknPI
1zl046qnjOBjkPPdgXjNDYV5DQDG3perYDgTTuLI+BgWubN2yF3lN9aruninwJAN
XyYfNx+1i9krrOuL07wLZXLtlkMNtOhsDc88xVWKeuWVrcq+bT8d3OLgvjOIqAZ2
+QemzCQpXglSfkmipg357+lc6/65RddXnXiVCbMv2ojyzgq8zwi0M0IYZGph+ooM
y6MM9GoHS8SOiJUdm20jun/GDpzzCyW4xuFjeN2d3uM7hsB41lR8AylAiVRrYVVs
NffmZVEMmSWXpZ6+VfW2yFxP/fv/Q/1WT2MdOm6OjhbibC3mWllRdlUmcnudOcze
c3HEkaw7TQCov/jBIyPi3rmNbvBjvwJlXnIASQ3HxScnG4DU+X3JrPFOr1uStsEk
b9iAwU0vN8/bjFQRs6nZthp8CUJXgzn8PrYq9wZsL4aIMj7RIEs6ltGDO9JfA7H+
vQCrINX2ovEZLI0UkiY881lUOeJE8OL5sVFl8hpbi8ar3tDXBaOiH7M/WNm75A7f
ZOLJI5oQvckkpWHrjdSv0WLdl8kbcxoGTMjzhLLu77J/vuxAdCC3ru7d8laaheKw
6jcHti5stDXJASiRjQlloV22ONjsLiy1qmH3VyJR/jf85CsJsZaLBQN/8I16e3fa
TrpvHeoLGHPofJa9D1bQBEzYHKKYJxow+Q9TXdiGFsM2cn08wIIfvZvljOzjvKeF
BmJH9HHm7DPi/H2uNJkoZz5ARSZO8FP0pUmxqkT0qTiFNaz4ZXo5f2n/64HpG9C/
QS5PccSclduxkLTsmH3DPvk1GBqHQ0rvcdPm6ij9Pll0N42GZ86W5fhPkTIfUb/m
bL9pJYYx7lvCWKeotIg1pqTzhhthpjmzhV6B/t+FXTGLSZjSqvGwXxA7xdHivTjD
khxhOgP+dDyvkZqjGhFtRHPUw+HbSrLEKO6KC4tRfMTSsQgA1kkjghplsGxrZV7L
OJe+TUxA17XShQ0HguNxPUd/PNjC1yHRT6YwTUS8x6PX+4zGEvRTnmwEs/CD+WxY
gXOVUl+7CukXzz7nXKKY/caNKHrnUl+pzmzjFRJlUBXM8k62z1VRB7NDzE/KIjpH
PJx/9jhFgKoDRBaXJRzess4glo9DWffWepv83hf+gUbV86VlkLoaDuaRny+gMyey
HJB4+gH83RV53L5fhhrkAxRX+2ZFyc/uz4PZBVZhfQrXapXDNYBIViOnNl71nFRV
lm9zpYLL+NzVAEIjnRkLTfDOV63O7eMQY/K3ai0GMMUHxPF75cIW1aP/FAE3ccw9
vaJpGUfZA2bjji6lSM7e1ardJeO3+iI4b5L6xSismxKYwRd8owm8uwLQkUXVjKiL
JiUiHggRepSxebcZ4o4Q5egV7iAU3M0sp7dM52SpGHoR3NBfAxFxObuYp2H9KFJh
ZS7vEBNRzHsLmBz9BnXwcGJ868tMN3KtPbFof/q18P+YNXMA8Tj60gbtuXh0wAPK
cG81k67SG62s7L6Uk0vMzARTwkc4/k8NSgoU+6gQLgp7+iyLQ7Na74PJB9FaLYJy
vikGmeqVGhcdvGCpk2lss+CdH4dR/PwtRlp7ibMFYtbgO+DvVJtcbGR7GEGA2ZOd
vmV9hrwMca7lzlUG/NyrebRk1cj+a3iCaX5g/BQGEHcxpr4zu7V+J8Xf4PaabCdv
APvzSV2END3PH93uAJOaOZIk88/1bgbhuzX/Qe+JMTs49Y8cBdAMemBzFVfx164z
aQqQyFt2dVDbVkh5nKLgk4TeKGRBg0Hs5FZ310TL8C3UxagLXS7sut1do99AYq1o
waVW3qMzRESAPuYP/xpR3GyWdEQHY3tiMyYjIJ1cHzc+S+zaqSp/1AYYEyypLyC9
HTHOyqk1N2JMIjaGc7dxgdN3kT1ZmUqBZBePByXs6eTWs4IaUo3VKytw1ABOko9e
SILidgj9eVL1DPLc/umQZLlfBmODU2xZYbu7/H161Ndoj4vds+FyBS78btfOIZCb
Flr+2lZKlUBAIULnIEP/SClwxfpgPEv1JdRtjYjH6C9WFTg1MX6GEt+AVomOOwpo
LD914x8asONgrVhDDNal6GFn4UOhRx9Lmi337SmExZRqwufEJiZaw+mPOBuYhIGQ
OroxWU7MAMAwq1ENBIwMGZQakrPLFSQv0qvHXP08czgj53DHsWNqyZCE3y7XYN/u
TP/U+51I10obe14YdCHRynnEnm762iv0+jsAtexCABnUR+sgsMNw9s4T0kzmalBs
vvhh7260S2CdkqeuRuGIIDFLrR5L5e2pW4v6yZOljq7niRlDjYST06GSu2v9bgLF
6Vpzysijw04S2mNZ+OzcJdgWLG+ha0Xidgv9z/366N1NMB4mdIwivWvOLzgOhVaS
7jFELeTmaJp8CRyPPL8Nkv3tni7doBjkDXLSCq+FaKO6+BX+LbBb9h0TaTxrkaVA
Y/W1vm0nhKM7ENpW4hBSwdB4nLeC3zvz2EQM8tHdmUuGsVxMp6xJt/UyegvY8B09
HP1EFsLxNsUqB0zDk4rY3bKbtRg2g106eI+JQ20kYmFfzpPJ/pJyoFwJphuj5Mwt
olE40UvVef30zUNz0H5PXprWaQScqYO2hEsJEbaEDwB3y6MBFQWwTTQZf60abrMs
aItK50g0EcrQfqYkTNF/M+22VPvnBeSUVIPcYsEyAbGVSxq3raASvb0ZUyo2uFm0
dexfkKpAf8UUgDuzVVjw3C9Ky/K2hsmAgyCUAZqJe6UruZvk7HvRRXRck5uA0YR6
MHVFxmimklEqGW31e+SMYpdZpJEdK6ZbmEtwxdxD/O3uVDrbKA0wn8BmW7TzrciQ
0Z7tFBBDAtGllY4wReO7rx2daRTu6lbfP3hEoIUxY8n5ttFl4v0f4lan6kIzFusO
WTBNoHM+1idCrhKH6vmMCokXb5JvXylOiSm5SUFWJ90Hqmcz5MqlRFgOXYBFAYP4
Diwj8BRtgv7a3q6txPUlyY4J+1/mC6wc+my0hLCWLJk2P1nJKe9SrmToy67O6tYO
JRbkYvL8EguDmeen99HYh8OmodMpiBdeXvsQahooX0+Ln0wXPH2wRqUQ2O8ZqYyY
4e54/q1ILtqwSOH7sI6Y/VAhMbBBY6ScUKQ3IOjCIxmOc96B23teL4iToQFiqtie
NPzIiIN/UHuah1Rc9VI0ctwZsH2tbVCH3kBHPvmeBCfsNXDfrkQI9E8gX0V5TS37
ddhmI+7F1z1g47ybBHvZwbILoofpvg8AHzvslef0oVpTA0lOVQYxeSNc/nj7tOzo
a1Ji7HqDM89/v918lAaETkNuIBMjqXSsGMQr8nMnX3f5IgD1ZWRAVtbmHuGQZBBE
AmCZP/90t8Iws9fw5Pou5LTTtS+aOHVh/8jWoIbU/4Oi/8ZU/rF1V8OWvKGtnYRO
MSfI6nzbHHjU8Kz+wBw5kKxV+iEvhL7D13eVJRsTF+lKBUX0UF0AAkRF4MPCKRa9
kwr3gPIo3z3a3sHXtsnJysoZ6bh1ln3L4ypwp+tlF2sv5EFZvFkBidWJYyvr6chD
tAZhJZPRAokJ9xRAizIwP3CfNFZGVYUjGuG0ZeWrpQVeD3SbXDeNPRitdhqZsrsK
IfskQ7oft9UgKr/1u3bWHRyJ0JrZ8FUfQnYBtSNiBmLWfIrqaPwHtxCvVk2GvlMk
nhEzxzJlUIhhQldscYj5ZnIN3WWzRRZzNClmCtQ6DYaw+0iU3N9UCt/FqO+2JrXG
Ik553CrJBLWjgiQ9ZjozDQyRVfV3t99J7gNacyCOKjdATIK/0NnQJeVmh1u2yH/3
dzVb/Nzl9nIULGi5cammeqlhNGTVM2VZ8PUxWIFdTiJpaZY19wfzotlNJJcpxIR/
z7TQ4O6XDMwZgGBUPbAMHaOH/VK2VQfOC+yMJzZUj4fA0wgl0vj7KDgloVorJ16m
zUdHWgVnaZ/WwR9u6NKaI3oxsEalc47VZ6H8rTUw0MC+BEPLwjvVlcuHKHYDV/ll
fHgel1G2bhmG4xUmmWFqv/O3Ot5x0Z77OnRuERVmd9jL3pzx9X/lF0fUxyxYuWzl
48A4Z7Q4vicvf86ykTlBlcBHTQqZr18U9+GwzBzOw3nodAiJYuROInwNqrjqJLMd
DjHC2krAw7ppAppyvtCYL3OVwLEnJw5WBSoQ/K5NIzqTQLdYgtckWHoeNuOaAWSs
EurLHDvGvcmuts3U3uYpkQuowWdtS3HJKnhsS25ojbwgKJVL4NtXJA9m6a5D6Pi5
jcONjivdmAcMWE6ZA8aR9u+wd7c3JPvuC3rgXAhq3S8/CW5Qh2yWwei/1JLJr4lm
7CT9EJcrConBi4IPF4LcWA8+7gHckjpah+PSVC9jMUIKR7xYAAKupw+o7Tn1/6CH
gl2YtpslHwVY1P14dA5nGCmkMIjc28k0FjBxJDex5H9E4Cb2J9jghL5mbEbV8JEu
VkU81AZeJzSiq/JPDWJS+295fRcAMNZRhNtdmEKESyaC3qyFtYwN8nz1NHsb2stw
6aYssMiD3pdsQXmJ4SirFShBEH+rmRGQXGf/IjQBCWWQcn9EFF4A9OqAthZBD62n
QRNBiWg1E+Z3ZpmsuqzhVSMMytk0qZSME/U7r52ikk+C1qqsqYcQtRW09pCYtDHA
1XKcukhlVD+uw6EhZtv7lxMbP7Nc+AJQuKLw416UD+lu8fjlFy4EhuckFULaBkM4
8o6x5uJpOBiKDJFbbYb5Rmt13eqJtfe7lrrQ+QwIJuLNZ/7UfuZB+HcICQsW8lS2
8hZI9Hn8KQs6qAwaEZencmreN0EoY5XRm8RNkTG7zPvm2sVCG0BN2lHzdFV5V8xD
UtPfATXrCANDXSiQ/7q0CW8fdxqzPMCtczLeFzRIZghZRKSy2rJn0FTDR3oFHk+/
OsZ5/FiZ7eBjOgP7MDgF00ckysWlESGX6ALksbBPksGOEvfpxB6K99DrqOeYFY5T
JeT91s4F+eTAcDUvYaAVrieByD+Fjdg5O4sBRL2Jdld65lHl3qjqlApZjXvmUp20
ims2pbVk4kGW9k2MgdInPhyLKx6ZjOAE1c8RDD2p1lbvvp1VuitqIYAzLwE75RP6
JFR+zQYSS3t6pQ9riuKBamA8j2Zslgd1AW+30sRsOhTCu0IdQgOHv6tNRLI4fZWz
bYB6zQuhyCH9XKzOyfOJ+azFiXVh5t+4ZSSo9PUZFvQ5lePKfudTQDEf4B4Z7jld
b+3ogqxbHGSrGWMkNoPGDowbCahSepmCQqFQOEaIb02mqF50S78GFrBnWCLSPEl1
EvHvnLnNTRLAQ/wqJ2kzTiG56KNapOFMgutKsaVQPyUpdf3jjwVoTnMzAplPV18Q
8U0waabzm2zFupXq+qf4cKsq4kdg+j5pWc5zGHXALpZupDGeFkdopMlRsSl9zPc/
SwQT0Yi3YRlMfb/ot9aaZWKTKPHHxC+PzZRo1xl1hb7wp2cU3kbKxdA3wxnqqWv7
Q/tcCoaKWP34iXRJxlwL6r4XKs10qwB/t8WkWqBwkWSrdW/43K2IxrpFvigVEf5e
2zNXta966gILNDgHUKoegb3AegpbFsQEwAFnsZt4y9eDy8RyrZM8UBLQmwL+1+3o
b13t2i5BaDXezTdMkjz0rHgbbyV3VHoj1Hp9lmFDDy0zUHBIlAEl389TpzVQMwuR
R+If82s6AuqPDpL1SQUcowZqqx+u5bZE+FgDrfB9mZvJ5ektRm8qIgeJbIt9wItG
07YyBrLJQg+AwYcsbEQIrm2ziCX5hQRtrveo67YFCKpEerO1OTOKpYxIvxGlvJ9J
2tGFJF8jTmPuMl0sWVWHtJ4fAnL9E2BX0Trdlo3kykMJkGRqOVYbW/MFBeFq9Zb5
7yveei5dLCCLsRseBNwmxcMUWIxqjbYk6R++eD4gqdRwAeuAioAU79jmQCwJVAYv
U6jx3F/cyuN0MDZiisYUv6iOt2M/Xl3YJL1x6btXm+yjRyor1jyD6pp5VMKiqKQJ
54CG2Y90PSzy67cu1DGnprd8HOzcnH91ukSKkVaeblYUJ6vqxLE55yN1DeyOA2OQ
qmdCKAVk8nbWaZCHNgFEXwQYnbsLWWkLFWSDqXqKUUlGqoQpFbJlNtn/T2VfLWcr
r+H6uQb7Hk7TE96rL/lvCq7vODFBpjjCrpSh9m9Jkol/M5Cfha5XtZzZqP+DYgp2
gzqT8tBLKvQko8d8WoO9QQ43E382jr9dRRedGIc5rPbdXsUuGXqJlfi3bs9MahwT
FiUIvvzdtcoMCp7ItAqhBS2TDrvMWQs0Ct82AU4RxiwYTUEPmpILHU0kJ7Jfl4YS
SBrZGcgt1drSWtTWY6UPW3fOT2FnKwmqPzM1Ui45ZTTCoLL4lWrGqTCVDP5/yTvs
6Mic77W/T7AUSVRyq3teRPxTpSD74RMh8VaZjBTBxR5voi+GI1+u9uV8yKAmigCx
/ulvsFUoXKsGLdHfoFhcIE3oMnzgngP7YpwOyUZ/LonBCU0rfkabfKQPoc1uL0t2
WlkG7hqzqPUBEy+fhEUxNt5U+/U8zbpd9HMd8IrBI5dusCqE1oVxM6yMSB0uzXXO
H9rZmGsxrP1hhiyqqfsdlfi9JKIQfpBf+CyMawY+RdS9NssWrk2n7jPnkGc/r1Hk
a4uqhytJLgxjGoxkLb0gCPC9IvE8Q5dyX+9V1cQKtbe/laNuTFeP5UdbzhdPEmDT
ZfTKJCh2b5RmqLtWWxZVTUVo/MelcKKVL+unnTfTdjaK8s/Y7fl0EvRj4yOJtd1p
Kl1BHZvJ5OfYkpxRigckFBHKoccfcl8Mah+YTm1k9wTy2rwH/cQJOhd3r0EbRLCU
qYBcibTRat1zn1ZsOFR2zmgeIiSbc68nOmrcFnMcXOXsO7WHg9I/igRTEDVxQz/o
Y9cOJ58bHOcn4ZecSb0YGFQDZLxq7jLeOjLO7zKUBrdcxt9tULHqDYuVi+A4i3Kn
j0t7xIM3LrfSscuu5Har2JbcjzxhUzQAvEJ1LTLZt57qYNq4AbUJxixm0MoabkPw
97j1GZ8k0lMtYkwrzlOZCHehv4SWCx2TPiePb89bnVEC1rVAyjp7px/ZUYeSsad6
7CXCYufTPKra6o0k20dEK6zScBczueuvhPV44x89A95rw46Y87/J+Cu2mrWYbSEL
rMLjnwA00kh0lAed9cRqkwTuw0T2oZBMP/3xsvjiTdXtO1Uyvu3xAwXPlXhbocPq
fp1bdDI72q56VFVJcoWB08voWBaYIwLMVt+XZO99jiAyWyomGj43avzmJbfimmDt
IoamC13ZTyF1QWHruOhRypqEV8rpesRdpNUa3PslznZ96D/q4o3haLt080cIQ3sw
eFNtj54foQ335lb6wvg8FwwgBgYxXbkDjHJVb6wJnTCmFOtrMuaiFFUc34XY/HF6
ybgEKl4heWpKOji4+WRspnq+T3+/xYAQc6f34nv9BHyitDuj4JZ+gUiyaeM8/sLx
tbm8gu9FpkD2hiV2oMuENvWEa6V9EOIKGNBnxmCjh97WR2Hg3KlUr/9/aWziuXje
AbqI2zr4gwyageNsCm8RPwEq0TnwkfA/amZAxyulyUOhWqgNM5tXGTPhrOvK5lmb
a5ey9BDr1H/5M2o5E0vQLuYRtFGGxyWGXd19caaB6HJokxkD2gqIHAu2+uq+z48x
HrDOyZfB/CFle7/Xj9MUafmkI/1J2uRnkrLZmdftrd0IfuIojEi+cWq1X+ywJGrQ
lL45dgewKLCG001qTtMTJKgzp4KZqqf56qo0oYx0d+cw/GKnthLkIYKYUEDJfdJv
uICOo30eFWTYiYelgxw+CGqxLoduPMABUbM2KncQsZGjNPOelJqt+RmEljQNgJgS
ZPTs5UgG4xpxRf/nfkIL1dPB2R5p+fdoLxksYme9vsGOphr97QbTj+0834qyQY4i
qMnqVVd5fXZvyFdktBOPRU+eRkAlK7PN77TJxoXN466MWdlMmEdkqQs6+95t7vSx
I88msnLI38AWOHSxiL1oRtCi0VMTrbBjaO5Q3iEaEY8HhRjQukXQntaw7aQ6TWTu
K+qkh/RcDV9RsknjwqPqykdlMuZnAdNi9L8kbwTDQJAoq/2ekogPVVGCIT5PvUgS
2S9Kz3NYBjgJ1Nahg7X6PzfVK6nj6zDia4HiLkOhGInOR4GbkbX2A0hOy9wQlSPE
xBIQbqwvE/emtujyI8Ow2AqQKPp7dio0DZ5eXM9U4rIVLNjL91eMJn86ACvwwUpo
lMxYicfrWwZxr+mHQ+cfdaJhQtQXAS0Dcwr8yYtvMNYavNkX87sbMx/XVHBCWuet
0Hz7ipErdrwL5qGZM5yRDa5ejNJ362pk5xkXcSY9N2IpP1vwvOaGWjYhINJbbKtA
6FCgmLJGLhYIVfcI/hKiFRdMMJOdP5CtX4lgMUNs3V7PO98rB/d7NTUymP01WxTo
mHZWhflnIn950dDW1eTUsOL0Z6DX9xhJRTwRbE6bIUMFA5ka8awpSj2XZ+cV5XHm
o7M61l/srovuguV8mZlwNKCKcigCW/Lmy6K7EzM6+8dCXp3C/mMTyBB5xJIAcile
uPU2FcHXGzOGVgYB5GgwOLP9uf4mjRt/d3yLHpSQH3geo2gsnUa1QhEe/TDQht/G
zJyv5G71pn/C6Y1Ng/8tO0tkDOKbxmZ1YigrwqRH6PaapLNlLvoiBjG5vhPPOH9s
orWcPoafYT35GfhzopSmWl0WCcVzC9jTkMXk7yzxwFeQuJd6y9x4hBv0xQO8sKnU
VjHb1kcqAJWGsaAQ4EE4dhdIBHzIWXx7arMAPsRmxBkgd/b5Vcg8Opx4VoDWaFu/
uh9g3RJxf1NPNtMxpg4KWS8E+MmUe/Ppe0vzK0Y0FAjGqhSwgMr8MOM+74JI1d2r
LC7zkY5bRiJCV59U7NGGJxfAADtGg4+Bu3bdZDG8itoFtaA7Se/UQN9nNhqgvSMu
87nm4aw85n7+Wv7a5kqOSkAL6TKd2WNVrdcVdB+JFj9VZYLui7Tr0LrAQo6cdKzK
Gjr1kxonDDqikyVckRwXxqdWC7GrjoBXU6DyC8TMIX+j+2h3EFM7d89jpTTLJX1a
v8A2/Mex3Lkeai7lKi++A+bU59rB39qszKNJKFm5mLxdIg2f2k8Oek+H+2bjWUsh
eKT8kz4kcZLQjKI52Phra1nVoSNZ1R2OTvMdtQ1qEzjKMcGxVGpYPZi7E1oJJ7TH
cDmDnRrDrMMJw32O9+pUrh83Td4CQs2ZtCbHPFPzwW/7cKfZS5BeFORFNucpQnYG
54OaYPsA6doT4+TjC6pa6sUdUQE7Rq71mEP8oexD1u04678lGtwMEWHBxeAKSdwd
JnQLUrANtfducw14e+4kf/42/29ldIoHsOha22GzDPXhNooqZHdUvATcTW+TwqxX
YPHOYH2HXzpZbiwQd69PYeP/odgcgMLiNN51Jk2G9A1aJ6F8UWJCUIXjRvaJhGut
Px7/0g5CtCGi1fOdJVi/VqZCTlaJ1XxWbexz3GinNscDopI4lOPkAe6jTRgfLVnL
L9l2N1SLgXMGFrGBBF1D0HcZOcAvOa5MXELdM5/jifyNhO2/UoegW9PCNCx8eXoC
r0rm7zwFT9r6XIZufLEXEggOb0pMIG1eY95h8yaZoj+raLsE+psWqOlCscCaYTH9
Rm7m3TyCzmh9tI8jtMfOKqvUXzNuKinkrC472qhVez+Y4AB6tFIRDXf0wZHV36pc
scZ76TyBmxxWkKniVpTfYFsINg+QQ8mtQGMGQhXhKFtCA/6qXUHMCqxCD5la7ACm
1nKOFPD/Qzt3xBIIcyUYIopxZqdaEUZlfO2LTYDlCjxf9MX6kPd+sSbIHtlez8/C
LFlnmL6F6P657sBBna5JzirNLsgazZsKbbNBMMYbNXNA6EXH/HYi3XNsA/NvC731
voC3M01IcVolJ9YoOgD3PFCseP8UcqCs/FlpBzubiFxPcMEo/eQ4aPjGEbABuNlk
pdVbaxNVXGHU8xlq/fgwQ0JV/oOeMm3ZGLKdT/JpMkQrVRdhORFt1Gufpcdki6hC
1zwFm3b3wpS7LMgP1z09tQt90W9pG0KcP08iPB7t2OAHwB2n9Z2BzlCmUOtiT3UN
5lGO83ZwMlFC2r5xoLVBbxtKMDO7vl7I28osyduPN8T5F3N6FxCHY2+/uRDXzyls
DRsR3uM7ufQXUSTzlSI3fcNPtPToyOE/Mkh0P5tvkf62huAOr48m6JgCCMsIplNc
EQm8Yh99mYC/GvqfHY26Z8vcJ1ddL7k1TO1XGlxQPKhXmHNmHKSzTr3Uxyf7bpai
abrsjPMK2AIosfe2E06u+CMkLHHni7ANAlG89Ov0m7V87P9PVtj13y4rrh5xPPV4
0XPI1cTuMebCxHalT1YvnLblhjKgZHz9QC4xNcN64zGIfA2XVHNuThKBsceSRCDj
MEHKLOteDSTyfPherRGtAhEVXuTKJTx4NCRtumM5NZz7uqLmOlBXjATL4AF/4Xg8
GMIsPOeRfdP852/JhlBOsnOl5iZRUNdcgPi0g4E/gtAlw7fJ+pxMeiS1bJdt6+9I
co4Jna7XFjQFQ2LuFsOFaNWZUaGAT8cUvdTjK+YkdZZiw1A/MF4G99+gi5MnizBj
nwbd84+PQbEunUtxZanJ8sBwKWHog2R93bfc8ALMUOr6CCUQIyf2MveHhNLdVVJ0
z0yWp+pAoaiMenankX0gZ31QlYxjJc09BeXeerKcMtyrSDqEbmYAZXibcYiWx8IS
vcrt9bVNdSZo6xNzDF3QQgyYCXV0AODIICNVhBYycRDVyC5b/L/VzmL3RjEA7O7i
qo9p0Yc/DAHyypyWTf7EAfbc9T+fvbTY0221yu9lukUAy5jzzhSD8s5UNKIhMLnr
a+d+lk8Y708mIYpyk/j7Bjj+eYh+1nZm+H7N1q34Rpz3ER/qVWublwLKmUUffgR6
WGFzau2vCZ3VXaJcLuSOLJPKjQEZQipoCqPI7nq6zJK0isloNBndNgEQ2t6/vkEz
XCqx2hah58i5BGdaiSfFlnc40kYqGslinTaZe+4YHm7oIkIG7FgUTbwpCJwlNJzQ
xH1TgYipoGede1hibgizBvmfRSnEDFn1Q7th+SPclTCo1lGnfs5BmIHke2qD+Khx
hDUIbt/pEeeI56mR7aieVopH4/sfF+cYsbu0EoCEHmVpqwjUhAzcvvozdMbBSIkv
1OsY97zdSq0OdSnZVP2cVm5g1W1q1TYDNueChW654TJnX0BvE5QY42eF+EnoSIpA
wojRxHnl32YzpIw+YiReH0rGAhxoWdbFERp+cmND42WrTGru3hJTU7inarc8gmQW
mw9ZVg6LABrH0yEVUALBY2H4SatiX5GIZafVlxHCbgXMO6GF08sK6CQUWbODy3n2
GKFXBK0qVoN4dLkDcgT5WsNEGbK/+6UVv8OOH+JbkoI7xhL23A0L3fzLtdp/xeU+
cFxrq4gJ88AqSErx3KQeZRAH18ThWmHX/vhweIHF+W6sLnGD8dip7yESzG5JqrXB
HAUP5c1ShKn2F3Yhqed4+Zw85/77k72ybTvmHADjMhIo3brM1FwBiKRI/XNTx1IE
9TgospU5iT4mVa7NGgt8QAlZsmiJhw49Grm/JbRoXhPEL2Ug8ost+0pqiscLGnlp
BF4Utry/EuhjRTGJr1NKWNJQKkbjKPLE4DYclsybeYvRB4K8JGIZz/X7c1V195Yi
e23qMzZ8Z9MsZsM06s1crYDh/HMBFsVlRurXXipQuwbWbmx9MQ2s7JPd2PwBrXXs
w1Vt2JHY285nkBMjBgiLI5GAGyMaJZuiSQPQI4PR0G8p/yVG02q1pNKSFgx5BRq+
G7h+FWFNWjMtKc19W3cYmbliJ5O+5ATR70wIClC0de0n9z1eL4yQ4absDAfMxgBG
a3EmPBDwkaQoS9DcGI8ens+Ul3LjJPLbGa98EF/ydZ7ZDMiZZ8/AV0zwzqOCvjJh
rl/tZbT/YDY9BeDE+AIPDK/+8lcr3NgQs7aNFLnvo7RfBgJNBetEEhz9GiuMzasE
c0mqvU36tS8wOw6tDL6ZkKbmJaakkrO4C0wygD7M0bgOEd5OlYkvONNtn5uVR/H5
4HExghbjgCPvqwZQJ/kyE9gMwN2rexZus7dmJ4jnCkoMvrNNV+A3WGoX2JKGR/MP
lrbq0/qNXdGJ7M+T4qR6LwHqOKFG7cefZlFU4S3JTNBDbe4Lsv1drdlZuSV8MGMQ
QxwiPhWgxtuguXajHS3Z1xtysPQhoAAiebyl6RTcN+CzUZn+f4KqafVQrTgdVaWt
c+44CfIKD+G5NL3fQPhI2WIoM0sUbaawSV5x/QtuiFOqEP3/ARsRZY0mc7dcTtGF
hMVRB1YbcphcizXaMm8BVgUaO88Tq4OKKKNI/hDk7AW10W1Pn9KEMlJSZlVZ6e0s
KqeX0TzKtgxzqjcG6gHn+wQLd72tk5ugI+WTRVq0WP/xxp4YjCsrBUbTDS1UVbd2
ZQ1qa3jb6T/m6LNjEr6Y0jLjMPjd+mxwL9QCzq4jKNCCtTDXqi7ISRPVHi0h2kJh
XvBgjJNd+yNq5DquCBsIrDtloZ9/MOqk56543l9CHrhzEe96C4AOcuKtlp5ox27X
gvFJmDnJaPssOfDay0yRCEOkeEZ+JHe7dqWVD7Bhxcxj6mgC1LCyhIqfCtaoy4he
lKVuGtycBhDGxmfVE5kDT/voa7iYrKzkzNrZQxKomSB/UjDr3nvzTNZ1TJ4vAgMx
vS6W2T/pnQ+SkYlW4rk2HikA2Jck3xIrxS5px/ILrf3lpyNMA1ixT5qtb5zZofD8
a3gm5R9p0gZNF4VtmFflgveHnidV1mROvegPYI4YIREL8WpdqvPnSxTqU0JyBZjx
aC0JiVF7s5hRbpxJGLRX7tP5Gv9+04b/ocXIz01p0Z6YQuzO/4rWhcRd120aFKdN
1ovdnCkJ5I3nVQCvbzSUkrJjskvpHhpTlUtltnCdfrRzCQjvtFnBouwyLgY/mEZ6
mVnx1ZTo1miwTEMwj+dm99loZWeNM/Ygj7qEhweP+IiQBYe+kx3A2nnrTPC+P78p
u/0Hrm5fNRQQd7zy9lUDJsdGdOQTN/Q0D4PN82TJpm+mI41FOV43S818aD5ShPkE
BknoCK+p55w0oKw5JG95K/JlYx0ED9w5oKOLcgvF9EUiGBlJ+BwN8woej+rfSTUv
jJiHOaXgz3tbjc3Q83wjEJE3NZfOnUUocRoeXahiNigLYmPXfbRSSHJlYgXCugoQ
hHjRGaXX26tRaPWYwEpMRFyu1Q02zKETHNVa/H8hpxCaB3yafok7IfvK+/WnNur9
vTk+7Ajc5/Wh9gE5EhY0AsMXAAsDTk4qidqpJlU5rpBQZv12NUO4bRir0Ze0r546
uy5FLX62L0H7/B3sF1Gsps5qrIbnR1qEgaC77AYE0UjZTUdrb+9Mcw/EAz/NoG4X
cmd0ltFDy+0HFMkuyw4rXHDdZOLq8GXaQYZkPnDxyOMRh8HZx954VxptXFJV4CJ9
MV2oNuu1dUOOZO/XZkt2qhvUGGeIK2676MPDlWRwWpsIV18b2jaaxEY2YdtovRLl
6c85CDUnuD4R3llrUDMjeu290YqRI894WdQwdeQFsKEAXqvzUIBrKYfBAF4NEP9Y
j86OWYbUjzYE/jO6dCx/51DoqnE2nedpY9iStQEoaeDwIgrMm/Z4MIDCLPOh+upF
wk162tUhcANvjmkG8uwVOPrY7O5idKfWJo0RmHn4bRsGg0a4uRNJjWWTXuUK2JAc
l3xlO2ssx/vzrDIyCVDkcaruuekJE5kS9lGStasHsDEKNTu8bllbmTZsxX+uHTuu
rWD3HqywsJYLVTWlmSrZR1p9/wS1NhwA2pWlRLs9C/cpyMDtyuSopwurD5bcG6zL
PxpzuBeCWdb23RAu5v0gn/EDg4hLE1T/1gBWxhbYq12TgO9W2x2vIcuMua2vRpVH
LT9DG6teD4+Gl3S7kmJvVm1y5EAMy79JxmqFpdMnG8CSAPUbitVLuFKMi+FK33Dq
RmEF85lIjldiiwhtkJLACYY1Tah/jwkqkuU20bIvSJyExABQqaysyr/hyIjjl7tK
vOY++pZmy9JWFn7+87ZcsLJ6/WiczCyWgsFkxWSc5CsGgYsk77j7HMUNoEOIwvLd
HyO2hdAu0zOe7GyaHyDH6fjDtIBeNakdIn+ou7zIceWjfWZgJPefFG3XQZKFw3hR
TeNWPoJJz172JvIt2x6eSA9eoXhzN0sDu/dnlMvArPlv2m5VjvdPcoIt4yHxa9FD
Hj0ZTLxocEMwWEc8bODsCdNmMiiOjbQGnrqosL5inedjUSpzctzQ1jz7IEsCmd1e
ZC1Be7dQf5+mMfxgX7fvn1ky1+ixYn2HKv4txyH8P+JLAEQDRzlbdTwOFEnagQP0
IsDomy7uSiqWj/gumcIT8BRa4Bemtez0kmLr2KdaniuyIts7yhFp9FRr+wiv5FVp
EnOkpB2LPKDrTyAclCm6+ot/5+OvFP3Zbt1hWgKTpoWs5ju9UhNgdSLJZ4PWs/B6
HS93oPxoIIcPecOIazYo1QB0v+ZeKhyXnYoOaA+nh2n1f/SV7/RJzTsICIqEztfL
O5f68K2fyROsMrW44EOCnGEl9Bc8cZHd+ikbk97oy+nHVb3846rJvbd6MpX18KY/
hsi5HEF1c3mE1zzT5AWSElwTyBysVt2afD+JcNRjJSpoSLpK0d66SadRpYHimqPN
SCFqIMVE7lJaT2fOkDjDqRjf2lARjc2+FaF3g6VWM9f0lglFYKsJZ18KH0qe2TmY
Oy8/hxUdPcAquCr5vUL9X4VHTRX9a7p2YMkYO6m66bBlmKRtnFQ3x0qOpkHQpIsj
S5Ju+4kMuktNb1o0uddksxEgsPmByi4Yd7jctp5xUDqG0JzIOgIOoiylGpEIQc6X
Re02O3yvbNNQqrpaKAT0WSrljZRN2IScp4SzPwGV8QfTR+VvguW92f5kppG3K48R
soMsBZrB4heDi8MB2+qeQCcEScZlsyT6RcPONmy1H45TJzZ5ffoOQ8GxCUF9+NjK
GdFGxv1L10S8fh6xytnMCRQJcaUUWIF4Gj/NnWDD2/tZi1/x/UJ6aCUIEbnDlAXD
lqX1fcOlTHdPcOBH8niC5f/J2Wbgs6BLEK/AFqMYkWUA2hmcn4vV79eoCCqcvCJA
MMRZLmTSqguhyOEFl38pIvOVbZ5djwGDAb84rAbR5PE0IAWC3NtnRKE72Di46u9E
ffX5yAY3zplD9f5OiwYIrU1Vf24RKG7THkWEfHZQRC9GqPikb8z4MAEawztQ1Meq
DM6uF5zVRVs3yfIfhlOfkJ+HCl7xQTgpSkDbJ+MCvMaPD8DK3qYDIQEOAqq3Tgmg
f6VRkaZietGuhrhs20WmT+X1LSjX4BB6Qgwgp96VjSMdTG4ux9eAqYMnLW+Hr9Ba
lDC/ETzhw/HAvt7ql9t66mxwaGW5sicj7aPL9yR2jVnl/L7e8vedFQoP/5aZyBc5
nswWqrmwVlJW0/195kQ8HRusQhO2P382EZXb3jSyOfexw+yIqLKSEF9+2dRV/LiC
2XsLc+V3BED+OBnhWmhz/P71sUjYvpBrq1K1q5DZI7TyqPuQK9ADTVZVAWfZ9iZ4
++Rold6wD6TGaFSZpQvYjobUQqS3Hc5H8bcP7MaMc9TfIB8kscSarfYTBuB6d6k0
PGumLtUiZ4pMJChPNEovpffK2Zc3uqcHnlm+7jLR/WFdjo/dQzzBJgReuDc4Zr4b
U5BcEBFDG33vzaf1TgC3VbXkYmgR6SCDY9X+Wo4wucVgUofR1pWBdvKmjAePRtBi
OU0LuOBEzuP7r+EzlGfGKj+kryy2/hUKQVtW93CW74Z65NZrA83WlLV9yxWqhXE3
WuK8gDMfS+VebnBCyZQ9LH97mdXxj8cENemEdloYkJeBMS2IdWxLjuBHIQp0rZex
On5Z9N1L/XO/KCBb4zv1uDVnsVYS2EG665Y7KftrqkZY/ND4RuN1M1Ru4TPAJF7+
Yu3IkOoi1iih9sDYA0U2u/LHz/v7iuj8/cyvHZma4TLPV29uq33iGJ0IA2LbcftY
BYH2IGLDfyfhiqQeNOrXvrmgZb4fS93p2n7FChf7pXetz/ftLjsklhL/2A5HMVXk
AMCKFv/KErwayKSb4y6r18Y+lf/SQ8YmJeAZ1/3dBtlXWH7/5RfM1t2tTn0sNzcS
WovFYO64mkn3TuXQgShHawlj9huO4j/Gi5LVtuiGmgUdzTQfSaTH28My6k7nIpdX
cLVK9zZ1AfCG39w/zbzQFNDWMjbf0UUgqwhFdoceyVGSnnJARr6TNcCG53fC+kua
TUeQDBhLVAbfbQsbDl4wDZJB6POa0a1IhcqWMCfwfV/oW8iDzvSjot3twQybE6Zv
GxhTQMUWP15RGaJ3ly0wCG1hullQNzENhKOeveyGDtWYrOhgCra44hjr+u7gAiPT
cIi6EegVw6k4ORPI25CGRel1qQi79BuphgVUOoby16hJycyzlfixPecflKOY0/Nl
We6o9Q7HPmoK4nmynd2cXcusflyqIsb2XcUWeFKWFpqA+Yd4yTj9v7uAD9C+iytH
iZDeICHMujTP0BDNy7uBzlLZ2a7R0/IKws+pIYqY5XWak+AxNWjgvpNmCzGRoUCy
Eur2H8H6WKVeHjLcp1TkvcKfLA2v7nyH2yk9wskrzvxrvfHa4jKQcw9WkI0U+lIN
fNDcrIdeWdzaObxN02uQAHCUUFzs1cejSMhIMxKp8I4PcmNsPtNKi3Rizj83lt57
jVcefdqK9jXUbqy/LceWnbOkhtHBAMZvsh8PhoVNxtq5wCAMCw2cSf3yT0bVy/6u
sMRZKVDKTUMwsihIqNTU88ri305sdKXjsmN3nbiZ2pb5cNLTU2tBa/pdNhEvIkgp
X+RllET/fn5RxVK5bb/dx4RXCaWg4XNQB4Zt9jlRN1V3sKnopStxw5Vx9eZtiiWm
jWD8PruTDnWggvGubJkLP1vHvLh91kP/LI0x2CBKnxFWoomPqjdTKfjviJCVradC
PdZdwHklFjL5QWqu70EyDn00befX8Isgbu8+R4Oo9nhmquwx62qtiQHClF+Jymv4
udfcw1TQJCdIO/ztM3XyUUJaftCmS2zPwSSEsx3wObp7mVU2IsW+zSiXBSgpgNen
eK+szXaSKOZstPbPy+OYTiZmV567VkId8WUSMRnhySqynmHiZIUfbHh3wR9NhpxO
cYOt7gbFzxf5sivNmLr8cyEcCndcdGYkBYTS+HE33w60ZPrISIBTag3JpYytm2zE
jOj2U9K5+HHZ18hVBgWtmqWlhsHoenks2Mt/+ZLR/+5Bq3Ej17KJ0SjDUbKykazr
BGfA4bfShvws4Bw6l5FjfcUC8MFFljjL0KZ2pIOn0Amwy1eFYM0HVQtQKgpp2YsZ
Tori2M4kPLDrYRANEagLyMhEjI8G5Uz677aiW2sTvQuq2XUuhPbwmV7ZOq7mznMH
WtfjdKCsdL32ankvpeGyV8jSDDiZrHQHMVCcd07UuaXXOOnmfwNbF4RkfxPfsbFj
HiJ/1NNid5+WjRf9iHv69DVsQGdhpTLE1KAqH49VE95yQMBOluJ9kChObXjY/V3k
2qzZPAssZZn0o9C/TCU5xJsJ5GoyTR/thNWJr8/iqi4A/X65QrmTgRR+cVBdLkMq
x1flmp6KPSAowMFqPrbMbN71wDG2nwTYWzw5AOJl3mkmE2n7ite3O5MS8nPsgMRa
kyWYfKMYQzQ/HWwFBJA8cvs2fog2hs2NdsERjSbVARt77krf+FhhsWgT6e19MlEn
YOs3H1nVBG/g9hseZw2RrFBw1FTjBfANOnot1G2ccJifRyzZs1k8k2HK88uOaDzB
MJOjS9Di0UJHHe0s/UPnSqvmN7ZmIZvRHHeG2eFJvKA1Xj0JegHe+9x1uswNxWyM
nBknNkrTrY5f+Gb9B1+oBgwkuQNLdx1TJYeCg8kuPjiyuw0PPJI0OXxCR+D8HOBE
XPWYZ1okL19HFZgydlL8Djg0geYcGj8fSdwOu4v5HRWh08teLR77A2UAVH2ab2KF
qIqGT+uBj6/S98SjZbYWZURcIr3ro7TfCQNxm7lL2+t3fzQkDLxL5cDcflilOPyc
7rjMrvLcfxPzscSDeE4GEAXiJ8Lp5GA4BjKUj8ITDSOBp9BGs1vji+7yCOyNx793
vSZzOoFPjC5yWhIpuCihSLRpSwSWJlhbVjBYClKj1CqdqiY04G7oS2rKV60YiD7u
BmZAdd9I0ikrUtZcbsMQHnBg1NFloKUPHLgBwyQgMCGv+hYikKmaru2EB1mKksQf
wmEioVMh50RkITZxulGSahT1JcbFcVQLUq7EkTG96NLP42Ca6H5KNciiPabKyCvU
DXzASK5f+v6MavlBLQ9swXU6ZrSB1rPvacZIdI4hYwkTCbVdY0U7RQAcCEFaDFRY
XhROtgObdu7Sv/s47K3P3AQHIS2tmC+OZV0LEmPdCupF52C3bbK+kXxNP3QvWhnj
lgRnQA/92ICRjue+tR9M9UU5gY5x6s6IcA4V1U1wzS+SLqUV8pUyca15aF7gPs7P
aZ9QiXRJR+eZvXf42Ru8lpXpLTH9GjeeKGlO3ggD9vhs4whr1o022gRwxKmMxg4d
z4RFApYbBafSUmPJr8iOGGlpBoDN5O2URHc5RKlTgIERnI+NAA3SRJpNr08Lbxry
lsn416wfuvv0gt10mREneM2nBqe68fQL7P2kDMB/2UeLXgwa5OuQU7PBqjbY1HT0
g+IPqWJkp7vaWfT/f1tnkqCDuZtBbew54luuWCP5cUl/L88cGHpCyFRXMHvqlmzn
yWHSVhcaWhNjNYnJ66wN6jp+VjcTGV+L7k7IJefTl3f3eIOwFOrgqlxoS8iYEq0Y
CdqiXLFSw8pjStOtCBl/X+5msJ2VgDC+IG+NCttinm2qulTjPlLXQVoie8ROfHoo
aMDhp4V9qT31sO3IQZz3vt2Lnwa/MKtYoSjjSZT9Bv6Y6GHXcx1oaVmKQplOSXro
SGGCgJHuqPbNHrj9DFZZdsAt1yToYFbcxNu8wk8YFazoW+1+DKUkR6Bu2M9Pf4oa
DKIcnrcZkuRmRH9xoSfdpNV4POvT0BBzrYDLcQwMFFWLYxGx8180zY873mE7pfa7
uMwyVD2MHbPw9E3ge4ZqF4UfVQMCjMMS/rKWaPBdHAS1GB5q8cw8Vdo0/lmA5vVd
C5b65/fMdUaf6aC9hZWwXWmuH4SgSv4z92ghpo4/hCyH9WWe7jbML/meZAgsM1DP
C2lmsE3d7ybE3iVpMT0T3nk/GFL1b81loftfodAR2pg6arByL/qUGbB5I7JQTojY
YDbQj06OTMGJd2+2Y8B14Kc6C1PEUX0ZmJ/3l3WUwhJtEpH/9dwE93Lefl7U2YA+
kt17CaB1A6MLpGmZhKFfKTHc5BQ1obV1NAO144zRtJ5WMx1jRWCZaEsATYGq+59t
7+TkviTP5CVT+1lzs46VGOSM+uFQzYUvQRcUfE17E315azULoYkrllwrCfeVCxsG
kdiR0NOVjApT9y0gfQ5NTjaj3WHlRSqEOEvynOMh60qMsEbE0i3o7sFK+hBCGaIi
jJ+/rMjlbwzHS9OyxoUd2K40rICib2H2Lm8lfIDlcP1T1NFHmg/folArJ2Zrd/wG
yIrxLe5qHCVuO3jKwU1dibGji0XhVbdgv/KNadsE8PkAlQC295y1/XSGsJ1rECrK
N2YyICaw6eYu1N+BJEq/Ik09BFirxbSdq32s4FyD69pFcneEkfJotreMqC9ovRni
7kYGCn3aAILSjQcOwMkNl2UeLGVjGlmEdgoCjUaOC5Cf4CVuVM3QRCMVC00RPXzC
kGlxscZVTJUENWqDUcnIR1PGvf8Rr8d6rloEZH4vXLPFQTdtNyIOb2AKFHndlRKG
ecEHO7jg5353NJKLUTGCaWjXosEKupZeTwaujVrUaHhK+SKWElD/NaNqBQuNrLpt
uZEet80uN2WaBob1piLMpEL9uGdogOgf5l8x7onvNAARINp4LavRj3/ZB+GEu3hk
2RUPcA+YzoxLpa3dX8ofANCkww3PB34WpcjQzFSt5ymmB8j/QXFHVLbiZrM1J8g5
oJF2SoSmHBCaL+qURxiRCSMxHfb/xwlq4l7JwVs+MaV8dVYHkm8LFg6YvK6eirFP
/2V/hdufmsKylF4UDC5j17kEw4+/KWb5MbfItI0nU5G+URDsf9JRB2PsY05w+/PU
r/AV/yA9QnzWEqq9NZPWMvMkKLvgdQXaF8Yp9C01B+4JPFkdA+7Z5/W+DPe7uXZu
5cqCLrafIw5CY9SuN6IKTOCE2R799gFy15zik1Rq4tt3WCDSENubZwmeMhZIqktD
1LidqWCQ+axq2sTp4FospblRwdL/jbLiTd0m2tBbZI/B6vB7vkw3rORAGQJZagBK
M6WQFqcYV0hrmy/Zwf+TQxM8KbTuarD6zLh+O8DGn8zpMl/gvyiqgEm5ezqO783G
O23IrtROrW3dMQ5IPcdY1mynYDIIMR/SAo41hrTe5+meGyPitJXGystOTzvdL1PD
IqIeOZvQK0USAb79V+iPewfPM8x/90FtYMdjrQOWpu+vizxFWOKVLaBG9KM5qRYR
AmxxPSo38uOCAEji7OI1o5swmydf1NgL4/GuuCuu+GTU4F0uIUjKF7bW/tHlsAT4
TUifgxy7jaUnv4jPTDyuufro33qD5AA9mnTT+mqg/PYFYyHsgRi4kSxGFiGkVWHV
9ZjuzLs3G56Vg9OWK4MfAy6uENnlU7NUdPBzPTQimOBYaaaLHV1YIB4CtXbgs/Ci
epqGxZbs2ECKNyGLK/3hq6XqZYS1Tjek4JoncnbeJOlXk6yz+nla2XShsaKdRMTe
YreCnTr9QbaNWqwr9o6JDfDenfbx6iHUcjfpdclX0JHg6vuMizKb/UHe02YRLIHy
eydcFnZpxAOW4981chpwKbLs2WhtsmPpOKsQbklbzluPuC4UvwoWEWvTGRGHO2h0
ZQnRlWNvQMkMM1XFwL9wQA4BvvmAOyEIaRWUhOTlOspAoBnH1UlS4iz6uTIAfVxr
g42ewiIQZywea/ODoKFng+/8Nr15//ib1OhqVLooyHMyLrk4TcTe2LL8V3C7vFWl
8CyjH/WJ76Gg758xsFA9gaOJP+yIXV683givwsbKR8bj5NEQtoy9RqiJTgvfG1HE
qhTshrVJ6Z1SJlQQEoMya1UV1isiJvCfLeq5ZmVu6IRWtbGbNZG4TAU+TVUKvlFi
MYNQL5hYd/uVYsQ8EYsK4dgPX2bRA8S+VUABo2373Zzwf8XCwUOqD/VETNOfA8A3
5W31sm8BQ2h+pr6OiH64bh+A1A5buAekOxx2ljD2/y7ygPuKSPgsXMGXUlE9R7TP
+/CEJ6qtSeROtrJ2tBalN4W+KkGMomLeMW/G7ZGjX7JFwgiZK/WOTejKGeAk8e2N
GnbnNkvbkUPfiwZHQniFSQXELHvwiFclyhvhrangpmdC0wLZVQEKNK7wSjnz/mu0
2DF5PviLlOBgFDTOsyfbw1AMKuzT8bq7COsROfEgVlClqPrNw5oMRtQUVo6Z4Ifk
gt2HSh893Gap7LKcIu5yFMVZl01ap2TqGazNNnxD9VNjvThThHnbuH1Ws/sEEc5B
ucjMFVj31tU1g/kPtLTPa0v2r2FA+r8pkj+/OBHv4/2T3ayzf2e41UapH45Jajb3
i3ywsF7TmoqzXVYF7djVyUEG6XaRbo6qBEUPuapkaSZTaZ2huXQaZZ5cKYvKLKyI
IyC/ZWURD/v0IyhDAkAfbw2SAziiTzOt5xRxqjwqHTZgkukNsqXyvjFJsVja74Al
uP0nnIM9GwDMJPCm0Us/QwqDe7x6Wqpvw5eoLRHDC4oRY2UVCnVZyEYYQI9YRsi5
9sytaX0WRmXB/K4a0Sn+/nTagd8hMslovImM4/2addJIC42Uu2LRz44R7741j24P
wEgCnVYlNj7/PGNHAqmr6Gl4okhnhNaFOCeL2NZ49BOk+TaUhmdEoJ28unheMNgi
TfKyoIKWaRA7lRpwdGTN3ERNHujEKW1RY5/vP447vvsej1eWhvwyu0V76GkbXOba
LWWQZEwv87TLH+gxzLgLy2OZ1C0vX9uFpsK4S2bwVqOxRzBwJp64vlDmMUfPgFHw
7Lbt6RZW7wAeYhzWQj3zC1XsMeftgPhTY1GVOm+ALtbGaEkMMTvPx4Cj2DNNVHf9
fkqb/TNG2gzrCeUERpkgxgocGnB5dp5jn0ire9jNd30ua5WsmnHlCrkYjT8miOcP
GnUPnV3NbX8fKlDfkND9k4rTru7HizeF8SpzNX2gBCiZPttCusUPm/aJ9Uw9eshQ
GJF8KsJfqOeSjEhYL2BfA2++d6ikpAArQnndHZ3XuMy1FraQvIZAHCvfQ6M7B2sv
SjU0hqJg82AdXR+sYoCprTR7uo2/5Iq1DjSnB+qBYIZ8F86t/KbTZq7J3uJjyFIh
leM8a4lycW8wE5HEcDyR8rsesSVk7T/yV028o7zO4A7lPFi10vnW/yAwheeNtQr1
soiS2F8xjIbAg2sAfjgVq/9AkZlnFEWXrhv4pvL6M1dBUW0T+lYkXrBgyh/0MlH3
xke3iQlDHeNk1kTe95B5G2tsRT03mOlrldnlj6dCAZeMiRfmGKA+L36aYERIhDKj
Br/dtzXONf4FzI3FR1admNb8yui3bOVVi0wyY58FpGSl4F9iwCdRH1rOKrzwNmKB
Sex7hWW9BqVRO0LU2bdz6gWxxPVkz7P9pxwYiHlB4+hEexrBQQRUbtPfldxWfm2d
9ldoqngmkULHad+kYwLOMGCnTh13WBBHeYUmogZZLYUPUw/G4JIFcX7XmztUpzFv
22Gs/Nrg5J3/jXQIsfZ7UIWNNgvqZqVa8wr97GgB4e7kH+RQ+7bUUCYqjvIJN7Xp
wEkP/z12tpx1CvcB8OV10ToWWdXeYMBm04MvlTEfbqW6N/oYgDZThQuWk588NyKg
Zws+0TXLshLsozTuLB2LWOGMOAAyXFX4F4YzYNAQ/RLrUWhtkSniIh+5UXA/+CNQ
iAzpKZLjl/D6g2SpORUxgoky2aN4iNyTJLA2ABeB46hAwhxNsaLSN/Hz/Hs+fyK/
BfVcW2rv9roJipIiMVmpYmBfkEy9wgiqb5bSl/hJjwrrru3ahUuAkeCpRsASKeBM
XsuxYzPjP1CouOBrPSKDJoOpe8UgR2r1rlV5j1nwMmU3bAjKA5mapYz5mUzXmax9
wz7vjKckbVmvhGnKFiRK9PBlkvopOS6mJE6hQgOWYsFWMjkj+A76SRIyPko1e44A
MUnOjGqv4gMbxRtMh4NpgBe1pupVsBm92pGCFkKYebgHeTKnOfwiSNuRfNSAFGTx
VPO8ryhKW1Iw891midUS3qTRoFA8hyZ8VShyPFUmJIirXxUUx5tnoeB6Y5eqyjNV
rDx6RA4cUXwH/V3klr4022xLbY7rCeKVhDgDug2kSCjvBe6C2crpl28/JqV/ufIC
uVUpXdHzDcAVeu22H1q0Nwh4/U3LGGGhmC9rQeeQ1FA1RHjSRGUR4/lmQHuN/RY5
ndEXMoVDbRdmdsr4YtQF+pXAESOAt0kpH7UeN+d7qjJndtr4MLuM9zGSBNUG2BBE
rzWe/+QZn2V95jWvbdkzgKpvLD/y5Wo4tQeMSFy/lm8FD7OxjXWKsXHZ6PrEfpZJ
SM/l4e5K6NXeZuqivFpbEgR2GsCy9Hy8zpewnQif2tRSFSvp2NVF/Q/Lm5e5tXjE
SGLAp3lowIWLzmMzAMNae3RtxWCLpUFO42CZ6/gevxXlkFXPtDeLe/NsKy6l2tdE
QfE1qU/vc/Zo+i3QFwxovTzm+w4HZsozRhGLOyJazsLWgxiSMcck+gHg6Aqhwiio
u4FR6CEsgeabG/mUOjxN2K1BszssgNEMulG6BAIf4+0i0+Gbioiw/Z+7AIMv7WXJ
P7eVWIsrRCFq+ZiQNZCI38YEIj/Jv+50QRztBxsJ3IZK+QSnKEqcocTfTKpTHwUl
iMlyzI0upepEwjahtAKEDloeuRyio89IEQ6RO9rUd7uN/+0HMuOXjVfAFzNflXfJ
PrBowsjsVcPNZxT8m2/oWyA/zXPPlqTlmmtmXKMpn3Wwml3RDf51krFDThNAafjj
k0bm+AjAHZIrkJAGaBQms+/HM5VeOnLw1PKFEUoi7wx9A1+pMdKHGqntDDUFtDYN
uVL+LaUm3668FZfseTQW8kOH1B9QINQxBn4ngsLk+T12pbmxugN257+DmKdUwCoU
jXTvbBFDBraIRx2rLeHOxx/alfzoue0SZ4gGgEN15l8jXJ6ebiPppx75+Waznsq3
BxEeff4DEmK9UK2NgS5K7/up5VtQ3PaIzEjpOmkTDoPDDh82A5DoXjXfkLFGQIru
44l7zesmvIS/MVNVfp61Zlqb9USj3YcPf2k0MhRukO9ai03xS1t/1m0N1IdBzPZc
IgQmO5War0VVj1az4AYW4vFsnmoy/TRKTeNA/ffpBXmpu9tYQbShHc1KfqkB32r4
lf2QAA6QblFIpfalcC0HUp0peCoYMuf5+UZgJwwECcvtrmzxz4PKT0c54EhQzgk1
CPRdCeatxfISa0nv+MYB6zAgGDwwYa3oyW0jqITd4FLS5W34ShUhysJWDiMpkEk+
QiLyHH7ovG+DBuYgpWlAPXb7tzfy/VZJhTBFYCPDgR6e3obA+XxEeStTwMwNOhHC
cM+aRUL8eHLRzmFwIIU2KxU1C2EihGK3H+diLHziDfXjG1VWjc5YH4ZYEsD+UHO9
ck21rQcWGoNZoRXI69X8LDVnjOD99CHdhpGuimgQYebcmpwO9SAF9k6ibTjcE/HQ
Lm5LNvGqRMQVZwHN6fleNRBZFGNI343dB39vqzWwwhbNMo5TjyB3IsmvRfKNKZHI
lDODD1aSjx4m3Wtm2zXoqYt7PWZAzIvG6qooxziv4pPtC7ypGOQp8Zg5prz3T1Vt
4D1w2R4tKkr+mt229Rjlf5FIx0ngnkkClvOiv8yuF/qe1Cz448SmYjVu7ZU4QtmV
wAC8HYrZrT/amzstmqDm6cNGGUeivHwV/N/l8ogBXGPXdhnHKaEUVc9+YjKLTM7d
ENEVN9VWWN6U368LBsLIAw3Q0ijmLsBvzTWlWn7BJCJZX0XonCyMNysuR8WynF03
vEuMJY9yKRkvCwsdgJDFyyC8EJ5EfCHb85AwLqPV4tr6Exnn4hCEgt9gQul8sY83
ZQmYCSN96XhhU9J69BuRUBusHxPNr2T3ZpgJhYEXG9mK0TNEMfYHkM1w7OdBFYUu
dA5RI+3FxVtmd0pbxkRURD0CGfKG1o+EaZgTLnLK27DpLT1Q8/xp7SYaYbmqVW+p
zcANiuToYH0ppzc5SnhxM+f7Mr0F73gBFDTwdt2ZYTPbkZr5/qbXyhwbWeaGUI0T
KI7ZFz9bZzcEU4Ne7CSAEw1wZkx7rNsSh8jKQluHppNpmdeKAu2Um6N3zaYIAEtW
RpchTT1a6TQnZXkCutTdO7DGksOt6Jl02k/x/DhfyvWLWBQZ233octWVbyeschHw
BUEb4BLVYU1UhL9IJmcVM4J5luUbPHwxZJpvSdmQ+WTPEksnTh+MDhrITQfpARI1
I2Y/OFy/jtyTKVpwb74gMRs8C3elO8k4Qb69RuvrE6ohYD2anJ+FaPuogKtR01pe
IizTkIDVOuBiaX9sgROrTgXABftNj5m0YmMKc3mdqB3FfcG+lizQ7MphrFQSdy21
wUVwAG4wGRBFR1YLR5U8bLuT+HFjxdCpdUYpdEVRmzR75t5G4Kjg01OgOsYuPrUR
YKpOMH32Z/EtjZZDnO+00i1baN378MB2dDXk1G5/0e6KUA4M7Q0pOkiigAV52hqi
emHeE4CvRK6LTxsfiokqOJozi/L7VlrVXrau+WfC8ajGPKYiya/yH92yGWH5n08k
ibMsIR3dXdEHQkfINA229ybliDUhyEwP635SxZpAvZ1kqyBL1rsY/mmY0PIu8WYu
tJ9TYQfLdu3eK0PgEi2DUHzHuDiNUgXo/7VwHVuujFJToO4cgIpjYqTxhl1YyJHa
ixq3twjGYHjg+W10kBCViDWapLoQpMKTgOc/exNiWKGSfJnREGOnOc8km1XZELNd
w2dncGbjYJ7VqX1psKY/eQ/s6rmef5gNbJoHd1fAHOmeCUYZ5ABDfYRxt/TUYwLn
jY1Yf0BV8xn4mgQpBPBNuo6fSFsWQ6m/aM3uzC7pUK9rbRGPsf5i/yzn7llblS8b
QsURdX71Vu16X0N1mX0gajtTRdug+HKtlZdQvhJDubzdiHyoSY2qyAjThItWfUKC
Y/6dXY4oasjdyvo9tO7GkaP1kdrcVKjYFM2TnyC824v1sIjFsx/YvEEaD6TvmFlS
Xt7HKzFmWHf5pUNK4+OKQoqCFGCbgpdq0yKIOmqyk9YUNxKnM+Dg10kmnNjBlrrL
UFD3uJ3N4ChwG7z9hz/exlbs5rkRxaSXWxgXt2AnDGlwRxEkhdIup6RDi618NaI9
3skkGwRaFMXOYBIsKWxGpbBDzRewACYkBotlwPzsvIBkUP1sjLSKIz0aoWSytBPI
tJ/3L6jeQT9Djr+AL5Cqc+O7kkZ4mSMi7Y79es3Ud5AyTOeSN44n1D6Pd7AZm6ej
vkVN39JmT9LDqRg77u5Z07l9vZ36lLmNkxbpehaxxYOkq68gErI+OlDZshlXiXFo
j/JHabFg1azu6CSMGGY+QNN9aN+ATtL8BP2Frio2C/f55cU5DrRTAKjEhN0wFcNT
QGr6VBwDkAw4M8IA3hEFpK4P8wUeJgdrndDh+AK4fj/l5d4XlGonA0pHH1EAsuU4
NqdSEUxF9Ahxvc74qo91VC3Ha4Go31DO1oyDX4dkUIDmerC9Y9ax/shS9exqaJRy
A6Y8x01FggeY+pAH2zv4pwo8jGCjm3zB2kv/AGlqTwgjeWSt4E9PaZQF4ulrD9Xd
VEgvUg92HrgEj4TITwnC+G1ZYWWqxJmMqc7IS9r6luRTV5Ak1tSH94i4DlDPhpEQ
Fq5JPOflzTzw8mZJBXTy07g9VGhs5RLEgjFvUFJ12yKXWhiJDgnsR3hA7CZoSHDP
+A/x/QzltpXXN5yYyoRMx00Fbg0I+6/JMoSKaR2wQlEjlabAgHjbAYhPC3kAzWIB
YS9iyyFxXzh7jKU75clS8wvJMogQG5hVLUQuKzNxuiZo2ZGK/88rBweHjf1FNAFh
DuGvutDJtwy2EU9Oegd/sMRgVgbg74HjGwqWYoDvZTwkYdA0JUGt/af4cWMZRatb
EEIkMiI+q6SufnZfPERAcjTQFCQOS1HnodO1n7204td84sxo/kBS9uD3Fcx//KnP
nOWyw5p9XWAVXxN4a0Maiav5RWycZO3N2jJ3vvEr9bDN0FlPeG88dEyRL+c3bfBL
bYYGROsIp2O+Vkx5v1FRvyzR41EuS8LjxQVBlMdo2TDRvEJF3SLdqDbGeBrMgW4n
bIZacu5wglsdExVVKo0XWKbPqoucqU11uwoi65wTZIFQARcgAkiQzgGLumQuXLS/
Vn8iIKm7+609duPn3oXJ8zyiGV9t1P/0kij7a6I1FpcQwF6SBH5mzVxereMTZ8dN
hVayhaDFia41yhqtkay8XJ1LmNpxt2gSodS15LS1628X2f2JFlBAFGjqZd36dC1W
zybWLf0GtK8LwW7QMd11VUdMdN5DHXSUu+T0Sj82nglQLyXJlPkHV3WXDkjsUpHS
SxmS70el3P3b4SAuQ9JAkoRoXlr9DJROEtt1YF6yO//IHcaCzIoxm9K3gKYCLz8k
ZS+Vh7YB7EMXHx/Bf7qQRVRb+OBcQdfoIeTmyFERAOl0Tha1JhMRil/dmLHgmWo4
BMURYjyIk3d/UbvU7oxjatJXLrLn0NuIlqxTbkLbGuyMve2VRvhKDV4XcDJkRJXU
xo/qXNyzoa5uW4LINGctTjsCjc7ndHbSJ5SCzq5lsXfp+HEWVDmEFdN4tE7gYk3i
sKwQlBY5ATCGi+88VAPovXPA9HPrTjWzjbdm4JGCUDUnixMxGZtTzyhMVlM/ppnd
FxXOc5LDsemFtNhFgoRRsi3mPx2jcnP5s+wWI4aN8Jwlal9RIcQzfS1JcQjWzJUi
YbiQr5pE9QLakMXG+JPUo39NEexbeQAKP1YqdtLA8HoFwq5SR9hXkTErr0K1Tr50
UnqbOPZHwxt0ebrTQFq9DyYlQ7iPG3e3Rw9BRcqlOVbX3KrfbJ/QfWb0Ygu8MgjF
g8GBpYBYQdT25KRc0jOpQnXSZtAf7PnXsv478viwd7bXyxPn88RRhzOR7C3iM5u0
wkY2NluFmi3qo+P1BiliwfwMr9FHHHDlvv0cOmiEHPDN4xSjARNLgj9iADwq/ucH
rGCUTNsoeEpVPuigVukyBr+MJtDTgyp3ijetxLGicBZpKvjrgPa0YaCaOIbqjU3i
d7tyO9rS/iSaEIQrE4bq7ORQP6wNc0/NHtwfeC53UTJ5dlw+oJocs+A8xJ2muAQ1
u4qxaB0o0xg0ljqsP8kiQNLcY4kjhmcLRS0zamDb2UWRPIMds4yo32EHdVaVR1AU
mNx2BCBC0iKbIWOvflaQkP71Pd8T9pkxQVQyopcSzgjrf5QItL1QeDehRO7nDkxB
S3SqWRe+0Y+jdeu+1ie1QM78wDcnhpi2mkyrcwdp32YfAQFi87rd0W1VgUmi062O
9V0vmlbryGXroiIB/uJGHtl55akX/WrynFEAs6hNg/D4Q3AtSfskocHXQ/UYs2Cb
GX0lwFhAttG9XuahpDCW6pIer9MWKOKBX3+9Eh2OlM8I32/QyicNJuh7n0iS6ZEP
ZwGM6+GS5eLMw+bFklAfWqHP+iJHxwg+6369j62KBNjpR6KwgNHljbYhKxr9cAfV
VcUxDRHA9HSAxjQd+WxEYobx1Pxfy+IlESpeTksqO71Wql19bK9aGgMFFhyKVLIX
JzWujkgXkvxUFROXwQoknGiVHGI1tiG8JmXsofc32dbvH9NH/RibXYzsySPfpt9C
UYF6Qila7X0yjh5WK5GgwUmb/ObJALKnxjX4HINfiyevxMKRu2I78KwMhesVV7pa
KOaXQpHytWlMZfFlVYbAPltPdGT8/EVgL+z/tZXfRNm+YdRJHFPwpenXd8QyuYWD
QH5JeVzAufSqL4MI0NqC7ryUWOBN8ip50XCSXOnLwJ1in5RG9b5P7YcASViCjh3n
IsPXLN1MMweRHy5fioCQzbZgn5E9247ffmS64qK1VRTe3BgHvXBOVVmgITLkGYxc
ZepOFvWIk9uiHXo+s8ZsO0x348GDjlxksDeUUusehLlvUs/HcuZY67lGxG6x3fez
7rScnAoTLVtMtZpv4xDeJCw9y8vmmlP5tfQvKnlwFEu2xcUjeu8/n6ij9jRYmxGF
rqfbXUx1iCx/o9vRC8hsSoO2OX7PA3TXmxxKlJLQxlD675RttqoeWvdd4XMbQPvi
LsSqfv1DDKbThF/LheOEAUEL17iDUH41jc6lLRVEhW914RSNBCFNJjCscfMwnQ6k
gKhdzoTbNxY+5uQABosiNwoUzFdwS7NjWSrWmivuatxe9FdIBt39ty7eBqRpe2pg
w+nG29zugfTfsqoZlb9qWBhVnolGqSfHQwaTwJdx9aXxnDEGA97e/We+8/w7HB+u
uGLj98CH/l1jh+Crw7YS5vWNXrSyCB1l5F8KzROWGUXH9+a4l4QToGBjOq2RczHS
YenAXXdRf3uRD1OFWDGSYNuJzbVbYqcNwaOkohFRBj0TCwxvbGwdMSK2ltHlfPg2
5lKA8cWNJziSeEgWlM81FAjgsy9b5+W2S3YkdqclHs+W/ykv+caG3w4fmKyvSR4+
8Jxr3V7gB7yYIUWO9nJm95EThYW9+863kDPVAtGHl9Oa4TzGC/0OOCuohRIcKXyM
rlcgGBTwn2IkX5fpWIh/Tg5+FcHBaXK8C/r60uWlPXgzvFr+YqwWwfYF89KoQnPb
b4V/CVmKJKK/5YTS5O5nK0zdGa698Nq8WPPfOu1cZYmIs9POroIrn1/v5rfg/a+Q
YlLKw6TrAj5iouUauxwycOy8mcMBAEH65BaSBbZLuVEmwU+pxvLhuTJFp9q5BeHQ
iXKAMnggiu1OSjIoYPhLfc4N6Oj59NKkB0dVHEwL9XYQvVcvxgQ3bJ8VchiD3Qnc
dIE50xjGDOCne+eI53VPHy87wdsIxF/TtvQusfCNGKZ0obGXgugTrL0374OYHPkU
ge2sRWM1xinNb+o4qi3TZmDiO3xU9Zt6K6Id0ISED0NJX6z6aioj8/Ka0BiF0n5N
cjlzZieMlF4EY1c4TLwB56ieDJsytd4VDYINsf05P5XXyDKrvPyoit90GePVeLsU
Mg2t/i/dFxiwN0xoYVrRDZLraO8C5Q8xcAkMMJnwrO3HqeWa1kDjVF/P+RffSyva
2J3MFEwTmH1k91Zr0KFx91O+HD095IzFNSJe82UizsCK3MYAJNz3HgiIqlYDyRiQ
9w6yVU0uNChjIdYtjQdKl68aA4+BRmZExVSkRGT5SjDZoI+5G7igCBVa9R11xxmm
C4iqTASA7Vj5taSoaKEQsUgQJIHehqOelSbwDRTQImSgLnlJgepS6MeDZoChEh2p
9DJ53O43X5YVQa9BOw/IA5sUOU+w7SkY0jPjC9atkRLh+gq102dSf9PaZg3hlscz
bFEtC62Og548eDMX9DxuMfz6tM5PR8wuOQvcKInkblD8vowoILwSxsgOFtUkqVwq
kUzRbvrumXWzUe0Dy8GNJColvJqsk4u+53ScC5zkQLm+gOKssEOTfpU6PdkROyGj
0Gz0jc8NjRQhso/v70KA/1Yl6FfCl8D/4Fu64xkmHnfd/RTIPGZzrap9wQD4fVlW
MlrG2In/0BmUGPwQ78LVkfSHns0X/dZJyHJLdBa04EnGvgGJbqe7S5Cyk3L6Zw2U
2JtjS11rltGYucfa2RlEGKc4YjH4HyINSe5AVGRxAru4qnm+wxohPvYC5pdvRgHy
j0pDu9yVc41JUzGhvZjUin2+NuuC/LSoiWErJz6nAnDsuTc089d024cdmAAdD8em
5SH1u0VwEj2NMTr8VBdc5KUpHoDwdbRb54zMyr4zedYJtRKw0jWe19Z5Ol4aJKlr
PBFDQYzEmTQO6V6DqZ6XtlC/upRsWf5okQ2dgrbGVP00ULoMfY25fsnFgtLp7cWx
u6LButQjHaG53ofDruf0hbF9XeDUEYbIwYNrSCXT3U8DCXB+1UwgRkrLOkMqcy0F
aJ/tefHESMUZRIcMpI51aPNEJyuP7XNwghTh5rEqn7ZPlnQfwADCLAMotej7dY2S
6dAcL8eW3wBXVOe9E14WjxIr4txuWZlU7azOtooh1WnEqNW8WL8q99kItXXicJqd
PFzNQ9Us5KRwsUvxbgAWCLrwd5tGmznBxzgsz663Gycq2uXIZ59xuYUG5fQmRJuH
/SKXO+zvS2x/PBIggeai9+SEmzc4VcBu3mDAq0DJ6+S86NkFuQFIj4IgbR8S/1E3
kK3jcH4E/kGAm9eY6sCydp8MoPj1UKb8hxZBbQ46G9rYcp5iv9Osf/vLMMnbfJ6f
uPMPM19KWiHlhyc/1k3batFDyGt3MNhWWuuy3rSPQ7AuOW1kyAHG+9bguPD/lPC1
pH4w11zDmZZBrXqyPVzkFisSjHTRCRf7gDLNSK8LEP86RLvBBAeZk+qliUoqtHqm
uetEe5x/+A2zRBidRXpiItftF7vzME0RX1OIWbE6pSzLhxW/eLedgWt7jZ+rNeLd
N8k06RH44w1bYMurSs/LOqRNAS5Khj/5sN7d/04UDgLZF7XjNV51xusFA49Ghv1W
61i60xqd8G0mOoOiPBDAAYWegX5J+epAXfpmEV9uxWoBWR7dY/cBZN1IHNNFAI/E
DBXtBB4Jy6QBjGn8nq8os2ejU6RTu1Shvqt4Se+xqU2P1HwuXoBiOFjgrH1KiNuB
iQgKhwCCfQ9/x9SoPzr0GeO46pHMHdjYJJN2dGv3kU1qcVl+wAHvq3dPTfDYTKdz
erhQDPdNgjlT1nn8C7y/ppnzfp1Ga40kMrAfTKIKgyVvdKrYm+ov6aaL2gZ1Vjvh
SVbsANwGpV1xtGNikYiPUS0HU45OCKsxchsP4CNTM0EltOchKoUWMycIa9C4hgtQ
U4JqL/EuoKneBI09b+IPOM0QD/EnUm59ZJfcjJrHSNZ6XrtKn7VqkTXqoZBoKOmI
qTpnSg/47dIbnf4DW3o8mA75No7SN2uQcUFT9dgPJLcfaP7bLQnmdgADH6ee4fNh
xCnc4puLlEHs7pBDwV+UZExX5a9zVWbe9pEdXQDNQwzIQVIYmQjRXYie+M4A6G2s
exStMXeriQXbKNqccpieas35d+Ocdjx9cp3r51PwQWt/yzyUrtlopYFm71sRfiPq
EZmrsZo6NcFymp0X/56Eex+gCnEWs8Jo3tikB3riv0HKwLpBPKr0M5Nul3dTh7x3
EbTcmWfTF5L/pc7ZbKAPFdvSKHl2hqxjPdcZusRzJp3SmJ9LuI56CZemSz2lKz71
8Lbx9vX0mMnUPCJcKty3eDdm1xud0rU+AkLjTKFwJEqtAwycUA/2v/mNWanIvelV
rqbvPfChfimrWakSH1Cqm5nwMrs7Yq26SKyrKjkQMmrW207JvJlKra8dk6/Hw5uo
7dmFYkPtUcSK/IAjnAQpgBtHIm+h6boDz1NDXNpmZIFwoU/30VU6Hfz06AXpUWTK
KX+be26qH94XQM2jPLn7DWj/9GaqnjKOSefoO5KTsGsXTY4DjbtUuwYI8UeZ0mcP
B28x9cQSzM6tD6S6zL4UQVhABzlGVtpjopLVowSkqQJeXUe4vUsrm8eptxDS6EqW
pU34kEyklzOZp169Ot6a/+jOkryieUME5y7B+fjsSFyHZIoTdLpnRyglO+rwDA5W
tWlLAwOjO6gB7SMnpFJNWzhatFFsi4YlTQPfVn02E/sI55MHVM5B76/a9iZE675a
Eqkcv3bLauDC764f+QNID1zPonM3pNmMFxvjg+Fd2+/1MPn859AvnLa3EoL7j/VP
ZDysJQ7lAE4sZKm/89glpPGWtJ5VFLTSf2Qko70aVLD++FvdbLJiUMtDIyviGnR6
6HDYa+BwcWj2PikzW3pjcFiPq3JHKUqLI+T1SRDf7DjwDgdiPv/1P9Y2BEogX1nh
uQuW+JhpL9qXkAD96piqQNe5sdvigAUjCmY5ZcK04HHsXwpvyjDadjiZSdCKsMg3
DAAKfOJ+MgtjQymvULzY4KHyZ/bNQT1W7oNFgg70y33MWSrl3wxCD6vuvHFARVB1
GjR1JObJ7aWvNWacjM0csEk8MbxwunMGgl9fk3R2A9OPz1FGOVrhY8TFDlSDufW7
ot5LovkKnQBcDFob0f8YRiKoW5eOGVnPnvqvFJgLwSFDCzu47tzsCbpl+syUugsh
6w3Io8GuFJ8U8yijrovMOBvF8xs2fUArR5RP3a6jkDlU2tiqZfb4KIy2zLRc6P0l
cX7DgK/mgYk/IVM/tv9+47/WjrLTjT7b82/Upw3/nj2aijx6rXet98OicF4zwmqS
OE6NJTOgbA2eWt65c/t7LF6XtxYCyfeOEH0DpWbzjU/2YQn6Nu+kU9dwr119F8tM
RP8r/7uAAtsEPe5/vtXsLBKrb88tbvsYlzCjsDYTDdkgAn54MGfjnJltnOeL9r3/
Ay0vaP6AO+P/bWVMMjbkOmhVgq2z44iEYqLaEBStF6izCHDvUdT4KMwjnPhNtRQT
tfgnUNQZysn/xBIQT2YXNMtDrKDxL+dPtHdH/C9Hj4ihoEZb76ABRi5usgV9xwth
qho3En42COyHbbLsXm48WAYbdp8trCl7H+PmUI1LsKyVXNAzv/4+P4yu4enOVZGv
0guU1rAp9a8nS8es84XZXDUh4pod2MVBo5HJ9a0tXRdA+nO0gL0MiF2AMc78F4xD
6fdAoCIBpJ4+VhTzIcQquefKV8XsOi4VBE4gGVIbBV/TFcertLJBKAhxPHGfOYwO
ci69NV+mi6c5bfR6UBu+FV+g+QvS6RxOX4qZDAKMzP4JepCLI/A3E5jrbP6+If5t
fhnBKRRGr8qfZoX07FQjGlH8nkc0e+eTY7yyOAodXdmvsvR3gbQNqxhVUcetxrQV
5zvj7V1I3eJC7bmmxgtQLL09tlhW+yK4zO7l1hnJNdUJKKYAZ4n4FqYdWG+kBPBX
TIitV4WQ0oLYU0eVg3lRVM1BfCzEBgBqzAz0PhoBTtpj+RL2iDX6ImVyKhNyMG/T
Pi8feVA22VHhJoA6aim3Gtvzu8cey0sB0wV29PEG0d50nYnAodBaG0kKHbVq8Jku
uXwWaG2jDWbYaZJ8haFzGJSrcKjy9YdJNm8NCxQty42LIzAxbAvevZy5tFj4BP0y
jHT7pGf1xq57EdZIgrjDaos1nnmoGjWtiOf1PpSQYerI8WPMx5eRzzo83phWddDQ
bWhuZL5xD/o+4+TRdT41y2FTODuIID9g4W9tA7Mf3wE/pTz0zEmXEyRxA9Lkgo/5
5oFbPaHIFNEz0YtF3abNwM95w+O2tSb6Lcda94lYGdcr9hFcgAuhY1xgynIpMQx1
7JnA7nTqFVPGkIrkROHYcXrnFs3iUuNHt8QRVlCFrIOFW6rLWAjLH/CuGKatCXFy
U9d1LFvPdzsV7rudPvJ/GOPjTU1kxOCpoa4jFnJkaV9iLJXOmeSeFHFRrpLXyN9R
Owe5lwDDMKt2OwzGYFaGKHOGQRkOVa6i1DbXj0SJASboZUzi1sbmr10oGXWIum2a
9Q1HqYd0BOwfWAtN447kqvrY4fEjYtgTb1dPL2p1P6KAkvzso89ssjrinpYzO7Vt
G0qf/pgZG3g0+RfDOSYB+6jsgAlJcEHUuEnvCLuzhAcPNESPCh6n9FlxcRqV675g
UZ2PweJ/QHhLLKSUIxRlrMhUwqs1zIHc20YrQt99VY031Ts1cXX1nd45q3poI2R/
6L9IlXN4b+HeA7uBWIgg009rMFfLH6pXZ1H/X2+/gyswYGN9HewDivgTc3gJSG+k
xGVVd5m7mlqHs4uy9iqb2gL7vpD9X7H23LLVPRJkMYgjHXMdMy6mFhiBVTw1+FdU
2DCdsODnCn8PbRBWFk+owcTYgvWrN0fzvpwiibHxCtoa3jNvfydKbTcRB7gsszt8
AEzozMlL7jxssbi+NKNYi5vPCxPqSyq/g0MQJV4G1p8UAMPQILVasd+RB0jLSdSE
/qKDL3ApM1JTDKpmRuq1JWLcrw1Pwejm4oko8JhSPtv+6YLWSJSI1acQeCVpGWMo
KvQWp2ofu0CLKiuReYMS5ZqECSSnnhWEzjff/cUKrDoI7voGtGnxJAjVV77Wvccv
Btic3Or/lEUtj02q4CdJDxgeJuWv1Gr05wkajG5AIp9NhxvcWmQL+dRZ+3nyTmTa
66e4Y25dpniY4TenzERwP80OsCyiS2xBTnbWWTtipCf3hZ3rU3D6/uW4yzwaocSF
swkFQcWO7Fd0UFi0v4OKZ1uDx9b8J84Gk+hhE/7X2CU8jPzT+wNHT+C5UlASqztZ
YIfGH0oMW5YaRa/SeLrcA/KUdR60YYRD42tZiOnldYjxSFWAR6Yjw/O2Slsow9HN
d4Cp4xk1K1G7k3WpiRpnW99ukGEWtf3Te9yMG57+KhpqieOjJtI/l63yE8JO15G0
2RIrQ2CS3QYUTt6xVVOw8UNB1F0UcSQwdYagHvGr8yqNb2HbRVuBZAPoOBAKzsUN
O2x7/TEyj7vCajAN6OehURteAgBiDEKEBodugVJ3piKtpcoguP23etB6zn6/Nddw
tDfKkFGzrRk22RAvkZiRA2PwZUn+gP8L87vN5NJB5Lg4fKY629h3kCNQVqF9S7HP
bS3z5bsSAx2SweF71r4g0fUXKD8NB+/+8shDcRXDOclkmEy7abD/igzALnZ4SAQp
KCdGs36Cj8eSyy+1CzUMuChaYtpfFXyqk4ZEm6OWfjo4cWxJgzNR7v7ebwGsmRoK
XlsWtej66h5EzPMQ7+ep68uC5XMXReEYVkFT06Ve9sZnFkvQo31sG8vl3bKw/V6d
8CpnRHuu+g4Phhd6X95z6ml1713vsjKF8IpWf46fEYutvS2ljqJvlqt+U7VR8FJt
DAMrxGYzN+Sx+Vv4YzNpCTd76Bx/NNdhOaMOCXPMmHZrtJLg4GJeQvYilFlEtukO
XLofJDCtsClD4n5d98ukf8fm4pyjfD4VEzakKyg0qY3If7bgTfNcJ0KJmAWeMab2
ci3YsCFMf6IySC7St7Qe+v1b5Ni1ojmuvrAjVOOrzJmq7fvfEa1OEt2w8zZnXBW+
v1G3u1S+YYIjb35+C+FvQfn6EoS5J7uhPO+hS9N/2f8E+PFMqU1puhcgIytTYbii
j7QkhvaffY9cqYxqext3E5WIShI+TvH7YnYJe3El/zciicoAV6c28GKkWfbb9lti
VPDmVgPpacX0rfhz5koW/X9YQZQX8a/UHSK+jrLDeSsUJSXlMEqNVI25PotvmKVJ
K/I36EPXmdd/VZGHm+g9jkr1tRYYDZFzeHim8cCBHKxg+0wBdDQYpxgMuQndyYh7
/fl6nptpf7gcd3TG8VELDBguZAIPCCPXM4m3oQUb/UTkzln709pd2vF6bXqfuIHI
pTqsNFrsFjiTwp1OJsYpUAk8IdpiNcDX8Ks1nhhjtTJRk7meaVHtPykUmYIj3gwK
5pcgb/MxEIxeqlqDK+JOX6tinbKdfis4hHYVUMjVRqKnFE3rP0Sopa7EKJh3HkPv
u+9YWozOch03L8h4GZBgU3gO3SUQ8Izj9FqwPLmt/yeDofvEj9SHiIquDc8MhVah
hJRi5vWtvEI1zxSixdGb0w+aXMVj60gEaDaFfN0ftt+88CSMtpfpkDsgOA5UAzud
/k2jYaGkLYlGmas4/IuUTdlO4mUfCDnQjWj8VfV15HIjL7mlksy0vR5pxp/ywc/n
h+9gL1vAEP1gSmEA5I62xOjRhf6y/khPrC9s0++xFLZaMiS52/ajZqMkp6z9H+S7
o0FSSk1LQwbMJNeMWzZ9YIl2782WDivyqYzI9MhYVQC5Kp0fxJ/tu+GOJaDQur5s
MBJ1gH/ncCh9tr8Gf1KVtyhb5v/Aer0+IYQ74ksY4wVKak8vxOucOcGro4EtfvLC
rgUond6HHifmfYkjgxw4o7knYSj0cO6/PQq/Qq4CfzJCHnB7GTuR3Kwfz2up51/N
o6iFndQLUOV6yK5uoj9AZhtJiBfFq3B16U6FA0JiQ657tFWwsJkDmdgp9vHRW/bT
2Xk8qq3JTWD6KJwd8FJ64h9x9ERioBI2A/cLDZtez+xUSKvjgZQYcsGKzcHkLjn0
PpJcCmkvJDdoRSgWYuWLAOVxJODWWw4SoWLf7mqtAP2cFaVYzQhZw+GUN0mlxzQ2
TjbcEv2xdsYLYAKoL56V7vIglj9jp01uGNGTzZKsWehXu5gsMhCQVSNZZMfrYafu
+z4bWuEDugFDl7YLstTWcV1XWl835ZslZb2oy5OVh5klj/cV8I7O5WrN6YzsXY/d
LUypWeK2gwgEFsNLP4zqt+4ZxEfBSSQsfKAitcJtwCrhGrB0yNHeftnehYa/Y+xz
hGjcz0nDYhaGG9RVww5xowqjdilwK3kdgLoYvsQzzhosnxCutJlTPvhqIcCotZ6r
N/iV78k3FXCV5BVLy2DhpC8IqfcI9nduP8B+XqRF3/u+gjjI2h8MImXiB0nf2qLZ
CEGWM81ef6fendeZovZyi/oOQFIG+b5G4zeFf+lWl2tTiy+Rq5SvcNKZCHK18ePF
bkTdApKIvBD7quGj0FgvyaITf5YmMt3Udz6Ek6sCdjxSk/9xLgPRLi1XL+kWz+ex
KSIc4TleMQRwzWqmVPVcQvH3P17NW++WC8C8FXnwimrrejaMSIvfrQCJIi0oBqq7
NkFf+lWlTQvBedF9Ra+4YAL7AKshJqpwWdFeOR8lyDfo02nkWEKgMo3xUsVDiC1r
BXrhqcmpevFOqd6772ufu2R463UH3jxwPHXzBPNg2pJGOtsa/KqQsqNTuhi+0VD3
PXIV287UBnGphzTIboQJz0XVkXk1wVWkJE0gVl5mu9ToTsusa1Diy3u1ySICWhk5
o/oO+mUrotzFY2Wcr0JyN/2j3owLj3M1UN4xiZtzVWSdZ6+Fj23/gr4128s5EqWC
Wa173AusgdLSuUIqvAakTcEkITEPkKm5cNrQf5Li3CJoIgkIYVAMnO0YkiWho+VB
VriFrl3lwStGTGkbwM7+EakMTOolJLE4dcTPmS3NRp6k/O0ZlfhBoKjO5hVYxaBw
76hPJ16EdRhZXpdgOSf+4QGHdaI8c0xB1gzYGxsTTw441+bIEfbic+W/RvjV+2C/
Alyx80JXGlr8lrx3I2fYfJP0YQMXoIMi9tiTEINELX3ntlNg0sKl1oRZSsdrtRrk
udUcnQzfbw7J8SpK8Cye50yYpF197pFT6EjqMvhqasZ/TWHt7RWXAL5ZxALDIPol
IHTq0Q+jwwSAXr1+HK+89o0a8tq8idWOvkv4n6CSspO6ZuInvIg/ME5akZQ7b8rU
f2dh/3ophcUoZMJDFMegaiJYK3Gxvwx1JHGYW8y4rjcTm37zYELIIxk+qfimtyMq
AAs3fPaLRNxoC6eohTCm+CsGh/jBQTJoxpFFc7dEry9QGkgThY/6qi3ZdLOPgnwu
C+4dUDtWb11R35sby+ltE1cHsCQteL0ikiRuIQwXV8EMnnWn0aEKrNFo64HBCQcs
bkoc347lUfzbF2PEgvqbo/Aevs5xONaOEHBBuSL8j07Dyl0SmlOeedFC4ELZ3m4O
0Wm+kL+mtfAzN7/poBoHMzRtOqe6LfjpL4lbHYcMYekohWjvICETwzV3eu/q5StK
rHAMhIQaOHaPodn/MREF60Z57FeL+NcqNKRRpYfk8TlL0y/yfd9D/bEtRvCxPW8/
D66EdkkeeqRvXpommHD0WACYVJ0A/ciM1d44XP9Wc6P6icRaG8ETGWEVrX+/agmp
QPB23wuJ4vrMuO7a/OLQuJTVrZDBIq23UcBQlcyFG8Chcw26ZUc8v5Xj/y9bU2Oz
opR7vfVWDTCVxHQUHLloLZ/mTdd3pXURRg9MJhkaiQzswIuwkbIJQgnlGggYYpob
kiohF6SXVAkmA048KdLicOY7BYwcQjD5AyoDFYBteIUQAr4lktzRADEDw2jk2iAQ
d8BdX5Yna+BPzo4UhCew9tHOPj9+4m5q2CftPZqOQ+IxhzRe78pJEdnXQwsxeAd4
kUAMBuK3TRSPsJd8W/iqyT1cTSGnGgaRyKs2UOltaMqmwU5XtEsYdue8Aafs3edV
W7Puyo76wIjdiUBX8UT6YnoI7f3j8O0IYZUPg9YLhi5/S3CVutpSCUrRxcsQE/pM
NdjRWc6CoNKgdSha0ODhzKMGjTzhNpdrZZvklFFTegtsi+7ojZHNqf6dhxjcy57R
i0xrZ6e9GDmrXt5b8mXJh8wLrSG1seQiBiEwb+Bl7ozMzBmO6Qux+lvU/NNVj2ts
5fVgoK7xbOtbXsebzpROHwgbB7q9Mhhve/yaZe63siff1IoKzZ7KH6nvEtc3JqH0
bXpeE+mD/CmU7TBvJmqoYpOZeP5dI6+djMfmPSkIjkK0tHw0atVVGYQeP5LInATh
XFqhb+KbNrpikF/dRNeQrGevmAhSGfX+eiDgM4wnKfowB5RvLh7czedLZ/AxlKh8
llgnC6Y7EZikny702WWo871hbPxhGZKgpZUobDmybZOkzyEcU0ysu5YYPyUEAOr6
R40lQc4zt6ewhtBXG0/9k1hEXPaSmBL3EzQjgZ4wWkqyJoWTX8ygKImPNIrGhiwU
fbkPCKzyQplT+dJVxpHu3gRdEYjkKYC3M4SV9QfnxR4ghvaitWsO0wLQ+rJZZPeZ
UhStk+Z7IlRPp9wi325dSrNyTiOW6dV4RlxBshbg4cY2Dv+jVVE9hk7onaWliEaG
mhkIQwCVWmVNNbWWjGi3sdaIka47tmi675XFpZ+jj7TAH9uDU+0A+YPUi/idYzjU
OIV6VSGARO7N1mAWjO+wr7w8HfVFmFTjo45o3TRZEFNKCGMrXTCM2SKDhaiYjqkq
NPSb+bgUclxRiZBl7A4Xos0i9Pgal0G0CIGlXPcFQ1otzsqUdfO2M6jNWnIvCBnG
bGL2rCK5kaUZZYNYvURduBmFR6BxNvcqhsxG4/salYPAUWPK9+Ut1mCuK4Lqtqll
UGwMx4nlA9fHFI0Q3KSZRLSydZK3WwfbWrL9P/8FSCGA2JGv4blM5hoSnlS23OhU
CrBbVst2or8Rkp/Nh1Dj/O4MjgUG7/yM+lolN65+7LIX9PIU1vXn3FqFH9B+rdUJ
9oHuraX4sRqvIvtO3BWdWbGPS17VCJ6V4dUWG7w0QCTEzwfGPa70GulXrICepReL
VaihIdIjO51pgcrdUo+5Fn/KUVqZPjcy4pStsXu5s0IljcFZ4HnvQ9Qkh23gZAyt
X9tOF7jqgQH108wIBDK/SINRM1INgvyRySBFNfHylUB/y27FWZmHuVP3C26Qd+XI
s0U8/SGCO0xBvLQWbti5oQgQCwwU/2iYppXbLLLfWQgaw7h2b6E6q4E0qOpFnj/r
8ETQeWorKVENcIurOYh9yxragkYUcGFAMfOCxlfDNyXE9yPvowjgFGOR8U5P4AiM
OLjM1u4qRVGdHLgSACd5kiq/IxAM+Lxye6cFBqh1S335POpi6+yIDz1NG1+dn/UT
8KQA5dxT3Ejr9D6IqudfnCO7JvHdS/A8ZBCTn7Uc7mnw4yK5Z8ggB0Qh+NMtwLnW
1TZfB3a58ggjYKA3iNK8uj96d3exdPnLPcK1rzjk5L6/VacVc5qw0EPPcDtTaV1o
X5NIG+JcrHmvQSpTjIwiw/ZTEypQrJurJJHoUDR60dPBpuM2L+VICsu88t/xdEcd
tu7HTXdT9o3d/PiVcoIF58J4r8q8/DL5XALWRjYMRjJNhTflMMJMIOmZbnGnIgCI
hneBiySYlT4Xt6d7c68pa6OI83hhp0+g91vYRBWiPUqr82zC6we+IlD/o31eEJY5
loQmYqAmAoJHYEEKqpX+xXc236JeZhRQpPMjqraZIS2XfmxhC8bFptVSGDr3dhXz
FCMaaVHB/JOrgB0595jA/bGfsTZtjNFmoRqmghEP5xWcB7tcyIX8VCRf+6BGyJK8
p8jayzqduIk1kh8REAvSU/oB9x9G0G/y8gJiyP9yrt58c5GgTgsc9w22+WtUBoqj
Xq74B2yxfVYZAdSu/76fyz7y+dbk78AJ1uh+9zsJ6dDmSE3A8xyNZ8zCQceZ8a4C
2znk2g6b3ZwOOvsoAVlk5hLpbkSMc3Ax5wwEXshAG7Csz7gl2YkKpqLSehE3LLoA
c6w8VUezCdaL9fiJRwIWj5JN10VA/Io8AGcgcV2drelOiAUEUM9G96V6kvZK0Uos
GsiMAI/z3d+IAddhkXM7sCu3T12OB/hJRjiYQ+2Afm2WsyF2k8kKDANLRC0MY3Mf
ZRupLeSZBfHPwHbwtx1zKCFRj6iZxZVfNWkMTW+k42CRfswA+qjSt5gcdeLtcUqG
sRNVKVKb9j0S/7eWrqwySp/WwhklkiO2MuHftpGCFrKSDNqJgoxu1EyCVWFSKQaW
JTCgx5pNzSBffJw0XHRZnl2Ct4G315sQ/JXANgb2xOthf3HPeIDOIxicCEEep8zy
IdPeMGjIEB9PD09owS+g/wE89huqHET6ZcC8WONHGM8nbLlN8jPwEMfwpywI10iC
FUXPkG97g8VEiRi3cpZiZPu5KrYOC+BAtX+Z97xnH3X8I/P2q09YtL2qhGV0ffA5
6F1fKCTE2YQb992OEZDGcse3e/TM0f8ZnMIpKb590HfwXd7CH1JMzA77UXW9eTjR
o2BqQRtGtAuVfPKep9MWnXReJSS3w7duU6OUddmtQgRx4U+sF6KC/3puFV5nIwiO
OmcghovsOf84ISGmToRDgKtVzZPeo1iJImMamM/BNb3CKYWNxtmaLYidIn58S4cm
T9rCo+JvYdQ1Icx3Hn49RrNqmlib7rlL1LQzEI4aF0JhiwsnKfXNsaQw3208q5ic
D4m9D0Ye4K6KwlTAAV/dJZBzBsRYv8on6jM2jSB0CQi8vAC95uZmtR+dsxCkTQuv
hk19WjPnVR+zvY20+mAbkj43ciEYV8vIsO/xOLiy3Ci1O65+es9SXA2i5926fDsK
JYQNTZO/6jZm2AbjyraHYjcsdAFAr209z25u6xvO4zX1U34Zmv0y/ZD3HGO1kkGU
bt9sQEvtUAUdJaLy5YCzo63YGjHp/t7nANjbQDkXtXsQr/2EV83gKfRSxE2nvAMk
jjJy57Az7CihiCtx4sCTLC027k413c5oN5PHXv8XTMPfHYUQB6Q748aEhthauOoE
SVO/+3kLe37Uo/cAvUhaAxT2L/jZU4vyi3eQY+V/IK3tLkEHzD6adlRIB2qGMeqz
8yBc4ptv+2FWkTWTM0UjW/ed3UEbRrPxBGe+IQr4Hs12xb52paKRDcuiA1a/9mXi
HJXcagnXgzBQUFKlp8f7ZetZgxjqYxK6SPMP0Nb3ZylRJU6CsT668l73KnrBqjLk
2RrfMlQ6D/VYoEW05eTOp1W2M8Gl4Hg4oateNeWfPD2adEtAN5MG/AygrltnlZ3P
WmP0c8RKvv60WHUO/lluGHkYSF/FwQw0T6680ThKLJWD3FUrXmfBPNUykR+3YdNr
r3/1OyNcSPX6x/ine69JJ9rEJZnEXVmqzoJLEXNSaobPf50t9BTff2hd/rhjPsqF
Qo2ayBQUsnvdMEwYiocXOQs0lr5KNiEpkVxMQ2MlZdqoo2V4q+sc0UJYYYlmZSJw
YU1mzLkFxEc7LBuNOifRee9u2ARTy4dbGWfqEphH5GsDELFuMX7mFoD/q8DaAOen
SK76nWKs5cwBmJaIi9vAk5ZUutNlGXk6TgvGs51k+ZPFQN8SBfKtBBwp47rVNUq6
3vPBkOdf7DZsDMLngMCoIKC0E9kH+ufzdFRAjLfRarD774mwo6NW6NcoRfGhTiwp
yl1qRIlauRFgiGKXwqkJROQETUn9rNN0ymoAj8qKTjLUpBifMOLvqBlzBN6ys91J
cwPHBEoIXzquIfR4AwdVNRqZOlYoRrV8wfjMnLGsvtdoJbXS3dV0IqNnF2XxZIvd
riYN0TINQm8xE6jrPioNeUbt57q5NAswW6ung/Zhri8IHDJtNh5gttfw7da5iLgh
2tznAvt7X3btCg2CZVjhDELzPLFSJVjW2ZjvNd4Ug1hjrkw2XzgwEQuUz8yA9HxR
zv/1BzE+bY1heaxHYMW3GhV9j1FDxNfXYtOrYEqAmp1oyb0TUkjgWcxyzVMcM3xK
7vAHVUpiaVy0Ev5HtO3ILENuJ52d6eZbr1viOiuO7nP7PWptuKel1ubZSyeJqLjA
Igb8GmkvMfjheomlbC/dMkUtrJH+0JqPGAsQkUzpyV1uZvflpQwEAABoTCIMs/bW
CFEs00pf8GwCrKWwYMSXwdAoSSUhaspfidp+oF0z7FJPkjm8VR0xvSkHAdyT5NMa
l8sR4+vU5yJfSdc8U8/pYHAEGizJUosLsfULxZ7ywy8cNs4D4qWY8QtakICGA7iO
6NLDATRadVuTipS51kz2zTSw/i4bicaSNpPnkn6VvUmCSdD0v4QV3g283cop1r1j
mEIbl2yM7WzybkceJ7/CggEo7Nb579S+GlyHU44FWmXIvYtBPLw3gMdGgRY62FVv
jEZnCmMC4zbBSJd3Vo3ALYKcVf+FZWG2YlAGNolKa/2rxsEnGOdCdmWCS+TbCw4r
OhuQO529xAWWcw135n2cqJdDpm1QiN+aXiAWyXHp5sNbvJWgVBJa3eeXuJkGTtGx
L7MBRk8HhM1igZqYxn5z75qY+Cu2lgquUn5D7matM3QNUxhx8WjGG6UU4Lhi4ZF6
4H6cIuAHtFWBmjuz/6f9IccOxK0ftv4tOqppdh9mSrmg7xgXPAfRdH09aqzncVJM
c4gP8/zQKFcvVcJ/BGIt5GmFYXS98qyix4cn57kJWfdLvhxsW62clvBTwi9bHYMX
zvvpyc5k+zMxuNmpAj2bC+qJT+zGcgYD2uMVYsRdun749lWvHX5uL8Ub/NWyxjTK
FMvwVF0x6GLUU9rQwsMwtEZHN4VUiQSEOoUp0d6/Wq0J2aJE+neAUYPFbREmu/Ol
hdlQtBIgesF8T0yVJJo3iT4uWxX7UCiPJOGlBooPrM9Yk+ZVapbHk6R0YZAXLE5H
ijQn0OE7l/CF97w9OkvEfRpsnnEGLINoXSq6gJZ+q22D6qG0N+s3S9aqZ+3yY2/m
bVJyOI8k7FF5/H1ciXlenlE8aizp/xRqvaaFDtRgsYVMghAcEWHc19Y/5Su8joqM
iArpdF5rLvfqHC0/Bvrjxo8mG0dsmweqsopMXsYaQEM9vBv6iu67Rpe981B+6vt7
0odJfPq2otktJJJtPD0tHFIdm1oRboHLoEgWv7adfj6ReYBblmVxKZ29vwhMcmmJ
gIVpF51BSWMxaXEv89rjENq5DIZVXzSLXHYGrQqLUy4uIt4Io07WNwBm9GvavCF8
OajDvaQJfgv3nya5tazv4d89VZ7smppTEBUIfraOcaQ4pFRWjSk5jHfrIYgM2bWu
i28Ty2S6Vw0qX4qLfX7w7Nni0oVEMgVcoXgCnL5YQj/q4H/f1YzcxY4XLU22ZQog
vp5ZpU5gK/PXqEXIHkkSKwvilLs15Q2vRe2++9vJ6TnHXpB7cpkvcBvlKcIsKaWL
B24w72KVod/pGr9oNCQRNCoR42LOCInhlAA+pksEeBhhzMJxFUmWYIXpE5ts1+/g
QVcOL3gJQq9PfPfU1uB27OHFCuDOdssNbDWgGec8EpkSSySSlHAQH36t2Crhg05/
w/tsmjnbiXjj75dyi6Blb9QvSyoCLTSUGbIsA9W9Vg3Smk70T2U9yygD79FNrJJ0
XbxwdMFg9VUbGsyPBUj5SmHDhUU90g6noDJd1dc1WzLBVNJ2KMFwhzjG0ZUI2Uq4
dUBEL14Bc3+nabzOdiCPuED/iNohxkBB6eeCha90myc9jJyXNkZPxcDQbD/69SfF
n1blwPIWRc3+CL5nEdOZcN/KlQdaBKYrYE98TIcyef6ZjcYKISKETlnPqiNr0hhf
n4SDBmWPlK/RpkHAM9MCbmDA+dh/y9IYrcDz1DT2+vLhKwmS8yiOnwU+ilYsfXdC
O8SuSgPa+m39DrjRMwBmS0MSYPYgbZy/WtmecTTDErvGILWUunqqIDzEaLcZjVkJ
TL6z0pdJY8JDC0o88l/0rY5UliZ+/8NFYZkRQhjt95AtaF/KvMV2TeJ6+PYfVciF
x8DwOeGq6VvULICFaboXGQc+aOmeEf3PFjk9ngPQdUfAJI7bTqmAs42a/PwzQYm/
znOO7fb58/Nwms5ratQu8lFn65F3m8OCFYebiLAP3iEY91EHqWUJu5CHEVEYK5Ru
JhSD81Mib7JtTRia09/c6g/CfQR8lxDHS2fZb8C+1dCTjhb7sctf9bFdcQVMwxga
ku90UNUntrXiS0ym9lbhzVmI9s6rU8s4qaQ2BrvaW80MfOdc5VPDqLJMfh1Kf4eW
gRBdG5tVyvlz2eZJ+asWtblvBwU4w4o9PM7WwsnXLzlX8nHYcD9SydRCiidbO7rE
cV8J5S6fj1YCbNcmMWlNX4NARe16Z/6vQpl5gwc5wEc2ZBqq8v4e5iLKkmSfJbXo
BxslaN4CEj1Oac3ktv2DKa4GTUOMmFygDllV634OOEvvGy9KiC88enLaR3w75Pf8
1YeNpxutBGfTNz5tQLhTBqma7gL7vjk4oVEmCYxV6zF4bas++WKMGZSVgdEg7Lep
Jk0lU/fJt1qtEtbDUPvRixPTYvJvhxdj5FVL02IJS1Jn6E5up7ePip3X77xnx+LD
qvdw9iBxFCPM7zdbU5sZgtcLYskbsUa28BONnmAZifkRtr2AZ3vm1MeWyKNnSF7M
VgHF+uM/Y0kcqaxuZnFF+ut1j3gh2C+qLR3klaIK7WEqj6Fuufn/4HmVYcDToSry
GRJzFRieDpFomm8HZLL7iq4Rx5bGSb/LYjshrAzZEc2fsx8cLt4+ri94VOtIWDC9
CHm/uqyf7B7dXdSRSD3TN1bVDoBei0WgRW+If6T2DEwwrf9y1gNLj1gSyojfQ6iB
lu0ROhHyfpArYPOHDOerWN3JDHLT4dq+CO2gGvBodWuk1N2zTFx53nx9oyBLRK/7
YfLa+FIF7coOmCRFHe/zsko2pNSRAvQqQMtuSd9NWBOUCRpBWC3gMIdwBOjzwJQQ
sFmsPfrTmhuxdIWyHlsdYJN8PNPxUxRWrvZxAYh0TiPC8mLB7Ify3oQpIqBZQH1l
Vgh5Ouyfgz8uxgZdnGFIfhlhlpp6OuqxswpD5XGRwm25qW5x51a/Luiyy6ilUBeX
9qwB8LG31vdRL8LPnLPKJVRrd1ED+epSne9fj/cUEmozxJ9dk4vQJpJ6FitW75aC
jyy//Rz1nPP97MZ0eK+K8Sjaw6B3MWPJstMZmBqDjwWYSRamYlkx3190TMZn0QTK
pSvpYYzaLnOIYvaB6AhLMpw3ENotAFhAf/Z6/8CyvSU8R3hmo4+2M/O/leDQI/xf
qUTp57cI4T1VyYUlHRRdjxcyqQ8kG8unKgtfgHo5rmQCUhlGsIg5KUG1Z7BS0ULt
AJsvADvO7iMxmrgbbk3jyY/L6V8alJ5mak+6k6oe8+WRKFNwJk+S75HmtI6q69ml
CQNK4QCPmrVILMedb1BH3XIy9vLjS3In7obGkSVCfM/qK0EOzrnWoqcY7+AGv6/q
cylhlG3sFBjj2U/g2FpLEcGqkUOpz1kcaL4F0PX9bUUZA0bLXkvz6qKzSGdkcZMZ
GXYnWdiCBFYPQbuajdMH1bDLsDc13q2LE4daNqdKncdIQARHL2RRZ/wmRFUkZWoY
d6UB/E2fYTNQhbLv6SShMZgtt0M1C4Yt61I5G7U5fmcZyWVnrWhYvbnobJjtqj6I
Q3af2jc8sBEmSzjfBdKU1jtw+W/tnuYtWJlfUv3I9KEtPVdRfoBPWFLZ0vwWek4z
8P17V5mnEZvYzgBVE7G7SB0sFlwFDXnnawyYYgrX9Vj/nP6zE8IFO5AJ/3rs0gUi
ExvBe+O3RxAQSUYZ33J41MyXbvCLQwCqHIZICY6mHQRLR7cllHXEhwTRQmg2Fcrg
9wJ7ZMS/08H6XjK2npNN78vVC2VC1DbjHKou7rbZOl6v16um8C3oeS1KnJ1JgdAm
Pd1wJwZS8AljJkcRVJarBgE2XjH/jKtpJRvmUlTSzEeDbyZFtgutguDkmnlS6QTU
FOmcrNqqnQ0WTBfHSbWUevE3D5nHePNxSpiyAuuYABaX4YSj2NUzIx2FKSZ4CEfB
W9sODvD5R/00rW6y9sz3KOjuq8E1mClJVI+nQSePeAxmd43l4RhfM+v0o6ewaQcn
yaoQzRug0U6vm4RaH/Z26B1HbDR24fqYTdwOhcSHH/apHPBaca/XBJSPzm4hcjuG
9QdZeCdAz3+FAgdR/gfq1fFlS/lPxUVjmHD0Q4+yzfxE6pUg2YzMB1hIaaRS38Sv
FP4akq3AgIYdoqqcpsNBgvLRrPVY0Nr1Ub9J6zM/sbwA875l+DBDE0H3aAC46qJ6
Jk698PbKC0F/sePPewUpAYlyq5mvVg0wh+uPiF9UlwK08kXWHRrtNcIOPe/V2sLg
uhGv3QdRgXmB/9tvu4lN54j7+uOCIqFtFe12Qg9Ipyo2iBwyO5rCedEaGbXbNXZu
lHQIac4FzT5CIzQbzh9oAEzy6UDZtHPGITwzVlgTSDG0rIj5zT19F1//vGKbeu9L
6AtBL7D4c0oVHbzhpWoZdeTfoU27cOAEzTQ2EmMDZT6PNIkXKyKmQ/myXLWlSjbB
Dely+l43fXhfH45QckzwoBZM8ibfmrco7Dof10vSL+ERWjxSA9/E5xIgyjHt4Kx+
KByHehVBNjFVO9jW9+FWaMUIDpWZoCg82FUt+TqKcxtJTp3ycIa9zNtvRV7zqOAl
9zrLpSQRTFpxjUmLQJi6wGuDhn+5ame1+Yb0P1EzwQKDm4QO0Si0V6+2rDL8fnkz
Y39gLekqmTzIyJq7CpvTbtmhP2M1Cu9q2B2G2yWO1CQcY/XmdrK/44Go6rDrJjfG
q2wxZWxGCALDAh3+pcaKsT+j9CyQMMeeOJELIxZa6t5Goz3tmRyJxhzAgMqB6rCO
BJ1g/DyJZZGtXqbzgp4kNtt9HPNyN2pp4qo6CcV3278QTEto4oBrU0UtCUzNk8zZ
0WAz1dqCCBiadUUqh7hRkXxLRN593Ku7Pz7LnJ06HhnvVO8RqRrb0I8c1fcCfFhC
64j/c3uhpW2VavPoyb8GDzA7xJSbwzpS5x3aQ00S3aAKSv8LJtys66eT6IPfmeOf
T2TWRHSG7Zgvfc9/DK9VC3gQa74K32IYBzGDED8/EjfxKmJ4icYSW3RVGuHSoh9Y
t9MhgRuZfhYbyGfjE1/vk0RSezVaYG4XW6+b3ADEPUEPQFzCZRQsOMP2kuBebrGf
ZbG4ds+/mDwd/LuXLcB07+mX7GimmmCYas8gNYC3kUWutaS3HJvWYMgIcUCh+w+d
in3SEl8Bh2ABgkmDPc2u599pOTlo5kfUeD7gaFMZRGG9+o97h6zLUtfjZG6M3R0S
X5MQjXM7c7xwKai1mVnjnz3KOrx3ABgvyUxOO1L+V+p2UlE9Jp1OT2D6EPMZndiU
H2fFGPbR/9ThyRTH9FJ8QUwEmNQYwF3jcSw2QjddzXjUoorTNN+E+tecHd5BBJZO
fUR365SIF1Zp/WSP2pC+b8jQAvRmEbaiui+MVS7DFKaMbN8Aa3fsu+YnKOXeurMg
HTUYNvDeAAzG0dcwP1+v9+3R0JctktvagDQG6VN2xWRiVrPFjBIoZFg3B/OO2Sc2
7Mss/VWxGgq+bybYm1Rcs2voqvNfkh3XQLPr6o0znpGilR0o6weMDE3viPboRTAL
L3uuedVvmCP4hFOLROj5gBiuAq3E81SR77lhShB5EZStXmY7WKhKPPmU1FWPfNMC
jmWkeCkndhCOUkjYppB4Z8WZ3QTgQvPp/WedjNGyhMtbKzxaRIROw9x/RCxJ+PlE
2gHuJihWagLgy0kOrWr2/KMKk/B3UOn7gH7Gi25RmrdCCaTMOqKzV7fjX2BJJpVj
GOxCHjGcKES5VBX+0tZ5tZ9GnrUE32iNx7bjyrLNfImhkbFnYPhYkb4haCHs9y72
09tRbmE2XozXg+eRLMP5oiCELt2txa2zjkeVxg+RKFbQX0iNtvgb8wP9K/pltJ9e
U3wWY5PlceVCFl2epcsZnPmeh/LalAyoUBswK2TvzCnUSNarig9gmJeWMBpU2tuc
wAL6cgtwYtazBPVAxdc/WxKxMw9LhYlIP+IHeUK7HI1v03tQnxbt35oWwdTOpjbD
DOqmtyaUC0NtsK9nxgQz1Kt0fkjJWL5YqxiNtbuO5W//cF/YQAO1PmnqTHvizdz1
6j3JhbTbkvbzUYsq6X+rqjc3dwGDTNeYYM/OPC9TFNnZZRSEAbxyljFqbnigraAc
4lU1Unv6GrTbGIaQm+T0JvzZD5LchNDKJjVuzcMjHCPesaFQoF+nYSpD6WPZnLzz
j5vidVmy5qWFn3M67NCzblJYDPKgNimsXOTLTEJkxtObS/eahqslVCzCMchOOoar
jte4ZsxXXCoSlk/900NUQ41ZvPGZMXbSsjT+VuhIPsUKkRnjhWL20JoYkyxaKLuA
DctIULO6z+3OCPQUOall/cIWgPJ8B871l1xMdvAuM887Fx38S7MqlONwq/AcXiVf
C1RtC6ruWnnflneNm/yyODgMwaWf2p8L22762m4vtcj8bIMUGOF2+CO46kdrPzBj
V7zxbyhsNz9ADXwVfFT7YaUuwZ2nmZfN2/Cgaj/gOwHx/46FdxedXfKwwsEGvH8a
mWizk9mqU9cJgcnhoD2z92aTXqR7azbhU10CFYra8+DyHVnZeUYKepaOfAkgiRkR
Xe896YD0Lg6cwmujmTLmrUj9XP+32beNVMYguMGpHk3DjKUW5YZzfS4jxom+c+G9
4Q/B2JrugxN+t5HeGczO8+lBXbs/NsHQvHBfPCY1PAR8qqlzAThPsvmINtyA+jNi
gg72wbIzGuByFMu83aHnoslKvxuEjUtm/F21zWBy4aqhkl3DabGqnfkMf6o3bROZ
IePeB9X2PVMykqQXBg1TzhoXw+wUwBKWTe2GK6JUhY9un7C8WIItpUIuZkd9EaTH
XQIGPGXG8H65ohbAVYUL0/ptIogKJT4fpu+ghfeptEAMASmilzG8cJWhHp4LoCdl
eq+qWN4n8NbHGFLXeP4p8NH0mTbEWOBLvjPXgDrmD0CrtZatJfIGcG6lbQCkgJBU
z+Ji469cU5WeqbZbBtTlUUwtQ252TkVzB/3PhXeQCOV5uG55zAs5coOBwJ/letxM
YAFLWNN7CQVQW/pfMsv2T2U8rSQdwO0Sz0GaqIGinjt07hm5lNEq97EfY/saZVcg
bOC0NbK9c/zHfpZdZgPOQ65S2+M9UBT0Di52tYzcbZjpV0qRk6to0kdb9a2wFOD4
K2wICE5OjHQruMyP90+ojOeHzaDWMGANAj63O+R1icON74qlkhbX3aVKE1o4t3KV
6J+XHw38QyPxAM70N5gsjfCgaWFqXoPNeSJPdDy3hau8xACY82p+w3XopvWaxgJg
Xkjspf2EECXiC/fzt669xW8DUPg6/PGDCmGYACPLacwbBK0MoG8FlQD/COy4PdBB
a8KyQb79rwF4052JN00+PP+vM0SfhsHcLis2pAIMpVxMcLqxXEvolKXqdSOrc/zR
Oxp+xPqqO1PbKaIumXUg9uPdJu215KGPJ9Q2CtBjnYTA7K+thvPWTDAq+IPPRY53
2nN9s2pc5VmeIDaHXd/WoebpewZG1q9NnoOpZ2+S9tRIVVcIoHZ2OmxHqNUH33Qi
sSS4liD84V414wUZtzIRSUt7m5VzfuUGkgwMFcmt38LwwKJ8F8HQ81AKHRGtq3zc
CWEzNcWEHdPhKZrNOq1WfFXPbKQDMq/L9Vopqm0x5y2VMXO8GneJinLuF/SuUxcm
0HfYQOq+sKiqvDoZbKZ/a6J7gwp8Bl3+jXvQcp4+yKJgGi72mc0jf3VvsqCRl4bS
gcm/96F4Rv+4H9Q3Dw8CKiQQhDGOHzxE5vshKsW2+SPjELUcLvFfvm1WX2/9zEPR
hmzBjdmVDMUYoGQS/Lx2CTJuRRkmt7gNJ7nHu+yB8kkrEJUHP6p5R1iPPnQRK2f+
ndWL1BL7ifaxcSOtmQvUKpfctKHKlSvIQXwMXXxbLN9T91Vj4s9V6S8heeODRHsW
KAyl+uUolWIaPOPEVKFdruAAz6W7jmMOfcVRv5GiS0z10oidTGw1QRiXa6RICtE/
x+NkFhlJPJ7pUWeJlbdZpPAPeqR5oGmZrwsXEDt1rhRA5tnSMMD7yNSAb49uO6DH
QXS/4fILtAGT40c1Ig90dxszGUSlU4+DxOK9M+AMWkJmcoHX+DR33V0WzPmvZA/+
/jlRoCLY9WFPqMTne6cb7RbHMmtUDn6yLbmw4o25zwdWLpluO21nikFyLnN+jprS
jaiC0WVXA1oMLIe9FQZy+ZM0f36agQpOPpfFNcMzcRZmpBwiO5RFG6UnL7BjPPsJ
nZlSBlQv5mLf2ZvWAQ88eAnb0c5eQRgu63/FeSBPz6dOTTEU2O+L2F6itey/aUq8
SplIXuv8/RUka7+CtO5tkh5RLKztgGt9yDLoJWzFwq+nPfnJ5whOXYYD5HNiX5zT
cZYSRkJUCO1CjkJ2PrOgFnfOBEqcVntF0cxME1pZh9srvYU0WxX1uvcoBp//uuOf
Abhnco4jplJ+Z94QEx6gBL4rMDgd6JvxFG6WFVsAEoNfja8TvTi5ROFG0UqpvAFB
g+dHFnJJSNkIptM9/iL6uy7MH7zgBsL+tgTnKepnL1Zlqz/iDNoda2Y5ZqXy2WdM
ZUCwR69nd00JJd2tiU9q5yhisuEgeuIyZxw0Z4QbSo/IkaRfA656Cmn8xYJxfxzB
eBfgW9PZ9NZ/gSn3u0qjwRbz1NWREu/Ls1AfBW0G+hkuODg100fAksg2IeSflpMA
zlcCPmFIqFKJIS9e4wNG/6u7lw728btQsJW8K9O5FVPaIRtr9wc0LisPht5JuLXZ
j2MaRHx8yv71Qs9r8IMZkJuPlWrgCsZfs7t3qWryQlu5xYJ2xwb+fZliFsBGflZ7
mOw2+Uoolh0Fh4SbeRj7TT/SvMpVFvtpXbsGpkgxDu6dBdpOUq4i8x2vYLRw6+cx
JW6O+rNVvkkay8G4yj3iu0vrFSWDZqZm06Q0BnjIgApbrp0g35y8zow/clq4iH4o
PGFWh98AS/7qAHiuKdpF2uudPmTG+54e0xVCrFSBnDNJfytTApMbMcMmG6/GghiE
mYyKNjW/NPgTpthMwgMYgkvbTjHqJKOS9i1tZhY3dTiy/pejPgPCs9+Qsu2adSsK
xOCh9z8iP1G+NNEh7+D2jCcm7yxAtMTRFkpK3XcyJ8PgCwKkFhWKBGbeWhbTACkn
bE/3pc4KHAvcILX1JOcSy70a6Uahmxfm6vpHRY7mNgglNdvoI049uT+vW2Iv+rPm
mFLB3ibRhzx2pcnK+xNEwDJdBsX3bEU5c2H4URP0OwFw5MPkVetcLI0bkWg3QOnN
UfHbh2uH9D8i6blq31Xs6bsQluLcCxshiGG8BM5mzpcfLTLtZi646HTg0wfb2Skl
RPDlZpKZR6axi5BzxOH29MEwsaqiiuEtebNnLu1XGglUETAWgpVk2FRKA4cIl3rM
uRBE0EqeuuotdKWgOAtRxxSlZy8EvK0inyuEcOMC1rs8TRJplpC0uSf+FnLOV1ok
OQO08qdspz4RF3dK9cnJZlYBFsrKg/Mz9fIjFkN4tfZkGOnctdJt15utYhD08oqG
XulgZ/5bIday5k+eno1givzRQCsL1cdphs82U6p1r8ql043nCQv+I2pWS+rmOBwy
hGyf65ebp01gUtOmCmhpaCjZ17acdikksQ9fuSBbDWE+Qjfon7ecMi7+z8e3Wg8z
+wCDiHkELZFOskMMKaEkh6VhViad4VBNxhFJbpa2UIHwMCIp/YxhmuwfUhB8ckMR
Opt6Bd30gA9IvzaEy4bTs5YMgIqTYSSkrzzq0zpYeuwvjeF/1K2I5OnGMjKqO4cp
49YiWqAka6bc/+6W/d57aDrC4VL6xwlOXqOoXHVVvAAzk5SlWlW/PGzHxhDYJFhV
HypRnxXizfT0fPH/Ma1es/zSIQXK4iPxTmO2yelthXN7kO2LXSiMkviFzJcnKH0u
9JzV9IahBeiM4k7JbmwhyuzJvRuNP9UlfUnDvMG1hWLJpOs5R350y+nlqu3xPiwS
CDglhq/FiRpmzmS3Ct2BYE08wQP8N6VTlhi1PfFjlDmmt0qr0nqR3ZHsi9PKdvCs
RP/eO1gGTHWpMBXZJculC8/EyVyBzk7aXUyaHFnsrs1Nkhv7c0ZMJbOomvG55Zyt
Ae54kU771gao0btT5VcdUceynkvfr9j0EZqj7CeCsqBAf78s+GYadfuypRgH/R+k
FDrSrkPX+InQ0Sy1nDbuOXwucbEc1WH8wO9BETEdD5VxfFFM54pvnxHdq61IQ7vQ
LdkvqcQXOUG4FAecYKr22tq1xv0vUPr8WiDxjnZjRb5S7VxP5mQe+XBqE2+IdJlT
/vDDWAbP84eHlD/RdS6M54c5AmhsT4H0raNBYypLBu6ib3k60sQa2OE/sLUlYJmQ
6gts0HJWnMmern0sAjCFizk6bQMUUw8OnyaVIy0+G+JvzljZkn3aNxIY4KowKxel
BSXgFFhxJLn3r1DXMod2z4QgnbU7V8JWAv+D9TDUTDvTkTBThGGB8fbEHydpBbY7
XdFhzzeVQTd59eeaRaxFbwZYyhKal26yd23JvLF3zIDHnYaOpYHPmIfHZPR/tQ1B
6yRh4/4Mb5RfTUb9gOJU2gQ1sutKzOrXoDFoGrGsYXEU+ttUTxCITQ1f5GHGsdQy
FfuXXLX6BB+2CPzzvQ46GumBFLImRxykOEUpaXu5e8CYj7nKdZvb4W4bpBMp80ma
aC8pwAvbt3LDvWZoGkQm2l8WeSyH91wEdXiYm18zkxrnzYbiGhLhdrOGPH+/AXaU
Mx4bmmnZb2BtJArCnIWjMYggsmNlmilIArHQnRwylvVxUPPS1YGblBitHj/qXl6C
FIhgdLRFEVjvPrCKuPfOrfTgresFd/5o650Xh+0RIYB1DspJHn1LZx9GzVU93X2u
1S41O3IWBNRiP+lIsUVdSGNg+K3X7gHCDEzWmYfLFBcgRC9jKR1NuBgqvBwgYtoj
xCtJklcGROPMYgowg2aPo2uGsQiKEw36OmYrtMjMDhu0MXJvYs7dTtCu8R3g/dI+
M3tzMuup+2PVXObpNGAtvPyy3tWJRcmH1J1oYahl0ezu+dorHY69C7tW5EaoUXNc
7sjhU2nW7DWHeJGjb9GMsM4Ph8GMo2PP07yhPs90DlnjPtRcbGgo5MgalpsOOop9
6y72xq3jInYig2HxoUjN3/FS2Y4/FPC3amZ+9b6CDf08r34ZPaWo/OT+SNGasvhn
LuNu8TgAGXGX57oVrAjUUcqzDGtxFhJF534SwkWycVgoFbqT7w46uIqM0/DPYrWA
V6U0EtL0FB0W+QKcWIP4uOUHvLHKNsC2Zt/fa1i8zwbY28KyNg88oTB6+dSzb5Rr
IJQhxw1StnRwEPOOHNSgrEDOjmiVqtmjOrdlxbpwO7jj8HOxoZemVnUzUBtCVJ2Q
J7NC0har2uxOjI/ynXnso4yjSXelPs7RkTLMP0hYdGLWVAJGJx+wLzqV9Dwyt8xk
YXQlhHbkrSYI4uLztSDKX4E/5HrFbKfGRjqm25I5rlpFmV0l45Z2usdSq3kCfar6
VpYIjvaSg6XiyNIr64HYbIBrZvujUGzTqsQXitv2cZ+fQfKNIqkOQ6u1hyl2vfrJ
o0zwYihv/9+7DsrbKloJiSzf86gcn0pDiDLSroNpa1SryLc5HuIP6xZE1LEuZsWh
REXya4Z7P/1zc7fXV0pdF0REqCQrDe6gsIUsmMvL6da4BAvPrsg2TeAkvYNVcjHC
dZAOyrVafHCjOHUS8q2LIuZJTJjU69XV7mzvDZIDKhPWH2exbxKoYfk9+fl+eyCP
3/A8xHmWdsZh1P3HHQcKayrdth1GKGK2yFpJsGBJkKNRwMgj5EIzUUoGevNJpDnJ
U4snh0W0JzTXAnwNr6c6ZXd7W3asv2BRdX+0N1VFeRWTrx+7gEU1VWUWRGZaj3Ij
+1OLqKVy3AFgQitTW3RjyphDZ1OO2hHAzaShm+ZpZcYnd3HsldUgOks2NSbnNljY
fIYT3u/zCdDzjk22yeZ+YwV7p3ASJS0sJDtnhEP5PLuoO1YLmQ98uHWCOVnsBgYp
n84GZWuBbYm/VgY8TneT786M1LbpWDxmIc8x/n+Gg8/DTVmo6hPelXtiFFWOHNVR
R2bKlnULdsx1weSjmPkEf5x8pIikw35VmQ7NrtN+ep9+ZgZu4j6zyl49seCNAN2s
qxVjqfI3cnrd6hU4OAmF9GKGvUPjromm7rtZ+PEBKkUtss99adgECz5B/APmgdXx
jQbjGrz6MQRalLKWFiRBuSX1CA/WWc0vwaqdi+yAcmTz5cln9bhgPam08rag+4AY
NorD+QeRT6dRToDkaJlSKu7oj6M4YVKajmS919/7gmo8PHljKjwvlOLr35uhCwbw
OoehksCvzBQ3QQvMTjFD891cH/+advOhCIlLos3mzEpnRsLe3q7Uv2WNaImRpjqi
h4c9I4PyOKfr6GjZz06PWJzYHJ/ZW1IKtsIhTyG0UKQnT60x0vHjMBtzHUNbSYhk
nUZu6q7VzKE33/TCoVctH+ZUY8kIB5v/vONCZOp+wqT8FfQVvb7CdU330ckWZxaS
1ORbMopokHMr4EGvtdFXXzRi+8Y4gUImyQtfusPRc1uBS4x6GsNHkliIITJedFLc
4P3NtR5GyFb8KJ/kM6hWulfOG1Ml5jx7m16EwEmxJkoijbZfL5nl9HejT3fMEr3g
9L1+iKkqOROPyidvwotlcooQKWhQp5uMEHx4q5r3aOS1WB033zqaeKx+nVHqQNG6
KsW0s4a0DMn46xkZgCkTS9+MhIO3AROMLPBeHAw0Wp7nkm4DcesG4XE5mlCTDEaT
NxqRpCvtJOg9XFzyRt1/jwZPyZdJoZDRdSxCsFsxlH/YEjNmPezhW1C9IO94aTfS
c/bqYs8+URm/LAuvAIqf+63Kv4igi/ocAoSMaJ3vSIzGRQG81RIafLODq/LErFC/
CYd6BYmho54tHH49LfCI5HxIZuiEpvg0eEPqMUAMpSI4QsE71nbAZfd7qIIGg16I
vE7S/LP3G1B/GfMWeevkOkNMl0JXIjyCCUZeCm2egsd2RfnUT9+OLG8mFco/MKXU
NeFy5YgjbZyBi6/hkSgW5tbJ59vVFuwgoVkammHq4Pka6qGQuKbpFTP+2LYrk8Q+
ryYs1f3oPf7vyrcNMhW/AxKpmYtTYjXPSu36CkuSO2LkK5rbLpB4HNrt8fn/W0sZ
qQ/orHtZSFdVy92WPtZdf+isa8gLwcj/8X6PtOHRfGX7zJJAhASMHNTeLbenrp8o
StX6S5jjkg22ea+deDQYZzc/fzv8AGXF+RQStbAq8xz3MMg8iIKyfPUizkC5qYao
F/Lb19Umz42bw6st5IyUvEtdc4GqWMhNNGyX+DYz05uRjb4xMF8FNWfWvpWxZDdr
BerT5Wc8c9IoY84MbA6xWMT8HvE17e1j4S3RY9ERqo2EEeg4BnKC4Lvisrx04qap
gQMj8FwYQcaR+O5CyA1g+P0QWGgfVxyx0s3CqjkAbtOV+HsCMtOq/3xRHA/SYefF
75trkqiUJuDwGIYXptmGeLobgpwxbisSUldfLnqPIM0aNl51rncY/IB8nccYEiF8
bb0W474THhRuSVwDzpep0AP/IZhp/Le7nwby9yLCXUSRUS1SF+f+Xgm1tyBSQ0eu
u5RCklg7gm/Wc7QTKI7iIhDmUUvF2UVHRHhJsKqSDm6QsliB7flmm8I7++foKnws
0RbP4WJGVybLvEnacoao5+kAu4ow00lkJmNJ7k8MeQ1C9q1tZPj4VhSRdZ2FGlfV
QGq0CoK2+EexbMwFwZEhwL6h7CU9na70svrxhDXrpmV8F05vjkSEbdYkBw2FD8zO
C7oLylStunJ+JYLGzDLCgfN6fJKge8mUz21oUJqn1MyGb5VjGsY6sYHHil15cM/M
qq0k6kd5iLV9eDoVeHzhf4px9ylWYcatSRdoA2MZBgEhgbvjuT8FkKgrsuQIC3el
QqEgTGJoaVf/h+rfU7B9iSpDczIslt0kkZSFd/8v9657BBcpb8bG6cGpd/e+Y9iH
eAP8lv0ck+9nsiqnOHJ5jcwY412vbgXGcAAPThLETYkqNfnHafvvZxjS6SDzg1zA
T7w3tO02xNlC21MF7nab5ympUS+zbEZqdYTTdvfusKcZNU6VyoWRz7ITEIHD/ZsT
Fd+Vkf2GTazH3Ea0K2ckPtfB4IEQwtIeqN7FZU8QKZm7W4+9/bHSkxk4HHnGJoTX
CGEsxG4wMO587cRoBtJTG33yEeQumH6G8OHjyWOg6ebXT/i8LI0Xf9ngwEE+8ME/
KJzAgaEOQHZCfW7h2ESlOiLcxtjGYMA5rfePWC8zso1z76U5LSWoZ0BIg9U7jCcR
3kyq0rVh4oSsFtcYU5HYAqAiYxjLJgPR/x+OA4ud2fYufWTYqfvnC+ds5Z0cHp5D
yauTEiQEmKn8A6IIYg6zddff/RC/QoLil7ZaAGKPh4+tZEePFTMMH3kVc8OVNn6K
duoH1gSlA+lgJ2hCPpFZuY1frTT1wwfU05iw2zK8p5nEqq2IX08Be73kDqIucv29
a3mg32z4aR3Hc1A1V2AU1AZXw+1orFqYulcj1Oqo3cvaKUgN7twdvMuGsnZhRHlN
dyrAVLyW8mVsoEDmYbLSwRCNWj+JGgLLx+84Je0++uLS18MxVXnw0avedZOJ7FL+
aU6s/fvKFRxVcKlWEgwnNIJJqMU1zHB87v0RX5vk5Ta44BtHOVD0rP+R27FqrduC
uTpSJv3lKYG2yZxEpZC9KJsbtDcfhdLqLgJjdV0oozX8f9ec17+J8ZABugdjgrNn
/61NyKJCP1evksTBhn5Sb8VsR2J6S87o/HiPLfAhJQ5niCb15ZDTt0XKXumkTbN6
QOsqea124Py8eS70E3FxgDta2E1+4PfMbPndnvqgxzstt+XLjuHDGItRHbGtC9zQ
BbCwFjX5sgtg52k5AJl3grFCDKAiwa/6GL0wty8wc1cuIiNQKlx0H3yaFKLhoSqF
p0AJ7uA5VoKcyNQgoISJuEUHp7CrqE5H0RJj/4FrWbLZw/t1c5BSn+8308ZhD9S/
iGr9xtHhWXQPe1AYT9/dEqamjGCfrBZKuoIs7SYXEyRd3FiSx/1ahxxol0HiCreO
fWf/vja+bgAhEnPbE2BepdMH9UUlTyjrHGya6iM7ZJcC2E3JTyJ/zTtMvUG8YwxF
VmrBfsd4ULb5TOfFjptz4SljXp/PK1pAvtYHGowXNeHmFEQM47vPpTCvtxiqWonA
q35HbZmsvRyOA0X/WS1g1Ar869jtBwtzq/yCOywvhwX27N6kL4rm0P6r78COHQut
lnsxFmyaz/zPU+bV842IkxNbc27lLbznWfjLyq3PWD6B1452FL3rprZx5i5x4tyY
xXHik1CNHrAj9ZwSKJnqMIalMNCLt3ezuHM0ZeO9ibW1bVxZN8T98W4+k92nI2wv
FhQECA3x39unHiOOQIEUjd2qZtLus8HJ5oOZll2prlMeDMSgClp1xFtTewBWL9VZ
gEjXWU53hJNnVh/38nKsWNmdQX/Lvc2spGSrWmSN4MqgeJz75OMTAPGZrNz8yDte
VsVFNDkK7L1aR3lB5qHrvSJxL6J8fHVMMgHZntQ2XNhxkPTNJM8lB3QeImGb6xgr
ex0jXmhmaRbVd9ntMm33RkOZ9eLLPgcd32GnkRkTbCAtXpS0ude/MzwwOb+deoxj
PedaJPgR6JYOuBFt2ZaaPLX+RCNydKXGmcUpIhR4xFjFH5BCOEpejj4ykqOPbkOv
oaFVSzbG9v4CZXM0Cd20WFdgkqzYnR5qqvrv81KpH+rr1STYMTShlLsagn43EnJt
fF4CWlIXfi/FY2Mz+Bl4A5opoYGwZcI1mroLzGX6WmqOTP4y0hIUI8nNEvgW/Oso
AVZqbICurq+eYg633V3JWHMZePxSirgIYKors1H60f2IUpT12sjHGAoGx3PKwGjf
5ctQvDAEu4zGiKhwFQi7Xv8YgF08q72DiloYU1Xd/JfiQ/xLFFbn/hw0ku8BL21/
4l5cut3F5gR02msDEtKnrmMLqAx9bEcGmHlYs96a+IrwHIRHyrQ/pxxd5f7S3qnW
2wkYIrVa+h4XbR5smsY3XGDDChlZWZLh/IZd0L3vsI/bxETo7o0uqo+/yD42nkZ6
7knU1U1fwAxJmFeA2M0ZgLFjhVsig1YNgFaRhWknUNoUCVKHFE3H7CEke+fVRXM5
G1yFFV4aT2OjoBu7uPj4zCbrEgESARih5jBHScWqlKVVSBD4BfR78Lm9HVHBmbn3
hfRcQmLg0P4j5CJbMiNZxsvemhGU5MSqfTWYRJOVVazeM3gX8m920hrKLOGSRL5h
PJAwg7tKAh9GM1d+OrFHkScuO38URlDPD8OCGpD30d2RJ5Fuy/SGtLlHQXEfGyuw
gz+Zy1yN8Rfw6YLQK87QU1HF9l2gbzcqfIHJ57uaC4z8m1P/ipo6vksaNYxpidw1
qZkMXpl6pomvrqG+vyavQyYqX3A4QvDODu/oN0LXm+JjK74LCoAjfd2ZGdrbcxiq
oXDj/Fe77EAxTt+B6BY5eTIgJM7nFMijvXybXaGnLlQ+skcJMmR79uKkAht2EC4X
na+0yZk+XYXmouVhIH+KwpBWet+/z0QcbGeJXeyONpTO+U0xXaJNaNZNZsgAsOa3
o+7dTvY2PPiUWIxi8CuhWynrscHhfCMc18INCFSEuQeRpjehpzrG7+SBgW4z3En/
tC3GIcg2KqhQFXNgRgljmZ9xJ73xVF0I+TOTSEPagJZHyAcQmqHBJYQ+2PEmoeWq
MHUuJZX3FiNy57qUbzvbv/2AMiGP3WmYJE99kfPmNbRnU0xVGHAhLagiAwhFdSvo
EofJx6UjN6A87gaFkGOEmcQlznhoOj2DbZtIDV4u02Qo3eCe5DEVScOHUB5Nd9eR
aEtdYDPWkoTjI5aMZsxsY1nWox2bYNvPmaVF7syEFBGe2narEQyR32eAedEUCK9R
wJ8fhZHHaWF1PjOJiFAUeukkLA/pYS3VbTqid811TN9KiMNQNv827dQ12E+CxPYF
lGUa9+WET8qfNNWrA77kWM52A0M7smuuh4FbXTiPLjzSmQsCzgiyWL5EucGrlXlz
azK8LRB0XaIbYpME47POOgpIBZJhXUFAQYMfAFKc4hphWh+T39btihVUoDOdE9o0
DhWs6khjRMK57x45K3EyPA2X4wQlLuu6C6dc8q3sJvXjNitKuiKBPlgt1/f98pVc
nM2ztOQe1momjpk52djNrRL+06ZhOVh+0FdkF5YXpyFPNjC5GdMMZcSOYCIqWX6n
wzLmbQ35rzy/zxnQdAQFFgg4LOPmJpT+xeYYSbqjZJ3bjeLBaEDZhSeXXT0Cz0a7
uCm0mY2rzGrRHHHXX26N/tpMQU+RMmKC/KW388wh8Do1gFiJnT2XLy/BGPx4DbBV
L9nKDLrJ2+Qfr+KQ3WxWSLmH6fXqs2VeduTvpKftk6ELDNzkjlrJUSWLa73JgpRy
xQlIFsUTfLvRLTKwneCfUCwFU0E7KAdbh5BbAWa4fxHPbzzdr/sjlNPjiFA9lMR5
5/Of8SdExRKcu4QOzw8+MbMMV4t2wxN1ZUicc/PVfmE7eVl+TTCh2/OANuWO8vGH
jn27hrD93BVOILxaqc4vWog7OJcNXiJ0rBoPKh8nWQ4BO7FLtJAGmUp+7tTVoH4x
YEvsHA17p8+VGaCpS6gMca2q8DC5vacwxwJWMqCW+QoNUlyKSVpj62LNv5KnImBR
zDxHkJm81BZdODG+3zLbVmaFLcqYNcZ45FyQRlNLxBPaNnzvVPS/SUD168shOPJt
yJubkIN+5MXm8NYgamaSv+ARobboYMHcl8OLzLZc19QvgJyYDZ8fLhSrjGzr5Ke6
WdQlrhaCrTkRLkpBxWVAqBpUIveouGijS5RgMYqRleevY6oLd4MPPfYU6s2Ve87s
PpLJH9qLNqtk/vJVEOW9pj34qD6r72+DL4gXgg08fZ6DgIo02AYG0pSjnkGcjRiW
P7BbIM3vAc1NS5gKRbKCCQxaPL+TYrn136UfdPXYA52Bd2R5ANi6K82P7NhJVEoD
aXvNuGz8eWATnjfJCOtBYkYJDBaymSSTXbWBCTWK78NA9jYLEdhtWzmY9nxJS5tW
si9oDMRbDAA+PCHrlPU5BSuLSJpr+oH/LJorbkmq+HaZK1DuwIi1kzS7DnZaQt14
ZfbYnzkfKRQAG8KEW5rwVhfi3EPtAa5cw0hLvx9WwPz+o9RGXvUAazWN1krMmh1q
Ba6J/E+N32Q3NPFj5WsPWzoda3E83GiAoncK+IWBcJukRm8BhCUvvUCmjrKGgC9j
6BjmC6URbmgAq4bAMb46Yk/S9TuFV6+L9Wkl0ng4GEBelNDTKYpOX2SDIJMqG+gd
vQEMX/23oBB9uh+T/7a3PsbnP5rn/fDJqPcwuwPqyy/QDQptLjwYiX32H1fGYbIz
/chKRXqtQPYRobdz9goAODh+YKdJYTJMyDBZR6jqjm+/leIuo+BiM7+ER8bmq06m
UBcFPHAVl+IHcyHnE1KSdW8LuMT19n6eLWq9oTzS2WYwWGt1QxMvD4frmPQTpTBy
kAehxclrXltGCfGDH0Rn5iQqt2ltp52y8eTk+gd6WAln+GTZhNGZBuvEC/UbbZNU
7bbr0DCIB1OmioWrm7Q8r7ShG9Su+L+vpO75qENMyDav/RBinUuSpdtVxDLpytsU
qvLZwC8UYEqURlJNwMv3Ow4+oPIjOzl0Gnb9O0Ii8myizrvSSRBI3PqvaKykp/Om
Vm6ffr2DNZB3PeefgmcfzF9qMDFQfpFff6vwXc5VZlZRXjcFJcvEhSLrDr7SOLUg
+9uARZnib2LSdjFATwa+zo3km0as60/UGTRFYzvtvRZfpFIdLet4bkv1tI/YlhOY
N4k6/kzj2fbDWFfH9QDHYSCDCvpLbEos/UA3MuYwyo3ST3OlBe9/aAgRpCNiv1yJ
OaGSz0685+2G0mAs57fj6f60ZCCofXPoUw0pAMB3tVhNTvWacQk5lcVIn45GqP7G
JGPAkR7t9XdAzN4qJKn/vdmrJeVP/u806M3TKJHcpC5SefqKIbIP73NT5wICbpoG
LYoS4B0GS5pRxizKQ3n+ZB9BBnBNi9KuivAyHSC3S2lu3RHbweD6oigfZChgPub6
kb8r5qJAF9+cU9vJDeujHXCXW2C2JqHAS8hlEVQNSNONArn+uCIwrehkMDtxKyLz
mTm4c4IwpJq8fmhxFMWkbUR9eYHqYU4q+wi6G5D3+mXuMwKrgGfYWKEIIPVUykzu
Jcw2NZuRwi0N2IhBmW5sD34SL6m3QslMjqLaTbR5u0CZ2wBCmqQFdPsjNVTdZWty
Y73Tk717VLdyGb0gXmjGslNjCdpF2vDrwEfLlLN0xpNzmVRuekWQMEbiIogE6mQG
V8yk9WnBEDp2sPlF3rcn8ucZtfhifdU3BdDBj6ux6pJHr9sJW9Q0+CQKxPjtdXvZ
Y6V5baZnXpYl4scKKYEbsoqQdR7DNwjATRg5yvQbZg7TvNZYPRIgyS/P+rR7bBco
G56fYTQgYrJAEMtZJP1CvgpjsAwjfeJ5Sg2Sc8jqd+IC017VK1bt3WVdWWamTWQY
AyaoouqziWixXFjwS0C781/DRGlnbe0JALdHOlhtDwgIlLw5b+1icYyMYGMLcUvk
DA+bCFZ/VuBhw5uM3FinyZ4q9bvir+7+03dXx+ju2qcIYb10I07ctlSnE8V/qmkD
UI7jLq9QVU/jSjnaMHxRUfkRFAAHYlnahTnEkRaGZhBj43bpEz8NbcuZsh+r2n+9
B42BZUb7D2UN/ytaKqv8+YnI5gFttIhydpnvbRSyxG11sqcMdv+JcQb2szri93PD
/S2RUaB2jkYHJQIVUhsaW1R5k2RiLVHh/sA7PumSSjmKIq2cpoWUR8Fy1xUKXoi3
dtlpeDza2QpjaXqWxUlJ0U1jkDPtCsQx6tSk2nrnvp60rg/zPfpLjtDbeW+lRGeQ
iG5+mc4JwTNFCcD7E/gsMufUNmF0aQSdZJKVyF0m4iaIFlIzgw06H7b7Heae3QIu
5tE8L8XSQWkya/YV2kWz5BepYnrpEy3mS74m5KB7TXx1efpsTxqJgEVFhzH9zzWX
YKu8tn3muGQp6ex7t6eBdBpGWw+B22Orfk+RlhrwjSVdfqaGUgm8pMI1rPjLKFed
HZap/r16w36mTXM8xQOFWPuqrinRQa7eo5iEVaZKz8kzctTQs9tT/vMxjAKhFw3I
KN5B244vqMUB8+BBtL9VOqbBO58vzwNg1tNGoF6uVU2+iwYTSr3jv0Ktc19XcJ/R
XNjgJSwLAI9A1XeXxXkpN/KIzxN9e8wqa/K950pRwI8GOBOpMOgmpHq7LKaRGGhG
2A1nZFcyIpusdtT78vQhwO6KjkAsnIeG1wiLWZw2IQJJrjZpm0WumqEB7jYd9oKJ
fU1rb4NaamnwZwlrF02LW8xHDO42fU5XsTK2tPXtjohVdGz5xunZ5kjGt/acsOHa
19iJOezwDE8hTMi/sM+cJZZ5P/ObSEMxxb0ar18G0cmDTLzAEeSpFq1X2IYRsG38
O6vTqc3b0Raauxltlf+kaSiXB0YNSy6EOHDqctmwmhF19jP61NfHBOYAIzyU5wg/
ZIzdp629RQ6sRTtIX+0tfX24I0/UXWSXtGD+yrv8+dQUjokgq5scfL7XhObhaGzP
jbmE0mDzMXypCmM1igA9qNTyW/9GodlRq+QLHV7z7ySvjVIQLsG99lnz+Jt7aO65
S44uBiDl1LCwwhX0nUigL6a/2wEI7XuJlIyqzOJakzerMN507r4Qf31p8QANiz17
mGDDAspYOPEbbVGlvbIyOdyIS7oelOk2WyDrqFZn5AxW1im+hOF3YFgnA11gG6hr
Y6qwzLATN+U+TWxWPSe13ZJEfefC3UZ/9xD4p2CNT8yEzx9FYW8zDxuEq2My/zbu
rkoGJl+W7OTcIsL24I/rJG6TD78cYbGhlKVHS2QRxVeyJHzYE79oxQ891dzRlJfl
5JI3nq/B27tcaueUuBl3Nu0XdPm2ill3uxLTl9n34M9fkizkBaj/NXc60Ssmx15r
F7RKwB0V8UoAlmJ5+7y/FQGB5KD+gJPKoOpxdxYqyt7OrI43koc/uKIhhDms9mWb
AMSxwR+XHOd0k5UmnFdRKRNsQhUpLm7uQTKJhcjwromzOzxPzzN4J6qby8gLBJP1
BRD30/b+zGtw9rQoOV3BxUyDOyid+RVhNVDVseOTQzLX6YEwjm5J8WF7/1cUXU6e
vfxc1HqzrYMl56LfQ/1zRzaFed1IqI5LkunMSzU5oNagU9W7D9h4cHh/2nY9qLL1
836RQ1sgu1EXjWIbDNba3ciRs7IklD0brYBwG5fTTffbJd5mPsYMehWHZ1QWJm30
H4aqaTAz3j60H/SDMfDZkHAJHnwDTTyryniUvzS/EH999edNXBtA8u5SZi0uoJXA
n079m/YEQYFUDPKvR71N8zeD+v+ABWvkvi089GdlI/zn6chysj3wvzvGipaL7g3H
qgakxEmxNcnHwTbeKA9kKfLe4Z9DdPEnJx9cKVS9tOETz/sWnx5lKEwYInWylH6N
gyk/nHa+u9KkV3MZ74IhEPYsUtKLcn5qqqFJ5xZUoO+T9uwQ6tXBHPc8BHfpmQ2S
f/oIQlL9Xuls7BILjI8M3HnyQgy9ELHmlV0Zv9kCkOkUwpYrTMPostR0DwyOz3Op
jx6ZVf2XPOJE4ZnkSDfucU2WMXGnYL7fviCGdfayeCPEx5ZrA6FaKt8piMrdOFUU
gORCBlENTvI2kYHiKYTK/2QIBg+36IJ4Zj06gimXwi9gwPGh3I8JIMwMUaitIoXi
Rsh6F+06ScjbCcam2zEdkZJ/BIHPGlKPVTGFqE/oWTMv0x2k3g2NSzWJEOovomK8
JH1Tbggl78aMMTJ98ZuiFNg3+TVavEMWpU9CcHJcsk5e5Hu+GlQJlYjRfzdfAJtP
m7vvTZInwGdiM1eWixQ2LTdNsWqxNU3T1msJh4E6lNfGymbFyM/TaIzpnOWQpKc4
agc6pSFMxFPIX+UsZyDh86dOaUwPE7vZShbsTQQn3Y6yYTlSG3f67UkcLQ087WtC
35kP7q1pcGe+0DlE8VSVizWSN3GtIaBzjw97DxTmjkbd++dnC4/CHQLZe/ND/ZCv
v6tJ1reN5ozjm4duQ9iX9kP082KurBFGt6fNfSZcmN9qjJFC7RBE0vsrZkz3aqJR
ixbWrbOENRZMNAbEY6osSbJP0Hce9CD61HdzlIvzBcpVHyjRUYckxSi1bsZPNoDg
DaD/jEXTq11EXsL6jLovIF5M0GLs1gBZo7O5KBzOvSQyNNwAsGXwdc+dazqKXMYl
bDPnrGqURcjoa9qzIS4bzD7u3D7BOcVVx+4TxWgKncwaQFOojtdMjtCly3nWcuYs
7DFmbzPlpHVcBaMkhf9d4/yACRSxHb28hGtEAyLyahMltLDDzaOlIYX9/TygxJTe
/zPQ5lwsKCl67aLGbQ2gFj+b4vf3FvVqK6OtMn7q8jTylCDk8pUPCFBVEJP1iG71
qpoFtLuyEb0FUkNfGjq2FJX7vLs4b0yEM4cgai2mGRnN3uFSitNG8AMQRehqyt+u
DjR7e9bfogumFP4PlkYFo8FY7PieL60uf3VJllzUUf8RhkPu1iYjBbAMkgG/w5eM
TZrt0BMaEwspUVQGtEhEmmy4vAu3fgxWAIuWT6N55ge6mveC3O9/dv0XmcRXrxg9
1WdWkunwdA9rGzYpDYSmXPe4hW1+Pz5pFMJRpVAzilS+4rylc+5g0La6Hn8vD4W7
DXUsbLNBAxHjEJYp/AvFtOQ96DZdYLW2VTdXyVDuw6vnvHmSidBISp8rM7P1HUfo
1EL0jXtRx+i7cUecLOGPEfZYDKkONFlIcW6V6GEFTjX+ANyj8WGm/GTBSdPCCifL
NgQ+V1YJisM+vcPWlrUDN+4jd5/JD6NenOL74DARnzG6EFnI1/xrxuWfd9fRwXNu
pFezHbtZRXL0ZrYB/DQ8DWek5U5EynQk9f/C70gRDpBwesTHK7RzFnbBzEdDT9Ja
5i4vqUqvhw7cvn3yElHLNDzm4O9xodTKCnbFNXtnJEDy0xzF2DsK/XxrMu3aOlA8
4jSyQW41GBEX4T40Ud3eIvEHP0dauYpCZHGIMU4snbr8w+sKrZoCjI3Vgc1lwKE9
p/noxqBFZiGE2a9YjkSfOu3WXXO0h02PbdTcDnLdGm3kBpuDodcNh2Mc0NiE5m62
DAxjzTBBJVZ9P7HKaKO5O8ppuQP4oUOhgZ4y3YAZYdJg3Dboe2K5rSJYVzn+nQDs
mUcezaOOBG72wsuN955FVMWtvioaB4vlW7uXI1nKfKxuILadmVq9Btzb7QFDD30+
il4DQoEVW0kLRkN8NLsWP6fR6vrFlcYcgI6dHSqwF+pUWMNn3izp9MCkFZeIZ8Z/
G711C2xMd9MAVHCcFQRElUIvyq7P4+CLFoCiuRWz54iMQpbPxpdaAoixO/0XTiKu
IajITpp+K+n+vl7prNduJCY/HfwZGee49bK7VUozo4r4GcYy11WhAl9RhkU0Stm3
BFShVn1fkufpGCyQTCQfZM6KFdg5OqlAHRjqBogq2gNP2TrwCOKc1jLfNYN8f1tD
m34nU0s2f8JjsDEgDDEFknhBF7M1PMwm7AGeU68zsoD+IN13S98+NKrHJOFNm+jq
IBEqJ6At47s+Pr1ayfcTneEkJuXRWJKqMqUGC1XSg2TvQseNWucwDsfjWmIJPJ74
TZ2oNGOh9luajFHQ5N2OlYw2LJqTAZtqDN6xU4E/xApnVxQEfRNhPVJinkaRV3dn
8SF+4tNOKIZJeNh4QCvWByCjCr86BH+6U5OK8vE2L7Ws26TCQos3PEniRSc0hCNw
C7A4DeaW0cQw+nUch/y2PkK5grwCXZHiOEsCt9D4Al8ZaowzK98zCOH9V6IiZwhN
ylF8ozyjg9P6v5fBLO0MjCf+QueQxIYmxBwJ/QBtKkxwSMiXWXxjEFWEpapOnw3d
w75/j0jmalpUws//0tZEGfwa9CSAMd+a4u52VHJnoyfOKS07ylQLCBYPEVA/3XrO
nHGwOE1DG6OnvMoDy1s7yE0AQ0l2ixdgOHr4EIg7WvDEk2qdnC/F41jtjU42iwm5
J5msOS4hRMt4xncWMc1U2SckakIjlGeckmLBN8V5gd9Dcqk3o3bIFRbAsGXmincg
Do2x+O4xtd5m4H1e4xzIcXFFO3cSF31sjVgkIWpsYOO11Etl6osvS6MVOE8+N8VD
G6iBK8K6SM40GPKzGuENg99R4UsUS3N46KEbXHjO8TNvLKKaP0G8nkbHBV6C18d3
Y54ruGFAKaLGzfGA/PwuyIL8wbqZ65nceWKDIGaVNqCNeHaOzyvcbBy7uESsmOLD
KcH12kRWWP50Ynnd1K2XWAM8vsqrLvJLNq+ERFkm9FU7azq93B0nIwndRk2HCkNY
VrLguTxcJubgm1Pb1388jCOj7L1vk/o5ocs1Trv7QveHtfHokDGSMAlyvL+GF84F
xLh8tR32aIopxTFs/aqqrb1itJHnE5P4row2sIvbb3o439KP2dD2452DNox8srwD
Y+xBXPmKDP2SESWnJKWmWyzBnw8epzbbdtOf1RXcR3hpCnBte8vr8HngsDwo67Su
gTN73CsVHsuz+bKAzk7CK4KnHQ/aPhLEIRGRBGpVj+LqAFxflcJV1+KyRsqLnhMw
AQ5WgpGJYWu7xZ8Y+eCGGVVmO+0gS/MNldEF4PeN3EZyCA/5PRDJRLnFvffOtJRf
JcOW1/xLd66+35MHwnQ+dzKQ0lvbMeCb0VgioPa2OJNZgQff8gfcNjd+Gh8N/Qyw
kaCNAczpoSeEmQDfzkhV3uEe9UNyj0YPavyVaajYMbLUcJYHuan6Pze75s/xXfcg
pNqINnbs53bX57U8nnJLOWNvaUHPC2sHsA25NESnAma1GRHYNFJL8AdFXsGsNCop
n/MY2FQdtxQmswc1z5N+ci2UJcT1rJ0uwzksUfVlbbTWU0EsKNX7p1URoaftD34S
yELIGmvc3vFZqZT3mg98NeArLapUf4pZA8zv2Zwq6deNS4K9y0px9/oMwOZBukQD
7kGJBg9djQeGOqiO9ew8yL+Ztf0NH0Mq3WHH/FJRxHajtIcuchhhH05bkOBzeeq8
uKh46HnwdbWRGadrJiw0MAJly1zk7x3sQXsPzEsBQFHAiEMH2TyUoj7jG2I1cKMF
HGuu2eavl3eF/ozPYSNSXmzT/q8qOpdAEHprMscD22DFylFVzhNy6kE6Xq6YNLY7
i9g0Ue5oEswJid/RFJ8IvHDn7yrUd4GM5TS9VXTsITEXEm4DccB3aaW1/ZK05cwO
ej4Gsqw0iCocXqqJYRuDhCO/RJhVzIHL3vNYhC3z1tebbHxonlHvnzPbnhbezWul
QxieNe4aDYJ+UkiQSJbStEW4MHUsTkWX+8oxbC+/ISGps/GUg3yGB/tdVyLJWyBw
D7dCdn6ZegGTM5qTf/ZOq7g7lMm5krlZtF28FDjX3Udds/91RvYMzwn3HmagUXIA
Ul3zH7TNAuHfGtmpEKi2XQyFiKzSaNoT8XDde5VFofQ3GNAl3ZZQ8ggFTcYXma3e
bWhre059wQrxsors2nAT9soi3WD3MF6bBleynNSlM7vMHNqs3ReHzqzdO7UzCqlP
T5gg6Zo1z/Wl0yMYIattvXknTY43S0MsojguHq5VruzerbUBhCyR2mmEAh6AjZXb
K3sPBp+o+AtEl4siOplbwxeoJXY1ajZCukMP3n7AnzyeLOth5Zqfm9OMA+p7v8Kp
FpJNQHKz9/zB6sFzvnc9ygux/gREcz29P1zOOrWIZryGAWeIIFvjuSGUhu8842bu
NhpK9QS4eZ7Z7IW3Uvrr4/PT+Nl59ykmanzBoL9yMPIjDQHfiQCrFRS0rk1m9BIx
I8WXn6891wBYAmr6TnDAgIOe8jaVoIXRkKJFBMSS3ca8B+Kvm8eoTlBw2q7v8FYt
JwF5tXuEYkbo4QusyxtEZBM6rOqm+AcHOkKkoEO45xt+gla91U0JdW7E3kx4afgy
KpYHPyYvdwWzQdycXXYOp2rY2WYIHuBI4EfTOx3gYqSLo1XSQrAdiSMvmcx0QWaG
NrQyey6KuYBywUsf+BNw47tYe0a8MSpELZvD6adThAx80wLFvQxcKmGJmwRQVEOh
kl42E2onxgYoszJmmFh67ppclzjLQIRfPfkzUz50kanprL/p1uC3DcYGE2URibh9
o22DlbIJuLDS6lIBL3p/dywbowjKfqilGzTTtooi1iXF5axPpNNDSXgXCFuF0o1w
NFV3mxtyKpj4k+D9hlnvG7pRkZCl/zP790G78lESKvv+zT35zgsxqvI452u7vQU7
FQBaXLH6qbQssGg47b7KCf2S9L7TJcrEozBr1oLN8Dqz9GUZZc9sVseA3kUlxT6G
0yG8E3WXL7Lu6sKPlo+Wsx2SDoXJeEYMd1LXXgz4ormNaeMjKbub4gRCSNnaZNUZ
K1ynyYFGgTURldMLXnto8EcU4CHNK/sf2iMQW+nejdznmaOZ4Gas+6f07mjOvGDP
LvKjzLgzBpJMe4NkhMkB8sfbedn/DSgQbXNVcg3V3KAo3ARyoAhErMDVFYtkHESy
nP0J85j1jQxaaR9hqLNZR4CBLy8PguM7StlAFuiXohIAK9S1YgNmpprrYggVENzh
FYpShgGnbLytU7GLxobt8YSFgLuHxvJcmRUfKJ+UKtpEI5B3iKF4O/9Cid1SdHr/
5REKALqM1bjAyc/EQxZcJc33trlPTnnKkquy4JhhKUcuey98p7cPPkvOTDSKl85l
2w5xKGXXgfSt8wKpbyPv6L17eGtFjTRhWtfdSwPoy9IrESbsu6WZ00ih94nFAqJH
TY/aEZiYWfChGxCUfgZEs3eJ5wk8IwgssS8A8WB33tivPXAmdHkOX/v9R2qARsGL
GHTsxIC218qEuni0GsS6ANwmoOhk0/iHjAHgfqpnqXeSNYYwxD/ezDOoT7tBmZde
8Rh9odSmkIGiEIXUow7JdmZaRUz4tHPMkJehgpJIWa2QvVV9hJLIsTuRlxPHIbS3
MPqMHSfbHsAIjxOnChP8mhZIq8YeYc0/NJggSekt166gcQCvazwU8bBlsXpv3OfO
fDnMpwJSonkBwmkQhRCp5IjNeWdoGsGlcYpQ/dfhiSD13z1I+jK+h170yCWNKFWp
e0FhdTFDLShKbjyI4Kgn2NR1FjyqD1cTNhRxGY+i34cFEh90phZ8Uwr43UamzLQ7
p0+aDd5J1TL9ont2ULMWf4D6uMceoPacA/bbhGbMUcv9vDqFyEtjQoKZLnLuE3Oo
hwX5Xz6V+PsG7A0hxyTqyMDtBp8COUwG8RmUtcgYUGi/ojU9r/Y7Z/2t6ED/wV5L
+xavFE+1L3Z7HUxlC6bKhFcbF9SKizkHYy1OApGJjbGM7Iza2YkqrUauJ3r94gw8
5CEu8hXBeRVAFKZbo9lIWGCPfn0m8hJYpXqbV7ivJAokpEVo/zbN0bTmQlUQ44Kc
lwXfHVNryjtHDY8178+kqg1Q6xqa0dAmFPB0FfJaA11RrD/HelvUNdzkvtJSiWOb
rmNTJ4LtUvH9y0iEi1zn5r+buahb/W5EtLypUFyZA+r2l4aECarWZbShqwZekM9f
RkB90ihvWSJ7Lhx1r+BZ8hi/iXJR/psmPcTwcm/7KEvcRpY/uxnnyAgywFrTK0Zl
MwJItaMhsUXkGJJ0aAWA7DHw+/sYKgUar7yVQhJOfex6VWYjR8sCa+RnWlF58VXK
UPjEDOCsPl6pNg9zGbLbDOonfgPs7Va/WkhMwkSTv3mkHbVEkKOgpRLcP26Cvuty
DyI+Z9ifhFG/q0yN/3PsHAEbVPsEmidIz3Yse5VY5Lx1ddBFsVMSToi+/htG0J8o
Yi12EyRIZFxd6NX3fDJycQvcw1urRT40uhfa/hpiFwkE85fgMAcxaSm6imHV0hwV
RWA8jCaK4Tmw0OWsKyBpvJcUBpaIGOS/VpeOn9mre6rvdvSTor0a4LORNAESg9Tv
jyt1dpzHlLRRGn/lBuWJHHFvbadkOAQiLfCEaVt+bu4MgvX7gZv5TUzKzfn/nPNb
8QdncxuL3iCWkbQHePQES9HS5AAI6hK+WQdrQNnOVumyq0GaklE6j+njtNfBGBId
ExOJJgxTKbqM+IwWqDILYt7y3Fbk+onyJ2F3oF+/HEZ2MGRjhRW9PRgnx7cnz9s5
ol1BZjEDmZgOeL/xYAowNwf7vQ0gAc8Ym5l4msRuhm4/HbDfUhkPQ9ZB4eOFyn/b
5q+s3U7eVDyzKkRFzjefoTvZHY2Gjvex3tTDFtoV0m20HinAj93Wg9CKCaHpKJU9
2jU3fbe4QRZA/2tBSxQuMnelp3gT6AjpwAJTCaQg/aPNAQ6Qn27BsCZp45n0i4Hi
/bMDXg+Bw49q7hPwEZ8VhEs5S+9VoYokgqLWQpVetAJNI20WIqSY0vIQRoHlcOUO
F0O90fVQv00qEe6GgB53WsSbh/ADaWUc9Q9fIlPuMsxXTXjj3qHj1XwGzxDbsPTJ
6Eo2GUjvS/Rdc4Xf70wH+/H/qsulqfyk8T/kGjugzFUudPk5TpYVnL8D+v/pWXCb
cCj55OpCwZ8+KDlb/UqQKNrQDmCIA/H8CVCrsChm/exicZwK4xRcW4QzyQ/awHQN
xV0IpJHLjRVaigsz6cQeEXYeiJEFDxvhPMPYDyz8TrLoBccK2qR3D0hHG0bV7dzv
K9g+nGYW2hSlM5qYAUp142rd53vcphpqkSklfeQskV2Nwk/wPP5W5nPEW7kJdl2u
KP51Mmtn5gshjKAeW4K/J10SGNQkQDwADIuXWDMHxUm7OYOKUdUl4WoroWxXs8xi
W/nGeh+0s01WTSL4Oc6LYKwEJGuTY1sLAOpBf+5b4TLJZ0hcIzZuXIC8DXgRk/qx
b8vb4OK4djjHpdKe18Ay2W+J1VY5OAX63SCryrjKKY2jJtpjgoRTAy/XWjDAL5wL
4GgiXkibCcm8ILRZzN5PJV8N9DhO7zJR7RewGz5RPqkVtaaQxyjpVaW/G5cwehCx
2St9IUEhKackbMF0lRMxtxz0oerBLHQMK2I8dQlu/5MFfKj9GPsSq+EOY2dTV1+0
9fEV8e3YbhL3skGXIxa7EzItjy0HP7Zyc4UmRRp1T4058K8jWBsWeQ60wYo6FOXt
LubT5wnfUDLnxZGSVI2sF8gAH2LhKaBLEw9ulxHtg/ddEK7cFPZKZEvaxKv0UBVM
q6PZaQf7NMpyVndGApn5yiiWjVZFTweks4QbIaL8KTrhe9rU9qDlyqbTYc4pOazp
2ciohIpYFTHv97eFLxqZ42CsnEI96A6hkg6ufLmDPZg+aL788tDl2+qHF7huajWR
eKiAFj8IhVRYtg9bL/tEi+vQmYDphKas0JZCoz6doh8nYCmmVjjjvsEfYNSuORJP
AnLavKQvXmxZYMcMCc3v+jpqjnqEZmHaIHoaeavXfg+JlnyM7bQv6eJ2LBzvTKfd
GErexC1Hn8UBlo3RwvvLFejLXgv52XpCVvuOp4z+txJf1goVFzQ1fM3Bu8wuHRzC
UkVV71hoX+h2ahx2HHDYDDwQUqoK9+zY2o4dmd33ywdLn2RmS+EpCmqDKLU/e+6B
VkyKUUBjJoLDq1B5WSXV1TZBBOenP6yw2Jf+zRF4wE0XZLNDdAlQg5ph5ITsGUWT
ryZaxgVN1GPd6pDGQQvrNIgzXIC6212FzOFEh8TvxBfEJIdq+2SBQeEZxvi7dQIo
dpa4pJ4UG8Crap9k06ewfXDUxUWg9yA8nnZComLoWz/pkJW2QkSWPKC7js3wsGrj
31qRs+o2rF9b5JeOpAcQ3rRqQ0GZ2Ew/cxaxXA3Wa5NZjXgvtumkKgtI0OPw0YdU
IHD0ny3je2iihXD6slcqweFc+yZRpR9TYAUTkNpl/p8V6uSQvn+oqhnL8TXpe+Kg
NkQEErG0+MrZmIczrQIWW2uuWG8C7gS1xq0I6q512L8PBqO0/p+VlVPkiSKn8CHj
+XMhcyF7DZtb5VQsfHVaC41CICTd5TPZac1MaIhxNjX4U/KvpwU00obmn1Hjbefl
BK3D4brWeYAC3WYKMkMJoSJ+YStZfFThn/6n3f29j3iJDHjclkvr9r+qB+Dair5S
ea1J3wmiVCcrFydUTwklI6+h49oEjhLU7atp9vfT7Q4l2gsTlceD/E9NZ7Bo2Ejf
Dpa5O9YyCAjc/UeOYWnMWCKVllHs0a6OghRMRACBh8fTW5FxvPXbmLSV7ii6suWR
wxtDXuKoh3VPOdgurRdKMVphaqFFyZtSWA736F9SIseU9rj7CvXzz9zcOqw+KhjM
J2e0D7+NkPc+8eZWAEIqSrpX4d25t2IYbHjQCKjhWHePWJacQAo+YhOU1R7PjTFV
B/SoFDohQJHmqkrpnWrl/Z0zZtqMm7+RRhJ8ykGD/Z8OKSNcKrtJAB10a78PEINN
dVV2rS1znWw8CJgLi1B7aDKXQJq0dFIAAHatK98x/Qltm1Lx2K5Tj2xX+JiB8v3Z
D+GvujnuTAnGtC9zcqtzWnxmzvCJ1rVkRnDUXooyj//sKEA6VTyxTir6/4XLtKMz
0tLVFj0R4NM4ks2HN5X5+T1GxQw+Q0yhPqzHOHnZS23oyfS21Dpgez3jQVx231of
QtcIJK3tgQXfh2acchPgTCLfh34hHOAc1J8Rs1+CpEuwYhuavMQ6bmyInkKoewlL
Po4npp7exzkKciOW3sUdNevkA14XA0EaKVZ6CFxrfXjmegFQ3FzUvvxMAPBdmf01
17duxg06+Qrt1AVkKCVP56UClwiq2lvz7i89FTDc+FU1oRlNDh+yMLSD8HHKPVBT
CX79xOWsmE/QgceFM3HB3B3Y6wDzdDREvAifWjpaDHMblqubY8YLL75midvhkrQ2
e/aI4hSwRUPYMM0h4k/npFUL2CuhG4uiTpmR7VcZ9b2up0Pw6ixSrHeAC+9h0fly
i0kv0tAfesokgC/KaJYurGP/HTXJyXLeUoAvQYCcvltbz06U2e/BTbnDUBdcA8U1
L5KylhCux5tGMj+zRtBXQJWvqfpnZWsjrPxjfsPGaiAC4CSbZxb9bnrJ1+d9rDZB
F6PbCLtEbYQof7PaBPc9w1xlfJ4lLl26Wk+XfCc27Acdd+Rzet2fr7Pa+GIc5GNL
fw5V5Tp8Nfw42DYHtIm5hoQy0VxGuxCUMEfgEvn8+nGJ3BAffGAtJPKtV8LztwAs
GZuLG302xuhN3swxAbillj4imabMhvj1bij4LPFllqtz1BNf3/2xBjurHx8Tt+2h
YJJDyYE+i8T2uhc/W6AHE6t0g49QEI1xl7wwVveZjYFy46jk0dG4XsHuOkG6EdNW
nz7hLrDQxAt3mqMK7GA8Mt7bxfB0rmoiI7ImSBXp9aMiicDJILpWBBQ8YYM/KzXB
0HAIFL4oGgblOxTVkmY6zhvbC43MKeWFXPrjkHHL2OHWCJalkKdu6wP5+jBCv/8l
9PYaTkDrHM35YYCPDG3WIVSFC01HorYaFI6tb6yQIvdajCi6DtHiGcGVGqxRUCXe
I0fxMAU5sT1jLmcH14U5H0QZzKUpoLkoU04Lqd3BsEubQhRUPnzHresNvSJnhl9V
zixKs1qX3iZFcMiWMwSSH2tHV4/XZVikpwMQtjxhzW2+EPg6xCELeRcwuN+kE9P0
h8eluUwg4vBwImvwbRbk0mIszp/7ectLBCqSWAaJ/QRBBFJ8A7TELyfv8Zwgg4gG
7wmzZa/zoJ7OQixCLLIvG7ydNpO2UHHaasNJ8LlTcRmWuNrhxQfiiOq+biioUOIB
erIyikRaxy469DRbi9UhoJt4Q0iYcu7KGd0B+F0/0r5siZAOWOmUF7jbVD1G1EQZ
3XriOapTUUoPZG8LebzDaXKR+JY3kS30LssXihCfoCTDYZxsHJUQy8vbAIwBBO4b
ajiXN2SS5b1LcqLQSPuTYBQojL628EN8IE1GDMlc0w9AeiG50hiTTzNZP3dN1Sj0
MYPBaO2vdNguiaJ3ckZd3bz58ERtp+kge9Mndbae/GE7wPgGha8z4wP07jHiMlCA
yVmHsH7EXZNj8H2OglAARhmrWcqjNseWcQfft7K3JO2aLsbstduRplfa/U5bxNNH
pC0sjhS4Wb28qUOLC9DkNZ8iNBtV4Dg1fs8d/q9hz8wc+OR3ZXQ0jUkSjP9LwyZX
ScWgey7PGzJGWUgxeIbJe+vEJ5MCWt8obhFNdMpOULK9e47GZGCeETYff+HMaovc
1dFH/D5EOJP4q/sN9DrKyxYSPRjGLjvGvnXarL3LwPFVQmhh3kQF8X5pexSzVcCF
3wHPzquTusFcgbQNspBO2fkLpWnPfeZwk5NQjD1VZRGQaSghcu8RZkWi3t/OsR3v
sEHNr11h+PTIWCSFWqQUZpd0l4/b1F9UBKf4h4Gyx7dbSInBh+y5a3XhMhhCf6PS
Ap3kLJfA9dppA17yn/htU59BVdHaFApdsYXExQtEi2gll3mvn7rxACQMOAyyhsZJ
UeUy6dN1xxZU+Hxnji4SmbmE623IbvPBMDIWz3Ny0erl3ggfhKlkVXo7pzE86Iaq
+Gesl3qqsjEZEwVNA5vLG3MoEdYxu0c1eihxe0NcjvjyZhjyokoquwakDaOW7Oy9
9whFmbt9IeB1p10jaioIAFbiJUuP78HBKbSgobXFzDBfKXTr/RCahm7sMvmb6rG4
CLpAlfY5UJkK3y02Er39Wpn2wYIYzPVGLiuiwFH90JKv4pCUEluGyoUnQxrIbl2f
uQXU8e6nAu1KEJ1P4BtLmj1UY8NTJlnPnptoUoYrtKseLW0K9efQD3GJnTVNCASW
tfEQL9wyfpRlb/PThq4dttP6S5maXpdZjsLITy7IlxJoVDR9GPNOcSPIXvVhC1c2
FmBQzeaGtVeypXePM9EI8Y39PsdFphjLeCYVy1Xct9Z+asQ+qzqTRMlpG1b5dvaR
97EhB5t3WKVzXnKsZImjENMS72qmEzzxFMvw2u6JKlIwMWgd7tlneIPLvPyzqyWC
rtf+x/65ePelMLXGJW93zXGLx2AK+c6V1DIu8gL6fT7canWdAEiYwxhq28hGdHz6
ISZfyMwV/nXbtAgv/bbtLOgIo0smfD5HBpMLdoIUgfUlrEf3oQYSAEYnJ5d9++eS
Nx4Me2VITVBHcYjdCSYBQc/ZOLwpY9qsePXSq8D5/vTcrXgdQ3Km4CCI/wpy6OQA
3i27hdu/7V5Qy7u4OtiyVx1Ql0ZTOjW1MX9z4tuKVzFnczXZguRy/mQtNxEBRu6L
hNhd0BGqMW3E/YWE4NfyP4ddlH5VMxv9L0v1GHqhp35LvmvEwlkV8sP5ZIH1aS8S
k7WsCnEWFGHqPZ9OlVxU+ze2QZxpGDkXCLN7UQr+OqAKr4klZ/wj4+xjQBxmz0Cs
FAAIto5MXjV+l6wm2UIaIE9EjFPATcjQy5dvuNaaIxYVhJew92eXJSmPRnyW5g8c
wqdjndGucBQWtRhv8sd4bQcYu+ZckBicTcrWXuhhOlnQBdJtowao+DySl9lMXFBb
CjmtSRwgdYV0q1EsPJRj8/G2nUVlhOlbLhy0CKLfo/ZmOshCVrdoH9Zrn9Z9dfQM
MjM/OwpqJEHAnoLox8X1m9Gay4ngQ7T9VeCBKUHi43RlQlScA79YCuFyXQr2Yws8
8YnNQ7fUAlg9hP1qEqoSAqMxGlrCk5Fcziv/5QEHyiWhbzznkwMflLsrk6P9gadN
yhARjRxNbXtGsfD4P+mTjXJWUutV7AsReE78fj6qX+wr5swhMFA00Mt8wfkx9F4z
FAgUbVHwjinqJFAoSsm7NagULC14e4lapKII/4rN8+oaNTwwbl26uSaLLctugFWO
8T6FFsQ0w9drPSyxIoUSU8bHB71gavaG4BPpnGTP3mhqOQFrBPl79UpkEanhpPzN
1Z3CYUjIVJY5PM9cnTqj+VfLc9sm5+CfKGFNLAaCllJdocs/vrIgF3ZhHGMqjYdI
j/oquOd0yh88P0jJayY4H8sl/O0oAK3Dd85zSKYWMDBTIA6SLpS5zvE2aMHTZCeH
zmjuhxGxsdTAR3GG6Q4DeKUqqlfxU4PZcuu4z2trUwsCouG666nKLb2krGMl5tnJ
6KUqv3Bmkjso+5wZ8S2kL3t+IgsV/YRVqYFDy+CW1PD9+KsoCL/6YXT8fbOuOW6C
wA+tQEAS+j2fWfj4qYGvY7gSLUc9Nqo1FQbiMWG/I2H8EKiQ5JVTG7ySHxkd8gdB
z23pFagtSshOS/A4Th+R1aKb+FTYXiotljoWqvZIaCJ/sJopix/z9Y8XRo3la7Ep
snP4EpdYSlI5YxKnlTcvrAeB1ITKkcqkHVu5RUM93vJTkpWtxm03cNnndNlMDATs
5jdtldlWKj/ikyCMae5RYzKMDapyrhZFEpi9NwqmBvqv52Rc4/OK1pht7XaINSNl
TSRNsZXjQ0Fm8YfVtzbjf7SM9/u6s7ZPvbAmEbcsOYnCgBBGN4gpUWs8hUzd5XQN
U4wYyqBQH4WvAuiHJ58Pj1I1i514V1fujzA/PVpeb+xBFX+h5UIvww+d705jO2D2
DAxRUvKaSwMBIb+c1PPn+mC0Dk+4VHQHHlwkyQyTQkbC2BJHh15IqH8fV5CADG2W
8QI1QPxvZ69UwmwrpAjKe+jmbiwyL4X2NdNSEr69GpXKOfCFMSwDYCvDZV0a4LbS
cbuqi39FapuZpfEliIds0U0CKSFhQN59P2FPXH6jxWrFHt1HL+zSfSZK6yQCGSeK
uhrpB0mmTa2woRjLSUSJzpu7oZ/Fpa6srD4GBzhfeVbFflE8+9uEOWyLX+cxYhl4
5sdkjtERWL+bPAlLyZls28s6e775TJ8Zq31/vHHoXUX1+kjCpAnmAHiq6pL8KlBI
zTnutwq+j9mzvH/VDIKkrtfHrKwd+WBFtoIw3NAThrnBBY2rHILCB/FoxX4F97iH
XQrzz5LS+1/I2AbSf9bRRwzdaBReT6KyP1oGV5yR/FGsN/M3VxLCL/fVzixXTRHX
8Xu7NJIAsqaYlJW0CMXJU1tx1g2evhr4VzDHUvs7yuJ/Tyb/ZgjQXKNydCmq8CFa
rWAOQ6IPTtyw0aypXaVYneugvvIKlMJuynyhBj8wqNB4LbO/bpzRiDJGfpyCWDSt
I+ERYDDLAIFZELI2LA4dyMAMBQ9xbs0plq7h7z5zubIhTefAZWYrPE4HFMiP1gYd
bGpmUs6WaBbopeiw7S/16shJc3cJZuwnA3Ab953ZhJ1a17ORH+Tkw6805R4bPc5q
yacd3f2vjNcHuqsZjYGH9rS/d1PylKN3aQDa/ZpnvEISE7pxlS52tW21l9FQ8TV9
B1jxqUgjrsSUPc0lyknyuYH4IpKnnRdIenNHYYrtGcZGkVsRsYyYqRu87vsgfas1
FcUl9IGhwH1Uc+BZd+4d0wkNOQnqJH9Wv7OQmLVyA89wB4E0IXDwey6tsU+wwR7w
Bq3srN8oSMCHeqFTqgwKylJZCqzL6JCkx9UFjt7qjjwbsPxQHymtTzKZVi0sHpSz
cQqe5GKiXzjqwcPY1ji1uQtyWlUyvhiXOIT01R3o37ktBD3lIhxR/GRzJtOOUcDY
8E1ZbPFMa9xyOScaxDp2iFOzG/mgaRzmdKMCWmi+JHkRqZn7lnld5x2c7v/a7W67
e5vcdFPWSL6+IZ6xRF1Bq0dJU25fFovaYmQEUfVKlqAYyBcVglnEbvFpu8ip7lrc
G8FJllYWRAf4+8ukCax4t2hK49zASIgmr4mZfUjH8HLbIxYIEmkeEu6ihJMRw2pN
yyVZ/QSL9j2KK6itqUYGUxGEBSHdU3iZ6ggnN5SGjyRDpWBslrGtaHFO3baUkt/c
XuxuD+8mQO/vn21oHtdM4oNAqoOV9YWdmeFbMS2Ao0H0d6gZTnyD7lFizPWOGgcS
Ymq4r8N+hgg0i7gTNNgaXcTrkMvlc+iqoV7PzvU4kjFilJd3uEjGskQfDgUno0Be
p39tebs0BLzsT0sD6Q+TOpufdKQYD0Nz4rw4ycFZctiLJg+Ir4cptueHrExYQUU4
AWtpslb4iT2JFa5VA7Uwom7sSS2j0pxdfEhAFseVvwR+mIVIFAhy+8BSxvdFrTPG
H5YnIkjXaa4CEoI9UCnfdyZPEgl0dxuHoYxOQSJaOmiYEfzRiWF54J0ItmxDS7XX
sRYu99ATkkfIFrUi7wptdKqDKYRtJlsLY7XYoEN255CsnaYrZ5loFEj+tneeAnNd
QGzpzYkDKKMTqQBGl0H6iP0EqErFt2tpHVz5u/H7SVRd9iNes9K4lFnUBqeC2rUA
b7LYxAXi+NnXD8IswJZC505ONzg06PgVuBaj40KZV2phE26kD+FKxG8h01zeSXyH
9LwJe1UUM/p+h7KLnNA0NViitAICGmvhCNI/xtiCj5vA0IHZUYlJv2KezWjK/KqD
1Jt3s7PpeBdpJEtG6AdmwhbzupcvH5DasrDFz2covp2Gt4F9uDEdLwYaHXSuO/fU
shhgfoQtUVmSCElDFhUiD0RoUH3YdfZ/e1W0lrJRpAEK9HSwdw0keeVCsa1YeCcC
gu8ammU3KuVDTisuBsybCgNqip+1a8SH7CAg5305bR7wkVk0FeDDYX4L/xcIEupi
ixqAJvQHv5446+pC3emGW4f995E8pAe8SWfBdzVsX2ZS21RoGG+23q45iRjuN2g9
yY21RBdog/1kTYiarOxNaImT8ty9A5hLQ+4DaO2gHKq+SdDoJ37pzjxhgLno9zIH
ss9jd4JQjd6pIuc6MZ4+iFwkG3ELfzsKQuMARqDXKv/9WUamS7ZqbsTmG8voNqdr
64HTEIJzZyFXxG4zv5+jQkdmI/CKHIOgHEC15eNMNUi+eX+ehgcSbb5jlMdXoiw+
vPood4VOhVPL9deM11itOcqLUUyH/4H5GZNq70/x+rYGIWJyLA3G8nzGw6zBioDi
/Pv31yR0CkZPb7T1btdccJiuBljb5rjFw8xuQHlMch+Hp3Nso9otV5gmcSCtXjt9
6u4y2BmDf9ZG2cn3m3G1Tq6jb+dUM2NqSydsTNuR/NK+jEH39QmAfpcoYPDxNCiI
k2zguP8HS9IffToA+PxgpH2t6NRNLdFBcK6y6WcmzdmujaMjgVYc7beU95/VbrYr
c5mEVeBDwrNhqOEHBhx1jk6Ke43j4CF/WnDdHoMwvY3Az6TfYPaCy8VmGLOreW2F
/SllmU58n2CP8k5eezZAym7cb2Nw/6h79wBAZsp8OSwJkYgDwdyBY7dxgHXNAjjC
sZB/BCA2JimwxxYMF2+MEn4xjF9fuuTJnnEWv9LvPwF7X2xRPL8XAWN6WI2JlCUS
NzMB6GVpEZ3RTGZQomykp53NSDGSIw2Hb4LIJdRgDX7D9qteuhST8rytoXf1f6aF
kYnt7ZJ/TenRFd781p8KvTcdRJG2qPxdV3nuLv18qFt90/P+XUrq3Ed2ctevnjz6
J2nw9lhO2Gwo5w4moBWC638Vw0fFyuVEhBBrvPeKxQTKn9+krzzNkcPnvOEBsSaF
P80bK8oy+l0V+suZ5aBqbb+Pnl4/Guc8oWz0S81Ye6bwX/Z8jh7fhhFoUc8wG9m8
RdHZvQfFGvwseTsuk5kzTV6E2HQhtcEs46rPwiJAKpHltIlqZw+ooap7+s8V0LmL
t0YTjIbi+sfzjIwCDI65T9I2I+wVHrHnrqVtFh45T3CD1gVaAvLWE6SGVlCkPxiA
TsQq0SOn/RiveLNfmyOGSx/4hvp0wtxLhwjfb4eytkeWNXbRivFVp2qNgB4jaBkU
5ixxSOo/qbUWP0ZvlboRTSqUasuyCIaTfpn5ZNTSi81vlbVVYBXkNoCcqphI81/7
LPPxtov+fKKvLUh9uph2Em0vtkkmuXI0v+2oCxWmGy3Oi2k0i4s3vORpwS3pk2nn
gv9Er/Pq8gNtdbpu8q1iFd9r+aWUG6f6lw3OjvufaWHgWljC095YWVME3MU1MJ0U
t/yOQeXcj9iYErfLSfDsan0eP5qB+v+y1yIrKVKaN2Ea1S3ZW8dDU11qZlIwn7Dj
KVl24TQ+ze78lzbHC2bbbg1HfV4m0Gz/G1nWNvP3UTrAoRfa5dt05dggyxx/LK/r
wVSI6cEYTSM9Fgu2dx6+idOcGXYLyarvWpRCiR8sFQeLp95fvqFeAuSEoZX18QMe
LkWZC3fcJNuzmkFcVafgRVht1pxG0WdQ/gDymuaEXSLoNBdtUsc+wLirMoegbR1Y
/lWvKF3cQ/3jNi61+XWqpMPI/SdQspcYc7WmWoPZhCBOG2KGBHNJ/doYzQKGfpfw
2nUFdoowcx9RRuWldPlxtMJYz3EDvgd2xwfVez4zXQqTlvNdoFIQ9yqtv4GEKZdR
K/AfI+tcg5bH/wJDLscqZRYX6lqYmKJbNlJcAiGcPfcYalBIDJPYZXR9kk1CW//X
YeSmFlKD8af47QnYBILZ9DSUv13sEiFc7I7Bla6wrcFNM3/GGe5ILdqt6RqtJCCe
H7S7iDNsMt0RQw4Es6lWiFRbZIUbVEzKz+Rpp97+SKcUIIqDtP8JwjIsT1wCU459
YOJJnd7D2CFxLyMBMXDUCDl6sGDVcinRmjk0z8n6LGF3iIdceUvh0UpnLefOAoX1
KUKC9caxfE0DRJ7pokWQjaaPe6hD5O6Ja9DUGos/OSmnoj2zyldIZJyLLOIqgKj+
uFntAOeGZQz5qoAxAyy+zXLdWmqJWWQIaelkjxEneC1k5NsJTzq1iTj18a5PhyXY
Rbt4QlfQb3hjdBTEr1rpGKNV5u16fU+fishRlAGZ+BngsFEf8BVXbum+wKq2J+xN
Wo4/y93l/HoVabb/baVNRpfq60jA4Bm6CeDUW5GK1gSQ0Ku7wbmjnNDpiAZWevvO
5+7UEDC3SMPXBa7GL2NQtDME+6f5hiPFe7+46CJ68HA2IizfUSDgAX+vLTfz5hFf
2BEg/iDS4D8JJajYnAfQBHYtPCMxwCcNZQTxQ9u8AHBuymTPN9E2kBOeRubTGSIo
7BBpyDn4vyY0dQaaqBinFMROwUK13dCbZohFvcSrBQqkY+CxXjRcjSolXoAyeGBM
6MN7NCKQQywUZRydbl/4klS731ojWLYQK4I/oqjtE88ZXmiWvgznyb2o0ZtPJbpL
r918dV0EgYT/V8jKqgDT1BMCxQ4KVNXU+9A0VoRuSuHwg5slt5dq98uT1KiTqrg1
r48Qz11/4xnkR2b3A3yqSg76801Ra1pKKihODiNawPwp/CUblux+/EQXvXHtSG/b
3Vba7VBfRu+bGfMatva66ES+dPc8i+61E7DM/s0HaDBs6e52yt328GEC/N+cA40w
P7uLZab1GXIX4BMf/0eflwkJvB4GEWTX78DcGaF8l9ikRpN4SMAI9oTcxQpYtw4K
LCZwWPAb1RElF6fPpe23AnT0MbqN4vRzdOtIBcYQtEhfm1tsxecQ83i3wPPaNovM
ZnYJSrP4gTtj8wWZNmq8nQDLzP//Rlun8WPZuOnR9LcqEdrhnnR1gHOQ2m5yqASU
XmCWn98W2F+IJiu0EJmWnHsV4IdiXyrNIlzy9X6jPge8BdomFTpVvkgL2v++pHi/
CAwb7f465/OnFNBG8vHB1m+DXMwinkVs9hwkfjZeAj6W+sbhFovUiKztKxJxQO+1
BFAvZlOVEL9HyhnWPNRcbwZg0VvGCcaf7d8jCLgl1YBEvrdl6JsFXu0isFUqVguJ
F1oHeO6m2Vjp9rOZqkUdJ8qS8mW3Lj63Z4PVQZ4Bnvii6NhY1sT3kaNIIY7yju/r
+Z449+oO5FnlKzW0hG5u2ClYVR9/jeV3f4EmFuCCE75UfeeRRTzBaNrr5ShUEuBT
wrn4k2JbDx8/HXZSYs1RuXpSsRt0tYV4CQFlSPHH7efBsLZxuysMm9Ui6NSeOqeo
ToDPbWuONHVUKh8rkkISetd2EVV969cmvjvxAGwozPKt6pH2w6CbVnw/8SeBR3zS
JS+0zYtz5ARRoOeFVWipC0V0KqKMkw549Y/VFqDv/OuVhx2pnxDmodfMh/JJxEY3
zQXxPLSXbCQUQPrH0AlJXuUt8nSgydaAzsNWMdEIekJH2CVtDApAAqUgZ73FM6Am
hnOrd7q0ZmmXVurc4f2UCyvFUJxmkpcEk8rTz/h4yMzNZ4CSgDf6pjg/OAVXj3Uw
MFVvVyehbLSX52ko6ffhvlar78j4JBoWs0RyLfqx9zP0/XisVTjx3/b5wQbv56nz
tqDKRf/lC+05YWUmxye22MXtoPZKvQxxd5RDYqRdk66OhHhp3C5uL76Rjzsq0Hks
TzP7lSXQFiXJTRPSfYL442jzYo4vSPvUREZSVqycIZ8MdSQIC0sBZyfzCW5ab+Bw
9PMVyL5v/G7iOU/JRaGLgWqaswHwazhKSvY25x/iFN38yLKoFxCGCKVpEHFYH/Qg
oIgmdWiWvlpS231LeKLKfqRylQMAGFErH49Sib2YuTYIe4qm4D63qgS+7LPtS0Az
+gRAoKwJSQ8EbmvmM860lwS9WWw+TC+zWYky7f4n9X1yiGPN/SaUuxMt6MwT07ju
xfXGc4ZaoO6CYB/EuWKSfiVNOT70UTTDS1TwoDn+gjwS4hjBqgoFL1PPNNYOUQBg
lYc3gVAh26ZMHdBcenLXdQX6xltpCVGibgmXyWkofcJBps1AeptSg3fjFlN2jPPI
T6FRHVn9jq+oSLv/wcKfx6KX0Bj/v8FY4q9xROa5RuQdqU9k4DpZ/puczcLdYDTU
7NK/eUDnm+tfKVcfITByROf4qkqX5eJoifd71vhRXAmcTzgUravDQKQLq15j5mrU
u/HafK57ac/PO8xcWKvw4g7MfsFGPclCume9h7Y2idrb5ty2x+wdpCQeCzEhTqgx
/a+vOCIOzQHZM0A2fDxQ1BLNE+4RoDbXW1JS5C7DoZigZ9dHYRcXwgtQreqgv6pe
HTObqBwF+jtsWFCTs5gj7qmAHO+L0kOOx3GL9LjCbG58Xi1gkadqLxZNmYb+jVZR
h4cNFK2GEUT2BW8gar35SAA/lvlo2lWf7paWCjkrpa338HH6XlcDZA0ad9eGFu89
k9B3zHr1dVgbViExVEMNPUyMsytwcwOiuwbPW3VRMceEyrFflP65tuOuC77nl1Cw
ege6Df8uTA7UIFQbKLtiwQagRihbS/eEMHWxDKksCipazCMVrRN0eQmeIZcJVClJ
VYD+rTCOee9rA4d6guAzcnIil37UlFFpzCAPwC8xD+cNtc07KVVMcIKtm3aMilN7
FcFi33yKFyTlqb7o/ea/vnLk94+SdOeM3i1Mu6spA59NHFL6o8mefcwCiYQXM32p
PNgOqqP27jVSn1VF06KpPtT23/yWcuf4SmYv+4qqNiFZi2NKq6xB+toaWPg7a7yi
mqbQFyDZDt0aQ3zntqdPiXvt+PuKuCcmFmSAL3Wd8vgC4R6esOLq9VaxVUU1Hais
mryOaINF0pHsFbb7o+oBM4r5TqGGaTVYYd1gaxhii1vQCXYe5ceodyanQgp0WPaY
RCy7OfSp1Afr69s3ZO9BQm/Y60Cm4Q/nh14TFfcRSXWI6z3X+zkB5J8SAhWnpO3r
wJI2dSzutU4fPyw9NJ4bSnri8uM/gv0fD6OH/MwGFECtp/dhQPHaHyFFQbic/F6n
1HWKNVbp55JNACjvTZT1oBrZVY5rRPU5+MpCeQLqvbfEuf/4Ye7JBTN60Mfx/FvD
wxXy958+NMXoq2LtWURsU8YpMc47LG3JC4lCXzTdkPckKtcoQgG20EWV496AgWgV
PFlx/khHkhZPmlo9BxII7o1EranNwy7l6FikQYq9UUznC0cutuAogGiaRiDqQJ8m
oycNL7+iZZ/nqunHgDkn8Owuc41d6CX/kPUdL1KI771oQ8xNMKib30bFAJOVRaBs
FNNCaVKGJvTFySGLI5URswvbYVTjBkXHKIN8Z0q1nFQKCOseY9sgdO2ZmcdlciVy
sc7OL8/gTgrHkxjihz5vckWIDf2yZMVf1PtkjJpWxNOqPLPLpEUc0gueumFOYsMH
iAqL5yDI6ydy/nX4XWgE3v/Cc9wOXtv9h1M/SHxUZJz3LDT4TWxSoZLhNCsV0iMz
7eypRJGuW2kQXHaAZzydg+ieMJnJB6KfrrIcLMDP/PLMAkW3YhOyhQf4Lq8NXG8q
tgYXtK1rbXbryVH4TlDO0GjovKTIvqR787AoXgQHL7hkbd5QKxqe/gUkmtrAmffQ
Bw3KshC9TWcJ85Z5qhwzJByXNMrFlikLb0fAG0/iCt3yyeAWQzSIjnbO75whd3dM
lb9CKiVKIdAvywYKYhd14j2X3kT5+wIkVI/KpkMZSXXXe9tSoabfGZROM/PmARU3
qAyUm/+F/+xAZGepPkt/tpGWdMufGHEdo1PusiL8W1K7jbQ5nX8hJHOPaQSNtx8e
r2fWY8+orHjw7Hyv/PK1RLLGcBNbjN0ey79gaBs5Hqnz3ttKwOymfJW+dJ1xhO+/
CRzLgsofjeg/NQ1lFNI41A2g6MYDptE4kfdA7w3yz6cDnM2+WFjC72KJ+xBAYtU0
R3MHde/+GRP/u4BthaIF+Mv3ESV3iSFun2T2XorIJPReFZ/2N4Pc9YMshAPAOV8B
SIS07Mai+C33VQiRWzlBb499pyY//y0GQjlaqwSJk2Mcg3t9U0Fkziya6N257VZY
h78SMMCIVZRITPMP91R057ZdEYqdToK9L2GlMPJplzO9Zo5pDKLTQlq2G0mlf+6i
vW1rf/HZvH/TzFZ0zLSz47lrFHAckig7V0lYZgm1GZ02QyAvqfusHWcg+jkt3Ra/
WSa1dlRRhoESYzWUoCVx1x3D9pg3kNmcgIUAdeDxFC487yfah5ROVQsQDtzEGGLF
OMRcH3heTaEsCDqUiq2xnAD6P3WqRT/JGCdfYShSyinElVboyvE/JtvkTE57Ihz4
6wHXKiGgfLG3uGsycZ4Ds7NP5mrDRjJxHZLx1NcevueWqTwieRkwLUYyAro4z9N6
qv9M+iHIm5Wt63WVPIVBUpDQlfs4hjFDPpnIN+82bIF9CyhpKz3xc69ofEWYP9N8
fPnWaPq9mRn4pxDowQ6HctuVHdRmHOmrJU/j6hKjE/NnutSm+cOQp1AaA5HygfY2
BfGqHSzc00A21phQBVb/Q+hFNu210rqDHCs3RRQ+gHBhk1f0Pknc5CrJNQQikibm
fPUktPpHpQcimFjGKKTAW/VxCTbWcCIv8MiXD/aoGADNaRB5chM0EcFNqriFHFEK
Y1+aDJX55aylSqjnNaZ8bNzZf6T7vSD3DCfPvbNR1aRes5w6sWCImsoLcEfcCnqO
rr7ZprroUg7A+9AywGroI6rSV4EA0AxjywwcV/u9nsm453XmYTGWehcDM7nc/s4s
Xvf7i86BHrdC4y9ULkISxVo09XrHDLoJTlNH3IHg/9joJ9fugGfVL28ToDVEOUdB
JDkxx2xlmu0qeVeGE+8dv0JetVWB5uzuAd8LrOXKThkFvXi1PiP2GHHYdSoN7Ag+
eKU3nrsxK3eKbXTM2l2gSzJkZmUISuSXcpwN/9fB4Oo15HZ0N559Oo/mXmVCcx7E
CJIDbeZwnG860j1BaE/rMj+ogSexm2GgXMRUpHtt+dm4fvsxYYfn3DQLvmxZFkwU
oyrYDXZ+i+H/khDHvVYH5pP0ceWxe/ahIcB11Rx45ORUc+kuHLl6BUThpA0ySuxV
/Ul0iPWuQUXHK+NVXagsgp2J3A/fuR3vCso2JxhU2QoDDkJLz2fyh4Nd4bwc+JSH
pN8m6WLmkPO5QyLxt+MoyQBIkeQsI7gQ8y/o7RA3dlV+YYF9fg7g2x5CoVb6EOTH
A8BgT5HYOHR2JRDK8DQ2asCyNX3O6LNG/bXhGFwqQ9NNuHh2K4aOfVtm0efwMsuE
PEla5APi3D+x7pXw3TaYc5T/+j5UQuoqMJi64leEntBuqfoioYIXbnmZth6HFrQE
3RJE4Z5m6xqmh+9WfzcX5Dp9hJMuVUrBiyINvsPg7rc1mix2C50tVsBeFswEP81Q
PzaqriIfHDGvzcBl5+DWgn9Exnvr4COCpGCCKOgAoHyiJbH4NqWl5h+CKc5M5KFa
Hq3oxCikAjQbgJDm7/lBMJFutgzRB+zkYowEqNtkRTfJqdD5msDUBBgRvXZjjBC2
qc4vk4eXxnwnTAH9AwSlBdp9x2pKTD8sFKY5Nfilxcc8/kG3YFB5CUzoBw5tUfln
Z4qOvvuSydwDTty/D/ZAbgWLXugmqUfIP3eAFjEsm0+9yQ0eAx0lWqVeJ4teP3vR
8PcfAet2k3dKHQdBVhtm9znJVf8E8cFAHUktch7sl2GVAYGyWEoCagDZv8KlxEa3
6lT+AmZloRioGbXldFQKiTKK/M4fpoTdfvIFAQbwcsaeSP9G35jushyCWewQZTcO
+Sa5ZxxFmg9vioKIRifUln0JEFE0YI3f4HivfqU8Z+XChlLgQ/ilyAGRU0XZEIud
ee09G63Z5kmxB6LXYIfQ1Ah/41ZOcV5ybwS2/AJWh6Pkq2WRts2YdUxjpyiT7dto
LizvDVfmED52gVRmKtuk75lk5dw7ut0GoKME+aPMLn1Fk4GqGbJYPdgI6ZEiv3FC
9HLnW4hRpPQ+lNP7wLiGDmGcgGndJuzHSC2vfP7JkfAbQbYMc9uzAIXY+4XDnsUt
U6AUh/YiLtHHjJ4Sj/HvpMrXh4xEzTZc1SVuvmlb7ZgUrkx1LmZcSRuuOt1dCIo3
N/sOh3SRsc4PWsJUGdNSjvB7gzs+10xKBXJgD652Ptldbo4sDNgbFIDKjaH2YKGR
H7k1fUVd9UnTw8Wmq8lQN8REYA9twgi1toNRsApy9iMMalQ7YMv7u5soxP7eAkbZ
nb07a3TbEQowKrUn4/D0Vvdyg59EH8weR9VthdafqGdIYBF/44yfd6PrdC2TyewB
DZzENNqtBOesOe2fukcJlm8j6lLOHzKHWdVbJx083ipTLh+CAWGxYlHxIaYSbwpz
flAOkMwbI8tmiVu7U7LiHN7vWgR0T7mKr3hnNRYbnxPIgly3eK+ZKMeASzzlvh+o
v0j1DQ0tpieZYajjITRpSPMsiPX8Z0ktgX682iUD6whC6Rz9hhAD3QX4p01eZ/nc
L2SAPArm08yzaLd17K5bdBt5o1KjEAzdF+2tSzv+/Vr7jS5ZxcC4kKLSJsZdGnTd
eE8PJVPbqjF78zhu+8uQZxNH5aHzOYJOVhc0UhN14xzltlEkHTVvVeJJRb7IoAWA
m88psNzPZp3TeNOVmHpg0rgCMPFvz7zhJtgfjW3cM3MDznQdeGPRuaKDEKSdcRVH
J0WohRCNoxu3r+XWSm+pes7AYfVszA9liQZylJKCGRNvhSylLmOOBWJS+wBdjyfP
SxBJR84WjdSjwskYV40zhrjAMPtj1vMS3B4P4wWy0UbHp333oxeVp6AhOUwGKxmB
svBdEhOX+UQrtyVqa4BxSgtSYl66qMNfG3TlyTiYdi7Ce84a3gp79d/ATESsnlB+
ENMpjzLY8TIHYU9h2BE41XkD6MKBQtqEw1Qm79Q6fSzFeXnGalw90Zza5f56Zf+0
mPPMogAFqlY1UA7Zt4Rg/74cOWWzXRWeehebOxZEhxDMPvG+EQvLwefbVRd/NxcZ
WefNmO9vosvZEbL43T1EB8K2/0SLjVSRbYx82Y4K3bJvKZEONy3A5qBX+rgPUzDL
+o+YLim8pVLFgy3+mtmV9l/mOvPq6yXBw1Xrua7cFFcuy1kVlxf9OlpxDhtU9xWv
5IfqpOviK6Y+/mrT7JtBIfBWcxGY2Q/sXveohYiP843H/wSy4gXQ4aqyuvKcBUuy
tjtsuLyfLyQCETLTWvsYKdOafo6VUbMlTzYkWoS3gVD5Xhz/CBjn95QShGy5ZyTS
jT8lSvd34HwXNiNIX70nuIQCUWBFcpizIPxsz424PiaZs8vyF0GPTraSrcCyVPnZ
tmrZV2rYTPDmNhkzx7XYSHrOZu5DGcDXA287axkNjYd9cssFABWXk0QMO8gfh/Ix
zSnghcxH4ehDI7xl5xQ4J7eCPEP9VZB5QPP3V+HexLrz4Fttuz3YSsFFfWKcg35v
VVbOwzox/7UnnfuFiAU12k4Y7NM6KB0DDFj141lY7b+a3OJ+Xz2xY+DolmkuEHz5
StuHtMGGKlD+47tAUu/Ir2X5Ga/ULUILkiCKQPFeM2Q90xBEvgXx9YBeooCWNzCX
9ipZg3UN7LikDr6/oIwGmLWNHdiuOFKE9bvu1XlJOUhTw38Tp5P/J9pRvf6v9zAp
2jEPDvw4AkXsfSabYzB1gSq9VjcSOZIKRhjQB/NRgEPw3LC9Cc3jotit+PaitAaF
Ybre3KVFzI8mU/GEpfaOxVXmNZlLwc7kkWJufPZVbZnzOu6kTk8YDCScEBt6qIFs
cxAe596j7cieO5F+BynbL/LWH/A7e2xILcTIQtjo1qL1K+nFVOuFGW7Q3yzYt5pI
IXpj7nzSpES5yDRIIpIhVcioeWEBSNVBgIWNwHian+qPYuMY8yoWwtTJvjlvq6D6
9bps3udIKY892O8sJOqtwSHYeVb/szUxqIYZv6X2bI3TEQu977Q0a+UqzOzlztOb
w9TmDbGdonp3Dl5bykj0t+LdwOgpk5S9pKxc2K9gcgrz2KlMZnyxUJim9Inv/LtZ
6NNIkqdVgdmtlzKj93/WFavF+QznAbyH6r0Y8MXu4674TLV6ZcuKdkUJ6oPtamwG
nU1GDsFK8YYma4NEBG2ZzqYCONnDyAra1Ci+a2FpaFCy4umAT3PedZ6EMuT8U/KY
8pTx1MoaGRKN1krVU6lo0y4sb1YwRjSXVd+FZhE7VMPE2S7UdPLfjeQ7TpReencO
dD+oEniDm7BPCQcsewDeHyjPjyQOVaNyWfORSiFhXeUcQZxVvLmMeu21hxIkr9o9
ygycpFGT1gbgH+bd+d2aTEIfBbPX12Jj0gK1c00RyCBvTeOMrjP28HtkjSgRKkwd
gbtScAh6zfo9yjtKTAaMQVyKQN6VT1nqdsAXOiGrXKOWvF0vpSjqbRJWpOASWuUY
sO7nqrI5ANcXHwJDS18ogNQSw3gXh9fSu4Jypz4+loJLtSH/6cmXfmlnWnDlK6Js
jQW9dMFaNaqaCwLwylOD8QTUpIYNur+4DVkgestc4WGeyTzELh0NfhicSnIcNniI
TiattY5qz/Xfzqcr9CMLVXlCscOh49VVI4ZjaFKaPwQYQXvqbmfNVinsTgeQUjeR
GbOzgmUcs6obPrmFOyLWMkBfj79AO8FT5E5DD0B3zfJ3+1uRPkzarONyS8UAhdPN
gCfn/qitEcGS/luDw5KzxcRi3/cwmbNFa0dMbskIYiYBH5r2l9fueHZE56TVAmdd
VKzcw5IW+3Mfy2OPob0jakeYIlw0tY5xAovPCITYfXYQ/R2obvPrtdxBeB7jJfGe
1cZBIBr8s5JW+dtIe1Kn2DuKv4N9b0plsF37Xm7DgIhGQDfg+3IEryqgu2HKzX0S
9sUWv2Z/pXlpovv7eoqZXRigU7DpXRB8TeX+PU9ZHgGCTZjtWoiFM3hC9gCvTW9K
sp5Zsjv6JkuF7/g1HKMCNelurNwRaPjUxRg0t8ZzQcTlFKWue89r7DH+jTUEWm/N
yZOkiMyWvE17FG0PYvodffy3HQO5DQpaX8OkZVobv1IXivdj10Scg2TL8IqKR3SS
fudB+2HHUW8HGaf5v42faVF3C5VyzD8lNX2xLK5gB28Pqzq4HqfccMQRSuZBkELC
bRobSK/qieT1AIFOCJphYyMIIdZFkWb75G8YZF4Lz6xmaY1v+9dofEyX76GHgKg0
Ykc4VlixEYot61nIwXzsr4dOBfQp5Cy+oTQqyHjJYg4j9NSBjc5bWZnkbsm5QeLb
YNUmlclQTHp1g8yWwKYQPbEj6dfUvvTB2E4RhBVj4FCeb5IbMXBwLm3ZXHtr0rxI
gyqfiwTtgoppGbZsesxdw5pzED3ibVmHXp5Y8Msz0bs9H4Lz9fNaV8v1h3NSA/YS
KBw2yQ4xAvQB5ZA16NsxszJUVqcEkHcTpN6/snHaqk4Yc1zEjuPuvwFmil14OPDE
Vs6WwLZfmsJVzIdX1kr5Uhf41HfrKAY6xesFYy/qHboJHdTwp5ylczoayWBZlwf2
TjaDngPVzWuXCbUv5dwzoKsLxIFa5QCtlBTZTkhSzcEAaCbq2GYrpr1mrUvhTbnk
vcx+O+iphVM5FouNSwHs8rjAGd8CWnzRM2E4f9OVt7btQ4xe9iHyKgo9g9FBEswT
RlPln4hcW0N1m/vIuiyrrK4A8r30z3dqlSK3LVhir6xJeLlZINfI9dZFv11NMna1
GalsxhHkohE65z5PVlznXfMrYBGBORj6xWvsIomeNuzUAa/dzomXOP8dz9wFpscj
PtuC14BLoPdJ3ZKuz43UccthKMPPn2TUaqEzsFh96vY46e4Ql4L6WNm/IPw9sovr
NbqMVhEtd+e7zVp1G7RhuxEIx1Y4Ph+LMGMOUBAfj0GcqiTx1ZxO3MYLbTdZxHRa
2sdIRXG7WnD89xHSoxGgaDFfUjj5/Lerg1JzWQL2ByLbWooRKVnPofwi+gY8BBgc
0l3hZdlaLnoBWkFxs1F5dzJrWa0w3Ci+wpUL+2evcVYfYD1BKDgzF5KFmgXP+jMB
pEC/LYA+ZfpOCA2xxFpDY8NPbLyOWTlxNxyN3OGisVzXOgJleEJT8cUGIvjsIg2a
GnxHX/IFam2RDihPPHgmoTLqtZsENxDg5P3UpEZGZcZyokaa+0ceSg3upVBBfCAM
17f1rjfDPJYMVwh+1HB6vnBeObhkgX2uR9uQnyikTwfSD8m1Vg1enMUSnIjxRPQD
cm8r3haL4w/w9eKxpMT6zhyP9DvyzsylTlDh58mrkJl93gCzupijg0jdaf4O5apK
T57Mu0QJdX2EzqwrPOdxY/pD/nfuSD+AlTJAOeqxGbLVKX2iRrFTa/ZgV3YCv/+U
X0Gy21+YgzFtglMW5m+E/WCZ3ISEou8kPfaAEJgXvaOoHTPm4MutJfn0e674n5Si
F9uvP+MLOeD0jh+qczD8IFma+AoWdQpvZwqyplV10wbo758Rw1eAzC4dPuYHtUhI
gOk8MfNyFdjQ4b/CrFX+mpiP6g+6L/BH/+hfo/y+yDWJUXK673PAiL7CAN9+Ephh
+LDERdRCL/MSRvleMh9x2UNOkr7b4mqapDriRL4wWoqF7ewzMa1jZPlgeU5xveu2
VSZ/xNWf5DXTvba8WvmFVN03RunM4BmoSkP2Pjd/M9z+Huh8TQ4TdaOL7hlcTkjV
tuv98bqtkGxW5l76i4uI9SvD01w+j8xA4ID35y1+qi2JfHXKhDosQJ9u3/Bt0mEW
aXbXGMFeRNlZfTVfj3ijOrwVB6UVQ5PcQOmPbevDOgF7rxBrOIx/gKSX7u0WdBtj
J1+09Y5uhkLwafOjj+ONmq62Jw08Xcy9W+IjkTGHq36Gcyd6+Vd7lPvV2vGWB8J+
kw8M7zA1uR/AcE6GCtzBAR1UFcmhm7+HWqGFXUu256ama8kwlJe4156QUSQf5cBG
fJTzvy7ZEvQjF49Ezo4djpS2A3zl/o2phPg/qB3xproOmlFMx23qapMjzX+90QGS
rXMBnL24TC8N/n6r1is285rhWRneyn6kvQ03K3k4zQxRQOUKgqEkeE3QDVRf5nYh
F/tX+QpO3DR/xpAU0QCkQjA52OuFgInBeDBAJj9BbbwcUFiYBPcdAWYB+53qq8Bo
6NJHkIXMNpq3YznW7+rh4Fe/K/SQuszIXtz3+grk3kCKNssii+qVGBFsLrjeFn6G
gCm2iVLteJWu767n2eq3e9tF/dxOVEGUW6I7wjUZWqqcfCA2dcgQTiWxKI0zt+0O
4WvVxAxX52uVSXLZb4F23IhCRwt61vDtPmACs3IL7k1A7g/PvRnr5wgVrQALKFmj
ZEKxJZHE7E2GrvzcbJ/klEB/H1iTeZ09tMKgRiWPWIXDsXFmkUp30OzxZUs+A+gr
w8ty5ZSZMOH8+4xyIBm6lKSBTxOEDJFmtZlXLnM7AjmqzmsuQLYwO4gXQhkNxpus
940Dn86HIBdmEHc6aHk7Eu/MfIHMg8n3XBWTL6Ya2XC3Ie1wwPaCLSPbxIHvOcO/
R3QiBqMKCrCALCYyLF3v//+xXtG6pwLtaVFnSdKfY7U6fJ31FaCfqcjm5avKBodC
ZsyulHfLHWfHcIrPTLUEodNWBfNx2erQImIWHxIu64lqyEAHCfS8UvUAXfMj40w6
LjRH7irfvo91WxRhNaOUjmJ7mdLtjQJHsdSf7fpXCSPz3MI48b9zu1SS1/r5lz+b
QuKCk1+7UdRvtTySEiNHNNO0CK9XPVJGetW06cP9VVDg7S5fiMWR7dyfjrY/lFnX
GomzSw7B8UR38owDkh707PrygFHHL1VWprOTYQqmVGLyaJo5kqoxPC3XqVAtOXAd
Y22tYwCjY3KRsG6ARJOlyfkaUkUxYX0qEVKjq7Uv/0bZFzLoTEWkpftRN5mLeUnI
1MhE5VKiS8/hf2+GrI5Ae2DzP8bef+eECWGROdFQ0uWf8XTKUfuU+CjoVc3a5qLY
Tud6Jib0ASfO4Xsd7HSYfpFAtHvSl/emYoFU/U7KP91VSi1mfrmzyWqWoY+BBmzi
kJeF/g2hI3hs0XAMT1X4ELir+wjBc4zZPJzjImBXdG+XLN9YeUw0Wy6VVHHqnWq5
VoCN4NDCb+JYdw8HHWx+1y4isDd6J3DzPQl4Xfunfia6QZ5QnvDgQVheqHG3pV+Z
ecZgXJDUut/OYBOMOyuj3gNEmGu3IVLXGF46AnY3VOjd2LbZfZ+hYGGD/p6L1gCk
598S1OPZkK+bmiMpd+HG2Gw3fUqq4bzqOVk7Ut0uQb/ltaSzdy+MpIb6UdQHZhjp
IApk9Ns3VHHSobenTAwnnTRdZ7UYjwHmWCuP5CNnmyaFV+xJB+TauUbGUZ9PE9LR
nBbJObn5TUirut2/ZGWeIfME8IZqfWOb+iBki7+oNF9LjufybNMSCC6qOr+wEY7q
LTznzhix5xT8wOtVbEyr8p1WCi6DhPSnGHs9IGYfoATziLVI0LuezU9/mSA/DhCc
1tV9/acnvpbI4jd/+XdxXg7nooeQNMl7mBEIv11XfloULcj31krEPx0haPDiObBx
m5n4IWjKWtPql7s97yFwndqHwyPdi++aWLeZD9ayhMBZHuU/ogDTzp4DIsAuN4bu
HDF5DUAs+qeaFlwFCH+DXDSOr1PctnqkETwNDoG7VtYjQluU62qiAYczpkZzmirb
239bY1TuRqxdatoQDtEYZ7YYkh/bKsS8gA5bJxkC1UYPccjRWG1b5Zbhbxx7pDRW
ZygZm9obNd6z+9cXzGDvfRrVJiQW+vODTmuxcxqa+D+i4U+t6jINbpr+lCCo4Auo
diisAWX9DDvhWRqHzx/m64Chck2I/QcaYgAweyrI4CvE3UbM4dQQ40SSDm+dQCD3
4yRZcpS0RMiu67v94ukHASeUTfNlPhAE9IvuiaZTZXE6EQlhr38OjFZA2dj44GNf
XXKLOs7kRCMdjViQvwl21hHIeicGsTyYnNRyBiq+S+auXTw5lRamb80OWkX/zzjc
6P+a/cTXqedZJ+wTlTE07WpFRvilTUfuqAuUB0xqtZ/aiI74RQQU91ZUItahta44
pYat5gxQDky87SIXULAeUT9qlfmj8jAj63VWlh6klHI2oTTlvL8FjsurFQKB7REj
hyE3WlvipBmW/URysvR8c33ym4Se/wPx5igFshE8qnRF3BpX7gtp530sWfKFkB9i
XvcTtsTZHAucwZdLoxkVBcewpyKXedx6SOYwLlaw343MsquDScGRM4v5PDYEuWM2
vctGbh5Yw/rTfeAI8h1fWrMEmbgC1YVWgmyM988Ssdj0LM1GLboXINwu8ySArOA2
foYeAcVlCyhb9tT0/Shk27SGo0FL4mb7E2poGckUwll2LAdqFkVTHEuYUiRaaEl5
0hYvs692Uuji6/IKdpOmzwHmypzlnT7NYV4deTYP60rqbukFoemMlNERpt9rDAPs
ZKsTaWmy2rqaydFfoslR5HBdp4c/RQlUGjfAg16cMyxu0C9ur+JByvbS5GO+JukE
5A73pPQUulCEWdhkqG39G0cmvYamAx6xLr2tkJuOLzusYTqIBHIvm8XgdykzIOdX
0R3y9C+wl5aEEY8RoHehtn95bgeXoGbG2DRGLrPO49gps1ysq0SK71fLfNFiqAxD
e/urC0BR+Jm1vPfelYo1qo/6PBQppFzWj6fBD6+ry7Ek66ZE7CtXVuR52WiXB2tk
ZEa+1igZM3STmA2YpWxH3KN6EPseGRSdPpMxVoeehr1ih6OAbxgI1K1WpVZbaCLK
85bvAu7pnR4l0n7AkHZvt5WcT8Jy0uogqrqIReTOy2LgZunRzKVH0SLxs/Je6coz
LL37zj8I+E4yjOyDvHR8zbAjbI/0eDD8lPntd30REj63jyh0/+IB+IBZibHeG2mh
kctGgCtQI9GTW7c0iEi2MnKKnStwe3rIrkJivNcjjVvPmRv0adk0SmYT+N9oPEgZ
rE7RAaQxO2GttnO8h7l8IyvvzWii40LYJDCR9HDGE5OdY7+gRF/tSenXFko7BSlE
inVGGYOCxzrsHJ9uw7UxKBZiC+iwOBobJTMCBv31B+ddoLkG7ptje/j+PG5lTYbT
8rREmo3r9nR+sySw0W3sFLOws58pJ5yo2ZsGpKCJcLL+Z5SpV2RZWBypHw9HVO6+
4PrsucQ3/+81J/vkHX+JpODrQGIykAhJYeUiB4FxfsihJA94UrkrNkkTmNG9QC8l
2nApfPwahm4mNInxFvQrWY54ADJMxPaL4lxfRq1rzUZ0oJbcRyaB+iUjbetI3xfu
Ae8QcbTh4vyJynAbhbiGfHgtFkhyH4mhKwZdxWKxHYxiQ4vmnbrnUPQb0F48AGq6
HRJ6nugoSxMfT3KInz1vW/g4pSnT0lx3hGa+DtBvFiPh45lmbjHSBivwLmxmrxOx
2KOsAo5XoEysxi8MHNyZrULfYjQk6MXKZQE1v0TERogNvsKRcnBps62bNtukw7wh
8BK5xA6wUFzlSHNw0rJt/DjdQME7W5vlHo86RDMy2ypCM3+n5Ol8q+8HeY6tF6vw
3dedILBYXmOzDoD0EJpt3dcBkWHvGndSUKPnk4mSz4sT+i8KVX/uLr5IGkcl8cLf
I6AwkSrLWyjKLHAkWopvW9M/wzexTIgVQZKtg7sS1oy+xwp8njjpC1MulQWp3nYq
l4c1hztSbNSPUZ4WbURyiffJ3bRW+EWFHr9DDg5j0AU4xETkF0hmAmfJBImspexf
1s5KIzHFfjJGkOlGJojS4VhVJjfDIPCz8XV16yMfZOXBlBy8W0gTQz8rKijC18GY
oQ9b1DklBBG+B9bGa7fRVaTCWm9LFhsNIV4UkIXaR3IlazPR6WQrmLk48+LCLB55
qM9lNpILGx04ZyaCpD3wwRjY3oUsxaniJhzDIGBIRem3XpjheU+MZi2sVysSZGiA
tL5dMZ5omo0/UOEBMX4SGuHdinpw+65HMYhDqyVe1SD1iS3oimNJsxsTRAYK6ItR
PG1Ht99r/YomT1Jy+5DibJETa06pHsjfCMdpVKX9B/bkwLaAtuqraY79IXqcksq+
r5kGeIn6o32wnB7zyy4kBSHmKCk1klZYeIlWT0OH04ybHKzLvO2vyR40kSJNi7C9
a2CRB5PdyBZoef+52t0EpjqPOe/GfnwKqjcT0NqrLNg5kNcO038eb/+Egig5eTSY
rztseKjrIdDZF9k2EwCzTpOwr3IhndUiX7iO7eRio6LaiYeo7f6J1uvnbR7ZgZgh
dR1LOzvCG5HLprm3cmZkh1iI6aIhj9m3vA76PjPo/zocuXPxDr2atIZPWDmV9ULP
TkjVqzLhicdB+WvDEdo4kXEyLVQj9vQQGmkYEHT+tTBL35pPlIz1FlRwcMPIN85A
nA4l4Wqe/8Yzx/RhbmI27SS3DLB8i3PsRTZjNQUwlij9hSI6J+9YIb5QqXsvppio
Voby8tt4wLMDh1J7QdeTBQ8km8JvQ+7tqgeK+odFfWAiiYt65hVo0KZ/DUHHebKT
US3H1uuaK3slcJyEADgruylCTOWpnSmQo6Z7akioaehEzpb0w6rMgH4Z2c/Y/fTI
uKLfZA+5ixFR7tsQlpeRfwvNYeqK2sTCwGplJPGdW8P/DD13DvYd4frqHUXMER+W
aD3tdyW5tYQHn5NVbfqKzeglg+Dn+E/lIL04+LS4PtXFFOWNRfnB7jJwilNBLBqN
b8zd1kQLXXylDeTshQphKJuZawH/+g+CTUMK5BwcVtZ/pvIYZtApQtAyBuFoGZjb
XYmbFfYuaC764rOJgBrOqPoNySyqIHxhzQrQXtwkzN0vDbGR0gVpqEg7N0BntovK
BUU/FNuFas+U3Hnk/XEb/ucuWyO2mgZ6a3gYVHgXl4JppYRfBRlWQSxzC0TyEHBL
/U8P3dd1cmh3uuSHbqwE/D28PUnv3clJki0lEkDSeMPxBXIwIibEGV6qnLPYqgz/
gMBia9EmYR0+cjDFESlPD9bs/JFh005JU5a7xX78qGXBgaBrWnKvJLHOay44ne4Y
isrmcmaQdiH3RWXPDVFkBMUn19Exzspar2GCFW3LHjh8a8tBWxM065Fyxa0Ws1W2
zmoCtTr5VGir4beBqAEMTvixhf+rJAMTXMVz1cRp2Q1QPXkLMwUuJ/ZrBKf8Ud9d
e4rswlgIt4oRsnOtiqCNA6J/8E2//2TkfKrCUSQl6iRA/Rjzw6dni/RWSCcFvxPa
tcnl/eD/3SIMxq37pVvHV9/hNEF2NozhNCUNunadbSY+BDmdaUvxsOx+bsG7FaGO
EpdcIZkVq5zmcKRyPTYFySIpKTUw8umvqpmRfek+VnPfsAswe1Q+DZnrdJQA2GjM
+57sGsTtjAcvu99rX1udXzlqtnGxGnUrlCcX1qKmp1YOO+55BvQVvU5/6xGmAIpI
ZQNAvL9vV4fNWUFXGyQRVA0mGI+3kA5H8VitV9O2v8CkQJsgXKL44lWVzaL2QuvC
5kmRPpL6V5L0paLcWmjFqHCACjj+lYcD0zTr+E09JneT7UtBEWrr3zvdJUyZuj6u
3eC26RPA8z65NHCSNw4/fs6srdrbEN4BfgbxpwrSHrL9yNVD1lg7YSzsBXwNxe0F
5xwJBUGcsRRrt6ATC9atz6SmmOK0N5/psG4aw0EJxu1so4WupBSKP6aQOE9PiPJx
1d5ISS/8GscW4cpBUkrAdhUeSLb612Fy+eAL03iD5lVtIWnrb/niQOrUcbKhIOOc
ZmJyff9moIpnp6XB81sN9vrJ0WOo/xpwOxOkOF2VI1ZPpEEm/XIK5wu/tn97/WB5
0gLKtJq1DpymYU+EsmHhhC3NENG84HaFm4Ey/FRdFikw+4r2R3CV7+i67Fl1gKiG
xNeHogxUcl4rOnSlA7pyK39oMDgLKN4EE/zMbmrht4ZOAYd0CO7Zs/1yNg68Pfv+
k9KIrRlv28AFDxepuGCRFrkLHRiXs3ZyjIFTUH0FumTbW3LIAc3ymcz9oWJLbO3U
LXEaqj3mpJHDeJbTSa84wI/tX5EnEhiOaLvEYTXLkh5whd/7f8UgJy/XCEi21cZy
OyScFAajbWC6fxURYSiYxansJydYeX+BMtvyR41GvZRrd1jcPqVWNbd0u7FIPfsB
O9zOSUvdgpBBZ13s4I9ARQwwPYKhyUBCW/CT39oBx6o5rdXgLslpm6sUTNO6q90k
ND4VC+HW8vbudJ0IJo4ayziiMOI56gfF6f84gf5/Yjsn9bmgHW7cJcz3iV/lbYgl
CQnK7oYDYyYzZHp/5N7vQBdpRNt34BzbUxWQl8z/xldT7I989EnH7HlDk5oqs0DE
d021ex8AYuDwsPR/zG0pXBzqiywjpinhO7mSSj8/ZsBpq8hKooAoh1vSuDK0nXiP
UspMIFGE5FjRy56olndvzWl+5Bg8+LHVb5APavSqlWzB88lHuvmnt566KnoqI/2j
sEPVGBRZI449F93n9lM+0yT8epKG66qxAfPdg1PyNSwfRl8ufmdNxVl5dNlNbDnW
vAdqQhbGeVowbK/X8rgct35QiPxOtxDkRAQ6mx4oQxxv/Wg6hazX6AGVkdnpZMeT
+smPTZy0LBRyr7DEP86wBafJMj/2whZlsFWlr637k6+Y9iD+Dg7dfGkgMAxeeYE9
LSSsYs6iKdMLspDZroxPU+fHweDeEYXw73CS9CAZf5Q9jG+NUXls20+CojS2WPRz
AAGlSPSrpnT0m5VkWCKYe/TvGkCajKA0JFpZ9/eMRRr9MS6PxqpHZCBsgMEzCnS2
WFp5plve4aPqiFnXIppnq6MZckoFm8/EG5hYWif6tDZQMcZwBXgn8Q25cNOLBvP9
NCZIs+xxeaWu8SORCWLCUDTF65LKT2sPPeT9Xw7VInZNi3JoYlk1R1CVjQ+7Yt36
4vCt6kymN+V0YQVZGJrgjwrAl5pAvs4Q4JLbTjaCX3Ndnmw0/Rh9GCvvAioijCHK
Tzrma/Iew/yzQpasOIdBcVfY3KiQvxqwYExv7Albzn0wQRL01Hp6dhXwVfpQrVw3
Pd31utq63UYbJtr4Eg5k9EZeoT5VyET7a6rVUZVtG2OUUFrn+wJ9sogb1MKR1BkU
nHsNikEpN6Kq2az2CkFmcWl4Of9SfKJsWx8NJsndpnGCCgvBLvzTbPfs+8yLQ/Qp
XsAEoHqeW9QOGHS0pn18UMiZgwV+xuH/siqjVOLiKT85Sue7cYCf+Sm8wtKKW8WY
P4iKT+SvFl0J9y5HBtSEHEmaUq9m6yILhfyP2UQcCl19P2PMEJznJFoKIX+MpGJ9
d+KqLTxDYjKcNCnaegFRTKJYPKlQSmnexKQ/eQQ/S6cZ9dT37P3OONGbi+gIE4kT
wHk+SOQEL3q8p7jtlSmuJB3RjoK5OEOi2MmGzUITzmlHAtCKoGZ7h/UDqPC4STfu
TrXwd2a4+70+9M/Ip64i0eJESMuI1/4L13R7X5/248MxHtzmH4h+MveyavALXLty
zouh9oHctMa/3WgBhsUbWaMoZd7ZVfZ2gkIjgpf/B+nVLHEGYP7Uh+bFM4+32wdm
9dwSN8abv61KX0au9lgdceSfy8hYOSNXGAeBumYN24VRSEqTs7og8HA78MlVl7la
WaftUZDT0v7gcR3k1McZEzx8TxiJ8ycSkYWOSmvXnWqM2R7me8av/MEXcRfWgAuk
q+U/UwLoB1s2sOfGgLm44c7jraA1IKi9tt8EAK32i0pox8BYxSCdsWOHPrTAtgZ6
vlR7JU+BPZ8KNiWhbVXNV1Y24FlJphugaCjcwoafxBwQ0JEXrYj/e1EhPwTq9Qor
Y9jNHO09V9zT1ktGm9Rlt6Og2huvE12aWxQj5x6XT5W3zMDlaGWuFiicDXWOGMCF
x/n947i1zTIw129PZmkxJQ4bj6DXKTPpscEtG3rmtCdeUPu70mqEhBWS06PHaZ8S
ope7iZD8uPdfsHIXI0yEbtFoPN9nKTTkvIM4Nqv3oLAvyv7EalsbsTI5xnPkmuNX
rhvr3WCwC7rA+JMBqyPz29OBpB735dw01uXAokqUev75VHBbB351XbwD9umUDVWC
bEGH6IqDHKHBS/ImV40h3fCj5EvdJFboS/Mj25uZuW1o2JJoeB8231DdcJgQzPtr
0hJ2GyznJQNZY49UlsPC5ooO+mG604Utaba62iHlwe3BWYH/b3ccbNw924VX0WX5
GoUvALB/czIfy1KpujRN3FfuFCvn0ZNJ8p112tH2j1O3yF8p8R/O3C6QeIzzTqA8
J7a6HnLoan+YNYDoIWa/cjtCrBWc/Qe374TKVJeUwdnBeex2gLLIjCEaZaah8zJy
h02Lg1q3ajZ8HFHVTVY6WzqcMmiGDD7zNNNTpIl9FpALjTMLT9i9UOt0pSPqOGnq
hpMDdtzmFSpBcH5xw2L/9FaZq1eiqUqIYzg7nLf7PmuEsBlxgayjFj3ReYe20UL5
uEoHMGR9Y286zdJ4rYlaXOT1KeW0LUCbhLePzxJ19iwP6wILMNgrVsg7d/GTNhcb
xqW+XPR8iX5EKlwq8Twn4xURpHeGXWovZSVmCl/1BXACkTaRjMu1WpGPTfS57yVQ
IrUVV7gJ3kkhePPPz/axoBHa1IZgZKSU0lOgEQx0BZ6R49xo1Fdgkc0dDwW39IuZ
QaUS0/USqPH7D5Nhg5WPo4e9sBDcalEhRCXp7mO/kiPTK8Zt7UZmx5hHKRp05zUc
hf+6bFHVPs+wgHX/YCU27HyBU0SaR3qNEYPDfrR9L7R8wwFwUObxvH3sZAiLmH8X
OxwjSV6DHS3fnFUPSYjJ+k3cjaYyBqNBwlOsWuAmx/hbR45YI5TyE/14wcije0Qr
35vsm/Fjyr79lN9BkU/kYk0HcKyWQYkfn6Fy5KyrXT0qYgFMWEKRg8YMyBWTOTJc
rnvsxramwJO/cpvtFfj6MSbjFF7UQH06Ih4S4XyhgxeXxl+ihw2oZzLMWHH4/Or7
KVgjxgibZUPW2alELw/arjs6Lsm7vRbNk+5apUR9D+tPpyJfMS1VQyyqcsYdGuSB
kOWJwyfyKaauVq64AFHXpeU6DMDqk2xUyC1dsSJHPoElMXyGZqHVbV6KwLym3D8D
0TvUiF422ucfp9/XW20b90KWlsrhfVXY2quEmQr8nak7X4OSyTKR6f2a0LGFnmQ4
QkdJ3cTpWIhofSLP+iSEPDal0d95skdO/L7rKBLdQTHgzMyGeU7zFs+A+6/G7XV8
/7RHKYVfPHIUWKXb2p+ymy+Vb/ziIcrBb9Yhxwd/qMbW1osWnx3PWtN/nngYs4Dx
G4B1UrefVPZ6CdiuAnhcrEzlWkyfXw4yYMMkXqz3JWRowSiTrERC0W/rCvn3uYhR
Ed6DWW6AahhRW+iyMOYdRnB3k3mS+7D3UtGQ048l8cfZvlWuv+XijQ6NQaLEDBov
2+fpYkPN1jLgmwQksA2pm8enRWW0Xc24TQQqxwxfd6qoYimQDP38Fobby1P1W12/
YL8NiuooR39Eq6hp4zihC1AZyhAAJeUAf1Y7IO7+r8nuDfPZWwS0clHNs0xrjCi0
+anYsm9P/UulV9UdFeSFswkBMoykuGSLqS0rSsm4BPtYl77IpU9jHyM/HZ/Ge6eq
iChIXde4F1FfwvtuqeSY7oBsrTsROh3jeDYRtgJC54zMmCcUJiGaibN+SFsyDtMA
YqqRIMh975r4G3B17pS/tbpCHTKl9oNyiM5OK2fl1HeeXIHEkTkmSwdVLSgBzWjA
tl3jve4ilNeyvQ0WkjNqwM/TkxufJFI3BVYwfJIdPIdBUrUGXyRul6wLNDK4Kcgy
60FKnc3P9A7KQHmJHmJiigLhCLPIc9TxGtnJXcjGTDvajW7Eq2a1aaTmFEhzx876
zb71grh+ZmZGlPpWT4L8932nHbUSceNaOqDKiOrb2dEBD1jxalYMAjkcojO4iRT0
8oY4NGvGV5+KtTOcYqBiV8m/ejhDDVWVv1HfK9wqk7Mbmh8JYxmcPhJbNZWW9nC5
YLmcIRvdp2zUzlrYZ8fnK54D8SZnXOQKzJ8SmF4TMYcerMBlM44CQyM3vbtgvaM9
DieAwvRAc2peruiTOB/e37/2AK2e16KYL+Ba3AQu0Bsq8bCazKD3AEHPSyRWeoJX
arHAnUS6JtYOk1Ne82zbwKpFppOsfknZzu1T1BFZ4Ijmjz+yS2Bum5xtscle0TAw
jg8c9+Y3qlpwmHHRDS1bWDV1NLAwby9etWuwDv4S46KYZPq7WOJvhMs5bvviI1ai
50lkpD5VMYMy/2POq6IhBxPIJD3CpdtkzSkTNXzldTOiqhWE8kN5UgnQl9M5kbry
RaTcxe3FhKFE7iXg4Z5XZmhl8NP/+jjRYVAiuoKoiRCUEJnxou9QEItE+ePgFz7C
65pzcNAJjT+0mcLegJd4Aa2VuACa/xrfLHGjYPetGWWC4kPPWwQ0dugA3rEgX2or
JtP+u7UHGGIF7giXj74m2yK7q4LG+u9WBw7edxv6we2XIxTGmSI+nCo4EGbwF/z4
xy48qoR/uVLndHj0AEC0HFLiOmiYdkd4lLAKEevVixLiF11LAPmZ90l6J6j/X5t7
sAQ7AfbAZ7YLtiGj/1+QERRxV3BzKQOERtMFiBfgxvFahYNa8vyJX62lzJYad8Et
eivvew4Fwt3PNY39g3rsh2RlCVZ7+x3CvHI5d3u1FO31eBOwHO0QgZYV/wmn9xKT
Sn6o6sGolc2x/yBJSVFk/NbKcsC2pM7v1liHwMz4HMQ3BOMBwPQi8BMT71+gtuNi
WIKucaFAlkOL1t1mk0ysejq0W9Ay7WOE/fi54ihXmpri7H7c8Pye5sgoSaJ3kmKE
gxOXnxpeYlnOHzW/35sT8GQ3Z0M/vSCmlD3X69S387zyX+AFGYs14VCL4E0Flzl5
FrqwzNBHUHP1Hy+FOTDSL/6tV3nXZDqViv1vW+ndSVYVZ48SMrjM0hGBE8/3kBOe
u1Fdf36m3Avs9vovhVinDxWtJCXaNC6e1gdCOm1yFpip5TAmky6C1koAZe1dXnZQ
W3Rm+DAY1cXAMWUbwdymSwH4+kjuqDl9njpOYUED2GRfRv6oMRTGzOvr9RI5x7iV
mk3Tz4aNuw45BAQ/Ib0S4hVZ2H3Kd+SiWNWpS4iR6zQ3L1zwTUGJ1VeFGqcoSnq+
BgNqHEQ3SR+KmtA1jw6tOza5JSwfcfaLOK7apXjyYWUhj4bQmSrhdzG/8Nluey1u
QXdCoZQzaiRVAk+iabm1MAmUjDtX5TDO2EeM33XZGP7uIMzRZi1NvroCOLUOITqd
y5X5g5Fh27275oNC+g755ce9S4/ulVKt7uzQ3BVKXqoc/uOBrGlSaJr3buR+8vgJ
XDBkvXtLqpN6KzYuhb/+bCHsJkCf6dg0/UoqoXczVuvNxMi2SKB+F3tc31yHzQRm
GSzdQWVIvdsCvXYgq57owBwLzH2VZHe1eo1xK7q2k0ImxKtg99JKl//6mSXLrx5D
wqu6bP/OMcdJIGXWatQpxPmQgVLa/HXNWlUFvc0PnndrvpVwi3EV4/5bJFBbhQ57
ZQMPajL5R1nBr3D2BRyUAd/In+/7WlmUBlJf4H4pHo9U5NuM7X8KGQEkzpYNpLbs
9sex+k4O/tEFHpp/+U/PHNSJ6Vhl0Q12zSA6g8gJxkfrubiCSqHh4GVdlrcQRWZ3
SgR9dZezzJymWOzqlNOd+s/zT+992HIvN6DllYWEJIH2Tffadyqro3Fph33gPn6j
hHjvx2nYYAcox2ECWdefD7wmyeC90t41Be+8cioANRLRWVxRYjEZ1eTD5BrhZToD
39mLqrn5mN3IKqiEiYIZdnFv4wiZ6Qadu2UoOZ3q7TJN49aZqMufwEp13evZ09AM
5/P1zMiAmZBDc+/t2dfIeFksmd0ZtIOl4LqNlx7PUhXc357zfcv6P7G4LWvanTrA
1gdp4vWMKc50j2jn7EK6dFQ+7YO5jA+LRthFmySfxnjnDJrbEKw9Vc2bVWFrSu1N
LKEOJwi2LOhJnnRVA9drbPoZfiMb60to+LDYUETKO9KEgwWJ3qFpm9vMlMITJ5Dl
LlSYHm2s/rE4yFwnZEfi+BqcgYXBfntPw2GmK+LazBzJU1nhtPYt6arGCeqvIH27
oSxBrVPeM/+VdONEJ01YS+ZA+SEp/M5ITFGFbTvWgxJvvQ1C0tKPXYTgh4xlAiBv
+ECIk1UzvXiWvsf/Ln2SjJg/YE9X7DdaALn9JPVrx84afq2OzksZeLUDX4+0vWQ1
7PEydpx/QaaktaNkbB6tm0J6xSlqoWLmUg1g4kjjMkRqVCgG6Fpuo57saM/dL2Fm
aTO0140bt4iC0tozpaf0HVCGQskUAV4quFUJ1N8Ny0H+o4pJi3eogEGv+6sBofUA
gT97Jnv1DOYjOdC3jQDhLAYNRGebj9a6tgeMTDm7arjvPeg+OQPDhOvLv7lFRKTj
0i2G+QaOXERnhdzBfLNYfqcHm8nO9jtN3Deptob1xtFatARN7pU+L2iePdR437ew
qOBooiqUXrwu5dY+LH65HMvHT8y2I6BGbld7AVSEHvJMHawlOQbgjwqE2tMdkWkH
Qol2I7CZ/Ih0QOLNvWEjJGqs/Q0rx0wlelKfCXHoL2hXBl1J94uTwP97FfdVZjZV
J7TGdxxmbms2J/lwyVU3sl3G6nT9EXUblL7ippUDkfY0X4YjAFxzky2KoA6+7nxO
IL0SlaUbobjf/lFDAVh6lKft+Uju0KjYyR2EfjNS/FUKbskY4l1w8aY9MrRuZldj
JNJZEDa/cmslvgz1CdsIm0aRuLpPAvRHP3PdDdUXi5qWYX+eefg8bZ0+kafWOmDY
Xf/BrL5Rw/HJBgY8Ss2DNL0B2xtO1BHDCiWFIF6IeWKTg8SMBsuvSdIFCMoOU9CD
qR6j6aeFNWzJCDQS1vkn4cGkfKbjTKScGerU/z4c52F4gk9vweP19PNiCOr9MW6G
rg5EycfGZjn80BZLgRpTe0hSOhBxQQpy01PHwwdWkzWS/CfI+Bpef7balAcFjJ8Y
dkvJR0gxQDEUaR0YN3gg+6/OKavZAiJdUILMp2CicJdxoILebqC89TuyXTSQXcRg
IMHYZq5WKJePAFSS2746WffJpMHD/Th7ePiDmJhnpnvHBZot0Y/gncDln+oiWfMq
NvEUOav2daJrkPAX3eT+oLJqyfcDk8J7j9QBSCsAz9Nx4gELXXiOLJ1lG3alROiO
BgCMRbF4EBmVkM6LnBHQi8zo0La2JomIMxOKpxK2VIEXcpTvNY11nUkyTgmY1qtO
d/EICNS65UvuBA/0b/dnffFc72g96dRYBdTtjn+0NgOupIHe83m7iXuopwpMnZt6
SkrcmedQUNg9LzRAic5D3O06y2z5Zny/RwmthYzezQyMtOW5ZRI0xxQqTf78W2cx
CVq4Pmu3ib0IwZiK3OIoGOJlNHkwp5ciWQHIXLWsRuG9srA9L833kU+DZ/41WdiQ
3IcXYWcDibsmiOwGiNXrU+idUytO4Ee7r4rrUpIvHHriI1KHRLCKEDB9G/fKxvFm
/M+g66YXvnD0e/OmFui1gHY60ZTvv/XSWEHhFcX9K+XVoXy9QQPUaltWrzrB+g8E
FhiX6MI82Bpu8dibgm879J89UBI3xmYk3imxjI3z9B9h9DsVbGv6S+xhwhFLLKzZ
FgWIJ5fwCf3EWGZy0mwhn4hW0DfBOg7EAdUzRboCz8k0oinY4wKYJWeaX0vs6rGo
hXpXerJon0TI0P9kBixi/Fkd3Nx/XTQB0SK51B3XdGKdcYKUPaRz7H8C+OHV9S77
TYg/JkvwiXfwrEgf0euQzeAFbwlD0z0IrX2yOItF6+EOprdgvCe0V6Ob3rGBFii+
uffJz0QMbYMOwZkgl1QNdLsGO+Wftptd2pBWAXgBpyIeM900fpKrnbU060dOXpdt
Ydkj/nUoRDmfXBhG9zViQIzc7zZlTLV8iNx5Eui51GpacfY9gez2qO3EolrvG4DR
nWCXa+sZlUyIoBrhNm0L4XZC4yHTrYG/J2ojORlAByrS30OSzvRXx3j48FtFkzmW
cUA4QceGRBr3KFx+5ruRXuy3eX+P0PnZnrDuFNdu35P5qCvurR740PN27BlvcsLl
eP7xbtP67PfDEfubR+1F0mkegdXA8PWaRsXOuK5Kc6lixT1rqEROYFrv3J5HnOU7
X+wbImmhZAKkYENgAD+nMEFKY6LJ2QbJMdWvH4bqPBgDBpQGQyGzcRP1CyqrVCR0
lPYmQrP3zfMU+EO26xk7UCutSKPbQxyhNCD0oM1Lq6WyUH37AP5xQUaC2XSF2RY7
VwS6EUVJOGhkLUx/lkvB6HfiDqful0/KisGfr0h/gAJsLhfECCmvwCxt2KnVq7dX
jfbSmGAlri6G4MLMTytydpjvEZQFzFDBn9JD5B0LETw/v+Y6tMwHA5Bjcqrnn0/1
+G2usjlTyhupffvfacrMQyDlPnPTAd7v9pgAUyhuje0uMLvofWOLRmggAwpedO2p
TF8L28aa6UMQTDT42AdmGbAz8P5VJCkT0iHj80ZHhUNikY2CzO8TsukJ8TRRazCc
1flWy9l/KuhjlW4f+sBeyR/OkT8l9CZEieIM2X8wvKSW/13dr6n5nHvD4MOTfz+X
CP84d3ccFR5dY1l11JCkAJQbYEIVltudp5WHmiRC1UqMgFebTaZL7Zylp+tNDhEm
fluePw4HOdlcKWh+8oth4oWldj2KGrkk3rUh/ATz53gZv/fHfzfZWCXtrpfPdMHY
U+iYHeEfrUBVefciuKT/3DpNhmdA8QxaodWsPUGFvW4BXalRXGd8GPcvkYviCzBP
BqKDxtoXV6T1+TOiaaPWYJvQb7pzS82nXow5Ld4M9jXrHQN3lx6HAvbbOzqwoRW0
E8FtCqbVAl9Ow00RDW20OrbcEhdpadTLCRiFsx92tHtKnlzlikSd3We/oUp2FnEn
ovUSXWCPehhrHimxG05C7ihtHtU/eC3Wq/+tN5w5S4Yhhp17Gnguv6cGBq+sOldz
OOR3m6dUFzSFbGXzO4nD291ULMeTG7sjdTyXPkB2ST3lQpmp6EmrWwz7GP3i+ndZ
lvLZCSlxacRd0AMc1fR18pbMhq558PbgKWKR6vhE9nnXICaGaXavRh3/Td9EJzA+
T+61P8M0VE8hm5AipHX7wTWXp8xZeNoQogTXE5J03NP+t3cUissGM99Z3kRgmvYV
yHLnV5XE2ACIc1407V5XWLCGKB1pGzOiL9V+9HRQuLyZyGga5ldfRExag/YOZaAD
7qvas1zKeV+u4DTe8j2BUSxCHV2bNrrTm3oV2bCaGbpdMVGH8QPFfIl6XsHn888k
V2X4Q0ezrdDJQPnehssAbYiAjzUc3y71zBiZoeEYJgyb1fPsH4FUkwYUnVu8xlkq
ZR3Krkq99PCUzDRFiLIwY+i7B6zWZRK8FuSeHFrvWyrW+hAMQY866WlCjYmP+TbB
Y6CwZPUzpv8rLyE76L1E7LDdJmmYIQszoiUFiw2YUPwNlMbuuxeNM8JT9lIcMz6H
0PvovWz1JuFkooPjF0M0BMCe2yqYJ61e4yJiWjSczLaSz3U/DnQZS8hOxzcSBJ40
84kV79X28/LCA1d0S0MlJiRIcbFSHuyDAHxzkUlDkA8we0TQban6lYG7moWVRJ49
/2qSdjoSAuX3p3V0WGIn+/qK2+gD0I92YLmkJv+3tXEKqT30nX+ysicYs6/CGUJs
InTDp/96QRMOuCP8e7BWYMRCrtt5PbKZ1EFOBEfNX31EUhB4ZcwG5xWpPd063Ted
pb/OR/nSVtDP9UIzwdQI2B+7isUfsVwcBnWjrHFUR4e1lK+WuZgJxAjpuvpuFh3Z
sFGDr9T+xX4Zkj9xos4PYdUbj53NjUO/P+/IBaAF5TrBZg6ze/FufCJTFTJY0JVJ
dYi7Qm/ExdI0u3V2t6idqq6zX/MRwlxoYcA4R9HHOTLEhhnQWXvXDfSaCj869weD
weCH2cOIuox1pF+0ajp6pu3/WCmyFrPkF2dUOgEvUhZsJQG/KLr8BBUEXwIZbKY2
qad9f1bLhiP3sv+qpEib6vAXY6A56GpEkpltvCOq2FVL9MQYUemzI+XFHZiC54Kn
XMPEokm++THO6NYffrRGYlK57O1uYTzgVSf6neytojQVwISi2rhqJCTSWtV5O6aq
FnTohsk2QCVqfrTZJeLSE15RoXN9cX6ZFqsD/O4JUzahkeFtaoqHsZHCEpW8m77+
xRebXtJXANGdGbAQdPmr4rpFq3QCrSCYjwHiM53X9SpFHPG3aj+aTs9gPcj5XdNo
N+eiwepHuUTYNd0HZMqj+5D+aItyHhmipoAhAIsejvD+Rq2hAQR5tOVwoF+1mLaq
7tOpTtMfjkYfs8GpggDD9nwTlyp8KWSEIJrEfYaUZ1ml22BmQqv18PlCY1UoZ41B
aDiETpvGnemaRFt5Nd73nYbul+0oVEOZedr1XOkaXosmRaOFGdHW6y2iV7wPRUlj
EZHHYRd8YYknROuNrCHA1gHHCFCwkWb2dxUdLJg3R7isAloAQh8t5xAxNBbzo2uQ
vsQn/AnDOJ+GvaeXWovZo328R34tMVLbZhVAvPQO9qJJwX0pag5KB4u8QPXvvuNA
BIaVusPYdQbrkd8Of0lbF10ukgmQc4h9QQSuxqlBhlyZDKrzAnl1FLgu+viF33ly
KTSwHkbCapGvCUtwIR03Fobec25afOH5eWu9V0qZRPGFPSZUbLx8dx2wcNmo9LR3
TpXaCJbIwvtbOaTCmERO0t6aT/A+rD3l/V3y5TbG5+PMTIfnvIQMKHijezt+W+za
QcXgKf2V5Rfl1dyA1NXTXBfbR7t5U4kmzrUsTnG5wHQOcgtmr418DKVwmtjnKFPP
VE5qjRRSwu9o6Htaa4dmaYFLRY59VB8+MeMUMH+lZ+s1zIth9jfpP7L6vPzABrcw
juBXKn/DibuhaDWE8MsLvDNAnahsNs/yomIy4I9jO1UTFKJ2l3fjcN4zb4w1MwI8
WVeY5BFAskvFbuX1Tw4IpOwEbRRWzJimGgVTdAORSgrjMEvfaU0Kgouoh90g+UK8
2fj7zGhU1WdteYs8hHBwzpGaaUvA+BSzm2vFbLX12hZB4fKVpGV3pEhPdzBVj8EG
OePexDP5QJ5DBBAQXcfpg5N4bleTYFKiv3uwFVqWoMqTatRbTAKT5hkEKcb2+QyG
IBIeHBZ7/pt7GeicjbXWHav5DuOi3uYreB6wL5ZVwuhrXD6uQu3dhsL+Kpn34Abz
oyy3lEhzKdvCO1x/cWaMoVmV31OgPp2wNrLSl5tM0qKCduMB2wCRdjPM1oHOov1L
jKPKZG2O4QyWajmS4czLhwO/UTmkhqYaKHPuIeJp55xub7DvQXForcSnubpHJA9N
5DAwxDjidqYW7+yR9LH+XusjRh/F6Iq7fefjc4/jITfdyUbPhZW5GllVNI7ARbEF
o+rnkfLyjddaYTvT5GLVZyEW3MH8pcNYVKI2WqTCKYizVkourQVVRtjiDKi/8FDk
li0HhXxpgrMQYh6iRTP7M21+nuwtSx1IcY9b6NLFjcHjSCa6segBOUCYKczDOIc6
dgBtWoSmM+sWWoFRGg1g9l81VcJUCvGKwo+48YnNZAeDNqxXdH3djaMbnehAdDHB
t/GwYmk60JtzCuWwnckQrWxxbSw+BgcijPbnmUhQ8z3AaCbNMCYtrE+d+toKGHOS
R+x6KHUvaa93crNVxSzOoz74axo8ptRIeXI+g1NrsZsng5pWbP9INOvfBYBfDVD2
+63Px04Y2ornSFekDUu92S8SGtb1ij/L2i39hh4qmoTLpfeQJ04RY/pzfVYYBBB3
62P4BL1/OMJI+y5bg9g/zNm+fk2YyQsQAQYraNa0IUTuqd/u5B8+AYyr3CRY9aBv
tAKST0mz28TNn98lvIx1Z6iNXFA4Nwy74e2JXV+vCiIBcoiHxq6c2Jdmwl9tIcsX
G1bCa7/6Akru8gf6GDYxvsf7WyAa4Mc/0pXw4sV0w7+HEflnnEvK3PRt63CGW+Ow
48QX+HX/cjtN3V3PuZxS8HIAvY/exsb4/wXnUWwBtMLx3x0mmFEmnkYJu03vwhdb
WQsTmLyIHc9RvqmjUmorRbAXV59MuoDb2p8//jTqBTpazX9RESUx2WDwmZRQQ3aK
Tom8ypfxrEMObZuuhdLoer3TVX7otvup+RIjn1zrcdRCGnyrIYhPDdyQyFMZc6wc
7c0EMaNh9sK4bys8zchaYUid/Cz7znSquRpgxA4wB4Ib7XaV80pYrlxbIsKtDJ4A
pDbOLWKxoBFwXrhZzCWOR35XmC/qHWI5TT2VVH8yD8muZ5fklaFijBaulbfQvkNO
1FwYuAqkzo3gLsOmM23m+aeFJV2YM86gdCZdGU+MoYTkY9gLPqndd/TiaKz6Ltk9
blYnrxd3nk/LG9yh7GcNaLi7DIr/T9icHOSWfDESo0faxiAbsVqoDNJ8IoFFk/Fx
fav2WBc2K8o40yJAlDpn4G0q11G3W832ubPLziQT0iDhENppRkE5aVQZStGTU6iQ
1FQkT429/L+GNYy7XMGKdkEEBf0CBqZfYt88plxlYtWeBMpJaLZ9yrxv76c0wgPV
S+Rw7Lx1e9Rfn+YulEjjB5oFK2R59kHai7HWpVIibL7pjwrvNvZjQvHgdbVCNFCA
PxcC6f+HbbLJreS7FwV3tRUVl/Sb3OZV6LhG4D3boibXjYQmCvZgKWDpjcDUf/Kc
V/b/p8byWUpoeWMkc/bblxFa+00IEQG4oxk/zGTaIP7g4LYzqPHiTfKwmcbvvi8+
C7Id6wNlYQr1iwLkeT4i5Pz5/KiPhWKqYpaowZVah6M8nZoXuugbHPcfjxgvw/hr
/IiosM1YjvC2h2jW4oCaJQ8Y+QRO2UYkMXSOyP8Q/Tmps1xA2OsVbdmnmy7YO3he
ow+5TpNTLL4fzEp8SzUaHzbJYUHFda6C6gw2+05FHOjrmVdvKmd6C5VFBjMdfgrT
qVc06w4oGoUGa+fwvGOVaRn7+Plrzg7dynFZ+dGnwdaeJi0drWm4eP0pxOSAseWb
omHOx8/gXVFugv673M2fyeOPwssYmYGJOxz+ojEvbTTYg3s5EqnJ8dKT6owlBkOZ
XoP45wbk+cH7dWTeJ40zlKRWKyk6wM5ou6TnhQuf2WAXt2NOOEMICfYCRxIulWAV
9v44biUZKIGYmSrZc/I6FomfwliNvj6K0sJTmvg177djNeiexIFv+w5GrQY78/z3
nzo1x8TLzeKGP2nQFBSFNwYgHdYn9hQdJEGeoNO5c7sIhrO4nbJnjB7KsBMlm28T
hvbH4vtZh6aawBzVzcxO6ByNy4WbT7hPKkaRPA8IfFFGHafnUcdhy4cbY+S3Y9Ax
WBEwT7CTKaC69fNmAOo6MJDOYDAQAj2/+JGHCa2swY3HNfUmOBa0XEPm38KhHa07
1QWTQLPcobnhZ+kGO4UnGP03n8C+zMOhSmCFtIYg9O3u0/cjcFee2Fm1vN4NdJyD
09ojbo7xkyvxRJhhKOomJqIHCrYS642+RNgFqBHPUcjdjPJDXs83/yrT5vIDSkYo
f7V5OHk0smxBfmjdg5yMrUyUdgmRJY16egCXNLbwxKbXyakul/6na4CdK05WG4yz
JDOfVYSKfIn22yM0WpBt0VUYCe2qM/M6jHUr/LUsMTGPdAlo8ZzdWKRB5m28Y+5Q
+f+BRvVRjJVyeCijJKvy0aT+oHpt0JtMg7jKPZU+GRQ4qnn7koJh9y3DaS/GWKIC
+9tNpGqrRS97p3mAOHrWyCZgh9Ls5Wm6i2CY0y3z9UKOsa1oXKXDjIrnBT7UTDVN
5qz/7Rvy+wa8IOu3cy9XYtohncVBcTPsSaMtASGhkFPcB8ZM9uiVoSypc2yElh7u
FMbMup/bITCI5XaBnca7AS+eZ3KEn/2grAv8nbnfnlxPis6kfNYizxCMDRmu0NO7
w0hGYncVyR3eKYO1tv6PiYxGnAjP8umdSWFa7Nd7YdHEfG0w1BkoVDEHa5z0hwyj
cJRp3Du+DatJcK0Vuv37/cDIcev0a/FaLAU8LG/YrurCmziu3X3l54CCT8dKL9Ed
5LV4jW+o5yLWFeZzuQFYjaj2RUtvbXYz1+OQ+e7lZvl24FRGb8d4rRiu6x1bYIHt
RMT/H0tNHtyDiExPCAd9FLO9ry+rdncg3J+fDkQ76eJ/dWDVKICjKqPtQDquImV5
64YS3CC2uzwKaoisRH/rHoVtcIj+VPlxheow74FnEjGwmAlyTI2lCNrTq2NGuhNL
NYPO+hRcPkAcQ3GcC4AjEcvL1hQEuYN3YLByOTpzd8Se3wXBAq5bsGkSyCPC27qK
zvs3nWe/vGnWMpICJFBBuZZgAhOk1jzzBMAd/Kpui7VTQ7x9NHTm0f1ppu5F53iB
2h9E7SWQ5CGZ2WfgGd/at5nZJuytuZA59QU1ISmAEQb0pVO8zbbiRQ4Djkr8QK7g
GBn1cNX8rG3XbFSzL2qG2VZ+r4v2Wz84lsN7XgE7nJX9QVqkOgSbzxiux2ScSv8O
Ro99dy0yDWxJmIJC4ok1nLLocag2j1qLFQXB3F8UiYws+xthxWz6yslLbZ0Qslef
tbr57ULMzFrKdNvFYxYYG8Nr2T9TAhjoVD30FlPecamNvJVGtvq8sfPX4WBRhpIQ
AIU3ISOKu+5b62OmtxqydOu5xLFieH1BmI07EsWvmZRYfIuQb70tvl9raEbxNkrc
Paj6XiLcDaiYZt0RblvS2MptkviDK1546Z765q0cJBkHgV4BW/oxIPUgF7YZqMul
LSf9wjkOIeCj7DzQFUgKSzg1LznUYXexsfuHSJs7mLd/Zl+zGKAnHEbX3BqH7iSI
ORKbJFyalk7qZEnzss3ydKSRoLaydoKvi+kLIp3d4dHhIDGYtFcRwutXYOKvW2GH
8/lyCx9CVTSGYY7F8g/Kjqo9UlcRAjJIGZje6BJ7qDPbjh404cCa7avLaGVewT4T
kSP4LOYgg6jhQPkZ6BnBewBe85k821kIscPys7ecPH3s8LdZbp50mor6EkZsqe85
zp86Y1lRZipGg+OOshcQoPm91SFJRh3guhO0l4tkRIGaB/PQcyLd/673+WGqnPDq
WnxON1QdGGE7ZaH5/laMRu+W8KzO7PsdOoNgZHOYXHzY9Mq4WUJsfnfmthAqFo35
JUxxksq4QSIMfErfPosTcL8Js0ZgUcKNNGPJi60R3R8eaCGqvkDkDn0A8Sn80MAL
zy6nmP6u8c3WZrkTpi3qLGcdh7vRqXLkfe3T4iz8Rard19PRwAXutPwJjAY2ugzY
fxq1l0afcKQ84Xd24KwrGxzfPbIIc36eNsKtRG0DdGI60HdL2kv7Xwf6ipZXpsD8
yfC6ZYphF1uNTfNxowPMMvbWCBqMn3swG9P9YYAgu6L4oiLzFfR54uejqovdi849
sxPnRE9RsDr/k1sWycQsAkcfmMgv0rehwLxCNQkmRdDjsQaLXyo2ArYgXzVZM+Fj
VZgAjNCNFgbrWPkbpGgZyax5YbhZyJH/j75tQmDz59tew2ZAbFFMvBSbbx7zDq+K
7FMs5+dNwkYuBiNnf984X7MTGQhrDW1EziG2h1uvAJE3uxOfjDAjf1HL2HBaJstN
vFLjx2bfBUZVRoKxp8Q/JefLK0g4MlJwTTwr8BIc7+m4VeTqOzR+4SyZAgoYjP7q
8RzUEvnDycmt9GIp41AQeZR7r9eLc8S2IfolRr8BmiGLoyI1V3UsgB6P0+A6Je0m
yPci8e4NRar+t/5f07m/kTAU2NthQG7AJCuwOeWmGhdGkr5qi1HjJhyrWDMyyVnU
+DjotiGM+4NVa9C0DGFpYBjmd9NatoJ6o77+n6u5H5q2FnUNWwID/77rze9zL7t+
cB3BYIq/zKf0WbS9LRkNIPIZ4CyxlKFmp6Ha9YbPt79I4aW6hEeZ0qI4yFpmhgn1
JmebH6aa+WhbHAbb8kpCh/ctefAc5lnHba8SwZeTsQ7skTXcUUrJORpBOaLksC91
pK8ndjqgSnKnvNr1phOxUUI62ifLCQfZp+JEgivFJG/q80oBjrS5w75phgKgNCqb
269xx66BbtNHMdCxubz5+zdCzXX48uzrtxoerukztv9v+jeFwlZHFuM8wNgPf9I2
HAji47ORlikJJFsF1NGcMHRxXPEdJj3zk9aRKKuroz9aYS51XNpB41DGeADCUUNv
LH8XJ5oA77c+eCXmBzP1uACVk+feBz2r1DPvlE+NCw1Cn1gdfejHHkr0x8kxEHQD
+JmRU70wdqUHFvEVXLfkqPPMsplpMy+A7uI+/EcrqKFViX0b5fG66PflHN2SSq7f
1D0jrBHgbJuSnZeTL+Wn+tOuIljrTVTUxyWtAaYZ7XFFceAZgcPz/9g2CNO+5Ii5
xcbbsX7qB5P08qmTfJlsN8jCFOLvu3TH0wLik2WwLlIcBl5hVWxA+82ExilKWNjD
qjhOgJ77MU2gSbT5z4YHOOocEdakDNyWFsw6RSSWeQbwFn0l771bWWcbzQxtTSiB
zcqIwnNUEBmrvNnu24YrwBMfOdxhpDbSCJUXyKUuyus3pSVPvlOQM9LchCecW4Yi
tWMPeg1j7FH8ljOsJGaKUgv8hvxq9OAyYheZehuG3+z0Ol2Ju64Uvx7GgComrVai
lwyqTx/IErvJL9TKCyAnUAHUIxO6j8aFyL8fhYz76uoDR3gc03OBWU4MhlLr/XUj
agY05g24QThUENCPAMCNiFM47vV7qgumxMFdm3XG5Zrfyk4MeC880rCc7M/NGQXB
qdDXcqxgXWkgYn8yVZyXhNpYZ6ZfjHSiApt9vibjSqLNr/pMZSQPtZtwMdWCNvnE
NhetBsfNEPxnYBRqE3fkq5tHHxqLA3u4GiQHKv1wdZJaSHPHX2p2NWSf9QSHAzSS
cLBcmmIp2SYfwkxK5KHsJV5+ypGF2CVBLzUbvAKQLuZYn9LZqFyUKhTpoPcTFFbn
NR+3j/fzXns1G1ZafjW2TtmoWzVN+TAYkEuII1SA7XPBX3g5mSjyKofIjnwovPcS
w21NsDik/FnjvVFVSODm5skUh77VjF8zrCtnEE6HBjbVtIw2bxTcCOZXgEidl39N
xvmUmf7FzuvtTlAR+SEhARhKsze9w+/wLNIe2fvrLWWYzUu28OTs7SdSFfaj6c+Z
ymZz2yAChF7qG1gkIv5vBJkDGKyzOXFN60mhUChXETWfNpTDD2flrf9r9HTfbekM
Czbw/dwjkEsiqKJ0hf0QceEXtROy/iMIYFzJ82HTgunFbZLpl0rPQ2hjOXP0ORzh
8CigkD75pZgCk2LwVY5v4QrTNwT2CdGlxOaGF7H1ZHZmlJCuztNIFofKIUeF+99V
tbcAUPx6MNmOe+tyY8XDas0vOMcHn2KDDxlSjQDlvr46v4RfrgBQxUUTgzQGNts+
1YqcZR/NDHI5tqoFOQ7ySWthhVdi1bDfPaROZ4sSiUiXGGUuWYiR7rB6tE+L7JGS
/caFZaDa00ZNxaGC2N430vQTKMpijltG40rY6vYGfJriyYbE0ZYxkteriWKe/Cum
EYcukCQp61KXAnXw+UqO/NdbAHYIuVpGseSxEFLDcPqZwZI5RCkZLpC5S3WBENxm
EI+EimKV3wIylKgjlqd5dVhvDk3ph6CPnubWfBVj0Oe/DFIP3tIpXlLis1GyomOU
6gUJhAS9Ma3T5AM2Adf9gUjaTNk7vgxdpG8dQ/+wzYOXLEm/suyWq7ApEHuVnBux
2j0qbpmbDnSlDHfEMISVyX6EPz5rLVsXe6fG+bTYwe9ergRetw6JrSkneTskU4MM
Ih3oOtBwIsgPlFETVaRYWl8K8ocjVyDUiDonAUHPFJvfXRIpUDrD8aTknra/O7fQ
FiBSicKo6PvlW7cJXrVJIEAP9WRcJlQChMerItwcH+AgP6fu3Vlu6xqfGH0rUHkd
R/tRxcjMAFSk3r7W8WlZ5Dhz6qXjYa3cOgeeTI0QmXC9BSQTrXZxNJHlgYujGJ7M
i8hRaLIcWq4V1EduNPorz1Ewl3MRyiayTcSPePz8LyjlFju1Uz333+I40o3MPMbx
htdTchwYe9qqWHS0PcRm9RVU/qpQ1sg+WE8Fz69KcZL09m3dHuKHQHhlyTmuibFR
zjZiS6ovScst71h3BVPpdmWsQxnYIMU4yq4sXYSXUvLn6mDPrjL/VLVC2fxyd5oT
UOZJ/54WeaRsVHrR0okXHTkwjOGJQAFykZH0HJKGn33RN/HS+EWLQWnCSASj1EsJ
Aq6Yue/uvH18/y4g7JSvidbTlpiBfblhWeV4WGP6RmFSN9X4NUqBWVo0+uJkID/X
pHr8mixFXFh4d+8g5XuYb2u00LKRTbHG+eoRPSEk3mXUBfDKyf6z/TFu4DFRvKvU
enlOvYJRefECh//UoQ+WlUP2nxD6s/SF1FjqfSN4iM2H+eUHo1Q68OUU4bdB4iy/
VPEq59pyGeub9O40Cx/4HDqrVtvkeILYVooCaQ7wHprk+zYya1rv0EvwL1Fsi6xM
GJgE8w9hyIS+KNVsCgb76zaPlUGK64w/fTn+heC+kaO/AKoNJ3ev1VZE59nDW7bN
nS5brZZyudCXRiBTJTC9Mg6xJGktCQ+SuIu+kD0KQpSdooTI82QhA6iTNgCpY7V9
I5C1X4YXtlbO1gvwyd6lljE6CcpX+Yy02uzStzymaIPmBqkCQAv88uPMh2ffcdyO
g9UMUfKZj99UHdR/FwiSLtcoFVyuYb/uf/v7/QG3gBCuMB/dELgWaEesiVPNYubd
o48v9PK3GvjZ1/Z+oGy0Qkl6LawoziH32urEO/qDl5F+oR3BxrYur2iKtJc/0Woh
iQyoQIUpfcaCbtvHNBi4qu+vNtB6yldcaHfS9zNWUHoTTaLmDQOc0pYBCG1ujIs2
Xqrdb/YatrmboixsKZKw+7PeYDn9TpPFXCfqnpDCY/8cuddde9Sp1n3U2a8a9aer
emgrlwVsRtw4MgBnupNMX75rW0MSCX3mkT0FszcmDbj2klNaTUuDXXNp2sZTLPib
JcHoH/oREUxkLpqF72IG5evGBFORmQxBdaJISHGSZYVhGrB2/Cu7qMr+ltOm6+UT
96ZL3FmMFP2QAU34/eL69u2/6KJyEpfNqZDQuhlqbK5mhPEB3nmSsEPDmRHXw3In
Hb/QOa5mKnvFC0uQNgJZT+SyEnOcbQGMY6qck5dZZ/tK4DJ5kbVhcjJ9K8Z5qdXz
NKFJ9EQINCJAwPJB7pcb71CLIB+57wvzOGvw3Okh/EuwOd34YuNxCXUgSlWFnBbC
ZWuoyivIn5wVE+WnVXuCKdJpZNUD5UPXdkvIhd3xY2bF1lg+0OzRtfqBG/QMpmBO
SP4n31SuJOFw8lrRD3LPwBohAE4sDGx0gh7W2qCg1rWnIfcBhBNDFW550kiXHhfX
J5b4Q5W1uci8LBGbpPAkl5qAJnFNiOg7I+0WK7Cb8p08vdKHoyTAwi9RhY8+NJPv
WSSemmbbvCULRnsPG+Cg9E5SDy+x2cqf4F6EvjeIk6DVdssfcV1P0WAZjiUa67Vc
L/QEXVbiKGjK0yaigBdXvwL7hghmPK6sXpYJTB3h6RxIZRjR7FCztcXiFZ8cPWzS
0wXTVhc7V+xYuXIUVPr7DdNbQiaM8T4EdH/SWFCUThxbBnvg5lwFLqM+zVJHtqay
+9AXhaUKtk9tl7/zkSCnykd/QIyA3MwOFkyju/S5wQmPfvQtbCyB2YLD+XWO4qCi
oGlJ1DowS8SyTbwIPUvlarVSdxE7nIq366NCu0ScmiGYa818ypaq9jn8v2WMvvvf
C3yn4qAOa+pYnEowAi39HP0QmFQVdEvfd2V2iWfUNbg4xV/Xtuxj9Ze4st1HZ3I8
oFGHeZR6zo7wsM8gNfo81I5QGNlbseJK8enw9COg6L6GrCSRHng1r5vVLSV7EWsU
oHKg23hPG+4bkMleGsnx++XOuMqYw0dzv27JV2lzrgU+fFNk8H747jGpH+jjVniM
2o/0TjwkevkCFWh/vXj9E0iRFjrENa9AS7PFfiITVgZGCK/RNfOeWV9k5p28YNIm
oVgTpoZ3pYOE+PAEyhZa4uLEe/8hh5BBvFGyG3mf8iqgGzH5oYrLoV3hreJRjTts
WXeZSQ9QAj4p7oCizF4M7HTxwBDHWvG3ttspZ0W0/t1ro5yemZuVwxIUbIKMgxZM
fS2m/IxV/ilY3M/6/DJnjatGI7QlfMR6PCa1FWfrJ3U0bgREK8E3h2nSp0ySzGhA
xzCyw3cwFccRrHQuR5GP3LTlT+ahkg2WwhZndhih6f7iSf0l8vo5r0sSCE03lt5u
/TfxlXebrKex7H5Qq2jcw+WjIZnzd9br7B2Da6U5qmrgc72pSQOpbevM4N9/762r
d3+lR2neSeIZCKK1xpoM/fryncdzEzbI1SvQY62Zzk+phNqT27rsTVeU4oo81Cft
nRyyCSTth821oEpvqtg8rpUY7Ky4MHSTMu+gHHG9DAonWZqCwuUZ8ZEfzMTRLNcR
hBTPneRREfq3XtzqF1GOe6glTF4Ls6P607+FP6797082daWxiCsGLrL++9BUV4/U
1D5SIQ/jKqKkND+FC0OLAAMAj2yd7hXnkKrH4XKfyeVzd6G5+vQkalEEjSW58a8s
SMoi+yctUwoflZl+kd7LQ/Uvoh35/6jfiXYQcCCd3PRI0i3GbtPSs+dZmieswzRL
Kl+091IactPCmddRZkhu/nuLvWdpjVJj9EZToezPemzNIaANHVhMX4qvYzbbWXI+
UMX9Pwlg1iOT/ZJfo+EZ3Mk4vfTi4RWzoXXN6jNM4I7EeAR3g4kkkED9nnX3k3DF
stfky/olh9M2oYH6UosviJJ0kzTAMh2KXrBB4vNgWBx27IW7JEbOHjNZ3Bt8w1Xq
szri1XssMq0zEu/ylEmtIOyKpeYgnUVtSUZwC2lOcoUJgEeUNdG4Pz/sVUNV/a21
3gtCzReIyAF7i/BQWFkq1XeIGoTySEeshIfjkodT+jztlia5sa5Bol/hvrinI8Iz
5I65wqgSaaYWVBrIDEiGFEIG+QC00YMOlpvYPYlt4rmftOF6LORlLU+B5gM97NxP
7fVG231Wrpr2Lu26UkdKPAnZLlrIyRcLGiu92sSRI4FdTCE3M4wKrcNxkHLQDCJb
h9z6Rla4dn1QpSt9QG2VPMOmUAwyDTzzBbz2N3Y51ciEfNUpwWVX/l846Z4x8CZs
WRfcowLVwbD0V+xfrKGKg645IJQjrMr3Jz44p+MiCTUUdRJe4p7A5UbcpHvABIFH
oupODfxhS9VAISxzq1X7PFEASEECgahguWMl/KHs5upsHXFAU3ut5Icm5OtL1sxE
2DJxHqKBlebZI9THtTp8DxTkL1qogqn36E0GGM5ojxI9jQn2mzPdRYapOXEATElJ
MQKu/JBdlj2CQA7ipmyJxvXWvyLZL7Y7QpreaqrWRt5zwROqbzllu+CLDI2Ktucu
J0RcdBdJA+Nl9soXPTdK1qUZF3MADqrSynnqiyq7XHhzb37TxQuJ6tVq4ak2gZqv
1Sn0M30yFBFLkCr6IXcTW6zGhUy71E43+cncbjVf9ttRanynGcEr3eiyUvxfRFoN
aBiOJMIjkJgmyY0xPe/wNzWg3CT6MMEoAEFd29tQpYlJt5qH68Kt+XhHyGURgXUi
pxUZO++IaOz11UT1OA4h/bYu6LpjLteTzc83gg7Zp13bZakNJbkrU0ALcFGlI52p
0k2wBuHFEd0kLNL82GoBC3CoPuWGpgWo4QHxyhtJYvNEjHb1+9fRRhKsgUFf1z6K
h2PnmrybQC6jB+IQkwUoYNtnpYpcjVJOxO6r3V9H6dAVB1nl670x5xOun1Q5agLT
iOC8m+/jAYZnxF+QxwzwAXHjYHc5Qism5CQBnq1Ygryiu+MZm43F0d3OfrrOo+tn
4ygTN7YwMXWAahTvLvRf1w984Zt8pdG+7vrDMgPrqt6fqAX6ZN04YLI8VlmpwOpK
hKNgZXwVkcwqfUWvnFedVZzgrfYQOXkaoT86G3bgSlr8i65s4gBaiMJtsBwOz055
zVZpY5WhyUgIWRILrIxsra+HFOHeTcIJcsTYqHs/hZQ178bOgwV4DNiHlRy9e2wR
T6VY16ekyL4v4W5mS87kZIS194N/Xj9bzqdjtUbDChTbimBk5t+qjPuIKZShSvKH
Y9ZZS5VEsBK+MxSilXK5F6KLyxZtyxj8pIo6TWAT0FVoeXoXZWApylgMfYomN/d8
qSFxyl9QCqqrygSKUMwHBSe6Ils5sxHZXB92t2K3VrTTXBgMuLLTN9DEg+7IWbnD
2KyW1xvmw/L9USf76XIItDS0JmbmjDujCbzvOJZcaSqvD1t8FSXH1KgA8CXDS31y
ZR1mYqEJO7loblekCqP8gMB4cmNcz5zhXJyDLzrauNYDw0yAbwsPOmUCY7GjW4Zc
eRdWCLtAvIo87kzFHaViPT7CDfeff8Jxxj0yMNYyG40P17kJdw9ip2EE9im7ZMSg
nLZs+ULYmkSM2jQM4tGD/8ew1LFaF5OYG5o+w60r7Ndiv4PzWA6aJkR48qI2GkU7
2ChAhCFHyUVkQYU4yODog96Z+C9nrkCnuRF7p1ZpbxFXkU5TIlFkkp1yl36Joy4e
EtwMPG1ALIR+ovffTpFzCBlToXb08C/B7G5R3iyHjZn3vGjQsyh7WKLcMrqdWMLl
/Fbp+J9HIp/oCYIpCURaPKDsiNIfrPAfBHpX8D7JlHF/wsWeQOlCLOhZ7pEDPuwy
QnoYAspbgvy747ZTl+zywE2pFaQvt0o264etfGqF9zYhO7IbLPeaZM4IvMe71ZyK
dtpj8zCxh6soFalOt2GC4hDiHysnAeHMdQGqIkeEqZe+viLzN+EB0m/m4vgffEFR
E4bnYxD/OBOxOeKO5htYTVuIAEpChQcdyEX0IZnWJdTsZbV7Ouga3C4A6ZJ/cgAw
b/W89xjunLwI8JQLQ1shzTLiYWmC8jM2W6n988owMP47uBCk0/QlunUnAzg2Pkpx
v40Rlx3FA7mL+M+6gel4hXccHjU2/YMekWy8reQUVuMjO394edAVMlulGZZujm0y
5+srg5iFyEGNVyWtxNijZP/UkYM9LrMsTu7UNzk3xm3c35VZ+/MkKB1D1h2waenY
yukJ5XB6MFetCIuYuiCtdwMIpOXD5efOgXkYSWvQHE3f/kvGaKdPFY6b7RCmklBn
Nzy3umhdmAGk6VlCD8Yr0sp4iDKRQtVgfeN5Tye0ZpZ4SC6CEhJ+1ADdg/Xq/7TW
5bp1ex4JbE4Ql7ZHO+NgDf/7pcZ+Qmd4UoOJcQkk8wnNJWX8m0d9TDaavNwmK3hL
0YCbTKfSA960GY/cfsW5pPUjkoWeMkZXU8i+H3GrdhqsLv7Zd++Fohs2EjbDnpg4
64f5nhn4CuU+sI5JgO6AQNyeBEMMOvrmuRbIfi5q01rrELaIPh0Hi0fAX+opHJOR
qO6fZmLsauhGntA3kN/VspNr2/UIMBVNjQr1EsaZ21eF3ChAeFlW5ATmjcJD+9xt
DICCuUWiJeP9kg/IX9x/3gt/ckoMS4V/Lbu9y44pMXBSSvwBt6EAStRRFAUxvq1P
N4KskaDzv6KWO8UGG8A23BMAv2RPrH6LOZ1qYYfsn+vDxZGuaPJW29jRi2+srltV
GRyk84OhxjqyY1y4H97NLsPRcOuYc7Q60LOZGdSIV9mYKvJ/ZjiH1G/MkbqNptsJ
XM3qnJEMaTWPfXOAZqp0QaIn04iAi5axVDBmTk3ozsvCbsO4pL7Gh3gRixvohElY
yk8GuKqxKZk8A5PZVfrbYCPEwwLcxgU7jpPkPeramu2RZgkWr1/UZhfiHCcAiuaq
8kVyalFHqWDn46H91BE/C1o9MhoQj6QcwSFZHufGwnVWfc4bnk2mA2tm7ewpYFee
vc9sLPHCE774tQ1JOmOSgs7nOUgWyODJPHEAgPT0PrWxupvSpsuy3rIRloTJK3Wb
WmjgV2gRKo/N44ztRmTur+tGu9tkAKzS4CNaCC8n5MVWtiEJ2Quz4T3yLdy2J1i2
2BIzpMU91DCNYrM3InmtcodI0zGs/c4/Ur2Sd7NcBIdhodTEp28iboccdiMuacvu
9rWxQUxbhbc0XhUDpPh9ZXsKD+rSKFzOFCOUrJTKpfdkvL/RYSUOUcltfc9GQjyU
PbPj3LByS5CkFf31b4Vq/zi6ZBWpiMjSGgJDku2Ek4MxUhW5CGBHVW4DT+n6ljCM
BlMzQT2H6NQG2UtNYB7nudEFiXg1IkirEUMi8ydZnAGAzDxjyG+1S00vrC5gHQKc
6rFKZxqfcuktusLLih/gT22Cjxa9r4ziCeKOJTHnUzyfklQQ8xcRADclejh0+k4W
8FavX+zjXIJXoEGNIBl4z3g9IBh4GiL3FtD+YSQJOHooottTpm9oWQpaRaLB/pvD
wSx+B4HzdOS13oNL4ojYqCSlHLMOvr2DHVo1Uloso5/IxIaofu6wiWTbc3b1l01O
9Em6vDo8oXpEpMUCbEr2OrDTigWhcW3lUtCRzEpiZA+t//oclWxPE5V4e/1/pm2T
VQbf5n2def9GmQF0kl6ML96zv3EYimmzd7tBjPVZ7vt4i8AfOI99l9tAyPnd947x
vXFB6XzRPu115ARtzeGYlvWWz8Tckb9KZ+SV7kml3r9vjtX5d5/HqXL7GRv/QfQm
jJiXhWQj+/oJRquig8LWfL3WAZDtOs/E3bSI07B9lHM9SfSuHJ2EdsSChoV2N4Oi
61fjAwICyruTH97bGiznzwRTqDeW489KpuqMPgaRdaRi9W1S0mgVJqLdjytDDPR1
JTt9UweBFLuoFfURGv/T105KkO992gluGp2wF4OcQ+5hzQoixgCemANm505/rWwl
jLwRbhYSMenWzH5PW7ilhQGQ8XMIxG60YSDaa06eHe5Y9BcIOLUuJyw70c2KDy/m
Ay9pvMReKGyEcocDd4Bq4DxK+Qu7K22udzglOQTmSA6ipKSqZSM9SDTYK4576X/4
afhW+D7RfJEnJzcxlyRx3+mawELayunebIqvli+2VGNNW4yzuPfzhm0zvJpUzKu3
dwDbFZTSkkh71nC09wmHSHCA+ayvYhhblPzk3lFghVa59z0ipGIqwcpEtzrcaQ5e
sT2Gt2kWQfdp1QuQ2sE+Xv2YJgjjB9OIwwZYwk4do/nwsj7cHOsduvlwRTg5DFN6
XxC6cv64sPefUMmrXbT69a6Qw7c5vB/cH6yGY/wHtN6/Xc+RR46vHpZZ360GbWZ2
9IU+YItOd2oZxRH2hvQvL9mGsz/xMB3ZHnnJ1EL6VrWeRKk9ZIFTDHoCfLUThIt3
625QOLusxfY9DUa2ZQ/X7cnmZGq+EwUJznhWXL609u707M50ZO4Lp99u84dldv4G
UgqxYWN2l0j2vs+ZbMWUArMFehH2oYxDjlJZTeBlEvt3yy3P3CEh8iKVW7o3SU3B
hR9G92cQxj6Ujq/aG8sHsNhNygsQWSHVJcCeo5cCNYbvyMdtxDQNTymJHO/dneC1
O5y+iqkOg+x68uVNRP6w5BksB/1QjcxT8lQU2wRH4kFNv8bg2Ta1Me1gyi/iFcQt
GYyvQ7hx08iJCZ+tZkD/PAYBLmQgbO4FGSSuvUdUtmZYtk8aCqk1lVkC6Il5NHp2
ZHaqn70/m7hKZWsA6D/6USDAaNxNIhMmhbHPDruHBiuiUXxxy29aRECwxi6IeENN
XysYysKXoJK8bxMGKi8Yq0KLC7dauAZTrpW5JJnCeHvTvlQtCmxdRu8vtjcbTObI
kuDcNrnL0tha+JupqSNnY+8KMxa1miIGOTp6ifYwXq5OMET6y1HyXa/jU/69K8s/
A0i1GJJN9qOyzN3sAvfrvxdyMxM0UAe7B5b28DjvdT03mVwJpdnYEFSMBu+lfRm8
5elARVtrqg2FDGd4ckJwE+9f4/tbUFQ9iPRLOI6Pk9ba+DCRruFgMcRclpEJqG5A
3jmR9megHG2bVzmt/e6PJPG3vTPHICZG6/NhFN9HL/lPmTZDsCga1v1vp0trsxEu
zMEU+AZu6/thaPXlehwIUK5hdBexE1dy8GOVzfDJJYOEBtgUqxhgkHgwx33lQ03G
fRH6bs3uOf1XE55yGAtAmHsoWkP7OEETh2NK1upKMVIEp3GchuyJ13JawHmmMB5I
vbfoJYI8fJEy7jr0RxI/fbrCdVxz7Q/8Sfb7Gl1eFsH1BQE0ZuZwp8GDv59UYsd2
1Hhuq0sIjgAaSxNCUrZF9dD3xRkIGBRvPSQyALn8ZKTrr8/qI6GO63X21qIvRHyE
u6OxI2XxTP/V55VgujJnxaFvdhCE98Bp2P7Y1tL5czjp9qMhyN34uA0yvH0gLfsu
uqbXpp/OXmuDVjKe+3A9rrpo87c1bAD1LEfzzvHcAjZ8LkeLWV1H4qeDnnL99rWp
sFzbDb592eodyTc4YrF5T6TL/5UVMG50/Au6wGxmV61SvoO0DFvrppB0zVqlcqd1
5+h1J1ZdSOJZUKEXkqHPuuwJKLE6RRc1HbYxBvY5eraBoPBjHQIZvspz8G9Cg6Pm
/izjINdhrAXTPpKfJQRjDurgDUFoE2dfdX/d+Tdcb5U5CJG74k2OHjhcZiQDqMuE
tmzCI9Ej7y+qZ6YB1rNOeJbrZUoOSy9RuEbQj4tyj3zWugJ66PTLIFqsACsQ54M1
Icx/Hfy94fYTCFoBT3+r1C7ZbM+HwsbbsFdTj5ZGOl26X1WiFtnO0qy4I9gAPw6b
vMv+IRIjpVt/JSmT2gX9w9kWBBKf82Ic6y6Z/gOBAyCoBNlKKCBs+igomhIPxp/3
JdiMWnM0EPrZdJWOOWCDcWFqSPfscvLEk8qI++VTKb1GwRkSSf9I13IPz0tNwO+X
yM1/vw5LtvWVxgPGdgjtNrW2ZKzij/XlBzfwAV6cJPlISShLlTfMaUldt5IM6AQB
QY3PnpDBAwZ45qqisu9SJKzkIoIhq8qHsZe85B/wJlrsJwnhwpMXN1s9u0RF3YZJ
yQ2rm5/NqwTib4bBF+9KyjpZwU5hfp1xhWQJYJ4adsL8SlYBZ1rkCsKmOy7L92ry
hN0PfeGL9xJ/YBU4srh1xXDzMQhPU9gm3GeJ8ODG1okRm6d5Fptr5GCOI0PprNsY
J0OfqZ+jo00jL9+0b0j3YwG2POlUD7jjEp7hlGdpH16HMtJJSD8l3OQj+pHdMUYv
at1rnEbdAbM3SCD9/Z6eWN0jOYhVNay2raF0fA/SLEGPg6irhKtxTzsTnnPHf8nj
S0NqGqKq2X/NQ91WC3LBsoqIW5FdQqMTxvdXc4ZeXHQAH3okZ7N0fHU/NF511uXO
dxlL9Me2j/qLYL4l3XwItLkN93gIRjy4K+flXuEWoo9O3qJBycymHi1JAR1Aaa2N
7PBYk4hHr3PSkxpoNEWRGauJ/L7+cnXY7oAKaLkTRdamuKPtm36O4cr/0yoqZwdX
YZl5QNSeJ0ILkhuw7p0VjbR8+PnkJiaWe2OpHoNxW6P0/3Q9UNRkd8zUJSVi9LDe
mVSkdUCGk3D5Q5iyCGQAQW3XMlL5lMn7iaIwFxb9CincEO+1ju9AywqI6a4RZ5Md
26yUePacmlZf7a59ekZYMDOfGvVqPL4nrOC57udMIdlrBTu5U5/CS6szz82vmLed
QH7dWZ/0Bd+/CYITIrt8tqLroexIqQCrB8QXVP72H0sRbs1DkUQUQOox1OqRrd+o
yovE8hm8I7AHi4OnLFLwwbt9AokmKo3xGYkchBbArQlhLXNRiVsZoVqK+vlVWls4
4uxn5bM69cwjSMs+w/X2GJ8IiLCNjOaQ9kBY24kW8sMiwRE60X4AETimWSLfsrBR
WRCEJShaoSGBrOdzJPxdoa4rKpcy/TtgeOArXNSaAKlsawzmsPa0mmEr7Ho3a2Va
STlWWmsXRJ/ahZblCFkRNV68FzRL4ipyjtl/ZaBvzYKoMM3rq9vSBbtK9j+Qq803
xyNMvRkRRp9VvUCWt6aRHjc6BjtYbCrI0b8jL/2ZHjjX7HVHX37F3mtQvjYmsmTF
ynnBsPa+lssu5CXHQ2WRWCMzwXwuWI/8mIE+wKSOxuemxZSLrgkbJ66pgXe6bjqS
wzPYjrIokRn4WMdh+o97DOj5RZ47eY9SKOODBm8IknQBuaNKXZkxtSVcqp8bJQ3E
EqGbCWZdsUfx3FCVHLm/tt71dL2l3rpkVbuR+m4TY6pSOqjI+Pu8WHvJ7+kTB41n
zMe7bdhj48qjM/STM9gZGEIgby6OTj0QV284bWyBHuIOtE9TzYYkkvL0UjI+McaD
t9gHlouwWsrWt91luuCgr4FSDUOfiZmtm+DQaOR/7Pxy0ldcFXG8dnCt6T9ACKTp
Owj5ngovyRbzMctoFZUM+5Crvl0XreXR0xTs4I7DaoVHhstsEAYRR7kr6IaOnlrN
n0uqvoLKFU55d6MvTl4Zi+dC3ela94U99PYbvBBzpK4FWrdIvwrq9+BC0l/M35RL
pnp8Pm7KbXAFv8FX6i9dkUL0Ca1eG0OIB6jd4KPgAEQeDB3jraF8dIZVZd7IcL6K
KV+Lww7W9vSdM2XZObxnxyWoz6AN4QtVr8LvnHReoTisqDsCwQnMvibCYiCxuSx2
xtJPeX5dZXkNetyOIgJSCaWVN8aBU9C+BtYYbacwRQMJz5uxYDqrdWU/HLoinlRV
GHUeRxwFUdme1Rois08+uEZZ0y0jxoXN5RqxCYH+ab06ViKHukLLl1M9WdkX9xHP
dmkR/G3JW/5tEcYwnvZwlDuS5yh9WbpKH1JzsdymNVFqaph+gLaWYm+cFVTzJSpm
O0ien2g/IsqFiXPdV+LNenBazcyuA7mUY5iOuL6Ajthjx5FznANBrgYSh1j5SIBf
LFxPXPjWS5Q+sjvLqzBFvRfGiZa82p8EKBNN8HKhaOr/XET5eKf0HPUHn7nj+5Iv
oLiT5CcuYZDzToXe6s803GwtjYOI7liGwkx5VckQPkR1xwxNq2q+fIMOQXbWsbSS
KWfyNbSx3Uv1rnG8GgtPAxjnesZ8nIOtenWY52/f7mS2H9fIRViLdygMQBp3c3OP
TQexQEF+H+djxplhhMbVWJOLjNnchR8y9ALDidQv4kCMAnkzB8RdREZb8Y0wq1NX
4Pu9/1befTvkQPMLNve9kDwU4SVY9IcGvuw8cIttp2oUFCBO8u8dlWeYsmQNuyPa
s0COVLLZfHotpzrPCgIMmk8yPq+kLH9j/MUFaYp4OrWlTAwSfYnRG7qm/PPDSiuG
AsNlEYH8I6fHKLUMkmGkljI2VTy7nHCFS+f4YcOvV+1DQIeDHxuvKmGUF3fiAYJj
bu6PTNOD5VO7e8pS3XgFunaaXLBEVi1WQTJxG+1i76/0UwX24OzA+QTTE8nQmxdS
e/IN0R4QeDvbUhDHDwlp6sr3N5DIPsa4YVIgYJpgovXUAPuSXSwsbO1u3RcjZJrM
/oVroihy6WaWCueCDyEFU1Sgk0lbUTG33Rk1Ur6gmg//eZuh191LvEaqGlfExcCr
0WK4k0G2Zju8F4CiNlF+SIIn8KlBhYjG8ED+PhyB9kk6dWHVMGX66p3mqYc4w2xl
IBTBqoQu9d6QIhg3fBpho6EUsAzWRTImznbtcbUb6Cgp8Tc1MUnY9ZNHK1BQV/Bw
vgK3oWWAgnvoHagIXZszNdLnZp8fquJLm3zgfikCaIqeJuzBTPKvi5DTcf9Y4blY
U7xhb+jh744GYQe/UtYBilkMhSpgtH7q+pRSsi8qNwCpsOUz6zea2x4gfek/8r0j
g/3RHelo48ZrMQJ09vjn+hyBcXXZcoSIMKIahOlSz2744KqgRQwuOwXnLKvqRARh
Kv3Hdhj7w7YJfoQZdBdfseJ1w1fU5QwrH/H+C3QfYzmvH+4gi8CGuM6lQFupvn2/
g9aKSmEvHLPBNmpPUnv97IZHnPXtGEhF8Z6TACZXJ/toUIbEL3gIBDF0UoLrFSDc
kFpvVL02kO4cPnLZY2zi9lpSm9PIB38zxHVUeGaQF3GFTgxxqZqdU+BfQD5l+Edo
yD8LvoJD/sYwVKqWiQY/G9D4P7lwdvDocsYbUNmxEamQuWqBGv+eeLcu0AuFoCM5
qP8FIQYMOfaZq/+DP9LFr5Tb8W5t1e53VJMwuG5plWnvTKyCe+eWs0A0bjEXORJ9
hHh9SDnswtMT3UEA3P6oX/Lw5UMKzDPhN6z0AUtAlGBMNxm4BdPeu6runIR0k1pA
hmeZA1RT2sR0jenXdC9MazxBjLtK6GpQsAMbvW5VXHSw2GbwLyk1+kKrKhKWC3BH
86B+ry3Zok8MQLTQe7/6mnGOcFy/DyphwHOOkyGDHUca79RoNhgBvO8NqFk7EE0e
fR2c6ZzouK3hphWgLncsjn2DhtJBAxIVodUrtpA7g05ZTBfDlxD45pWgZYLDn49m
jfAD8e30n8vQ/4NDJUOhpHX0Y8OHUOa1rL/M/g5TOckIBMHRgZMNxgpYRos4ORwE
LZ/TqJw9vDugLW61K2ZqzKARox1R/qVPkV+f3gCJFTbHXry1Fvy0ZbGou1sw4C/M
MNzddemo/KVPcnQFQMwGNBn3fMynvd2nLpfmfmHx8KgiUQrvNxkUBp855TD+Uapm
JQID8Ci9ts6YvxPmGB7KgkXRsXI+VTpCbzNrs/QKLbryW1wsp5lWZ6aGWfIsz4N9
0vvgkbyyk9+NW50JoH9PzBzkwY+CiICXM0HkYc2LpNm4+vFBSXXPZJURcVlfrzvr
dcTVg6eIAmt1VtkfZkXg2AwCcyOHouQXXMIugiygnqa6FNo7VwTlg6NxvYE1hcV+
PdmkTpnqATB2iws1D/fbZ6GQbngV8JyaRAAs8jq90M+wVQv2L+y0WnNDEltqnXAh
auCKflD/S1UvhWMGpT6Px1iQwHmf9NVSFSAsGKUSUW0MRKaDT1JQkE5cb4ZCgz3W
vm7VjFPbmP0XwVFVBKUs9YTPB1bjlWPZqg0mN2brPVmPHyvvs8kUxCR7sb8leyD6
v1yW8jN480uzGAQFuboj4syhBHUNcm2n+s5Lt1jJHZWsR/Kfd2FjIXOB2yEnwFEF
XsSS42IBA0hWA5JsLlmhIzYGqb+4m4ZBJi+SaPJZi+r0F8OCXgzfabaqTY5YIy+1
5ag47+8nSXY9fd+HCplrMsxYRxa+4dlej5/Mjz48TsWFCj4fk3qJpBeTFPjK4a2Y
xnO8JeFEKey49h54sCZMRQljPiW5IlGvbI0eMH4Ei4kkvA412ySrn9O29q/wrQHv
nT2HbX9/mxV8uSweShH5DUO7gjP6FISvFqiT8N4Zv6b5SfYjYwFjdxGoChN9bKpf
Lj+STkwN/TdRmzxwroM1W+lzL4sGAMjNrR1pPOGErurfAWDWSNWo6SpxhzOXd+jo
ZoDI26t2qUwGyR5xNyhHvHjxzcHryVEtkimuPFpauSrEqHsWr5K7jjRx/ysUf8Bw
w+EigdkmbGOEmcEiRd74LQMuCsXmLTyYecPIbrkNvowmT7sKcb6zQpRuzvyjevrh
SeCoSlG93KpEOgs1TbQwUmzoyKPEsX8pI2qGV56nLANmZNpUtJJnPO82gv3xYbUQ
OqUinkhbJY7XhI4OurrhE+QdrPZHFClVwqas4JkaXaLlEaY19EBeaLJTzbH4e/Xj
jKLShZ+haNhFdhOHTaLEBMfvMm75sUQ4pmhkByindTJW477pX4KpK7eUN5Gov7vv
PK8MkJ5D+viipqcpGQ+jyx+F/k9tryl9S+sbcxZTXLEeUCg886ZId/MaDQ6x/7Nv
aXZzWsQ7Fzw2yCxtIDZrY/JK80t0KrKN+oPygIBCGU9KLy9DsWaohyZmutjAF9zn
AY7ejcONPQoqqi/Fc158OYudkIi4naHy/A6Me5cf5oel3hq/9eXHNKpMG2GQH3+z
9k0WAXBfyvUskxk7DMbflApcaASRwEPyzK9gxzZUx1PO9jA2ItzJRmable70QIfS
gdrcYFY22/foaRqKWsycj8kG1WIB3Y3skwIBGjyjCbMxJ6bL2Ds/m+iBzvxf+97k
0yWGzjNuGh7YQicfQzLg8O00KTMUGoa+W01dFnEn9oYnCDUAaOVRgUyN/v5lmhgS
ZsfKwWvyopRCjlKXCNDWUwzZJ48way7+4EdNI9P6geZLsnGtEhAF+PCT6orAjokP
0CgUOvvyjpK4sg3Y/BNBIEUK5dlPviHy5YJ9OyZ1rPXBS1qQXPmz7sppMapF2FT/
2auDSZks5Qh07u6tURFxpIoKkneEiLDbzi+t435+HyGyRP/5/9Wdu8gWaMN519WC
jPn70VB80BZM3Yt2jNXJhOlgnlzLER44DW84zBDNZkFH8LlogoS6qX9QTDLhjF4L
6PCUbkWRLEcnc1EXRHGjZcBxjEhqRfImhTX7uEY67QzXqF7C5wzKi9zWEkTzObaf
yaop0quemIJx37IfcyGROvmSZJhiwcUOum8cgX4GiUcfNbJRlbeo5KHprYnInpsV
ngym7svBm97ma4H/ioS558pxAuY8wbd7NFHuvfDpGE9AqQ2UHvFKEg8UpEGB+x28
SNXT4sckONgxSsckPqXnyBbixojUYj0GddXc9RcvB7yO9u0/alkVsvCvcb99W0lI
0TB99neBajXhA0qeKYdjcfJ5lsLNr5pQ7QLYAQ4XNV6lJ5HV+2g9+ZzzArIRvfnC
rwnjGXM7qos8po4pSz0+qCupo0MTuy9YccOtRfjIQGjLRmcVq9H5Eda5fWzQFzN+
xe02vb0cxBcTIUMtqgwGjGQN9DszHWVJN7LO/ORqmuKKV3mA26JmDMwSGVYlHHIs
5GK7015/aVSJUa4j1aQuAhOehoaGlQeh4Lac74OsOF7SQa/LqdM/cp9Ak9eeVA3U
EI4dWU87g0wEgZDOCgwD4XZDY2p3/MHWykVnn46+9VWnu/TQATMLBApOI31qodlF
QnshuVwRsX6fV/EmL8HKY/9UAuE7nUSqZJrUQhuJzHCg6uJsbkPaN9qmPhbyQX+s
yKP7E7PE/GxlN8LBSKKbSrMT5l3OCncJ7+jq3PsIx+HfscbU64KH7SdGnxsmvEPd
BUzr07mI7AQvDxqrXKFncHLypcum42RVOm5Wq3UD9D7inWTPTecuVYyEDETI0Tqz
08114EuzYYyHA2cEIJeEHPCX48gzYYvHZmfIqyMMbr+GiKw4tTi4FL3lJi9ZrAyE
K8a8HlapQLLDwO37SF4GEYDyoEaVUMrF2V1kOATt34lZQctBJ29YXf2mETmloHvO
SYFTCPW+wuVZG/nPIhWpCVzvQduoeYTtZW8vzbkHZYsglQ0AWeREzJ0vTGxeCMVD
XnuKmysbfT6evnyj1tyLafzCyRaaMMOrfJ/KvOxzAADqW3+rhseTsOkKp7VEvaYY
ZGe1ANsnBC26C9O19oY7+lRI3SOUlriUnSGa5A2LKa50m1DD/qp0NP1qmCkBD1cN
QQbWtm9CP77YUWaIUrptpWtYAwZt4K1tojOgbUIBOBJAZaEQ3Befn4E9z62bJwAt
tfJDOBxnMWflLpr7aLgaG9vFgFtc/yNIzxHuAGbzF5OzE4w7hEhZjzIY+9kESaGx
Z3Dnlg1XHxMRP8tgQbOdO0PWXMOee5u8K4HYdb5UeLKPyycqRWQxZ00SIvkQi21z
4hI3umrE2DJn+3aIM+RnDHI77/LQaZ1sWtx4ZMxQYygmcNUOeGoRYHMcs6nSuAS0
3/I3T7j2rddc8oZuYn/dAxcCOlodvK+KJbtbTnIGI3B/okiMIDpvaIcTZeWGwzO9
72X5LrTRDGdBfJWqYDTo5dGIatBxNFQjYPiJphye15oBb+XKWR2J66rFL1Y9pOn2
FWNf7DrpO5rvlXVMJ0GPeq64R+x++od5+Jubcy+8eaxFL6iKmS/LBej0nels3kbG
2cIvRALGOqcyi9+OKpWOzNjZhzLyUHFAtQ//m0mjSvVbZhhZoptQStaXb6QTs0Ti
jFl5+rSlKCJMWnbnFKRgE7aVA2XxK1A3S12SzunnEo20iqWUnY7mn4HmYg9ocWtm
99RHHhthGbeN/qlV9Z09/gmWiYyCcR0+ctu25Pf0Jf3w0KYvwBO8Cc9XZMB720bf
fgfejr+z1Eh+yKsiGdL154FcCOPeXroDBwjJv0rOIWMWNjvviF/IJdHVUhCjFiB4
ufpHmi5pJgNKOlmMqBhbUGfQaa3ksjYL7Xj+v+4eoelaqsoQnh7WwOYvnlh57hnN
hyB3lsIQ2P6Q7YCK/WyhMAAEduwVBszoVRDfAnTLliR9eVhW0x1HOjmFBkvJosmc
c3zSO/3n1Bry94Hrs8UME4ZqvdDky5hrxivcnu6J9QscTvlWblqty8Spe3xTWDlt
/9OTxsqQP4QYpLMm8Yxd26ecNxnVEqypFcKs/HdF2tJE6QyJBs8Q+HZ81Zhp5Uuq
TaD8bs6eB83mxu+bca4fbXKFbOao2Z1OzCQg4vI3YsZL9j2zERL5WHfCWJ5/0CGf
G+HgimM0KXborQiOUhUuN9ia4BD+UXE/ZIBycXPbu66AVjlAMLqVMOu2meNxQvRl
93DVq42ZRoVOtlpdtye0C5UXHTdb+krZkI9LeLMDddLD+RbFF+pIhVnyrk0iIFrV
FpT24IuDVFvmoWTbuTE3shLm+WBuHchHmvp7sKqLCuoHf0Zl1bpJD1dlrvq82M+5
/QLJHYCZji0N81S1A7oYvDXm/3ZjxhZERRiwQ9F+/FGzMMI/V+CccUUdmtUzBH+J
1PzV0y6ISXDVOxcZujCO38XmxIlyNai7LJLLdUQwixiI3NYDi6gEcQK23vkXHI68
G17vWXXQm/6fGOHTNJfyXYuomJEoKtmfe2SNwmR0uw5H6MajAXUTdcTDIcxj9zKS
A/U9brW27ZIPus/NB18qMF9XbhaOrwm0s70QUD/7UFbRjDUkbWYsqNNEn5dTX8G8
VnrP6O8lRifz/TkjzPEO8iQDX1/Ah4AYNMatNyGM6RRz5wB9kub0sFln6wy0mEhX
nfTlx3gOp5eysfi/qWCLczTnNS17atGV1ykMIYlru2jE/wCty9Yh6hYPLl/9nwIe
bYpHeKp6mTulkJalXwq59mDE/lslRlCkEybzqqW4hMAQGCXqw1ZC9peD/E0PPsTT
vVeCuVSluco9qF4hIzp6dtj/rv0clbmTAenoyZsIwawdQ65kR2u/lwnc46YyVRxx
40h0gSArq5cDsyZOZZ90QTL6WiWlLkrOTPLvIoAgzycjqGusGQsEdDYhzP7unCUz
8BEWmIr40RDD8AzaVMkHkWLnYWymbmFA7GV2LMbPy2TwihUOhNIfCG2NAcYsJ6BQ
S5hZEl1PbbntU+MwV0Qn3RR0Gt6lyVxGypm/60Inb40nZkFiVR1ZU0Jdmpfu5pon
uXK5IFRorD4IrSBXfUVJSki4nx602cn2sMyjgNZbGEbZk3zoC0ZWMDX7zhzUWfQq
OxZkjYd10kxrExjewhoCw95kA5ENdwN9u6ddpYZennyvwDvuKRcUKRMg9IYYcWmH
ktrnJurCDPKe8kUDIW2pMtqXcn+Fg9GmTFGfyWYrmC36HfNxXINs7qOERgLVY7tQ
MOAH2yhXxbViMKLXQT08P76y6GmzhWcEd4Ge2idOPRkdPtVcJdCSdBIuP4UQgHc4
eI0oX8cr1E85mfEzDtgti8Otmc96NnBVYttYDZSJKtfAqxk5Wue3Pft4yWoNvLwM
up9VIuSI8Okn19cEeCt1MY+DXNPQNWYAgptq5+IzZhvo0rVzk2gGT/srsRm/Y2lr
/HNS5HvyXJrPGdPMz8+ZhSNY0qOj6aIxommQJW/KcQY38+bdvgqPprEAG3JxpCF0
jH22KiIpF6+rAK3cKDT8KieuVjjZjS7xLriP0EVhvQzc6KOrJjFWO9/6WpNR8VgY
Pfd/gdGbxsvHX07pWLHzcg5uwhyBIOoGJmdd/I84cW4IAEF2efEv57sW/FMpstEB
MXO7gNAMvRcfN1s7QTcYN2AzH4V0XTA6Qg6pHtKWsEelXcPFbmBNTuuIRYVz3ZFO
bU0wjj8DM3alYq11d3Vf7IXbbLr1HvbKDRZDTGKqPuJikUkLWtB5bYXMcB22QLDu
wleN7eXWo7wfGlg9GQc2x13owR3Q5etSpLKGAkuUYVVXNkOyU25FjxbA0R5ULy2u
fIu21adJUkJfyFVnh6WQiop2xk9irp8llmKrvcmsNzOWpCFZguRO7jtrWD+MOvYm
KesjHwVG+Q3K3utqZNsiKZJWY0xDDEYKucTE/uTUkKAwSve/emSfx06iN6vS243G
NVZ4CkQr6NSaaeE7qkqHSmIbCx0QhGE6ac1iQiTWCNcqsw4KIn+BCpEOBrBorHYE
EOzuyDbjdItbXCIpZLl2wKsp5YUCCTNd6bn7OsVC9kWNLa+0JUdlLUwBakRkIEVr
mhm1Og1/gT5VBtMrSEBoKZj2FL12iXGfhs5r/jyCF3xqE/DP83JHMwc0k3Kp89Zp
pab9GOAURRNxL6YLe/Me4V5lsJLijZFql94tndNh2KwjCGC/NGUeQlVRlgRasSKo
5mJ6Kfa1q8kZ3roxgDInifijqLhQFm8Ed7mycMecU8m5x7FZupJQvZo0IGOt2llx
J0OMPiENaJAGNqAo4geQRDN0lb3a21sdFKFWemb1+moUgbibNQOJOcdSmPNZ+D+c
bLaTIl52tYdUWpT4HBvO/lwf7o+7FU9NROnlt4+/OoM+tnIqWG2OVtxuHYoJb6n1
lKQxQilQLMKr55+zf77O/1EHzFNZR+zlsX5JTAqEybj+C6mLRR3YZC0YB95Bdj8f
xAFB01IKmfWYNrvd0Ju2h5GQcmUxiwp8eV4aHlb+6glMWqWifgHW9is9yl67Tq2U
KojLauaVKrIyTPUcVsIlxU91u1QpeMuNE9SRsb6lmEGRrmYDyVL1SrJAChq5T+6F
v0xbNqKvqYYvSJShmDjrX2HGL2AQwHpcnrfe/nXGGrBb7gI7gSsg6zAxr9BVO3Xu
yVmBNVOp+49kPyDznHo8g+henMOILV9pNTk9E5BGIv3vdMIKsPQuKy9J3Iooo99F
6WMlzBCrhbDE/qvTw0sDTLPWfhtPSQPQ04n2gCLeBK9JgMmFTVTtuoO91Sm3/LyI
IgGtk1NEiEApiuSvgeWWYyk7oJ7cp1iSvEDTWtpTi3jX9eQMu7efFFaYEfh2c0Ev
TeNaFOQa+ilVRN7OZWRjyYaC0Dbvet+w7ZPROVMIORMQL7q0uMIVmH4tlmvDidAh
G2LLL/Z5KQpE8uJvzQ7DPiljxHG1OMO1H//tvEgYcTBn0KYcJ/y8kxn7a1NjhipE
0PmlAPDJp1aSYAoFpP5Vnp9VkG3FcLLh2cbNExtfhXe9l/1SMIxjpJwWcS/XcV9P
H8o1v2bJOFclAFCcRGIHcl6qCGS5P1VPZWKxyfHrhtXqrJnJd54vffJfF7aAWczi
1lNw5pQ6+hgokx59/R3FCDES+NO9SSfzLTSG1gh1+JUgO2ALc2qV5N8EmG2YrMFW
ZOStxnxMZ9kFzK3B7RrMqu7ipigmBLuu+AJP8FKlPl0mZhXj0EbIHdSUHNrLcpS9
OAilMV1MmBlhVnLRjBCgaXrgkNyElUhaG4j7aoQ8WHFgOrGnnr7A979gHjF/wZxa
+wP1zREr/eSejJ5OhYOJJNIdSuGs9WEoxeHVef1AyZTgci2H3s38NhYUv6JmaK12
UGofaXDzhoNckO4FvBXJD0nj/+kpM/hUgLMQOGYDib2ha9C05V7ua7W822zjLlnK
cX1/iWRr8KqyCo1NnhH05Vz5WEozur2SLT9PKDyx/H8iKb3U0u8skFp5WTy/1x3P
fyImDsrXORm35X+d//t3yd9XFccUgOn+oWl6Hs/VWk0cmUiYJUsmirYdKX0TTQty
msJ7lg9GzPEtiXWzPR2AJJ/dsc1ZTpDJnBEmFQOC9ArwjAsmjO1HSi0PKm3EncGK
XudeQ3lpXF4bOktLINc+2yIRPuDNpySPSyk4n7FGc3EssTWYC9hnLX+0mUlGeuAa
zWRkQmmNj2jlWKc1QlnULylVhQ52q6oRDxhypEAxma50/zyxHZj7GRRdKA1Txw7/
70PWPXSm4MEsLdJJIBr53/384HxlEf8U9zyp3BzkFmSpn0V/gSbmz9ZoVU78QWxK
ZPKaNMSOPA8r/1l1zmH1Jz2HhMwavYgdvbYKXlorvBornZuRffWmQNPOfDUvekfI
s2um35LibGC0m9uYCkYkkTNf+9jGdZer2JsU1nDXBAXZP6yIdKHCT48keNuMGUUK
UGSCIEdI9+jL4pkE8VwJ5C2VTYIzTYOxeJXXzueUhYledMC1wSgUNcEvsJZE01N6
rKse6qcX+aI7HUVvNN/uHoYFhNYOH5LK18O98S5rKVQsjDJ64HRdCbiKG35CjANd
pX8xFEEg6wM+B1PnKj3wJXOls6xiiqlkWc8uxQVKOAouc0hT+dUVib4n2NRHdgP9
kK61+Fbab7AGvOYc4AapMHqkWgYCyeGD5MghgZXtHC/siNq9b0A4UiLOxYjq3bPc
KVL/uUCqErlOe/h3n6x3gvFqZN9GxSVMrPRNFSoMSHg35WTlENPPJXtGKi9x0DRp
PvkH70Bh8OgHQCQfk85FZCmuw6RDZadEJhLCfG6tpBiEY1jr59HL+IhO9GvfX77p
1QAF8hLLQMwbwmhXmslBilUMm7HuXISamFKRkHP2JvuZkxGULA3DhkVjqL5JrScZ
DUn7ulcnFyC9/wvKXJDEgV+id8kQYD2DFgPw90D7gJznEuYemXBgiXpuX03p5tnl
cAcBEUkz0bS76yEsXo/3z4IyBEYag3EHOowHr4p6Y/BZlBodhbGFEFYHZClPddTW
qb/zwPR1G4phivHWcSbqr4IPQxp3si9RwD6l9SA2+sk+qYfQHnqFFqmnJKeMfsME
oeevdAjSuViXGunV91xJqLS+JM/CSmqgPp80rVgwolZGCds7AuVc9YyoRn1Ex05O
i8z6Zcw1iC4Oxv308XXthBcgZZEI3s//cgZbRE2taq/Z6ZTEo7oVTTFqza8dXcCT
4W2PzvwZhbu8NVU5nugTCIUkKEPLWIMkW1W2moNC8vxxrNGEl4Wk6VaF1xDtHre3
KP0oYTceULd7C4DHDYjniJAItRhWOY5J2Oqe5/IMYv3pLXZs+gWEesEwEsw3pniW
mTnu0dR20th4uqFbeymCNGfzSSKb2qkIj+sbd8hvyd3vddUHXhilgLqy8/rRetFY
ytAoC0qvrtHRMadpOQdePc526L01L3UPCMp27br0yp/HpjxzSO/dUYgp9yD37syU
droNPzthCmeUyEpVHBDgnoERRX09aMKI+HJzynLKB2mopesj5sMe5OCZabVHW7qV
M1vHWU2YWqJ6E46Xgfs93zksJwn8KDuWpHhsQkirLU4Sh3I9a2R7Lwwsb06ChjD1
6GCSyuYKs89OyLDg5ESHm5/qunFoInL4aNYT80Pv259NhCs4oSAsGCYmXEg0gKgZ
Ke7eIQBlZCJtEiyjIOiCbvXq/JOyKg1pmfEXOntJtw/FRsC+7Sg1jYgkFenaZuGZ
q5FR6mN8cpN4ABg/Rf0n0GDXXwtUav/s1ozUiVMtkMtytnspvGsm1FhV4w3mGz2s
3OEe00yhX4iIHykytBZNiXfabeEXmlBk0awLbGP3EQkgYMJ9LUFPlOyuhaPT0xpN
6dlPr3b8ZQsmlo9cKOK10A8iC4LfS5AP/HI/R1TXwvOtuAb0I57H4hcr51Vnfhu9
i/B70thEcS6I6JuwK4pqsTfsLGLjILGUjKkw0c7aYRHs1HbKkc0d/A4JK21MKuiK
+v7c+6K9lrVLWXombzvwlVoLk3+HPe//fw/qWQyVdSyZtGbBzVERTRfDCKW0s//I
yJhYLh77HeI7YE4IKMOlKOAgnldCxgYnIQBT0cfY8XQjxoK7KG+rr3Q/+Q18dMNr
2AkuIf0ZU86ijjILUZ8F6iwIeToSydWhWm2KGNwLkOVA0wIkwPmPn1MOyv+uEEYf
sGLAe0mlZsvqqVGOGyQ/SgzHge0yO/2YaxqpMxZAR9F5wsqzDq+wGwKNKPJHfHoq
btDIQyhoA79Nwu/XND6un3KWpNZziXqvmh461WoynfUXVvn9uCMyBPEeTn6TvT16
OlyhYEhux+WusAUW9xuUHWk0mNSKEoiAwEzTcEBHLes3unnqgCHygIoBQOAFyD71
5CFv+kTR+SuGe/wipmUmAeJ38fSdylPY7/z+jsx0V07wjlt4bXmzrcOkkJc/WHHX
U3whq6RF4COac7tW8fcS98hCoNs6LRkCaUSeS/Z+o29z/XB/hSjPAPIH1bmNCGRO
zkF12jhtNKWuGNqDlZ1E2I+qgPrbsydWmoHOzLPeadLmaL3sy87gkEgWWzibYiug
kNv/ba/n7mPxqP/12AyaXBG2tIN4eJEj3g6T4J2Dl9c2hZkPeOXaNJ9wDHqtb5T7
eXs6htnfkCD5JPu9k+aJKFc3cFMnjBMnYEqrEH00T0PnGEbONdYLvM6zOIHxf6Gn
q1VECg81HFGLBnI4VOiCDDxPE7XxESe5T0Q2DOdcm6U3gleCoGXCIq+sJUsvStCx
NsO4H2frXDR78BqPSL+DoCS1SkaJTCHpBrK26N/s4wAusGrmQbvVQISziYb3Ls/o
YA3SOG9no4jZLKJj6+kysCJDENixEV2MG4wOEepvWy5zzIu0NlDBaqUBPAr2yH0U
bz8li1BXYKA2Z/aK8nBdPs9lXMMQ40gQs399TRVTQKsrtQbKXwKz3Igo2LR3W1v+
rK3L4dFM0B+fveOdXCcYneWdNz682kJCymYX0wVSfGjVQIVIvGnMJfgNEVQJ+WWI
Pl2xn9vBfEZ0BT1VOKY9TUErc0Lq2W3OEVy54+whZvj30nfDeJzI1cp19Q/xr4xP
8vNmy86Gg6BqRJIXIIkpNjgfLIyBftEqZnErXUTa8D7oGE46WnrUhjLcfnHCzmmw
2EXTETRCgypWHxUjMQW5LqzWarsdCDAk/sjH7x3qTG9daB8ZJeOxsSDkLLqfhW+D
AmcHc6qb+tfoxJQoS2KyA9DB5bp8OSRotgu2YTVrrJDANvbeKrsK09a40ZJOdhah
cjbxwZOiu/WegQiUVLvEEU1A8Gc2W+2mV0+D7jmKkwskhRTTwjvckVUovfpDs+wG
aB2anBWbkAwBpkQ4xQ2TCU2nIhqRPARW9OH+3NkmtcaiQzLZuYxqKlmu11BX8KN4
Hf7/tse/Ou7dSiLu1eZ/ZUJhnQ1oHT4H064LPHKxJ3Jk1/zuvpURbKX0NqFauXgs
A0Rp93DJqJ4gzVm8dYZzVF8A5D1/l1d4nqNss/Lz5uJ8hvRe15J0FQHre72CwDKs
A/PJw6OjZaEkzUZR6WirnxqIGhZ9PZyYWhA3a+8dqv6817Wizxf5ZN8D1355kgSs
Y2m2EW33UmPxr4BrdBGJiRre60ZZAx4Sb0O8Jo8kQuT8FfTMaxJjVDiYRQUVZ27u
hg3gmjY+T421R7dvNstL4qSOQrHjrbRPqm2B0TVOH2M6311oQ7A7zF2AR6y8FfQ3
N8PvIkXCURJ7Xg+9kS5oYGBPbKINkBzBBWiVpEYnTQylmJsKP2ZVGH+oOUbceWas
uiReD2QS/945UqLTHMUn6jnpfbNWjraAY/vu1dJgXlRfTSlAGARl5a1SCBphkoWj
v7U0uMXqEQpzIIobTpp3L6iyZY0SoXmthcHu6QnHYSeNm+CtfWJAVFWZ1QarlHHg
B13AkVYi/KJM4OmqRRGRCDLhxqaP2lzdjZBctYjjzkmEvYDyy6BLdyaw3YudzTBj
y3bpY3/0WKEnOFR3Vs7Z+fJOfYOhPWAspz8j+/uq//yK2ri0cWyDfbhqF+sZspdb
iJVqHYncrRpUcwRy60byDmYs7l9NQCE663uvj3Vrn97UqdpT3rXcr2IN//4oOMzl
L5w8WE36vISZawEEMg1sIzn3J+MVHznpoq65O/bFPXsjeIkf1gr0wd+TGfga3w3Y
P7NJDscb7tOZGYRdnE479TxfkO6ivAQh6JpTXGU5NaXFL7Iz4KCg95yGkU0wJUOq
nPpMuudRwpQ+vH1AVXJ3vX1Qp0MHu7ckux3Tj61UMbAiSYLjTwpLuX3xgkjQsWUg
h1j4a3VgSdAP5/xINFSuLbiCIyGUlZZJ2EragAWaNwsJuHuPgdX5qyUR4tuM2zZ2
Cjk/RObsZUjew9mMf04TAMtzL17/2qsZAPAO5OPVkq+toVEZVw6zsT8rEUeXb9oi
jfy+g0BPqaLQK3U36MOBwaUFiEBZGduxzk01yV/as2mtMeU/SwFEwnbk1oEw3dsc
70lzd+BHpSVdDf7nlDGS+iwSAGdZdVG38MXQdT+rK73WOcnegTkVqsdvOPjpwORa
IDZkjeQ1KaghTDa71vHVhGAQafSAqz5Eq3sbsE8Vrt6BgQSOOOa5+fDH1tvgmPwn
Wk8YU6LT1K4uaeD0TdOuoYZmJARPWJybikAtqmuaQcDaB4RdxcFu8k+3iJKIg0XX
jVb5tPnPSIfYUsi5aA4OI34CNY5M3phvDZuOGCiOPXdXsH2cpZWAP/luIz8mMb+r
wG8Qpllz5l5v57jY1fdc3GxpDMXmYY6mbIoKaQ8PUK6QCXYDC94SueTrZ9Z3PbKN
mvWpkdcgz6znFNmOVuNuLpQfk7azGfluxA1m5b2EyfRkYNxkTfQ4NFCF99b+3QuP
Yp5uPYOfS9944ntzv+jlL3bt04Xsit/YVHUTxKHbfrhk7xJnNEeflr1kz2f7jdYX
XSULIbw4fJxuTBaYW+7v/hBybLtXjEfEiy74it5v/+UmEeJkTwamuqmJEukslOBV
i6qxazygUuG9j3aGpvdSUavcuzjiuq52QE020tsd0HCO2Q/+k/QOy+o6MovEkSKN
k4AOM/KgMXjQMNB8WINNycCsTBo7hiiJhDzc5bv7xP0hfWey4ePuJeg5sKQDuFEU
hlL6dWxKDf4HRPK0vLAtSXEKiMAnqYSr6IirlmG3mLsd39qc6bc52jpNZUCJ5MHA
cONJ3TyGWkWujAeWn2fPV/ZlgDOBT8iX5OUkc69AGgqwkXd8dXyjrOC0iuS9ZhPr
XRujXfV1WkfOkwL1Q10ptFcFhhIZlAqYsYxSk1POfR6HG2OmCuUAj0Bw+8yEZ42U
rkqMK1LP8YXi3dst9SW23l23hxs4RwpoO4XyQZq2jfGbuB+G64sHiGLVrwRYQTq7
RHprrKht5G8lfjRb0wMr5UZpYCLcGRMIo35+h0VclPwFngd/XYctti4QTJqBKCtD
QJmpUD1yPeZ17u45D0vlAnJAY3UgUhcTD1iWZ5ChxWzxnSOVYSEcgTXG1ryMZN5M
JvJ/KFaxK/w6zNr5bxWwhT4q+OxIXL03xnk8kIXtaUZQfHarlRkwsSDE55PP+FGg
VKs6ebT4OvHeij9F7VUPZ7LIZlHlxaFiPYGe7SdtgDub9h8mRSjVnv3tOCzPnF9f
LA71K+iSeU9ZSRFnPmFX9AjHCifKXylY5Q8k2FktsFGN0agDdsqDDL86VKqBxQkr
xHzrOGHz05Zn5utGn+L/uX/fJEyE5feYnX1XDJOxILBwVa8AqHzqtSdFGdbA5hig
YVFWMBRw1p6UxpUi6+p+ZK/jVBhyHs1jh+70Gk1t/UjwZgyo+PsZHwSAV2pM+kdc
W66+hYes9ahnDNDuNATuGYBE4xIl3EbupUNai9A+xn8hEHfavRXZPtWmNOBLTsie
8VXefee8U+NsJHfraDJzmEzWldcSi6gk/W7yD866WCnhPswoWb6tpdH0LK/Xn3xh
mfku8AjPuGX8iMbsHtquNFu+Y57Ao7XUvKcJ5fMJsXz9xIL6Y5QJw0IP5LayYyzr
dc3pRk6I7LP7SWH2/mTTnUaxoz1/84AOYotj9yahZ4Xm71O1WG3u8WE05RrFHCu6
yU0sRdoDsmTqy9YkqC4Xy7whJ47xczv4wC6k22F5nDnEZ3vXToIMXBPvMQwXDmNo
jJAtpTh0HKfVMrTHup2JHpEHIP97vmmNkFxsWgobJq13+b2Q/G94SWRe1kHOBKkd
+sR0h/1ij0xtIy4Q+rdIiIStRVNZFtYTo/Rj1L4UGRYvWg6Xu0Lx1bBg0pcPjj3v
frPouugu1ys6fo9cZ4zfIZRzmkpc7VA2cY53GwIb5C9G6rBOZkWqbk34NTmrGGhF
MwIpOSaZQIfoOwVl1WRcmGPgsgXYJ6JBb0sYzU6hq7Y9Kq9CBQ3RRPhxZ1VYmwWu
EwQdrNNPljGlrdDT4TxVICbU9ikBJnTDM6U2H9NqXVkpFVcLYojpBteqFRNrIP46
OCH9T/BbgoUR6zWAw8ztuxf2irnoPIt2iJVgCr8OLnhWMucYQnxVxRTFrsyB927o
3F6OwM3+fohvXFwa4clA8Pav7WgELPB4f/YrQAm+PtkZ5t5f8j3CejHVM+cdaPuq
Jz0AGZ/pZnnHm4DzBNKWUjrbQ/o2+P5XP8hODkTB+0RZvuYTI/PCTvxNTX4Fve+z
8NALdcEM+rsW3JhPxWtaAB9Et2nE7V/SeFewdMq0AStrPuECrLQRoyjIfVZBLtEV
3cNqnJs3Ycoqw/glsAz5aAmn8QnYAhkNfZ+X5+JJUEvmqSWvz1Oev+5inmb1/Q++
SAvUys9NFFrVPtd9V2oA6KToavzhcGVjYAKMksrvJIrDjvsbw22L17QzJUf+HPWv
Fu5MuOdu7I3XaDyPrG6imqL5JVqg8Dxg6vE3XaF8Bm++uXWZxp84sPq1BTc1rAV1
bmY/pfobZbAob9YF9VuWZ4Vp2DgdXPAbjwd0TGXdY8/0k4LB146WtFaGtfzyzC/j
tSviThcK0JTwU8hOxWb7se2CAsOm/qbfr1wNOQqhk9VepErvEyxDxr4iF94RuXPz
kNOkC+HPFZtlcbJS2Mug6E8OKgU67CDA9Hhdr3ImV4DuqxJmq98bii3512wpdtUi
3K2EfRh5Naw9JNk369aNwNu2bCqRDawsAfacS29FvtstIoFw0doJbxxcnCjB/L0W
T42NY9y4PY/bdHgueuNCyTYi2XGftOBIf4gm7BS02DkGHcm1cPYjYur1Q4riaAw8
lIs/9Hte2eQMXskqIaZY/X/JMBzwthSSPKuTEcZf4BUFoVlolLY3IVk1vXhW8QGd
Vwfofk3tehXb9YMyAE8bh7YH/+o6dAndWw22kZP+hLDkAdY6/KCkXrWcBHR2zY7A
Rje23rUK6KPn6SPclMI5eSh69ivViKpjUYLirOp+yC7fOygmiYIBCObUYVdnaPOd
EMMPJ7gWvU4I15633zIe+KcOK51ON+HY7QLDRvbXDOoOdbIEWS/irTlnr/Fwn/VG
lae2nacY34D2znj9cZWiiBzsLiJlibMVyoOHGZLYNsRsG/z5F/Zc1bPIh3qMZrgN
Zv5Z88IiRTeeJ5KNwr5rD3UrimxzwDjnHLLniU1IB6DuXRn8cMcBzj/6WrULRkU7
lXiJxBxUO6xnvs81+C5WkXb9ztmL/MvONa8hVKvMggN98S1iFuseOAWMY6uRbIyz
b7LuDnmq1LrqnoTiYUuRfVIB/CwFy1yuzgiGEM5+BLNRqXFZzADcYKyhB+XEJYpb
jJrAZ9B/rxAQgfEjTy4BM4xT82tafqKHq1ckaxqzUKGawEblu76wkleWQDemaBd1
d+fMXzRWo7RoxpY2Qns+qIY82stPokXyvX4Dbu3i2ZrMygLrn21LD+6L+8SYCBFv
FfyRzbLplxpjJEOxUQt6aK3T5e1aONsoMmYlC3LqaZo2ZZuRh28aRgTauvE2ydxW
wvMnNckGjtydPHyesAru47ueeAkbh3fN+EZIOlVji82voaCl0DqlkcZ6rG4s9Ghr
CCyVodGW8V67Qi3yB1UvcDRTwCXwBpwt5No9DBSX9XQVdm6N2AuMKaL6bUFmk1IV
AjHBKS6Edj1UchMvKWwiQY5oU4NkgalU33SMx4XO7dJB3FggJxM1VHaYwMBEaHVu
ST2wm+lWCYo0LQklqpchbc90Qz3WqO1p5b/Ppsuu0yUK/3w41EckNHXsOXkL5Q6t
Avhlzyq7uo0JwBRmwxVY8LgSZrfDRTkPoRulvilSnPxbQtueJNJQb3gsFn9HZUUO
sDr/ymN1DfFhfZZhhI+ml0xvwTGKrKATnmR70KkvfQWYUZIaetCubUitJ8SFXckY
w1fCWqBmlAd9gAdMwG4LZzu8B8eUMhbboK4GM8dMBdNv/8srC9JpkGmdj+Hn/XOZ
eU9IDBYBr0oAHvlzfaYJeNsCPFVbd7cFehq0gPvXU0UyP1IF3U/sGkTg5Nlb/1Vo
tetdJkdSYoNA2RzQG9HrRUEDp8jdpB2h/eHG8MWJlhWOc52eDtjCKjZI2DIVBRla
V1BcBpLqhYVIGsvqD+Y2z4I23WvYc1saM1F/3tZjenbJe3YCHGvnctn5At7dHDHV
GvP1v2yRFnEGGWOmdYtbIRigYeBGUH5b2UjXCQS2Q8MBiwKxBuTOxpkLcnkMowDI
l3H3fMU1ReQXQCu2msasORj6ag860KlQ0oo44F5iK/dFQaBgoc8uAPU5eMjOkS3h
kruKg8k4ftBL5eCqlMIXpEnN3PjnuafZw80zrGUAiWa4/BoGp1uk1cnFm7YCb0Lj
slEk3dPZJzhgaF5ugRBg55MSvSmP6maYmcz88UO6puawlGYsv/AqNJhCgijmq2Fd
BV4T/9eNmdY5BIR16V+NGG/rfYZcW6AcAxPGQ9C/jLcvbW1NoXG2FISjzzVJcBWs
/IPx+s6BjmiZKf/X/DbG4pyPyJXAtOBfhGu9GBc3sEVXZEkbsHlQ1YGpSEiIgSR4
eGWtmwAByQ6azkOT4zNTqyTrKlpGiY/GaBspP+z+xOCCUcYXzhaMnuKHtSpYelL0
YpdABQm5jpfmvmKvKt900c4jdjJL7TKt9bVJL1cgteHi8iND4zm02X4TrUr/UQE4
5jP25jy300AokL5NcIJLkH1rhpzrl17S32OUJaLlxKI8nvuFE8aDy+ymKYB/LBfh
PQkJRjenLADR5Pa3zJieSDJz0kytyUf/mS9P4dkI/sFE029dGIbKIziUrbBA4RZV
CWzWs8u03O0BFP85BXzhVMBLUVxLABjnJBFav2s5/5eGMhUansPoQYSRFqtp/pbY
6bpIKcHedRy5kpEjozvKsTmncdTzT3CbyLc5mhZ9eO2cR3SoYerkc/t0LROvkvGN
RG8PbxF9bLKzoa+R8Yd9LLZ1iptaMa0ZCwqWDfP5dUWrKe/HucwlAaAPQEV5QNYC
/5BZOXNb5Qq7NjLlnR52gci4g7MD5gfceA/6CT4RbKlbmawkBH+VM82w4Kh+pVps
uqzXgx2G9JC3LMjp3xkkj85JBsR3CJjgIj+q5lzXIEDjZ/xSBZORQ0pFfrRvSt1o
URr0BHJeTjatRhpD1WKzqx0+9i9/SoEX5ay/uKvG7y/HJzYJEbn+X/HtpQQ5wAJA
1VeRRNysCRhB31NEppNZu7cHklc2EoUel4Ycz2TEgzMmD/cCbrNa16jySqQD/pBK
hnKYJkXmE4HxZumEf8oaVyu3NFAJ7kSC9M+eFSoEPmzOSRlE3l61ou0Q/y+/oBF6
TjsYKIjwnKOTkIFys/40x+ZLpJjJ6S0L6JVKR3hy3h6rWfQ+sXZzg81RmoRrl/j0
AWiAdFzuFVwdCvKqXq6aD8+RffFRur0lUyJHdJAlHzaE9onWAynIyYdzh+GL5iAf
bTNXOyyUgqN902w/oRwlv9nOKH9hs6iSxmxC89CatwukCFNWqDJylw7uIFBDgjjP
El0Zl7PotHI89G+1DVsoSCUkE3AT2IFAgqgyBTlJGuBdBtS73tFqUsg/e6MgjB2E
53YU4TQeF3WLWpgJ9BZyPNYj68JL1Ai6d8xbvpgK+lDcafLtJd11rYsB8vPQEOob
NOTqBQBM16VqXOMMlIkluWUlMxND2xrq4AgVBa59OLsO+DzGlJgOJ2Qe/FFxBbpU
8f/sPCBD0sEP6Tt+ve6NfhlmqLEIVGHvwfqqz4IWFRwwrEtN+R+t+0rhluByYGIJ
VHb+e1gIqWt7MnwipXbATwh+OEREdV/O5kRy0UzoAbxzqtbqAp4qoXEj9r4nROd6
DiRcGPQr0ozNIbwM8SEgS6VhYmaPBYfOwXsl31fQ+2Y+xYG/kr2J9TeFqrYK3Goy
5gUcwrBu+oQrZk+EcfTGOC+dDzRbNz8cxMRFI4DOaBdmYMF5dVcaLcwMNYYw+j6t
e/9gXWHOm1Ztu7ywAkKkXCdGLR0EGTTtynHWuiQsfEUI1fLNRWsuO/j594Y0S9dA
TGgKqnaFEUYPlOm8+r1CxedIUybkQJ1LgZBS98M5x/WY34i7yHQfKlO11TN4GdDb
4/HYjnYPZCNq5aS6O1p/bXoZQNaFMMy4D8efI8ZtACoOmbXPeL9Y9OXPTxnG/oFO
L5QfXTh8bAxaexK3hJPYuUayyGqM2pxQyWa7fSrb74JQ76rQsVY7Kgyp4q+aRcGR
nENl46RdPDS1YMSfTbOWLWaQuI9XMdABlaTm0RGcVKa2T/WDF7DYeskJZbGTTO8g
zKmBIEfos3u00ZE8CnGxDipwGLtD3huD3aqzpv9RYZghBGUe38e6Kncpyc19JiTU
jSW4L7b0P4UJDHYO/t+AMOnx7ESgoRL6iPN3FAyUOV+gyYgdlyAO1B6OUoGb3c8V
cgr6VWhnZRRE67m7AjfBx4s8KV/cyhbM1oSpsiKPAzbQ3vNkNlFQDZDWlF/1rjg8
covOgUwuTMHTRyYNQB1Ob5pCIOedVRcEWTG7qeiCEhU18hQoqYhVHdXXIlfOpTSs
5Clds6tcHD9qnNC/84fMEHNqbDk//aUvOABcqKJIKQ1zK4PPGq+fyOV7iHCPfgRw
Xbs8KnSaWGkooKNmUeRTzqVVwDqZjKwerPuEtS/V5HSmjSgILtquejXZtuHlX0u4
fpLMM0yiNdRbbOPE0c/8HEPj8JZcDpmO9RG5UhFRP+GTBsN+8OTJcoDyxy8OSMpS
zb5taYWHi0vLdrCPDjLsP9TAT+rkdfzxY+43oKNaXNteE6ymsLtvgmEobf7vJQDH
+/4Aq1amDYD357LhBsqAp0NJbwVP7YCxyK6EUR8Bze415RWHnvR+sBYWFi7quFcn
+gc07xeyA/zOESAMTqwM7EPhTosrHOnbwJBnx8H0ri3q1KD8YJE/lahO0ldcPuX8
PkyIl3YLvjsZRoDSx6DvGXmCHhNXp6SGGqhbXtltbfpNMIIf+9EIckF5PV8194cV
Gfmd39LmCWXj9v3YIdHySQ9VXtpyNe4WqkS9hSWDJJn8edt9rtvPQJkTnhDFaftI
Vb9QsDCwncUEwvgLwF2TKmmRxL9pJFyAzYz2//X7ylWkaYFeuDJpt0io1N/duyEd
PFooXichJD+u9ldCsz9GVU5HnHcpUvUjamqRexFkmWEnHMpirq7OZ5/KZ4Q7Vf0r
zDHZ+sNRybJ/GBTRIu+XgTK4L4F6BiQ9U/tO71Mikt36n+S5jgzyrz7XPFqdOM8l
Vjt07scZ8FdshpivyXoTCKIV2JnyoSvGPQyAKuoDfD6MoWjkbkKK72wMH46OFmis
lqA3CwQHi5MM3F6lhJ3BxaLp+a0BzrDDjWL149XxUoposf6wC8EWXueMdcha08p8
kDY61iLP1q8LA6sSemrQjiZ0PbZzVyASRPSZ3tKY+Z8fYOaOX+SfYpgvHN5qSeST
WKKw8dTsmd4uNmPESneZgDLJScuM7b+lcGEDHULCnhMjt+ZRNYdl89+/gWmbgNCm
NaSPJJ3TJmZPVWb4OPnnsVddCUy7OdQjKM7lhTz3RPOoDkMDtkqHt1yMMKeqf7hy
fbhgT3yFJJJSG+lqbzBw7u5+uqZVOvGiOSoAHQLrA8ihXbZNJXvU7CUXw1acW8yp
XiZ3GjTNLdOpHNByiCDWPLSAzTUGS7YT6Ao80TB5wtLR0mtQrknFrZ2ZktFJYATV
IMvlci+wUYPD4u1crg4U/yCmfvriqWsCfNeTpu0oPFGlQwcJ12i0K0tLYpiLt47v
8o7JoWUqjXStWnsJ4ucL7dLVyzkYL252VSeFDJl7/wOGUlr950ukW2vOkuoCJRxN
zZySA1tqeQLfLagkn1pZtBpl0oAb8hlpLVe3nb6i/yyl7LF84AX/OH3Px0n5NkKF
PU+zUABBiqg0jMsnfHvQlaocY/mPFacJwI+3Pn4VD3qolsA1I1R1lqxt+C9/WiOd
jx/tkAqwoLuC3KF1ORVliyT7027+lJiSFUAfnxUdGjgIzQ5hxLdpvahbVsu/jL0q
OFnwKYr8fYY/TJ+QBajT1xhyOmhedp+1dVoVgfkeOhBKDYznTH3nSle/mHPSPytC
boBsQgmTeymqXIohVK0tFIp5pG5BHOrXsg0iwvnotuvGJ07zn+id2rrx17Y4OZOq
axiLZP+7b3MgGzwTMUmCymMilHEwnSqwExdiRM9PzxXanbBgjYjO2tLSe9iBqyyQ
C+rEO7+z38cxkhV8u3GLcYIu0L1zxzkiPLR+BXoAf4NCODy/DSip1bByFyM9EpkU
/OpPhFMEGyv4NmXXzM7wOW1IBuqUFFrx/O0Xt+It/ylp1sh55F80oW8klOUc70+j
+XPdtmPmMgB/eU3O1vDRFlhfTR96HJuk0Gp0hrg18mlMo5+0ZDkYAbIJtSXignJm
hV1Ui+Kq+bVXvTGowUx4ng1D5D0a6nSstk4llDlrJAlcyeQ/fZGQbrrmADodPfWo
/CZJILmH7sEJ0afxiTKQkS1NCAe71YFZI2yr6DfCJNI4POSiRb3oYYEfShUsW7El
565zY+dAdUyDVT7i+4jSeu3jx3jAMszgj8pBamBOrnflGBvoExc9XPDo+K82Tfe9
Fbssv0GoFywD9G0U3cC5VRKdjKkNQCgPTi/HPTtHEP3maeny8HPVoaE4L/Aed84I
GGOzPHc6fSjsxOYg5ExBXjL7/9KW/AHArEoyKrC0VRW3cJ9Bx5JjTwtwF8D2bWPg
3AdW6BXLyOgzek44wZfMKyV+wnBtXBLAfJpeiI/gaCQf76OeacXv/iRx6AnXoohA
9o3LsqRYrjfHRCkWJvW+WMFSdfsg3tusBMNMschdOFMXbEJLixhPNxHwuE0ApBYS
IjdZIP9eE9xBfF/JdOVfC/kcI9wdQYe8eHOlY4PwirYSR7pr5Rob8DGiGKeT5BDS
T2Hnmp2zh84kokSf/Bm3hc+3yUeMzpIIX2qihZmv+++313Qvdz5wTYpCg1iR/2Dm
gJmzrw1pNH5aR7/UZMG7XWe1kkMm0syB0S0Ipit9sGZczkOYXabQaDN5w35D55go
ILZmbTt+idPNF8vtepF4Twglwf4An6p7A2Wscwvl1hMzq6yJ63YRZ3qCiO4PFQEy
bQRBFFM31IZUEz7oP9moMS2NcHRBslUD/mrB6aYdIJt3Fh5uc2GdhB6OSTwYQnp7
rHTGvjpfQvJpwCkrx9M/1VHLETx1AaM+6ZYrlnkYNGiKYaXsS0Kw0dWzTaMtnquc
tfL3rRaZce8jXG2qlyiEnitwPBo4PulYbmFeeAge0kZH1UgleTgZEerbrVsIA4nV
HJhu/PfUZSFzEGz6VGKeeBybzQ35uzwEubRWA8gm7KoCAjmn7CBKSU2nJVsudDxT
YWUQG/vDbJNwi+AAAp5jAeYNFmPv7LiLGKeJ4BAs8K69C54kO3afQAH6eL+MZX0y
w2AQO3dpyQjhFbC3wMA2escsPsbsaq1/aRAAwtqmZi29r4IhRl12auoibVcQEwP8
TeRlofRQkE+vS34ZhDVPfAEauALtHVkGHQ+hqyeuilVmIwdPDWqH63w8G3hPiEXt
HzD0niNI0XLljilZo7KF9/fzDZEocRckgwbjAqEU6dTsa3npkvX/Nzc1wtAbszNP
mTBAwG3XZjS4QxqbYAkER82lYoCaMZtM6UsUsVj0abg6bphLCq4w7sE4OG5dor/1
G/tfp7UCVQ/oCjY/MKfHrX/kczIzk5MysbN8j5lw0p5JVMnI7m5HMYw0Gm9b2EEm
Gly6b/1k60mCzQFNs8nKw7otz04rrOfSLxUcgqZPaxzs6Lgoa/TT0iooBnAEa6cm
IMghtljVyAGT9EmxOoefMrEOcwb3SsGU71ib6eCHN5n4Yz6wkwPI+3S88YVyoiIj
1xM2NCqtxXaEYhrLLH86wVnN09NhI/aQb/Cp8QfeOS7FpOYJJ+nv3dxne8ZypB24
6HHeq7kNIaFGfoK9A+yGJz/RVUikpptinNR8W1Dp5qSd9IyadEB+3d5nydJ8CfLH
Qg2qBemrq/XoYwS0z4v4KH6dfBAoImkrNkD/KVGUwYTi1uvOhw/lUckHFWfPCpD5
c0VysXflK8r2YKTVAWtfcnGrqW4e03lgojlD0ptDdyZSkKNrnA6us/f8AZtubStA
pmZdVDf95S1TSksoJRMGKfaRkrGoNQkYfAVauav0zrK4fksaWeXRbDiUUNddpVuN
W1D08yaEXTCk8seqggAQRIXiMDBYXZA7pyQY637dfzIVlVgShnQt85nYDkGX1LeZ
yFt8FlDFrKaUEp1DcfFMmkqEOUu6NBcTvldOK1jj13XjWNP3rUIIPJ3QLJR8tk8B
uMivmNe+jOtyYDNSwa8Op64wdoSdU8wRdBO24RyIfK0cbbdTH1Jjw1LfZ0KcjFg6
BFELkOS4i5XllmufSnbNUPmcNeBaLSFuvPoSieCBbztVy3hrtsQTYTYpHmsbchOJ
Bjh8+Hv8yyR5ZBO3UtA3BMvJBxHyiG1EZuknrdVCaXtfuTfuG2AuKywK6/XqMq+4
8XylDBXpa6ucr1DAKAlMEk12/7xqHd9bNOZevKYb8kFSMhYK3perUIEzOT2+JnY5
Fh1qhSHLLQK52Vu0Uo2ZbAVdf/Ws2oq1eth5OT1aHi1yyTYU45RXcEXKSfpnMRFn
cRBiB0Axxo35r29ZfpBXHcO/EsXV1XTPYghN2fgF8aBK4VeWYDCnW+hz36I6JQQS
3xbyOartkFG0TKAa4AoSo1XRlpjAq6hSMnWa/2fa/ZqnQ9zRi9tt7HS/7Ch8dqj6
hEooFjf32fMeQSEt+uKpN+mF0S5ZfngKHHLyKK7+jQ0MJM2UEpwUJjnsKyzrsNcY
uK49ZoRvrY1W2JIxopNKbyHluc+GhpoK0h4CPwnuTcwuiL5NzFSDTGDmEJFj1fLt
crgf4FHeYyPiIqwPD5EY7RZIZRzdagU7U2y2jMZc00azfdtHCozRQ06en22eG98E
9cKDPDsEOPRoMO3iRSn9Jt8zfPnP0wr0Y41M4d2NTRiras0hIxIH5Dy7EKINJ4XP
71PVUTq1nXTrvf2EofcSMPctLt8gzP0i3xGR4HGN85wNtAH4Dwk8eAf6Tdy6o7Hu
n0+Aw63U80ljbOS1GJuPSmseE4zL8oxjgRm27VQWe3A+EaTMnYcGBwjoJcUX1fjy
Ic0vkjGUluysIFmGEhBu6/4K6JSBmXJQqcgXIApu3Xg7pn7NPlZXShzQOrqZje5F
yQ027ldzCMN6r2B8Bmo/7DuB8R6XRpysFAtBfE1T0tk+oi/g+My023Av6D6Qg40o
/GYhXqLL9hJoDycwMMVlwArlgfirbG0Ld6qViOE6YFj6dgOcKN8aWOK92dxowiye
U6yiHy3kDE8W28mgoYL95u/hi85kjWeTlaCKO7DoWTw88fr4NFdJWPjUh7vtFWUG
fW/5aTsragsyY8TG6D5Zwpmkomu0UrawpYXBq844iAijnci7Z3bMFnqd+d/slLfX
Q4RRmIzhpkT8cRb2F3DYdzrPj+fNaB2yEEi1VCu5zDYrog74gCeMaxXc5H5uesLA
Z0glDoiaWThwd04W+In1tTlzfQQQBVAK6d0A7BH942nVrm5TxhC/qpyPnw0yUTGC
KX/umbrCr6twZVkDMd7ebcil9gkbr3dzHjrnY/OJ22zJ501RdRfLUweEQw3PCR9k
kyLaCOxuvuTBKiFCQm6/GOffNgX0ySCAdtoeCozB1Lu//FA9nnf8F0hpk7zO+G7S
x6aSU7Dp0LzWH+/4CPMFcdL0+I4olkdoZIA+TcjtT2q8pfygrjLusdLql7Fuh2Mg
upP/yl51J6OgVgw1+1HFZ1oebDsTinvCxHkYRpy4FL9OZHho3KlSHJgaUk2gXER5
doEQdIkyCMkQtlut2yR7mwNFUfK1ryTnu3RdJF/YVVkGwgaGMFzbzPEe/wr9doSG
GSYDSL8ntPXTFpuoZvGloNFuuqyO/FiZR2XHGifFnLB8l+yV+ORsbLf2Ju+VYZFh
3NhABgVJ4eNqx6CIe3pfv2haHGnrNQc//rAaLkrJKrG/rXHZM7anjnrhoUUuF1en
DHywvoJQodJ7HcWs/X/taaMiODCzxvN4VjBzpuKZ3elZ1/tLU/X8N4fKD+LDomh+
aC5nm1dVnzU0+omxvauMBedja/pc6IGiR/gUR4XE5l2JGPJ2UW7liphLhEe4TQxt
hStlpp935XaCC+5K3wcgGM3QWKA1B0GFSE9joQHOrUxvQJauAZ8+PWBXYN3lF569
4yGXnQcRjgYAdTAMyz5ks00Q0qb+dQKgAu8wNtCyS3TLtE0vOghbjjSj8RDlXRLE
Vx9kwEQQWEtcYSi71DoieQICmDlNGjtcfceldB1txoxqSPPmkcMJFz+UlZVgbhn9
aA53AtGnG5ZEFdFUkWGve9Ai1gnUtQnRDilPC0f7VpJ/ApExGNDYKhOdCcuzJaUK
7lXGp4EavnClREvmYavjpG04OuV18hZyb5nN9MBS6nS/v28UI4s+lTq8KnLYv+wh
WmWy2ULLZ7WUiVBx6tb2GV3sjEyrZSVQA7PNmmhI5TShuRaRI+Kcq+Er1HRBL+10
aKtrcytis8bgb8aExQUyyadC15Tx9ZFtr7NnXrHBVYsSvJgDJZ7HReZ+d4VVU7gV
RwEMR+CHd10/7GUjWP92Kzz0iyYfo1GQ5cZSp0jDdPhA6fKlHXFuyRH3/X4NaxRm
QJ1NbMrtfV8vr6Vyj7rTOjzUln/E5EFHiDpA3QxbNmeHLMlLseavFOXEYMh/XQZI
R/CiKydVNOTNrgPP8FobV29w0Hdf1/2uoUr7EZgR/FtVfE2zIO+A6lCZlUOBKRG0
ZI0rNqP1VFDKpLucGwoWiqm5LIbxf78sP2ivhYGa0D10xgrRoDRn8RUc9OJ4FAHn
nmDsJqjfbUMKuBvwkXPjP4BwQFlS9EXy2P9I/PpWYUlubWrRPvbhM0zL1M4iAI6/
2G9NFGzF0SJb0BrPjA2eoEWyUQs9CxFnOt4TsG4xf1TKukBoRHO6yUAuEnNB0IZ+
fw5qWIuz9CBH16NcreIP5ufzHaYCsCW5bWZAuF/dMRcNaPWUCI76mJLROwTfmyLS
uD+7iOqLjzdNbi45fm/bGcm2fcfyoAOl/IVoI/uoA5BLzR5Qtmu/9ub/1bZ0ll+o
Wb1R8TEKsP7iguB/iaYfDZD9QedpW+SZEUSoRxWdRkqtXuxhggmIOr2Ka3CVwLp4
DV3q7EbobXafW1eyQ6VvZY+s2Wz/FNro9zBOr4UkCBpD9KJx503Zt0XVC+h2crgX
5EWcy7ufe+DppQ8IG15nB1NdT/Z5eXYKc4nLSQl6aL82O7evNoFsD78BVl8TSbFw
iWfXotMJX7e5/g0ojOowf2Gi4VdlmbwqacA9QHgXmFZlHh7Wgwrzh4yHbBP6D4si
IpeED5CYU74YsQoi1mxMSo7lGLgeL8/0dgbHVfvH2gS5HGI1xz0Nki5UxrMXKX7t
pVYRZOotYLWhWv4HPQNKj71mFAFNU4JgLzk3FO2Mm+XR8zUTOb3FE9Oor//IuUKn
iyh4mrTZMENJlrqTFkB15NxcfxrywCCzdjJFrY0MBrqVB3t3EvSROKZrlJRwHedE
HU1GAhXR20fvGlxAf7C/EMyakwYncxGDS10SzOyGrV2t5AJrBmo3okMNK08F/i9J
txHTQqQeRPiUgMd5LbIgrNLwraGsWyJxRLTL9aqUDMYn3onlp4PIx7LrDNXhcv1J
K05oVMnD2T3ixLVUt75RqqP/J9K3Y8GmxbCGQeyZ63SJ1qkJhcRRcOM/P2XT/a/i
Y/1l/z0/3YSigUDSyQBt0tS4AkMg+08f/4yk3C/z/USpepq3O6eh9/W8T5dJL4jf
FUFa26cUI9kKZ/2DlMmcI0w1rhk3UrDPZB9hJhoJqVJ81a3PSIbvJqper6quWR/J
yG9uThiu3YHmWT9m2zhGPRMcDPhC6YMQaXXOCDELH6f+8oRjmcbl1iCw90HkXFGx
68CKq3bmdx3Xd7vQtKdtED2W1s03dMM6Pnf3PhFpFnBAkXNvTrprkwBaKsBv+2UI
miOgX7baUZg9IalzmAMqAMg/zlehZJovQ9H1ig3Ne3r9xppRorhMZUPLfLZgwoZj
yyWFniz7QypzqTYf7TTgAeI84FM5j438hS59RvqCJtYgxzoEyccUxDVWIdH1uUYO
1Os2BO2NTZRPXEgyOQP6rOOcLMj1gw49HBbyvzvV0GNeRn+n07F0hGFnaIMnVWrY
8grut6nkrnD8beuuVCyrGyUJ8Dj0/CPG4vs/d/Xcj6RmwZA1NLJxhyAjz0tSs/Xz
jNWCCAG2C1WsKGmMPvgsR4avelxljMG2eDE1zt4OEl6O1UvQJ+0uTEyqF67iW7KS
WXta9M/+pIP5uHir2HgxbHB0F4c+RcGglIaeJ3vy5vmbQgvQ+Zt3FdWAh7g6YY1c
vGs03HxOVwsT9y/lF4XExkS+SFzff8iMmRq2eoPI1qcUvrFIvXvvXCTbdxgVok6M
e7OYPtGr6ThsSUU4VtCNaku2QbB9vhT0wkQa00jbr6qUCd0QbOtUj6hooCVQ7n5J
0eZPvSoQpRBSedNlmX1w9b4H8eqet3J/9+Rk/kWb8wARpyHjCbi6R8Nbaqop6hyM
Xt6yAT9213oivEcmqf3+/f1XviFaYxBjX6A41ctVJZiN4rESCpeX25vwpjwre2VJ
BlykFV/7HB2G/iELts20Tc/n122qLPxwJ4MLg5dV87JoSplZQwHC04XzBWzNLWYB
cUvJdrtDUManBxdZOvnVKKf7qhLYvqCUq+i4flTLKfbj7+7buKxSquFW5Mgshpsf
yDOhLcTwHpuhbW2URYBJryT1QV4HyYezgdPNxTtjt7XXy3cDb38U05VOQFVb6LBJ
+WYHQFqshzFhRGOSWppcWV2cEjsgiO4DGqcKvpniJXWo6SHhisgB9OFCRgaVTPNR
T6AlIBeRXPEnpimnHzgALC3TjzY9t8AFv4LjzHhFWPW/BP0VbltBX0KDf57vruME
VeqGnRD++sRlilto7zejxdCgatdCfmJdNkn2bLz7gpODsQdBTzy82kUzZuVEJXY9
sXKw2i8GnnNfHyj7SO2G7pfnVwe6PSjVvTApjY9W1ZnCST8wCa48DaofEvRCB866
eF9HdKAY1RLmoJFhA+x0oBl2RVpAPBmtw73vnLgmLhR1sxx1/8HYbXpwEcaBXB5e
L/M2adVDy4UU+hEOmd3TBademIe0I4DHZcOnIkYbGsLubzVbeIrSi9vhY/8nA2Eg
3zMpXyR62CsWGTIDGUik4gQzWlRPiSkuh3kMc+Hl7BtfxExwiig58uVARElmuFJx
1D56ZYnz1Dmztico+9fg0lX1vwu0x0tgAbGOpzIIkJ9rtTmiyFK9Kbk/5FmCl48U
9bgYJMdLJOD/9L4NU/T99Mju8oxgHU0Ev6VdqPfCRUoGCeOGXnkZSm4He6W2bu83
Rr+GuioRNHykfaGTbjb+MHuG/TELlZOKVBFwMn0UqOMrCHiSTxjwvIxPACrQLnuv
NRcZoJiPxhg5FdU1dhJbEY8PJ5/6AXVzJXIiQTzpjDanK5ohsbMVTwnsBg16v+6D
8vrac3cBIpmddxxtplQlKO+1cDCBBiEOctvl8Ii4ThjYuMAyFsINSwRi1KDU77Xr
3LWCUlwa9XttCpl91y7s7mkMy0Y0Pb9W/8C7iY/piVBpVBIQJxXe/0mPn4ySfRTC
dTDbCY7wGTdVfA85xfT+4bHkb7eI4YcaUXX7eyjrfZuiiVsn4K37EG2Dz2HrM1ZE
0u8fa9p7jiGqLvLdycJfFrVdekUcas/krKfV4hjdU7bBiZVnSZeICxD15UGaTZbG
sLQksxQIb/AxlkcNPjnbq0Xj4vir10DwtKPFWVpgE2oZ3311162z6o7bZ1817aeX
D3Ks6FJiX8Wu/sMfhQgbDnLO6UNbd5FqeyzJAZ6ZOAw1bmyCP2DewqDbpr4cks64
eMeTQFLJmhDYWuvu52rlDkm6ETdG+o/EmNTFCN9/Ow9PcgMeQwcGuwjqoxyXwTnt
cbk/lfSSlR4L0Dh5Tgjs3sLTZr3AOVS71CxEUCJ6NaFwJwsG2I508203FZ1rPsMT
MytK/eP23AL3R2LkGHTyfMt3cfTH1rOr1bnBtiph8rArs2LZjTr7Ng8AMWQH2NEG
jmSyl+HrWxTd4XDgpx9ExO+y/H6LMnK3FOub5/Q1Xbgq+9ktgc687aU1r91bQ4q3
oKWBLjr5Wd7Hk1R+WGKEYmkZ+BrD0u+Bq1O0k3h94sdiO9ak4EFQR8kOZl5AvBck
Nj8Lq9/svE2fyKf7huXxl69n/tvLZdt7qYnTlcxSmvH30oHAdqzB56xGd8/e0I5q
cQh9btBaojI0nuKbJMJAWGJGFtW2aVH29R7/GJo6S86RQD0SMYUbrJp/VVzKc35X
J8ZZu7XtIb9RD7CrkmHFPJ4e4PGmcvfSiiksgyYqOCVYmvbNg4yRiOU1/7ECzY/P
Wr5cWWxy3tNvbvlkdnUsBMRL//pJTAm1HWNb7VYvZwrGXIwMHc8KmvbhEI0f6/FE
1td/R3y76gjL22ehK2QVjr4WQW71XWZIAn1CdKk56whdfdux3Y6+931QTKEm99xk
fgX8Xr7bitELCiynYy5LW8R5RlGMq9i0dCm7Ai+uO6rQTOKcr32ccU3Yl5B8sBRZ
HucQ64pJPygT6XjLYaSSmhxGr2EdVO5s7RNKMaWqQppi90nzy2WzV9ngeWeXPhrq
I5ZgTF1x6pS74fNzn9pLfJy95dFpbJ6BXbVYCW0mNZrASYADvqTF5GVOdhJxsp3R
kcqZjgRzkmKO6rIHbc3wxu4DUERUfJOd3JTF1Beu4mkanP9b4tAQWnqsa6L2Hv2Z
q9OIiYgZnUQ+4ZtvGGSML/tKoRPpAUBsh9zVyOTlWRuNKPPa8E+aIRXdqzwR0uI5
PYJWL76vnS3FKwBgfALdV/xGuRQti6Dd9E4StjTagR6qx51W4a1mu1yd5kkxrKS7
K5d6CsXM+RLLotAEzBNzSaZkGWrvTP+Y7cnaM8xylE+qAhO8fkj24Ha8t6sDrFAu
/WGkozlVYBB5MZqViYWFDjbz99OttdGYIqq8PVM8iN4xfoAYWbVP7mJ4Rms87Oku
60eDvV3acV5XVG52VLCBaOgndqBNzI5fAY8OIBQfId98wRg7ULLcvZv8xdODFXLb
Hui7JUUQp6RHxKDu2cZgjHFmKPfTbrj1ks1xa3Xr+c8+rqmf0xtts7ZgXE2FacyI
PGBLcj0PDUhZfrqQSciGZc1lBTlV1uJ9KcYvJpLz+l8UAOCf+E/5fAozImjqFzVL
ObNwbxlU/kYyu8P3Pb49IOGMAv0v4/rLxZi9VgsRhGgRoG4O4SVC6bV9msRRKFzC
psZ02xQjs7QUETVqFVhBcB8mg/Fs9Kuy4TAKTVRoz5IVpcdO4GR5TbyAX+i7IVIx
+63n6ENyNK/UjgHAe332CjnKFcUvH8vp3PJwCC3TswFC552mBS9/7zpc1DgZs5ZM
gWYRb8aAQkOeYS7SZi8ndD1ShRZLxF1JoIjhoxFW/ek8nTTfaUfjFF6h1n66+g6N
ktAZPrBOFJaGohYUX4YF94IGqq2kBfQEmE3GWzBw4+7PwEqWab/nlB1BGzD97BTk
b1A2yeyTjrH0RzPO095vg8YcavMe2rx/ULflJSnEcqDs4fymjNtFq+PKAwLhAWwx
YuCsIJr4NxJ4GK6ESlNNZmlaaZHGgqNJJnx+cBGWi0l2rFYz9LQC859V5JLEOuW4
48M7FeYkk69jyJ22BX/SY5Aa0xunC9h/kn+roeZCldKjrlCDZLurFBb+2T56eEl9
0RAI1EzaqmNWjAk6BWelcmwBgQL4BQY2rO7rYIdYdpez2z3WJCRNcpf9alNLomNM
OeLsI6pR1LaFrudT7Ka8u96+XhOwdMK5XA+2GVddvpAn1uuG5uT7sy1bPkPLPZC8
l/aOvoTfXZTrtqHXblAlRI8ci8yR0XRcuBkV6Ci6KHM2gpFeneSDVndmyx+BWv5Z
9FPb/WiCi1BIPv6wvQ1bw3ciFZXvbRTgxgbcMCxw3fRkr9dDJT6gyAe78CvUM3MO
ppaA0jkthgtAhRjggcercJzFK29XrswDnB3SvqKHGE7hbStwwSFbdibU+LTMG/Bi
NNaSBN6hSN1Stu1lr3MpnE6mwe1R/UdNllzPLlKG8F8PVCwQbe+GKn0an3Jxqbbr
ant9Qt0aNsdAmeca5gGtHVqMZLtop3WbItabypbHIPSnVYahkVhMMa+Hk51FKOWb
dSzFgodjUAtRZOM2HYjM5CYKR2USr5GzjN7dgR+/tQoUScwKwsw9KwfdUXZSU7cE
IKvccNHGyA/kM65oqChleuDBdCxBE0gKQl03MD7EHJreCm60Em1j6f1RZyg1ZJ06
cSAtSRvotLVxFb3uLHic6fAXipBrDH47Ttusyw2vGZ5K8roAb1ZaLnlSGj5lepGv
FEf2MCJckKchj5qkzror02aYOLITuvxj2kkxzDRGvX1bVTvo/IxBXL+eulXilkeA
0a4EhntvDKBAw62pJTwwEr4YwGxG9xUNL9Jry/bQkOt5VwcDxGT6Ebb1mGype7es
1NhewJyIuUj4tchlbrCX5v82XQT+Q2CA+kKL7w0Imdkwiv3MNuKDrLiIhLCBR6Eg
qy4ba0GHihBJ9kklMOUSwYJLNJ8XSms9eswHbO1NuK+vgj8sBBrXtBBMp3VgIil7
WlRGMNDEXzov6E/y84+V9bxIThqKb9ecl+V/uKoN4hy2LYclQuyeAk03GWkslgB/
qHP7wby1w635boaUqtxwPUp9//kqnyEkXSVQPuPEi6eeLzsOtbzdULBVDpaPdH+3
zg0gy7THs2N1euJuLD51oiIq3hasSQSfD2BenEpkjKVemrB3tr9rB8hBIwl2Z7kM
+kBbzhZ44yJcijcsM25g3Y7AB+vLbEQwoUZ3TTlm55Ie3oZ3GGIJRGtcAv0uMi4k
YLk5bQUwVOF02Si4dQGZcoOV0pp0PVRz1i86cNjGPcJimwS64NED6/PxrQoXmP6U
jabr9EIozGQutE4nG3XFXl/glsozg3bi8r/PhcuLBzWKQP2YH1+m4PjcHgfOyFaH
/OwsuAB7qRH2fsnBhNtywc1xFdzQInwUA8iFiYE5FM9AZJ9Mki4DDyGNG/fmcByN
14gVEAsvDm+74JxooJYT7dzhHgd117XrQQKChOhAFYhnvHPsdbOcEWboYrEx26TR
2MRrIAabw8FX/BTQV7j2au8hiHFnc9cNbsZ5o0V4Q6CvtpvS5MLwV1A48XSldEbG
Y05WRjUvN/9f2ZJCvbCC5T2RXWbHFUQNtDyw8/XeoyCRKhY+W4Sl1XH9zVZUC+6Y
8lcwzPCHziWh9wN0gp53iFVvJbvtwdswsZBVA/qc0tyC/OnIKL0ZoqrpChyDz+dy
bMx4UnXvG51zQlkLn/eNxTQ+sA5uynwhNdE6lod2rE8syyiR4KfMI26yzf7QQEea
F2bbKH9a3SYyTTI/qglV/XL4AhN0duUpiZHHGN4eZrL63JSdGvXIA/5ZYgby3vjd
4NDicFIS2dOhKveEaYrHpLMkgr1JlKXdkhODuTppYh4c659SjPBMM4H0dO4uSCj3
4jOtqFWoCVIwBDNSGn0mGbmDH95P+JfgEk6BQr+eA3g1VIrnVDGSdUiGKCSRFgjA
f3UsY7vr8fafbh8YRsp4rSWTQh34glTEfeSJocS9BA6PV5cnx7rDsFLQNJ0YFzUB
q6qalwAlpj9ZDvJhu5ZRTlf8m1VYkPaJteYCW/wvT4ULASDkXYMRgbklJl31S6fc
tYzAlvProbFlTxgURV2IZSun0WceB0JO3Pnq1pFacIUYiKjA1eGFifDk7BA3xsX9
ciWQQwYFwyxkweruNJRoCwKYbXyfX7X7zPdCVubkgu/jo8beTLsDYyi2ujUpQZxp
L8OjAFzLhrfI7m0BJZ5MxVDa+GkYavCJAharoYY2abVpbuhynLt/61Vwa1k28wzs
gGqDLbUK/fw4m1s8Li7g3LYGnvAaRvwDXhL1vJBA0NpGYQ/jOqBYleOLHOGc59n0
u1L3dgD6j86JCzkkANbXqA9lAd37K2tTJEv1dpttlKAM62/KhqieElUleXOd/em7
+TjLoz3/4yz4ThtYjXUPDD/F0/gZQ8Ykl2xbEjML6+2iABdU8D3FCFiL9ZOMzD3W
QgoD+D5hjWwawgMJl08Ko3D+Qm1r+VzIMk90RCt4xtoxBZnEgrMYJ/RwnFB1Vxks
OGLQtFWrqkTUa5hGLQcigwYw7qhmeYgv/CD4sSEtejmRdp3Zh8rzPMAJyV4LhDpa
bQrE9/ZZSwxM6H8mUNcc9OHA8tqk4HXgteAEv322vxGOvKTpXoZhYJs7Q1KzueCx
hgJkWJtXjw8XbwdQ11jkT6rB9IJVnUOjrgDapt/Gk1GJ2DSTYHZWDNFt6nCCIPpM
fLDhRclqgshkBwq+eIjb+Ak6oReAbZjbnP5BYhZvxgs6EbrQQRsFaUblwVBEdgwj
5aOjnHMXDuOhXUuhoSFyXS0LpirC8MYYdJbV3u83eaiUCRvp6PfCYfvQt9hlF/GW
HnuG/4DOOG6wPQKn02ccp2rQIIN6UlPLltHKAg1rH7qHgvEXGxFMX7STKTtVaeOH
e2+H42iXUrKQBlsFRd2Tfid4tSKBqGWOqpLZ/MRExnaOiV0AHg36Q3iDohJlfkIX
5LCHviQH7FLLtzXJXr9NSmeuWTaQQH0XhbqdxpCdkdNnaRQFcIWrsINJhwikQQKp
pvgK/UbIvzPuuLlQCLwYv3GW4V/4/oBsrCCfiszAHSl6SDlcewv83585++ytdXVl
eXnUlvE8QSJD1oeACLk0sFdLC9PnTeoUB2LHB0dj+PP3OYAUrjbQIHp1drgbEkzB
zBc4VVj9eQsjwOUCUjplUoU1U5WZ2dB0uDlACch16Gz9NeIAVIBE05wWemNzuzRI
Jd3u5uL8unBf5V21IueBEZA8iAbZwSohkfqRFtWQyfftSbKgbxafradjYSHGbFRX
pAhAfKZi7QApLiOksHf6eqmKVWJaTUcxfGfpmvcRzB+jXD1OblnAUJ8UCUbfyGih
DGSEKaBkmdgZQXCvv+AynKwr9WknFjidlTfYyKhZG4LS61P7iphcx8vGNnULAXAn
MpdmA4mEsbxK70QazjCX9lFy0slfRP6Ae/xInOBTsikhacAKxUhcx16gEnrfoleG
XVfzmQJL6gJ9Sf0WlsXmTa1ZddzGyqS4Qm1jAQBcNV65H+hJ15FNRjuDfutGkov4
2JSxYj7opfjNNKhZxIoB/L8c9AO4o8mlA9IPTlUNSKuDjyAefQP/ptk+dNKD3Kzi
JB6AxPPb6+cousSKCg6p0fEjkZ0trssCfWTF1/7gUGH9Hxymk6MY4w3WebwGDgep
iJh2OyGc98o0+NKkzGPaeOqohs8jSegIjTCp0rCDC9zPAvXamUqew2LciS+5iw80
mlY9VuYB/c7wue7jClKnYtnWAC+EpTYSAQ34P978cfgaD06Xl4Wip/xpOjz/03mV
wW4QKKLatxJHcDWxq5IEwYjOk8m1rrsk709pklNc/x5n7cb5S0UCmxWGnMJ8EgG1
aLejfVgEKpKgvEHosg4E8YunfYE7ahSXPtpMtb/yCCxwWOAHPAJxRc76dsTFVIRe
fz/aLfwI9DSol1qSJbJukdGWd6MTARcKwfoj7uHqnMhBrwDD52va6YdWRNSP/kMj
ttMB7RQsfb46zawzpcinrn/mME1vn6GhHTlmm3bGVwsEr4pSqfptBeXI6jgf8nDc
77Va3qpqcPr/4fjQW9B2RdSxAUf/TtQPmljdOd3b/+ffpotbXYMRWeGijWwnrRvB
dI3C6un6+4qFc1bedYEPPRzs9KIcCPkznYLdljT8TY3oDWKpDDsDO1kxUULGww3q
el0H5ApvcXA93n82iytIGZpQNYtl+WnjUvJnI3FMn2aU7NAl+7JoikmgLzTGV/au
H2cpLDPpwFNRi83lqjJIEQeAHd90xa5o5GfaI66Pck0WIitJ26ixJhVUn5HWYxqa
tEY6G1KBrO4GTnF4+AWG8DbkbFljphGqdII53fArIea+fPrxIFTVJtdISboNBP6z
1f6G0MKX0z9UGEAwI9RQ5JdUFR2ZbUhYczRwn5+Cdt49eUtpGyK5mm2cXbhB2eHb
1dnc5JDS7zrHfBCfRB7yT1MXNigrybqwMaPisLQb1g4o601F2pI1gDs7pgD/yyR4
CEsce4Vw549As4rHalx5Lu/OEW2ikT/dFa8TK/M4vBGl6akuQlMQXz6enwtQ20o9
wOwi11wge2g3x9VJgwjSe8AEbUtwwHWsWs1W2YLwZRDrYsycTps1/8v9h4Egoi6a
C3HdJJD7uAnZWR+Mi88M9ievdvwyPLAY1Go4eK36NdFJrIqjp6WV47EnYCeU6KtA
WCdDZsyajR3IxApyT57Pu1uiwQ8NrsRCGw6Xr9Wp5s197gtNEj5O1lDzaeP+Fbao
fSA81yq0HTAWafhQbjchp/A0JR1+Qjg8lTq2EOBh1mqZQeuoGHnYMExEmv9m0Gqo
cn9J4czpWli92uQgvFzHs/8yUfCjAHoQB7w4DVp2+9TPNWhCLDy17kKJv1+JcPqX
vweqhvfnpNq4zt+RZmS7e66s7pyKqnKkz/Kycyl+IUakacw19Iew4AguLkmcSUxw
v9y5mMJYfwUnQAuaJQMBa+Qbf12J22HjhcojGOLYZqEw7h0p/jd9apokKd3GM2eA
eTi2L+FhWZZTD6mykMaN61JCmuYJyNtpuZeOG6UKSABNfLfIHHled8DA5S9fr6F/
p7HzLxhu0QTF5P9LZcw1eQHZCeZMI+mYykahfFyF1g9wgYp7n0rZYKMbDTtmwkyr
P9iTM2mTojI3X9fAQhAEuatZ7nGpzem3lmOJzLmHNVYOiEIq57/Td1+1CvsqN2Q4
jYxECu0/6gAgZTddRwI9MOZLfPEp8x2m9uBgwP6MvSD31SmNtJH09rfkMr9eHEU6
vVjPEHZ5yO5lbnlT2uGWih115AcR/6XVepzUc1sHBr5O/DT9Dq9/BuwBlq95Z1yf
KYcMH1VYLznrq3y3OoJ8UYjAN/oP7bIzqc+8aKC9TLI6rGaOIZamjO9y+EyXSdvA
evCQlQwd4b0Fc8eOsJqLpuk/jjgCMhaA3Gb1ny5vzh6KSpAU4c8j8KCPfxrk76vk
e65x0TQFKqya4tN0/YBrpEXY1zw41x30UjeRVtCzzCM6mzo4x2J1c9SZZm8g3s+a
QsaqqU7nCy+c2ZO0yAZKoLBLstqRQRkCPoaMehT1nYCDK2Tlrm0bON2nYB+7/tdl
RVfhaf+g9kE6qCRE1m9ceFWfsi3tV59H3qAyaPAnMfmKdH5nFhqWDCg+UZIeolo+
4I3ChTgnLgduQ9rmLY724HmQAVpyz2dLe38zeQLLnGL9sF8mY4fTwYWgqBVQ9Mvz
Zs33+uuzCAfeGx/hJjYowfu6zJQVzpR0kunL4/wcb7JgfxPuT+vDikxyqjkUfuri
0qV2f0AmVsThzeKTIbZJnHoFEeTJ0bWm4q42z9pNjggshV7A4ty5rqphHnjPVsXy
+W+HyeLojEJ5jRB9CzToLLmU4n+xNOyYTGjDKc4vs08kYdzaUZjqfvp9mhi2hBEP
DDes54P/5rOVznP9U3jLhfFsAl9xD4wsr2wLe0GBOLsZUGVXbsIsRUaB7G07/2if
Hjen6HnYK9DfbHKfwpRJSEzT0vTrT5KnXc3SEbwknnyOO+cGT++u4+zcvFD84wxP
kXYq2thzryEhJLhCzdkt6hLKZwnOCSpn0tfSSY8GdIu5CPGB3Z+IiUm04U9qNV18
3rkDD7kwZ8brsC/UI2JBuqcCWEg7YEvRI1TPlEEbKCyeSBoaaIu1aq/IP0HCxA3C
VOmD8TU/+wApwznJvVDDUnObftC2f/opAnEv+JQ7OFzOYEVdf9UHMjWAa1d1H/Sm
8ZyjFZDCRRO11kNQwzfRFsl0WW+tHVr5SVHzApcQjLP5BDz6tW7Y+aDoLkAhc8WQ
9vFoq1xr3/CN+H1gxeGa7XCbKJ/M3SjBQsWR7vxbuHtorI9EK4AxI2chEYTCP2zw
2Q4D0RftWIf2ELM6hRY7UGW0mzpu+2Mn6IVkqsV4i1PqJoDjsOJ4MyyGQOygAbx6
+MIuWiUK+njj/aHKW9Ag3nMS80jzhvQm1x50q+i8+y/C+zJPeJymcJS9KI12Y+wQ
OBWGO2nMLPF30rawlZ/uZdFqh0Ar/VeL5/HBZQoXE4Y96LRWxFi7fJLRCrWLc32f
jqmbUPJg4vqTCqiQfk9D33pZigSWaFEFyTxGmYs4IlYALfZ+EJcnjY+G7LOMcHfF
ID62CKxB69jq6twqik/iDQHxpK1rTjVwfohkmzqet2aRamyZ3xWdqS6DzZ/2F0je
NHNdInrcILI41kIbgxUiOjb4wlQRXqiG2/OCX+ck5xoDYRRy67aapiC7Sduq8KQH
1nRseraclZlT3euL/fptX0U7guGrFcxHCMe8g+YPEgH1oYEVVcGPMi396ZxQQVzK
o84ds2eg9A7EwhLFMmCirJ99yciEGLZ/gBSKXVJQ5S+kf7DitFYOuhSKFbCwJa0L
TZuRkLgzGsTb4VN6aY5mESWxk7/P5p7Uw5lySRbcnA4aCO0ppAgaGmsZiLsvtZZA
tth/dpgzLShYki6E/O0UPiJlhZO4ciCVSB1+GwrZ9glHvxAOdE/6RqXINwQQGTlf
5yD4Dok2shqA9hYMIm0gna4vycdesGTBX1oMvVfFvNv7/Sg3w3pa37b9g5IzxnT+
A+9HC3uoiFW1jZC7igipHGLUBrqZ5iovdmetVSSTuu7LarohJvnKLrGXonq/mEeC
xWVEGFNpsq2TuJtuH/VStAs+W2SmGg591hKX8RZVHM4c6fer6L3bpSgCwNcV7cTr
tq+q8bU4Mkdkd7fDROFaVK6xCD3JKpff5q6P096WfcwU9Z8NGydLvy+fvhPiHK0T
xaBK9MBRscWgtrA2lHPOgUpQQEwbpfNuNFIdZaehBGthnqYB6yDCOVfC2K3MCiy+
QNhQMu0H7HBwsqsPay2hDPeuw8RZSHAa9niwQ3j8Ma/9IWPtGWLvKt3MVd34Jn1O
tbfv2cVom4walMYXohNxXeYjQCIdzXb8CSVHqjzF29kmEFc+26if/HIw6l8wB5Uy
qOAR+sFeAVH3o1OKUJNzPwS1E10UHk8asetsWl4h/KT04fviQdqvFesVn+hE8YIj
cRwMjhbbo2zib1pCepMf8jeoylAexqMxEAHdQHpaNZ+xh4C5Kx0WtDS5BilprL8R
V0n2GkphSUsGLkaZd6aOTxWTFhUVCbGItLcv1Osz1kUUJPqietq0orBrL4Aoxr+X
7gKElW97681LrLiZoRJCjMJ6KMx6Gu2RTyyq/QxnLK3qhP80C7cYRtKFgEjcHjCU
ei7j0mY6UGNL5m9ehXg5SvLJLX+k8AivYBjYfDDM9ZL16i0RiO0jf5l4p4GqL4tl
4TMWpK6APoT/qm33Y62eiy8FkdtKDswthiiaKDFpguoya9kZrsKbUmFXU0WHRooq
1XTvOvx4iuzGcjbpw/NQMAkMb1UhqRDfLBCHpuB3mXSBRLAGm3Lddw5c/N6DZzLP
vx/k+i1rEBrdugzB5mLD46f7jFsqknBx8jwcg1ddDDlGz0nPPXmIIo1ZMuASIYTC
JDmIuNMSImB3o5EpRHZXg/SRNCgY3AykpCG68foVgGzlPm1BgyvL7c3jL/k+Gnkc
mzPJEGzXvNqJyanmjA4GEFBCJBLgSWdmDWCPdQDDeek9k76h/uyQAn1GEAx5H3Y6
DCMycWqG1NmzISyRUnQK2QVZ4xE4dXb5NYmIV7tP/8QC8Vsn9cFi/p3YRntWMLSa
z5wh5At3hkNNkICG+oM9azPVNaB5piddi7BtoeA0i040bJ2Gp9mrvOsFapumpOcm
254jSUkO16d9yIUMWfSOuJZO/YYyVkkKmhmav8tkST7YtbtK4IftxcKza/EY6nX0
ihRvk+xrjr386jQQ/UcTB4I0MZ1O9gIXcIQUgoeOskTjoZs3g8bU0eFUPi4L62CI
ONJ/yXD/xR1nC03H9WoYOJzgK2Ym8iAsMeouFgNYuc5FNQmkTx9nteGOa3UtOoPR
bMVOtUVs8efyGCT23HfWrfFQAsLfc7ZmP2q5QbbrH0V6qD+Jk/q0pNOEmWkfwVrr
hHF37omngxfFYgmnws6IZjGXOcMmfYr3r8xG/kcz+A49hnTgCry9rl+NNhDboQO+
+a0KYiwbvFgeS76ryPHNT/zC5pF1n5KYyC8Smne9C45xTFTrfm4vo2VXmpIlnNJr
lWSEhEMT/S+LwWnxpIl2MZfVOeEU1F7t+uuiHoJ9Hg5kVKX6nxIRKEzlrEO7838X
zBYRb8d8i2DsWEC28VhZNG4kvlAIPuUI938ds6F/7dc8DIS1HJ9BWuMmtonPxdIq
SV0TgtTKKNpW3YW9jbJDEanBMogvxQM5Zj3MaR8O3o+8Bj+lMUNtjtxUQwl98g4B
VcvYg30Z5Risz3fw0e5N6+kaQ+fDqbnSLYUF9Is5XjFZL2FKnIiFlZiFPi9IQtMJ
urt1c+vshdvjA0GYLuTJ4dIajsUM8sO++KIUYZPYQ++Tze+zHeLKPa2Fk42o0GeK
n8Xge5meiu7jjroNGaOdlShy49Y6CZeJb5/AdGUdLUh/YyVNJ3HI1I5VXxX6Wn9w
ddbmY2BOmNaNLvT3EmrWCNiWEhEJATQtabvekwBMDIBe00mQ56Mx8h51zz0nkXxJ
Fg3WFnTVCI3U3ERr6dD/pVecdFyrI33KeAULPbLUonih2mumWbwstk8ZIa7RFohj
1FmKpuY/iT2n0a1GFPIoa6M69x81mn/VWOmqfFN51T3rRjNkRN903L/Y8IaTNZq9
/ltRTZ5lBo5w0pHSqsphMtodyYsG180aES7y1u4K8qoOYuUglHdoDfUWAAQ2Rvah
9hcri5rW/M0fBshih9YNjL6LeSo8Yl9a+y0DEz86t0PEHLy38WEys+R5Mmbahq94
VgHYZopl7jCuUTabGrgThRRaOU2Yf4g/uEa81ob+QgbKXqkkwpEBdvL6mSXJ7mHU
OaxEYw6z7CVhnH6k6JmppXxu3b6njo1IcY18t0lXX2ljuNZ2n+yxIBLWZKq32YP4
rBUmwNVyHFWKHYxE4LTilm56Lk+wbKJPeVNKCfydG7RFbs7D/kx7/oS8iWocurpQ
VaDy8WkV9kwin3jCbH3jxeojqH/MZPGrsStcNwau93LlwA1qrl+Z7vWIUHZkd6kT
H27he/LZTNNvsVXgQiscF6+kcQnogJh67gAn6Cw6Vwo6nwpSSox5X7MnGSCXfny6
V7KJUBR3TPW0XJEJI9zxgLxf9z3H6Y+n0yi+5H/pVafl4u3riaNNdxUKY8ytdKLf
SXyfh2yzv9lao0DSU6N1YSZ5gsMwjv2CinkhHc1Hh1UrrEwvVGT/48hGjGuf5Us4
OwzQG2lLSS/PkW9JsiWSXdb6AzrTbYl7xuJujwq0XAmy9jjmBDimP0cn0O4HAFgV
pZlSrYMbAG0MhZt/i2DYCaQ/TwkZzEEmR7FZC76hzmFgPezukGc2nN6d7UxAIErU
R4I79Ykg8l+dg9XbmZvWFE0QIoMjJ2tRu0uUWW2x55iHueRSK2gzD1c0Lv6QQDd9
etKwc/I5LBUcNq8FdSd24nXcBjsYzUs+qlif2v8T2E2fcbCjjxl0ZF9PTNok0u0E
/gWVRP4pMLjQG3a3teW9dSisRTFkZ8lmS1/8901cXQR/XL/3/OpbY+6c4JigTdwI
5veFQJrwvmxSFnMDjTFZR50z36BMHZ2ZbZZKEccKIJHtMvoNc8kB9dsXC2+uRPlK
B4PlcZYz83LB3XuQN8h6WED1aNDfflzRUnsisOCPXQfClt5LKMzYLsLUJOe0g/ER
4Yh8SLiq4ejtuVa4MZoHyE6V9Qkx4+jh5tkMCjuuLWyYaR+v6mKG93Iu8hY060eS
2cAG5ZyltXojMCIwj8E/7HLfciorwnLBToJV20F5EtzvuhrrsykJiGhO8w+OylTo
cQ28df/gWgf2jlzpG0ksZ1sZyngfM/fWA+Br42MaK2mAQLeSc4e+QlmJ5IuFwGJs
2kEl0Hh7ajSsXE3EW09MTVl3hCXRknGRj3uaBC5uAhQ7CJ3cJXJSF5rSKYtpskWa
qqRmHQ3V/DcK6U0MfP12ZFGBoxp4cTBci6XoFiMrqNJXpvEUetdiJWFA+jWYYeHt
eQ6jfr2xgVtIU9tWVBxrOPhs1QoiUzu/QVX+FogfBnQWVeIgaNC6uGINbehYBjzk
P9X24SAOO4XQTmCup8TCQQwpRMiWQHwRxZGQBmswX62t8rMUAZVh1tcLt8MWxlrP
iDUOM8DtUpXOCK8yPXCEEzJd/SGWXrmldTBPYoN/f+bO4b1eRXKcnSd6kSWXH+yz
dFqhIjL60xctSfzUKXkZYaFxodxLta8fbsnKCaB/zd8jlt7c8MR7pOtPb5RuYTEJ
LLmBLD+fKLSBMVmhpW/fBoIEFsf7ZT5jh53AaMvnncSP+ld+DAFYUoXfSc4e/mjC
xdtmUlHIN1sxOB51z5TjSZYaLm/xsKHOl/VaNOBTRX56VL6EvbD/icqBn/XcBRGU
hrGfw06RMc3fwrIseAUtcFzsTyIMHO096Cgpx2AoFMX4lpqPW0dCJJX7mrsSKf8B
qyS+36gIqcs9HZTFED4A9L7+ioyKQl27IWUnFghlZ5WP4Gt7MCuAs0I+NB4okPbc
oOE0g7QuxHWBjmpxGkgQ4rheDiKNiZcwmC7EKUoatYPqRsUwrI2jNRMJjMDj7w4q
JSsryXeTrz9RmCHTSphw0ewe0/t9R0XgvtAT7NN56iZYS+7rXG9d+HWaNSqietFz
6p6xvPDaojfAKAGGL2pW+8tUpkZq8MhLNSEUbA9N0rC+sS24NJaIIQwhVpzCBzG7
TXtENmQWjRXqxpFzu0ftYRM4liGxGfsKAQmxbqBsOmUKIky2wRaEv4D1Jb9Bbeyz
rhJQoIlgqh7imIuiQHork2WJUJYbU9NOGJ8Nts0wYcnEEUJF2cj4f1VQqimIgUd7
WMbCk+Cx8eJFRNDAp8XT0P1Vn+52p/wZ0YD7Pu7aNRor2WOizUh28Zz9V7OkfaUx
1puZTxLC+9JIUFA3+Lmwr66tLKBGyjQ+GGET+0vK8aC9g47qskmwGkuriIumelEL
6zZv/V0inzkMbsqEx5tLi+ozfMRg53r8CYRyF5n2PSU7Kr5XEn36kFmCobqunClo
QcGq/cywImWX6g9soaJO7J+hoVbpiMQhmToRSKmwdfdkHzRQ/BZrDOo0vfgX1RoC
JsjR5WDVGYvBhPQR0IsGgSFafPsl0Yus9qNRbWqWb+XrG6mHUaIApthHK6ZlPmi6
77va8eiTS47uKeYFUoaXchj7zlB3XnnnGnevNuKHxTNTJW7oWbEbhzuIzydOhp7F
IdB65pl0vnCXmPYlZVtUFtDK/ZBXZgD1LJw9UiW3taPCij0Q9BHwoD1Pbh+DPtDD
QNiVC0dJ7Ke63oo92jfmVY0yNHKtEE7zhqvJfB/Cu89n1AckozgjtxrOaCj7XemX
i9QJATdMKkD+9VY3sWmMrMqpiyFr9a5TA5WICOq4zkmEEpPeY64gnoLe1CG+DKYV
hBvi+leOpT9QJcur+SZ7l6OKxUFisVqR/QiW2zdXy3kLg+AYBGVZDlBs64piwUIa
evGHfRpNs22nyIEdC0CAf79e+2LtpXPQE9Qdt74m4a8tZlFMKuJwfqnBgkqwifo2
+VqVg14aeUGRUgFur6LKpkm5DZJKGySqz7aQAcZWHfqlJMznlurDGofEPC3ucwJa
gKsMdkmAlfUHq5f7kQlXKgHommLXxLfBwuw75ChJkOLkwYA8GxdDDOUIcL3BRfEy
prXUsfzPexl0QK0s3Q+VvRMOr62tMcnYN1p/aIbvzahttvF1Vvfq1sk75mHUMdcY
k9E8DWUNwFQzx1eIVVVfHoYKfdhsj2K/RiMxGsao8QFU4bZQemP1cREeQ2wAapdK
Vm+8819/Wc/2Fu1FiG58dlRJ/cw3iH8oRehAG8QB0LxPZC7QOEvAxKagWuEQiy+V
XPN5UZXLO3TJS0zLvK8cN2zdw7jyUak17QdTsQtZ/LMo1BC6Z+GgGkyyvKalRrTz
S6LHr3hDwq2QQWINhlf3LpgxRbyowFNwNyE6zrytfm6P68HY/4zzvwJUqBaIXnqk
bIfC6hW/5mFZEZb53KH8U7gosJx8SPtTNLb9kMAnouSAFuSrTTzZxkcPUbfbWkwJ
Xjl3qnmoy+E+8hlWWgriFDUWpJr+H0XcxekvkKUbl8sxkJq9cTJoRMWTZHtnkIa4
dV+uYWigka8YjTcA5Zzk5vJCsmwNd7ZXOepFx84GH/rnY2FvH8RtNFfKs+gDj6RJ
RMwZ2bDUEn3Dua121IuIIkBjbsr/poJKMAGvW+WjCESYmlS5Ewo/GL1o30SNPwMe
joXFfqEsrX4o2xLoER4GYTiSgPMNhbMmboVODWRHyRsU1mDdXLXT/anCIXRieGR4
TgO6j4fHsNkI8QbvHlhXAoOX2J3yTu0+/fObhT8Tjc7MZZ0QHX6w+6aJ0ocJ80ZW
EGsQEdsUhyQmu9cEwiT7unPN13czoKxa3b1ENd8McOf3C4a6ZIk4S7NMQ3jI2165
dlGUubCFKITGKpPNU6qbdntK3uooSDrsmyVEnPWOdddUpAQczaSKTjHysCjY3SsR
6FffsiADdPOUQvZqAfP2Q3Z5MfYsDivaQiTn7uVHi3buXqByH0Iiy7HU9d/Ka+p2
hKB149s6fBG0vdILXOOhWw0w/RRRPw85VBJBHzNyZSvQFnsCVA9A6ZOTfeDl35rs
pUE5jlKsTmGQWpDiK+CVQJyLAy28xwmJ97jvLZiqmL2nlKGeUSut9aeYn1tyuOiA
cCHxvL3kdH9i6qTeYZJGkTTjhqstOs7Yzy3xCLjjxIB3+1CfJbwqShjLVpY0aKtL
gpWrRNsQjmGLmwZNfR3bzaueTVSTGPnpmmBRGIMkDToDWv2Xxq9iBa6YBPVoBykx
PxVMqqJloBAWrFFY6ZjSpzUkr35Bme3A86wPOuzbbH9Yfb3Ttw/v+AicQtbMCfq6
t9iLdIMyr9iWIUqzHdY7NmcwUYhnmahDYfgE8H2cbEgXgq/MacIqxOVEq02IaVa5
GA4So30s+wuO2JAMpIgnL9dbYQF7EqZHWGjCd6O0jAidg7vH7S9gyslLK8VG8Pqj
btGwrgIuSOygeDhLryf7+D0+Ha9V+NSxtNuf3u1N4VATup1xqrLEbmRUFcy90Eaw
FvQjakVIeRTIR/t+O2QqDCxtsRduLXBcT1OfLbXHsPwNDkLYIXx/hBTJnYvxntOu
lRyxgFIEIbghOi0+iD3LG4n7xcfw+AMRBKI7B8EnjbS5Bv0sfQ3SaRjHteywILF/
VZLJbIa0bjVDVA5YflMnUhaKhAgrlNPqNqM/JG0/js0t1Wk37MHu7Lm+o5RFUXlW
kIATLd7VqoQBnxHHw9yFKHS8Ungka+PxISeXTWPlTtb006tcPqxCZWxI65OOIAN2
XEP3ODHq7iMX110xKY2PtNETDNy10+z3uuXKljUT2dX8+rFa4FSBmGbXd3flqnyv
Z8EzagoI9TP9fljoYe8Lo7fLuK3G7s89GKjGUaMpfth9zL33vPG8QGIiK9zijW27
8ZQ4v9NyvZs1tXuiS8BnndTV+XjkBTSWNgQXGemtyo6vhkgux16bGPDUqxqL8v6Q
pnjwafMOA9kMbv7zRWCoU3YTi3bRZSQVfL2j4ptnv4H4zy/0PKSSKDLmaTkxUw0G
a8YDXRoVpcBT9gXjlSxRvC6UQTD1IJCONOGSNBIp+CI9E0Kq8Md3SmSKsmkne3xt
2ailE9c8LS5NW0qtwjNY495NSgr+TTOsYjbnNR3hELTcRYkE7UqxFJnAZHoRByD7
CkbBSWjPMQg0jSqT5zN2lrz668NNtNsVoWPVb9FYx5CzMg0BYt8Nvd4dtUeGXtdC
YRX6j44RzAYoiXOttsgdb1rzcPMED9KN46492XVClcTogq73R/m7PYkpaIKCYFnQ
ClxQZHizh/VYWczgi1q4UqGpiUQcZBUAmyPK0KbJtV4FsKbztyY31bXhZbXChA6V
6U5TUwddq5zaEtDyNglpcrSnx0jFMosPObfWEBRT3UluqFcQFLL09eL5F3EtzYDy
k5XQ4BkORVYMPg6RpO+C/OUOloYV43L2PXMgCE1bMnZ/vMwHBpRqxfYSgvOpdYPM
mIKOkT3b83fmfYLvOAYl4kP1P+cF2ZrvzadFArU1AWboSQD10ojoucf15JdipLOL
bzG3pIQ1fkuRd1JhTpIc2L5h8VIL13lHrU9ODP2+d7kqxf6dCtlAnhzFgnCV+FYE
I1GccA/+8F6p96q4FNSSZgVYosIbzUUU31mWR/jtJg4y0fNZO7PF1moKM7RsDMMp
aoRvT6cLHbXJofgeLRC0EtQ+Wm8WaKkdo0IivU//P+B+bxm3p6fqfO8xg5C7K54y
KaJPTeBsrRhFYYepHLOzYmMv+O/VvTQ+/g/+7zP4KShstf2KxVCdAwPOC4fKPioj
RBirTOKMdt3Wa7JlfTN//A4995Z8AG8cbORkzJkueCW+t7rvMoPdhAnUcjF2+5HM
wTtZL4Xaa21I79/RknvBSYJTlCMxHOFPkXisf7sx3OpuMOCRwL1XuTS31z1Jld0c
15I2p0OyccmKW0yFuIm2+v6C8E4/98oEdEHDG4kGA8IoeXIGluptYod4xZTNdZLG
pv6/3hhmat/QPV2TydgzSXhfkDuiiMFJDgxxiW0s+gAgFvtiU1al+1CGjpXl6Wm3
rgpy10udhWdi9CCIix+35UsLOyY8iygVOS7QlfEMwcW9VmQ+HmyPEpQmZ3MO7dXq
+sk+Fus5rbGdlhoqE+ZpSrkUNixVsKKZmARv6Y5AehBxwx/VJBeftGK/wAwuRnvx
HSUNSAVrN6sbPPry9JKYlfwNTgzOvKXwsv5+e99lQeeuPQABmiSpP7uIEwf4ePO2
dv+CtU40YbKFO/T2CZTx1sFNIJzO7y4bp6iNe6LzJUYY+s5Zmi2dNAfpfXp4IFCR
frUVym/wzq0oJwXWapNfhVR9rLDpSmy+kFGFSV7lZFNnv3ajVi9EGJgvrF6lA1uv
Acfb/AiBFGh2d5n1MW+EkigBc+b2QzRnOr88jNbETv/ueyhpB99hn/7jFHEVKH8e
3kYZvyO7NYFJI7maroZ+bDwO4hmdsS2KHvDHD/aIGFn9Bk8+nQfeWfNQ15CXI05E
dgAD5/Y5xdWjaB7eMrZNLPqiXGeWeG53hn1IN3O6nSG7oBHAtOqZIu4n956xaqFO
51e5q3GlbucwsqXEVZdWONecqQSotlMY1Ppbi67TOC/0pQVxbLhMoHZD3P/F5zKe
PvO1G0r85lQ6CoYpjZ+zCHvOQ5I4ciG/PTPw90RXT0iVrZBB2RbRvICTryp2Z2Mr
bmMjzRcA5BbKayigWi/I8bs7LihkOtez2pKSwWzIMfbVfTrG+HDKK3KjxJgLE4fF
2EgUDliKqC4V55i8RjwYuWBLRH6Owudk05wT6DezXajVAyj471Fj6e5pUsfG78rY
PBzyfpg+RisJiy8GtbaVvNoS5XdEKEYthQl9Mrfam2D8FvXDcn+qNANTcRYePwX8
fzvuS42EU4tDWcTnH5f8AtZhu/s/ahLKjhtIdLYH3ritAy4XUhZFvt2IegrTa83h
BRS4XFKfXopJmtua4U20Jmu07FhYwS5Ny6RAdFlUiV3SqMWpQgz9IrLI4f9VaUt4
J1r48StQiU+Uzkuvv+S8W5TDItONWhzNvoRTQJorRv+3dXVeof11mGyYRZdzi49J
liEIu35jA/7TLS42csoJvTCkfVD/WqLA7clfDkCGUn/P9OHB70ku2H+UKocohJat
avVC16Na/HSeJm1q+OJqzBDjIb/GTJb7G4qr3U08WydumiNU/RkLRdYZEO6eRrhe
50kdxSIy/kc1B1ZRLDqzdXXrI7Ta2y3clDcEGefNhkZEkNZx0SR15cNiydh0u3l9
GS7deX8aNmz/AH1Wn9og+Z/S2o7DGhbmX7A492z4BgbxJIfRcPzVNKRgWlNp/0lU
ydlT4SmuIeSqlVp5/COWVpG5+QMKBIML5ECOQownWPKp/vtRyEpzTw8f9sqM5jwG
yaAqVt/oXDMrt3kZ6nMID43ku64NHGBssQUhBPn57HpYk/iksdmmWADzXUpe5dw4
pKUqXBamcChHzpOghXuCafRgRtadFpmvm6OSZj0aGMv9dymAze/9lkb01te7JNDc
LZpE3k7D6ypOwRHh+X4tDRi+UHExN5HDqBtp32/mQWMTPHz8r/RindaTYNBW5+NI
jDYjMWIvoYz+HyrHnhUNgjxa4yz2VtsUxL9Ps49tZaYkwsUnCVOjk45fitYXvdx8
IetKybOa0IhYfiYTrKPAf3tS8R7D5Dtx91BIkDZul374wkW1H11vmzlX6g7BrMbb
/qClPqy4rnM2kiBGk1ZaDwZfuxIMqmXcTy55GHTMIkshe6aQKfsUeyZbmBV1DyBC
ZPvc8ozXO1rMGUnLq1wkcwdEaeiBsADt5dNs9g6aW7Kaf6Ba7yQTla/hD3ssjZjE
RxreI8VYQB1dSZ/vLvAdICfoVUeYB6EVWCSS7BhhT5kwjIPZ62AtbJiPVvQclaWQ
rSgphrQG1BeFsc/0mfUwlYyxPd2LZhi1bCx31oESTytd9lOKFv6SpQaRrADlakYe
N1Ptwx7p6iShU41tQrGbLSrjQT72oZh1GtYYRd6UyjXIPtCDuB2fd4jYt/rMYYK9
mc9Mw7l8fjW6l2s0ikt+9/WWiKLpReHt+qjw2sHUV6p5tgawS/d+CCDLAhlmpcpS
iO8RGHlRFu28+GkR97Mzkg9tCnwfdh8zpuwyET+i1wr8rL2sPkgLnQP/tri4pe+f
f48GtuJkfqUi5L8eTXTuNnzFFyZMUSikbwrp2CHMatfNN20dUfV4EZ815MtdiYwD
CI1MDBCAdT7UOmlGKu3Hmu+YHyd5cn15H/ioaN1mNCanVUSkxsTaKTvkjIBhCC35
hkCzMZKPcTCtngoc3fu+7MQWdG3kx18YQcCd+50pPaq61SFaSg63zRhu702nxUdW
+wrlBQLuCszfmQX4hBdDQdYkrEjnV3BZUcmHW8geiHd/a35QveIVCTI6iNBLF53P
ikic9j+G1UrmUd5ijSBJ6BCCkVqECQ/zFsXpRZYjgvJMhqVnGKIVVhyhgAKsGd3L
WQW4sNo40A5PXYpJ4ZgH351pMUX5uzN+ggFfm/fIY76sGg1q1O5Fu5ZPj/UhjIKZ
+Gm4YgpHW3sNiJh+bL9c/OfNjD2U6SM6qetYgs8uDYxlu38H028y5PQ90swDxfJu
dn+49IRqU7pROTqAN0X7EqHXoTO9BxtNXGzFUC0T/cFR7N2VuZnDnnL8babatCz+
AvfL102hlCWQh3CVcK4PDIcJBV9QQ1Mkxbjr1J9zjDw6/7OlE+3y7Y98WYMMFnDV
+x8caGntLrRdGx+YukY6HYA/5XXxjovu8IwuMBJCuYrJYPBtvF5SDyFsDoiKK//a
nCFR9uUtozqsSDtCrZQ9gNRO0D0K5+9yVy2CwtGmIvOwIB8VNMgOAKgmb+XyUjNi
Ma8f5ZYWackitgXcVj9fmhsLtKbYuRKo9iijtPTuk+4Pc8xSt8ZV2Em1gn6yKfG0
B6GwNTMo4viPQ7mCn3Qf7xrvOHOlm5QdW16mVkOKKZuhk6/25cBsa5WtnVXi1VWZ
gqk45fVTm8EEjl5REbfdKBMlBLtvHxCMS15sQzPAeXhiR/Lf/txOjTj4RUciHiuj
6KuQe5klIw9p/Gf1Buz2dEAd9evoteC8ZZweacTqMR24IFkfZiY8ZjVIYaJs461+
5wQxtgWobygQouUEjg6pNSQzkYCqEAEnUUNIrmJDVs54vVwiPZYtupuMEwTgwGkx
Q5yLLE31Ii6oVY55EdLhUAtNCvvw1+MfU+XbPVqxW33F2Ofk2aGvDBBKnip4IuGd
4HzuzdFG1NhaiGq5YtxUsO3x/fah4R6hkIT2qOFFozlk+F3GCq30dM3yMIaT4YII
zyRhVqsH/07742Na8aSzrptIIUqE9g5/PCtpN7r2IHE6L5/lkb28sDuCLVYLeyme
eaXAO3SUgugnGoURAnzTsVnzLhLhHF9fskvBprVJY9lVSwIkCuqVD4LfvkpJSfVT
NaYmyPwxlCxASqjWNgw6ivwR4nhVUj5KaY01SVMHJXv19X21m1oVTBjUCeGc8uZN
JqPHsebU2OddRp9XX0mj2l2aVwRsHX7RqzWhBqpvxVM4TAzAfrpw8Gnu8bah8b6e
2i7YgN8lHlm9QYZ2EdnKlfshoA9Kz5n+9Q5DbhMt+TZYN2jHhh4VmXF93W5wHHTI
hbzfLlSNCpx6WVw9vSKdQxuL1vaXwTv3mnIokwxmEb8bHBqBRU08WKiBSFrCojwC
jtW9EjNzJ8DSkH4V5SwNzFwJKc2QMTnwmD4WkQt3sa/IQcRpDxbqfdFxhiqyyqUB
SPyP83aU0IY2jJSlQPu6FwdXZCK+ptJYphHTgpEtyl4O07kLa0/ZpBQdp23oKs1c
Ov6tofVxMgZ8xfj8hCvHTkgUs4c6XGwjaEKbsDhbzqatH/8w+uOlBi40+Uu8QOMl
X+BZgho/WLvICvzQiKU4HA4V6fERlzMW5BmM8jit/Um2JWce6NtQULXujE2QOIml
rDl0pE7GcP7ZhB/tc2kUmEopoMuK8ICTssK+JGyJ7HifT7I7JDIzxoyZ0MdaLuWd
wMcP0PUJ0pbiOFUmCHAq6Voc8uvBfrkiRwaldQzTEprtI7GsA9dkmg0i29ko51ne
NCYiRJ4Kw1XIsyE2Ek8qGkhEvq42vvribv+XH5A7Ux8u0VW+WMFeGJkX4SAY5JZ+
7+jITbDTB3lI2bwOOOhFbtFFJobUbc6hsS8EamEHUhlwt8WQwu0srekn2zSpH8HB
AW6ZHD/1bX1OfenyTjCXYJxU7K4i4BK/157wJHzi8yaEfwQc1NJTOHlLRtLlhMwA
TDwA/NY6BGzyWqsjWoBwxrrNZwX/w/lVrv1+KJIrRIfwP7Vemr9VRI7pqVLfuets
4fjvKNxWhYRmJFnsjIvMrsyfsO4ji7T5kxKQ2G8kz4HyGgy32zV1yooDQgowfVKn
FNnfLmIlAxdWWAR41vkBz17KMVwYwqi3dcTdrbAzxIxtM+n/hsWdVKAVvLJaaf4t
VyXzW/9+OqJD8EWku4t07QF1+CjygxpwkfOjwI4j4rjmpF83IKJUPr+SJNDkZ7/+
+cK359y392m1vHuqC9/5Qb8snSIM57eVPUQnRlV+zeroAKsz+/7S45elcLtJh5rY
TugpzBc0gc9BNXUThvlHa8HtTzQsYaR65owO9U0BqBjhSroI/l6OXbdxr5zyN01f
iT1DEr6Kk0epBeAD9gE6V8PoW9IBgoFjv3daD5gvRczSL2dkYuqOaC5rWBfKmiqP
Stla9yxA8cjNNUwZKlHJogVExjiwgVlxEymGjpv0D1U/nWR+Gxah2nIgfB8wc/gd
LeDATVTUAGkEtahPd3dQIM3/RERA0xWqZcmDxknZHRmiCKhhk0N2Sn+CBKs+DP24
XY4EDdOOwnO55iuQpWYGfHuSQg2w6N11egnl98mbY9I0Da018wdaBgXCr8DQuoIA
3r35XH9C6K9qj3Vbd8x+q5TfeQpn/cBo3Mn9d+rNFkTRznyqeitIzQUQYk+kmxR0
UzqhwfOEix2epHOyA1VTOHyDXiIPEGsqDIj+cXXgxLVB51IUMt9tZJgx+bOO1SmR
CYYuL1CrucYbNZBw7x25xUWRpofzz+j/nKDUOzIxADyzDsw8TpGAj0+RyZPUKwQx
nZh8OHVRa4oWTmkfDpSfJUQSCr+F8Hyku9UFbYxHw+J+5+99v9GQf9GdFQvSdWQv
U41eUCGznXeYBN7zeAGvrBSGZXS+bMV9cu8gPWiwzpLubOOfizzNBQafeBBrAqK9
LtQhF/pTWqC/bxO4mmMawT4gASFhpkwB09T0+YzApASBlsc8viiUbsBda8hZHCem
Hxep6YO+YZwyCl2/6layDfAifOfI2vlfV+Z9hRbZrVuxUs81167XTX4SvFDjXyvM
DoSy9oTI3z0AaM2J63wB9kE4tXfCb38QOhdrQEP0usQGNP02hDA/uqHJ0AJ0NfKs
1RM54/0icYq8R3RWN/GvyIXccn2JHEDJzkxMrjt0m8hLG41jUBAJshJvcX76xT56
TjYpxzb16C2Ded7ATlwNNlCrKxrC0pGi3uqT0JW0P8k1xjDmhhXDDY5SzFrsPbmI
iXQjPNiaVAaczvlIeSeBDVTDCVgJYNKm8Og+0DAHltJGBw6CfQ0ILlBGrUiL2Q/U
CuL+8oa7I+UP4e1R6UJuTHWWJocDDCj/VCV+7u6Us+xaYI4aZpE9qiXA3c7z3g9A
6SIhEI2JtN18YoK83YUl/VcHJAfWGg7fFedj4jjy1TQ+7XHEAWzZifdNvCqwl1hL
jLeZOkx3Jc+SxET/GxMDDvVSf1UJF9nid9FaIvGVDEV0MV+M8lIPFjUIYGRHnIyG
SGtHc172N9JcmBgn4gPiL9xC/2HVeyMc7GMhbPjEy2bkRmQu2OZy1XvKpMcvQlAv
1SbI/hOJ/JNWxT1dtT71Zy7HM8gcoG21YHojrNgH7PU4Z+L0uWhzrUVcXq1rpwF+
p720AGfWTFQyaRikrivx6l7Vs0/TdehMyzuIIgjBUp2dmarLMeX3ICdiHAqOCCTP
cjZfzkZsPi+UdO0TddmsOOBfBtuGP5E2Yd+vIlQ8fYa0AD8ki2UifIaoUXIuG8Gl
TbM87jf9lxRMmLURoaMb6XOz6et2jAty9ELv1tZ9jCeKsM9E+t5ztCOmhDg7Zhkx
TKWBDJutwE2J5UGrGqfIq4eEH2VV/O9lUicAXTOqXvu85+WXJQQXD6ohYy73/Nfe
6E/o0Era6iSuAYQfIaW27dz4asOhO0pT3u+xmN0ZPFJ228VXLBl2my3KFptV9FFd
16M0EEyAXUpy1EH25fYcIVRY9fHUIVfKE7suuy+k80ReKgyHJjC9n9MdiNRK/iRk
r0xs66IjZL8LEOLHJgGcNw5eTJ+jYwBYigmWYRZzL1BgnutfIEZPiCW/JoWuh1lp
oskNoqCPXpqgooaVpiHn2LUGI4RNXo+FoHSRLrx+HpMMiVObc2Dc3xBs4gkchXiK
ZvcVn+BAXhRHWPTzx3kl3Nbd/y9UaJzOmFm9A6hLGjW+2jDh1n4V5j/odrNWnMdl
XUVUF8bShNdtyTXd7/R8DvyyofRoR8dFB3zKwgVtU4kjVXX3auQnV2gNmAK62Osy
JOxmo97Aregft0LAt5AjTFzn5J5Q12T4F+t9f9jxhTkx2qnLVa/6yjxIrjKmMRjN
TnpQZ9hOVKaRdwoHD+VMMG/p+ysdFpogL2NjWE4NZzxFRJK5kxM/lnMOJXxPuH8C
hahFcku5dYf7jnb8RuuexN4mNoV/BFb6PbtDREIldeS4MrXBeQVDSV0ZADR2wRBb
qrRXJW1a4iTW9WonDpz6jd9rH4N4e4ZcKOhZibTw39H8GY5c9xIyqRjOTD/XVq1Q
ivOU2FTIkQbchvplKDtYIQ7mrnobwXvDoyl1yPbCjovXOW2CIMmhtlAIjLk78uQi
Fq+tnoCqpiESSRjRgNrp6aq5uPSA2DGdbkotb8L+u39UrjJ/1/HRRrPSk7yiItzz
1nc71cRssHKPTQCPz6uRa2DrMB375RAC+GCZUhKEXEgPLuBCiFr/kGVYDYYI8Nay
fGwcbmDG0Hb3DEMVeg5wLj6GygCJKB9aWiXFONht8SuijChmksupuEbjElthrxqb
3IrFlPmzexDiIkR3nlRLUmqU+FHC3n/EHiKlrunxHPfXZjoUod3jwHS60EqY9ek/
S3LQv5SjuRIpVsBzdwh7/UEUXqecWGrZGp9RWwYy4x6mw20I//dnER40NJsAXyng
C3bHBGZZFRQzNOqUYF/bsyEchyYhDuqphCeh8n+f+ksq5hp+r6fDEpa+gPGorE9G
zFjpzgxAnQ8iiiCJizoZ8RRTbKcPBqgzoZ3T2utQMYDStq0sf1/jVweCyveqHdVF
ANSUQ8BVI5zTO4dluFAhVdgsgnLkFkoBqmlIoKjx1lSxkCgtsX0ghNWgswbxv0uJ
YVzqtWDZjTTeABw8QOqijlgtAEnJJYUnDaj+gQxWMyVWJJCbHWDmslM2Hx8HCxzf
aWPJRC9gLXGrz6/z/lFg7MpEchCngO9UQOcDf1v/YrLWGb4jyxFIzsaVPg9cCzZg
wxBYSfmClWgpym9jp5SWlaeoqPN57VRv1do0s6JFgSnD7Tljpf4ehInmroELtzOa
lIatJKL+B3RHFWpk9IIAk9EuZRamN3kpjzW9gmfA7d6PAMOWrcZKTw9U6cPpSd7E
axOYMrQHvHTwb2Fcq1/bHs2WUtNszlIrQ7olZXSKjz4SOdkbKs5OvI5DniXv7Yqt
R09HfmpYZUZM3FrfM2EF5MiucghB6ZfVDNfRxQWOSFfghb1QTobNYj1l8n3gVjv7
LI/73ZmS/vxY+WIi3VIVFWfaLeRLQ/6i1Zn5xaCCE8r4UryULfC/BLfmLPVz14q5
eeNpm0v3As+yCbhh0aMUQ9XfQnHrGgE1fM/OTBxlam2vLajksLL9LgSb9HYQWrF/
0HBZUp33tjpiL/ng2RR9tTFVxoz4llpuo6e+1EAVx83/kYmAPBC4VKVNJtSICLId
s3D5GLnLJZOH2HUNoITr0+kP3GKwfSiW0ok2ivaYcMmD4Gy24utuijGlxLwIVn37
naZ+IOLun74uQ2BkMpGwroY/1m/wNUKDHY87cYYeQBq0v055TwnZopZO8GBBGGbn
Y3unvOdxwoUpfB8xuZzBhHuu4iDATe1aGCdcvmv7bX3MdClk96OvykFPU6/+fcmR
uqcyxl/vDN65wHvBpj8tx+y1Ga/UuOUtiwuCkphyPExdZgjDWfQbQ2/jzMWmLLMH
EjXstyLWDpKsIEIk6hKegCTG59dwK8DDPOKzAIjo4tgdf671dMu8ZwncpIWWmZLO
UwbUu/oaZHeTzPqb+oGw6Sn4ND6Z6qLxWp93Vbha1Nhj9lZVVm/eLWp24QOZj7E3
E9KXrkUgK4nq+W5oUKQ+nKdnk7g/XMp176toHqGDPSsNlDF3Ew5QOuKvAUQTPuk3
mNTzrXiE+Nk/t48oELl4KL1V3YzrKZoxOIxveWE52eya9bwQ+7ZxN1FQDzAXqb/y
I5QNix9QAd3CzkRKaddt2+ceLsZLNZHoa3fUT281LKRY84TQnDOyDnXlVdwNNIG8
JZEisddqG8de3vs+S+h35yuKOqNFgIEjxrHuQD/NKSFCfP+5S+dCsZbf3iEsgKMy
8syiVKZBBwMOolo84d2VOubGsivBZiGPFwrSBZBNQ7QTZumnObXmhocXV07vho7N
52z7vS3EvY3ssAFUTiojQ80inASo8UtTOFQe1c5vbL9DAQ2lfuN2hzcWTgv3jglF
92cBxOTXyGJ72shR0Ph5ddiJjMsLarcU3n2ifxQ/snl0sY4l68gmHTQQyArq/eky
r6qay8KAwJAW0B3+jJcXoWYRa/dEeBzcnPg6+uVe4W7iUwNmS7KakSkrMMpVF2go
/3JBPD9zHpPJzUiM0TwlM2wPG3PjSokAkvC3Gu4wHBWnm2Gm8Krzfn+KRxz0XdcH
G664kB1LkqUEa5LQsq7DH0GrzaqF0MHIaIQlVDy9pbTZ6L1BIvWOIAGco+WMxSdi
+k1kd0QMgYxC5I8h3EESAZwIqv+njvxrT4NCGBD1wDNwgxxYurfMzrFmwwk/rFZe
ns5hE86Q9reUz1pYgXfM+O9g5/HDTbkkNaAIr9qWLVcEnpTbnLRMGnfVtXbkp7de
VRCGipZX1ncOIJuBMKf6jmuLaX8DZecexd4btZtfnA4vtx0El0D6gdS5e21Yt1D6
oMrSY0ZFg/BJvdpkfo8vSEs6TYNNtP4g3Aa+xwrTOPMnhCjEWxElk1Z9VG5g6SOM
rqCnNz5eQQj4nivlCpQDCbz11vELh9OfGlGg0fTwGJxTo6PRTVvzisPe6f5ratNY
MC5Ua743r/ctWQ2q+go7TmK6uYeOfEkJ40SVSD/Jjl8r1bwDJcJ7LIOcCFJxCmsn
01Y8x3gsY8Yc79Z810z5EL+KG5XkdTHLPocqnMniYLdpbezqWJpoDYZ8vJuvVgJz
xdQ3+MMM7HNiVtfZgTaRV4PcjlrQTSKZ+JyoB5WMwxmdx0QudBlag56AV+yMvlaJ
bMOkk91juHVIKz9ZLr3C4PrefMy8ppwb1OnUZYW3lvBcL/1uS5F2YYoXYA7mx4p0
r71UW0NsZQ7zM8y7YhjtqSnQJKhcw2KInHEVifJBaBMeaMvXyCqR7kci4DdGgF5H
3lcbkn28A15N3Rjn5FgSzX1eiofH37laFq/2m51lFHS3jCsZSofahsPDAJN2XPSg
o24gao063CwpUCo0p4uRFMGeIAZnrr16RrRvKCiJFu/Q5GlRfvn66Kq5PlcJEUE3
7yL+alyddqIogQxTHqO8sYh8PCNiz0r7YOWOJ8jmNFmEdUnZAeNetuZnrwkBgSiM
8dQ90AfE1YHWgLqMYXPnEbe3/a1xKZHxP5m52QEPD1e3syVChjHsNw2rek8kLo+I
foojqQ/0JzCYn/d4O+JKCQiafRwh7Ip4rFaYcHIawKeZhFa8MQ7NF8G1Jt8rVuKd
xp3WevzadTjmzQht9oaoYy2Rt1JW426uwtFTRKonSn/zJv+DlHtXApgtJGO9E9Zt
BsxxhZJFa5P6lDSfOGfY98A/J71l9mE30Pfl39lYi4t+4vV2WLVuB/Ml8prVzX5Z
StDsj+yPAA4+ei/mXRmi4l5V/ep6vGNJ7hEsDHFhxImCQlQirmZU+vO4XcpsDgxX
jrpb0do9G/3zGu3fBPpVt6iFOVGbtiGu5E8IiXVEKc1/9LeJ/Kzr/irxGBjMBaCx
Ruan+BSsVaW33ihhFzLj8wS/dpvRTom4W4rrffNhAyE7OSfFXh9I8+S/HPdkVVgG
FeC3e30SSclc/F/Ua/y77o7r8uGBlO+hGsuhiPnBiuAIL9jxVw+rxZLB8swtlOYE
8LqjT6Lu7kvEHqerVhDHmNjvaESl88wF8Xa512B6DDSA/IdvvMJY22K4Xamkt4/E
OqkHS54JMka2eg/61sFsQ6Sq68WBx33XSJDyJL8Z9V+U284/ddsswuSSk7XNAFWH
pjOAvIq6ehOBwDg1//a+47qjBlxv0MZHo1mjbporumV4JhqaxavRUt529FAVwJmv
hVWfS5Ga6sv3nJBj6p1uBizkEnnW33F7FtrO/uYCn+Sm7xqsFcaI2kbSgjV7Oius
zMf0g79zMNm42fSudK6c/Yo6aUP6ZF2G5aEeEtn3KQyRE8p+wwve/QGudkAzeTdv
tHmD+xcHtxiti0T7baqtkpfqKZ5hn4B/quEzQlkYp+cRf9slhY+UxETSuWv89yro
dfjOe/+ahkeMu4Gbr6cqAlCtDChUVOTPUp5BM5AZwqEC2SGuTz/hrqwYc2diknHk
Xoi4qfCwdrY+5ZRRY2TXI/tqLT9O+gyMQbHEA1dcrkkut81FQU9Bwiu7htRp/YjQ
jXfZ3RwbDFDs/mBbYvAs9EtDO1tFXEVZeZUcUS8edM6Gv+h5cjMw0v75tqeH5Bki
cPkz8ASAXJI/+Sk+w0uvP6Yc7xKiv5PL9lYy7y4r0JzqO59+68rQ4gF7kDcHRDW1
M3vrbYty5pSiTxoLCXsswzY18ktkcIh94uHNsXKaN9lajQttT6/8Gzn2zTPfYcr0
W/wMVTHP6ATiwpMqSmQl0rO+MTrLczhUecCe8hNT2D5GD6UX179XOcxLu+bxL+3x
lgGzfuFMPsymSsKvrOnYqz0/kjCEMPRb/QsgRpLOI5Cek4Dj58pMg3b0LMLvfzFu
wVJTaUhQAe8cq89/a8rAxY4nEWv8ftItWcFCyV/eJogfPqPy3wDdYfjNMv95YUdO
oWd+/FyWAmpcE9oeilMymIUfraRkLZey4IDzqFnm3vhuduYoExr4qbvH5UFHInjY
CFm87hQDE3kfOUuB6YeV4qAfDvWmW5zArvHJn7+sMC0JUfQ2sJVN6b/+Eig31K06
S4bzZ4DLwni3dROkSFfcCj9WPpx9toWCddJjJcL4CK6pXYrQQ4Gronl4qvdsMXna
HdrmIF5SqnGC/ZZzf3pCVv4xYiT2VOUsMtMnHzqJEuHgbJsDbZcuvGT2yYus3rl1
XiOiBeyE8KsSzUvq7EEOrFdwEZbDNQd1IZ4L7MDkY2k8Kj6YBknEAN/EonCcFDeo
s3YgQEoQkUxlmZdmkVocdXcRqqv4yIx2FB8SO4eDDyJsteKSsuGr6J+0i291cuUA
tSILwMZtxN6icAUEFh3RijH5aB06NcufBsABxDBV0QL27u1JlVRnnQcndtiLBZhO
K1fhsFxt+8tKve/bQHBV/w8Y3mv/8mzvjmCrxNC4ySfZj0rrEyKF+zZ5Mag2ODCX
1qwXUUxi8pnCFmbR2zDnKw5KOFHkiqJ7BMC+KAKZmzzuISljg38lS0sxYFSagpPJ
zxT+AWiNkAmRegDWc2c5LSgS7WKioJf7z+e5Fue+y/gdGsPBEYTYY/meRDIADjf7
POKHyVuhBqTZWAtpkvCDLkse3yK9Vwxxc9VP3FjyG0jUGnjfM0UST0bVLRG1xtBT
ik+NExX6niFLFNKJH05eiU5pxdkeDTbEo5QeiWJdEsBf1BqALaoA8FIF9b+aCyNJ
QjmGwgL1Vf1xDQx+DRXwYhxBIrG3sRssZCHPZoqgpZlDElg9/L+0jp9YlBibgcb8
RsOVztj6ZaKPTsJRCONoMurQIsOpVCn8GVdOYJ+BOOstHi9kObBdFbI7wNK+Dk5j
ZN3VkYcUmc9dMIfZEHgVLDCtJLaTKMps/C6kIZ7Cl3F0WP08TNE7C6PjhvaemmDM
L3t+rMCUwn+QGK3O3A82KcIxa9FlnXJG6laV0Q8v4FVI4N8V4uvi/D5gOoxzgG6/
sszfJ6Ir4s5CO/FThaiPwWx6urDCos/v7vRPOtnsyYI5wvznqPUi1FChoGQivXhw
VKMG2yqR/DvNoWBIbn2W97dYcushEY3S/sZtbVmQl3eMC61faGyZgYGU6Sv9eLJb
1akzoB/CfqOyiqgwTFlZoeKBeiB8B0s3MDSxXhXNwaK6HuI4j2pAuCZQGdaADCwF
YeKObuQOvxtJRa20FSXZWDzw8WrP+N/e0XZ8DxcpEQjh63Fjf5UAlI61jfcH4lPU
dIcmzU5DIGoJATV04LbYylQEklE7Qfb383idCM6V6gEuyxqE6oNF74Ldo4Kfp3wb
4+bq8CC1DnmlZnQ1hw7TXOCJS0CSVW5AbN6gRBYjWeA+IA9csh5gvGeYYoezNafK
h01E9GI3owfUvnnK+bimpvBGR5bU3Hhd70mVwB+xPYBVoP7XNnb5H87npFA+ae2w
F8AYPsoW2JTacnvEV4N5nuuXYTq/J0CDIb0a37EWE1sE6xN1VKUhqpnUc+xHDr9Q
0C+WfeV3vRp/dlaJ6wEU04dfaguoQi9juqPSlRJkyCG8LWaUcGrDeGkxFb+2jA8L
TG4jkqIgpWAAB/H65LAGSt+7koYkfFKL575ssLSk+/Di5k4ncFbRanODCZV+jVjq
kAwik3snZWIL0HjCIH3Ec3/BenQcBf7O0cUlYsfWxhAjx1Uc4g84NhVnqfGhwy+r
DIBfCKgXG9VbTv0uIg01v53fQQU8Qdv4Ekf0tCs7FU+95zg0H5SG9WrkLKjaJuDM
dBb6dvDn5WqoW6Re5mBSldzVyL6vAbsXRb9nQYJ0dauyVf2DskQ5xrkzsyjFziB6
tfONTJ5o1rCGH8DABKNXAQdVz4WkQlFAxEWw2ME+QSiXmDD+cT4EWYhOfkkw0Rwm
WnpePzwsjHPt3QspeupwBk7SzMbaPUoNKTUCIlfLZVdXkmLuqi3+X+939xIR6Rlt
tclL8amOOyJbZvSsS6wUv8lN0+GovbTrFOTJ0peNL47GF64tFzMzDiz6KM4N4q6w
DzUgsJQK7ALtX1FNIvO6t8Lb0Sukovju+HW2r0h0unBtbZioXr4D/D8N+QY0ltw3
TwNO0MuV9OaGpSlHSOP76Xgr/P/xQLp30F33zeewC7e39jAdoOC3PJ1Ux8IXrXk+
hO3TPoUBPKOKk+yBHtZAok2BrHUhJ663UX0/7dvVpjs6bxrOsxj89xfAhREPcCcG
VM2yBIXQJeUvODHpYRbPmo+K3aXE9expr9/rTA5mhbZY2UsRAfih5qB48P2MNilP
tUoIwWS2EBetLZd+ltCIvXp7Feul0xBsQjz34EJQEUITZtTQ3SXuKvbano0hhkgZ
pqzmeGN46ukte49xNdqawq3v7DL/ytwZ9y/aWA9dACN0g9D+4WUSbgf/pUgmyZX6
p5ksiMza31ACpNY7euURKGyBvxhKGl0dBfhGy31h2wLB9uMidquJxRRSmaeR9WUn
hVpTonbFf5nHy8MRTQ+xiFlBPPQA12C7SoUDzh1YCqzbqfdGa3TFzfVHfgbCcny7
1Du/lX143OLi2JWQFmdgWI7FTvWFBBncvZsRhHkkeeJxMLeagk1Sv/Lk/liNvt5V
dKdFohXE/hKPY6EbuGPq5aYOmZpH9JUUFbtjxDDxNIGHxciGPhq57BIeZ4dOfKg8
EgqLc+XhTf9YTm2DcfRtZBNHdpTv1poTMwpzCDXKQ8VkvflGJY6pRbwualVzhAMN
7NXJXT8GVzQ73uhfL34yBW/4umcYlXVBkWnR0M1FyfldLGwA4lHcbTwEHUl3BZBZ
AN5IPLvSRalF55+7B/i8xgExfF15f6YvdJfwQgJlygIG4PIEVtuFaY9dRhNrQ3hK
G60WynruAcyxZgrBB3MBXsdyNzScsVLoe9Q7Lp+KEZFi8keEUgrLjt21NPk6tYS1
29ffOdfKzMNlF69seGpX3bV8jnPxmwyqqB3cBGGcby966+765kUwM1yTdOz0VuXw
xtsUZAZE7PShbA1DOH9LSlSMuJrx8lKJsiddcB1oeQkmogEfRmHXGEQaEgnCDdwN
gdW1/9oyuUfdBvij4o79U6hFk6sIWy/v6u0Hd0/ff0+ZpwA3gc9lU/q0tx9fNAMP
0HRsXVrzO6aIdxDLT1QUE/fTYNeNhm66UwjPHN+HJdj+/w4TO9gOiKXD9t4yD87A
+75ZzXtpzq+VS8ESM8+Btrj/XKf7GlqiFoBKh4hrGYEZ5+pfQLOSw4haSLIPwKm2
cuyd2JBHyLw87/jeeYaolIfs+p1RTIVabzJkS9oPmnIL8CGhRXF4pz2xjNrxuiCY
j2pr0C+8i3/6cp5bfCDfjFj3S1kioiMA7Zh3pGgylKS0uOGIAp07avd6JavDDdA7
teJNXbd6lPWilb+cqoTtEHzFrox+y3L+DY3fMBnkYeJ2wehWkIwddiWvfRTJSIZC
msAv6J5Rut6xchhvNae1rVGw6NfY5+KGrMpMFAwl66r3Yba7h16xySJKs9jwvL85
M5LFIdIVCjID80ke7zyUDRLj7GrfH5U/PEDa13q6SQKLZ9Xeo/O/QOtMgg+18Pma
Q+j8iCtIVENkKxZ7vvh0ZE6bD/2pvrrPFIQhf7vwAz5qPc5VqjXBWktrT/xjVzkL
5JKu/X7CnuGYNAeGtGQCFNLLXjxj/IcJF32Vw+6bcEyzilU9RoI0KeqfaIanUzFN
aKJRWcf3G8QtPr082g19+XGlWKuAOaBpjab3V8CE8KKILbzEYD/hZ15TNvwFpPYF
YXXJy5YGy7R6sfWX0lzNaYn6ygp1fUcV8aaq6LywCRCEpbl5H7L+0I9jch87ge2x
0STO9lEAbbnUgTjZ+cQkXdAMIdOBPmE7js8OPMJYHYBx5TndTziYkmeTVbU486kb
zLh3S1TaAueBiYmkw/VjqY2HU6JKLnnNHiQSLdfGAjhW6ICaSEefTFn0nTjl/sK7
ad36sviRSnLgryLTcB9OhcJtczzI1k7pwb/GpYF6j3H+4azwdmfOLa4veWBe/rs3
kqY1qTHLYv0i49OGg12pWTyvVBvBhjdomglSLqVv1A+LRYcwxbMX4zG1gnPuUBQ8
mBfs4tSYtYaJIrqkU7jklvwEg1t6Q1gI+n4yqXdakcn/KZKT8JGyh4cjVnryyHtp
PuKtmX6fygKXsmZqhDJPEwF++EgU2sqxf1eUoSkG6bixyVgtxJd28c4gjhXbIob8
9ByRVnmNg9ycmpbpnjfKQe/lPlHqC4sFJLDPSq7Vi6gvO5J3ePBT3rUo0Wkl5e8W
/+hfz/QaYIP6/qs/4ue48jFcnpQBr2/8U4e2u9b4NNFGr9H0qo89aDxSCxfYbvh7
TnWN5HMbzF/+yMuJBHRXPTM0VuIGrdLh0Ph/eWkFrOeY6Ue9oYw0zlKw7BRcVhCO
6Mr2lTBkkD74PcZa9FCEhB00aZnH5HWp6daVOVYQ4HjI12GdqoFpfI0Z3U0kzmGQ
Yse43c+U7o1KNF/xM3mSv7rWTQ4pcB4PGPQlNuDDSuVCOX5WjTIwlk9qtzsmR0O4
WUf9TpFq7ee+NWPXv3zL2FNw7Snb603W2DfihX5R/P/J6YNvrAzcgWPtx9VbGcEp
tC208wki2Z2TW8c7H4WHz95uNSzSqzbsZjcwMy6k1CHFRCMwr57zUKlbWoVlt0MD
BrGchfbrDkb8YRKkSkpDCMbiSiqLzLicClszTWZju5uA6b88mFVeh1fgMULdCNEc
KHTn9Ki+GFJdtuIdfkbuGlxaGlAzfhfpT7wnn93LtGdSe9pZ8IlyAXLsguxHW0y2
UpCIFKlskHM4LjfXgVvcwGb5UsGp8gcUxamd5+JP3OnBHVTX6ghkUePQCX2eTGFz
PrBfQIR/kdBeY3+2SKc0ttwMskBXirzpl4+s5c14s8YyHom9rj7spO3UZzi9WapY
GlMu1jh/8B7fa7TOp0gvVczWNsRQDhYb/v5y/RzWF2U6edzFPN36vPG2F3ERAB6M
An/fIDr50kNiIzC78Pawtl9be7MryVwAj8UyMaeh+9bHBZpxtx530FYTZSzPis/J
1VYZ/hAwMMp0YGDBC5iXjqsidanr7l7jkWluO+tG/ikwLfSDroBhYEdZN++ZsSrZ
wjOz/bE4rLTeOTeZtcnkVaiF891i8HnuSSfN/kfdGLzWziBAgn35cK7Tow1qaEqE
HbDlu3BwvT0GQxm1z2ZJAj14q/ZbFGDbfsbQglnrj7/gCH+8oucgUeMkKtRkRcWT
coK8w3mWB6urcmbHiZqRBOkIswDQ/4qhD9nOVrZKXPJwPzZD0qSDZgkWTP4/iCXu
n/BtUrmVkbBrZ/1i8RaR+gvroi2Yc4fbkL1DaBaGq92SOV4PnT54jgX0y6wRsY9B
mRijBLniCnp7LDqB/DEdKmag2o4W8sTvD33nQUQXKBD2ERQo7E8q5y8snStMGj3h
PwignLGJKk86q+7WmXghwl5lyDw8EUEirtC7JKJkJIX9ATL2m4YFRqoMyRrTPYKW
h2DHXtgBFOpv1A7sGelekIz8A1hWhWlS67j0S38QhKHYr5459nb/eMw5b/Dli4Xl
g4rHbr+fvypzdDkPiqJCwJFB9XddthEoyjxD2VljHAQ/AWIafVc63/WKhFtRCavU
s2J3PSnLAzUKMig8gaj2qi2bM7hzcOurcrUBBPeGvOtNKfRU13nSP3jR20w5v4Ev
uSeZfFn3Rq7SQzvm1+CU4AyGC58Y7jEOd9UqFuZKiaU97BrUYEcC5xQzpRhlU0GJ
rDnKuorfQzT+lnjdzFzGv9iHtU0VL4337fyBc+U3A/RQv4WpNupJqf2tteFqpRuI
nb9HXxZu678czAk6pIAwwdcrHujL/utoIFCXGhyc/vg/cNhBhLqIAGA74gjHy0pz
h0nFjTabvelF3NlA0Y3qDeWAGab7jbKjtjkvaRMv8q/b0AOuU5w+EFsklgFDglx4
8CSFHeZLDFGZhfCPTKUEc9uNM/Sc6CnA+gBEc5tyf3fE8f/+PF0svOhvkJN1e4/k
XCAl3AiBDZX9FX7Jn9ZpoyeGgTCYFjOynkyQIRu1keUpUe/1e/qrZpeUqq2u30VA
E5iU9jIP9Yzv8gjSYypM2VTWrPyQ2Ojd/1wb75pzUF+cf3/vo+6p4LA2ZlvrprCs
DYpbQ+ShuaAIMXtTARN5cDqB9TlxmYt3L9KE1Ki/5wmoHze4JQ0Gue8ONkiFFgPr
IM8Tu3JZQWTJ1w7OThhhb75ocDfmnXvwKjAfm5plIDeiCsVe1yuurcuY8XejT8pp
kQBA+2jUEXgS+5Q+NIIsVPVnAIMq3FFRD1/8685DQDuidNMO9DvtRtOUiYo6SIZ3
/wXhm643ndf0n3wXKPWbUI79BBU1NYsfG9JjSb55p/BTtbaThdaioJT1sAbmKa2j
PVjgI/CRVI9uNwPvvQqu9mG0bcNScp6m0vpdJCjmB2RHF8jhWGD64K6O+QKeUy/1
pSyJRARqemQLffOOMi4C72jy77tV9AkBov9I8EKSXM7HSyI7MgEi5jnLitYwVbGN
kp0aY2ds3PZq0K6aoBqiz10ReMjUvW/grPcC8jsIZgyTeFqvP5yfqCgp+EWIdopF
dZ76DdIbwrXwsMIoU/xMwkxcX+iikW9cLWBI0qV5H+KXDkz1C5IrVucRUF13MjkI
s0f/IjGNQoGepS2tR6Fs1eT297e5t1xLZGZ6rJNGyS668XEIfZYWt3UzD1mBFiLu
kFuD2Maq9GWbQyGu7TK4DAzq4/SFxU81rJTFFgn/1Wa+9hMP4Mb5ZR043udT+Bwc
YMpJuA12a032oj6I1CTHA7n8U4flEN6Q981nJ9i/A+srqUDxLCjCJ6GxF3tIEYRl
D4DrJ9Dmk9qRGirjTgZXAdPMY1Zi6h08wQ4ZXvWtccds9GZvuN8BJnGcPup+UdgV
TY2FcdsJpeud4fRUFTjJN9xQ6ZHDIW5SeB0lfDQU5V78RhvzXvrLRrbGN1OMguOz
SDbkCM4bqrjYslmhtxAqQS5fqGzU5HpMYBlibr8abtb7Bo3BswIeNcGvR8eCsyDZ
pJpS8Z+Wkp47gmtMS3deEkjiNzpGJO7Cakg5OJoOEQghEyKSE6DVP/jBZGmK0D+W
/v2+Fk4ZSRLgpIxhYrYTQmzGJZFWZMiQoLdPTgPaY1su1ot0cGtq2y65/L2iwnfU
jsATMMnVochZpn4v6JCfZCJj2eFaLWJioP8wvzkzwOqpzBW1+Y9hTY19xHXNNplW
CRK5ku4kERmQYma0KQvv51S+1PLKx0+1RmiAdx4UPmlLJ149uJnc2dawpzdZXM/5
KVcy5LYthLHunO3BxUnKRbCcWCThw0P0LAFvuX3mA5/CfM0iIBJL30Ub+r67Jebm
+JQ/26U2zs3lw2DFUKzE19MCS7V0N2Mtema3FjKwcfLztiaL/Z4u/I/IMEsePldf
Q3HqsejOG7m0mlcLbhu1hCTY9wLx+ka2O+GEL1PRPpK2EgLVLSIQcT05T6YCgkeT
3dEcbASdUXH5xVnWFWK6k0psP79DUbt76xBAON4RwoWjyzygcxKQEIyXKe1uQaod
ZVWCaxy/U38ltbJvTd6/rG6IfLwXbswBjBP7nIC3tm4hniDG2+NFeN00UbfF6fM4
FGLytIPfMkWSSKba1rWz3+BnYHeBQsK7Yf7hsvvolKBEwfbJw3SxUAriKwwDMuoa
ftQfrtkRPivwjXz6E7b7FTZ9YMs43+1HMhxlPHRrfwczKvUgHjPSfNsYNAXnd+0N
khB6wSUk+uNHYNEZlGHtVQNri8kRz/yZZFkYkIqSy1Mbxh7AAWYr8/MvpGM3gxX2
PF+HmlWBMpkGa5eOjuJjk19VuDyBhBXujwEZgEyVXNad/P7O+jzoiTNP93++hs9p
N26fVyM7ZJme/iOR2vgunR7ISMxAHyHqanEO6y6FAK4jGHwCioVhCFQXsSOhdt9b
EEWQ2fsJ9f5ePhe5LrtFeZuA3hTls7xenGtrnFS8+sHdMLiT76Ga2U70USd+Ep+F
dYXICG3JHkNUngLCFJ6apv9Xwo/lA9C5fnp9cxNXRGwzDEhYKmwRm1oGvmtVcYiQ
w6cWIsSt6UgBtwMnHB3cJvgAsDLblar7UScxnPHW9W8A7B0Bi5PhMEEuNzVfba8w
nWQRj0ddFlIw+PPHhcQc+Yuww1CJvVdrHHKD2hT+aGqtgH3M6lQsK+cczhH87zWg
SU5tQ/Hp4CIeBGTzKNP5GGSbPZXHUthL5eNkOzBdTB6nBErQe7OBaEHatKtz4e5z
r/d6broGvyqYKrhY+9UVuFRAVjPBxfimrlUFailyEBabQqqvu/zntYotjfGhDI9e
zLjvCZ6lpdYcv+qYTt6vEUsfPLerFLOFkAb/i/cYu8rq4vAJnXnCHKRUNOkD61xa
HMFhB5ua7/2T32z4Pofk7s0+vkPhaYOKbP2UMlTyk7PB9PJna2c2EworbtTyz9fm
9BkrYjFmOwNp+RglcNrL/qDdieudSFGZzmQjCNLhJ73GQyUGY18UCBELcCih6Njm
HTtFywi8ZXsZ7bH3PYgvpmjSfN9KS+mVh8dx1/L4Sqj5IE9VE0/NKzBvWlTb/Pkw
fxRs8jgBj/F7i2wscLD4yj9ztlDkF5HXEVMIcynZviBno36pQUq0XPNk2OqWxUV5
UvHNqz/RLRQ5YjS6ZIEzx+eCwQ7bKHXiptpgNcLLAg/c7xKMqaFniynwQBwSl4v0
bNKs31kxZ68ym9/bDavg8CmhTgdyzE+i+d8nUovBg5mQC0sdv2E4TOqTxZ/EaLBH
uBowBs6JdLFupp0PzH8kGGa/l6xXuNsh6uUiV4XpDubCbYEPGzp2buqNr+a84PT/
t2XTeIEpJtyC4qTKpGzH0hWlrDfAtdLabCotSHZYzITgyjon/pNZs1wsdAE+llYz
vkoj7J5PvboLu2EuIOBuIvjl/Ox1zamdHnO8r2E9Qkg07tfL411DYg2P+BWLi6xN
sKFEytnoMmJ3UkGGDWFp7g1vKI8FQVo6sLl6EXujWzWXxxQArM7JSomMqBwFOZlV
PB3mRBgRm6Ln1T3gcqHyzSY6kNAQs5pKP429Ek/NbCz2xMe5xu15x43GI4nysikY
iW6hJOSiHr+WVA0ybE2LJyb19DIk38c6JEeSUwb/ag1S9Wj3nkfUy8sTTVSTA05o
SfbD0IuB+KwLRgrhfW9R9Ifi4UK0eXPNuPXwTDgFwgD7RQZ+NJ7thkOapbzuxK7z
FEwH1oaFD34+Uds7XjIMsv05cZofBwtVwAeoMvLz0k9dnCKSTd4BKhF/+yWWmi6C
vnJ5bERHWBwmbtKIre0uCAZ97PTV/yiPV1mwW1CFUYLmYd8kXnk9xTCTE5rXyYDB
2nUcqBlBIOMnhjq9QUjYOZFQa8LCTi9P3LlPsISaXB8jpuXVKani96WUldfe1Evz
eyeviCPmRdKPK/NITs3wAbAQKbm9USTIcjdXCjjC078oyMwHTZXzhWs6/nAecx1a
s1X0gRKaO2Y2Zqx0U6x/PAp2F86fPXWlILJkZJYHPH1v5MfT1mAa+Zm3ehuocVvZ
FBJnixIc21LCy6Fle67pEDcfciBBrsvQlLnApJgQOGRD7Hc58Ljt947KbZXNn7hJ
bJbG6rzQsl6wI8Ek6LAADcaAWCSSMPOb0na9JqS+/npqV8Whcf7z8i3xmn4oTtN0
HrxPOi9ivHhyQKaoBH74D0xFTg31C9it6mRHR5gH1nmgADhbz7/PFOZkpw888nAW
N0mDfm0L2GLQHGbyqwy4dGhgPusbCyQMKl1Lxf4yOcXwNMvFjrmHPLVqt6ilr4jN
fxH/OVP4MvKdGQ0EZRXujf9r/e3tbxRebKmu9jyacQ3ynK+y9KCAKJlVbFC7Zajx
T0sLh8Nfju2UAHwRA7IRhdcm2G9eBHFqtuNWAzH7SncyygTejwx08sUOtQtWW6MU
lj+I0gO9O99mItIq7gypX7hgJjFa9Q+pXxAo7eyyn2vODmP4tqc5DTlnfKfTHWUB
iTKHpg8Jz0LVH4A7fQClBWojle5eSGWUH2jqncTX6MeOB8rCr9ESXJ2QKANy5ZWf
iTfPO9OBxMJgd45jB2TNZaW5p17nVillKLFESD6Bihe2UqMC60udyzt2j8eRHLkA
vf7IgxiX/u30SL+OExHQB1C0ZPv1F29UF7wWK/Qqbim8Ba4ibZx10UB5BAEnka8z
lUgdQ0obrsnSfI1RWurg9f1/XjBymLROcD+/CZzX3QmJi5yiit72im+YO27CDieB
m8n+1+SaluvwoYfqSLkx1eQByP8fNwTsm+cekEuAVGSsImw4ph+EVMo+6WuWhanU
4l/7YJbEuLH5XUJd6cgibY5Va8PsK/mbP/wNFmCWw9yWPRxc2ay+oZ9PIWvUxuEg
uxI7V1Lri8gR47XZn3kYVQY0+Z3Zk2DMT3ehW64LrUAqR1U8JYEnh9dwr+olz7l4
cgzVVoc06vHlKPC8d1M/Vj2TkUm8KHWPntbqTx2YtUCxLDLxgK9OgizrH/Oybs+U
x174ZFdzWiYxharuA+a8gN/t7s6AwsekqlJxz7CZhGQhX4g27p2o/DsjFcVW1aKh
JgRBxfDeOw1cZ6CupsCuzaDso3KaiRLtg89la6tEZpjNIT2MyydeD7LYxsSZ58DK
zgfRGYYR/lSot8cCK9yOAK/65RVr1DhEu0HzeHFAM7gHGxHQ+oNKedAVeWU6etL+
nZooz5NkE0oyuMcc5U7kbyV4Apg6v/3FC0UGaor75whRtvPXurXCv3iXOzOD6079
SiLSzmwYYkb0wWRQ//jcIBw3aCL2Sm2r9MUMSRNNyWU6B30KtqnEJFZpjOeXPX2T
LnA+Uq8LSKH9zeNfTN5v5kNpTu0BTZIY9hJrRwhUW4pve7sTfSq8s5L/iLfT3rEY
WWuS7D3V1LJpUH4r5034K3JYU+i1U1MZVXwCUmWL3GBkaxJzh0E54otpjl5xOj1F
FO6vM+o/d32SWIg2HkApH6PHtHKsVUDaxE28+jCX9LDK95UfdTthJR/me5JAk9Wm
s+7DuKP0cQwDi2F8K/ForMDcoAqLXMQV+HhVaQ7qFw97l9k0gZVI1RD5Hy/QLoWp
/TX8PQA8x2FIhTPsz9SZ4o1S4CFskwFkgkpJmMBkDyNiIkxy/ogp9GR/qvklLxpb
DG+Ud6pa0mSuG9k1iFeU4i9foORmUAE7RZyydUv+fX7nMs5tTJYdDrTKQ0PxBjke
u1pakaqTom6LuRsd6gskV7v8kv6q+vt+IchPZFSBG8vVfu+f4BPyWIa3v58eTn9i
o/ep5k4poi4mGjQp1SM4Bxpzk9RzPua6OF+hcPPHiT+dEF8wM4xL5/osfrWXGbzD
Pru5LP0IOWdKaxJb1bK6u1P7tUUs6TtjhXrqr273FIbo9zGOLYqcWP3/zWqsV2S6
9Rp/nsHx4r7X5CqrfY/fDqYdtZ3tQqeJPj3kO/xPN5UxQgTJ+S7M9qJsNxUndhE5
jdnGMKiUhA6jTWFRuqyMvyTXVvFvkYcNXO4fvTRG0hserqxNB+NhWaFiHOqGGxmQ
+sQKr4z+bTcBC5pctXARlumpYmoDOKEb+zds5rpI09dmfbk0ohx7LTmfIdGNOb5r
poWihBA4is9RrL8DZHyVTliELZ+r1kI3CLYEI/DxfhYMwt2j0mzVyxiIjtZgAl0c
5vSm8NPIZm42lSUUdflYKj7crtVu8IcYa6BE1pHDx1AH/GAJ5ZMhlh86E+1J/IGg
6LKfNtBCULYy5xTOvl3ZU0jAa5KOaQfx7+P1D214R5eSOMVbG138MPGUW9uc1ZK1
vJkQqa9jwvJa2bHxiGoC3eDUS6qmxYNr0R9WXh61dH1pUIuZbkibI8NWcdRFueNa
+epo/zCVuoApQHi4GO+9sV+o2pu/1/SG7rfGWgj9tuj3KFqRitFOyt0B7VhCKZGA
ko2dpCs1rxQexF8dMN8gIhzA9YSMmkedpwp9XOJm7VZXGIJmYgHUTs6kc7ie0s4E
+8rfryj7/JNng9SleWGF2r4IoV4ehgocAs/ZxijlHU2zt4V2ugSqPidpw50gMoVO
+cGEeBwp0oypReaTjy8O2TUTIOVh2wXx8n3l3pUaW/qM7IFKiEehAvaU5ldc5XxA
iqoYR0exeIiiYsRNYVizXHEQFrIlXOlRVPQly5TiyFZNkMSgu/vNUAUKBjTaM0kg
o3EWvhyQP1YmBCi55rONLzAORq//X4ttM/0TwVUItXJT/qy4n6oUI+6hHAnkehFP
2m3bM+Dmy9O/2rBJriaJjTIENiG6s0xnIFm9NOfANddmICZrI7222km1jn6qNZ9I
rk+tJSS9Sf7nbx9kRA5mL9gy1nFp+8KYq35AB7Ud3Hi50vb1Q5dS3LHCSoMOqLb2
23135A9A3Do2pYVdKYLjp9Ov5hdBayAYWxp88gMXjMazXCT7aLLN56bvlZg2CM0I
qqG6NypA2AJlL9S2z60NxvAZWZEqU6/Xit6sWhxoLM24fMdkXKTNPuZBsY2Rucqs
5f2iYF1N5vOnLnb2TK9JZhX+YQKj2weBhNaXWx0lTGt8W/SD6xO2VbVbeQcZuEPF
64UZD69P88iIPvrWILpYfusFCLu5AiLvXXEFMW+7ETnh06yj7s5R/iGB5RSdvxY/
LFHHBx55WTEdC57VKIXCWF8CGYeh4veYZG+MlF/vQpPVSX4BeGk8KmOX8/07unwb
2x/gtNJdQ/HwqspxgPFtmyeOkWogEUQ/p+2wyIRTinnZjkEw7oGZ+dCCAyxC2ZDh
OZIo+TtPM9r2DskWTXryHswgElXrCjcR09bWj+/qAHac69zEeNkbfMM9i14JJ1oS
m0LLRKG2gdv1tdYY4Q//C61o87OGrQ2qXOkGr0fJ3hei1/d/hOUmvp74FkFdjApW
w1cWFNK8JY0w38oxEjFy2faOlxJHAlx2/EXi5RXOx4RlnY4kfYB4sAyyQtz7oVju
31a8tsL0tWV48skJM36xcptYEhFHiyrC9f5exntPAnZqJIXWuqjFOA4cBOXtWod0
6oTLRxqOGGOzqw5FcpDJzr1uRjV3tU1dmzeXP5QAIWsC4VK540ZSlFj8OINWjuVZ
OgBvv54rrfcyT6wLyS1kvdAnbESoCEbE1lrKxQrDDZFWPO7w29NwkB2A1N0OF+Km
xT+M7hP2l6QAiPTRNy1JAcPDiz26sB7QzMytbdr95gr0AoN+jcLuBdpZ95Oy1NDL
dM2u+qxl5QRBDLfB9MfUzbO8IpF7W1M7kCw5UJUu7hKAMKwyTuRC7IP+6evsohQr
mlK1Z8rDmqy+duT1anzJxRy7IqTKXYhZXktIh5aLzjaQZIZYdMXn1swQzD5RQhQF
2/dzYge6AGwMpJOPLzc0LeCOelvunJ0nrLCwTc1/c9hYEn4Lz6G+ZtIf2ai7W/PR
TFVVVWGiSf8eHsSBAEM7Y9xjTpXmon1pXhgRiBsjTx4ykbdJoE3XxhbNImSPveTz
tz+USP2k8LcnoPaRn/o2D8osvuCfCUjr9r+KQH5ml7UArNazB7d+LHv1o//2CFHl
AuVqqFkdXnZhuM/rIWGJ8pA5roCet5itaWGHav1445mOCg+BIQGFZk3ZHvKMPant
9El5M8nPDO7FFRE2YOIRVmqpWmzmWJWL+ZAQMv4JQlDdYIUkKzNfk/kSdY4K3SRb
w5ipA/6enay9KtYNaq5nP7qM1Jbjcd5pMUAg4YIkvNoPy4PqvmjoNvMk9h0kfg/R
lDPRwwTdPlG57N6ssi/1rnWLBFU5RZjgXZz80s5zduUZnv3FJ6YhOXswqGffgWZj
1lFspwXBYgIaJ9yakeV4NCp7Nj/syPOOoxe4zmdpKSZQxCcfebXaE16es8raAU5v
qghpDkr3eyrOHqChr4xOIqyEXH6xPc5C+/pJ5auoDxo1L3jShVUcnr9pGySR1o/i
e7w8hzjbCJ03OTiFX6e6Dz5GlJecRo81aM7Z4H90Z8zIqFEdcLAgVFjpzHJ0wqnP
Fd4sCla3LjOkN01+24i6WHElgP6pgmYOFEhfS5XBVdBfPqUIXZ1eyn1a2cWOHJVE
BdWd2DeT2Cf2ode0VKt+g5bw4nD4ac0XyQPy686VCQpUhf8j9gRxpxuIcGaojjz0
zlpv0bZGXR5esRQUzR3/4liKA/k7NKXP5XloVzKmX/L3Ys9t7l4kqGkiQzwRZRaW
Fox2MN7JOaGWxyHxztgvGSL3LAhqRaIDwa+BUTk7LDNUfiZ/Ns9Mx7LSYRLkAlPk
Vwmn7XguWX5x/v0jOpvbSpCZPfWgdrRDD1WYH3D9fdYc0Ug85oAwwNpcTNLfJbuN
5e2o/eMvyD6zrehixt6IN9owDc7AEgQrv6zAbs+r8huUQqLdGtPvwB+8vE8/NZGP
qeDcUTbdGsh+oHejTz/YaYBRUD1OyKuXZp1gH23Rf6lSQQ3LVKehWpCDMeZXEayV
x+0aV4E6g0O1Bg66Q/0KI4CdeXFPQE25I0eATtdK5Yb74YFGJ1fXzGetOaxg8Yck
28ecVjrO2fA+6Y7+JCir5MPK2dvku2DG+AQWOkNbkeuFNqfmt6sf/WBwLZmyYBih
3CCjlkJ6AOeNy7UTodOnXoRySkUQxPxqN7biONJaIVIPybWyMRIaXfVMOwQThPFA
aoZxTpS8J6tvbxtKl7Wu8Qw+y/4dWIZfGCn+88aYeyX4Z2ubddB/AkeCmI0B6nRf
lDG3eMQ96DOdDWgvyj/myNUuUy2ZsCe0ofZ/fY44J/NHCZR7a07Abe132zeREkW8
u9P01LzwUVApd+ZDgC6DLxdrVXq1yWu44A6QO7/pQYDRn8oVqEA1k/Ydy1quWdx2
TGSvsxcqqp9FVgROALSynVguLx2/Wih/LfSlSeuHXeOTViKajSbLJzFH+KrsJIQ4
i2CX3ipZj9n/Y1Y2DXKtldkJF3sdk73FmsQgOXmPYN9TqaU9hruen7UK185LZO/J
egEt8BAaUDmrrLG4QdxmpxtFq+yMXrgGTSc3CQBykMZVWO1ApO3TJcZXbGqYRE12
R6Puflogz+odjuww5TujbXIPMJRPZWCe5u5XPckxe/qK+Ykp/BFqSS+/a6rkb6ay
jUWqBAOl4h5yW0vtC4Ppq+X/IHUIm5WGtywWenbqAX6rug/w4j1mWlitVlFiP97W
bU/vq1DFWh3zQhGJ94b2TfsIBeHKmp+NpXpYChnXy0L3x3VEpioCiwi3udpA36bh
hva7x7+hUr4CdX8ESZ4QnCQfzXHTv+Jej1bwuFXOKB3Pl3OIR8KNOGc9sU9jXKrn
6bVcT2LpfuaGD/gkbqtujourxS7Rt6MRPxVFrdvX556rDrQ+Qu7MgfYQfsbITe8z
eB7TLCtf0g4m730He0Y7URtQmBw0FoQojPBb+5Va7fhiLJDEf98SfHt0QQ42k0Hq
/tk8MRbtF2NZIz0qOZVlqJrXd3WNsERWa80l8GB1pp8lfO6cd7oLnlpHhCz7igkV
ZhJdCut2lUsU1y455UbbuAW+5bUzJxXHAqVJswojBfu5XnzVCAZK8X8j9Co3mrwf
asVMOfT7HE8Uv57FhC3KHp0HorWsZ1RXSicA8Bd9B3rZarqAS+UCRmHxRPmewgJO
x6034tMP6aT+cv0vL1CE0D/+40yAqtAUgYiJFMgZiSpd1fr8VS4phzD0rzuG25jt
x0DFdknnkOO/4o/yEquGnS9JV8E/HeAOzw/dE/SRXcbmzvptHQGNxk+hH8xr3+Sw
SJJjvERpNojbD07U1aCilTvhDbF2Byue546Z3a2jztfomsLWfIiT+C5DJrv/CLdD
gzIQrqgOpxfoBcEGsxcvR0U5xJ0dh/WNftAn2cWvTaIiSb0nGvUnNRAuUnxfVz7Q
SjHN4dEadNojkwSWD4JUfKzLyh+Y2xSF4KPJIQOJOv4pqYahO0COXFue5SSCJh73
4sFsozZANQh9b4Nx7xFwvhqjVEbVOqgin/BeGFVs2/9fivfesWPaHtMEEqiFl0jd
G5K8tksFw0E4X75xpmgbt/wm3SifUJy4pZXu1+JkTbQPY/1VC+hc7XIqxeBYdYYg
AGGCq4FpGzRVCHoFJuy5+Otj6mhLavNr4qtVjrEE3U3/OsW4QPWJdumBP/yO2CdA
UVLLDro3IXpIxnRwk0uZNvjy9P9d9gxVaTHoJzfsQ2as8ZbDoFC91LCgQpVV3Vnz
H9Ij/BkolpjeJEJolJqIszF42E4W5cI0SeJ827nFYE5W8hVa+pbMGMWd87xPZbrW
Px6b/TrxEgyJKi7CnNXv8rp4qstlSsNxRNeCA30nVYsv+QSHTWkiwA0jJTcszAaB
y4Vo/HCjOPJqc89NKQFmk/6z6hGbkdsp5de6b80+o1xkqCPpcvP0v5aRX4VoDNyr
9YNrpRxP7A4pcOZZNp8sMzcddW1XUO8XSgfzibCenNtzGb+Tj3tEKik5b3KecMxI
Vr2cQS2rsd7spKRo3+rmj394dOG0nWmm0Q0Tj5gswfZvVKO+OmhVTgKfVday1HqP
/UTot1eoNUKYnwPWghMFR1kjuoj6TJX2L8/NqGcvD4Krc6huNpIAn8tat5v99ctd
Kbrw8mVYvwUr6EQQGGbERfK6Gbl5MawBSHczFFy5WB5omgDZ3qE3R4m3ETIJS+/f
I02/McXkW19UwpLcHoM8LipNshcslPGQXm1op0IY+c/bJJSG7CjHFAV5toLbmtvY
2mjrX8+XT3Yi+jSC2ICEQmPO92cy4hp2MizyEY0lX9yGzSF0BlQXQ+P4/kipiyBW
uGcqrxusU+HRitlDB9VF40c2Dsa0xVaDsuAGUTqtEzbXicpHV9Mr66cmHuVV8EOr
awObmSD9CCjX5clYmfvshJnojUMDi5i5nO7oXRUtp/Svgy8ypq6ERa04QL+gIMX1
osuDyC1ULWuyKN9W7nngaCvM5e0DTrpLIrgLZnPkcnrflB1rEvCzy8dwCGny0m0p
OG8091+0whr8G/c30+c6h0JU9li+DSjtUEpzxPQed9RGT2oYdErfA0EjiIatQZem
ye7R/4DFVf9OlCX//eYcZ4Dlu1cN6NTbZynI1SEIDgDN2q48c8jTdkSVKEfC8nZr
B4uV9rJKN/D+3xhHmKc6A7kVhwEZGmSYgYIptqfg8O38Sb9oaqPMGO+PmTrE+VAC
iOF8kCe1TNbRclV087KxLxWVdMyRzXdjoa+Rb1pCOWPA70ueRCGOWJwA9Uv9iWJU
Kb1BJlm3oItU3tMMuaex8rFRApTsG8fB+LSDAb1dcz6ssWhjLomT7cwEVfp5p0zJ
BEwoCJuAntlc2uXv6xUow5i62Fh6S+170SoNfsEpKsZYT7DODcFYX8z4XB/a+wOv
HxhSsrj5r93rQLNJH4cQw9MtIfa22/9eS2R7h4z77oeQidBURzCuyPo4ggzcDvKl
km3tw61u1iPMVsB/gzDp+bce2JMH9HQJxw3rRsIjeC6Ab+pajo3Yq6qbj1XvsgA0
6MuWo34FX6r6QjKSsDumXODSPAGhg8YG2J5QirYDA29TMJavGSYjqr3O1aBiMcFB
OnOZZsmlTG90c26XPVQ2+NHYc/uFYk9b+8+2Nr5s1kmME6/S+K4LaibogOYfueyg
XI4WTyGXarKt84A69Z4DrhAhCjaabVdq6Cv//ukEsd13BZzA791vDKdne7OCrdQI
GAj7/ZYOzHB67OX1aeCCrGhQXUZ0w4GxGX+OjPp34xdQuQGqud5BYekaVCdp0fAS
CDlMJiVleHBLCuSMGHM055NBfMrXSmCX7sEBWD/zuBQLL4jmu5+5w1mAW6/MpxO8
Eg7rojvZMXnLRGWpQss2Iz3tAAq/1S1CzyS/3EPAggn1hCQYD7KkTDP/IqNb4xh/
ud6ACe0xUY0B616JQwtQlZUNROmLWZoxN7IkObbZshJcYNk1Z5mGq1icrcIlwRt9
0vznOAPsE14gJeFFfG48PEeGPG2WFXGMzIBgTciyK9y+8jRmWZuTtdiR+S/Neweq
KxZucTxRUi2UlxixIrnvhJs31C8rP5ryj96sjsHnUxSzz1ePZtF78d5u32sSYJDx
HHyFcwuNBI68m6oxn0aQhFiMk713Wc0Q8zUk7SX9n6vu2BIKA7TzfoBaQbSuxWM5
Y9s1irdevuT+rCSUN1aZ/Xjs8avDJPKq5iWZ26wuhc41kCD4PAkza/U4p53/dZ56
aG6IymZivd+pTfFh2NfYvDE/yKVmibhPf2bR3zT6nDdXDymDqZm0SeQAeWoJ0GxX
UGnjx2OQvDyGZYKCpL4fxxcks8uGu3QSE/T/5AY9lCm55uXQoBtJKu/CbCWBdeR2
7re53Ah8pXnC8RMJ5B/xRloXtT3tBrDeGdZPFV0dU2gPG2WBA3W2sjIivQ65/oiH
J9RNIFFY+Xn9B1Tegj9uV6hB9KuYihVeOo0x+7MuSh+KlP1fvsaGY921hkQLykBM
zqSGqPVAu2hsYb3/VHa32DJoZxloE2d18k6ddaibrxjh5QXWhCuArxVlv7T6LBqu
cZt4VxtoLvM9UE2t4nGxiIEyBUIja1+yz4v0tg6bH8u42f/DdaKqSloTCeuXJs+b
VLOQe2+Pg9v2TJPuhkglEeH4TJbgj0EM/ARNh8ByTbHUratTw+hqm3PXCjCdDJ2A
MbI40UH55v9SVuNURti6mUY51q3ViFsvA+3PYvV+DAqouQ9MV0FPPUvHm/WToSu7
cFDRsOBqdgYVebhRHA8f7SB7u60+JXDhrc6/Y57ax95GRYbTZgd4smUlvfzTo5JE
DyATsL4RMrGuTOU41ZszqjVu5sbO9Bnl6HL65sbMhAK2W3FN1LNEC49slVwo0YLH
hjluMVCFEngKnkjKE1M0pocZUJjU4ok3zZ8GlXukL8ipCuj7FPk2H1fYe3HS3LM9
JVhd89aa8UQUfyEKMKfKAFKSDssaZQUx0ebgkEpm6ailmpUEy9XsY22w/dgefgMd
SmzGkKARthMoHYJulIRmhbtGShd6799cKopx4VX1EaJKeVzHNuEdFFrPxTp6GzLI
JINQercelUI3hTtUUifz72qmFHC/1tq2VX7AsxjtoBM5Lx0eqFhu5P0bReP1z7Jf
lZjds+mT6AC6PFoM71sL9VRDEuf7FE+BPRLNNgtFuNcDXwGuUQ6M/m24ySTCWHEV
hfsFDlU2iEKt0Y7A6kaaG5BS2p6ee44YrOAbPmdcxhaeivQPMQEs8HH0D99vNOFy
j2S9LEiLE0agoiqCN5MfSgbxVnkM5+XkgvodCEZslJNFLZPgmu6bQGpk1FA86bL8
hDOwwNRIHB4yKAt1NkzJ6Q7gEnhAJidyZGvhpsWrjM3NsKOgTfY4zk3DVemqI0rc
UPPVS1qK1OUIRK6+1ytvCuue+1c9vQp8BJ3kO0K3/ue+B1XOXviYZvL4rawaIDOT
RvJIvUeVrC7XBCPrN4DHwb/fKVq35UojA8Z4sCWgv+/kTIGFvth0wR+VxseSqyqa
gONKGeV84MKLj63HMEqROkSJdpb75z6/8YGzgGsc0eFUmii52KQb/wqJ0Oa1gB+8
LD17299w2IUArxqcvHqc/yUMTXFRdYA26pRVoSHAKrYI/nUpXHfJ/Y7PlMT4wVtu
R3qWOON3uZBruG7OYkybAVHhxFpBmwtI/sOjq0uZ7CLrJVVyqvS/L+nnM9AI96x1
dkxVe8qOr1qA9HCFsSCLt9dhH1gCPwzG2W+Zr+C5SYKGfOZaM2BqGVIGTTihzZP4
t3uhqVPt7JpK0CphrDZyJpqBU9bhAv6uV+c5TBsJXBsfdiv/lmMGt/YgO0cOFOSZ
iUFYy7Q4+U6cXEE/51CJLA6SQgABg2KgMbaDC4d07XptNzCZQmtrlzHBe/eJ42ZW
sw6xHic/Q9fU103lNNPJlMHuH5I6ER7BXgZ/CJGJQjZo6zUzR2d9eauDCxUB09P5
QIQAdTvWNqlr84mDoQZmonADczTQbG7cQFH5ABhyebbWP2NAupQQa6HavLx5JUHJ
IF1Wrp3dlZ1cWUvCx1L7/8JhFUO9zjLfcVt3zxTVfSvv6Q0A60SVepRXTy1rj9YE
EYWvKQuHoJme9xVVaVKOuBLjjcteiv6np6ZfQMwTJChBCSuDp7tyItg5aiNpztpi
/c5hAv+LNyoBIGml5WNESIT+McAN9jnn90HKBB2NifIlJpqEKXmstDGTIxfkk7W/
aJGm3G5qDAvdii09lcBrRMkbNUr7m4MWKlDm/ak44JXg73OZitVpiRXABVC76Ckq
Y9W34SKaTGol8PLKbQjlzW7yNaIJ6t87gAqB/a1ur4isEqnoYuE9E5jAD+RFDyTE
mk6kuq37UPAs/coNUFI7AGai0GcM18SbMmUch5fBgLNySAnpEmPdZGzBTckNQ8Ns
HkNLxZc9ivR5kFwtlVwocIlSSxu3NnXWcjarwLhVc7Jb6uuhF/NgP506cwVnF9j0
vsc76jroJiW2IJkIOo7zBIQGflkyxoMtyYwH0TffNZC0g1An14E07vbQSuE+IxSs
slegkx3YJE20OLCxqXdSkRu9eqzmqGtjnDyWUhKe6u87zjb0Gu1NafDfOJySxMBu
ZqMPctHOCUVhVA14DgGPxaD9VUMdC43hbe2VGwmtB9MnTrJ7aOlKH/nD1q1hOnYR
kRY0tV+J1fbvtX6eZde1q/EFVd5Cno8MAxoiVS7wkFKGAh4KyAMhpbWaTn+DjUT4
MIg6GFURz/RzBz4RibJ7BE6K51pPSf+haCHEuub+fTn8mcb79V5E4plrOrYLCTkF
tj1kstGzvnm96jkt2bQhnS5Jfpjx6mz0uS2b38zSiscO5qEZziFuFUrGKgNTwFn3
2VrxI8LEqohkh3Kdhh+hU2X+KEthytrc6+E/nkQl7vSmeIppktVzckGYfg+Bh98g
FqG2IajfAlys0hNklvpYHQCAGZXuZtMiZ5tQGBAuXySF4U1y4tIHqYokSjDchAlr
rtCgboIF11OO9hqh0ysazzIEhgHSO/Ikmi9hihbCOXk3L90ioevtlGzqQsztDawZ
9kjYPfWneu6Qq0rTi7HHYNGYgP5cqSJVKT77pDtmxY2ik3RSpcsq13wGnCrEqmFi
eUMluz7J14ZRfs5VK7tM/6TogWruZl+h8re3LvV/dgh1bI4tf2GW+oEUuxK72Geb
vdQXYcPDcHofjy2EKT6OQ+Rr98kvlgNBmOv/2Pi0J7SpfK6B8xYHilCaEu2nOxQU
IqRrVmFoQMIS754yqab7vl71iEmlorLj7ZFwgaSkTpl7Xqzf6HspXdHfA8ts6laL
UW175yBG+sy/4Hjox+69HvRBamJk+FQ8SuQTfuYecelNW7w39KDHdb0V2fipWEjo
wsLk3/XTPifINmx0bdNPVcAPWALUu5K/QEp2TkhV/DjL0EWXo2XnqxIWAgt1ggKQ
z0bQ2p9w676Wn58GtJ+9bSyava2WsQTC6k5Ngbw/vAyTCSwVqEiUFuFCich5rEdp
pZ9LLkQcT6pAhaCVDui3hRkrF78arddphUvy27KMiD5VuAEMmEkF0xzyR7qI1kBE
lPKgaRzhKdy/R6cRIu5vFHU8UCeoXUTBe6JIYEFdMCs3t+9PtqOkVN9/J4VNQ1i1
2XiOP5EUz2cDHWZ5yqaRWbAkeprRrYlfGvuV3SfSGr7oGvSPIxz/26TQqjSEcCf7
J7FoG1z9iCcYoDMBS3IIFLuZ5sLSAHo47onvQr4sLs0lR/m4suzc6pmc6WmTvSko
gmAKZz4kRyobgp4HQjtdeLKbGbKkiX6V//YjZhWaamkSImbc8qxV5Lr45fU/fyPa
CDIUsJ3NkGcnJf96dETgsJG8EYoIAV2fYeAfMZ/TYpB2vXF4ZfERhUZ4mpLbG6eB
Pr/nbl7lgOk6hCzn2NXK9yafIdP5Q/I1gdVTUFnakJhDEZiSw5djSjLO4l+EitNL
TraeTX/Fg4abjda62H8mnKmT5/KzKSeFxJuTmOlunXgKTtYnQtRZudfItWQEYCyg
kxagx6vML6Rg53YmvAc0NaJ/+ElhwbjM0oYX+2ABRYPjofs4GjOXkOZBYLDRHFWt
HU4EFBPUNK6s01koEJ1K6U8brArQTmJmzqpTTA7Qp/3ROhlRDxlpjHEkkzbGl+6Z
ACuFxbSSivoWaQP3xaqgyQa5Su2ztjYMvlJvhSTYV9mUHC+Y/Y1gmkg9iHC1bAxZ
mQ7FTXmGfF1Cp0TWVGEBtCq196H9zbmUHeXP0QxgLjKAGxAcmN806/PgEZgkcT47
3AJR2FbkzFkcN33jZR0VLx3TSZUWmofeyq9c0pGE9rsV5nZ+5ei6tIHanwmylosh
cSlSIo1MV+vh3A2cx2xL4YzjbWnQH/04+uPtixGCkN8hvJMxb+X7xbOBsSblCFzT
sxXel7ohdIQyLxQrNlFqQBZ8ce8nFOWHU7DQ2TKeV/S6aUV30EcbJ1aLavq8oklv
8UxXJlZkhowkRnE8VtgkJLwxsn62oMXtD8ccKyDa6wwwNDram2XT3iOvy51j03LS
VE8Zwv6Wonh+w03TU0idhSsjVU3JeXXgIZBKNi+YDbY92tUlt32nXhduaQMLQC22
dm6CWrnvuurBEdEhXaBLeJN+De8vAHa6HGuMWM6TCxiiBWYnT3HEaMVw0gux1mW7
7vokbyzq1k3sd0xApkvit3c5UicLAQV2PwIhxWTg8oPHrD8pfcT1jl2cLdy2tFcs
O1C3Mj4HRYDcCBkjrXAIubK4chpSxoG+nJfqaoOJ55chk7nI2Riz9p9xi9m1Dw7H
LCv0GnAiec5MZc+u9pmqYNkYfM4NquW9v+7RtUjh0+pF2pE/dzKkUNpjYBDomLJp
zk9/vWpB3/R4M4tJn70oh51PUI/B6VjM3JJbrztufhdplf3vPOkKUdFzys03MKat
SEcnrJ1MbDSXanP1zaD8PmMXOxFPpvbxFOuINknuzxfrjREr9qsn4683l80YMMX0
bEoI9fjz99i9MaLwD8MkQS0nTLz8kFCFRCatiNf7GXHIa1rdymh6E2QGF8qCWXxy
Wrpei7JiOssXUrO8GEXpNk76eULKehVz87C8G+BmpbI1lEAqxDO2f/Avjj+v7Bw5
3srjAHqCFGcbgMPLYCnBVoRv5aACShcVEIbpVG1bwuqyRc/vnmsLFjR9yRo4QkKC
kj0bGGLUd2bewS8yWLcT2/jdRmHr7VvodmzL+MYrLgryVlltcV45APjLgF04AOVb
Kl6qqvhEvHHb4CXrYrPbnNnNfvFHoxrQkhtUvL4tFqBzp7PbVIYiZijOrgWGIGko
2GuTRuPKmuPkprt9YJWcnX76Hwy3lZby9yo6Ln4nOZ4q5+ZPc8ml1OA0Bt7Cdwtc
yS1pGTRAHsR7/dQquc8esR4xLI+dmRpBfNrXdl57s1m5AcLCHtWrOiFP7k7hBrwb
M6LSJ9pyST8q/VzIP2IDLPpwa+oiqm1qveCL5paH/4Z3+tUVcnGdk5/WzbarqU3h
AwBWwXQazhI5VFf5dcskifxbfpILcbZ+Vc2ZOvYzFh2aRsZAdZgmN9LW/7rh4Y6u
Pwk3f3sJZnxM4XTGUSyJPW+Vstw3VvkrGsWNBdQHd//ncZPLijdSmjL+Oz5QQeRz
v0XSGOP8zP6WLFgTw3E1LLJAk21mu/yuEf4i+zOXrqb0fZBlZTqKzzW0YCxfsMsW
1PaEgzSeGE2jEIb83REtJJN0MnXurm2b6xYxoTMd10afvsrxt4jRVHuPYA/pfQGa
9sGz/bgZBSATxqATkVnO9p54bnWrgQkfYJj28E9MYe64LD5kWC25th/gbiN/hsIC
XlK02zkDZWoATSUftVG78yRqNrkiRqWe4OEwKotqAq7og4Jq9fYQ9ItqLbT5GzS4
+QRzN32EuVPdJtLz98kU/4KAKapqqOo4/qpbRHFmQJS67l3KyAGSzzvOBbTqee5N
bhBJA4jqO1F3Sg8FtazoS8wblh5QEbxssuig0j8WrSua22476ocL9ARJleNAyY8O
IFY6NHZAaTRe2V8ZwQkRXkEdj8QVE/tvtCX7n4TGQbofaddqIPhX9+iAQWZ2CROM
xanIc6txR7txZP35Q13JApMuVcPKUipOCGOM+RtuhdhinNDtaDYT8wj6pxtUU08h
Yr6DFo5LSOFRYDms/m7zA0JR70Gth9dsVGeqNJqwv7/nNGz1jpWqGzLxnadN9PMB
4up5RsQJjCGoEWCaZnk3SaHHXCtjQHvQUg9kvOu1UKrapq+yvZeD/b9cNSAcHk6i
Q5BsX8HETcweJfZuxR9VXO9rQea5z9VUWg/Z1sUiXMGEnYClSSihdJK5u+CQOEvG
pymANSkg8pwKB3kcMvFhj30ubKEX+j6o8T58CvLaN66uR404gFs34yxvVdy5UzTV
gYIEQVY6CNiWzrckiJzVmNy4hPqUnLi833mQLvx0T+O1eS4JF+2u/2/4vCqXqlOP
omzIlEwePClzQQeopgsXvXqZmlzyYXN6dnCktrwmV/P240FD75KS/IsWKGgM8X0n
vGsR/bcF7Afa9DunxYI+/krbojjy+PDY7BkFisEfQ8HPqxfWGTDD+ro0svEzok4i
Hd/aEAD8fk/z4d1OAh6Hl75DdawjPZXGwgpICGuvkr4ls66TspeGUYpv4C/+4Sm9
EUdjiIImMurRuIMmuqIjRYphwXcnldTzuGKYEHNVfU+1oD1hRcgpqCf7XJLWoiTf
dmNVCL2i4x+5NY3yFowkgqnTApaY9rSzQ38TLMmfc1pL+hVHHAe41n8e/17zahd5
48J8T/Zy/kJCboE1zf3GGMYVVpC3lDKIydypOUrDTGlmTpUJKQ/pe60x9cUJ3zI7
lzyk71LnxJaMM6VTqmulGJfKMwZYR/2QmSa4mvNSUCsaIjYVd0YT1xD3v62CkYKv
lUEx+wkQ40SOxsluXhcH47eSodfao0qw/N6HEgQqW9gWmqvnCl+SNvwq/N9brf0j
eIHPWCVn3DkyzjDJEuz2Isbi7swovURYKEB3rhi5575iLNv8o5Ng1DSdUy4o8lZ+
i9aLEVmoOR52DhnPRIF6UZdFS5KSs3Hm8XUJskzb8RC54KyCUZ0ql1ngpM96QzpR
bcGxnEc+oSMFMTae2soeCBuiUiLoTLLXDUCYVcBk468UIhQ1A6C94l5H0lqcncdV
m9yL6f+Bagy2hnAn+yGpBKANHMqbVv/Ytr17OvCG+2IgD5oijLT47cp9XbeZt/ig
ZXoFhm2hbKVzSKQwg7E1k7oQi6ECYRH2PmgAKrcNMCzkyTAY/FkYh6m4DPCLBdJM
ZukFLMONL8jySK/sRyyG7wufzzN8jW2GMuJ9H6vwrF3BP14PbJl0SchcOj+QMo8m
je8nqW0hhPnFRMBEs6rAyfeJC4s9tCc0j1wrcveXUUmoYw8VTWppc0cWcwpmo+U6
sEyz8ulvgEQe4RiHOTt2hdvsY+kds4HbFGOCseVQIXTfZHZXBygnloGO/43gsA/j
befT4nCID0/z0ag1MLoaO0ao7A7Xl/otJVpbgjyKynjCVDck2BTimZdPkyrynAkL
tPr95Iqc3XXqZwYmw7NP4T363EjiWNT9sO1NWQb4cuTeFnQuf7/VtvIqdstq6e+y
aojIj3sJoQt5g20f8PTO6WNxP+KZKkRRaI5XR84KVZKSll0SmPT8hOif1SzWtPJb
SOqD0nO/1Bn5Kw0KNmm/hwwn17T99SjjnvXlfqFlVd/XD9H3AAM9zwC1qwFFfTua
qMqyNJzH1EdJhkjNfoAw1u07ZlU4ewgjAZqGgSoVImNzv6B/tGVNtZ26b3GhRphG
YI9aVoz/4vQv3lkOE8UwxqnTlVa9swNiHomRwtEi1vzkwscJiQmtHPpzyxRoOXeM
0w7xWrvTu0pdMYrPbOq/1tfUiHuyfiuSU/ZJNsYfEjDyHt8VGUWDc1wS6hvkHH3f
svwnEYDsM8UeHCFVwh3Z52lg0I5o1PSADEqoQcoJ9wc6BGQ6SXuP0R38O69NXCa/
DM/DB+y6UFRBq9O50GP2vHpoDFa4NEP4QQ+u77L4VTqko3J77UC9b6kRIfA8wcFW
JXclmfPVZoVGiD7M5kqyofFQLLHfwP9erZjJMQ7Ve0MrjVWhkvWpDO5h1hNVz3ds
hZhH0cRkOBnaip7hVahaeObqaSte5fhZ6M11xj3TyVxFShDR5UAh7hSoqhzw+nw7
1Xpu/D2GmqCZqED3ayb8STZKy5+d0hvlOD/6Nx1Q9CRXYgLIOYBPb5/Rz197kvwK
dTV8546ywzdkPsUlKM06iHiLSlHCc4tAcxTzWOEJd3oNpx5tZD9oc2WKpi8QhkfS
FH3BSmoZP8W+2FrAPZhW8V1X82TMIvaIXKSpRydkrPgUC4fTSLW9OepTu9Rz6ngh
FLwZ6Oz3B9H5HWPY4GQ1rppXhuLNxywGTwYYycUuWIsd24lLBRgkL60gjSBSzkG+
XNongpG2tkRgs3+Zl8Dy8nNd5C8G7oElUkDV+OWWkbCpxqW3sPEH0lc3ee9qQLE1
M/PA/PLgRX3l+fFUL9sOT4tvtKLQBbYyItgzdwpKTkC+oTlTuE7vZCtWCRAI4K76
coAYTrfDM3FSewY9fj/egnDS0MWSE5YgudLOXOWPzIf9eao/AsqmrMh+EcwaASB6
UegABhTpDL3pLMCW3gAObh6kAHAZDPEf6gwBIYO58uYo9IUnmbuKcL/XdTlEsK8e
Kfzx/81kiY5dGKUL2GCD3W+TOGyLKFkcV3GcrPw3U0smd/SU+ZcWEcMTdOt/8311
srbYlpEp1HJeUxA3gmDTLYrTAUo3lWEoL4PCjpbKKBmCB0c7x9IPSO57cX4E33Vi
CUu/MRLdK17cIreC3fpccTf/0sJquqr7mHgPtqxlWw4fcN0nDvb9Q/GZw9vCsFss
vSHeh1U3in8eW7vlJNaXm6PrwWnd1ZF+lck3RpxuAbzq652rOYZTt1v5gb2xE0fR
1cIvvuEIXUNN0hxgHN7yok+LWJJ7boKY5fb0/emArKeUtB5lajR9URoi83Nq5wZq
yifpEkxXAG0JeedMFvvRmXNaFZ3hA9AFWzKI5BXShW93FVProNd0dR19bGxw09Gg
pbCMxfzHpKTY9zHUHDfowFOOzl24Div1B2DzrpwdT0D0eNoiTQB160/rMHEtw0LI
aoo639FhtJXpgtqyzanGfFDJJ7zJP8Tar3wFUnLMkRMAnwpadvNsxq6/Javsgs1d
iqqFtg1gl2uoCo+WZVyWE6CtF2/9c0fPpcCJVMvW4JKVwkZM8Fp9d1FTy2rlq31u
hK02rJARnPEeFOTnfXagZMXMzJuv4FI8HNJMv7meZeIFGLbG4Rowoo84F9TGuRdQ
1xyw02xXCVga0CX/h6h2i00GWa7XpS1C0MpWNL8muTM+4hcwefsqj00ZXh40guXS
c6ttd/pSkI4GTKFkUaHKjd5G03XGRxBvrk+Rk9RNG8xkCVK5o8DYNYWzgYsd7eGe
e71E5kdL1WrlzeLvaWq/I5TiEFQ9DvQjGqa2AlLMx+Wt683TuLzW+QkpgbubRwLm
cQhUFIAhrD1RCZlauQ+rvj00qfw4s57fT4ZrYccxmzuHITFGlB+AwsniztkS+3dL
rx5SiJkPdxPoupaDwk7Q1vSI1orbT0VtK+/A+8VTWvTFtDp8W3GP8XGALrdbMfOk
6fpMAD8vZ/Pri0IBl7u4zJ7wgvJ1fFKvVAZcH4i42Z5LIOKFJ0kATtHQbwCIfOlT
dasJeF5u9ozVhGlV1RmeH/WaRg3Zf1o+X9THNStoyQ8vzP1fFr4Gft6FwLlyOK9T
v9+ta2fs5nZdZiGitseqP9sZRfFcsuiAWB4rSTe/4APYJIupg6+t/QMkxMl3yXjh
wMZVt2YH7WqvyFIORtIvx9r8PnlFvAO0BypCpyCyFS1Ax++N0RQYeVYrMjk2eJSC
o3qDI3DApvc9pu+wdFDRAVq3NeAdO6pljE30lDEuCXn1K3+wSLPpl0DTaR1J81ia
MSZqQHqEyNcuUQBCheVThR+SZoDbaBV3q20X85W1TLm5Ke2HQLKIuETN0rClBxHj
EM238xTTxvzOeyKl9Ua4ZiwoI5m2FSsYppHgmm8MZRRcFmnOMVTQ2cmfsBcCc2dD
b1Euo0BcPAjPmKQ47yT2iBxgWxxj2TlEDZo6ZcWAV0rVpGggjjglwi9wRSBX3dDm
eWVB6IGF1Q3owsnnQ3mzNlMKfYMdFZZufxSehRVj+xE+IAzKxStvmZXnENGRyeWK
UDav4rE/NB5I1+d6A2FymUyr5bYL4ZjTPlvxInY/tpO/THZelJnjetgom/1n2ucI
zzAVHDBEwe1HuRKmmL6Tm70o5u6LCkXb0iweRzXjpYC2om6w/MPcI6c4GKlc+yAC
+FDhFwVgQjC8FAm3t7UtIFsQCttEZo7dSOJUmwSCKI6vWG/JRWW3X4DfqGj6kQYa
imPBN8uXYVYlaiN8+1+wn/vnxbf+5IGLGw5U8Cn6g0D3g03AqrnPxmLUCW7ZnxzH
eL+BYbCE9QxWnix/TU/pvQJgbcey7hJgW4Byf7+E94Ep5lU7g7fv2aCnLFxYlCss
5tBPDD6IaIgjKYPGRuZlMlggOzyxTrCJLgfx1dKeh1mp0FT8fES9YYOQrMtMIZT5
1aEsfbcTV+cxvFjhUXwgnJ6D++WOuh24gB/mDTbOR9aq0VWfwvKglMPC9/966Tjh
ktfOHPeaJ1cebGIwt8wLJsRsG4V7LfYPZoVwN7ldf/AIVIK9sa2OcRh7qprvlQO/
/cTeUp1rMJZCjfXQAKKLgqAyPSqfWjmMM1WlzqmU5oi//kQ5jkBp5ydXGVCFFpYz
pQVEpxlw5Ynu9NcBl624NYDNc7x8+MiCzn3AVnp9Mb7W/W83cnFubh0U4lY21+m9
8NUSXo2NX2538EuP6RTYcVsjRC2LZ4Epp1sHYFWMS9bD18D+aZxDUixc26QBmyJP
UnkU9h93Eggh5FQedDZLsdezJKMIP9Y6oU25gWEX/RdU91lvW/3bSnpzqz8miBb4
c5hjKWtavkWizYFT9/dlJ7UHW6BSQRg0k2S3lw1noMmz4QBlhfYgiUMCeQmBJqTh
ezbjyoq7I0xQI48S0xGvzauZJkG8S4rPfmaMBtuulVXY076+JEVuYY/dBag1H5vY
SOBDSDzdjG1WJC/YW4fswireDjV1VLgkgc08qsjWbE9r3lXD0N7ZJhIR49Z3spud
DHZC8HMiy7IRCoakx+ulAZvAnUAo3Fbfd+/HK5Vrd49+HtlbHJBD5yfus4o0VzdU
v2lvFoQ6G/Rhn44bqeyBH7cAQpxfCxSZtSm8xVd/DWEGgfLg8QtVusVgmIpptLA3
x0Mudssd/MVXxhJ5H9IGFaTt/taxnkjwaPVtfig9ueUAC/B/7naEUD0yPWqorJ/n
l+nIohVhH5SAJ8CIF1zzW5lZs/7bd6QYO/ww1OZl3BM+cgZRIi3O3Ksr3LzUt29I
Ho71jWyx1yjAFlLJFGgzH96mE6K5gR83XS8oVCW6y7e8GtyRSi4fhjDwwsoQ/rGg
/hkA0ZXRU76tN8a7arAtwfYYf+ypMcQpdm7mQ6ymf5tXUoTZg4nQ3yvDigT3+PfB
xSmhzTJHS4FwBvXhBTOYh2+CqdGQIcQxtJt7L1ZDReWFPH2pmznhz5kGRWI1nF7X
CDXCn8xtpatmeieLc6eVgOl1tY8A2jxT+Nirv8x8jw9oiGFM1DTnHQ+DZ2GIHa9B
BPHHaSzmv6bXj5ibPWUG54t+smPYI+VrH7OFSo13Ewjo3OSz6Fh60vfHK4OeqgfB
CHQtkZ8Um5WBRULIZADHG7a4eRMYVRsPLrv4jS7K01jRbW76uRX3AbOeHVQdo/6B
y6mg2hjf1MUXv/Fa17UMtiz1cDXQgBaFS8TWnIWWPGdvxS0cxPS4C6s0oauhiT3J
UmqxoQU7usAW9a2DtIzZSSU/1r1d7gGz7vRTxqRAAgGOHoWvG4+K8qWQdRc873BU
G1eVHQDw9xUJ147g2sewbR2PIHkFY/QIJCV/DyCKUf70otSmpjSODhJSY0xgjxkf
kdUxwl+w1zEaNjAEh0RYahh5IDw24YcFsj3/jXlqtLSCr2ZOCZ4BY6dgna0hsdAs
Za6eHoy+ABuce63Q2vQdcvjxdUj1AVWS9nm5wAYflqxiKFdg8H8PD8XIsC2eywgq
FkJbfdSUI+S+kHgNsfV8KFvlB42o9abuJ4Ur9Xsd6DQSnaa9sBleiObWkASCRLJ4
p+FIDtZ/EtsD+ZlRCkUztFqRkOm4/csRSD1jw7TpsR3g/mVO1WBzSyHHH7sIV6HO
aKUlaGyGwE1WemQaoinEX7jmWgp3RDJAIjtoGH/i1g+ZuztOlIcanknV7IB2Nh7O
/hAVD9iok+Xnu73MK+fW1pHncG+7mgQBIzcZ4zpKHmKOEpdh7W1p0c49dk8w2PMd
6AB/1/0lBffW/xRtpAYMZaqM4/pFStFFNws1+dVrwi3KpG/CH8kDQXzN26zHFiyr
WAgdv9ylHOK6kSJ5FzNS7pG6c2r7cYFccsU3/DhmYDlMN7dStV7FtH6aCR1YlPPk
XNbJ+dNH1EvLmqFbNXdP3wzl/ujAcN5B9WIpUMrUAC1Jio2HY6KQXf93xcSsB5Ov
M7jSNMSJUd3o1mJ7/erm8YaFWVnnTywgTwttBvsC4EDTrGc9XS9azdaC/mBrQSo8
MSAmmQshCn4EUgQe5BcyaArOMzmQ0XEl6l5DzpUvCizzP2o3kky6mIefHP4X+6yK
C2yCXRGfauNsnHN9U7oGe/AW3c4cy2TlRNmvlxVWU4cnIZMKPWPSwmAxPX9f0q1W
6mF6btZyK27tyWzWr0Fwik8VqYd+Q1oyyhVpGrs2cFikdsTU/Ykb1nnRRxS890Y1
CjY+1d/RGjFZcTCm9WHLQgpCBlakwaflbnT7+w28yp/zeevcep5iJ3BxOdXMdsyZ
+uwzhjwQv4oQbBdTu7hh0w/T7S9LI1+TWNxCk/kM/sJl/qYnBvYMNydnsILib1Oz
e0/IHrwK3EwVDBaUOsMEHbhs6KR70FxI5t3Bl9tKyB6urvz/VT6QfFSfKdb+McWw
AsNux7pPcNuo22F0qpKlVJCnJqi2hh6wasAeCkcpRbRSUwWMbz7bJDEyAKJskxvD
8YhAq0g41ptN7gR6eAII3Mb5mGfyvIzcFu4xEqhKIud2lZucbdzPRvaIIVpV3NUL
STwOxWE31qWaScF1yde/+O1QbQP3et9P/DMm2ygx/fYyk2uvsWtTyyg9srqfyQDM
9D9C8mo0Reib/rELdqMhE4RRfQWRAXAm0N9HOs+7ymcUJBHsF2290eZlU9CkaZM5
IphG7KB1oIZ8TYrLxt+WLpc7zMFnVblP87pvfA55pqLPxdfeIiaku3GAw3FSNxHH
71e/M05sZCRXrCXUXw105SkQp8VLDDqew9/Ij7W4oSKt6XYdjfE4nElShwpbRza1
NBcBa6ojJjuWFVQNmd9rqWiZiEeE+op2FvzBwBym+QjWu4zR9vlZy7ckIHZnm+tq
m27i5V6AQiO40HtbRNrJcBL8r84Fl+dV6vSqvXnSKk4PvWcNBF6Sbsuj+HHefCAw
DK69GKYeEWDErYZMNX1LTSZAjdm45BEcPqmHpGKdz62bxhP/xwR2hmB6xTiKbQI/
RVdyJafPpnUWL+ahjWWLCuXGfOM4FuwqbYTB9gkDyqOBSNlyxwKfBnBbtFI4+QK5
45Z3tZHapaT3qCIFswsuyWYQHjmtw+xs7D/+2b9Cw6Ro0p+aLYjUYfMMfOIgOI98
Dns2JB1d4DUtxNJmiZ/gE/AALNfWgrUsXw4v03KF6I05y32BIxL0ReekimrDxodu
slhrITNCyNPzanzlz+FdTHhbjAG+ngw4Z4NxK2V09YB00Xp9ytUahFccut3AIcWD
v1X7uFzZxaPeAsDB3xX1THq6TvASzodrLwpKCRMfIR2Up0EnWPMnaUP3uWXQOCkQ
DF8VEgeLeAnSMOjQSvaF6zgXnyHrrpNLIgQyvBPD8p53cvrI2pUcvLCjX+SDK4/D
6L8+7Rt8kBBwY+Jemo02ZP12Y+UuL0JSrRQD0pSCrXUVN1/FpnYGr0VsC0+W5xh6
src6iHARyrnHTTnW6rOHESRKg0tARYjyMV3L24OGlhiRNwX3ojWjz7ZPpEc6luQs
PDldhLfCwhrB2XPXKhhFFTqiqliKGOtrK711+MEzWi/ftC1zdhUGvUObGfTbtxiL
6/WLuV8lHxatmlKdUmNd3WA4PC/hrZe3cPhopfzhXK/5+r3PInWmqk9cnLEUWLj/
mSG7yif3rDL6JMQ2pdgTOE60i5RH01F2kM/iC9Ew7JMQT3EI9EfrR3k+XLr4hsHt
CCIo/0DyoSmMsi9CbdzFtLm5G+E0D8VHLppUAQ+imCKSJ4bdP5gqVWwoBWn2jQXr
RjVWxp5v6kgdStof4ReIXVg6C+xFJUT4sthMKe88JL9uOY0XU6noiZGI62Z/6uOn
f5tGcpZqyuZHRKck+Szj+V6Eop4CcsgLNIaCuTrVi6vGLvd4pmKO334xcrnKOsSd
FpZ+K0K+Xyk3ydoOm/4SIwkvvCq+F9rzm6IsOX1re5NWV9zgiLraPYpvbx8mUQ94
zacTEhJI7SjxBM96CU35ZKSjTCyOJ7XrsGJqRMDy7t1+NDL3AdJjLFSC86aJhn5I
RzznKc/FPiWi8w0QgFKqVjI7V8z05OnLGtvP8ip0HkY19AxxHBm77fXNN7bi0P03
x3759m/Hj077uTOmrQY9qOr5qy1uhe93N5kEyaIoE+2hdlC+YdjBQ6MxOKyQMaW1
+umad7Dlgwgs5DL3SxkEJJaZTzIddXCXpQdXhIxcFlF2LqgRaNFhSDhNOzOormLe
oRTAphDsUoOSiFBlgpmN0g6fDvw/3w/yG/twdozqWh89Cam8MLhksIOwo1nPwzY1
ccU0BdvD5jkqBUzvUJJDvouZdyz2mEJpmZRUYg64QrQLsBCkgtBz7MtbEt1pESeP
PXWQZt/dpfd6Hc0nn3CDGWNur7z2Z12jwkUGsv1QFWvZMVzQG2/S+seOhamHvdN2
6t8IH1sA7CETux1Vnfiyo+UALk9jaJblWyl8K972h5v2XJkAVgY3t2nxU/9THcjk
CUMaT6vtHP2FWvIcyQ2ejb45VZBzdlPJ3GaJTjtuVvCNpNxMofczopWiJmAG5I0P
BHD3e823lZk5A8kJ+zPYwxyWyRtmEzcRZ0owEsy4U83QCrQr2WSD7u4KCmfq0ApO
C+sgnWAtUcz7pFP13SYfPsEPj0dzCX5Pz7sOCbvwnMDh8jzTjncrz4rAM53AKVOz
wTH2mx+8o6ivY2Rlw3cyINTqdcGfKaBiK8q7LbZkTbJVJeLnldTX8Bhvr8+YLsr6
e8P3es727xNoCCVD3iZcOMC2xNsiinyiSt488gKJAlGybYno2c21Ar9w4wDOPoXo
pvVYoHSBTGIi0gtU/VTpFxpD8rS5cKNo7qQi2keMKKxHhQ4QdOWubyfjrDvAh2qw
e1PqvI1ymrn2GV0rKGMvVDWTDmYoeLI4arJ3otKps6/MukIPXDTFYoV8gkGuBC0s
vFGxNKhwlMCywy6z4r0qxGrF/YFiHbZlqvNsW846z2VJEHS4E9rbQyJMZjur7nY8
ErEAwwQWfZ7UfI8T2Jl1oHAmlXvZ70Olu07czSzXMocOpPEU5wqGRe8OWD1HZCes
OG/OLJcATtnTDX4EWsuIkNi5+qyNZdzVLNeaAhVFCJdThn9sInvHsovRd9SDh4GV
kp2Ej3Jj4VFwfQrrByadbU3PrOB7RRhEKlHqL4+b0ucmo/McWo2HcN8+FYRIG00y
k20OSde/feBtDiEqTwTRrxpqmjwUGsHvalsKb8QIY3asKiUKOB0FQCoGhe1yPz8t
1WFmjelsdaF+LZbJUa3Z3M1wmpn6STmXirqxK7AZ/XvGDhISdjQghn41PozxL7RY
1VvpI80KreVC8VUluf4n8kXn0+XLtpVgk3fYoh1XQiVmUtYRiJtXKi+Eakijqvj0
XHcb33ESFcVaoN7S1ul+e/UCoi3oVm4mvbG7aujYJ83gmP2N1M3yae53e027RsRQ
wU5c/tIimRY5v2aKasyoqLomxm3ZXhPXoJP2DczxmvyP4J+dI2Cm3QwA7wMxeiDu
pAX9ygeMC1m6SNNIu+dHc/R+Dheb7D9TpeFlS+OgLcrmahJz8eJ6a66B12KHdlO/
uNwPfUIsyoc/uVWXufSx3YdjyorwR4TbhNciAPeXHyHJimmqE3Y3vgtgx2aRs0CA
0fWrcy4FZ39nBe/jXBBb6aJa3Pb02iuWy6tYOrGAwjwrqLpwkwEVgjOdf9fGMQGu
KJ6sIIIXB3SEoHAVe3nrNWMKaHX6Mx3r03e4OJTzUog4xNC8fyUjIqlgNkoLXZ+r
0qaPUxsD/kH4n2ZfJYfD0SnuWSz+p5sRSBP/Bzu2Xpt4gFxcEPHhWoh8kflc75US
UH4Cnkhgl2GzHWBZh+mSo5XcUgyeBhTbASxTADsAmJwncxzi+xFKglhUo6x6vnzY
hlpvsW9UCn0hpwB6uDTsrnlWAH0Q4hxciu8y1wng/6aOkev3yAbXilEsHXp8aDir
XjvuICAjoKKKjRYXEXeSdzo+IP6e3ntOOIpnqsAmOiNdLfLOjlKouZZa//0fzivS
EJFaZgs6AzDaW8gHqltXqhUc6iDCPrLQLZI8YtZI3muDt2LFbbIGpbDGVwOnBr9N
7z4P0wsAcDzv+pQliB2vQ6VFzvCtzD8B2hSbN6rUGzBmRrN5p0N/NS0Zy5ToZ1WG
9AZ/n7MLTDAmAtP4yPg6llPN5n9In/S+/3iztExvj1uQWogjOh0oQj/uZus3IBJ0
f1s7378YcxsK90F8dmD7kVexWqot7qY69WZoxptWYX4cqXj6aq2TPA/Th2/ywe/a
vH92lIef34/DEV2gtJBOyqq65bJMbhAnlKOg6BHw6Cs0+kWbDB3Ecfuvch3l/qZn
4LK50PyXT0grxp1xFY0kjLOIevDn7++0d39h0Jx+auCS1pEP6fvxEx2LULngyjGS
cH3IFLDRxE6ELkfLZjNoChDIo3y+HEQLAU3HcEwfkFH2Y8FchaADYnlqAY/MAomO
EZ9WUKwTfxbGhuJdPgdMG8CqR1qY/+jkKNd46AE6qOioHLTes4ZzhgzKbu7kyuYf
cgI387kPlD4eL+RZb7VLYC2gW1YY1ignKvREUMhqx3xhcHTJeyjtFi78IpquqdnA
3R+1jiJm3mGmJOxQsYz4CPBsWTMgbqbkmiCAcd+Jsyr8rRrbkbF5z3/RcXZgmc1q
PNfwETQ6sHSq5jSeWZlzhCZ8+D6MvcDb53kbSFeU6OeIZyzW8KCf9NQUTH6E9B3W
iFV8IExV5iSe1133FHZOgYZ8sh4P0PI/b+p5Q4YZRXOh3bmN7WT6gbHRFPWYBHvl
azpt8vxWZho0aJiET9T5irFIqiKAC3DEtSqPNCl8aRS3zTYjvmCSP3AkVmfOILGr
f6+vHX/irEOYR5iO4+3g3uuXOtHj48LjRUbttrJGgdt1ZUeha8e7aCg9yo7USfsB
Vh3s8/tFTJikYVrgiVJ7YOfBRWaztJxMXSCDkbS9UUxVG+lTSO4YWLbUss/9G8t7
Uz5oXIKI0YAFdDDsM5rfowm815um+/ikc70r0kZmIsZ0oIO2RMDyoOQgnflABHv1
kPmlpGJjBNHnOcdta1h8ufTtSOxrLBwwjzJexDa0NP2JQ/pLX5Nc3yw6LxxLAeUC
F203NR/LOZ/RJ0r0+MNF6pVVLrP95s2TcYslmbfpDt6W+VloObL5fXsr1l+zYDJ4
ud0wKre4R8OvOX4Y50gae9c74aMejO312HmZjYwxMHTWHPx9m+j9Frtyo70+piQC
gtd0As0YkjuoaE0PWiDqwXjXL3+qf5pQFyKxvCH1JgWVjbcpz/Hs88HC+kxNPnmu
9ki2tOWTBPo/lK+aaIudr9NTpZck2rDFo3ufsd0KPZzPPdkxfuc+AD1oXULzxuPR
4S3f4ilX40NKagf7Q+3WambsTVsvy8+nWh0i3ak+b/des1UbR2SbzVAamsIR2AiS
Apgk181Ps9zGbjjnr4q1Ab4zwTnrglPS+o739/259/YdzwTjCK4pffiFUeQ7YEU4
CMVoX8CKdMDu5x903l/GWGZHxXaGOfHAweTQVonyZno8u9Td4Ptj5gPYl5v5xSjK
nS7iVMJB1VL++HDZ9J8Z0QaPoeC/NqjLmDAV8tTRMR03TfHWweaNdjZbfQpxoxFr
TIB+dgYwEGSUOJUhBzXhmk+fbS8k8f35/5rzw/J9PnaZXLuoQmqMOeYy6dFqbze8
kSMcsVD1uXZkKWttTwVrdFlCLOjbMtwLG2SImA7s4krY7gRUWp2eClh18WFBTBPG
qTGeYEs9w7rojhTd7BTjPgr4ULjjOlXRt2L7Ooqry/b7Io+KIax/ZK78GB7PsnC2
yQy3Wrqrf6EjEdsdLyLz7ZaMciv2ttYQVsDVaPt+jrRu+BLHbHI7okKe6XwJDy1/
jXj1HjxY4TKCAEBYRp/OqeqxmKaI45KCuRZMzIUg+FKW5TVtvorUv+hJ4Xiu2rFU
WtWA06R+mAJGaAiKvqyMuLq67RXg/D4FMh5rOcJAGIZ0HVrxT3zijGff27ztpNOf
FBD5q13BngbAvmNyIn7RpLVj2vxRDbQjBAZX1I1SlTjYbkt27xU7D7AcRlmZtZiG
JHooLr56+rSx29dtCYkn2l3ETWY/XUTSByRlNKf1Ml24MOLx34Q8VkShYzjYKDq7
gpr1lysv9bo4wqgD+gPdPs7BFr6YxOZLSUVxOgIxLRkbAdSGT5542o2SgDUVOn+Z
9h25vkQs4O8oauLZaLFVXmSznBx3lcpKhlSusFnTziw8koDtip3TCUz2TAP1fHXJ
180fIELp+VH9Ytzbc2wPYEfJhKaCjoIva1XAdT4gW8GvpdIti6asfRJg0e11oYPl
uf2kSkFMg1Sh+74EP3U+dbzwCoC5wBzezC0yX5voQ5jVHb+uhgwM30OKJVTZ3401
cUPPzXJ6qmvYgLfR3PGmu6CQeSOQ/yDtQg455Kibet5/TsSn3dUvEGXXMPVB1ZfB
jl7q2660PzWCcOgfYY5Pb6MvMilZJfdwV0sB5/OoMiejuzGi/B+9dDuQVIbwjSGJ
Ejwa4Y/OW6abieyuwffqj0lEStxM19K8AIj4E2jKDD8qzvUlpfbWwbkvOT0vzuVH
FtRyNeCY3F8+SmCjwKqHpGp7SZWDgtei0pPIJiMiqWHrb6f8d+C3RejA9aF3Wc76
m/zfQO5KgiUS/GytjHlVuf9aOaN9p3wZ8ukwG51pyr6vov3QyngMLNYQ03ikjBb0
m4dHNS35fc/ezZ4X74qTu6sVdPIkn9S8/6OdigSUIQtLewjBVjz1LsAWPw/0LZ6E
ovcVUyYC9ThJoB/gvcDNxZ0zLg5v6tCHaqRctNhtA2Nmok/MDwYBbtyGl/j++NzD
lFu5M/IL5rMyJ542HmRXcTNoAFRVGfOr/0B+U/uI8fpq3nwklI5nVaX23JojSf+N
PJme43dJq5R8cYZwdl2gRxUzsD1hy57UqaNKGiXTOGsSQYCK6TIn8Jd04iW9bGb0
S5zn56syz0HhFa0tTeCFTbWi2Xp4UcxNdWRt5M1M1sLfXpF3z/+txo4DZplY+XlW
WbLEQdRSDQRnXOHQSqPy5ypYRNpii1X+zb0pfCLfpyNNhqKfNcDTOqLlnrhMpbtN
Rk1fvS8jlMdzE0JweSXsO61bAj6zx9I0HnzoF6QQ8b1401V3m6Ud79+KY6bnyWlD
mNO1OBhcNJdbnXQBxXZTwxvaYB9pU1t5/d4UADtvJjscawbJyvodOM/+EKCgFCnY
66fmVidEGBBe6Bt9R0qcYOOgrpqHcttsTkRL4ZoBCa9LsnhzpMmtfWNBkffXgifl
4lqbv/t+bbjsPMnKK85vkTaanYRh11DfjLTEzK3lA5H7TBY2vGRRdZ7tbRHXUnf/
21Rp6SCrJ0IGjFI2gQzob6aZDMQSlOA406c3dfvisgjQ3VkW0slNbc5X+1VokJ+/
2HV9GVuNcWQbPTNKewmXbql9NwyGe2jo6IFXHynNGI06+nHXyWwfB+X5CEbW9V3K
KA9kE2v4RwJtYNZ5RYWVelB/aPuz/iiO+1mB4RhdcRSIiujxYCjHkE50ADjOrFfZ
QodoSTjeg9h+6vLCY/+n8pP07vltOWew7T6+Nbywn5wScTrxsdCASgCo8lFGgiAn
WMFyLCS2+1P6KbG0OARHbiTpDOAow6CLgAZz46aKoNhcV3Ijs24YVXsJkv2jZNz6
o2jrFxUcB2RFDiCM3edo0+OgqPiObcB+nxj3snzOl7ZQ++3EKd29JK2VGJi4cHcC
5eerVvHcUWxnfq3UZpcozKxiLSIoCjzfSkqNFqSeNY/GAETOB5VJ4Q4zaUFka5fr
YRwb1YhhSl6m1FchtM6G5eFwuL4kmt3KQhW1ZSIDZaTYKPhnJw0iG5mQdw9e9YZA
t8eGWNhZW9fzqeYUVoXeAWl7EEZke6idCQA6nDRX3e9Y6Ut86ypgtiTCM4I9s7uZ
qAoedcG7/pJYBkVtpuOA6sk5ZKiy1MjUaXohlv5e2LWfuPm6ROOU0QAQP2Pm6x50
zQ/jgXox2fBnGoWilyxzipltFZGbRbBcZTMbLimmSYfKy41U4p05byURetu4bjYX
24bTS2Rf3O6ljb8rdwiR7zz/J3DDBgtF5mQtGyPjlBZ7TC1MAjLh88AoiTMgZv/A
rLxZ0u4Vfvfasvw2WxjZMaRvshYGmRq7bIaR86TtEXmIJwVpOsQrBPiTYjEkCnLN
f2WhqPnQTTiu5qedDj5LLrXbHWZy5viU3Yq9uYInI0jMPc0WU6iCHrBZYZizhk99
Id8869K/ADgAtLO8IhhHyQ/5PGQCsiWJZyK0r7KoD2+mNtX0z0VU84oVkX3OuPI8
bUqRnEq6BUfRjBJ8aAY9c/r1AG5NewTBJk69QXPKO4jncKgIl87UoKatVoxnrsco
i/nvVLqnpsbqXmNfrmGgOTl9u0aBqvyrBl7Ex5VSd49Rp2PUOrWlaaP/vVBl1P+L
Uo4DzFag4nH/1pVc8uIKm8RByhNba6ttbK4gngDklqs+zaOJM06neN10fPQ3rqtn
KdinuSu2gTxXIA8Sh7ULU8s2Va6a1rgRGS3jYtewiKOO/pbLmhDvio2zyYqyW453
vX9rBz6hZ8kFDbI8Tt64tGrfX0N/5IMB7/Ce4kfr8UhXk7JQXsMB4NrC9ZRXob8J
qAa29UMR6uAOMJdTHTfVu8jYzxiEc9lVgipUFW13fGnXo+INRL19wcsRc8kyxl3F
PCSEZKjJbBkF0oihEKtMAxGQWwblD3yaPdvYchPwIrvrS9cixNzbZA67cbZ4mevR
v3AFWhvdTTj9oNMrpDnAQI4hE3qo866TK3e2CUNzhdLwICayoa3rp7fkNRJlABVX
gfCZh8iAIrqlLavWbu0pXzcveksvPqnZn0Yr/VqaiVGzwwAtL+6fwzjNDuJEnrhk
gOIQJZaRS4M9naZsPyly3knBuQVOGf90EBVtJqNt02sDVHmbaC4Q2Ny1BJwKjhmw
7qmomnCdHWK7xmavObMh3H90WV6HAzmAi9xW9fph2Dztm0wNFHKQWrrkuCV9VQAX
nKsC+FBINu0PZbvFgRV7PtHpttPJ8KrMOhIHGRny9XblDgvgaZ+7OaEPZNAZdwl5
O5dwSWcYYrzNbxmP6Y/O/ILcZfzIEmFQlvZdl5vxmG0/FO22Itc89AS9hZDAGzH0
kR1ykT192aWXaoKy/Qrxd6vLKq/j54S05zqmFdkXr+TVvn2gOtpSNyppZ2S3K1Lg
Pzso1bbtyfeUAQ+j4pSK9S5KmsRVe5Mo/zZRDFWmvpRglNGKJivTwmCpc6BrzE5M
nAOgtG9B9F/zFgVQRNMYzGY4hEQsb4IUtUl0lnVJyNli13w2oHtB9ySmGlOx4rTb
0pPuoiVVLbhpxVXC1F3Y7lxB7ht5CEo8JzFHyXyZ++eyw9nu59tv0BpCBiqNWBUG
8gXe1LWILxSACf1/tAAHRUgdVfqIhC41J78LzGhfLgtOvYgCyDHW2XzEOFHU54Ug
yB7Sy4p39tA3QziobC8n8eWVSbgdC2b4NoLPWJIqBMRju0oOU9ze78hBog1Qmf0r
4Qj5G1U7OZKBQyhyG+XQlznQtKYJHvrXBF1HEcMHNl/hC/F5uDlAeKK7ajnvnRFB
11eQxGNsBBKvx2yONooBPAJ0NYxR1hIA6o3/SFn5WfQuvXlEFkAOYpcfcCZAhr5f
DhQRV8Co7e0likyThEI6Ghkj6jTvJ9YZeiLgpivT0KtVblXUFmRcwobmElUIBsE0
BS/m1IL8jF4TSS8JQ6pIsyz7Kj2QDwEaMwopSXBVfZYs54hSxQC3b8kA7hsjObhU
RMg4Ile4x5thRW9X4Mv1dWUIA8LgEU0DLUUToiqoL012kaFnx6JLkKt+gBwvruCr
EhkhEjkNITXtlCsiXV9vzcxcVof09H28JVbTOAS+N8CmjX4d+YWv1sG4qJKFlH+8
OAG5fX2pdFxfIDVo9wtchs4Xyx91M+0R91EI1TRy1iTMoiYAHq6QoKqp5hgjpKp3
HgBu/oOhqr5Tn6cvePGrUmGrKjRH72uPNXoWDsl4aZXgaYhMJNS+b1bPQAlHh5s5
QuiF/r4zN7zApE/gpjJTpjB8Ga4gC6VywgLvWNnOCmXsigi4RygJGX9Y5RZ/qnTq
GJB0YZ95cZ6TlRmZWjdy04zQVkSYtJDvmkiz7nwnk/X0Lhp6A/5hcKcSU8GiH+Iy
J0j+CFeNwNpe529nyIU46Qc2TDLldmtf4gtpb+azMja2I/wYfFkMsdJhAWkFfNru
X9LbTvP3hJcPPlDWcPhWbeKcPULcVDESBr80bIdvnESJWJeFPmit+osr9+TEv0LQ
jPt+xe0CuzQ4j5jH9ETGsn2e6WQ2VvLvMe+Z8Qdy/JMSBFjYEztBiel2G8aYHrkL
eg6jcOmhhBrMmHfAH78oH6Uh+SRn2ysOa218nFrJopHRaaiDCZhl7Cu4Vd2+x3y+
cPdJFom+hzvJynuIdffJ8pvE43OCGUfFPAd5tl1RpAujXxrOENH71OknAKV8T2VP
ExblcJ5/I7IyR6+rU2DJEWKoZI8U5zE8CFKoU6KklAVVAjcd4FMbjETfm7HYjJj2
UIKHRu0NroMP+eqnpuru50+lvW3P0VwrMFUMkjX04TBkCqt2YgZRBWFfQDF/AqWK
0kbFp9EsH/CXL+G0bHGnFpFh0reigIME0fXfycaaAKWKPuO00QwLCnbRgi0tV+Eg
6FI2szrZE+EbqnrNu7nXNjbQy3ukd5hhvy94jFyDvVcisTq1DglsJSDgEfCxe+wj
6vtVUQxGiGd0wUaG09vdzrCmOL74nQKG8U9E0E2SMmaa4y0g9VpaBMFu6+BrEVHh
adGGu4xmQG94foW6P2OtYktcBff4RmWrhSfjAcvYSPq0E+RLv042ecIedrPk7Zy4
apx1U9/r4A9elMNwj5pv8v96iEHpAI/rHVoYQcapzEbV1VIogfZiuhf4W0DJL9pK
f1Ch/NMXqrsZLyvcPWOVW7zk1OdnQsNDLnNU3rfDhZvUE0veTSkjbd8zDmWnCVb4
LBZvh7EaWoD5GUPse8NR0T00F+7rmeewhksE+FygHvh+YMs5zuwg/j9SDHe5pFzH
uRKnyhZZPKO+ggLhUV8arG89RCj3yrywufMXfU95Z97Jli7bL0MxeDKHWWUNjDxw
3AQHfgnJLfVux5Wvqba+2+D41CmEuTBsRCQxeExWTT3dzH8gw9b09X01NavbLxrU
PCJYJAAk635cWGH1xTsLsb/ZDmNl7vbe8+fqPCCCSOANqR9IavzmfR0iFOVxfsSf
K7f3viIWcro9cHe0lubmr7jeEkTnFEGDT7YSwdjtubAr85RKEe6/ZX6Jy5l2Lx0a
ysM0+sUaPXUKIJNHGSE03wqW6XhKWuNJIE1nmUQ58MiPqLQ2nsrWe+9U2O/b9o81
cvs/+qnLMNp07Y6cAlMFIpdKuihdF8egoUm6/VpRHuSAKN84x1b6QQ6nIITcexNG
SiyQLvRQGldGIglh/Ss+HuwVil1kjy8UQ98DMrfGoVArcjC89/x8uzoDDYr1lDhm
s7r3d2hDcUGL6Z6r1lN6bZ6E7hyB0gi1192S1Z3Wd/kKNYKbZNGKPqB3xJGcmhch
9pS5vi4rqTQxxEuwBnFiiRAs4OuLZjOvRPXCIDyBeibsMQdBdlWrAc0hO+jgcnkn
EUFDXbKM+GUMrvHb1Jin6EayY+yl6Fd8uQVjTuweJbzzR/RL6Ma1B7fD3fRnRsCQ
DEraZXj2SmVDADQGGUxdzPjr5x0PQm3yTZ//GA848aF89KceP8/HQNAh6L3P98sc
ml3rZF7Qv6v6VhpjjpolvblNgrFOFw9K0vsRRU5o+YbV9yTDWe3o1EzL9ICOl4ui
oju27HzQDFDu4qXgUqy5J9oMySs8Qxi07rzbd4Zji7ghZqVSv2q2g4m3jObuIxsQ
Y7hsOceZ/qCgsTR9T55JCWRZ8VB29K2AxdWxVcUIVD9L7i3WIIFdDaS2aNuGeRS1
5zUgiEaFZrrcQ9AqNee6iZyClTfckDEkB7PaHN5wwXis1gpa4odekK6ylR6MAhru
NQi292xurWVIPLNpyPj+A7G85kfRZz0kSLtQSJnQ0RjDzg1slT+YpJY4MY1gwkZn
fx7tQ2q6n1Y6olM+Hm8HxHe0Kttj9n/69xPbRyO/eGb5yaFmbDEgMUNUbzWCFxys
q/VX8S3wiD/AGqUr/c9d9ik4xgNGZTr2Rqcp37VMeeoUpaIJoqVA3w7Sy9wJU3WS
toK1DsQkS3D9TnkA/WFu3Dvjv3UUpb0KzlSaQuwbeib904H6PdOA5+Pr516WELE5
H+eltPGgsl6q/Z+ekiLmBivdCccLoWYpVoxgt5N7ddeTSC78qg+JY5Ouz/xpsC4O
5YcMTVBAASOF4VFG+riNPc91ks5rL7U1J+DLI0ClqqIEd3gVfsaOwIUWGycPIUAE
Rhly4RWFyjlqu/VU3v9WakJwmNiHjODtLLMk4IsbzB6jamHl5HvfXusIEoijYuuh
IxObIo40aW5gEYqTOPBa4yt3WgNxCpFuBsyJNUFRsJtxfNnrPGFzePNYmQrQuy5Q
QkJu8Baj8StRFpDB9jWTLmO6/PKa6bhpRzulijTQLUTapteI+XpF7BMFW1tTsnXq
ZKFjNd3TENaYh9LRqLqqinnkStO7GjjedbbS3dByrFzFjwJCWJ8OFAoY/qTMFOQI
W7YiIbz7LJ3JPYWEhnoqEiLMZ31tFphuEp373OEP7+rk8Hpz8fdz81ouF1oI4xDU
/sy8oq3h96cUXyL3bab0fx2wC28zyAHZnSBI9Lm3IXVJDLJXYrQHb5Svm928u70Q
Q6otLxRwu3liVdAAqWCt4QT45UpoJdGdAl/XmFNiYwgVo07fx345xFl7G23C+VRc
/GW7jEM8Jss8T6QS7lzLQgEy7uK/y89MgGMLO1GMwDkjULcmx2Z+jH6VGgJYqUdu
GWRZi/IW2ibo1qhQ2uZsdGGVUC43cz0Btm1LTZ/5a8dlg+gaglyH0oRJpsGPaYKw
Fb4sBF8H/kwFnhUiNvXkFa+ry0Y4UvU6iRBYYjEMt+4da75vbCWiJ1SXR9onVfO1
XpKAftX7EeO1pNuBjIs5p9JCEHc3p7pX1M1FDErCRgErzEEHiBUQAV/7cPmDWdGc
rSflD/uRVXVphX4OnMsZJ3MAUQ6hdFOK0pbQnij71J8LZYKWdYYUOo5Qg7YOLUF1
Rf4rQ1p5OAPTcOb8tsvNl9XmubS5GnH/XVeW5LlcvCDMbSjk9deomCC9EWf4mjuH
O0eKUWeOd/FIb8btzZ7fUdCyGVgZWQtODC7x1hqyJEA9U+Bu5ooysmvE5pUFBRzl
RsiVxS95Mo6mvlWs6qeAj+2dsVN0/uo1YNhTI63+avs/eRH+11TVX60vR/r7dPLw
jCNMlO549/n7lLGb8vVbysukNs5a7gWKQcvyck/4PdgWlox/ZsvUUZGPe4xd5b7P
4LLkjDz9Uzea3yhnrjrru3vyYMuyC8scu4Mq8nP17qH0+SgDoH8pYkah+nyup2Rv
DS4MOg4XH7h1w1at+aCDvdRusJu1qIEIGqtGEg89hUJLGUuC7i4sjlsbLvy4kFGl
qX3TWVsw58ThJtRGTnQOnyR1pqg1hCbUDtyguesZvnASQYht6HRwMGdcUn4hcPdG
AHemOU6r+0ai+VjPJ8o4+3Ik0JtNsZdtefww3ydv3G039rRZ0JI4T5c4Vc1BODf7
SPhRLK3iOdBATa+IAKSpB1DL11RjZE2f6poEnz3NNVxm8DDcNcwsxlFVl6vZPWCT
+ov+3FCJXNaJJkshuurCbBFx0yoSq8yLWB9R7hXMe5XvNDChXmHYRNSMyPz3Kc5/
S0EM1O3lGSmSGHEl9muqJGMUAT3GSJ3zzvmZs8iq8AqBVM4jc8X8bwcm49UxQG2f
aYIPrnmoDCgu6SPTIeFti820sQ/lCc3gypxbFgZ342sVoy0OPJPmOpn9IQR/0gYY
G6ROzGzgViwQtMA1Akp1kGfTssjTyAhNaAEgPmRhHSDrlHOwkiubYY06YB/FW8KE
8YW0Wxj5B+kWVcmoxo6gua26zSuUouDdYTmusvzrWzrRsNYrSola1w4aF5k5WbUW
j/P+NQF7FtgknmW/1BdSGkdCnLdWp4o5LIQxv1lH2iGQzVlmlqPgWgBsawUzl9Db
RJsB/8rvqgX/JY7oSllslDOEeb33y1LzxP8o9zU1wRATz1pAT95dHejTVw53IHne
h1We0WtyyTpJGPJc/R6AScfGA5wmejgk51phtsV/Sy/T40t2RwuVX9S2JQz3vRzE
G65Y2B6ie2XATfdwEco0tg/7mvuLon1TBJZ+o/kMDy8JUaOzleQWegvP3N5nlelQ
qG8rRWOwPHpttxNRbe6cN3DqLyYfcAN2ac3BztG1jrc27XLL/z3KM6PRO3xOCR4K
RCkmXck93+kZMAuQA729Btafi/XaYUu+fE5rOMSsLLedMPS3k5ZwrPTxd18y7Lon
0rEG0WTrlP4hqNz5InzU5CNfIrDuY3gaTqVR3t8ujhq8n8ABNWH2Uf8NJj2uDZ9F
GalO5qpkn29SXy9h3OrSDprrTorHJHmTs+1fJ5PeaAFmX/rtYPtPYHAKpG1reVBT
x4iPM6tHPcmRgmpMC/O182xmJqiZ6qDH5b6MeYwAnBmtupLyNkxaV4/eB78SeqrM
iMO0YBZjAoSuk0QFrd0Awm4RcahvD3qidyT/WZsrJVvJeBRAZsVmfDohpf3tTQwC
Hm4zGYE8suOR74NXe/mwilF5J4/GQMRE7H2SUyjTffJNz8Ici+uKjCs/OwLzFWSN
Tw7c6niZZ2oJ8As2B1QfFnsjiiUfkqRNMXRSihTj2i/TGW7ODXQ7VCz1IkXwA+uT
/yOHaRZ8bGuYOR/ASdLoEgwYb3yce0vySiPc79wrOKCMgkkn4B4Lfn+c4uaj0cjV
BowUzrk0A9WnTP2xzCqaaM5FDhvCoSDOUbgAhFcp5UqvvsJ4kbPqa7iHYxiiFw+e
xVmX26uIZHYzmNmKNrASRdAEmXQRZFUZGAVECLUWvXcmWZ1BnCBTXnaEP0hftkgK
LGJGVgAhkNtldhZzvsxLEuz4eA8KoiuCz2EpwAy67orfTZDk8ucxGLUSeKrRc3ye
pgPGQG6MBaiXnVHd80lAMFiVr0RWV5vZ5NPfBovf0WFW/bhSCF4RS5wgPt+ljQWb
NI/NQNUPPPBpVws2rOCPTwDMIWmE3uE3PyeSiIS4CiLovoB6MS8OKd8gqSGdc7EW
IvFMO2r0A45ZQHrq8nmsgVvNvLDyHAUSzLKpxcJ7ix0BW98qV5LTZ4sWA+56yr4y
kazzdoPPz4NrVkhhZYX8G8LXXi5sJbuIyVr0GR66TYh2PPt1fGzqMiVOjITKE3PR
oHnMw7LdXbzEIQZPsSogxkE2LOtXjXHnBudxKczGAvjLWjVhuTtkhOmo9pl3aAGv
L4KhHhhq4BmlKGYQmtOzJ+EhON3mWuN44QvypiFPpDm1vdQFe7hvyXMpAWXpU0pH
aWnWTt+6LCZVa7TQEUg2cD3BxMfxeohdvLo/HmP2qjWcRgMwGWpsOUFjap3pMdDf
5J1k/ScdJ/gFhCB1NRlQmeB1rALj2ABQ89ySmGExJu1Hpw/818B3Rr427gFPxUi5
I3S7SAmZUK25tw4x+sY5AsDAOclkYXErDFyYZXM+o/asgJ1uKhKEDSmY0b8NWgpz
FPcouq4AKUD6dYle42JRI6IZScAFpElQWNNBBtOveKbDKgSAi71FmF5dOh8+sklg
kRJSPmcY2EcvLZVO/qkWykiwnjOvI00pLnsJrAdEL+8o/kP8J6o70PUWgAANTX81
H0sAnEBLKPzK1UxBkwsLMtPKg/vJSyurcMdljaSjHriPTerRUG9za+IH6KjCQH11
0H/q5u7YtEhCEaRHDvldxlfQ/jvQvFdsomsXg9gsU34XrQCaxtu5HJFRnPxL9G5+
wDgs/Bg2y3XnpWY5uHoaG8NTzzQjXbMcHdkqWTjpFetHGcsYNFKZNhW9FguUbIKF
CtWmyvr81SFhXv90ygMjyfsiQSkjW9vmN8l09bBiTC7FX5oLxQ8Dl+2bpvzYJNPE
Kltv5URXs3HHBNXbLzeJA6sHRCxpPMc0R4+Ay+3ZD4gOY82THulPHZyimuE+iY2y
bVFn6pnmkXSTETnCyMgvOjnUbS7BT2fssEVsVjpfx65hRPZ0bxQEo7FyVyQ1Gn9D
BzaeJfIeYP7tisPylQioItNqpxub6iFEVeX4e0LeXwFQq7XZ3RL00vIZb2O7U6pX
M1+maK5RptiPv3/twtjU1e7lrDKrUCFD0ErtOKddU6+84KWzhevfgSdqySh4H1CO
qrQ1tIW6f0A8x8tz8LY+UGhGraLTxjKe3oC8/YVjV3PXq5gi9xV5FEpS46yqz6oK
O1fK/6Wc4+MUulKT2jouGouQCC3sh2JwDKhfomoz8+vBhWZnUB1ficb+vo2HQ8HY
gcR8rM7BMgDUd8yhmNUKI4MJHFjDF1nv2/asIe9AGEY0Xbrj2FNlOdrsnFmx8UYN
zzzJjR2HDnnS7bIghWvFWxDDSCB5qSGoUn6W8Xcx7v1tse4ZUdzUsmP50quvh5+g
Mkz+1KDaBTbZj5Z1IuG3ZSraN3sfdqblIbmm/7Gpe/robS0PIqfBqD1Cvwn/N95/
XtUaGCU41XLjbt36+1sjdyw7XBhINEEnRgPX2giCfcqi0ex9K4ZzSJJNG3G1dY5X
WV46eFjnHS3Vcsy+I1JMy2cOzdegHJ3E/JohoqwmXSV1rSnCmyBEkBCRBu2d8p1D
5bCAKX6rOJHyvrpsUqRkt9jQZJweT3tuwqaOyTEs2NE4uyxwoFryhtS5MWsLc8cz
AtzghCfGpRI/Br2l/B/wRdvf/k3nQ8aIzIkEP2nse1vv92TSuhu2wm5cYFTUShiN
OVa5Y2/yVQ0uPmEkCRuAnc6FWZvVVqz8ORzbzCVazZl0oI6NgGby/tRe3wWpY64X
mCb4nK7EydCZvjfrDQsP8cw/sBPdk5IDkv6g1wXSEoKD2MUoc+MmKEGIQBayZCoT
uf4OJoCQh42qYjaGzJF5tzOsMgHP5bAtljCtiBkR/6q3ANjG/2ArjRv6ULFRW9Q2
ni270qz2N6pXoSbfYJ1WTQVJuYQagBydduz+Waz29jeOnb1ZpuScmIuV1MAfC7lj
EaMpUejy87ws8iy18xDPsTKQjhMiwAfttNSMMgSjviu4qWyH8qEDquXG11JbVPC9
+KoAhWStz2qdgvnt4mdE5BRYC71sIBCXmhYdM+p+mBmlq8qSBFEhuhT/eQRSNYOc
J232HyHBsmvmUbI/XF+h2c0S4uiaGDQUF6ucNFw4Xe/6cfOi5jzGHogv1bWmfIyC
IqMkL3SdamUSkNQg/8QiClbLoAjE9F2yPHh8o1wEh6gh0oM/XgE4GWCEskrtRa9b
oVKTFiTP+5fgIwK2Z28j+54oEtuPmdqgB3vRMctkHyMPzA5V51h2IW7q0sHcppQf
rJ81URyaaTcVsoBZzxdmvfYT9CRcZq81/W7BFy8+M/g2EKkTSlTWgaJqIkbCR4Xo
e7JXlNOOIgjUYfKJ+sZrCOwM01zQ2OgXxLqKzntatOK2NqstWOswzR2NdALnQCFU
cwloLDpRF5qmNdEK5VJojNkZAF/SJEiOxx6nFfdGZqv1MSlQwYj+MiABRaKqrQ41
7wmsWvOQwGEJzlRZZXf/ZEJVApegdx2cejDOtOZTqykzeYTqKEOcMlll1MIkTN2h
OxNAZs1WXSTxXlqQhVRyr5HLbpb5821txCtP0OOTk+DztF52tWBsGfJbLoq2hn6o
m6eCc8nl2wNRdoeKcQskAajT03ENtCrX3ENqrqHevKPpLp14Tp9fTairX+d4kMHM
RFaaChoIUExZRp28RWcEevp4ZvqwKJxqUKlSV9XIK4HJ0PPW9vCzNrorxwH2eFhA
9f1WLPyihO++HdG4byizd0An41T0wvNO0UM6b8VWzXLq48eMUKx6zzaC4xaSddKx
cirBTRIYg2JNLEHaUIcyo1H8xAIOx61F3E4UeetlaVNsQR3lWPSYBJDqeR6OcAXf
+595cXsV9Ab0qYW7aQMrexqfiLUkW3mdBcVvrV9bLWpSoM75mKHsVH/1AGJa8Wfs
XTBNpgr9EDbmvXuh8QijLTgCwcT0i13E0iOcozQUwwzzzVfksTf3JtFgfB4dHciF
FdXq9JsFtdpxe7vDc2gjzT3CE4EuO9/abYYYwk4cArgI7PEnATwo908XsqRGjBax
otNu3nGvCMTK+bmlU/gI3phrMljISaj7xmiH8QoOTCx59lSwPLIMb3JKC/otEOXi
IaAYjp9fz25stJtDbc99T2vG66PuKZE9q88qFuC5Rdnxb9DFWXbujftIxTqqkR/W
lwJ90/5fsSmF9Y+xgInRkJmESCHkbkahISnEQF9ls90r8zH2Yp/o3g62boGE7+68
O6jz+BDWiV419+at2maTmMtghd0K8X7PuNerO6FCRSRaO/21eNltfjIELCQdVcBH
I8XGcWMCliu8rCjcns/16l/4xIrG6rFVgOjrJOz1ZeiU7HsZrG+7FIgD7SGp8OZA
eqMyE30RRB2lvssmC3+WJKYVQubH1EWJbwmy0I+Xkc4es9zEmegaGwPxjlFpT4nJ
oPlsRtbnxtpXOLVlI73x6MXLzYhLCCgpMMZzv5wwy6zWzO1paoevZRDDuYL470/t
NL6vLj5E3yA7/sG45MJlNyqPCzcN3DJNfAEJCHaa3wNYqOP3N7PfJnb/FaVA6POX
+gw+hXpF257ZXoowTzN1baZyR/XJF9GY6K39HWI7hn/MzDZ2oP7DytfA5u1u3AHm
nRMj0h7Xe0vFFhjvggdrpg6aJUgUmshwWyVOekhXahAqLIO3GjeMMenJxMwcLCrN
ha9qQr4Dkqw6hayV/AOnneruIqJcCL2w2dtTpuoqNS0zx6ceW9n6YRN+DP7uI5ou
BzI/xVsvJjcOAOVQRnFUTFIktzIGNiBxW7aI/gDWYPErltSMpyT6I+G3uzz2aPkr
xF/lHkgQY44DfH8Fk2G2yky6wU85YZdQ49ujCJv8SkQLSnmUNUNDbBJTOTBB3r3x
QN8cS4Sgu8wV0ZPy/tAwik9CzNvmtD3pNvzm325/rkWq1WDtm5dGkRj1n3hoMhbf
8wT85KXaxP/oeASKCniwHLoStAb9G5rfbW5tf/jNVj5ztCrfRgfFWbZgEFK0yTR3
NHT3UfC13mTBpCYSPc7p1JS+ox2mKyiPwN00RpGxOukzeCIpifg/DT6crPjbYOKw
EnAaU1VpPwWqxhOExyIwKJTKZoXmKKp9AgFakM1CW+R1/kOTYpLna5kJsFYqnDr0
gURVK/q/XJWaOlw7+O05/11JCddhFBOOwly9bBRT5yvZ7hsAICfi0B8amE1KDCos
mCqJfHrhWXHhbMagwnenCrkzTIgkWm4zVNpqnSEh/lLRI4tcxw/LEKxqHzLuQQM6
O0J07kFLMQvyqtHnwIhranAHU5HE++wVfcBScjDC/J2INj2MKIeDK1XEsWgpgY6E
ZkO+7+M6NY8NvriA7kZUPU236J5b9WhnjbT8yLdo9xyt41IOPufNbLpY2s79SjUV
oAMCD6TmVoz0zmmHFok5yMK2jucDzQLg666C0NZBPvDEcc2VAkij3KKOw7P4FRNE
OhDV/kDvIjYjUxBvs406/Y3uWL3hfXdjoT3OvBe53mUyvy66rWPkMbG2sB+T9ABE
R19k0XP+mLSHcp71rPIX+eVs7RCcyUhb+Zr9qekz3J+W0stmnqhZ7qdVABU2QxYF
6QQUPf+pIlMRnQZNDof+w53qGltavdAYGS7bDnW0yvj/7G7mbw49C5pEvT61cPOj
fWIupL/KVl+VBLRXerezisDTMbAiXxtclw4+ZELwDVgRt4m7ksqy/7u++KRdPRjp
6SirwKEgm7U/hrl9GbI40uAZGt9P3jo2c/KnQyj4YsmpMFAe2xfpIwdUyrVgu95c
VGo42yexzlvB2JRXlVBZmmnqSHO64Jax5Nzh1fHutGneKmjY4YBGTjVOgaquP90Z
JWW2oion0730KiJnV3zPgD+8IQ/h5IQWi4JqTCWZ0ffqUExTRmRqmQLXql91aiDK
pwUScSdzmHjvVG7z7+sAkCKBFUWQH0rYcNgyz4hgqo8O27Xs8ruNUYNckpgS2nFK
+YgThmMIbaat9IVVfUAQZo/HzpDKqsX7f4Tzsw7pPuMHM7nkvJNrbFK64KAK4/0l
xUSyyhvAHrmVQtQVm28amYDEFHXSClLWzHeb0I8sSj94pnLSaKRdgeMxcSXDsqp1
rtjTsdzQ9/kwBlZ0oqtryBCgMYQoUKjc6EWPUp5c1ftFRR2AGtRVvJy7c89+KO8R
dpZ4NdLuHEUMqfNK7d9nt8ge5V+LG5nnK01Zu1Z0OekQAmjy9OuhIWCv6W6JTQS1
W5MmCjLHM+P5GsotGA1xor0EzmhMMaiRYR54Sqk6SJD7lUPCUdUGZBmWeGcLY+nh
SA4uC8lis3t5oeemAz4AoSoOjW+IijZUqg+d/PZxwojA2GFWYTNcgte8KqbuNHJQ
H7JfmfHYjf6SAN0FmXevLv6Slo3sF3DNRCw5l6OzkB/L5T/YoA2zQCEGc/UKnNJo
1HT73olGKTnc4sKJKT4YmhqMs9qA1srcNKGRTD3ijcpSSYFTp8t+F//bXHCTE3Ho
SW1aEeaUCDyph8E4Lu6LQ0ugMC6+lN1qhqv4OQ5G4e/PH9e3mN9X862LcRJ65MBr
n6uVO2Vt69ZK86UqgqfyoLdpJEHyFs+SPqD2TsVJgkpKZKt76XwbqLlqzqZ/yEzC
WOk/5RPnTmgPY25MuafFEieZG8OsXR7oM7UdVT2RbQD56jcBbc4GCaJOvE/LhTvM
bYnr1H8m63vzMAPZGEIlcHga1BXnOrwxK5u0RLT2he1mNfYoHOlh/ythm6z3oYxD
TAHmZBARvdT2afU5B5Tw/RdQdk5qDNL8tATwpUQLcobPJ+ZByFP2100W8otPdHsY
CWI245+hPNaUuqMHvHvsgrj56gy2dNrF0qkTK3pkTw2wlxUzVrEIaEjGif8ATmN1
EfTai9CNKLYSNeSurADFZZEfTzifFuNnRuTdgSECWpZg/ygKmGHe0P7EpmmX6nSU
SkS+vE8AdBLVe7wuWkWYQCEnbkJMwnjCSwXsNHpjMNILZttDlf0+IUiXeWExNok4
YBjny39G/x4RqKKRUTzTwnIBaqABnjgPnom0AL+nW70t9IDijAYk3q53zvp2lOpn
BycwxfxvBX1S+H20Rc8fKRiWgZgtBIQBRGNpcafl29JXeEgEuKVlAIdEoOWpVzT6
39o9E9QR3xtDjgRCradOqY57JYANZFduaLHLqUbiaDVyOzJ6c/oOkvdUN3sGuTct
evwB31rlZh5sfS8K0Go12by9yceolCV93YjgijD2RjBJNzGpSmED2iB9YMJS/f+x
7HblwO4j2kq79LMYOw6bG8lVkqf+mHlq6VPOu4+Vh3ysLNw9yapt6ZLE19r6y5nX
UlL7c3NIzV3Tt+JPEw3EB9YwneRWKIwjeO4OFF0rgGKVdf4qTkPWPhA0lcYsknPV
lBxJWIdA2OaCdxVb5d7KLmpTGWvzM/EEW4ODlakBqheCkDSgb1s3KpGLJE+9BY8E
+PleaouSI9o2AihX4EOQhWv5PCsPaP5vrz8g7PcEhVTeq8WEGOH/fEcL0cAEaK4I
0FQrffD3cu6czoR2gCIg4YoyKi1Zs8WqjBWI80tgAzwadbdiiwRyKSeOhhy9/10K
PIUwlSuzUx/pvTgdUx1ycWmf0MfE2vrPzsOdJQ9nRlo5cMRFgJB78FsgmZCo3FTU
zmZnDgAcSII0dMtY7UVZpslzARL9JbbysBYbi2PtkK2avaIKsaUZxITOlr/HtJ3H
Tzo/FMmSo0uferLb/SkYxd3/DOPNajIWKecTzY0ZIjsnlY+QSr5/9uTJTaDOapey
kVoOZHa3Ae46NfxUw50vmDUz/m1VrEK4EGEMnM67K5dotMXwbcT449rKmulwgbIc
bxPArwiU3rB8z8YjPqJzI39dz9IETZ1ihwHLFbOv1O3XJy+q8Qh0q+azCCdJYTWi
1fUR4nJZ/tg4m1jScXBWLsEXsOyw5FyVfH87/zBfH7uJzof5OXcvppC8hbp9LT2U
tO7YKn2eNk5MUxwtGDy79V9mavg7ZsgM4iTpAMwMPDSUXClKms+YQYAsg2l/pgvm
aNYXEHNzu3QAibCMR7ISfGGUmytjDi0KxnmoxG6+1v1/51thiDzuDOQuRgFaja+U
o+ZxQj91DX0rnQX9AJXrmIpka/OEjVChYdjDXSc4evY0ZwaV3hMQWAlQ3CPqazGW
gyZbcBfWXvLD2865V07zRjYyhB0ybW2I5F4F0agw9En5vxY0P/CElwgxvd0FG86l
fC8UD/M+JR+MVd7aK8iGYBJafyE0MaG7+GR+l/OKDGMv9wHG+cEnFmiTNz7bolB3
+gGbtjCRVczolENFIpYO3LT7+dPTZq06oxfOsFOu3PPcu6fffz0iB2F3BUCY3GaR
O8YKOmNW/I9XNdkxELhOUzBu7dtPacOY4Lqu9Cj5ZldZXNfH1ftIMuQiGyDHKC2D
fk/J6+LcWO8YOiZDadjkX1TTOtt2WpQO+cwRcQr8CPn9o1Hm/55YuTSWkZNv1DAi
w3Hb9b9xAJmBM3ZRaB80XGlpsLyaxdw4FrLOPfiWVM1/+H2nxzMKm+IugfH5dKCR
qYu1LMbtHoaPsmChmnoc0M+4MQF0djNEvjyxw9WCQqUczWKCDy+LsVXYgc8P+MHD
KiCbvKTYJDnZSJaLyNy5C4NlPQUmrh1rtGhn90S/rxu78IehIUVHMJMfoAUNmRjY
dnT9xSD4GQQg9+uA5x16getw/izLHPCNCwJ076brBz797aVv25jLJtOcLoIaX4OC
jJVl28FocM5YdgOY0ANvpBzKRY/9lAg/8MwoV2vzgZQGTpWSCKt/sphuhckr1kUr
hnjz2GCK0yMnzl2ktRDDa27GfrmO+DUI/yJdXgMeuEjeAjnhpF5uZ/Q5qoAdP2ew
yf3KSabzsRw1JnWiANbvOij7mEKimuTJo8oDo1lv6SUqqjHyIw5inNmxSBCfIJg2
ic9/e3L1Ryr0muGtQMWtm5F02e2rwB8U8bfIVkJPZs6a5rdmnswEbS0hyMLrDEn7
cspAzGk3hH1ORUU7e0ilxiubmXUZvAlbxoeKnPkRSr9xlpVpUmLCkC3Roo5RKYvy
XdVE8LFnMAJdCw8BFxbNkVETJP1zGrOt7YOpnqprjDU2JlS3n01HJPh8yku+yEyQ
TxjQHshAJWMAmO0pqj74zXE6Q0csARf7wpnSV3zXTVlWeaQGWhazYxnOEPDbXigg
jK5I/Ujm18MxxzLczkcmxMAOJItZZGuzsbQ09GYgAQ5bIuc57hf/orvboKLqeoiO
ERn+vK3QqSPK+wKdGRSPLDUTjNBXgYmB2Rz7jNJ278ck/FRhNjcCSCsWF2rVGJFL
fLW6AtWrPUPlQuJn+Gu+Yl6CsLV9MJgsUmcFjwTATxXSVC/WcN6SH1ZdQKnnPUMM
tuzpjtCODJ0d2rWZbr4Rm4DsMD2O9tzZVXZTiF2rMpiYmCXETIX5ngx3AyqCfWzq
9StMSAIyfuIoHbmhi/Zg0ZRn9HdFWkvG1m9e5GdV7CECM8yiUaSBxLTonzYMaxhC
p7SFrreZEclK9sIhO5vh/d164DIMQmbFMII4UTbY9S5LJ2w4KIMU8nLMKD0jIVbU
IxE3heI1d3x5TFJ1RaB2VJZICwuvRVDXxwXImyT5ggrQ51a7k3MtUyEDKMc9u2uN
BiNPP9AKtNO7EjOJrWjgh9acskbPglFfrEQ/R7Ka9YqWJrygdvfiOCEscfQw5iyX
bLlQPhBbq3C6WNYCpljsBz5vQU8ol+5chpMKo6jEnutFGYmZ8vbuu5QzVD0X8B1l
4BM5lmTFISiBWFmFGeNyf/nklRfDa3hXz5fMR2zEO8WjQQRtawQuPVPDQ5ijxEjP
9BudYsU+zloh7Y+YM49w7qFE6BjQgHzCiVPPk7yWfvHeqtGHIpx3xHBrULPfuNHN
DC5ZqSrIv73Z5oLMMnrABKjOMflrwYg67wr2NJjCDXtVdJU7am9ppJK3JT6pE9Z1
FbaPLYu+3+ajfGzX9yAuiHdqCJyjuG8I7PmPnldMvJj/Dl4WMEQl3UzuckxlUx1V
V/IW+S/1ccwooLy2ljiCNS6ohH+IYqotFVsRr6yOd1wDE5o9hsASvJf7oUALMCGP
7IHEuxOGOdv0nLRa6k4K7A0D7IU/RPHx5MX2N84v+0tci0r5zIX1t1T1Y/W0DvGN
gHsk9ujbiFmseufa0las03yTysyNWaJzbRXj0QHZCtqv8dIVM4PPbhjCspRzVWqK
qkSj5G0VlK0hEw276sfUo6NjmMvlstdHvv1zUHaY3pjNXCMlg5PBoIKB7ps77vGD
AdSz8phKrLk3+ZjquWBi2tCbqTD0OnGmmmdRRMUWbzlZgYuKwlFtU/vj6+7yZHIW
fP1NuXmqnUDP8Od7PIa3bM8cSZMGkTk3Uvbu6J+yLoYDxuUlbxmnp8fvyJKrc6uM
yEBz6KO8eOF6JfX0kDHpD3zlkDcsxxCVLjsnOqkXEiUTuQawT8sNjQnEFwXUXuOI
Xnk5ktq7BIWXOAaFUBHfMwwRdjLQ/dyG+S4i+SQYmylZZ9uOK958fBFfEL+YPsOH
ZSNsqaxh4/2ZpIffQxsJLa+1ZI5GWTjkF6FOc3+dK0Pi/QNxOEjhl5OJxVc7i0vj
Z4JMRMITOLF13XriKSFRJ25dIhbzQqKb25OUIkPB6SDCEf2X1l1kTlqu9rnLKqFH
RJsO4X6f8diOd7KIJxc9ohuGLVWYNsXaiCP61Cm+RGgw+7nyOOIfNDO78B3p2qF2
dkUHBW5LF7sCSNmgbODAhIpCIBp6p+Ah9QgFy3l6Z8wSU5YIpIeax7HCWWSktoT/
5ea5qM97oJ7cYpxUHUX166eJXdW71B4b0KwZ63sJJIUZsoR+QkW/CcXaopSCKaD9
WCVdK+stZYX6D3x6GJHJUKGHAANXHeg6g0p1k3IS826Tx4MQX1TvUvA3EWLmtfwb
eEIX55IYdgR+dwevswnrafdU/s25BQRKmT2U5VIyQrPUHOk+aO+bjurpsnfuG4XY
aFoCnvZMszlBZ7BG6vwbkQJGy4bGtV6JKvBVnSoNntkAkSkH43Hy23CtzML+EHpu
BsqK9jdLfN8o3TbaQesliN8nywBxGgwbaSKIYDN77kxkZxATlum6VYRxq50MDVyJ
pR+L1/S1BtlB1m0UV/tTn6ClH+cT+LrVVJHbxFzZcNsvTRF0yPYd5FSU7VJRtWA/
/RW1oT/JyNcQx8xxYj+8lWctRjINtQSuxq3EQgCAwR+nI+JP/esGsEKJryhClXWt
WqS12de412hELJUNuVBCztt0IPD0PVz2WYqCCBU2gGGKHSZ/Mp+8yVnNIOSGMoh3
PcSApE8gsOqjIInAySa1Hh7isYBc/8kpTA2LHweuzLHWt/E8QBI2LHDTSOZSTmex
Ue38yZYDZirJQrLExxC7dueED5Nhg/cWWTQeQOue4iFNoLsOOTjNh+R2ft7Dwl6s
K8c8sGwVzAl1dvbXE6a5rDHRYNa66UREyQEMr8ALgWWs8/x+iSb9DphcWBEZ4FTm
s7geRA471TWzsQJdigGh5xhHHqOcly9r31KHPUAMXFFw8N3KpGrAcE+dFyUyrLZr
6Dpp9P8+cM0oxZ73cPwKXNq+fro03YrZS3vW//zM/ncz08YMj6yIGKSjyblOZv11
dGspIgahgNB1+CKbsi9k4BWNoAPg4Va3BuRFkGPu8D1bF5C+U1ggyARYLIK820m0
GenBLSCZfZhX9mOnpGg3fAWqyYpXAxPurRfrbiO/6U/5rxL4HqS+FO6E2JiZIROX
KgIJbskK2ieUUaB+K8J8HxLHruM6Alh1vrRIHft9vKOOMxfCstwUizxFUlYizcQE
Tv1ssX7xKNH/zLAa47rDsWO/4owhfDoko9RfFd79KkqrOScqa76AfwClyZEJC66p
Afl9JJPVsqWJV2dkVNG0n1hapXqCH9EwG9+5GYizyvBcSkRc3zK6NnzHv2iFabPC
c7A4q68kCvKXWLn9LizLgTYtZNTZIxBSS8Mu8on9JrSRhynDUp/40g0F0r1dvTLz
O4UhGxnJYH+Px4MtlDsvXE7ZgZgedC2zs9o+MScC8j3HW4t28KIlzgHrmGKWr9Ma
UGxRXGpjrdG3UgoCY1xqEKpn2/3oJLfBELKWMULp13lOn0ldqUg8oLNuqOFc6K/w
/EE7iIc4DS1Y/aPcZStGXaQ0XoDN4G4d788c3jx05spahxxKkUYIQd07FA/0ol1R
PiqHOTFzCQQem8Fbqc9osJrx3tPHgbDt7mJGBmfnbkClxlqTA6J5s6MEWCkejbxJ
3r4V2nzEDd8oD1kqUPE25I75ScMewvuDwbU8GiFHJW1GFh90fJlkeYcmenQ3RT6d
pm2qYWSa9yglIZ7ZHIrOXlJUgkxkZjJwdEqUxR+kWHjj3PKUaHS8zkMJBFVmto6C
++9XJ4hsW9l+Ng/IxPyRP3gIMb0Y3onKpPPP+4gjTf2t5bpZESv5//uL8Es37V2V
5BSTydh6HE1saPSd1OOY4AL+Jo1WthRkhnGQEqZM8TaGZJRDIIru8wh2DJ6vxviR
x9XD8ccG6uXUVyf85x3+96BNdinai4V2H6Rfv9FzdA7TPXChVqQz38zLcpGmnqgV
NYbty2Qq1LOyaeeBay3f2RKC79OHKyNwjQzIwXHQ2BznfBp/pvkeav3mvwQHWD/i
MChm2EIUDaNJnV2ZH49LA4nrQfQHWeIY6eU2lUMY4Yq+diiA1kzV6/+mW1iAME9y
X7SDoi86U97lk6FcSOrSlL5ZGm/yp9H/l4086O9/Uw46+fgjkSWqFa3kdzFR+qXo
hA+MeBOXgtbmsNYrj1KodEEiMqSvCyyzGtRS5iXOC4x217lUt2UqnDSgDKKmAirz
rcq0wK0aVRtz1OxLuHPokkHGidyeH9L3Ee1lOtnwYPdEHwA/8KSkXsHcfvWigfAG
V9s59UHguguvgScqojfrPIdKSrTbGGKZ2csWSVZk+vzH1FAQmKqaF0Wy0b8PxmG8
U/YV8xH26breDb4rW15PQdvhqDtGtAzn7OJh3GcRb2a4oB4UVa+CyJzJy7Ai5iYK
xUW1hbRoprqveUQkA9sGt6DrgxIJ5+/22nd12uXgqfkanflf6EhxECyS+tCxuU/Z
6pmmsPUbWJ3JjVMBTsLG9fOtsDm6jDCT3ieUPHI8VcKFhzDRX49sQVjYZ9nUL5Pa
gRojkzUVogsLkyD+PDYfSNNAGM93/xvAkmJVBPHgR1mqNg6t/kLIpDqhcTUwYHuX
GvL2Euu+Yj3zAX/C4JGm/iZejyIxSz4xQOGCbaCIOOc0Gh5XzV/0v+oCChNuGvXc
JZZSzDwNwmK7Wd84BbhFltS5c1rc5rfdyQeRdoC+n5p1JhK3ov2DVH6LZKcXHgfw
DExmyjf1g26oyWOk+LTywY7haxOnjJP683WbgMrWJbK8cdBU07UtzwBJDHyQRrde
CsVcziL1F8Pyujc6xdjjFsrvc/cWiehn7Jz2FAEP9wQ1Ose5rOvRyqBncmaO5lZQ
oYwkrzi58pRtVAa1Px28ccVqk5MzhAeAtyMhN0sVL7PHIBPohz8gPuQN1o+AzNiN
1uQ4adTX0Du/O4WyO7TTVib1nLgsXkK809VUBKZSEnd4mjAmS5TuFlqhAIK9GOIs
TY5fbpOdImW1AItIwzzl/aG0xrQNW6XwJjGpk6AOYCbodqM6HLrxzb2PrXWMMU6E
/vgBkZ/1V2nqXnaL2VU7+yYVXu4ZaXrGvPj6ZMCCRbOaI5OzkTIrJAJO9rBL+9fk
aOWkKCh8NXI2bcfO3r6r/VVTmQMzdSbtrV0S9xdOI4mOI7BosMcI9yXe+MmCqnGI
fPGYHHeDZuvK1VZXRG5JQg69pZiTuzUzYt5DNt1AFjO6I2G1j4OJqohxWZodug/w
QLko/kimrZPSDNeHBV9upaGz1jgVzaYFxT/c4VWS7hhd4agirqKzMoiXC5g+YuiP
8mYBPnSNMHYKJ46ZF7xtom7KSn0ie7sERw+BwC0EFr5gV/E/x17qNjsXjih0zcy2
UcSD0xeefbmsvJKqUMaoK3tI8clpS8EuvgD43uuZCSL5o6xippZZdBhNrpiZAl39
aYSiNzcqp88S/d0P/h6eDui4BrEXHMIoC+FrjWrlNxGio8J705l523lLi+UnhDKo
JL3Ff8SN9iYBCVQZC5C+k1PLhkImMN/njN0mEX+8SEh75NQ+9kz0O/k9dcYt46rq
B8YNWouHR6upTfvKvMdAOJBM8eGcH1Pwu2KRv1hco/AYVLwK3aaL4uaGCPqefO6B
qm7QcNM2LT4IcO3TE8PJN4aastT20uvsQOWW1fMzsHeU7us7/BWxskkjcquPYFT+
BAsUrixWSlZ2/2zxv6Hatl2s4+Zu1mDk9UuE/r9InfVY9p4FKLdZkTAUMMUivaBD
FHWtZpDWGbWee5f86Yr44+lFwdYEaUMnaAa9nElmqM3oVYp4TiE3CYth4HPIKmGJ
DhubB7nE+3CYlPqrnzycemce4dmooX/q6ejp9ajxflp5wna9TcOyDW2FvKZ4p/Hj
VhEdKkkpvRZlyMvj9Nt6hiRYYNlMKzGu3Z4UKHpYme80iJvQ6OW2EyL7WalJua5M
mrxuP0JnKgaMIgafDr6ws9AKUnVea5YnGa8mcglErbnPcK0at4dFj/EH+/GMO+E8
UVK062MQrjX9qyPWVJ89MYty8DlgD2fux6gULtR61Fyx79/G64fKdVgZx30KESCZ
hs/BctMVjtQLrgPSQcCXIQA9FL92cj/mnpuUENiEP50R13YByZaJdwQx9d6MHxui
LR7OMhse6bM5AD3NaHDJiHEi36JC1qZGP4eI5OcmcKD8Az6mneyXrBtDL4IWBQ94
PAdEplCvMKAWMSzFt+1xv3YwjLjQ9oL8eN7MPBHi5SgaPhSERdqecXGJCGqMwehy
N006clxq4k5TCm8XygQ13Xgwwifg3ovq7y4hFR2SLHohfn9smH6HcJPM54MLAeML
ZL7SGfYe6NOs4gThhdCU0+HCNJcuyg7OUusMWxlTS9S+B6naNgYnRDh98U/En+Nf
f9FVkdrwy4SUpSbFb0uFLXTdg+c3hrvjSg41ZsRCL0t3S1L3isRvcNqf1KIRqfV0
6iBGwtWiDN18ST+xFvm3hBZUZ8WN7smFdy7i8KJaqqhRdFae616dpvtYsqRgnOl7
gAtAl4rVtke94FarKktW/j1O2oMrksk/sXquIXg5YMOuQb8dVnToRaqcdI+hj9+G
Ls+djqwVmJxgP8d+toRj3DaF1Idu1KEUZM7W6o+LqWeqaZi5HpbY9z0yj38q9lTv
cch/awTDNFatWwRBMreQlzbfZZWsgABO5nxSPYCoeU4vVD9dqqOJdGPQUque15jJ
PxPO0Ml6Ukl5FLuiMkjkigLXQz0CLibMHHZcDuN85vsct1M8Dd1EYpZouYeQcA6P
U54qohNn7NAtyaOZWIF/IZQ/U7Txt9dyft8rg8lz60UvRfjR+hOTT1PWDhl5mm1j
BEa4T7+elaLwEw+5ckqZFgWqXhrbYs9agO6LlNWyA4wnTNwidYy5v4HyPukIyIUf
+oTmCaS3ge5S2o1Cz7lv5lu6GhcekZpKPj2sHqtOAUDDQTkV8FFKT0l7Wtg7SEaG
bIBNaXVlLm6Ev7L7PPjnqb2yKxlWBBGfR28a6rqEqD02iZRTyOieVT1kAq7YyKzG
UpUT0MlicJf/HQ7nwTtdLZ9Xhmbl+46hBpB5D8/Av80lMALCqoDvD5RQbmUcJq/n
/VEikJje6vCsTOes029mu9ze/T/EGU4RcRvKBNqnlT+KxCoO9D5fSYQUTbu0uBqE
paMj9ptWQd96kAXoMwUXAl+AseIWmoxrr/3n+BWLs2ocnF+hi1Qg+LURvVDPZfYY
6Ev3h1x6uY1mwIQUlByK0/8KPIGn8wU/LeycYHTnmoEkmF9PMaHF+UID+esm2F9U
rSR5zLJACbyhEzNWjtNAjyg63Rz0QPcngIaWMcly7sw4W5T6t/kTx/+xgPmZGOF0
d/Y+tKbuu0+UV3gLt1xhMRjfazFK0yMrijaZ+t9wlHUPIcFBmBr5tqHwBiY3WE19
WcS+5geCKbYKzU3JpLE1cUcgHePDVoe5k9SFvANAjpfjyvUXG832bS3xKBVX/0A2
4td0/PCD0L73jGTjX20wE/Z3k1X9s94JvKGPpTEuHqXevlkMst3tUtgtbd/7uSxz
2vY3sK14lyItY9zFjpUV17QXR7qZf5JCgEWkAySaoWt8ByORL9V5qBEcS8C6/bGC
fq/Yu4kln4eLOxZGxJkVVlvvhSmfMoZdqqh9o6JP4+kWRss04FRmHwL2W0c6+NK2
03TSAPrjytvJ/B+Lz92iNgsJ0rBPnGsIR04slqy4vuOdDw5mrfHunoEYHsqyVJvW
gtc7kzlntFo0kvKIxItDq2AmhLQ9KhrzEBexof5q/85ryedKm7XL98lPd3yUq/8l
f1JThkq4iWlqFWsaEN54pavXvmoWfLoxnMViUjtBt7EDHHYlMPamu2T+NScdjYPm
lw3yKVYRuaYzU4wYr6wIfbvWwpzFoDpShC95iLqW/9rVs8KBX65YYv7rrx2PguSu
VyNtLHDF2/p9bVu7VkUCF8U0lA1ioTnw8wfBziAEQ1qp1qJvY2IfUPiLY0DcoNQF
jCx9HBHBkwSVXPpdWoJBxb0YaB1zK2xkrgPJLgOntc/STNZUd+l7gkz7H8m1gXqz
R3PA7/n1HjOocmCO+MYLwW3ltr+l4w7nmseK8vaGEIfME3CQT0dBazDeKY0ofeAa
pwcT2tKTwNP4mM5fVjrJEc+rg2qRg3qBcLoMNTEukzTUmQ5EiYZsDane6edj5hrY
96ZGi0vGvhvT1nvCzktxTfBPXbe+P4W1h6n8hOr+aMc6+Ww1Z8JosTlWVaAKQ2Yh
BR1hLQIs0RT/R+cn4e4I+YaIk8pWxzWiDy+Ctw5enzmdID7YCYg5IO5IRXODmCSm
tD8Sf30chyKkaeVDcrhf8O/ggB9BCb+QMCU+RtE+NipnDt0a57k/bZVC4Ank+Wt/
6oRnmct2/ArvqV44LTMX8cAGyTkrzDuMlvsBU9UwEIJXC7YkeDKuDpWI4ueBt3/n
AXI3mQ855fUBcnVDYkMITr1tDxErdxl6k18YQuY6f/Nmbo5LSncsPjUePSbvGT1Z
xmkNzj7XKCUZIecC8hDARYKMkmTMivplYa4fnlTs3rrC6K33AuBqPWJ+u24MIVaV
ZsD3G54mG37OAZC4qKRUYCh8XhyFw0qApCQ+lWO48lZnjab/LSONyELJfULCjk5D
i6jzjy/xs8QB+/qhUdgaODbiveDfydMHbX12p+RPw0MP8FI3WcMy+fsuTFDhBMmA
/N0LAXurmub6maS0j+9ITXITsb8eBhjpEu+Gf8Y3CZjqrPVFIrUzsIZp5QQdSwaP
Y74CQOlf5Y1K32TQ/Ua8faF4fhz+I02Du+iIwULZRgClSsPJJfDEpmzt8Ycf6Enf
Zqu8VDXVpuJSISniBjs/bj211fH7w5uRNEIQT+EwF42abRizW2KDT4SmdvI+bh7e
iAGvU4wIFvNPjZXDp6w3hwWUpSpjqiaGO65462weouNiI/mM/u0+pdhWzAqNfEEb
kW6eRU6vMxSeNAnGKk28dTS3QZgFaMoN3CJqGWg1ebep6b2lumWsJ/iK/udQ/6gr
VIVk7W2Dx1eiTSHk50sd9hJ8KJZhoJEz4o1EnPHd5G6h9fD8LQiaXjBT3gR2bYBU
2wUYHOT9f20wd6K8r9PZPa042YPNIBBJF2aigpwdL1Wzs/amPV2W754lXljNk8fR
N2G4GJusKGhCcE5VtLqmQR/B3YR1N3kbWw2bQ72faKQ9MU73QV+7CkC1Z1/dQRmj
vLQadX34naUIcwt6R1e6bA/Rendt0dt+H7LpfK74DtaHyxkjZSMRtWMbkg/aqBbP
C+vZT/NgiSXvnNclIe/IRegBTSQxOrM2RPQtR10tlVIhbnUWSZLxlrIaBe8Wlun4
ErDEfYnATLoiMerAVhEkyfFlxXCD43m2QXIaFR60YBAA+R1xMP1/Dv7pecxnLd6k
YO+5ihi9rNBn41WpuOzxN7BTC9M+A5EKAY9rz/nIkHnoAmrmjx945GnELQhhc/7D
8+a0UVK22fuEIC1RN2K3gdl97dwDCBTi7xkp2vjtNTyZZgMaT9rfgUKj9yl7xg5X
fL9SXp2eTRpSMiuPTg6q5U3n+td7gyXNQAzmawLULgQvIwsAlMMSR8DBS74mxo+p
EkdvKEPgYNRlV5UpKKIgnQJWrw/awaGoU2LBILaeO+TvZKSP4llBNiPMZrlFgf/n
/VrHmAHdpMw7bXwaIt+dCwFXBxLIQkhVfIfMrnnHgMc5AjRoBy0lwSN4EBtUbaPb
n9XXfXAqF4ezfyZE6dpjDxRxh1f2VTiFeETcIep9HcwSUZ4wacX6At5ZWXbHAZil
NxtxIboYSgsFcxbRSkbly2QFqvuwwBCdYmKSSHAHrn0R+7c//rg78V2zA14+P5TZ
siWEOovz6Ps9tgjnIaYRuOuAuZ+P+xOBWqIASrEReH/vlu9aPOG/o8hxeCEd3wlk
tV2Dyv4GtdObhaljtE4Q5vbnnV9aoIlHszQAm5CtNYyBnSRM6TCGTikbDwjG5Pz3
Gg3w/yeO1xhhgYiNQuu+Mx56N3DaHvv/kjD+4gvtcIKq7DU34gE/EaPCtriQc43W
N5Vz+4h9UgaQ/nLN4CucUcuLNtu2oh2ejrutQBghLLWnJ2kqNgWZWw+R9+0HCPyK
1QGESjehhPL7v1mS1FdTbx2avVNkKzA7DteBHE/yaHIw1P2x3YY9hLLww8q/iBjT
tC+OYDOKmwijd593mQ1++sULm0BVKAc54GlO1nKl80Dj43U6hWAk32wLvhs57Gep
cqxOfDN5bQx99d4/QJrvyFRf8vY9tpV03LWY2jX6zk+0KtEPJuqItoQP/osgFOJU
hOXLOL+Xe9ucBGSbMrOACiaoyxPdZbQIxovrpZJKB578w97f+8LXGEeZ6IM/VxUH
HnLcOYFP5MOFtdVwv0JI9JkNmQYy9OW7c7JoCSFgXJPm9hcirQ/mh3WqCvoktgkN
7r8EyNUVPyV6qfYBL6ia9rVujQ1KaF40LH1uhl5FNxHyg9JuwMei6BOFdpe43qFr
dSNpQ8wrjz1AJRjNLtPmlotLeVRJ85/Hz7rqWS62aaprVfo5gOHwQU5x+tIOxBzD
4haWlJF44VLYi7ELiVtrvbgS3ZzeDmtBkReRIDQogn+vWBzxmkuqbkVxoZRo2rwv
e+YxYsoVZ1lu2of2wUSPBSSwA/JwphcmC7eEmUAbjtK42N1Z98EE6PewXyLoxZMC
TmLPIXP1tn4U/JJjImtlV84qPi/RCrrgITuGXgL1xPJbbJttmg0aFCaJlYXMMfuT
8Wd4IarQ3n2ayynM7D43KgK8R34a67j2i9IQYV0ljnswIKCl4DbnSHV2eOWuQdVP
8G5Je/DemqwbcY42JZquFqnG3fNdE/NZ2JwvyrUBy46r/S+umztN5MqhGyRbmxjj
f72r/EChF4xkCCDXSSsdL0z/aIFWSaFggeGsi+iSOmrx2Fjbim7mvjun7dnn+0Qo
s0sQmCYUXC8NcF/8o68CzWb3tORphk5pIcUYBGsA+9EThbVPqdwm+QO+4CwzFqJO
M04qe37aLKetwG+0Rc5dO18N7ck+zsrCM8qkDKaMeY95CuqGutf0OuqLksoPwHY8
fTo9AVSJmODFzis6z2SrFyWN0m8XXZ0zEr8UpLeTeHQS+p9kB67zFdYp+flcB8gB
4kv+AACX0wd4snuaufDu6HDXNoWnBHt1ZB0ffSVikugjyzfSYyPiruVeAvhSccbm
XMqj/uemYqMjLvOdVZXfaV4gmu6pSnHm/x44/ohWzP2x2ErAESC6+sYTWKS9ODK4
eUxqL9sb1+b/nEoh6anuvD12aQ29hJ6NhRJqeN1YTIVNmiKh42tQYrqHNKPTL5aA
0xPVDZc3ZkEauz4dfXqTNlyDFM0Nz8axniSBLZcvIbRR1GowMk4rCRhRASu4gzTG
9jldfWnfXFjuRv37ev2jJz+pDwUFIT1PilxlcKKT9in2rKire2UDVwIP7f4omMM5
AqNm7IUy19ELLI0HfJSjfgx2aibbLxfl3M4Fm+tjiCwoY4nKgm+2lw4aTZrqqF0d
t1lfz60LC3n87AxLXKxUyXu+erkZbJr9NwAVeshz6aCIWRbL28G9iaUeHObMWcU3
Ls8ZL2Pt7CaPjGqbmc+IAHSPffyh/cel/KEHlwpm4/vCANYpkW9ZEuL2uXO1k4r1
DygaCGqEfr+Ieu6g3n1/GT6LqpXG/YNRSxOcBif7fvmNgzqL5+REUgvPWHwvgcBL
JkYQzTqRZe/1t+MkTNg0uggFCkb0miHI0pHV2B7Gmb9QyVV8tQwnlb8AVB4ygYGU
eHkuQMkU8woKqff8aW/BJ/ClsUOt0V/5Ub0TKMFjpG+Ilwm47aapzWbAMQUGPjT5
cqaosB0n/YNHzVNHMvgFglfdnmzoRxPHpH6Rl0H/M0ALwdO9pq6INP61CMFzswnY
GxYPL6UPG1RlzxE1zouG9JdMGjqQ1iwZQev+c0+M/By3l4Q0pBa4Hlv9SNdziTGV
Fgw+AIqsI+wYB7GC6Wh3WMPfVKitl97pG/zmJxPKvpfec5uiSw/qL9BOVY2DwoUY
suzzDKDdmAzA99MSP32cH/WuBJdxng9QuumZhIzWwpO7oBudoM8plrAgGpg81FgA
g4M8FRpwSJblHAvSq8UJfxUUgeWtxQmI9nAxqtElKp3Cj+LubyqmbdsbDbd3RPTH
mBdoxVP67ZO+uqdS6F+ZmA3uohjoEfBdXIoEcnvDKJYfb+V2YWcqk9a0kq0oHQqy
n4uo78TQ/G7p2/NxRfoJ59bAFAhu25W5Z4MEsUIn/vAJdLzmM4IwxmOdkrBk63ZR
hqfgt4AiVPrX/rs0ADO/Q9logaDH/g+fedA8waduKR+b++G1ZZcHKEYfzMw6SpTs
7OUQXMAksQBzOfyrYHeaLYIy79hEzeK36perq4pXj7U9vDbbobmOnT5zyuO9cEHM
Y0nXU/R3poTBL32+ptQOPrPzHYhAdusaUcnoxgU9xlzCZa/4aoGTpwyeIJEjfj8g
Ix5SlSwvT5hbwk2EnlhSU02El1ENGpCOsrG371mNBFoCDfK7U2jFMkawdCNvttWl
acFDRyvhEiNkye2kwLZKExzbQ5T4LK/jP35ZX/i+ZZmZXW2RuSy3TiZSWNnAwa4A
XHGL9rGD2+Eix47UxgZCiRhOiTsSAc/GVC42qcY82aEn5wzspIICp1JT7zRBOLx8
p8GaRqy08Eifmo1e8pDnrgmHtRkKQwSwS1b5CgGfjI+cnpGZj471NxSvTsSQiApe
4UblKzaSkta2Kf0YwFIaDGpx7Qm0IGOZRPelnyC2ocgi9hQ0Joyp+H0tHmRdzlxq
MYwjDNS9Qcdsy1EwQLRz3lRHM33eVh13V2hu3lzXHfoxg44mkxvSHkbudIQAfCZQ
fQl7y+kbgXegngnHi0ALw/RTVxTS37Z0MFATaIYF75TOi5cA4neRfi7TVSOWk8Hq
ycBqpBgqhbgiFis07wyJ0o1qt9xzFltuisleATdXJgkxYREKP0qMCrC62sDVwNKB
fc3AcQJ9SzZKBDqCL2I7UEefYiAfqZSLb4fA98gcCQ0J+Z6/AUTTuAzC93DNF9mk
CB3adrsrJLdz57tD8C/FmcLiYEp6INArv7Auu+xoGiuJXTJjbi++DIDhVVRuWAet
G/4LKk6Gq+0EFoi0+9HLwYJsATxl9BA24sOko2nw1fhmlscCsuL0U8hdnODfOJ7D
N6tNydIXSoL7e69SSFKg6j3VFBLgyz023efqA5D44fdjbwhKVBGKPJ/pHeiGmPTn
sIUyOUVE3mW2PIWLvYxa/MyIG62MaBigk29EO0h0FrXmoMd2Sjx9irrZmI2g8jee
OdApOwKcUW3dOf15+qhfxif7PjgiKlV3gRR7QxNKKykrruBjfoFlJxmjYiiBQ1tz
Jkesf0CfoXtd7mb8GvVlhgImI88ZV1HtlehjLC/s/VqAAAets/CNmcURlkjbl3AL
df9wCHl3llRORHp5wGpKl9TykbbgvXi9NAjFP3j09UpFOSLTeSEYmuSKjhk/b+O6
ycOlyctGLjc5vg08/uzDwhMBxMNE7vUJG/N6ZonY7kfxpoOskuzKMarOuvyxAhJo
5HC/T2vWP81sqSHEGV4dp3VqGaYL23GdvJ9yrU/y3IwJzQfydlje/yDc5+oVCkK7
58JmJ7hfO6snHybqzDAbizkkXgBQY+jPdDNQbfhAuAYuaXYTwAE6f+8NouEw0vb0
lOS/ztXWCrv6a2hyWt4F6LcQYATuk0WvY/O4MTzsQU4SieA4k5wGKnqbmXovyq36
yu+BS8IAXHzae56AUTr8ey/emLncxZ2+4w5DZpbAGUSKdFxNk7XjPzMugMaFW+2+
HOv5ngjZ+r7H28sMkotQa/AbhHUMaHc/UZ7RXYRk2NaF2AIDSQtyBqPASWvR4aHC
Af2wcxLd6LtkCjgaTZ7hRBcuq2k+3qU1Z18HdkUDU02IEG2cgvoz7Zl5bE58JEuu
77feru/Raf4XQwSpZpO16Nb+aRK/n0OYjM1EpXzDCYlXuSRtKxut0YOixuYtt+Ls
fmVJR6DIW2jeT18GC+PBBBoH8UEquX9ZxoYlRkMFuGoUw86LITNSIW4e42VS66aZ
alQPpdm+JDYrXSNZYT4Sfr/wrAFRP89PMONNIWhYf+PTjjO0CpJLbXF+Tyx1eoyz
5BZpMKIl/2jZGUsZDK3McpkY7hA5wjSYuof+U+uIt8WD2piEMLfLfZZ3/WCig3hQ
EIWOZEgww8qZ0KMrx3gkuzIMS6PP0LQDEHH9epH3V4tvncggjzlQ5NVp+YEFjFay
PSSFVfPleU42EOupGd+mpLfsLOsmrT97krO0lnjmQZIhcIJ11AzCE68vpZlmwvCE
ZyCUpPw88zPfz0wCz5l1dRalp16xKg3BNg02H7XjZInbjczGmUKCk7Lvp2H5OdVA
BxoUMi5qtu3gwYE1vtF0E7bFRtiSs+FAR+T4DxiDBIwR4H9vLU+mmaTP9iJRovlr
hlAgiP3SO3aQqzYfEqg/Pt/9nEMiGXXozvLS4WPilQfsf8rOT/AoB93Fp41YEIqn
gUVjCV10R2V6vlSoGkYSSk9UjU8ULpQNm5n/GKcdw+tXDOldXlJdUNNfY/ga/ZSX
y4YjhZJWVpAst+eT+qyIduN529oZf1TXMWWuvBUuNBUeTpS9SXa7obw7xpy6fr3l
0li/C/ICG2PJ7mPG1IM/Hq4ZF0NooX0TJN77hH0p/xbShTZPU7mEhhuV7ilvH6So
gHgwajc5GqvgWvR8kqbtdUJRCvQmFqkK1W8FFiAq2rwxq3kd8Z+VYRXV8+dLjC8g
AOwDUanHE9FE3ZAQO7INwO9Ux6OD/3SjhBlyGxCwjuCS6MRv9Tv08QboOUr5f2as
8Rjf0nhI3QK2HO2oVbOx9I5Cg5hCysinSWv8QcT2sHL3zo/yQabu4/8lmenGQxYx
C5dqnPNwtEHQE/25Xc3KE3UACxCsom6p5RArx0En3kMNnogLBTLnI2ss4CChWuy1
JHL0oDYn76/jhyfsAvCNH+lgjI1JHbNxOo7tkcywwSbuN0s0KXc7jYq+MS/olMFe
tR24BQYDT/CpzS820eYmZjhESbdZKvJ2QkGcrU/NO1nDlJqqW7yZA4q9AsCrerDA
LmeLimFOaBH4wQmNaxwa4dgz032rAL7a2H2ND90jbia0HNtr8Z0wcETuF6JtaCPu
yiobOoj+zAxqx2f/6ffEFmZwp4rs4uSF+DAE0xoJJQiv7KW45TuG7Ow0zCLxl/oJ
60upTozC4rPC6Qd5FcJ/oKPDe/9t4Jb/3+DJjk5vfl810/59rGCcQXtX+fSm7Sn2
wdH/nDGfIhigpskAAHzo6lmtFylPTAUAfbbf+iEva+ohO9vpAZHKGLriZnadz3xI
uajDY1+GxTa3ByYmhSDdPTM/F7FbdTQPoYfKcj6+xammnjF0FQ/V6XvRXXEbKHYs
oecz2STUYXaNDH3tt4yGFHRRpLGSZUat2TopkMWtHAyZtwWzG9kkAAfvck3CL0Yc
kcdHJGYAShyxS/aaceu1PIctRzTgqHinTloFP7/Mfeu8zFPB14S1HKAB9ytaEaK2
nGfpAtwjBedBWvEhzFOiykPMMRdDfH6TQI1sPB9U8qvqirRgq8TcsReopcfxeYeg
SaNIt8H5sr5KH5k/oP4MvCDG1w8Ego2UvihY1miE2TYDDRoxJ4xYT+8ZgMIc0cdV
Ds5qB3PZlrjunfYy7ThGf7bPMc4pHo0GOSk36paaAO7OKEVnRQiPycV/T0TFv72J
hYUR2IN0IZXl1wJFkNbjevU0B5TC4XdCKL6KMaDZPdyUdrmSrBt8C4wrWZKy8J1c
cp/PJ4YFsBiNGILZp265hn9IVMSRGbl3dEUBhKY284KHSUtK1QOQ2cSSvJ7dQxyv
hl7dkTf7go17eDv+vHZCE+WC1S1NuKv04jOVcg9ahRSMzSg/to1ry7jt/yiB6pFS
0vF9Zqzs1QjY7ZcNZJU3eBvy7tq+I0V22zdVx9PvDfc1hRvAXI15lobkFYE+uUqG
KuqEtk2ntskQqrl3KRH48mnI+ntDpBPNB7juKjEpxWjLpa0h+GKbY7kKB8HDURBW
aauD+UQB3Kp20egYQQ2IJBichXA4lqFipfqQvtT8MAVnwQHPijY7S/XOokGn8zEj
qys6MnOmdOduEBdf+Ypj7CtSUPoL4ZTCsrdr1STnfTvLeQBeHESfNCHbrFJfdK2T
sx6rH6TvYHdBrd7ddJr8TxFhBtDhQENG4bwsDkn1YzvklKMrbZYYWu+9uMXOpSvq
/q0WhOoP9SfQHTyHmUgBBUxcNqxK6z6x1ocfYJRJFgYG4WnEWBkDimGUT5ZkIvF/
ZQKQnX1EOOVA5W5kaJnPbADp/ifMvhm4SRyYAkAsu9q2e0cxY/kJK6vVApdMJDV0
h1sVBpyvmaJSCTSKSnqjleIWUTIHjjKsipcUtyVcTqG7E3MV6Kdfsd6MWZ/DPuZr
w/fi342+kYZL9vKl8aJS8hWdgwGVVxVvn04KM8VoKPcpj2Z85BBFK9yxVQsoXJ5D
Wo28ACgWU9vH1csU4lNp21UQ0knYVpZyQAZT4S/dBUoS3CxijLctdS7E4yog5ybp
qNaMK2TasXFauFTCe+pmyiLA/lc5yJfTqvdogBHzUwVdvNHdYuQcN8n+pEbSWQwi
7W9gMw4cF456QSz0htI6M5aH7P3ex8UTpYI9MM0j+CvbNY7TZd8KaP3rjv5aN+FA
lMl1BoASz46wzram+916q1ELRU3Nb2uq4LnH5E0S7qCiuvLg9wm1MjXd12PzNROq
i5GLlnfwc97eSOOzD7By3vkstxUg4xofxW026PjcqkwWNRjGyaZvhZmv6i//IiLH
fLD3te6Dmt1wiWnlhicpUEQl0iOJXc21ST0Haqqypy/D/J/K6/WcJIsX+PSnNhJU
YyV31MFsrBrAZfMe6kXbEw/VRKw3N+5kXxuw1DKCFs3LHiP2Afjo/OX3Q1M3B8L1
KA1pD0BwwSoifA6a1J1GUeqwH3Wld/WwbHFFHmZVYUTt5GqEu6WxNYvlTcJOSn7O
NPt8Jmc8FCgKPFF6AoGq/Oq4D2AAo0JAStEX/JVxZ0NiwQTOJTwS56mDKQzjtXLX
79946VZu8JVHiaZX5VJSDa9AVfSFMRRbRw1pTu/PV8UNoDM8S9pBa3yIa71Iz6Fa
JKkrRA3CflAggvz549M6iz053y0cY1IeqqVFQXXL3miOa3vszoDrfAIV8P7fapg3
mt7B2YLUCGMDUIdRZAcrn7zKz9lonyTqPmusJedfdSmDk1T4PwXoTR/ej1dYA7PF
HNyGQxZ5afZeg/oiANlIY4N0adI8Qaf6Fu6o/IFMgpX5knJEsvvi2wG7uF1fJ1oa
d97GnTCM0VZ3Q7fFKpntqUCUuBB5jlnybAZay+c+MWPPTo46Uk6pafN3sxE7Hnbg
84v64QeCQOn5lRVwy2isQHuJ1B2Efpngqe9hUeiHD4muEVZAiD2Q9b3Pv63rgJIC
pCHC/Djv54XCpcZpaNUiZL5WEOt/V0hSnq1p9EtAhgocFq7wWvdpyvFMktLjqkel
JoNbfJqsgIMWwjC1iwBqDJO8rp8uBST2W1wu+SZxH4wVnhdZjbO3n3XXo64O0Mts
5Sn60gs0dgIN2QrDR7uFzMFjk7pPCuyjvRxIQeLc7VZmsa50Bi7qppJwva4sfKC8
nZEiuY2JYgp6ouGdbvrpd0m6g7WySnmRdx2R7bnoqdxvwoPUQJNxh0ij0HepbHxI
z3DfSb/Vq05Knq8//a1xNYJfYSZgZmkiQHkwbOmumGBk4+hv0D3F9DDxmUiFBc+W
2JDZZ1EK3N0rRWKrW2AxUVBRIPPncaoVvWeh+mARxxoFB4/jJyByvsoue+NlWpdp
vF+Axd1UVDS+WPofBg9C5KP0kOyZlUjOmdqv80RQWPvu4avoWIZ86bJ4CVFIoI29
ttQ88o8SKCKM+zHLd02MGBpik3DZzcwekzh7rYIbbKaWJf9UUJOvvHI7uvB2RU/R
6NBJuJhsvZSRoV8GAEgPFgt9Y3ExtwgjTtpnbD9VU22cSPrl91FgUkiPtTGZyb3j
YPO6jqHCFgOT4lZvRhcT4Lh3akja7wrNJfGtRZMmxPPdwci0LKsJ+3tnFtjAd4iJ
yLa1vjzvqaLtimNESlGInhLj2aYUIcgsuT7OgN/nkkPFn+mhGqWOm6pqvgbpUKSe
e2aD0MKF5/zhhNfJyxv1GOFnYNSCMUFiqPg8MZFHPx1kBpbTAS+2ilS+X18aoDBY
hywaS/RZVVxU2ya+qhwVGHHsrEcslq7MttSlMINsv+vG8u27mLlXledUc0WX0kZm
TR9BZHdKj8Lf5Gk9gntPogKdmZecOccyisb9BljTDPYSTdr+gqjojyH5tagWxoVJ
p8kbuziZXeKTjgQMPJ+g3mGqd91pKj8D4CL98fJqqdjYt2muQMZglPx8WSxUD1Iv
+sjW7M6LzPQ15bEkI11kKl6REKwWs7JqGZIvB0nWMvn4PLhKYUbP5HjrubE2YLnH
hNKHPRbKJymnPdE68kQAgvgKt/eH3yZOACml6HPkqio76O1FsRzDJViNs7qwPk+x
MZBp+Jw7qz9DtlDnivCDJOjw71AeMGfms+HnmOiY8WzPopzUgmuYzu/afFmuMojt
LFe64FepGI7yTNN9UnM+d3gY5FrhE/P+d4Vfom0O7Psb1xU4CAUsC42sn9PU9iKs
E/12JZ4oXzv5YevpG7XRw6b6+KBMvVto+G0WEI4x+TYIktbitDYn345u/DY4LYLT
Hsef1dbBpA+VbVS2QepYx9DQKHo3bq879eWiuITqeMGRSx04/3NCjv50xR3hgVuO
98ee7PzywPYV9+yWbupzC/FT8BoQyTKZLKuQCuU2l4lUFvvVK0uiqmyG3rM/bFm8
WsUGy9qBHM8YaJu9F/xiYNWgpRTdZgQQlZhSWrwKMJ0k3BaSEraZjp/n+aZGO/fz
LSTO/JsdcdkGB+gi3Mo37kSoOmn/x18gF3VrdDDwKladnGwWe0zmCACV6fhojtCJ
Ky2+PdQhwsS+cR2l8QcUW+IP074ZYUAFEdxqpWjxKiv21S/Z/GhU0157IUJDvmTb
2Ar9XFCNkBESsyCLGeWKGkjZRYh6S65H3BA0HKYAciY6OiclX2SqTLh9quyg0CbX
JYVDnc5nEy2m58ezp0slc/LrNaukaPQHszspymgewWYCsZlKim5lOmBjcfvZqAgO
zRX5JkA7MIao6VcfH14sLbYqDomvDJr1TH2DeQWvroHYmCHTx7cofhmnpUNgRoaM
5fAA+hPNowNJhV+mAXo55JS41i4sGpN9WLHJ6+fS0hu1sWwFB1rFomp85OwTLxGD
c4sTibvBwGPu9K4uDl4wwFu8D3XePLpjnIpmV4M1Qlq3PPwy05nnxL3boj2ceX5q
HgjWLV+VTKBOMETgRJwJ1gFW9AtDzF0mwuXCeXQbvtquXv84OtRrF7tQv6T9S6RM
ksrhxdplsPue1A/yKmudjKG9ITSj5oTBgpP0rvDanmkmadau+gSia5RnHYCKu+TS
HFLab5BSEsRR/kGD4tIi1eSAAz22CX7ygXmxf/3QvSYXOGIEQLt9S0X9iLTbsAx0
6u14uvml2ZO1bUWZiFZPI3lTDFGJttogTH69JXIGxCMjYlUyV7ac6fvvFkaobEQn
AsTgG3maG3Fuin+hodpPSMJt5rlyRZWxwJzSFRO0sy52JJXpCfbt5dHV6LXk6v2T
EbPodtb3PbAXu9+BeROkKw7w4vJOjEh6lxIFIjE5T9HU3IgTmg8x+Qnbk2q2yEXF
FSs5kdPJO628hL+65HIRS+/vZqJVg/R8XCqWFbZWz2RbE4dMXTUrryT+qQYuLhTf
qX+ec3luyACg4qTxOo7GEBbxKLnXIv3fXvvdaI9iM1mLx9SbPXSznc8zm2as5rDH
OTyXq/LgpFwRVHU5rlFt0xjcS/R2rDysK9wEZY/BfL0qj9ObvHCCw8kORW6Ex/fb
np5EQ+ahiEkEgfsU6vbVmHFjSyXlBvHVq0Z4VOkpoKlg1b/j+6M4VIq4sbUlRMzx
SJIHWvFmsf5kN9HSHZaA3KP9eaoW42p+qBQu1veUUDTCBt8DE03gYc/s+KxchVbR
dB4p50o4LjKm7uxRoVAP8IMkRcoNh3K/f2xeHZobBHqQeyZK2vixN+6hYt5wrzCx
ih5BiOgTQd4K1uN2Gjqgff8OSViAYdqJShyL08Xfh+6UYOKWblXx06WTnzERr53/
lprLz6r0DobVYyTflENh3IPN2yIM4nVK8mQvCXs5+9WM4M2JgvH0jNfVorBgufYF
bT63vqsHUCVeI8nILLghH5FCfbNkhEKfqd5ex7ZUCpc5fJY+soKmPhoMPQXvH1qs
GZTkqTbpK3Rb3R9wWZ0OB7gKwwdB/nzaPwwS9vE9r3nlRaqryyi17zjJQbMLRE0z
r8Y9Vq/QNV1CLz5MdRtRThmrjKgomKWfVd4CTlyV3Vgunet6q6gRRAy4JhMS/t2h
DslVJzFGocfY9Y/en+mAwkDj3zVtAl787xZ25VrybyR3U7bzLTReD9oinnDm73js
u0z57W9iGNJ5EeXM5+1rQK3X8fCLeALUtB3iWDKkn6emo+LNnavVr9TnR4knAPir
z6bHQydljZq3e0Kbl4KOJNgiCVQy3Qqkk6jEtqxJv52NAV2EdGwH8H+MfXblSvdm
uH2MRyx4WO7WLm3y20iGKNprSkHACUoaPz5rIZPdFXGVeIzo1UZDRuKwe4raUA8M
RLZdPzqBmGD25xoCcpm7GGKzabYZ9e+RWjZdL9MH4l85fUeX/j7wKxnSPKdhrjPf
s7lc/SoYw+mClnmHueGq4kTqIpxxHl5tZBJG7JV4j8woEqXsKZ8W2mCN8SLDZ3+T
QElDpe1uvKBDPuzihQoiyfu9DALlhngq3AKNt0jLIbpOFwsRKegV5kvQQIjygDtV
jS5OAHGtgmcapXzzehx5o4gGvZjqmq59nbXliUQOY5T543+/2rd2uTlgLPCuJD4i
gZPGqvyeowjO9ScY64uh9uGPRZMuOPj0N4cURZc6ejsc5n3EHMRYS1mXx9TPjgq5
3N75ohveWv9AjFADShoVvyUfHPlFtlmI9Xe8P4VEDqMuFxa5T0vj4m+Fo1WATIGe
ygp1AEuVY/aK4xGoA0sdRs4BVPgZI0++W2cpbh/IO5bmvLwtTali6iqPs7cCtbB4
f/+1YYFcU2aJ/nft06EccMMM112XRgSrC9SRwjDLIN9bi+z9j5LdLHbbuw5sZtaB
Iq/KQHOYr6JiBphPnmbc2RS5EfjO+cxqfNmg4qr9g3hwh+cSozkYKcJObh9VYWQ3
DzE0XXHV1h9HzNQrsOSD0WQhbI/QjjqZHBw0ETe1P6DMA0OBp/2cnccFYNpNf9yx
zwSBBtlZ6PSYgJl+2MXDOvkO9JHQZbsNcQCM2AzTUSOKhHtocrLvhoEfPeF1A7u4
PJu0uKKXmVxe1fClZwlWzZckZWsDqPXyoTjH+tRek0LngHeLOSxsPuHRF+fU8zl+
kdx+EBhzF189SdzORKqLUyagKtMSUJV7jGherEukbEhZzRC3EigYv7fTARd0Gq0f
rAvjp8CxgHkpH54q/Ouu2sFkVcAYZjvenYezNI/bg0+bFKFNX/fIv8zqCFZTDRYE
TmeDtgUv5u75VW8i2pwCu25jeDV5SVmY2krzXkYCqZ/S3MafkSj3nOQ9ARI0Hqs8
p9b+g/R/FgN3ebJlE6GFHXB+BkN+IWByK2Ntw2Uo/FwMqNkUVDcDdNirS5+XKD4a
oznhXCKuuuhkUgKeytDEBBp7ImTfrOUeq7K1cWcFTheSkZuwjD3S/xD3WnNvEVw6
7OLkmik/ICNAxz+WQY/7B6pMDvTuu81vr1zprGmFDDi4MLg0L8lw+UvBygRNuZsP
HtnmVpBPreE5t2f1BM5/FO+Cowj1DGwrMJPf0NvQbH3IL+D8uZtbz+TBrgRWQPpX
JkuJJVi3IW5v6pp8mCOoTXasSFDafoZbMRPD0m6CWA1EXnzjTaMRBc/MxVWLSipE
W/M5R2n02SJXJPWeZT9kLxFfFDzuQsNJfrZ5OWMA94ky+k9BrvqaldV0ZoN093It
nEaNgqmAdLuMysEINJ+QdTXOVzpQVEhDu04Dt73NigJRuhpQxnWOPH4Y65EMCjdI
2CMPlTliQ8NAvhoJsrOqwueID6QeMATgNrZDuhPWlaNHs3uayAzoA2IJbBVHvS9r
wBzfcxaum08YWtmsEnYkgP3hjtOKfMO8VFOZEbQw0MadTMHja4pL7HejrKh63sna
xo+HQnlY0/73AJH0jYgDynuX8gBiuwf1WRKu68b1bqUhGWtXlFvfRmaGfF52ciCZ
lEFtQgM7zvGMDCrc6vZnqaZ8ZqRznAFE52YsCRnohwwVvxAqBgfU6T+/mWuE+SHW
y/a0p2rL3zwwx3Kvd1GpjQK01fKygQ58F+ZjnESYVWZFSW13F+kS0btgsv4l9YWz
CvUYrUviP4M9iLJ3nLMTr4G44nZKgxIsdF1oMlUkJ5OnMmSSV47xDQPghakaYs/g
eqFgI3KSkeXos5bdZweEtJaKA5MAmQS0xp8a7yy1Iaazzco1p7oGV0afXEJG+m7n
EFEPSfx+hG6UON8NNaJbklNMVMKdX1xc+Ss5e2RddcF0gY+YQXd9tz7MRIL26W1P
XLCTm94+ErTK489/wcN0PQT4J3AhK5p4NFtryQZbl7mGQ25jHEAXovIW+fjFuKMD
D7q4vcuv/GEfCH06Xch6k7spmeTalGOlaLeApwwkA/8MN/d1y4cI/9zLL6TzeEY2
swGEIlQu9CerKo/xRhph4mg5jIZCxcaqmHnuEalAOckA/AIfQWcqmS6fTz4Urxov
Fy+x4JNdd4CzS3o1yqpDw0hWaEebUfA+bhBa+785pbyytL+WxB0lLm6HHHnC3vLn
niH9FY4LxfexW0jpvvrZ5jo4jwMtk5Pyyqd0ahP4nmciQqAj5mjvS+/Ap9Nns1yM
WX+6dEaJMtSidBQ28jpWG6xcxOywrK2qJM+koq56ohw+P0a1TBg3jm8lb0tiHXmH
U9nLhU41nIInhKqxpy+oDB/TeK6mVxPnH1+ac2ZqKY+4U+aZyxeDkC08mH1+5mXm
s2j3zspvsKD7BlBweUpuHk5RghiCzd8ttxk8L0YtAqooA5dfJEzac9vzo4h/rmnC
LgS3abiPKER60eEHAunkttt7NMslSYDDcUTKRP8+nr9voSkT2WR8u1garXOWlQfc
fzA1mVCxd5hYjBAicWT/wAM7aCZv/JBarNxBpeuP0090jKVuCNeHmKU2FAR9tHG1
njkAId38FF1o0F4g4wKGb2/cBBGVJX7yX0dvjn6DtMn55zFrJqR5OQsxftP8+Bdk
IStMX+9J0xgDYJeA+dsHRBMrLCD1D5xGqZ3LcaFE+ysJmETLuXRuIlW23exl9x2V
buMwma847BWAUxTMebaDo4SAbB7vQDXpUQDA4d6Jvyc5pu37re4668rbLiJJG6dy
FOPITdYpVFJpKEIaZJHyGTd0LhMErDpaEnzPdwxYIwC0v4qcH1Z0NMkrWQE01Von
jbeTlsCTa1fe2xf5yWlIfQ4xNat3ZYihDPb8S+pG9edUizeAhZbA/ticjuZX9NgI
MB35fEGATLKHiKRiz47wyjD2kxV+xS8nZj3hvmWtXLbhs2+mDKGgVkaY2Rn8jlX/
C2F5ha9jdmlBnviNfA+s/92trQP0+fW8p0K1lir7qc2m2QeS8DZzQqeyq2qwNiHJ
J8m8i0l9fPXrNpwBjEXpi3/Xur5Creus3kjW70QO9g9FZ/LPqfTvdzfU4UdI0qqP
8wYkX9HNTzJ3Bq40I7Q7wt5EuNRQIR4UcNO0KQsVKb8DZ5oHa5teXL38u9chLqFh
qg2qVwti09rI7JImudSD/+0elPgueAi5/hOk7Fc950Hij3UAVqXWdB5/7p2iok3c
d1AaMPmJK0iK7rFtKw+1M2EQ8hU5/4q40RFmy1kiHwxSbOvzDlSe7Pqj6byzu5ke
99LNHs0QwnKsQS8rn6QxgoyU+ZEuR+1iX0aPibFLpa6xljabw0FWCKlw6oc0tDPT
z3k+IzJQHhNDXgwCVg322vR6CWzP65p9si6g8uSmMl9WmjwDp0gPFIsy7y9oWBrI
yNWQ7YG43XyPu62A9AFtiLMGUqYxxM2lT1ULenwpxu3Lao5oNgTcmY0r9CB8O6v0
oJrs26I7Igzw7yObjjmsLS3AC8UCITMvpVFKwJg7C0oSZzWDQQdfOpsF5xsrCLL4
apY59csOA4J0zeYeA98ESWPP7S0r7IFaHih6tC7RrrYHxNNv7Cof/l2ndi2Ry/le
rckjhtR8Fp9Bvo+OJUD9gkqb3Rp87Ei6IC8JiVBwarEXzfRA8UBNXOfF/WPbjs+/
RCTXjTW6ziI37S2wxaE5zSXsUbL0Z2Ku1v/phGOfOZqfltF4Dw+OljMat1F+nXLV
b1lk7M9rYZKpQChHYbv48hi5OVPk1jUFjxakF0piH/noA+mfdGR1Ae6KV8rKMEB8
s6+CfMKVJfT431IiVkwf4eON9/G8pL/u3nGK66Eu0JLVc6AQNnVowqzrY+R9RXZy
94rWMvVI8aD4NHW/GAVI5y8M3Ez62/taG34yOxTGUeUhx5CNpe+nDZjMue6hsUCc
XeCP+/P/DwSPlW5MZyY5TQPjFB6RWJzNgsQaDZ+EHZeA1o/r5M4UXFft5/PIQwIe
EDpSg24ey+2p9lMNczKa/laO0wkWmLFXrDtuaNarwdDmkv1Nn4zKNFQ+6RPIee4K
TDwcnNbT6dEMx0MPj2Wn9Vt1mochNHRmwvZRjDMhjVbLIWeGHyVtr4En/2CvyU9y
dyKz+YhKZpyBj4sUuxwJmv57Cqkv452JsUWJH/VwuIL9SdjTDAekWAW820twzdMC
dBgOIb/ZxdQDnYVLGvvFR4AsltD5NNHY6EPqExdHyg3K6po+D3srJzCMPV1xKe7Q
zMVIyl14lBg3DWdCSnTAod+dVkj7wZ14xpI4a8GLsu6dnzq0lCtGSFHIhTJmu1Ox
j6XWS80uVs/bMjzqWVO5YfTsNSfQ5LrBdWkZx1jXA7SUy7tmrHveJpVt5AS3JvWG
S2wDsUH9xb6KkuMp6fEoCrK189w6S8vLMAPrAWOAGs3qHKmYT5Q/wZm1hIckx6Kn
BnBp++ZXmlfL7Go1GXxlDc9Vd/N9yVt1NKkrp+fZblcCZFdbsnhXzOtiGc/QR6mO
VeUO2l+p17c0b97G3j0ugXLIVv70EhllRtrgwmx9sZBg1TmnGgDtQBEMEfgBsOoj
3imR/MgZGA3wSM7BvxUoAPcbYjYaULsEmKUkZwi2gpYAruT5g26VNBoiKdH4q+rl
+25CflNOiB4/5oDJCCLFeoLslabDC3LHyWIZniOtO/cDCWsE9BizqfNdQMuCZEDc
jZrnA/7Q1HQcMcExmTo2F25MIo2XZXIsds6cC7z+WSfluW0D5YmYr6jhHILWogrz
qPVIGYtZgA7Rk8T5iCr01oVCyX6FD7adDT7/B9V2k+EvEO4iYN0sazyCegwvHhO0
1tUf6QiBqifgV1ZFbTnm0RpjMC2w9m68b/2uU2lC8lTdyu+sJlQQsBUIjMP81wBT
oZtASi7yVzo/XyIlhP5/7VhJ9ULp9lSkXYL+dF0LY2Uuz8W4BmrYCTHCBN2kB3g+
hnExedZ9TWepNVAIN3C85gQk9khtRIwfY7Uzjk2xYrZ9ixW99+eHmYGTyxT83SFC
xn3fnlWupamkei8lpb/c7AZz7yHyvTLEowq267Hr6Ex1WcslltX0ltm9oaj0a+YQ
R/Md0+WPLyo4/UAdcfGiX0rMw58plt6u3B7fIr7grYgrpi2QJnfqa3WmhvkLa/D2
efiM9OuoHNg+YmDccmyhLzTq1WA/REC9cPDnlpnZcm9E/w3Z89mqIdHArbvbJ2lA
G/iMgNT8Kz/73aHta4x8myA0g5J+izBF3ZXn5aOXuy2rgvVN2+8mY4ROMvLvDH0f
dVhmpgC7GrJc0uUds6fLxA7kTUCyO1di/Dp1tqboRKYN6YhCEBfZnjSPX4ME9MRy
h+OHuGOD4/ZUa516bH6HtPTJ8XlwBU+qIBaEQdNyUMJnBRZsyrhjMKTXheUbUjxd
zIftTwXEm+NawwFKs2Dn8QBZDmctUolDJiRocjHOfkX+xl1Sys2dG+RQASCCmwdw
uPYMFaaJX+sUrcDecfbo4gu0FqnZ3a3J/up3YUTUZ9OZREJSs8qepyoMMgMvxo7N
CN/jOLGEQ5zLjX6fdZzJrY52Xfk79fWLdxZqCH8LUTCoy9e6H0+Up8wTOpViHndQ
Nit1Bg1hk6RQl949P4rlF6fDHO+FNjURfLKpGUMBEYOv+PSc8zG0Sfdub/IGihHy
locL04J3X3jPS7dMUM4Kri6czndMF1zHx31DEvrvUFM/RKcgyfmh2sDR8SHdUaer
OQIs87blNNMGi3r/MhR7x+n6LD/C5qb4cu0LjfsVbJhp9Wemdagtb5gDHJRuc2os
6d81HBGySPs1Z6krK0/DZejLDLBjW74qfwdqcKnEmegm/5qGwxCmI9ZwVD6TR1CV
a5zaXCcr00uf6qjNiUH7e3JRAtJ6nHBuqpyMeehayCVUrmQ2Bi79tuRw7ry7ABNS
TzVZYVIK9E1tVzAfIPl/ZhWgFIfyfBBiOPebbWzsYRU+W6YLwXC/E9ADLmTwVLU0
rKROBK6TAztz2zngihcCJJv/+g0zLkzNQvjrO5Zh+cPOZs35JE/7hi4G+QGIlMyr
PDyEsi3GD3MjHkytq7y0rAIEyPhQEW0O8zLxOz2V+NvMismUOdT2Tj3Yo6vxB/ts
M8pzbCOyG/aHib9Lyip6NL0PdSBT9VOg38TouwDREOy5KUUrXtMJJnbJMS8o1Kal
hS84Ew4zOQ177bUBKBFtgs61az4x8rNx9jGHNheVkSIvs7zsE3MORxf2jNcZwgVO
f4OpZ9Z45854p6Gk3+0YsS+u+HXRTyU2sEFi5Z0A9tBulMG1aGz/9Lf6yP+s+FER
yNwXszvWkDEZpiou1HEFv6jjt3274Kb1J6QtjIj/Oq0LTLSiQEra3XB6ZNbE+HVP
DtBRHf5D0uV5Rt0k+WJ59Neqtb0UG8bQ7okTal34SBZ5LYmJCu7F8kXHdS/MMeJH
oEKPoC+eyESE87UIniwrXV8XX/lkNs+L+668v/3Kj2bvZlS2ZDLbuOxA4CsqwuTI
i/U365KrKx0OoK1GRdp3DxwO9sKYJ33nUw0Ik0W0DoxmEMn7wBQ+TizbIam0S9OY
4lCgto0/pBxU6WOdnIRugikbSE8ZSdVXEtkCkesbAF8KWE6AbfiZTJAoTp2KxIVl
MMuVY7uln0+R1Qnynw7IWxriXQ5NN1/QwEQ5LkaHjz3844ssBpiMUa0pGI4xyB6A
LqOele/TqanCQydoE4HfTWIvfTD3TRGnqL9uXlK4E/+mtswsQ0vWlGovwxcxCwpT
DgsrRQXV3m3BgOarOozrsM7AJZxBUPNCX6+JuWaSLOBOPmywIbebT2HQ2vPNby7z
O4JCUmg9XZ2ZBczmjfWIlh2iEl/HDzXygtAlOxtL+6InJbPI5T9vDe5VtlBhxOmb
gwXVAjlTE+t/bGTwBhLFj++4xPge0mVGCTRBrfbRbjHIbjrMj+RlXJKZ1T8We6Ae
HVIMnhY6Knl6CMPYZzN5umkKVRIqh+j7dzxss5AlIsmlz0BXUFTwIAWXX/OMIByB
GFb86/IIqHWNuKXUC9654McNO3ByThP7nkDiq9ubqz0UIJp8XCf9a8hIrl82OZMD
ZYVzf8r/q8rcfCsa4YC2r6L+2AMDnbXEyzBe8vlY8QpMZH0ujRmN3/a5riM5GHOk
f51WF2q/Ws51QPAVIkdoKbbzWJG40ploUCyfOF0qbHWU3QP+BZo7pJ4Or3kzTHah
zZXFLHqp7X0tW52GbUTErPvu1A48xshYQ7kBRS1/yk3uuZTCEZnHpAkbydu9pNki
Wz1KZqjjRRChCj1xP7tjRVuwwOBVavwO14xrPEsqhWtvA++NNXErgnQcsLhSet1e
yWNJt55xspBSnAfjgg4BQArIcLfBu4ixVkuV4CWHnWjQjtDQ4Jlw32a9ECdi/tVL
KHIKV9Vuipe3tk/lpFTQ9+OI9pwacXg3Nfg9nzDlpiO7E5j+sCC3TH8hl24F1rnt
we16ynCiik6s4x+VUc0LlZ9aRwg3kFqhcOsQWJ2+lzBoKEizq+gbL6X4Ly5jDot+
Z5tatRl/1vTWQPjVSNWvSZeGSQIObFftMK/3mUIXxcKt7FY3WgGnkSW2Alh/jfwG
Fo+QEdfNPqXGESnN7dcF/b9tIsBtJM1daBdYO7LcdtOBSCfMfOBkSHktp1EF6MSZ
robdTbPmjtlg2kxKTO3RAPRdlrsq3vDAfUsThaemXB/dh2bHi3OaU1PNe8TZJGpM
2GMMJFg4T3rLTi48OHHdeYEx3bp3ZVQqm1tVuOaNNmnN0AOuyzhWkD5mVgzA+1nc
up9MYjS6/xq4FFs0vkDfCzo1oA/VB1Le3QBWRSFacBg/r45VEmGgPQSx4JP8aTWg
dCgHxHAFu/l53w74KYuJ1ruRtdJEJXM5lFsHpIPncPVYe9yKQ8xu5A4Fcb22AqBP
5jM/cyO/iNlUSqsTEMxs0DjcgvzLbbWCnX8XSnLJul+RQEqY0QegimnkwU1sQVUo
GWpMm/MCKp30cEHprRHJAMpdBPSJcGVHlEJCA7J8L9XR/A+O1WC4qsODhlRtlJKa
ddWbqPh4NWnUlXvleWdzL4aCLMR3Ga2uyoQA6A/EG9rZTDXbKWxs8Um5uRaXG+z8
+KitHIkBAHu8DePtYGXcj7TKnEuPFiW8LGwvL8zyC0ao4QlL5DezQDVbGPUqk6t7
c78KNxMRciS6gP3+2M4+Z8+XFfNT3Qg+rWX/6SrsQbU/9r+8R0E5akPJs0lTyAGR
g4Y6N1OcCMz/aNR1NgIx6k/6VcVpv+ogclYWvLKgm/fKZMrZ2q4oW5elp/5hvjVX
kg5a3EbJgdE2Jh67QMVw6UZHwm94TEvFsTTnRgaYrNkvbIRGfIx4t0nRr5SnyunQ
TN+7z5VCRBlfrN6koTiz7zidTMZAkpsmzWcEawRa3L5wUTsC9kPgqs6N5GBiBkBm
KtFo7NR5uusq2Fv7+X8gF4/fy9Ob1/lKG20p/vkKFbUCTxTEhqUv3QrMCsdW/zfR
qTxAkqwYGJqSsuxPxQEh9RxkP0YQzhMsRFIMCy3TBp1g9jHDB/Uxz0PREskdyEwA
fs9qARQBm9sFo/gPeiA19/DBuqN45sBzd29lJJLNsAA0UyKDE6Xs8GNSLrv4HNXJ
Ytke/CjE5QlrwpeNEslkxQ4BHMymoVBvCO9StAp0biOGVm5/lSS+ovGHtTYIjns2
X9iD3OKePoOZBtonHKxIn/2F2bQim6WKVfqZygOkKmSm3MgYxyz9sqrliYZypZhY
NtFsEuG+NMfynaQejVTWOvl2O4KRx8HmTjPjz/cKVnSrA0Wq71YDovT5M1xsaUOn
9vhm4KMfGHqKlabeyxMTE5XmF6s5AtugGyw2ka6RYsnkt4P+tZtOoyuQEV0wgdk+
29keb2FVICIKhykeYY4yZ1Pmf4skD0maM8ycwBfXWRVJsrw6K/7p36RfxLGIDQ2Q
5G3jDCOQaaNN5PCvwIre3IW+5dJnW51mA9XJv/3UdIJBwohJpipfJU6KCsRJajJ5
qkXCz3AeqIxnD74COY8QqCfAa2iLQToswedhs+2J28APY691O5KAcbIm+sq9tW7W
IqvUZpsPXWrqSLCc5cWgjTd5LNLtNAYMbnS8f4UIHteRnin1kvQ0mU+nGXWGP5Gq
Cm0xynfTulzPQzxnrqWgyg1MOA2kgJsVF4OcC7o71jhHCa8EJdpxON2PWj8h3GaP
Zrkgsjw6j1xfxljhble8vK93NNvaULoiQjTbjWrojXhZp2k7AgTcfDIyB9akqhIC
RDiubOlKcFdMeH3/IpQ6XqDjC91pOmY6X/mMq65DWDXefvLnUV2+0ns8qry7LdzJ
XhPYoz1u6UMUVmeX4hvY2M/tjBSeioROOzreqgJzkuYn30RSIlvxXeSbKRZt+07R
UJqeNGa506V52i5zTmDbUfBgGVSuiMoLjjlzYKQnzsiVSotkazsqwITysquuTRrR
6gNq8oxpztQ7mXJzGpmzySpqvgp+HKrV2K3Pr7nOpqChwXjeLelAFHQoocPTN1sx
yTYgV0crw6CxqoiPTIKTciYTWJEIv9M88tGh0yy6SoAzlKdOyHSR5zJOELFdP3+i
jY09gLSZ5r01eLccCQGrzAO9SaAwEEz1i4VDd8/uAOuSWyveGBJDSxr5BTyzgZO/
oTzeT6y1aC0aOw6Y/npGSogNMYdfCv3Zt/T4A3qwbBviYPW1L2ZIRXwGcQeD+7rD
QHGaNbIwrQ1NsDniAyOXBPaD1ypu0uZtrEI8VtX6K6G1Yx5Ue16paCbffSIwniN1
nemPKo9WzGHEtKZTrf0HI99Qppof/BX9MoWZELjdbinMzu6nzPrLCG8O7KTrG1iM
/wVArffaVTzZhqUZfc6AqLW/+OKjeGF9nhQ290JuUqgGoSxt57wTAuQvgmPT0ZdX
TZ2Yn4A9wDHDWnBA7I59ffBEwuZSdsMTcHn4VHqXSL/y0oy8/QfvnzfX0F4aLRjB
4yawnAzfxEFF/ZA/IKlLaDm2jg9v+M9dQ4t8mKL4v2Rsjkg6DgSm9X0mtoUNIg4y
2z4GC+W7wkNCTJQssSh301QFsR69CneJ0ZfIrg5a+89kPSZiaaWuwwSODIRhL08A
1gF5/olcmvnlG2p5AZuFb6RPCcY/H2V+ommLHfNFGwgBUV16aXD23zlfyDeNFqF6
WgFp/I3JMppceEn3sp1HiuEwqPXOf/P9JXWaWGSVUCiCmOyemCMC5uBm92v5sBwA
52ICg7UWU3jmA7Ys++oWA4VmZq1MFC8MjtQWcizRWmT2ZyZF5NmnQHX3hyLJkiNU
ou8QYZMMxIhN+lfX0ZY10pd5mfs3dSyFhNAeeuIOJbHfRqoY+2AeaMk7SpKc2xtB
6BRmtUdUxRcMFy04Ii7zNxnzgPhSlJZpqYR2bl3204rosvjJysurff/GFMZsXZJv
RUNeX/G5pKYG3MAfuxuxJpTFeCvyIK76bg7INMyk2Ekg24A6sJqhyZpPeVBlPkl0
Du3LUuRmJk1EutsCosOJlBfaktecotTLj666fdeQH7OskEGgF8zLjH0mGSqMPa2/
clI0/jKH0l32QGSDp/ef4VHfP998gbhbaJA8UBRZ77CXDJgkjXmc9CSAY6WnWbvn
vLJjkMXsmp2Xp+ZtUrW9/NFsGy41vSSfwf899hR5RFBo1JGmh5HUgbbsfKQd83VL
rRaLT0GncSHv0XKoeEaXNJ5h0J0pB6bU/6kHqXIUlo/a6hARl8Ts8EThZAvOgvVc
dwVsDtkkB1zzekWWngz8b4ZmxIEkfqg8XPXD7xpmDhfO4mLPLsyEVA/2W/lRd4qr
2WcHxzmZjEe8apz5IPVr0yeJUTHVu3CQiMGz3PJG/IBm7DcZyJonasi11wTqjtn6
HuHhVWKmf60YbKKAG7Cfg/pCB3tURi3tn/LyVQeQGKKJht+l3i7Wyk2o61E7qhnN
J556cd4QBXikTi7Gm+Iv0/8LbOqHZCnYA4FnuARrwuB1Ot7kMIRSM9HrIzY5G1Bn
+oa7P1M//923bAZHlCtYZcdQ45eYJ2YW3jXO3gzGFKZ0gdCUNnGLGkaHucjpcQw4
YHj6ntvgYSUzjBm4mpN798BURzWpBbGSMGwEPyTs4IkQJmf/nGdckFVgypQzgKTz
rbo/DPmVFaTHzAaHeYjvgNFNQPNJUflhlFf58Zx+108N9aeCEYHuGryUyBSJ3INc
g4OvAwSxQQsbEdap3K/5fP6yxb2fDgmS1TRLXLp6OomNlskoKMddT66RrfI2CDZw
XuSYHIPjv95XHZkDlOpujmpra/Td/HJMu8MuDQx6cCxdnwAFIxOcVQzjUgbR1gFW
ypu9PHrODEUobePrkhakczfoFosyyEfGQo0yGbhpq0fFmpbBqEuHZUunLRojx+G8
8FrmMR9TQaINFhq+Oh+aPYsk/TUOaJKzdImOs8SBiPq8X682xVvj/PHc0kCmMMQU
yGtVtYfWs/pjsxaDbqNHNzeamBpKGy16RQgzvtXPedUlK8Av78Lez4wMS0JQt5pb
tgobwzQfvRBaj/mTGFC68qbTeXXxy1uPcxqHElZvXnFS7Kb+BZCVjYpeGTNELl7D
+V2VDixx7B31Xl7/lgOe+0nAB88dH+PxVXnkg2tClgIbrtFqLPX7egTZQAktbmDi
XeFl7gg5kNstLQ7sM74ZLNEsscRqNbhLZNTPxxGm3JOt1zPnit7VsBcPe+sLoCuC
PpNECoafIPKpLrwUM8jHG6ywZNr8U1l7uKmKgmZTQvJ48LyCkh4hZoMrUSu9zNvh
Vf+gItFI3F1i/FZYLMbxpKdwlNRGOR8aEzNO6PyZMntnDw5wGUQ9A2qnblJFOME9
7hZpBzyPd/R8jPmXUHkYrPJfQE5IXgV6QiUhXKfMdFVE2DEgiLB/IeRAy5Ifen8H
8ucQuGG88RjHeYVOgpM3XerzPustqarHQKulQT41h+PBBfg7J4MMnQIaHiQdZvH7
IOlNzVq9j397U0VxehVG0J1CD8E9Qd4zq1Yxell/FbB4yzHtFkgPSJsNQxLuaF4B
SY0IBU0O59NdDPInGWJPx01bMe7z+aHNRc1vokjZBf0qHi/tyHwjEyO6/vd5PbY5
ItzSLNKoevQG/U7eAgWW2w6zHq4W1fAtZX28HvBwr4qnbuc7//dpQq5Vj7gFbwtA
wrIkCABqR2egMABfeCYs14oMh7YBM39fmfGnuVVYk9Fr9seN9QAyC1fE5HZobSJc
OukhDNwHXaaPNtqqnIL9Vur0il8vf7Xq8Y0yrQW3Qw9zsCGaUc43GtpD/b9LEPNU
Eckykyqk9/+nQ88y/p5l21jqtl1UYc2tv8KqIg8nzu85YiCmj2FUr3yAKASU/zyx
6vNXydX97Rrwmn7MztSh6Wla0HCITPQl78nEySfuUqMyzNGNkVn7u7COlI0ztix8
VKCVSmFxOjpMPH9aHhihQkaRsq//EwJaVse/aR446d4ORjYijzeanuffHjDB3aNO
MN2yw0kt3GCs4nPR8B7Yw4YXH+Ij7AWOxe381g5HKkpD2q3nX3/TJ3/JUGwZBdoy
+rHcWzt/qp1zgzaFwDpbBGqdjn5nB9Uqlo2kzFC8xeSp//v6VB70r/zon1kXn0b6
a789WIleyCGOHl1Capj+ue9UVI36QAkqjd7WJvlwDSKNrh+MKQ9GbSaKVY7vs9Gr
H5za0IqC5caEYXjNhT8s1kTE01dPMxZkW2UhxpKCI6VeT74ra0YNx5kD7SMC47XI
ls1uaxbdqezqKB5IUYmoYkRPjrC1r9uhrE1c5lTmo79IpVrQwRRsRw18YMxQLDrK
9iv+j+qNMgQuXF31MGm5GBEBCMWtLGsCRGzNid1S8+YiCpDuMOkJP+T0Fjh/veRu
lSKZjW5S1aPGgFT2bDB0JNLIGicI4t/TM5AXwUrQ/fvSPSkoHxmAnWQHJHZ7k8Qs
jYrr6qH1dCn2jueg2GyUhrL/+zV5hdhLI//4C6No3qpVHPbzvGuhCi4COo6eyNdq
1peerVnhMn0RWrXdzYVhtadKVGJxltdT84NLr6LqPSIU0sknf5W4uVtSb/INShdf
qsCOfbS32WCwNjzDkRXB8nqXQcwhl3AxJuOVbuPLXdMQRcvV3Lp7RLNrnuXgrsso
XoOFjCRJQD64pr4kkELF6XD6Bis44JZ9urR+DqE7StAt44ml1HSoOGO6Pn8Y+AWz
Z8Ow46J0HDNiSeUwu1g31+WVv2u5ODrMQTqwFBcrN2GYXn/0DN7b7Vlpk7hWH7xA
TILi6P18BhvLElkurxY9bF76X3R/DMxtX9aNkfoKXa12ToiSHZ1NihE/m3lqx82l
FpkyCq5UCdFcPygAQZ31LRj4Cpkt5QzHn5a4rN0X8HxifioST8f8p6YNNgO4XOkZ
UKisM8AdY44AdPL5buGjl3b/XBfh9PvlNi45+GC9DlPsNMrePKASK8iumZH+vrZt
JA9Sw+0IRVCuuRYANSfLo4WZNLpdBIDINxzVQiHI2tDpceeM2RgNexoANNT7/Cx2
loa/T2zsQ80W4ELE2Vh5PQQxCC93yBQXITsFSgnZENzyuk71FR4reFUw4Qtt4INK
ueBvcBSLepUYuUy56Tt8rX5ZXFWIBu+V00cqN4yzYNPDY9sZgxoIbLVge5IbJFtS
hQpTQYoLrCLmvgoQR/DfKcIXr+oNWbRLe1+xr+q8KO0JiUuuynQKbRGdwUGmPPf2
XgOM6Do46O+3+rSRQEc+8Gm/3Bhyfq6sDv+7sErhZ0PtV56GR2Nzwafmgasm8NQW
Kuuf8cXQkD934eDkedBonlNWS6WgA7zPo5wkylcGehIvnSNtm0iZktD3aNc89+zP
S/lBQ1AmoeOyNn2tW0QC3jDLI5dGY2QOcHgsQhbVZvHdULDwUVhdQ55HwekIKi4O
siyOaerscEkFguW3VuE4JVEv+qPC9OfkrO+qYUeQw/hK0A3ZcYalWimg2/aaH8f/
sxZ7SsCpsl/51grajPCmHf0rePOEggwvcLLeFfBswLAE2TmSHvsnYiWtEf+UTjtn
bbtMRaH8/SA5blRI7+ket24HGPLfuCO9JeCt8eK9jeGIUfWfnbvg+2gAGG1BRhWw
htqM7odPgSply9JuVp1dHL1H3Ojkv4Z+03hRmwRMJ/7NmmVya2n3+eHL0YQZBDSc
WJoO/BD01cI8F4OamnDjku5nrayCfahBS9KKYy7uMrGL0mtMi1EMHHsNz7r/mRt5
/W7zSx/etVukJpY36zWq4V0pRKx+A20G5F5OHP+ZiABNwmJFjv8Q5jbU1s1Bkztq
NGQj7weokGwT2LrETXlVhL8Ni4/PNJ1jOc6NI1mlee+V7FNlA6JaRlrolzC4/62+
mf6fkBcdgBSZmUw/wRceCBo2LtkYQLYzm4iHmlU/GF2XMuEt7JwgQ8S+kLILfO3e
h82vWEjsJn4Lg8yxEMz56M+zf+YNRFe2KurTUTTMGdarGfSOegPPP3luohfQKE/6
pEYu3UrObFdl4H48Y/nDblV+ak4UZPc/y2JqhFStO79EOW5JgMybRj/wvnq+qC+a
3dWfcYZ1HdthkZVVYq7yjjuv2fgGaIexuOoKcFQYQxfcyQbN69El7kyS9Cl1p+yM
EdY1RpDcMFa0JUoV9VeUfsnjzs4gV6FXtKA5JozaZ54q2Dy8mub6KA1FR0XnlkiE
ibspaxaGwt/ZDhwrOJYuTM6RsP7hCCzIwjbKSoHlBvP5uaXubcJjS89CmQgSSkmM
XUtvE7BPWs87iVXcx5boXTsUmIPb7H3BQBO4a9Hg6Gp7Q+FXA2GMO6V8xs4swvpR
0s/HMoCr80nGUqzvYPAHD/wiDS+5wxh4oduFK3LzG1QNVWLmulvp74ELfOVE3Oai
kd0BqmcWNTmc+eOfWVXLTQzmpgqbYcq+dbG7XhcIEuHTRAUz9PpFKpMYbeFBThRt
AXovUhJhlOPVz1TGY2Aedws2KMgQ2EDTHTjHYtskycBMnu/NBzJlJOctMvn+Dil6
Kfkl3b1UylS7UpxjIUs1FUVGDGHco2JUD7oXu/qnG9LxZdH6GpbvX5FiVvpysLc9
WMNACUC/tt4X9M7q/wTz/0HwCQI0qOUggdyFScHWUAFKrovH9kgkMoHybugvQhPF
FLVrEve7rWAQdjvIKHnmv70j57FlGulag7dEnguvUUNqT7hTUsQUmlsFE8JTVYBs
jhlIbyYknbriaxCGufVpwYuxjQ6hvbmdy1OWgvRcQXXp7UjjRDzefRCEc4O1Nm4W
Jgi14u89RX08i+Dze5ux2+YSRyo4wdhNNN2vvzS+BpW4uOjYgB3AjwfOPPAzQ1zp
Bq+MnncOjfh5DVjuOK3gUj/dPsbRFACH8yY7ENRJrCCYbIT1xJPLRdIvU0yrB/nO
5gxkiUkeCnePMKvjmRHbZjYmNw7+nssseXfLUCO9pErwbFS/ajt7v+F23hIORyh+
og9DUQ+AizeqDu8rpqetSqWS9hhZKxFumIr5bgTBFli+4iMrq/tVtUd6FnNf1UJq
uE7xvMrT/nCcrpBbTHtpAg65hRYVaaeEoho79ITwNllDSUrhRc9XWw1LsRMYToOJ
T1OR3DZ1EGOjHMR75TdDfS+or8txWdPmCPvmTI1OdAKTHN989jmQ0hj8wu5079on
Ob/zYZ5+b5DM5T/xP5pGlTxYBR/Bmkrhz1nx6cct6vXLxxUP9sPavo5CPxmz18s8
rXeRBHna9Ncp0YR6i94yxOlTSpp0IjLTJzJur3x2M+C2ymffvry3MeZ1jAxOH6Zv
E1MNquP/AfTGXyPpVWJWjDIw2ABfaNQRxvL8Vwy9Nqmq6SrNoGet5zOrLKhoxD7O
Se+cxFt4TIdkax2u59K5Wxa1TX82ODeXK7NjVKjucCnJxI5s2WgwfsS7TlQ5pwc3
Mhj+i/2b2nYbTjSU1/XEX1Qc3jt0ExiIoUbClnfZuny00Xnxw0AujgHwii1dqmGZ
xRrmtC/da8xgHqQTkpB/YqsgzduilYgS5ECUh6rNcaV3A0EDxTUEAQO2EmFPvWnB
dtQ7wBB5LX84/Ab3VZ8+HNMCEZ95nYqEX9coVfh6HcOBbTC2SC4tCwNJEm2r1915
Z0ZyHW2FD7/WFC1AMvEjNO4X7o16/ZBEBx8ijRffOj+GeSnykaJMHCpmm43rYQef
PagiIQKMD7wEivw+zH762j8U6QhEP9Vujo7c9w8WbtJCOnNvenVYPIBkkcnZamso
CwxRXFpHW/w/cPxRc/jR954FMCU15nuODiSuSqSwXL8qPj2nrcZWBVSqaWzDGfhb
gHRG4yBykh5UiHN64U+crN8ZU0InJfDSc33H/DA+N799ewE7vJ+9Hm3GWLcYyv2u
jBcxD1WE4T+KOQV2f0ow1nSu0fCS9+pnO7xusjdhi7yh5pxSOFt/5jN7rBo8F2cN
Kl6pTXnFosGUX/M/1MnzG7QF0TzVp7Dgg9CiXAWMlBbhzOvHm1J8WVkpkXBaqIS6
1L7Z+m+V1aPSm/H7I5S3NBsw4rSpLpyeWd+FXS/9xuykD8aJ5YRgdjawmMDDocvY
tJb+ozNIUQF+SB51Cm9HaP6B8QVIvSjaNSCWQ1CSleS/0hvMAPL2MvKjmsuJcXqk
0HsBijrdYJCDeABdYCJzbc09kfrMCw/XnIXYWUIO/19KwakJLZQ3AgYskftWa/Ux
ZVzpiTGPKvIbosXiP0FOTV1J/ZMTB+2RM1yIPQMR7pPqSqsos8+rDKou+PreUfwD
SWpa8ttUkAn2F6/vVIYenLfXjcu4Qf+7Bk3BfWNANnf/Fb5mx3LZ30EZPCENpT98
sTYLqDDBBgUnq56NpGAzxKztIlQeNXUnKOZPyZrGc3Gyt2AP5wa6Div9PIZq2n8C
Ibor0P4948e9oVAZg9PIRNGERRsd0yZs1R1zb8cw3n5WNF+UfFGtWYOk690cybGO
u+3LOdbUcrsLERijLYgFyIFoQ2xg6+LG+oP+H9mlHB6L9O5iRmxn/r4jiGi4BtR8
MEDWt0Xjko7o0qlrogW1RMdmdvtu4J8rr18Wyio2vIW7yhl8q6nxFaMdbgLM9MR1
6J00u4cG2v/YfZzOYr3WMEB1/0NTJYvPmcebMABRlii9ZmTIoOHolfCyhr0HsT6y
rY9v4E3jcOQmkt4GXWySZ7OhbAVcSja0m5snAmCcB5Bhop7cWbheGIiokCBWx2EV
n9Fs5ILg6gUfGkAJwBZ68cSRwNqvaK7bpdo7MVPPmVbfjePJwtFuYzjLrYtZiYAP
9urjqVo+7gGNjbg4IXHzDq0Uw8bFdD/8Kcn6nKiNFRHLgY4E4/Rl9Jb8CitnwPtk
MDzxJxUYlUrmCMZDxHadzlJSJDnqMSVKd6CWTnPGjS37js498cOv9augFNoEiuZI
NcLfXTwYTshN5kBOp9Ug3iVVfwsLZeqAuDboskwes1ggejM3k6OCbHxP749HtscL
RhRxUizXAnUylT3UNHm25D9WRdm8KyKajQ7VeRIj2yL3ynBu8Q8pGFeMi0nEzo86
gpQ5azNJLryGl4hsmAwO9mvjc3ldIWBrpnX11iB49zSMEVz2UZNlVpcSHN1rJpeG
16gbpBvYaYb7zviUZuDO7bPjxrc/RCiaMX3j43EnWxbca7fqJRCWb9jBgSBS3JED
uoKbbUxgzGjMpiq8+bJKwlkT2seIfX8AIYVZL1ezDxKgpOuHlfz6eVE+Ct4cUKvs
sFfVo2T8GZXGM/2tP8lPE+AxJa1orBEutQm9rpOTO5WXAqO6EVfnJGC9Ycl+q/Pd
nRXZI57VWPLHXOT2ZIyRpUNptHZYCJoOw+f1EVas75RMvC7gIh1jAIzibmmv3SnN
OsNMVCrBt9PHg+UZ1s88flISRwU7F7yzPDb6YzEpp7WNyBNTgHP1jj+WbLrQYNEe
3JoNgg8bY1BuHlNLYt1AYLDSGMwuie9faK+7kTJ6fY3VIwWItRziyWrhQmBOTW9n
H9MpDeq/FguVdQvb+aFLMoukHNHIkYxdLr3lHBDBw9UIfzRA1sihRpQA5VqYrc45
bsWIa46AtDWPK1mvs+wAm+ZrCFP6DRVRPIgA6c6+85u2azUZ8GHCG5XBv5Mm7PPt
2FkJjn7sBdmwQc5nIYhrbYQhrKsnsdQ5wyEwdLVvb/zkusrCidQ0HJO8duFydkzE
rCmJZMlmmitxtxOzijRAhOgwmUd4joyrvhcEyMm6w7RCL+SQGOeGc5+wJIAWt0VX
BHb+tXHz8NzIVRFlJNcJ5GCO2MCOX5QS3fDCTnicKTMNUOQ259bKj9hljgGdP5ut
ssBJtr6JMAM32im7ifHvmlXBOs8E2+UxQ8BeePCHHROfzL7pOt/0+kCthjnbPtB2
fu5DM+hEcFqEaUK1X0+5yqC5nwVCKcM3qllLzjtgfyYiNpUL6KQL6cxHDQDkmlue
gTvQ0sRcRxo10/O0xL+1XshCnz1Af23bhEClZ/HA5oYINT+KpEQQUybXikjQj9+T
KmLuNwDxAZ50pChOXfp+o6nuBxTYSQg1hhPPd5maoPA2VdRfUiHr80HaYAo67KUA
D4Q9pNLtHGt5kEOxx3bcf/Diojq7hfHkwyE/+sSFwrHgmKnE0Fl28TDOiSmPrLrl
fg+HOGNqkYy1JJQaNmuTh1JnO6zT5dYzm2eBgAbfXQTMZBqcO+KT1GsJXqQVFOPB
LO+OTt/d4FMLBkPvDTt6jEz3E2w1OBGKYJAH9roz+2af1obTbhs1ROuCqYrbhlAk
mBMo6wCANScNO7KvYTS1APk7l0LZBGGQdgPGJPBUQVpQA/+rpeyaPE1wpmv0OZY8
gNNwrYRoLwOKCYDqlVVr51svb0VNZn+mkz36RpXqQU7hbucQis56NU56FFq0rAJa
lY95Uai4VNvunCdZVf3TSJCuLBGBwJcGZVoX3I0otkJxX69Qyy1APmoat+byxgYy
BKMbEGvU2O5Q3qoRQACEuOHAwb7h9LnQ58ZC9OPLzX9p8ZnDnJCApDNaYs+mqGg+
NnyH2MKm18M7PKfswlPyn790r63GuhABpuBnKR6pbRhOk18wvp8bni32DPTsId5o
nsdWZcua6ika+VQlD/ftVn+75volLRjiaHp6M1BiAnui0RTnj0ffikfO2M8JBA2P
Qm6sseer2k0+tmAWf7lQQOQdctBFS0nWsYQ/VtECEzXkH+YGsdS3J/2T7yiikrnb
HtX/tMGt4XQf/dM0f/NN5Pf9kEHX92PWvuIRVJsW9Dzhah0dVQjuZB/A4opshZ3o
CI+iN3XxhLOSbHrrJcZ7+9BgJ7GNEPd0/8iWQACsa7FlfCvFLR1XeaW98EnagZGT
99MkMl+6rb+3QgVzgqVJ0AFCNgNa38+2Aj+HPP50UoRRmBc+fX+0XjOHPbjEeypB
zIDinOx5qCDhJcnfLkILlluBNfdPMt4GjVC9niqDcAQS9La7iUbv32mn0+xfm/6H
cHY7niYAHod/AK3SSuTQ0NYeycZMYyWzkLylEe8vQVWczv1o9E6L94owZ4cWbgVb
KyCbIXfPXtwIu2zArnZgqGw5syMSgIW4ZUIhQ5usR8vHWjDCLaQ2PyoTzyvRnj25
92WF9ztuw1y863pDfUVB1ycE9udBnddLBh8ExiHRs/E8uN4GEXzA5lW4qvFMOi5d
CwhbN/FVifVS0E/4lVi3g83vyVeabvUXv3yjnoiCpiV92o7kvDtXE0JwB/jRiqAf
vsVVB1a/DBcd10dbu/NhAY9CiGdbMSqL/GskUO1yG6+FscbX+Pj5l5XYRF/dN2DH
uMljHQAsbit/LPiXG317CGinmAvnZ8a9mURZzt7WYFFJ5e73IBnyqpmLvrEg6Dnl
s9/piine1d15+w2Zaje/jfmncvy/eDSe+f7AudQabhMwP+6DrjwQH7dt8rcBDEyE
qMHcIGbwkJ8N+z5PPzD3/ps7frB5R5bxDEN+2hAqVPq0bGxSJsB2kZRjIt5BeKgz
ie+SR3C8nrwcUl9zWko2c7fM4KXfZf276umJRg8OdIB5obmKek6SlAIPjLrwAHvt
esa4gsCbDMmKTo5XdQ7+K3AddU8NOYOCekTAz8EGYTomtlQi5gXAWs2xaF0DGUWS
E2yDKg2ZokXEIcHoJPVZsV70y8CQIwupz+4y9aH8uj2FdrkUGQNZno8je8r1x+M3
kZdc0BOWDqlRspH7VYoFbxLDtcYXMgqul0d/0fmtnpLGNIIKa+91ZMuphfwSfN22
OQUrzd3C7es/OYDZ3Bw5uUTKiV9Sjh+ZwQUPQCykSsDVsjlg5yepjIDf/DIU2typ
fMbT3Iot59HZUH5yobgvsmcKHpu8eRyDFfRpi+TxiG9UV2x1b/CIZZFfTNIaZs2f
SEfadC6v2Txh8y0RuQuhtsmtWVvGbOaAP8+bFGjwhvDRP89/bsFxyQcd35uGadx8
VKdN7aicpZqma1KMr5Bk00F+C3n8tsM++Li7sKmwyQ3epWCbe/gSHx3/vz5xAINo
4Fi6RFTXOQLaYx1ayx1d9DmjuWw1+fTSnO37m6HR0PDpf1EumFGo/Vl0gqbpcCjW
SwuV/Z3o0MY3v8C2a8Ob7D2ueiZQIyRFKO70Hbp2LFynMOC4+DJIFpGSqF/hv4bY
XrPfBxkhUsLO90AFv8hP9OPEB1YzUe/Kcb2OGslLsFUaREZd2kYZmol6M6OwKDhc
ou/qWDIT3696hXdlqMxxKCbcEDibVEAG0/JKduZnd0eXpV7j93/qwgOlKaumBnVS
xYyfwGL1j8AhlU7Bgl/K+RdQpliPFBqHf5crs0IRUWi8/GYu4rHtvZul46/Mt8Ih
Sjqwux6akJS2DwQ1QlHHtD+OeNBwykTp1z3/l8DM2U6v1yE7q6FESBi6xsuSnYql
D69bsaaFvcVqFF+RK9QV8hJpCCm5FAW8ZuIjQFtnjZ+CD9mYW1LHeeGi3zB2VIm/
VrCus+Sr6ysaJ9Vf4yZiNMqTX4nNFBXdOtK4yykyUOXyIxa2mVw8XZa8BHUl39hH
81HIhwROXEkCBzxZY6KhtW3Q7DkX166ABgX7GaiIDeSQByg7tB7u9kErWQQVawAw
674pRSatakC+Th5nAG0NQakhcthLK4r+pQ6hhnwhR9aWy/Gfq+YuLFfBus1Ujknw
86JU4Kb3luZqc/nC261ZC3VShbSwBF785M/MwOn5fQFkREcfeWWc/+WilV6FxPXw
pKacqXDbxpVJLK7BLT+RRTghetE1Tt/mdOhhZUxszZouqukvIV8XO00/LpQd6trE
713AGB0oZWAkS9+1gNaH3FCKk1eOsfcA05mQXOFBlWSd2Gcsd2kfWuw1TOy+22ph
SCJnu/nY7cL8d8VM7H/hEO+1q/V9a8Fgs+A1WuVK5LjZ5+ojrk1dXf//i6NfSaUT
hfG40LuRBf+aO6Kg86CGN8OgZ+Wz5tEfY7qy2DH39xZA/LgvJZv225Srb/5UKcAE
V7BnLANf8Rb71FVpOMMym1rIsOymOezJ/QG+oMQtrGVoml8De4CwgL0AKWDpI3Dg
pcILRmcgPmR0b7681hQFwZtzdZi72za+WDKCqJ8aG8znI97ZMez4aH3j1IMaLNGD
no6ozXEhSkptjxNSpjDwR8FCHrSsKft5A/oOQbUhI8HBrm47/FWtzyO0WCPFZ0Jq
0T9kKNXk18u8jdbGu2TMswCa5FSllQMjZRXf7vYtzsO+yUSwU8NGrcwEU8wyt2x0
53FyJ6S0eeJGW7hoz6xEFAeGvEfIwPOWNTnETG9A5K80zHb+2kMYl6Muq9IqGFrN
+5+yoByXnVqvFMMstNBaNoaOXHXb2TOiZtOA2+1CUkHt4cyIoNjEODbUpBCZomye
GeoceHtRtqyb1SgyPZyeYJop5oZWu/fWIys3YTJ3KEfXvo+R65z7a8z/WA4j8HGA
cS30wM5zif6PrC8RDzoLtxfyMckaNm9vzJinQYJfIaio3fuG89WmO0alT+MmUUfn
HizUAYfYt/4uYvIytR+U5Z/1eeo1XMyZAJ3V6n1OnzXCoL+n7+PRmihbsE2sH/o5
mhbhXb3aLRoFEMxkMVOYHHveU4AD1niH9NchwaQbPIj8ZZ9KjlKqiWJYwPpgV+5D
q4pBhej8jH9e8cKYB62v27Qqt45XSht9R+KVo+FAFoBGztx81VAVbchJHHLlBfy4
7Cj+L83piPGsLp+dcZcA1ridMvA9qaDGrMLLTI6KrpKGG4L4XQpj5hN3quBKrAdy
FTd/mSRjjaMqQFUQzuGycE4Cbml8bkhMMf4pLmsj3R4SEO1vmzkplQeBpwgwWWKk
TVBGNBYj5BaXjhzeR3G07oenDsf/Xf+Xe/AFZDpcGPL7G5VbHe2EKDCYM3AQJWVX
8SJ8tdUdFdAYGIcGgPAd5Le71PL9WQtQB+diFUXs9Q82XjEtSs8dDIOqH4U47owk
AF8Jb1y39VmJ4hAvs5iK8nfTdpNAqpVBtmnYWwd2By5ei64otbmCFCXlHA5N4u2f
IUPSLJODYF5laYaMXYD2pdlC/GBe2J7Vu9BdooM0Ee9PjF6wsVouMdimTFYH7PxL
uBGAB6StYM1Sl8ScFgeMsVDC2Z1KPxOyp3SLVjltplk7KUQ/B6+ewiL7pskSEBGv
0EwyfmfIkwkXdXuycCBu+LOzMQs2Y+6lpcHXCdYBxUONPrtA1OSresOtrknOcptE
y8QQPwaJ9V8UP/evUi8egWS5GKQKU6BjuHahFuQDzBk8e4NB0PFaG8Dt5tq1luwY
rL6bBolljq7xTQ2k64Q5ycgPRzLoAhhMDKiQTtvy6YycJQDsdZ+22YWWjhwX3+BX
kPIJ7wNZIu822c+To/b5KTX5SwIepEJ0axrdlbxnaseaHAh9ataLjGKJbhnLQnYz
TLVDgj51+0IOlwsntJsUDLKDDqgUAe5zQcvJki2gXUbfwVUv46hEXAJLP1kYRTMd
Y3DD5ilHy42SLHuhSsY9nqRRPQ/NoWVC1Ht+OniX49C+LtWZRemVGfwLjjv+P5XJ
GEthax8pwp9YMQQhB9XZXSM1rPs5jWYyPCtyPsU1talTX9z+0++lSQuNv1h3zEz+
+Y6KXuq6Jx20p2MlDdxryQn0yxITYVYMo4OswidU5pI2vvt+YK7tROfRFsghGbOC
RplkkveXx7Zd+F+iIkEBVnLvfz6R3Y6fUuvdB3juUxMfXizMGqCjzH0nozJE3tLj
wxeRwTT9GA+OOsTL4b21S+9pJ+CXq83NPkbEIbHMzk9GE8qGAngVwHu6bPXavfrv
udkAsL5Kpk/tCyeeq4naUZss+KtbadTXfnAcoZRuJtdlGDVtVGeaChdpe/nUjq4p
A7FqfO/U9MN2weVi0Zo+m6qAUNb50VXCyUce/K9gZB0qeWxYTcybd6t9jnjvsVid
qYypdyFR4TrOTb1pgyxXSlnt/Ut7xLhlnlGzZyU7gvyERCZ9iu2NeVfIPne1jrJA
AgrApTjU3lgQqladr1HiS/q50WkdK6+yV2rdzi68iMPGeQAlKNVZ0E0KhhD2G9/n
RNHj3GNRKeqkc7czQCF+e3kTSWKN3SamfYxkPx16c2xtO4b3JxBGUNzcPaRXGnLK
K+XkH/J5Cr3jKBEamQTOgQDVWB/r5i/WUJ7Q5NDE374ZljfJkKdmbnpVJv9KZ7QZ
PpCzm03aWZaGteultmmnjqh1eDhWlxep/30XMme1/hn/hoZMMC+vQkzdSM5+URrG
WL1GNsWyqa5cVn4rzSZ11C2rJTK0DlFUIHB4VTejIFzPLhT3rzU+yt13JVboeQn2
HG2xoIpg1c6/mD7u2C/tYi5ukhyZNnyTTnOtxCgd2/8EXLUmCeD627YBaD6tTo10
CiMExvSfKDiKLF3Wc/jjAFeVZ7ciKouu0xKfRH20mDSTufakYGbqeoipIeLitxpX
uEiMOtj/vkwaaOkvqcSQKbxPdMCizpfmFhG0i3/wE7YOSih+dzU4j62qp/CEt90p
V6hsIvsvBv18BfEz8KAmKqiOG6R/aNyKJ8ZfQ2gFwLk6o2bmmIdRT4UCrkkha7DT
tdmccCoh3IDCLEIy6a4eqcYr7F9JYRKkZmZbyVx1cN8s338s4Q51NzH0TjOkqQ7/
RVz9uXSYRwGygahC/f4L2Iy4Fc3lq7qr9b6m+y+lpPiG2wxaFSHH88IQPrL+pZHB
sVWeTD2BgOGQR6PZuuuUpUnWB6pSqANAEPqbsvRPiiM9FMVykCNBhLRPqaKarIIl
1EsvYspIiA9nXomucNhWOctKoLNJy9BU1u9TS4IphQSNxYs3fVy2fZLRrnGUkwrw
WwBXY9ZP07l7lTmicXQZzeftoAVoxICAJBYAgqZXRiqfjIbHML5OkJ3r92FvYDnj
eFS4EMVYXhV4lXR3OG0F8YctPRXh7eBQTAGFkPNbHz0BdUUcjC/ETDTyUrapCNoG
VNnSCXtrdqFrnYSg9HYIAyeKxqT7ehJ+/gEDxN9mKUsEfL28wM/SvCBcTAbAfdLu
hsXFVurO6ln9/YlTrwU+7yHd9bhFsREiDl0woOKN96D97UD0IfqOBfPPARuxkv7D
f0nrLUM/rrii33ZBsurQbPGzzrNmwNsoGoMWiVqnIL3vOAyGfoqhL0K+ax3EjXeh
BDPQt8bKgjz4IxWR6k/9+4l3+KTLeJUGXBVD8j0drFSp//sMuhYgIFmFkHfBrdAJ
JLtr4qECrcLleJnrN7EvB7SFDp+og6iZ4pJgZbBJZZ1WWtGsatbuZje0q5ChY+ON
dhkrtE1zCKBH4Vlo9v7s7F9iSCtyv3VnGQ7R7h9xx3xsWWFYfS1oerLqhovsVklc
GFoRdMTxiBXHyr6Qgflv23lQk02l0K5+G+3QI3sXifN3jbRofrk4LqwUOioaaCBW
V6mVns40mEZAhHmg/xtEy63/C6u+QEw3Hb90E4dGpBI0Ycn+fncy7yJjx84Png23
hdFkwYaM5kYLKqKapBKcFWKH3mkG+fqXIu4f25vSiaRQ1pz9exMc9F7uabG9B7Hx
PSwCMnwVUpRVqhl2FjKhHI1bJMLP5Lx3job5s8zuxKx1FSpY4y5WudJte9JwaT0j
D09rk3jTotb4LbJKWJSwB+S3DxeDLrBWk5aHPrjAlQ8T01fzV/+1pFE3dfgCb2T5
O64uaAVDNvw6kr93LRU7TUZJoUsncfSUkfifQCmMBXcocEaCYgmJzp9bovHLapku
C0LYldMSFNGy7YqvMxdtP5SXlGLE556PCKCv5yOg1PNnqOPwv4OI4pXkrVqcnbCP
mBoFiJYCXI57Pp99LtDqZfv4THncTexnF8Bsbqv9ysYwfXMTyDnMyGlO3w7pf2bN
njgiTGMQnhYgsrV0qGKFQhAAJMWOh1UPvw//Xi272wGc0hPqNdAxPqbu+i0TOCjW
h2fexqbfTGAjDK8G6kipoICe7fZGYrmt2q7XI6gqibojY2dBOSnp4Q5TVkp5FV/r
2puPq01ggTwDwb+pr64xJDMa6BytgKLMpLlguhkViMNoRdkwMFmhheKZx65NwGHQ
uOe+Nloxhhe69Tkj9QvPncX/LVCr1pU5lt12iuzNWuueOY6cApwV17ZJGE9oSPPH
uGRNWLyc9uA+HLswWzg2NuwwyYjAwQWOK9jynt3UrG9qWFEWq44JWoIoZgQeHZ2M
O2GoOELhxWrSYqJRlgrWMqDKYWUVLJ8Sca/xB0NJMThGvdN7FQ3JOhWywUKDdDbV
sEXbpfkWRevkF4888vly0N0ITKzNXkpfFDYm1Av9U8QmiDuDgpWGYw9Mm4h86gFV
GUqfrc8medoRTHxZDxb82dDSyJ1YCq6igyy8RXgDU+PBuSxmgr2hakdbNDOcuHUh
IDYvC3tyU3cHOkawKFY5rvurQm8+5fcfVo0jnIugrJwV1g5ZjlayKwc4me6HK3vk
Gam/9DyRcM9Xdc4mUZFHbtipPAB2WsRRKbUEkFgO8x2r9klPqjaN5uGUc7O+j0Lh
f64IRzPXlixciKp5EeEagBs54OcFDqkteqqhyBOooTmCUZ87RnSP8+pSHMJ5u4rq
EHUgLurDxhmLi+rhRiHK4Z+XUjUdm661ME7K8e++Pzr4z11ECqKxbtM55zIHEfVR
tQCfDQ44tNAZI8T8gWYuhBAs9lc1mewYLjeprMhNk28/2A5bSoeljWZ/BqAIjHSD
tJmbZwXnqJdb1Y8tdgBMCW7IZMy6vzUoMMLnMkuoNyCb62Cqk9komeFSbt0JzhXK
z5zbt5KFLMSWPNBDjQEAM9Tu2RHga/8kVoxZdoQWBmGQZx4QlZqnetzzjbh3AXg3
/jwxXXqUKZIWa3Cy4C5MGy4vMrHH/EGvoTIcXkYGN90g0aL5+OuIXAGOKa4f1oF9
m4ZftnavxT+EeSDlwp0by6HCkJ6JsKUyvJhM+wAP1be3JuA7wO+L5L7nrOCr/QxQ
IpOMa6e02qDBEUKSeMK5op8YN4+cRpbr+oJLPUApGDrBoknjTYsiVJ5WzDD05PxW
TU7vp5Dd+aDcxp3dQFQwROklvrHKj1Z93seYxHkJS8tWYTXWPTUb3cvXxctD8U8S
98D1ACa8GFR/GW9xnwvz2DNCKrzM8uyutHJNsiAq7tZL4aKNETU79fFSs/qAkgVi
6T9sAfb1msQ95rA82er0GqeZfRjc5cj2LGWVGhYWBK91xqIb+xjEXmy6n5JSoL0w
ZXO9Ew8fXeFwVIZEXwDeSyeGCpSuJSo/ygVJfEqbKpFpDzaNQizSch4F/kVyWEm+
LrMtRpCJuh13Ot+N8XyyEQ76CpG7eWd5vs2BIWp4TD6iyW60xq+SH4Iq5Uk8jt4Q
ywjiOOHTHLcEMxSSrZlAgNX0FOjH4Xbn6tCTSpu1GEFZR5SmecVuDFmWk/f5fTuR
oT3MXVEpKuoaFGbdZOEyEvEFln+WAgZvP8EGnxsxS/pJx4vz9zJfIs3kIHKCydje
Jvxtfosz+hHXD8w0i7m1nYdHTJErmE3WgmrTG1ggtPFKJNS6YOioBfqpuhmg78mB
d3/VPBKDX1NSk3S17PTZclhuLdcONzpXzJ9CYkli6X/Wn8lDunte+j0sIKuAjDk+
LkMTqJjKdNM0mRz7eaKCFZJGcmsDHW8a6UeB7DggwIevW7g9CdKhsE7pfJun6RT4
ndBuWLtxJXBBd1QGg0qiVNXTneWCl7b27ZpgpqHgKejyyLCF54BHyGpPIIsJhJRj
j5vYAbWgeDr/wm7Q+hnCafnWZWJkiLpVofFe/Jjf1+6B6XopeOrwBPseNZnfu2GC
hLDlG8G4VqeyW27xgiVj8OCFZpWpCtFNgk9tI6MfS28lGg/BljQcIovq6Sn+gc9B
394D78Ri4Qp4j8VXAG+wm6IKWWoF8b9cWYXuUxYbICQMPlKchipJIyZ8urLbyQG1
+rbhFhNh3WoGlXkv5eK+eSQ7dEvKi6PXo3z8O8K59VbkrivaI3x1PoQ7HH3pjU5Y
7MHsvdtxHjs0f+Stb/MfAm/9BlE/6qvMoWRjSseGP1lKEtRgaAC2BEKmXIYvVI2u
IyETaTKVOd3iuuJhhJnSzJ9lsbk3dNxgpCgn0KZitZzbf2BItQk/3vRHm+M7CCTo
1xYWVsm6fAN/OCPsS0VttSSPFfvxpDkyqcsb3MiTZUTAYUquK3/mir+jNX8VGdTw
40QE8Uap1aL3PvQZP+Lmqj83kCyK5HCKWtiFrJ+zcVTL93PVJ/TL0fzVWOx16cDc
mRA4sCSuGU5PggT7EL2/o8qxAIqZFP4zICfw39FwBvRJ5YZV+HAIQIj2rkhBYED0
VwCYkE2kNy9R2CgHsyHDD/qrZG7jiqSrBvNXjn12pui9i7u9pD7lLAkg11oPfbcD
2huAe4T1QeJMEfN8zMSfBl7JZEvYQw5CkfdLyAaBLYdZhqgBQhzOa/QuGNtVX5QF
Wf2S18VYrKTbfWHdRPSO0D8QzqEAveNvgdgy4KHto8DwoaozvSew4AXtXIQJmT2V
W0ULSkv9kHdtUDwx6TsYI786gS323PIFtzGM9dDHbwX8qRWph1AipKGX9+eWLMyz
uJAh69OuNpnbrunH0qHB/VkbaG/MPSxxmBkGFyjkjgDFXT8rrHSrt3ZSoTIEmxdN
ffX70YLRzsaNumKiNBahv8lQF07MWsB29I7H6ApYICq1DJLkFuPsmDDeO0nADoOw
6U6EC7/MAVjLatW/qII30x5V69b0zzwL9/5dHt/90ooXarqCKtJ0FC/YejrosgdQ
LG/1VE7Y8/Tyh/AUVQXy2hbaPal8UWtmGuZc3rwZvsRTPGDsPuWi36rq1kKfT+GK
3tTJfM/FOYUu7BarZ8M/j/9OCBnnrYleUJT5L3WoRmLywD4kCHgGEWzXxWGq+x9C
msAyQWcxYGdRPmoA60Abz9JXx2jO9Ip6BFt4AVfFHGLexQVF7pfzPQk/SrQ2BIrn
WECLLkZGgP09oSrLMmx0xGkXPqXzAErnyDkaD6GEPSy3+ed8znb8biI0scaZwCat
QN2I9kRMvIuDCu1lI6vOv2ySR+Mt04JOAerTcnv8cHMDkcF8n9Ia4ImYnGukvmY7
z4i/rbv0FWbx3yxfeAWYn4WwAP+UXq0w7cVWpijYPIm4UpuAdCkcmiUVoJYW961m
r1R0GAvPjJZK7Noj758sydzk/4V3cUZMmrxG1PYPaZpxCh0GubmANCiwBpT3Qqer
SWoPTSi3bx6Z//B4qNtrGLAhLzScfOrDEIiJIvN47FUIHjJdBGNwdyUsLwoUc5r0
p54Pm09FmEPIVICQYRJCMsbGQZ+kWD84ehTfgLeF2YZ9xhj5uv5jOB6DvdS7PJvS
+aYJnTwBvy1SFPyU4LtVXJ1CdlCrjOJfBmkxqux5XGZkQJx+pnRIk4wc2KpC3UKN
2rJuzag4sYceWk5Xo8FkfaeR5bXB5Z/4KFYp4O3goouD0zdzUC5sQzc7c0lKz0bq
D5QSysQneXLzoAosq9RCmLbmH4am5FD5jNtRv0R96zIF5PFoK98SW4gfO+LD9Hdl
XXLH7A3GS+AT13cmFqX+zOJiPDugA7I8DDSNDEX1OZum46TYebKuYVtJX0o1mNFX
J/XhkuMFkq3IyZsW2gk6sc+gul3D2PKZzxkl6E3nRtyBZbHQrPeGmtNMBCsTyETu
wxVrRGvaWLWcN2Em975drE4XwxmoAQ5h4wKmdnkUxaOgtwX/BYDPsSWwlkdEAGfr
SN84vAdIxLxPLIepNQsXlxpJ0D8/H5fmEBNb7BAePErdA7tXH6iFkFkAygpu9PTW
6EGDpgOLsVR5vCmiML75yTuWwUSsLrSBomWBlu+kLlfThIM2ad0Q4+64D4yK1j6/
Q2IPCgHDF2rOcPBHgqwKOv5rvc2MPgNEvuSbhFEStuJWunDmzJcPb8vDL1xXQRbl
0npdSYeI2+3wpNUQGxKW37ameDXne0y36lvEoIrTxeiRY+cTsxlpTdyhtlFPEho5
QPEPTjuRsvgqJsiKewJmLZDPQTtp37MTSNiF4Wt35sk5Q9RL1kTZj25BlYzbIMKa
mlDsRQEGj+yYj6toJTf9feeCmdSRLqPB5cY8ahj7YyOSoPPWTGa7S3EScfld7joi
6MnFZkpW6M36CWGv+hUkN+dkF51F1piov7K2S88821ogkh0ICbdv2LsiIvI5QWhi
RMgekfGXN/Nz7vHzJJrbaBBJxcleeknZQupu9XipDvMwcEDfZWTBn1Ubzq0STgnR
MQWfvvtJ+S5VqoGD2XNWcnJ7t+SrTJSv8smb8DgnYS3p1O2AVk4whDX/0OS7Wt+1
GOLSr/W+qhgmuni5kq6WCVnO61C4lVpJwfzCdj5RHlA2e2NtsKFHAeKiB5D46wH1
PH8ttWf5ZIOW7daB45cDQH7M0gwD4o/8s0XwAClXeK2fVLgdC9UpAlITTepPiOVg
LHrcJwqxyQwhg8OGqzeNWai+P6hyhQiduFvNsBppNVUAHyBJeJ++fcICC/GRHRDl
c76uWcTP4RpDYyB252Y6o7tFX1kK7Hgkec5es1QMiBl/p38kaErkSajBUimAZ0Nv
rGOwELDh4jtUSRDyY/ndgtLIhqFDL9wAz07Lhh0fX4agMSbnr1XHF2mqKhDaOz1K
VM/+Hqu0lbXd0kIddCC0RV7CtgiqGvBKQ9PiNSrvhAEcZYtCyah9eaiGfGYGhk84
kaB778I+kiGvtp41DHpGCiU6vny8UL2JHD1V9GHadmftC2o7z0VGW7HHLJjd5F5b
KA837A+SRuVQBdxbAfWCQt5lnhKajF5IgxIHveE27H9YLtk8nU5SVsWE6inrI6Cy
Ysf73fVhXeUiu9YrbhwtgwdCHff2nIT3hgJbJx19huhfIwcc6DZfH+rV38+Xjk29
sEj0hYped7CqUngMkq8DCqGZrzgK/6gg2i4SACsAovtDUup07z0PtPvxx9M0De9G
eRXjwTOgDfiwoIAdrBS68umk6eY378xrgsoQE1GqeooAge6WGhfH0jRLOqqDDPoI
lIXat7nis7ZuRWT/oolTx9HTlInZsNBUevFL2rKOFFtXuUl0KBbLaP2T9R7N7X7D
GLjFMxQjJKGu3chB9Iqjp/ALFWIzfdmBVQK3GHzCRceoSGLlVYAhFGarXOhs8PkZ
VW2FDAA5Py8SZfl0tLa0vKSp3Pvqb76uY1HvytwDvPBtjRSKEaoF+OHYaVaf3GzT
MEWHGMeBOawfTo2cz3q3rccxiVET4j0ffg3cKktPOKGDjdc8F4M9LuWcrQc/lRTl
91RTXk/goY3RfuW7IrIh6SiQcXnK7w86Oh+85CcDy1tlFp5XbcOzTL6xRjyMDK+p
WF3ev0p3zic+WYJpKtCuVCR9kf84Iz+aqNb5TZEAVj9uNslNIPDUnxOpcy/ebf5f
2CfVQgrxSlvotVTPzuz9Vqv1RR+91tJYmtr6fRgXqdnSpyZ9NDhv2jKpPC+hjW3e
LqYolhCMfSIRxelrKTXv0SDBehZmwQirVCvz4DjLooTpGk8ipPgtlTOB0YYrd325
yvkrdpVuXV4BztlZ6PYtvXc2Xo1Uw6UWPSAwkBhEcFBkUJuGAyXbpW5X+T7nWOkr
rsKBMu8Pv0LECTRDYsitjhYA/ZxHKz7FlRBZY2ixyWV49SAVQyPeqZlbF8pWrqGG
LqMit0lhcm3URKA+Dm7Q636+p6EL0CiW+sQB6syshG1fwFGYBsQmXj0JU5TArkVJ
6+vSghSbs8p5mFu+SHPmibx6hhyhekDOfXKXsxjZOI4p1UrPTwbXYifNr1mJ8cqc
a55VHBJOTDodGUUvq/i+OyBMn/ndZfFgrdIXsdkDTwpxsCOZ28d0vMLGtDamGQB0
AhWTYTDP8P1nVI2ITHYdanrIuHkGrc2n1UXUR4QGkla2GzjLKZAuam8KeOl2Crc9
ICqS3ysKz+eaAYr7aLi/BBLADx2DZjrbu6TAyDeD1mxAOOG22nG8K9Om4ZUBQlAl
StP3WE7c+TTMTbRTQgf8KeS7Gpnn2SL/KS6sTLtc8ikWhSmFaEK3dHnTo3r07RpQ
hf76MtiDOa7MI/9UwOXZoELnBeE/WeOT0gOGmMn9XHP0QIHxfJHYaC7bQIiOFAlw
t0YRCbsCCEDsoeQUpIYtUfdLtAdbaOI+L4OIQ3jJmhY+U+qdHdkaZ5bwYoZ9XuJJ
U00CmP97sCjyLIEt7kV9IynstSgpSHAngk+jzzK2Ngg7TsgiHmBbfiQ/Cl08jSI1
i8g2ZoWc9YFBPlcyrsMaGZFx7PzgGEHdD0A5N2mal2oqF22B4DYxNRu/CdW+duE7
fSO7tiyol53dzsX1ebkHoa4K+dBFV8EEJH+dLWdkRveAx5RYvbupbTwnnH1FnFlg
icb30JTb7+4ssphkcQVUkHkHVN1n4GK4VX4mooP6eQiHDVK+YiS8X7tgJesA+63L
tqs63/5xToS0tmKgi384eAnyYJ1Vsi9svyR1APNYIMfAsEqzz26I4OGUVT5T2+Ec
WJa9AW442tcHwQyi0RTaHTB6OqFg3dUJr//xr1DmvfIJpyHFN6S1apZCdC21hzjW
XMsGviFFlfkM2re00BOWxBM5owz7+LXbDmmRvvxfRmH8A5JGClXXRGXi18GaFczT
wpGD78n3eWmWRHfTU43AVb69LFEstQhAiQbz3p03TrmVXtdHSddbDdZnHiyby0X4
Y/NLIgG+kO2UnyeZ5OwfzxR2lSXYExqLd6gI5uJDBkq2oKFD6QO01CdJ1/RwstqG
x+sU+oPvm0bmThIYVXRrBlsmec3K0CKtER0g5uECYCm5RCnrhjAuWD/T4BOIJyMf
fPpYK2Zm+RwBUjB2sNoj8MWGFOOHOX2Y594cFXRQECufAPjZEwwIbLIXfD6wOwR4
FSI4YS+quoYxH6/ipsD6i0ogfS/Rmoxr6Ffos8W5MfY8+a4ITwzp8fg+bTg22AC7
FuHsZTJIVTyrLfYnrrPoV73YkKiedOo5gaL9j4mxB1bpRWV2qEZlzak5pgKqh2oS
IhjPvKejum3MgaqaVyVk1j5HVA5JDZrAV34errGFJ2ZPflicEidb8bndj1cwkv6a
veox+WfM6migC7gGjN8dpzcopzRxYTobIPf44af2Sa8Y/hkqRR+Edw5foJ/OR9Kh
Dt61r830BUBEmkcjKPStsHpvS18ieH6QThDG8uQyYK6pNt264f2VZBVjQvuyzSaj
PsofmoTJT1gG2oUco1R9QaTVmkUfNYQ/QEBTp2myOfM9VbZb8mTk1qmncsgReD7O
ZTpCJ/1EGxFaSQ208VLYjlwOLXb7RYfqE8S41JdruiTJQJcrcijFUJp0TIfak8Hx
Fj4wUXfipZxicvQeAVjgY5aFFIzMERtODU5bEbFCG9DySjb2w/XLypkTifWXI410
BbP5rcBaI6iHTILEd8MOI8rE8QT194UNUWoUwwgghZzARLVqZvoUftyeHRLJSApH
c27AwzsNNPQUUfuNWY9tAEv693jk6mywTbARYBft+jR9UXDkDKdOpDMr1N0NHoLc
AwqpaVmsqzm1L8m+SvPB4+pXdoOTkd22RJnvOs0BQ0gccKKK4SdCXFB6uDtFxpAj
GnNi3+P5irJKY/TWHGKcEk/7waagGukBpxn31S/8ACoKS4rBM/fLqaYpu65wvEZ8
lFagWL2PPxd0rGo46irO30qGcw6uKJaZn1LXJGdZGYf/YMEbGnwn/Dt/SMEcboO1
9Yiw5DNGhENuWLLtoz3LIJUGeqBhnScCsFM8TCqUItIVmFUBzaNdece59Ix0hDWV
xUlAOr2/sA0U3FboeJkvalf1y2ukzvMr6ZKq9pbWJ6tZ/KErfWk1/2GGwn7rwkzE
F+uwA63nqV3WZ6fyGXACZnHvJhCk/ki/B5C2EzJ/NHUB2+wjXWP+dgNmf+bZr3HL
yF03jEmAUmD51IUPl15hK3C8ZKt6QgOFaJR2cNNZyCpZIbEU5m53t8B/2sxDfdHb
oDw+zj2thu787QJFocS52Q1Mofm+KUo+s8zfiuL5ZNFssCnm5wk2UYlV5O1hKyo4
JzLf5EUBzin0dLlvn702WS1/24nzd2q7tcpcyDeeXbiOYA9QrwuySZMuO9rtZY0s
WAw6v69aKMAhcT9C6HNjF0tF2ZxwEe10s4gylXdwsNiXFaTLaZTx/NMII8Fz6Llo
fMiU2wcPc8kyuUehuqkyRxYacHzXSAJmvpj+EmZrqdsuUrU1K1iVuSlwmv79DvL+
V1d/uAH/j6CiYrgpfkvKCNKnh1MXAIiBTwfQYCCKnv8Y360h7FZCyNzCDLeL4q4/
x9O0Xe7eky5+Y2onPKh7A6sM9Q5AVmM1RM+XR/HDNL3jnheE/kg+ucpAEtUCI0P+
SsvA3v/oLug7wVqzvPLd8oBVmP2gYn+//qxoEVe13YZX6jW0QUgGL6HJyDRWkUQo
WYM9jmJMnKV6bcInrTA+WayHhoDi3sFhBHsBRGfEWl84mKpCK6SeH3u4KeXRWZpV
BrbIKIAx2tHBrPHYKZFTY0uYNhEFFADX5INSK/5dySVjBqvW/1/OdUl3CT09V9dt
LbLJHjCW+WHofUnj4uFtX6pPyHFx8f5ER87B5VPdvNR56vXSOG8QEQuflOAYBUUp
/VWJi5U2vnrHJUmu4copr2/EU7q5d6Zj1ptDJoVvJmVVUV/pJOZUl0rhPHziNDhM
A8NVRTwUawtLTwrV9+XRcUel/SZ4aKM8V2WY+10/IikcQY2HpKRC27LNCGRhBMFS
z29mQNcI8mXciqKCvCferkJm2rNFh9zF0EvHv354+uuhg5j+VMMiyxo+1oZYaIPB
peKnCeR5T1YmPz0m3mtpGm4yGMOE5zcaErB9U4IxVg0xbU0o4bEbIDe4KjBW5k34
RhxHmLeJGWfcFnP1uSDTti8Vn14ygPuAeij2zRSZYyw7Zlhe/OFjSlquAlGpI+uN
i4amGhXJNfiGUF1us8joZzoi3D3uAiB3aVmM1zxRD8B8NmbvP9eL8BUnx8bAvJjY
gNl/1ZKGvm7rrmEGttfiX5nTF8Moof8qlcfs4Q8bZvMWwhAW+UJ4Ycm5oD6WErtq
e2D2rDv8ImZcW+s2DNW0SGAp+KSGGTy6MndWdh3ByM0oUr4dKgLrpAgWgi2f+eCq
csZCSh45J3FqUfiF8l58srFpTrTgWcUfQJfmb0I8OrTmjPZSTd+ubcmxnCoWbxxb
dajxUli6NYiTczLwF9YyiSQG0+nFKSOGjdhn2v2NXPnDRF6zm7bJg56OWcD6PLx9
MbppNEBfaDOBRXrPHXkIOOf1MhsDw4ckBj611lA++ZjvvLa46wy4pWL4BAPvcA4R
fBFP0HandLeevBSVVGjHTytJKJbvTFJ5UDmzYJHtAgYyQR7CiCkopjMiF+iJAQ/y
gpsGGL33HfCpo9o6z4FrkuGffR5K3Y+UnK6lTgVOULyEMgMinzvhunZwSU3yfDmG
a7FVLN9cEcfNpYfBAqvYjJZEetfAOEQO1TBSsLjNnRUAiMkCo6J5bxdpX8RmPsds
JMYoNjsi+wDxoKjWgCebq0Z1Yo8g7iIwPBuGB7skA9CBJ6F1H7t/VRPgNebeP6P2
IwwcvtdfNx16Oht0+x2xvPnlrmlZbojtgPKP+6V0e1yr4njBxOjNNu8IcOiXw746
2LV1BZitosCuEJOoyTSMrjUPUlo1q3VZDVDhFSz+kTUWdjiMnJw/wY+de24opf8o
jO0b8Za5pxjoQ9RvYLZQ80UsOBGEpGYOSMuIPvcSrwq/j63cG4THdr90mvCnby+H
/J4UGiZkvoD7Qzg6ItIWiDBt5FFxdCM4Yhg5swuBBWtnlbfzqeMSHEsPtsm+zGnW
uVHzmgrGpSb/5JzTwIG8J1Qa7hxcFL2IFFbw0iDF6ky5ROUQDNfMFv73VIsuiwHl
TYwZPNqnOcr1f4jdRcvE1p46ruzwjuRrP6X2rQsDU/7SL2J7q00YjxlTU6xwwlBz
7GoxjUCtMjcgtvWFDeQUtWht+c5/BeJPlU7Ifj+HDJGA7SygUlKymFykEdbhpNGZ
pfowqc85w/AsZIS3aoMgrLXYvHY11T0aT98S+lY9/qvHNNpyO8eXZ1NyK0brgf5/
K5j9HwwzTfpRzxr9xOI6shiD+XiyVSvgJ25N8COZkS7G8ZiTumI8zFeffE5I3aVU
tUyMQAD0z2j7yDixUqlI2yxY82pruHBydSUfSZStQWuMPsPqVe/3JGxTXrcCNXhG
+7asdlf+qQ9LewWNv6sIWhhVr3KK8awfw5264QFhhdPjeOYNIS6IpETJfegmfOpM
I+znUGZnTFk+HCjsz9FeVaajCzvpoHFr+sn5pRuurUuVIuRZh9ZWgfzD9XUvk9Rc
lV9qT5+XaYmkp6CGi8xeOj4MvKyseOR2Tj4xjhlsUtCc+lnlVu81j62B0Eez6xVb
zCWgldlqB1WdVrLdtyg/oxk1vsCde1f+RJBtBXQaplcIwGaBPrtYAE4fRal4Iat8
GeeJ8W0vLGulqglkIzKjQ9Xlm2AF39KGjKXOA1XtyICjQ9iD4Kb1oQObnLtzco1p
yuvQdr55vjA6V3YU6z+eNCXWZYxvUj1kfdZrQ1KnsKfUcOiXvTSKhaxjPSY6HHx3
ikLy2/iFOFlz1ED6LREp/mqPokYTnld1rYVdp577K8ZhAqAxdII8hm55tyJrL/oB
W/viDGWKttXcmOlXapBFQh7rJVldvETRmFVax9JD5eHQQhBS2pCBuyP7ryEh9Tzp
gdsWn8szSe/ipntUzGmKg3YSl2/uwF9d+11/tYISosFG3qGdsz3IvKX0aetWIU7e
I8rQjF3OVBlPS7DnJyAyHl1WxYIRyjMFQMfwnV/7MoltZ3cdoEO+fad+tLQOnQiR
GozO5goI/uXxjMnWb58VL57DZ8FC8ElRihdxoDIluPEgmgFHijFhDflj8vfhCXke
s4VS5m37uHyG99YeTgvxuXktgQjZmBm6SuWCTxMm1nxfMkF3SokT2KDYONk0vZ99
5fKkeMo+Md9PeeXV4yvMl7kKKbqpWkoCs55UIHpvqFukkt2etC8620OzoHE1gIPO
ToIR+kKI3RtdF8O2zDgtGGiHPxWy+MIgAEVtQOBbfmlvGGOVIuqmIZucEPJpvZ4e
7kguCpDCzB5amI/bf41XnVeafyx6OciYSTfRrWCHzjpKd63nUgBvg5tIjgF9Jau3
T1hKkv3tB6jTFBHvfWRNTbe20hWyAP59mx8UqRsPxAc1idKzR2CLO3ux4lJQD3w/
10ypfpxkEtL6B3citS76TfKCSfN2yapcoCuFSaqZ42yg46InB67MIB6m3UiWbmqq
E5iRs45Fr62Sn+iii+pGd9Dd5tjvYNKyQpEmN7h+zUFJXlAxxsn6JEiKbowEOYAZ
GpUVc66YvZDjFYpKStukgfLmSdr9tWaqe/IBV211An3/3DiLsE14DB3kamHGKKi3
jpxloukrgcezmFqoPMt8r7b51fxZjeytJ+JkikB6TxsPeKeoPaWmP1foEkX98Caq
lzOkRqJ/5XokY38FUnqLbTuHi+DFM1PZVJdvMqR4NGSYgYoLBWV+G4ybKZwXvyMP
+NQw/b+I0hElHzlbDSHkcJ6RkascspAuIQhsg78gWmpBBe9OfMG/tSppSKslZOu6
pj17taax85uSILr0hgxtsqTaYcPtsqji/DbScnAYGvqjGW9lF6+JlwD4xjoDUXNZ
Vt/62OAhh0nHzldb/b/OXzkKNb5q9+IKRXCyqJa6VMFmZwCGSgRxRr/6ke4gaNDa
Syc8wbtVP/TYD0Gjowu7cyCny+klQpu8WKI6LqlV9UFqSnLVJ2SjFnzHxgG5kSvU
KnRyY27r/ZIUnnK2jVnj9l+ekvLZEt/YhSGGpreNWr4Am1aUHPIwtn9zxz4aVJgf
j1+VqVnWVPRtycZAqZ5oOLNzVtbsOIpWbMG2cC7ocykmxzVbKS0Adxk5FNYDkfdh
QZpj965I6R8BMIpAjvcgM24pgcLBIUntqLJm/x+zdiEc/fN5ZPqZfF65hPIOOzi4
OO+enMXLHaN7spby/QB/jwwksMcZxW+XmEBNv9MqDlzLMzrN2x8EmZyTUDSjtogp
mGxcBEp7oJaZUNUF+iEStX04mm1lX9N5Yf3lFM/xcg1JOhx+c1Jj6uTZxASI6Di2
hb7fHKs7EdoS0g76JYd+cOOLx0IVqs2BaBq18hrdPWVo5fLiSFE9Y/UJwgfUEuDv
QGP3wcQS6FTN4peQeo+xqng3nTU6SSHcyVqtrC/AF6mC1tgOPIG0fOcI9+Do+VuN
I2icY0Ap51Uty6lP+R9nU14GfZ8pfwDtz9ouhlfj5KkM/SPwP4jpCikpjOzn9TGz
3saCg3nKpXu77lXktr+32vxgjKann9kLL6VNbCiDYYg+E3QQTmQldWsX3TLqYAEU
NhHDAv2RLR3xIQSIj/x4RD5vFvBsUUZgvuXwIBUn2kw4cQdujAQa/WfCC7prFo9m
cnyuos/Hq/BQUwwU9N4Af4o6Rb6dXD813eiq56yrj4vL6TfixnA9qtLRgrU6mKlC
7mkE4HAXQsra8dI7YEmRb5L6tz6aZ50Al/mlebn4m3u9OzdhuUYgJ6FxSCjD74Ql
yur8lIFicacyik3zcjHJzylYWfcFs8o+dJGRcCCXCrZbRGbHx5T7WHKJJ2+2FIBZ
6IC9/ddTWGiOf8eMK2kRGQ9Tfkd8323to4axqOt6lE+wpLfbPx+pemXmjXlzlcGp
3hS2iE4ij1pfZe0oYQSs8VobyyDFTtWoanEpgMSHcUeM+yFCIxSYuAp3wb9wfgu7
Jg84NtF9RLic2nD429wNYvYYyEYv+WWwUZ9nTLqJUra2FL8GlPz4DvbtQ5GlHSkT
kqbhoolMizzzKN2l19/HQspxEMWUuIydxvpnsG+8LBonZWou+rk5jR6Y7QQxLLdf
NbXPY74zXWDiXKbUxm3MCO8TXo4rcrzod3LWarGouZybctiBuyhYtHbzJh2DX8R1
RV+z23nD0c7ZYe3qiA9JyTJTbAHZXNt9MFJfUdSLsmEga/unYuewo8i6tCbn9jq0
6gn7o9hpMks0SV7Mm1pNqcJ/O4dIwA+ORmpULhmHilnVa6uHTG+DgUeUDZZGnkN/
DD+TtNfpmExyEpXzsfHBiSH3+Rfhq1C+PgDL8yyOf0Pb5znwUKy9rQxaqu2p4EV/
dQqr4WNN3u1sNQMlbrxYCDAwwYTU/Hd4jWCW/ZtE6t/lBZWmc7UQ0++rPa375ng+
3HKhmyeFg0jeOdrDzR2kbeUEXDKxZmetmuFRbhX0Y1ueoUVBCTQEcrYgZcwDsoqx
uanrfKUQNEe9DSppmfAy8ymd5ezUpu0WcHbm9JPJWG0+TT87Jrq5lc2mqn0uXsp1
30KnLSSK1SQbcvCp6GW1xTZntmFKUJVFLBaVdC1KXLo8x1X5HvPhtxh/T9N8fJ/t
8ZK9UPq0VHDZiFAmQsdqKdd99+qdP0kt3oDLChIGAJM2DgEeqIb/oa1PkE79LJbV
ui+2EkzPYt/E7OUXvTNDNPHR3hqQ9bzdEfv9rfCtP6ZdowVPWaXYGOhILMeF9Gc8
VWU+bKHfK5itJAXRfb56EMSUWP/cxZgqbmWZK7Qb1INENlwtBi7NTI+jlv1t5snv
3qLtnAysV6whPF9oK7BG7F/psZCFruABf09CYLu12upqrKmHf9JNZCz5NaFW8bJ4
ybBXTr6DlnMiDytqmSSXM5Sy83RAPpt/LWExnKpPy0jq7sI5HGM9AXWAbI79P9Ki
0gpr39yE9KPm1Wlv2lJHIq/tF64/agG1dxq6oLV61CfnEXtDS7LvzJfKLZeAJGGF
/pcUm6/895fPTWKWYRnA6Tiq73w+l3r/k2hG1VVg0lT8tlbk/EVckQVtB7XQPkGr
int6NY6D8n0aWGJDWhEnFOlkCc0poOWpcGy/u7NushApkFa8pe0o1SilB1M5MZvS
4zg+dL3XX98VWA7j022g7r9S80JTFPzL2P74NJq2fytImpbeGbKwjlxtCsPzXZ2K
Rsva58HDks7EJM8UONcMlS143gDehQxYfhnQtXm5MGvwa8FXLXWe6g6xRIwuxBCL
P7u+EQbW1uhkDt85zHscEjc+5raj7x305ngr9yX8OyXCIltAmmWHFcWVzjSbFLj0
qYWnkaI4kgB0rZPUnkbRuEn87ceppQFSS+KmeWCTA6mLDNo5aq5b+cDhXK0n3lQa
yc9M98mj1zXH5qttpxPZikomlpANdzQhUOq6GlSYwkt5qWOocKjVRsjMmxZG6NBJ
7YILJFdqxVeHjBP0etYvkNDff+3XlUKty8euR5A5nZxlxdNTMbTRwmXSGhpy0zxh
JJAj0DMiHFVndQI5TOntAot5+Hk2hjqYAoqFdmj9H3kQP04piKksb4ifZA32nwMb
oh6wbC6/AeR7Xi3M7z0VPvS82XY6MiEc2TGeL28dZBxxul79pKKRoRcFneJbWU7U
Yb22C2byNs54fRZlzPbZQ+ZSU51vHUSI8H1QoZvW0cLGVmxOQpAAQaS1Y2mhpDVa
ts0tZOENlh0RukLa/hipyAdgIS6f5J8IidAtVZS1TH7m/9pIwZ74ETYkvNZrTJen
lQajuspMRLO0pixNpRXO6FR8yYuLrVwJ/Xcr7/4SmZX2MqD+knIVgMiqA/yP92lJ
YUph4lR5RfCStDfrednGdFk9twQNTbGiSdntrzqOn6AcEj5ATI86QPFbBzf9twJm
iiEDy7arHf0eYFqesx0ZPCqkrRGEiqoe6Rg/XgVoL/fWDh0IF3WpYtd3FxrO26ap
3XqDiSAylPAu9O2/Rahuv8JJ2snq9/Ysp3bfC7zq4ISZ32S9LQY4CHKxq54HyNlU
0exB/7gQF92Fqekoj/giiukWwgcasSuaGmjO9tcD85vqK1Vgw7vh+v87gM2LEKhW
E2flFnRe7sWPz401gQDaCwrBo6LZ28ZfUJ1MAg6f30Qb+e5je/DZPTRyRqJvdHyi
tnWTKBLZ+9MNBxfp2/04vL8KDbKBWF7NB0fLQ5Gh9142tjA2allDBXEFw+uG3O2P
hjZ4PzuzUN2veyUQAYpvCS9BdXdHh0EnBkYOvkQyLCFLbxmVMc7uMv/bel0FJHzc
bKyoA7/EKZIy2JM0ooc5WhmwKGK9eAeOW6JcCrIbOg4800r5iJt5qKDhAwV/rTIP
n5ApV9SnBxRce+dYJylwq2SF7kav/glBk+3b2ittADsDQG3YJ0cHzp+cRyTXNkaD
44ADmD8X/vpnz3mfle8DoFx2xQ8U6bP8vAuYBBiQLJqm62NpkSfWZEV4YIzIY2m9
HPmGum7q2dUHYrz4pE/fyzfWyAFnxI7qLgQL2oE05ENERrpflXD9+bSd9RKDFgpo
ZSsOWjb7UIunh28L3xrEnka8DBClurkBoU2w8XWXgxAoMCc4JhO/jg2dwP/Uu6ga
KWgIrTM92m7li9i03S8DUeuUqXIFaKSI0U/+G5ruOSJJ2UurpJX1febvBGKslYvX
J7vXPNT2HMNfhjxhF04B9Fq86d29fbB89b775x9/sz4xViX1hvza5mjW6NVYvxUQ
b4bw1uWZ3NDTnMlNZYIRQ65pzdoq1LzN5EwRBI41fh6woS9hrUGjFKBlyjaEuZ2d
/aTcMdXy0zrrCHtv32Dx4YoT41/gTZh04hobs6q6cCSw0HQi3nVKQWjRARcdxbjj
OnGgyDbcQ68rE2zJx3OH+wrGqzWRqpDRCJwTdMjyQRo2Z7USBq+qfEFaC50NaNY2
X5ZY4X1fzpSlc06WtrkXVWBvXkq2FdnJ53C2V9y1W9sTvH1ROIEXbYT0jHyFjbMA
vRR8A4UWGfTMP2NSLugUqCq9Rgs301wZyVSLda6REwQOzsVstAj71Sr26azbpCd5
oLf6Mz9IEckIcVa2hS2GaJ9L7lWnF48qkFxesK7oWsdRJNtirRnaMA2Yprpcu66G
zT6YcJXNrWYzIr3MOLkQb5wUXQZ0roB1yH4zuYtI/r1YKd01dlGaq9PqtT/VouLQ
UKeE1R606SQjzpsZdvAy5WbAMxwXUlDy6gNDpLcngcv7z57ZAVZNFhSprP94IGcW
m1hLMQfwpoMwbUSyapYltnw4QI/oXpZPkx0jBNhTU5Pus+YV74svUC0EEOdhcATk
Yt5txc9TDD5cl3F0Zfk6pZ+vfGQyBXykwwM2ZPcXlP/bZ392GNtraNP/aTZy3JuX
Ykl3ruN/iEj82ldBP0KWJZy0YiG8inT6xpJsGkD3ikJaZjvXPJ75f06uyU0p7t+o
tU4RvXksN+/aOStvknTkhw15LnARZje3I0W3sUF/bVczw7l7SRoNXfjkHxbxlx/9
e+1BG47XOFQXrLVsEYiAzdvYhwbE/ggNnixLv9ZQsg69ZQgOJfiRAPR5ZAXxtWIq
efQ2DHVGSHt73F+QihWdhaMxAThfKaff8uMvHVP6una46xsevzEVHrUpYRAtEwcj
UMEBTIndgLyzmQXiHQUlPakERyWV1KCiYTSjQ1teUKFPgYTMFCBwGkMDuLrWJu8v
IcYkaVJx8aTnPDiPB8L3CL+AJ4gqIATuvfXWMNJZgCvSHgRcV7+BU1+Mc9XXQLQH
Y5dtSljHeB4ESidQH4wJBbVN40HnFxmft5x4X/e1n9yZ0/152jdyqXV595EHNjpC
369F/46P0w5ym3LXghK9wD6NrJXU/NANttcw6Z7jwLa/fzfE7+kpAlo3U2g5fYQK
vFDRV8ApJf1dH4EII7gi29sVEn17SwwGcjc6Mm8UBoQuxAAqtqq8EfNt03vkTKbt
KvPqSzIwUuirQq33MiyPK7RzarNvq/thxg3dxYwk8VvL6SWPaTpeC00lpqksPXZu
8SfU0Ye35ceXK4LUU2eV8KrtcH0m9ecMc7c/IciwdnB3Gj5/ZwGTsplr1OzWGhfz
8PXJMC6DNZLAVKiZvnpjD2M0wq/crXBzpYDC0jgS7ZI+ZEqVpk4IiwF/9fD3d6Lg
ZU7OQxmMw4BtSKRCSzL5E9NvGOUAGCx2o+PkBDuuNfGIgVNLp5Yv9EhveE+GlDbO
DIl0GzrNhgI8m4NBivOfgD4RcYAZiYm4Xt2o4FlHLyGIRrMlGhGvcoPcy3xi4asy
lAkGPEdIZU0g7Gln20SGB/fNEvmuR2M/k4WIDMMgI64zi/IRTGUTXReCoO6fm7Ru
vBjQb3tigNepfirbZghUVcFIWyOuykusmDwDNwxZnSM3+VwtjTrTZwVptNbNXz+W
Gy3VegnJQVB5PhukWi2FtyZugZtDzG3aH4SRlFrH53tttGQF1In9PGOlrgaL6Mfk
VMyxac9oZRBgC9FlDGaL1PX812OuRhofhP0aA8n4aNfl4qVAhS1PifofzEosjgwY
l4ISAxotLbQbFDqZ0eq3hv3g/r8akdsahuaWl9o8OVHEFMZ4qo9lxslyIfijZ3d5
uBnbTppfU5/ZADzPrNM94ZyQb7dmGIlta7oyqlOqDpmbN4gGb7UHPDjErIGzykKB
HAz0GSYQN5UltBqYchmSdLI7v2EXIjs+KJuw30Sy4m7KhZdWzq23wjqhwRptJiGb
RrhOBlzM40AePN/aBda95HmhsBVejEp3wtGEtKunWZZFpzd6DdveGbD2tHQ+Uqd/
BAVghXjmVubxc2mfmAf2gvPmEg9NI6HKbREAyo1u/MhWhcOnQQvTHsFnRM2AOUzB
dAbpTvc0M7fgIYQ2zv0A2C80qTnyyhN2nykbCZ2Fptq0HYK2fcBdg674cNQ/ZtX+
hZheOXz+TH0jQ4F26cZh3F5froW81JKfoCkqsIA3u3XKPvuZgVCrq+24DicfQkMg
oUz4qXVHWn1Dp2Me7y3f1B1JV8aLynEWpObtxYzLSZaDg4hlPkPXYHHQgz6eNx5r
s+PGbzNU5sv/Thv/JjbiDgMcJ+i9iNoIG7dKniArdreNaKNbLmyYGlBfbExWuKED
0eaLV9gA5JosijT/8bY5R/Cx5M8zWcqJ3BNdkuUV7D3Pauao3el7X4p+yIg9FJSX
IhqkpuNFQ7kY9r///0puo/uLnwZCHNShu64BfNc5XMg2qcIUp1yuZVOscJEMsM3h
yV5GgtCvBkPypn8JsLoi0tD9ldtUdQpmT1pYO1Q8jRXDOzdrNVjXKsMfR+SM2MnI
w2VyJSM/7Jb4Bqd8fDO8HZqPPRegX5icJ8WWgS65ngbxqYisti3Uu04/ptEsCUR8
oSaAUoYK458Shl2gZcH5ZXsHvxMp/xxo1fgqnclE39snOPQkxgytstdzKqgYN2+2
g9C13+ZYaouIJPi7gX/GdIJOP48tl8C31gNFZkEkeN8tn0gD3FEuFyb1EQIHkp4E
9wppPnb2zWj4VHzmi3s3Ia3lsu59rbm7atN6/a/AcVoUsQzqoYp1GWDvocU1KUTB
DvhYRESu4jGT5fx+6na6ooN7PYQgs4St0QV1q5p2mCkYhNG2P48fpicxEAe4rNSe
mbMKfUtjciKh60qc+DVZiH0hJTsulQyVr9GjWA7GDqgh55V1Jgb2zzd5vuZVnB9z
LUBVpktB8S55rKB89Y5qO2yRd9tAx/4RIuPSmU7+Jhn4KAwBG1UGLM5FQjrCxO7i
vxNSGe2KQiVnhw1nAicuAlMKHctqdL4DjHHEsnXT5iD5rsDgUg2QK4y+14zTpxag
E6Bcgaxf9r5sLpInFnObaIYeaKpzmWnS4O6GyKJfjr2c+cpk74phjZUNAizkFdAd
iiv4tAtWMheDfb5l1qUC08FnerU3ZW16DcGeuQ94lvbJgCi0L2ZeE1dc3biajW7a
kUZda+f/2krEYgG3QN0IOpDOUTTxEasThSGruL/HxG8s4B2+4RWRpb4PUAzoQtn/
zITt26twfCG4DJWEg7+dtJyfRfSHDGnkKGNxRXoBLyVyRFkAHHJZbUzNiXk6N3wj
6lVumMdAsF3OB8iz+Tm2xpiqd0vv3SkS3NDhZixGzEfumGMVafGv5t7h2zTr6RNL
SbjPm37bXEgMyu110rkqUogPDvuHhsUwb7NeLFC37yu1ZRA/urnmBwjbIYPFwBIK
xe1iQDph5lLedWcvSUQrdrcnYKg93+pWlXEl7Auet0dy/qh14wPuM5PmCDGgJ57M
IoXVnIyp50YcVpft1KHjCiCF4hyqrdxX+aN9PkhRjKqc3gVN1H39MkfYE8rfQ+kS
1XVTXoHs0MZf9Py3ymlaxUjq15t4hw2HhoMOGxBGWlCUJJRGGf3m83rQrSHNleZ1
V2b8+M1ANenVCPG3cNVR+VOo7gKeV1CnvnlmAXvqNH/6gw2gSx7iZD6m5oOCULSh
XrCvTqGmICBVzQxq4r/OkqnN29aIKymQfQaFNC3ntTwtxlT87ZHblGvHaoW9/3JJ
k+KqrYV9HBTLDK8ztL0GfpVrctWDv44awo5qPQdGalRIWaw7AAQHZKqi7HVXxXBx
MwDgkvMfyv3KPY8NAtGBa95kxEEyXhE+rcAai1gTpg7qPQlVh8TQ0mn1ZGgNWPd5
Py3wudnBrz5YhiZf3+RaAHvxG4Ynk0oM7e8TAHZMFFOGu+jIpmelDb7bfGVH2JIa
02zBK7Ccm1W/SCRURus4nsNow7tH+mQohc6F9ZJ/o4N+5HRPqZ9zobOFh3YUEDE3
UY7BZVQ/Tdp/Y1bMQOqbDyu2npaIdpgPwoCkaQJrnxk48qBiRnab8BqpckOpSspo
ZfAHBY60a0aMkohXvfCd3Yl33BmTFpKTevo0Sg9i0QqrVT/+legRTBwXqqBkT9Mv
JjdcoD/lOxI2mvj1S2rQbl2GsA4XGU75fT0YC8E7YyBb0dxVhY+ziPss+/kslY7/
Toahnjo+iGy52cscX/MfauXRONxX8nx6AqClWEOZhXDo4QJ9JHmwCUUqt4f6cwqo
fHbwSbgQobBo+iw7ZM4CaF0N7hsgEKFUTsWsIvc7fvxi1fRJzTHgjiaw3MXlTmrZ
8ULxki6utd8c+gWREw53fuLIpFqPjT4RvX+N6tD/Yo+ktkXDMJFKe9K2MHa7xZTn
7UbSDeZx6D4cH2MLi26uQe1r15uk4OymKS3quDgE6tVVLKyqcf4/kNiyIM8f+LSG
05OcFaLv+MTDclQy5/Iba7f7X/g9tCx8/YV4CEnrZD794UAEBKptHnzUjw5mOqFe
L35J67HGHTRqw3Zdm8SChxo5Gq0SlbKedxY9Zu+xi6y6wGVCweE/yIQzS3BDWyqY
jQ7qF5nCIWW2iOOVHuE31ne01Ua/n6oZyE0yvi7SBRvKsDTHHHygxBBt2j6JeY8g
1P2nrIORDtYpSyZUqL5rheZa83YXb47MIgqpS64FdHTRtwwsegq2f36O1SFBHG5Q
RYtlFqV0fGlhGP6H2f7ydsQ42n5o7x274uoEg2wzIoXy/lmkxkr0eGvz1FvgPWxu
BNXt9me7YRkzLMC8yMqVO/kq6HuOWwUC9SiRt1EV4ChbUQ8AaqnzO+SsYtPq6cmG
3DXWgImDvUEV/BEFZDTdx5ivmITxm7SjBjp3zsge4oeRtIka99drfQK8kDlRgODe
G5aEi3US/k9itHfQGU/KdBSNuJjcwze3BSwPBwbndcQoIQOPcw5PzgPV74oHQSNo
+GB0KnYaOiv2zJ9W+mE5DPYf3fqr3jaGg8dRUeizC3nxWdlALyCPbYhNwLuI5UGC
sSr2v/XaUtT2RNJCcVc2coeNZi4bLhgJ9EwsZOCKJ2gClkFMiaN7T7na7gG8Eb8R
GYk74IYG65aLPnb/PBRkY40kso8i44gtXweoKXWLDWWaM9/MIEJ36h/4RxXPgZsl
yNHtCHEad7rjxNnl3UNAk6+0HFf9U9Rhv0IOKVk5y7Oaslhy3L+UzrJbmIOk5sG9
Td2j89rQfHwQyPCuLrYRk3HQ/2k/3MC5srrC2WwtYKtElZWDdB6ulOk3qtFlLua4
P9L+9HksTV9yzgcE7PALmQgNGRHvbqgip+1WotH0iQcMdMlFQRFldXkW4l72dEn1
ZRe8D5LUWY5u9fooI+luXAuJpDcFDt9kXs/GrbIulDlLFQB0bbzekc16tAt8UITN
74qo31Znvm1qXdTMNAuLQ+Xz3r25fAwkSrGIQbuQJmRz38AbAqXnRuadPjeSSN8g
2P+Hc16hQrqwHuwNbJLb5K+WVj50gAdLJLcqanBNpjL8Hu32KJW2sUrjeTZldZ/k
7HVB3+ux5Eg6fDXF9UneIiAxDvtFlJv5ZIrI0/wRCZQYtb8mlFnywhTTkaiC7Jz2
qCBj5G7+/1YLdiYyn3vRqU2PUWNMJBGdLrV8mlmEEAEJQs1zK/vGdPcFYc4jdtcU
bRKm+iGc589Kfp8ChCZGSQp5jCgKjwuq0QZD/hFSDOWkTcryWDA5pAljlKrIDxMG
9OaGr4HTlRDnrGU+csby6wGEK7KPJo2CUyLh0C1/e83/ycRT+B146bqjpGprkHMv
P2DseV58GPnK0XgDY1OO2eyUtlAhP0HmbTysTwv0k5otKsf4wrKh29JWSrZQNIrF
r22lVBxqNhqAQNqwbQFeMdN/pNAaozVkPy9f7xmXLVbzocKMFz+BaJIaJGssNvNT
tSXtFvBJPpkLvNmCkRt27WuDUQPnfbjdWcM/Td1QetSlIq2L72ngVPBqI6GeadPP
8YXyi2wmdtOwESI0WTW8049CebZl1/zqWxapCHrnI7ylvcuaro8l0TpuoHUm9iKF
hPwCHgAbRqse+Prnbslr49AlxsWUq43QcJnr6v26BhvzfKD5sPcv/8RmAazc6eTv
YCeviNot3I1PdoGoJyTEHzrBAJTXE4qsibqTFl0Pu30baMEDaOH7Y8HFNRwrmbG0
5qi5FErbI/CRin37Rbbp41qw/3q1BjnhNfFZozUQtf7xoGzVYZRblOpTXmGwoW58
ITw17+1v9Uzvt7f0ueeh7X7MH8mj1c8xzab9oXHIP8bsDWoCDJtzMa5qI1yBxFBS
lOROikHZMT7a3B/Pjp7sxWIgm8Z5U4hsApKxjyRZEz9elTdD1gRzPdBsXGT+pnUQ
6bZ2HmUtwkBstE408683LrLEQXcYk1zwwWdOMWF41Vz66VUx8mZd1jWuXHZvpK2l
XpUDy4nILPQrWdfCkOQNxGFwAy5IcLZcW3jJ2+mxP1pN5WlnL3+gUa7QLul97lO2
RVhI1RXcSJFpLxjvMZehg7vZTefZtXxFf0oR4oHZFCq8DCYZ/L0wx6eWR+ZFc2AT
kjKKMdFYBbHlN3/6tb8Bx5copQjsXMHKtaRzkBwcG2LHXA21aJegmHgqSB4EwaLa
IKFkapjXXdHOTESNU8YcDa2TPIH7IIPUMsil9P3JR6+t2rvy5FhYDhX9t8g6iRcB
inqtM04jEkHl+15t42fsOstFNg0mPSpYPqR9j78JBdbBoCZNVXJPQtRKytm6YBaW
vNn0lkmO+6w3avMvgWyGh3ReQVF8z2YIouTNc0SWd/MXj+FyQKaxv+/wH+bGGUpw
TTOUqAk3Cos2hl0sCEPiB2OfNcolqUVAk/3w6azsy1yK8+SE8SNkDcHK4EsMAinT
UP7jkZdkxTpTR96i7hP1U6/ABdqJthD48kmdIRQlivX1+vurHi7QOAP5s57SbX/J
Xihl3gacdkTSCuHOe7YSP6xRDlXAJkvKsr7wIcv2wjF6C06phWLx3Ci07tCVhZ2I
P+amiVEeLz8lR7Sjck2nvK1dNi/CbaLinDvvOZ4jQJwdOIpuG0V2CFj9JZbvNEfO
ycrBchZwHvdURojRPy+e/gRRFEOtNgCKTz7MhR5NTj+i6jSsmkFbNDRXaB5Ch/FK
cZvkblnOT343FFwRzBv1VYiIMt9jwxH8SeS57qyDZLURuvhQk80pSL6D+tRLbHHd
uNkGwtWhjjoED1VrKro0IyaLE+/lBNDZObsCbmrNVjfb7IQmAL4Adk1fbda+Swxt
HoSf/2GdTt6GDJcDcRRxY0rlYf3iIm+VSDbf2BT4QY5cRKet+9SpjhuNjKzkBNhG
085RHCk2kLSv1Kj265itZsjBerzDFcZ5OxZ3qG5ABZxWw/eHW1V90wQuHuP7Bx55
AmrKf/aH7tsP7egX7a8p8fFRlRXXzhzPfxetb0DeZOnswqFtN71TTjBUn+AIiAD8
AB/cCwfgVqR1M7eRvOvOq+GLs8QNFlhLDNGVPxJ4X8Ativ2yRo+94NDbBUI17zuF
Hk9x34bzaxWZddbn5mVetmpTDqprjnVrui4D2Wxo9QFoaePbM98NEexMCIw6AuAm
5NrgOsGDlpEN1DQl8DnuybVEl9rrOz8WDtnDa9wskyy/JrV0eY8Cn4npyxU5rQpy
wmTSl+qvdi1iTfJP7Fy2kDw/WhLmyV9MUG3e4q5Jba7mZmmwJfGeAqSmRzt1a9sn
5l66H5JF9mVOgZysDgjPCVWbt9dU7BAyt8LAquqISHEcdGt/trOy85o7oycVS65f
VRQLyPfRCcdiakbvx7mrSi0F4OvQjznCOqO3FzwxWZquYyMEBwUVSwmkniM0Rgeh
osqAdGOzp5PTWJzO63wgD6v5ZMEdt09Qq0lCL5loENyB+/euxm9UNsY/SzVdLld9
L6e/lVxqSgOGmMbB+x9fphTj+602KSbgzLhrNDeZPc7of/8GFkxsj9oMcUgOR9xr
5geopTjZnPY1gRNpjq8vIY0ehny/lZrGSpN07UKqz26njPNP0F/HdcvMldpum65+
qY6oCW16E+XkuBExkFONBg9vaZymqMCxIzJSQWUc05xixKoKxPS9PyhrJt9W7ADr
X8l4qcCOQw7vyV+DtaGSLl+8A639eXJcmhmWDsvI6zggW4toyUBIhPSm899FSfs4
tvf4MW3mcGkfPBwG4MJqYoDeuLLpqOoj0j+dNukJehQ9m5NG7Y1M97i1oTq09rLP
CM72x/EqHhsVp/RPo14+RAieHoh+Kg2PJDIjmkwbc/Kf0KjKQYj+Mm9drVRN+Xdc
FtCpodo/rUUS9iggxu6FUzcoxMxA/DpYcX6RRTAOYRfTG5dsJ5oI7yCaaEN6BuuO
vH+zam52fvcVlop3qg09rABo44/DGA01VWPFNkzSPfdvH2yN6obeklEjMtI+ATh2
jLwhLAPx8+69nW+xw/qiwENpMLzOcxss4QPPBYXlCfuqEzGuWO9RZbrrrYk6bqqF
XQ8ALTd4Y8av3vfJlt8T57SBL3juqKhttcNtwT8kiNgojLoyjlRpfxXjYSk41j0T
BgxoPM/nJaxXKTJmLe57Cm29lfEV9+ptFKC0RTpTBHgUkFH+HlGbnUjdVpyf+N5h
GmOhptEqZxVPDfAyS/QNZRhqCyQSsuTNPkkQ8AHQbj5N3pnxYIw9321L6REZD2EP
UeS+ldZfXecHWOG6kE+A3Y0btOT5WEUCR09blBGzp0LViULISZ9N9Kp84PQcfwFf
W+wq21KfBIyzIhKN6V2z+Z6kvK+oL4iOkEABixqHqW2kT8LGrx4k8P8jKiBKpe+/
F7ckj36fYtK4SoOZfMgeYEcim7cvr8Wfz0mYL6/LyFN0okBhdWlPJ7vJ/9mQJKNo
cQGcyfNyTzM6Se+FtDz+XH3jif0ZA9lPTxCUAkl6V5pg7mDZ45HEVJwKbyKNgFcs
N4y1r4r3UJdmGADtflZr653hH6tE9mB+BWaU3D+gGcKdhsrxHij8aDO0p2hb/fMy
/JBBCIzAU9DmbFOIM8K6E747D+SVE2GASYEg6MvjMM3z2FsfRl2v5fYMbKs7uRkX
nzYfi+/nKSb21fPLqYdgkC6lydmeigqLFGZNMObkG836T2Fuk4ThNwH8BBXzDXMJ
A3OL50CTA7DrElws0fS7H7EEb/wJ9x/22yrym/mXqzwFIbIiN+yNAse7ww1kr+Yx
KjZHoqgZn1Ds93sSE9A961u95mAEWJBaIiVMhNnvBcZZanl7gqk7EXqBLYWt/amK
RxiH9/bVsiy+MiwFbbj+Edtppqt11ACZApXtBdEzB3hwOcSF+cR2XYUix+hYVwAe
/iUiTwEctdKUTAlzbNvcvi/dqwiay6op5su0WisuJKLDqNpALzjpg1dKcgKoIa0v
Z63VB45PM9acxPxs8QxSISdGB//nGTrVec+KtN49nVRj2tdaOl7c9aLhaskKeCR4
WbRbJD3KFxg4fQV3ZyrpzaO2LiiuFBU7tZ4NI5Wn+xSzhPUf/AxSGNAcXvw3c0Ow
fdupuQSKGznQEWeSMg+E5F1QNsVK0wW1S5NaZjK7JWAhjz1hQgrT5fmpPCGGyUSf
DUtirAMb6Xu4OBB2ZpBd4hqH4VsJdJQSzNPnlQ/t3EUZJ2KZ3qIGBYIq6pbaBlIC
mLLuaizZwzIf27vUhYL5JaTxS8JIVNzRDMnc9UIf+Q5zoWRChE5h9pJrQ/BDOktS
Rr+k5opq09nMGjffhj+rDOdcddJFDE7ZnL/jjmUP80a8J22UGMTh84I/7nCS+haS
hPJCE7/MikJ8UDw0gqZ8EUt3O9izx5Zxt6NluCJxamTDbWim6vWS5M1d+wjWYVRK
GhVlVaNbHUMSjWkbUeMkp80M7/M2aO5fUUI76wPg6YJ2RuXkO0UUgZ2eA2sjTZYp
x6BPjmcLarA4zMz1uzv4rqfeLzizKuQ2MTjr50bQnXI/BwFCWg89aIEJPCbqckLy
es8lXOIOayYfmy5MAE+8MD0Oizi+3/JT26KRgJSu9BbTZjBnfQmb5gjpmK9FSVsT
mtz0bY1R+G3NmJUCzEUzUNxy4HC7SlOYxmeog3gBNPu5Vy2CXZDXRBifo9yz6BoW
SEnTBhFCJNIn3F9PQMvWCsBoVrk+ME06F3ralWhEqLBlUTITarpVk9y0M2ilCU3P
p21n/LQ3I+s6ghnwT96Ots/lvnnrxaEg6KCzE1qZ8mNyoxOZh5Kpn0ir7eLy4uWe
H94OjVXSeK1vkgStPlg2uKbkrI6xJLCggOfMbGDx7v2dQ0QJ2R7xVoZ4RLt7It3O
3KAd2nF3cSVH/otZh4O34YilhU0yWF5+aiJv+ivWOTW8lC3Laur6egbL+bk+Ko8k
nMWXdRfVQPeRPu1a0KRP+VB4UYt8hmRedxcuv2z523V0oqZr4eiSa/JsYHGsjKpS
LQVqu0n1JYAtzRparql6n0wFk9LIcfGQ2c12O7VvpI5NW/HHXhOE3uKKPgGauCc9
/M9T8kMfR4KXITkeZSG0xMgY0nfnS1kMsSiSReodIt3zvClXeaa0vPNLYBxI/ZDP
lyAfGwbnjDylCSMg+8mO5UWF+Tyl0jPSE1aStSxYyeLOMDqbOCDtRf7pwTYIJFr/
QmU3Eze8FrKnBG/0B2itKE7qJVBKSizmj4mc1Kme26Ur/oyjCJe6DFZrHzIMV93P
d038K62aXR7y8n2x+L5TxLwWVl2l6VtOgnUWeUq+hbK/048ycUB++rJzSXd1+Ira
xGp87obt7sp8Ud05myuC3USljf+sSOOyNtvInN3vwmZEZDedAm3qdO2y8gfUwhgF
hiPWxqRkTSKqR6XwRrRN2hFFFROdM0f3ZNdBfhWjx8ZPaASAIHrBKwDJcPJVF5FB
bNrBJpN0+kmSvVXQmfcCnQmZa9zdMBVfJ/MU2eW0uOVLOPM7ZFkmaEY1VK5TpyaJ
yYx9ni9Uou2u4pxTH91uHRrB08PpFu/uquDaN7n1XeLe4p2ps3Z9We0BAkwH6b5L
1GUByMPQO2Oyn1gCl3lHLvybqzmiLUUCdT6aSVjxJ3zLIeCbVg0lQymStAD4FhfE
VGR2en7PVuYrL+NSqvxzja3+DC+yJSZxoxc0ClXWVB0hNnrQctMS51phzoWldV6Q
FuY95TvQN5rEArASKIYbjnr87LLOQDpZ96iQeBiouwku3mj1+o5AjZA2y/6hWGkH
FqJhWeQ0h+Z0kl/h3MXPhPTXICy2kH6EAU4ab3/AtRP+qcyEfZm5o310+cu4o9F5
rWC97NqwKJg6MtOT7EUUImvzT5QclNQQK2vo9iTwplpOdH26/tz3fGkM4jKsv8gV
X8fBKPp2BU1v0utsmD7XH8JfCn7BPO2nAGqvhf+MHlp51TKkJ8rprDsHVuVlaLCW
WNQ5GwfWzJjglsyNiZnBzdnyvkl9CBC6fUF7Re4WvGvF0sCtr/QFkbY79PDatEXt
6F8n2FLTwnKYc6s1ZlpVM+9nk3/uHahY7Z2R0OdhUhSCKowYSPup1RlNsiuJZo6I
doA4r8gC/I0vZG5stp7TMfEAHLNo7StULJn8F0q4nhZjjVeroVveKIugCIwnTNAm
xtI4WDPSLkYz9p2eb8n1/ogjsbuISu3G34jWtCLF2iowPkkQp9ECKkqfDnAf5wuc
Y4FdyGrVvTI3910cYoIDDpndYTz+Q7EOs78iO9BA9r0Ud7QpwvfXhWIeA/lz9HiJ
ewB6if0FPa9ClLQGM6UDtUjtfgdp7TNV6PaM4YSJH+x8PujSkxWiQevuSzCpZBgi
6/Urrf2lEDDdKZ4EYjJKlIkhUCbKD6eQEzBg6iZuN9mi/sJSu1v5e5nOaYesWf9Q
+4q+xEbdV7r6ebIxdcD11ya5BSior82qEX3TAtZy+/Vx2YiaIemzLq1YIU8hjEw/
PaS/XCX929UFmnHDUSB4Z6FtQFbbRNGsD1Inpao/e7Cs/tT1fYv08G/o7tv0MJ4D
FhLnbbsESWYFQwj3y3x8IWMCKyXR90YWmwr9Ao/6/Qjm+B1YZlD/b4LrEN1bfPfY
4Aw7t7pIJ9UNXAZDMZSk7HFdy2nGZh9dxpkKKuJLnp33SMv0P5JULvl6Cybqt5m8
dyxR+uOlQZfywy2ic74VhB14PRMMnXg/NzLWAOCywlMpUnElW4SmJLiss4XGmHTk
pAPyk9FWUX+kZ6Vm4cEoBScTsBY1OnLPtrs97gh4LwvKlJUmQNLO48uVPzoiz6Qs
39jyiKXBJtvToZ4C09Zk74T7vT4xKN9N30obGGyvG/qcNXLcCGZ3Td500t6H8xQn
Z2PLHM4pS9X/UWiozzqYR7PQnYVyyGR5qkpuQNY5LGQyYZlu9RCJ/xr/OerqxBis
dZzrX8BEmFIHnXh289ZH+/LSd3GZ5lqTJ4VTF+G63yyeUxV9ZWWGiJiXRu4tsZfO
5HQMlMN/zalBUfgiCZ/jJBG+aH0SKUnikR6FbC+JzaY4uMZwcf2to8wD6ivyBRU4
yCOzfmOKTVwgMoMkakuL0fMqGtx8yY3ps08l+A+EGLQ3mrsxwbd2gK75J9jBLY/x
SnmK90M+8zNjw7moZIKYaPoZnPLY/offkL7ltkkBYI8pE0Hux4YkYvwv2V2AmJmv
DV+aMGOsnqIItRxvOKSxLx6E3UAEP2iouH+GkFbkcILGIVNxXbHlCTxl8LGaYLWC
2QBReWo07/vJWoseXKl3YgrkSf8LMLCuc2qG4jpqujWIatXY5wV54/JMhhmEFuY4
ZsP1pr2lD13V9p/FqN5wJyMByle8ZMmwEb1/bqOGiaYXQDx6QaHbTMfOHapjE7SB
B2RJu0fA82kz17cBAtbBTESqpUaPI0N5ewUxf1JUtvX2wWX/w6z7Fi3YairNOakS
Ydn7ZcThvhGLhGH+h6ZoQlyr27aOYGcEyuOWs54udLoiUGp7BEYuA7KSxdp17uNO
zRvrEIEO11aiQLh2n0aUfYIZvdMyCiG0EK/mxs8j6bNI2ziDHgLBFyCP26W34YHT
nXm+dY8tV38vl4EoOqiObIMXkxQ68Ye/t5H8CD+QGk35zynOv14RoAdBIW4HjVOG
7optHJPA2Y/FEfy1Gz1k8SNOfLDq6/Ati9mypmvNXI8G9U1hH1Yf5lxN8CYcdEUA
btbprXicdFfwjOAohB30iXul/UXqeQZ9oLBlMoZZBLi+kCi7w9n50Bu9oTOOsNRF
g/z0jqokyVulSY8mWmkJkOdN7MLrsh4c8TVnfM2jEG2PjBmIfGmObbjwLeGYkhly
KRra3J0Up1mb7UApXob69rguoqV434tWP3Vkv7m9gTiCaYIEiGevt55cZb0vSk/c
YuhUuvd0iljga3U5IyupdDfwQ4B6mfJ/n/ofNyjz0JV/XgNFcOgwZCsesusCpJVx
qTZYGVZDdCLCSnz9G/nib9ziuOx3YBrBfX1hG8Bku2cTmvcUElZsJHbXPQ+ks0QI
YO9RpQJBl0KJY1i5JCZtRJ43aa201GNmAT/Ny1OrXFYHyQ3kShHAHFopQeMaGDCb
Rq5wb88Eg2orglYwSN+2dkCCNCsWEMETtLgREzfBKH1kkKHw9wv4TVat1cDm3h3q
zdW1bk6TIG62VY9WLJsqezLJXFrvO1vNeC5hpH37Jhr9k00hAIVvcskuAcwbF/77
YhqeVJ4EETt4hgWNPEKS9i1UaSv4k+f7G3sKrAa7REEoewjWcSRmysZnBNr5Gs5b
3WglI+caSS6i7MoXF4yU3KG9Ab1HcctizaJEHwqTjtK5Lh4Yld411SvTjm9S3334
2vmUPXTXvEL2E9VQoBbKe98AS4Ot+bokm+zepr/llDk5JojNsm2QZfinDDHpCKUU
iIB8vJe1adQSqul5vJmYuNaBDqUcwWiGyzRd56ywTP38VJUEHjFTuX6Xg1SY4iCd
OuuMRAMq6pX67X1yLEcVpsOjvRVveMUH2kp1Vc0U9ten6+MAARYFW4x1A84/3LsT
C04i4l1l7xlVnA0C/MTX6PDO1ZGU2V5mDzGTom8azr7Ff1GLpLuuOv5lN9MmbmrC
uIDHSIzJtj0L33Zqd8mvLP2o8Bl9p0A7x0PgP26jIdZNpNiFqCkysLEilK2ko/2q
/TWR7G2cRrk5ZFa+Zc+7+4hAW6aQAhgucFcZICWzaZ2YXVMEZcDJMmjoHJmABdE1
ItZOqoCdGgSSR61xcrS0Q1ECs5RfYtYhwWeFOn/nLcqMnbYxv3TRxmkd2x5abDgT
VPYJLTYWMGnRwE9Z7n0MVq/TSfHBIuOPxOS1N+uRIwG7IapbtKD+QodmsTIVKvep
viZi1ECEXKP0JRdRnkUpEdZe0DHw5Cc5fUQoUcg/L25bvlD+Zl7DYvFcfbdLxlVr
i1VFbrHao0tEvrMafOrci4gYgHOm4bMQ8fnPhnk1w9qZZxAggzfMXt7uDV3Dk6kM
LIJUI9wh+VC98MH4fndhPPKZEQdh1RO1RRk0FRDKOFqATfdgydOIagTPHiZ0b3hu
F8UVBQKwDfwbcmLVK5W7deOfx5Ew6bap/gUj8y/bRWzSK41U2sVFDE4YX1SyPqQi
1kwQF9roA21lGly+sfGJe0dGYIF3DHiIHcaqSVPUV1eFkk6qVrKOBHD1N4SsW4an
1Bs72MNKVr2jnNShL/UHNi8jRhRhT2aKO3z6Q8kaVb3lquaEiOfVHGou2mPXUSnx
/x65ACmbVnP7FCopX80SS6YySYM6T+L5cqQXgtAGtcJEaxbM/VHh2vwwCJe89Ez4
ypEvmZWoM2qxz+gyvIimIvIXaF3q/ObMhiPvTIoWd7DbctwM29vGpzVPKSKTrPqV
6tFmsAoe+0kXUqq30+ZOURFMnX7SfG2XP6LwE69Jb53PCpLnXu94V90jvOQg8UlW
9Du2d5ITCL+ZUHhaBZYnm59oZ9Le8AoCXggor5U1mRKrEGn4OPDVbmR6Rcb+Bi5a
4hw4IJmLL1FMph6k+/euB0HKBggFf4ZkUA4dFPPUme+roedEBlLQCLAk9txc6yh4
lm1uEtNEZ3TABujlONIADF7P7m9+n0JLPCM+Aot0Apqlw6y22YNVUOhNNVXevGyN
gSQedvR/EogI/7t0Q/O/V0NaWjPrIQYphOoMQ3NsSYw6Xw63MFFpZBaxPwaop0lJ
bdiEsCsscATgy84HJv7T0N8o0e+RLtI5VqTLskO9M87eiVbA04Iocfb1hP+H4O2a
RkcGAwny9XwEmwiVtS+X2JVhIAKg9/VFIFGaDT8XY55u3vYKgKfMkGD0ecCVjCQq
zsDKyVe5f1QFWhAAtTGFGzC6Jy3VYHuFHbSlqJD7XWHdJmhJvSwl1iwufuJ3P3VQ
hMPf3ro+4QwAGySc9ZnpPoWoPWRpYJz1mTLXfEpTaIQBWPondXVcZBPCcUEWaxua
xiytg3Ms1pAi2gkTtZs5VJoOYQcacJT6AEqWT5kJFDhE0mMl6/BGUaG7EvXeNP0N
sQQ1VcFhpGjdX6P3oVLSX4C9Pawmdc8cBlU/NsP49w2pbgC0wKRZrmKUpc90m3CR
i3W5D1oKoqzSWMwCQMiQGXmNiX8g76GyOd0uaiQ5aDZDOsg2gOT8l2EtQ6BGibF9
4u7d39WuGfnWi8fhdD3wyL44YIzVMXr2rq/iiUnT7ejdefCiuwX2cDtQUYGQCF+3
1d/lPn6cOZuN2DkOyb03swQIh8cfyoHNwFigBzqjGulgJu3k1hSIPNAtXV6uw26p
KU975Cp6GZCwO5GDRiwXmN1yoLVos5U8PY5KTS6BQ+U/b3WA8kD3luqAi+xMt3F5
vLsSDw3izleyJnojWC+V+utiwc/wBvwN9dr45FTfVeANI2p6Ycq2G7R5kGfR+UQh
NmiHMppWfnhrRRBawFGxbYMAutxxTCrKJjJk78CkR1VNhdWBQRsOyd00D+cuaozM
7EYm6zeBr4t2hrHIY99bKzGnkLnsXFAd3yeWCsO8uhGvL8kmQRvijBamCoIW/Vw5
oGbfYPoYIJc+xxCdvAo8VCPH7oQJmzOysqu4R36o/goyw7q/EODqMBeYBO9bk4pI
EJs0At7GHLOelNl5rtGJ+lOo3ihGw8sHFp8oid+P22hKflOePGBqnd/Zk0bUYCt4
rX8g677W27ah1m+dkfvN/R/EzmmF86umnOOaQgNx0o8jRyqW8Vo8QkOAiatJ/+0l
f5Z+i6NTH3tCfZDIKR03vki0hmeJfZDh61CYrmcr9r/o377rPHvPxv09NYI0yq1Q
1wI+EgsoOPGRvZR22xMBM7sxUKDgV3SlPMkKzL+iOX0BwGbpPp8CfthIqGRdUT0C
uXZlkTDM9NAKgGxHjJphgcR2etzzBScL88S2wOV9Z3bdJ921GUEmzVJdSCY22SEV
HRWkxGOJxJ8Q8Y/xmJVUKmo14Km90Tesp+tgWv8PqfRz9r3S9kMr0Of9b0bMlRVf
kFKklTS2nr/OX4ofqVv+M8YxDuwem/bM4mKR13wOoY0QgP1hDNlcqRTYXTS+Ppzi
5XPaJczYq8cx+5kGgg+vYDHmCT1/ju0//8XUgIMXP15WVcSt4jC9sV8qUdAl/4ld
1J6MhiUbLFY6GFixbdzDTV7MnZfrbg8xtwYVGUc9XSEZuGfIL0Jv/m3HPFNrH+KE
hwyVzVZ6j7ylBRsEAM4HyN1nmQhlq+Tmh8IehO4YKWVec8B+7cqiiz4Vxpn2x7LP
dkDHqpGVgowAi5MyVH6GiVzCTgRVD3A8qloeKFbEsI91h94KkdTjlWu8LiypnkgL
vlGtG2nUFSGZAdTIxFUu1swYmG+9DaqWPsTyabwuv5vwOUQzuMWQmxD4OPTwuLmO
Kbr6Lq414fc6UGWjxmTIVesSw4svmYRnF+JuKwl0gZZ1G7VhFHcYx2nu0uXzLCcV
NEpY2BrD5elis/QKxEM9JWGii+xhKUWi+BU9rhWj5+4MVFzvztM7ZKywfAPlDoY8
k/JExmQOY9wHDhYH0NQrZWBM3Rgx/q10vVx4hBqKbbdc2FAlLs1rV4HDVpGefr/7
4DwVzjld4qWl2Rumt8HXXL0vy+UxUJjVh63um3rnkx7Q3XudsvIKGelSyeyQJXyq
BhHV4BqG1RMaEIheTchFNP3yLj/P4KqWcUWknLXi58MT9zSNrm351tQpn51eKPDi
7O5Bcqau9yx5+nOHFP21vdjayMg79dWZ0T3oGWARvibleL4z/S6rSKNIV8PqyRR+
HXQr9mMn/Sgx6bTzxSCRgsp0yiR1pY+f0yTwU7Hfs1x17V0YwwzgQ7WXfJXvArkS
nWnraFkApvpO6MQy2DVAIyyzQJgX4G97GPvidztMEDHLDvLMXo+iFg0WzOEdGUKR
Q+Nxag5OXaxe5dxEilrkW+S6i13mLw6beDOTMryPaGVqPEFrUcGcAB8OHPQLs2QH
uUzWVtcP2nXIKnGlzgWK50ENzHiR0RfiP13VJr1rs2FAGCgUCBHkJHU/uDbJXfGM
m21Z79vYiQW+UgMDcohzKQK7IT/8Egre0CNeNjqTQWNhAfH8X9FpWz0hoa3UcPjy
zuSeAcpXn4Al2QRIijnJXYEYlrv7/D2H0nygV5t5OxQR19Qf7Grw+JiRacWEe0J0
G7Nj963wdJP6pk+21DBn62aQeOwzGZw0c1wlQSQHlP00Qqf7fSGDvtN1egd3h2q6
EpB/ZBuBkTvWjwxFeoXKoETNHZK9PxgwoHCQcCVWouz62gGxVKshCF4NimXzXBX9
2T4NO717e6sF1YtrJ9t190c4xiXsOf5pW9mFMkamwwPSwahB0qNiHg8up9RaDHqQ
OiFcbmlaIokreP6j+2xj6cENvFtmYwQHMjSNErDGtoYfQW4kVuJ9KG2irZYd+bEl
SxbJG7bpbrHTZeZ5dmr7AWrfuhNEHMAfWoHB2IM2LfiVKOu9rmoHfwj2nVEQ2Wfm
CqFPMi17U5IeWhrmch/2I+Ii8gEpwynyq1vgZuDla+fMCvgkcWMmKr7BnrPvU+bv
l2ufdUeqtlC6Ow9Odm9Dl/QH3EF/roUJ+I7DyzbIT3uDX/8uSGqala3ZfRuJVu7B
cYatGVMxlrbK2oE0gV927xN06yx4ATPiI+l75ZLH1krc3kRMN9wQqIGfN8bpQM1y
og7N7ZcVsrsp7B+oy1CWc1NOMwbu7lH5wxcc6pKL2GLIQj0U+35CJfFzhjCxCRmx
Lf8pRBs8kitYxRz4Qrj6rWyb7Ef3yzFHiuWJ+REzFRNI5eMyyHaP4pJLu5Z+dJyS
Fa5XYWGAEozQiqbNKY1xZdxGQuWB+NstGBLutPJOW7icy/rRJmkIed8sCd4dLWZI
onIt0hykyj+XP7n2rjlfx2gI6KpMoZMrR1yXIZnZMGdkwuGqyFT0mtMmy2bA5fdX
j8YQ27AzmBW4EeZnlQ6N4EWyefZRXWYEgbOXwhcehKJ3r5caQrwF3S04QdkBdMcC
iIYF9dxlAW4EInVaRMXbeLoHo2zNWtZtBC0YxiRt8a9bTsBG1pWvnrHl1UAq34lG
f6oBiFSvMm8INwPkJhyxfOkL9Itk9OpzkimNK/MW8t/6lSPh9LwtrHkQhFuzriFA
uzkJDhQaQtlZLG6wftrB+PBZL5d7RUMDbq1P9yi9724/0UFXdoHkldzy6i6yrDIH
PpAIW74RMIWNaEzN5z0HomZddCn5OV/hXO6zhZQIS3TTVMblwaDY8TnoXHtAJQqB
S3AZCOBQwvn7xrYG9skopQBUObN4q7a0Fo+zUFzOwwpSJ8vevQ6LzofdFmF7XYrb
ncCt1lpr/7Q7r6MJA2cQxyQKV4ZWmMQateNTDoHMF+W7zk0K4h6w2HrWRdwFGbhQ
M6qobiRMgzcNtj8vMVrvhOeJqp5Ydt1EbIz+2X+sQMYfYc2cTWuBhtWJ+mlVchgH
IgekoLa+ZxUld9sCqu+XSUBFDVjxyAmkxuiSf+McEZd9EJWHV0CVIC5YDk1UQOOb
F7xfJ3jDMgXm9rze7SaaypBA4fN9/k984CZ/mEl/VHdzVvWYhCkQu0gEqDGuVbzF
GnWgFO8WREswGOymO5S5wN9IM7Lx5lzIB5PSg+xMc2IA8fcWN861IzuaX7M8lme3
0Qp6CEkPHtG+4Lyvruz5JgIMBuRY5XWB48zMI+ACnE++lx1mzUCCx0mDuMRHlADl
eidVvSJ4dW0khoyuhILCh9FuX4HdWj+X9+z8u9xeN/QQQD/sLjMDz53A5pvQbfLk
P4IBLvYIZ2hBmyevcG5K3MauV5rkctzZfjEe0S+RhrTHm9pyFQgB5uMU6f1ylkCW
9lsHZ2L1nWly0uMScUP+FPZrHyvNaKU/+04nsBnWTFlFd3WN4V7uLhKOfYWY5p//
+h2LZstWiKssh0P0qtcQleEYM1aFQltlbcazvZjfshPMySn3bdU4nQSb5XaJcwJp
4LRGfwLlhPQ5ztf0RLEAcGOJMyXU+oXH6VtY/+vY6P8z3kpvqqTJ4ryNy1gD7HC6
XFxfQbaB1Z9213BN2EJgRSxS2+7ovYPg+q5JAGwz4k1rGhvSvUJUfu3rxODsn7kA
aqs0dy+0HaQAmqtMAv53gEg89fybWr3u/I9liSzMgw3xnvTh/uy2v4Y7HHM9nfN6
7pklZUP2qVGvlEJJhX9uVfeUTJ2Ax4mNAhetjVg4tCaESo5RgCJN6omM4B9ptBon
lx3lQoFx7Qx6qDtE17Qk3CdY1uzutomy/PgeDSJ6QtGebvKIc9QLsSZxRkVN893w
wYgqCd4jfDlFU2EWxNM1jIqcUjxD6XVBuz/yG+ZyOCvCmUy50dQbRlLp7Ss9WUG9
TQGlOWghwBFK1Lb8oGD8sr5zcou2B7PvT9XFypFsOOABVi1FybWKFeawlBLrRZgp
5DASy3SUsVtmBMdWViuPjYJMC9dT79ZGbo6U8dvT57gis6fkqSRk843S4HsCfP9P
noT9f5R0/goWa7V7jocnC2LXczUrwPvAef58LCmIqt1pHnlozkPb1UNU2QKIKV3E
du5EO6trTetrWOk62b/ifZBTcHgNyZ5hIAxbFhtVpHiO0dDdS7wY6NetUezER0Mp
HmTiW4Ja4Rsyxr7GWEPjZWWAAV3BYKskynoeKgGS9vaDLTb7FQd5PpC+L0mZFu7q
EvHzb/qrY+ovkPFtItbuUeQrjayw3b0xb2aFzz5wXGWcrwIRcQZV6iPZq+2zgPIq
NpzmAnNY3rH7gRjxctOCC77uNDFtndV5seA1wjRpvq9m8YLvsW61Lgt87K5jf0H/
B83wJZVbXmgPk401CulxuSX1aKiFXOk/Vg2MkpK/U8pp788Dl9IFguFEIv1OZ/EC
eX4299y3f+pTwGe8YsFgtU4NQCVEGgfvn0T3QR3wJ+UcFh4Nr3J68hyCjrVhwuXB
FP3Tb0S9IfxJPFyOYrL78ZuWNIXGAssvjDQRHLWNwA0zJBRLNrYn2k/o84Kx3O2M
fSX+r9D/lWbU6gdRBnY0N20tZjFnqsTbY0oeG4RREG7JMESVsHFpJ2WHY7//nTqL
QRqKbUSyA4ZPoyEgdFg/gtjiSljBxLORIEEHfvAT1ecsN4mRlhS4O6/w++J9x5xL
w3rZtfxdWlRmT8SaZXXCyb3Gu9cO3G3YrGCmJ503hgw6o6BObqPjAojSgmpnQhQI
/kzxmnU3rO7Pt80r57fPuCYU8beib4Ex2buXHmiDj///7voMjIC78A/uztNrDgq2
AZjFjfdxZdHlywmmJ14rNnVDothaDpK+HEgU/CrJ7KoGCk7FxbSexAgDme581m4k
Isf9kSXpKhO1C2opr5gniZGorIkWGeh2uC6vkppvHk1XxFkMsE0NTs+biTNUs56t
UI+0/+8McaJsD7TXQVKn12ONcTaSNYO7mABgSvrAaFF/jPasmaZjpNXwSGaI92ZH
HzI6VfjsNpeko4V4j9d1zsZ9d/AeosQFKzbPpIbFwjLpZwLXNADJ7C+O4Cwlf+ef
5aJpHGIbWWn12Ou0yZTLDHOsJdzCY5clKgx/5ZLX7sEXdWlfTv8VhiAX04PkfmDu
RbDCNE9UMYIyT1vRhLc5kudviS1CX8CUfzNfgv1DBAC2k0AQ45dEjtNSZ3Q/bRVh
N73yjDC0FXqqWavnSCde2/Ji0tYo77j8epfSBRccajIsjST5WGZrvOrJJDJIv6Gx
0LDJTj4idATA1S1oCCBgqT5rlbY6bvL1akOZGREgSUNa3I4bsshfkpqfhlLo0JRR
0iKmYCJ19Z+8+OtNd1ReqqfLwtAPxbCMZOSqLEmWrdhRExntd0rNVroHItRHzrzl
Tl9cL5ua7/tnllcAzwRMeoGU9TLRuf6s51lWLl6EUu1MaEpoTsVHjQeYHRtgn1vv
ewzdpuBVs66cvYIJFGvv68ZwhCP4lJ/to0ebjppo7yNWp/hyOJ2NOL9YUbfOLWPa
3krcg3mUQf+wuBoTw7G/ThlfJTeul/QHS5eUmmvezgmsnLq6LmCVnM1qebpzGSf0
g9CO24keknZbi+mk7YLhZ8hd7jKvCKbHWLjjlBhvYS3sc1/Zjd7ZEMvFWpS5ZpnB
SOWgIyjXUEXVN77jZ6i2rqrR3/Azqgcc69h0l0a8J3/4Ot8uA0S42WrPpiqpN+oo
l7yLb8eiL/f5fSDwJVDL1+dCYG8zt4S7KKl33U5WaxETTh9Cz8V/9uU5CEDHXqhG
dR64frwREnzoCCallSIYexW0pQTsS2PFplF+zZ9qbQF1k+YbVxt1yQ6+VHSu/+CX
mPJZUCT19EpVe9zWmuyvyBEPLqYp9IspckVO7jbeAeQTy1jp+aeQtjdsSAOFvSVM
hFd89i4i6dkwUR/qBuGQR02wBu5GyklR7wNjtnD9zbjBbkR/qioMflBOkdIReIpC
dmevRsQfGndy3JW+vzytiDYxbjnf1jffGjXIJJoS/MZetfTen3bYMK0Zy6Sy8+wd
6w9VDaQn+K0yGA8d16eKtrcH9fRtpttWUz9Yw6BE9HaUPHQjOEb/xLT56DJo1lpW
xa6/RFwFhw9t4jQCAW3hQOxkvk3EGfvxn80CC7gbAjQ4rVaR1Gm1S7mV4GjSz+DW
yQsFLXxKW9FG8Foq/kfPmFdqrCcdjCgfsLCFGM0T6LyjFRfuVa6ZbFRHpEhBmQ9X
p3/IUPooUw4d/kQYFkmBO0Zz2FtpQ20iKBCLQFZKTw9gudjj9kERXZKn8peEJkUd
ubrHoqzlCJ3UHFOimMYX2Gs5rVQfL/pR2/eI6SwNKl5XZi/Y3bfSrO6BgYbK8qbQ
hltyo27NsN+21X3tsNzSiKg/A39SLs9R5XBoxh4PtFSddXI7BiNhx2ddCUh/EOjq
hC6Uv7I3v2z7D9r0NXR0bDYvHa37oI0S9BFDw+sgfcfZ8aDHD+o0CTK5caeqlAi8
1Mo5LOvOrDXx8CbqGFE2qrhw22HiVgmOOvcTgSEqYdcr/SiJmNw+WGM0xXRpqwTd
49vvMWkfwbU/QmsIYZeBlCrTQ4kuWa9nVdxgHHK8XnInYSEN0uu5XG3ryCpqxzbp
l8OD2W5xHar1aV05p5NpLYpbS58qBqRHv2vUG1ci0erW+VKNauzLfZGA9GOLoiiw
LCQCz6VANMIZ6T+1hi8Ye9r249T3EEWqaS69GM6uRuV8TQ8QSVnRsKVh8vjDO57I
Y1d+QkzHr8ToT+S3ptRdgw6IcoSypAMbfsv40/zfScuyAmgRg8Uja6k8syVL0AR6
o0xumXdKw3lMfB6qv108UVTOc6AyyL5ypd5n0mbMD08p8g9HemG94evYyCMw35Bb
2kOEo/zthrGvSADPmVI41rsLUR5QG0okzSrronJatK3hPyrA1b9atNEONc+XFcMT
IeDYmN8rxxRF8SXt5kxWEjy69V1MpLE1TCpG3jb3Grrxnt0RU+Gz4BHEUuBwbC26
hqbO5D9ImDpYWFYRrior3Tb1hXYiJhX2gsv52EpG2L/BZJZN5ddMFbfO7KoxQRVG
PO+zGx/P9ZzlGiLA7EbnjcDV/MMlBmvX48YKbziG5XvHBw+1/gfuTLzWJV4Rfgmp
LTDrZmbZ5z3jiFFWeWhdsodFiupx1Q9W6Hrt+8CVsIm09Dia1AA/8pb8yP4vmH/I
7V2xEuh34rX8jaBz0ASDygLfdhBRe8cfIKZQGG+it2mMRStevyjaXXMlLqdpYs9t
5VBz2VFlBsxx18yckORQc53A9yIAm+qr6QizdWAbMtjJFgOGLJQcscestuGVizA5
z4h2XETTi3YIEk3iHq5aYe9niYniP6yrAnVoEPbaLroWhdPsxSVj6j4rVDoGkvi0
kbM6/IlVNHlyqJawLo5EKUEWfVyTeKd5JX2dovDNV+sR0YevI73kmMciOKoHBRiU
6ptY9hrsNAYSc9xK97ncHQkhO8e1WnShV80RyUCEvPKgyiXDV0Meartrqbu9yrRy
+znarJ9TVsF24hZQemAW2OFAMuf7Xc6VIGjQqlgXEFhxKYpSXiRchMBqfyt1nH04
hmoe6P7tk8EjYmLpPv1Ohqq5phv87win6tzFPSoPO7oT/HldPe8oFifVmxlGr5nQ
lYlVPwigq4jYxTi0jN+IMdQoQvW1v5UWMCl7CMKgAp4dfy0lyKuphWvHzrqeyJZS
yl012DqZhFNzlZuHhGCUHD4/XefATkBa4H0hly5xzKm8Sp4KYR1o36YE03VWOy/s
JGzIO7l32we44IlamlkH3BRM0SG5CDq9tWci1vYkxo7X6/L2cFNLzYS6JhHOn8+o
NzWGjsl5pJRb/7dc46ZapJO5UYaLgp/kLvQLWmMaY1PksbhMHHylnD4oMOdrzIIz
ldDK8MmiBpjAm6+eBY65jd1SCwUNvb2kIMNatFV+1UJ+pxgzIjnpFxtXrVpMJlHg
lmgN77fAFl0vE0t5pGF82AeMoIIiZd0ZWxL/xGdhZCVZ/86h7HKPbrZahTF4mD5B
u95r90bfooBE7Hhcp4xw0H0JMUSUv/CWuS3to2ViW8AV3MoSCdM7NF26f9d39lIj
lFd+y/vTJe5xP7KHteiKwunHHaVYs3bLsZsvCsU6gOcUFiq7Fyw2n3rLInB4yVNC
686fG1XbMZNvzNZoIyz3rEfG6dpiJtH009FrBQKdKCo+6Jcp8hwC5mI/3Vu+5EV+
dnvt7q3p6u9cnTp7AZqb7D63ttASTihuU4+FUfAaT+5yYZe/1PcguVV//Ia6Ph37
6a61KULrswHbaDgg7IvA3zLvCr2wQIMTOJvvFgrL/UMTHHHhoOEgqlxjivauoiI7
uAL78tQ45xmEzA+Q3K9sdxRF0lRl5v4DaT4sCLA9uEsmLVMVBVr5Zw//PR2T19lV
UAqw2EjlG9oYGeMQusrwY+eMPm3clpg3ej3yhGFfPzkJMSJEHtng4DVr8FIX6cnB
EFnduVBTkcmMEml0urN0j0XBn7S9oC+KU0OamwAcVKFp4B6Y2xCZ4+ppyWHVVve4
vHIrvLexjSvRSnfCC/gtNdpgjSVT5uOdqK/8dj3t9Hn1/BT703b3v0whNGfeUojk
Avcd75+k4Wi9kAVwtbbSo9th2XbpyWQ4FUf93otOvKBa5cn35q1DgEadopjc4+Kb
REQviBr9lgYHgMEgP9XVFnxJY3St5r8tAtgaz1cPXW7u5K9ZVT3hY+Rpy9otcR0n
rarPxBvTcWuy0FPwNuIfgzMUP23o30aBxUXui84kEYVy5rI7fSWMtG1J07l2nWmV
IYKgLzyisc87IUgJeObPTfPTGD63tF9uK/5lNpXXQFfkwA9Oc1O8uUN84KIGC8ot
bFoKcWurpYDymnaxRqgHzbgeVPcnoPBXLQhM0HlweNf3QPMEigr4onmcl3TGOrmk
OebvLtS0H6HYpYAmP0YUa04QVSnrqAIfpmYCSGOTwl5gbvYTjsja+QzjXS6FllZl
Qro4YeT2jUj8Ff+WYirSDTIPqQbh9gnsviu7CI+G0rFn65Xdk8o2C5f37DuguXDH
zsjSvDA0Dkl9njlzuYMFZWrCpZY4DpLAxq29CWAzU/fERVp1wHoEqJPdlKif2NKV
iwsWmwPr/Cn6bJltYYQMSmfag7OPlaah4u3cJhmNWv0ycPIDYPIJFLwbjrfJv8lX
PAs1qgwk2hfYK6zGym8jM9/VKPXVcVvHgrg447XI/wKIeNpsRUYU8GB+ObnMMXZB
CVUNCv/S3Xoj5UiwRCy26mi4F1pL/5emY4CrNIs23mDoHCV3U6c2BLrHvJiZ4QfF
RJI35lF+y1DShphdG9olcMQiAit6WJJ1Qt+zV5Cvy2pZNVG75STRApAhEY6lmV+4
7hIKlpKcvQwSnUoKjbIvh+fyHcRESX2zo1B71C8Xtbrx9HHFC3ShNMqRj9wDil9Q
HCgCcTRE9m/dVDqckZ70HzRk5VWFi2/AkymN/3RyZ8W1/PlPO57j74XgcVXWu7qm
uZNtCqRuHP6Zv5SK20rJVznN6juSBg2UP+LdLSX5SteZQCyLWkOGTxMwedm6AH4Q
3ww7CEm6lN0a82tdjdXDkjLafvJLRX25WGlwVZ9gmirAY8m/KM+sRZvM+lyQyKKJ
aAtJ1XFX4WRfwgFwku6DAFhCW8LoUNvAb1nwAnCQ5qWD19Dq+We+dEMDFNtyTefv
1yo4E7M4FrbQiydGBI2OwhJfPFUoAty5bSiQ3oBZlzZ84+xWBK7HNZoYChALz9fX
HIdDoMcoGUNOzfcnNsPNO/ciON04FQHPQptRT/kIG3Rz4iAf5xEI1M9PJ05MifVq
9D+Jw0L8JUMiYWyF0iwSTsjeYdoGQ4wmiaPUa63CKwennMrQU2xd4cElTXmB6b5d
G6qo9WrSnvH7zYr8Sg9SokDZKWyOIUYWGsyHFUDW4TShiLgXh9bNOT974ROs+qzN
zLpbBQWjqBqOfSTY6o0MeHcfZUC5pbjSIkWTNM0t6idKxUr8P2FeZhTiAoNbISEN
nIR+8B9MdgYFV0xgnxrUKa7hOXUclLIm85V5b8uG1dtKq/wH3K3aIgcnSD9yeuK+
st7SHhH/ebsz4UezKzoBr+NwSkdqB4/9ITKe+1HS30hbvuGFylGCoXLQlatetzfn
mZJg5Y8DwC4hLuYpDiEkyvWYM9/ciS0OdGLuqnIsaAxL179coTJJ80eWGwr7WoaQ
ZTyrMINljasBk1PfwLBvppmwfKozhdMm6dPrKSTJjxVHZ6C4xVK7YqR5TIqhbrkE
3EWSHa4lS5Wx4Yhc37MfpkqjsjVvL3A0Qg70znY/H+cxhUwu8JXyl13NynHy9ODv
hXOft12dXgBLBBQZctW40mqXCrz1/XQvAXXsl4F9mABa1IfZLrWG26DImPJSYlRK
4n/sFOUpxfuetPKeETqz+Flk9FbKTU5bfETvXbfwDDnhtoPPcVJMG/W7mVCUBiiZ
e69HI79oMKy6QMsXZkdI4u0JRZuG8yEpksXAOEd6Rxo7ezYbpoAST9FGD0xum8rF
mpJIeTNIgElG3azcJ/hRiz7jwY0UpsPh4A3ftd1EVzT03YkkN882xEcFSDzsAQPR
fKc22W9gUrPCnJZNvsD/HBuYVKfwo6sPb4p+5pFRNDa0m3d29gfYyXbWXbR2JYXD
szngLw1fqfbExbxr9pRFdTC8ZOOH8SQ+wzmuCjM8nNRzDtEOklMcYu2D9KeOI0+I
xAIyaCtFInWZTvnPRFdWCFY+YFxGzBaMtoTVadjVqKi8B6jaVJ50wtO7S43SR2Ha
UDfYaITTSEQ33nwswyghE8QnFzKb+0WFTMr9tdwuMRdwAJCVYEIc9F4ByfelhAaP
OgQjfIaAdpeYymNtqyEXTEMoPQaZ+lI1trx1nX9T/ytrF8jCop6ZBRTpPXchGpOl
tdibTH/R0xb/9midmDUW5c4j1YLSnjjTv+qBN2NGwSnT6mE/CP3HOfgJI4HuvyGd
1ZdaTlBaK3a8MIDD4PSs7taPhYnf1aLBpUs1CqTj1bhMTogtW1dEu+LKHsZlQHv6
kGvE8QJUW2XQ5H4VvMBK8VzLl6WliiaeE4v49T5THm4XqX+Xh4Zdu3/ZFgM5Exhu
VwsKMC6DhHz17tLUeSc7Ckk42F6mgIV3DTAQCdfwlOsXuFPptH2Ku/7r2wYfEZyD
BY9f0OcOkLqIeOfeO9XbEe5gGXgo6Cy0kvPpBMqmcdnHsqbrLZXiYLeIsSjDjEub
eBPlEnpEtuQjAmmfe0RkCPZ4nRfeOXEP7I9H/c1lflvXPfmQFnF3XMtICkRn2gGW
o1tBYCqA4Ir1n7184GhwT9lPPstQE6Ezm/MZQ4JXhGxj83Fdz7XTQ7JewVDAxDuO
+rnD1MH2XxNbK9HI1TE1LFx9Zt4YC3RGtV5HLOuHXPAnJM1JMkcXe4oCZ/E1aeeT
HwKP0odeNVXcDKbtlUhClia2urDcc1AdThpfi4szaJJDR92XWoLS82bjpT6WkcTp
S0wWUzpiifXfvNJvlkK2/taKADojl7uYBXRaCXjxD5kOSDtLQxHZ9m/uX36y01WD
O4jKBtCj1Yahxw+o2MqKoXcErrEqNFSIJBPn7LlHdu2vo9vy+6VxVTYKPGzZUT+c
919mWrq6qLs6e6DcQoIebMaU5L5Vag+VNvyzC4V4VDpz52Zj9lZjM0+arLLTXIli
lRex+GRNQj9XZFnz0Ffy3/bjDnLLLXLEqwXQmokyebGYJmb2KKqUVNBX7y8mP9HE
8IsdAPZqTU+kuGOi7xjfzZMbtVMNZMCqdADnU2LxrUtIjneVJNi/BLEAqnSNJbw9
cuEy2D9j6jXISLcrCK+uz9LjCI7MZGgTHq2ZOnB4MZcwYa1CD3JMUhH5DNpNFop+
vQFB7P7PEfeHe3j2JtN0G20addFEiuA7raTdLYvevl2Vgu4yEYmkGes5eSWnfA4/
2KwM5KLrPi8weR8XrGBup9VVAGWAhuZrTSAe7BQLRpymfA9/MUEtZ2oobDvsT6sq
bh/LEg13s4i/D943QPw1IEZlBZ8Lgd9eSXXCl7UGeP/jZhrJmh3brRuRQisaNOmE
NyUxVg6JVcLeFCzkoyvkz3wckeVuAHDhuWRzRBgFI3ufX9xxp6jgIzViHv16XY0N
qi2HhPu9+XZdeuQwP7s0KcHvkpOFDu+KUeF/oAxAPoI4RCl/yvPE/jKDEhxmkqRv
Ut7gUDT18VYfZR54KdPjXIexAda6wDbskVl1lqqDTy3vchTU/B/Xmuq9x5IopeuL
sfc6GBZ1L4vMVqNwPvXSxbbS2V3U4CbJHjMZi6CUQ1qqZ+wkALXs53zILgG4ACM/
hh8iITdQMWPiO7psrELPJrMkUnl8wSKxQV6TyCTHJHYPeiX+UjT5DyMto63DNPg2
rcKOuP2JvzBsYhlo5JbKV5iBFzXtvZtRrSarQUrexTwoqIhF/ACP6/EM2mWNc1E9
N6JfqCSZpeQmtiUv0lX9gBAZZD6TyiDCccOmQHDiRajbFgZNaWfw1+ekhVRnq6+c
FUF+m/kCBzp9jhoqgvFTJ8qYAKK2MWIZLuTTlIpUNMugrwHe9GOCMjI9pSAaOQlL
9QKKXRssclkW1HfAFwzup6qbrc89Oz16bJU2Bgj+Yb0SHrjguqp2KMPDqlo7yUUy
lqlf3G8h2wzGU2acDe2Mof9lvCx9tuCEuAn3iIjZ9ygBc9WssdN5XDRIPgvVR+St
pXgnJgzef+xGMyt4vmdjfkKtsizqc8esKBtdJxVnjFxaigYm00+x6b0WPOqQebJI
GBnFw6uHMvqIhglaSY+WAz/AOPJC8oSJLrvmdq7P9MhtpvkCoS2xWg/5mbOdx3Wi
0dk25wwzjrYTOOvlh4FQB97WrRoCA23Z1BeKXFQZJpDdnJeeaqWCoSwBD/bCPQLi
5QD+N6VCP3QQb2jSzXkCFlxH06NnGXQ3CGNYpkupeCUfx16UI4P0EW9A/zrGIKle
s2My0tnaGpJohbbae/o+vjceEA5iJOzUaDHJGX3fNoz/uYgDpsuWJ1yuXGYaY4Vg
kQWaN1FfGP3abkiP1Nx5gmOdjTPDWpZRP4UK7abd+IZjcqPBPJsmKroIjnpDmPQQ
tL7OMHB+9KviXmdV0jsJArl8HdaTtkrG+3kueVUwghujDP/aaUNmX47TWUWPKxey
Hv4NNNo2DTmb2PcWRjU3+Aq3a/ovzo7rZTeHP0tMxV9/eb6QcqOZba7CDDXUSwI9
wuhWx5iX3f9dmMn3r+QVVek2Z7rd6c0YbR9dCdF021LOYFMR1dYqHXexAvjWZlXA
+9VDpixJD1j27RmzJEtkGX2zjbeW58UDzSd2pV89+B2mtTKsfQIChdw3n8b0kxj8
ny6x7saosZD61uq/BHtEo2hKuMfJuz3yGA28IDr8DRAxStwl45TGCz9s/mzKB057
Dz/yCSnoklUWcMIxmYuKZncJhlzijpT18MIwFN2A8RQTfJ6+AbGhxxXUnZCVcFht
sUyrV0qXX4mLXd8PUhbJ6AhxYImBsA93iosRI1o4QQ5bJOlrWPWPmXwH0ngeD/if
ix+v49LB2t0llTw19nx2an4/leJH/9PJxUz5OS4R1QmocYFbLJ+zMaP6xd5NszBH
sY8hpQMr5MH1iWzql0DDGaENiDxMnWL35D24Mdxc1i478MOzg9f2IAYrlu5oT8Th
FJmGcQ5LqSs/zc/ixKbv/0WwfMpB6p3+CCZj5EwwdOn47yRiTQktlbku7UpP4dOo
dUif+k/IBCGfTjHc93zHMNzLyUN3Ui9hkgssHDlKPXtDF/sIaiYgzv/y61mvhh+v
PPvyWvTWppiKAE2G10aZXut1Mxbl66JpD5+HPxhOmIkbFoy8/wdamqzYy9v2J+Eo
BtWwNroIgqI9dyk7zj8VRUbNQ342kv7Krs6D474oCdYkeoQkmQeFGCW/bXnfnS0x
+sOMbWIYDz7Rcx3aIVy7NNvUCBJv6WoSYDrvQalF6UavXJi7Vk7nnZNQHiR0asby
pV/ULxNXJ0wmq10ZDbOdzsAV/O1mOQ5Fnd52ELdsktLC7Yo2ham4WqIYyNjiBex9
aLF6bYuWXOkqpMIELwj61mAFLD4RQ/PJwAaEGlgtinZvOaACma8NKTEsnS8iIZ0m
GvD2QYKtCg1wFzGKiPiOoRAUBwG+gJD9uAhefEafGC7TsuJ5yNuO/frQv7a9OOux
rvIlYKBMtjuO139MW2VwiVIN7cp2/e5nUpakMxM1piFhynBYFbD8qMPEPalXC9SQ
372R1iLiCT7zWmYaNNHG8NAaG13mLFOIQ5VAmNVld1X3TdkUBkAjK6IYi8oW6boF
G6+KTidnrtZ9Nb0b3rhXsKfRFFZcWaBfFKQALZjRe/YSREWmSVgtxZXf1zcXBh0A
69HplSfEwi+ZrM529UZtc9MK6YVELdSbAH6HPbmpEu2hRETEOr9+f0GiBxrbvVC1
draYOZ2raB2dQzyZ1LTjpenRpI9Yb/F7YVC14U60QgVYOTHp7/VpIL8uqAwd2UF8
AKF1EM2pO4Cth3wFC5HjdgA12pt4qcmhaXluRx84zCzsrLRIlrpshKzWp4YC559p
aoXXCLt6X3OjlSBwDpvGNb+LFxUj6zmeSy9w3Ro2bhUKnyP+eEOHfPb7Bvj2FvxH
c7zfqYzZvkLA9mmyr+EnduHKf0CuUaD2s5pSWJQGzHIyCtvBHsTh7kzk2oajGGNY
RkJ4bNFvIjWdlovZQLLl03A4GP5Lg1La9NdvsT+OUOzH8OsUs7DutV2Cu2lVDYbq
Zyrq+ciiFXVeND/RJBi6EIfzyqg9hXCTmVWZrgd+pIor+1agdrDWiusASabj83yL
7VklTu1GbvQn2GIKfabZOhHKYB3bx7xMaijbMOoCrH42uYHKOFX7hA1uKP41hnpr
Xr3waadYRmbqRcYCgYILPqWTIL84N8N7QCOzMMKsuq8kHWB5QN+2+ja4Rd9gO1MR
HFnJIW5DPrbmZ1jKuzlXI2EvsYTBgaf6eIsMXhJ96R3/Jjb0fbHvJfmce1iTboZH
iYDikfpLaSNssLEoOAaxpi/EsRUw98BYpsJodXo3Z/k3VNwGMvKwaDbdvHQQuOAL
T0kvbtA8PexKetsnze+3jA4OLuta10gmZMDhO+hvHfVuWsffDcDJyIWjtD4RITEA
xS1hpAHO/arDLQsB32gk3b4pz4qqEl5M++SA/hL7L/w9zdh6QX3B0y4tsRHww5CY
lOHWAUHoni3aqKQij3Fo6Izn4jy06HsIC9O+fI8gLk9LS8bSpmjcbK0ThNKfO/jO
lKbzwQPBBRPelf+ZRdh58VSqYrECepdHzYMqtvYUgCmUxZhp+XHs0gunj6V7iS3B
hqsZ72BumxEY162Hz/BFItA/QyvFUa580LIUkK83I4F4XqT/7Qo40mlIOaERuEOf
BIJTMu1l2lmZ3xWN5NsRq1F8ugWPHtRs6mIGfdJRPugzKDm92jeecDUsoclGptbE
rsKfcKswQfHZoq66QIvYFoQj7VyRVymvxRdMLPPJa9ilYTOfBVvRg6f8aqgBhkct
2fNTQiRwfeZSBGMEG+KJ+h4Plg2QMhhNpJacpUkw9kfRfAav+vgFM3m0jq5dNpIj
dBBT/IxOjtJ47ajWrII00ZSnkgGfqDPibLaJwA4/7NUa4O3ipo+/OJ8amvfSlUuv
jHmhY0W9lTd3IGdM7Z+AJ95so8lz1ZVYyuUc17JxW0PSxdJfrCHRzr6Is0fyFclZ
9SFUxEEh9gLlVwaN+VVCzVxdsCYZkKF2jI4BNj5dX0k29WQis5Ja/XFF1z4RjI6r
HNhj0sDfbESq2opfZvOhQiTEndMK0zYWInobj2sh05QzAnI8EXhyTo1AZ17o2/rs
wLAz5wvg/IA2N6CrwQBNGDn0JPXP6HgAuLWTphpsKSghRq6ZJqEYeoUkQo0dAQwK
wNtAEXw125aMK0Ruic8kpuIYJvKeNWpR37YJw1VZoZcoQqB0ItxVs7R5WWEc7NIg
aabQ8dJoCfa/fE1mBVbS88ktzt7/Xfmo1Knv10lpsw+djwINTzvAt+LnOaY674tQ
INt1/Ca74w6NBEjcJBvEnL3pxrfJaZm/g5SLUk5LrKwXUGpX9qeK5N85/eWekzi3
kpMLMQenD2CIa1H3N2FSeFhy1tJYzNYP3DgFiGm7b1CJQL5H5dhkArO+oC3gvyBY
5v9fOP8VxaUCMMEqzJcIee6yIOf+rkrLQelwOo8kHE113TZ8BVZav+vEfHuGmI0w
39grkHv5jC8qX8HY69JRFGDP4nIYaLxdy5Cm0m7wuVu+Z3CT6umBFCaM/W2uMLIa
/+kIVoVQXnaFB+8xpKiZorUTPW6HluswACRMHpjzpjt6qJyc0njm9BPenw6Lu7ab
tO2fJveKhiYT14PwQRaje02N3uoPUcW2ucMwNXDb4Gr9JwoJS5pH5Fazt1nXiA8Q
Kve9dd6WWy462qoKh6dcxDKRUYe0c0/mGs0EyXwTR14WfoD4v1m2hKiMEHxDXwgC
DLx5FoZE4ghiACIC3/sF0JAHHtOv2cX9/9AdLhK+HhzvdiCaf8aZNhsoNuFgaQE0
MJ8WACHRmeky8fP+W2wVh+tb9PXDOinIL02sV1CUAe1y1OA0M+79mV9vcAbc21lh
WogBgYDGAd9wK4uHqueD2lI+E3vU4QCub6zED85w5cL13vUZvE8sux7t6jPeSSW8
mt8mh3VNf83FjG2oZ8Eo+IjMwNBH8tHRQCCeHHmYCCPwo6I8H0QTFcLskGRBwNMc
NmA2btU+A3PELXOP67iCK0tNrAKeukylatRGH7XTaj4rGh9VLs0LgQB0fNIS8PmP
6FBxI5hiXne+VeBziVZMhkp1ueszVG111y90JHLQoMlouwKg1KFlUmkbaaygxFW5
+wr6aqiqJI4uzSTj0hB/CkYZqBpY8gGpkado+QD23UExOazjXDSI5lD59mAndqdR
8d2G6FLFBHq5+Nnx5z+iIZgL+MciL5ztRpK4MIfgSh57GN45l2r/CRmVL2mgH+RS
eOmJhA9qesAHOlXJxvERDEVkrKgTG56cY+Rjflnwzm39YM5DVq4gPe+ktBEvl4aF
TJ9sJ5QhUuzV3UrhCZ8GMHMkIPP0ifoii4OLSmwFeTVlV0ioSMc6LRq7/PUgpc1S
S6qpS1mLT86PrKjNgbN2aFggNsLu43bddfZMcBLKg37YfXToWiLsKziZxgsxkr9M
u5tOWpvbRqlUv6yujk0/tZWWAHcdn63Lcu3VZwWkNp2/ceMGGEkpydfegcyipspR
HFtpWkwbc+N1/Ix3wBKa0BKE6LTTxE993Uzvt3/8neOBHTiU/57dGjubWabADfAz
oKdUM3YicMUuJtZY+teiQhQ1v0qWVEu9q1WATzhotmwFMYJ8EGjpjBhH5YkjRbcy
UP76oIZl+O6Lk+w63Z52R8s/Tec6ycR70Hkhd7hjS7rioOpcsOor0GegI948++20
2a2SrsPInXcWB8gjZk7ehpUMdkCUi69QwZUEl4wB40+8JheJXJ1lldu7Kt2nbbsT
IUpqOo76Iv2Y0L9BaM/VQAS8gFQsV9yO5JYCyP1wNbguYW6Fq2HoY964Q3FlI6ad
IthvvUN0OpeKcmDaEzsC7alwYxZLijo4GR6Jw7holK4ad6ot3Cgne55FMIIiGy6F
6CZQHunddAHcTO7Z9k1TPdbHNCTTX3Fpv9EOgZ+62bBeDdhCXgqbm34s4lqtGTkq
+gC4mkKAxLrAwHMFcHr2G64dZhPa8Ix9+YLi7Jv4gfMvkOH2yy7a6+v7bFIOB18y
1kcDq8Fw1ez7ysgx/ZWP6mEqQgFxit7Lut5DmX62fnXRirzUaVfhPNPwVC2wFmKe
65G0phcBlWnTIm28IHF5GLA4U1rzHnXeg9qSn/UfuvNWIaRU+w8M56O9+/GoKI4m
PTVtSE8fnVD3GmE4QB0smvB/eakZiQWR+ftHuL3FLBSLsRm43s6JJsjziPMdcSCU
zqNTLGgLeLbKUsX+epa78dgZG95nUzHyVyMXVXd6RdPzutjTOQUV4naxQ9w7U4+6
P8hSHjEqRYoH3bkpOQtSh9wqO4nkE5Y/5Ng0+MF2sSvexLRPI8td7DlefXSzL6dB
AqPgHiY9isBX2YfTEVhFnpBHk3KTsr0p8rE+7zFKF95O6XS6pTzcdObPyPR6vLWH
RxsOoL87tMDtXxDLgFb611AhV6M12RP5Pbydqv6QsgRCDhbr9Yfv0nu3nqc+1nO7
TIzN20uJqdTvlc0yCjGHODlw269jRxxcAd+ovceIgpzbveBOudeACkdWWzg/DTiS
OuDd4+yelTA/PvbpJAkCsA83S3d/cw8PfHJ7qIljACSe8UbXo5XmrydwTQp5tKCC
ERGEyimdc6LWQn6/VYE311UUrMEVxW+DxBlA1Wm51/lcXXQjnhmK0lkRowCmnPHd
pTz4lGKmhRJ9DeoLTvbKMxCUK3sTn5TjqgUfWkf6C112fx2cU1hj7TIHwYT/day/
BSHsag752BQwyGl2hXRl7OOUCrVih4jTqq/PhOtXCDtrjGuDegd6r3I7gQGkXzrb
3Ps/Z6EEtv1+UsKhBXKKrRL7tBa6+C12tOs+QQJ/2Srvuaia19PuXnu7KP7G+QkU
ql6tfwWXjmpBAzvGAreM8Ggj+vuwJkATVu29s5eOXA3V2zhNXgUtLNsYbh0mv3Rd
UX9VJ8nMBWxS1LsLdXQmir97UDD+Q7bjxsbItFDakt23YTcqxh3I41UqqS42ooiM
HSf3GNWSiaBnOjJs1OJkT5URphungsiHXk0whIEtB2nggFg8PlA6CqzSv9eU65hr
PhuoMuG54RYvO5sbuNTa4QA/awl0SyOA15PPJZOVv+TEXKFb7WERRWVoBr7s4ezf
p2OBySnVeI0jMSz7dbNjtwn38dz+09r4FYZLZaJ0yrr/1J8j6Gty/7mOpZtToaiS
PBN7Td6dTUVrLljN5qZQAQkZpm2wfZxfO77Q9tsyLUCfLqK5z3MFi3M/IWa66xDm
kauMKD57q+W1FZ/PogQypXgLP3tEGjE5yRQ/TfimMlEpiUTFwY8rZy+96AifH3dr
T5W/Ty0UFrPXVEjju43Dkq7tZxkvMZ/5jvLGE86aA8jKawXZlHjJyfbzaQqcTBjI
w4KsAgd/1XkbK8YdpYuE3BaegVSMVj5fHNFrY8uM3iy4cKzYj6dcNdo+4cbzFqeO
glLmGKPVE+6VCZKwxliGQ3fcaU0hu1/iJoawg5LE1eq13IGi9CT3qQwPAhvDao+R
MFiu21qda1805CwL42EclE5RUgwm/Ue2GtnG+UrZfAoUlBBZtj+T9bT6R1Kojnw4
HrHgreELGP+zcbVFirlPMe3AuMM1hvs9BjLJC4Cxu9/wu/+PxFY5X6YKahgMe1F0
BHq/OQjLK/gsGz/2dCUqgbIn5/VsIEDDTLJ1jZjfBk3UXBxLh9NtObxvgqkcpuRD
bpDbuePSAf7LEUSqrsSnVkVO6/j2Iq/p0G7mjE5DrQu8CbYCQLtpyhd5qcrLICLe
b5cueNVQKcb6GE7MQkymOlP9LBjQc3ZkkdZ6zS+dEy1A5Iu8Y7af7rWfUXOtjQkC
ArH8mGztKfbsANfexq51wV7VahFNYeNFjswvbxYdfDh5GzO/Z6EaGZZ9HDPsZK54
2XHz+MoxRn2wSdhgz4F3HP/ltxIK3ggeSYXruHfzy4Ul6MIZhTg+Tj+zNv21TXcv
jIciGhTFyPsWOEMZwgyn1AS+dV8yzYcWnYuXLmWzNI5/tPGKZl5o2tZDaosXfCnb
dzIPmtvcDjYNru1MQkJthrtXdbWu8nQ25LvxeS+sgbFwdMsVUJ7P9jrWlp24nTh5
sUD+fPAR99tBB+a89KIcpp50jxsWUPK+6rhW2SfsUBcRS5C0wQRvaiBt5XyLapUa
4AfTCobtv8K9hdXhQFER1oFfKZmol7eU+Yd06weNHXT3ULrLFlPoIHk/aicqIDCu
wHEMxcxdWP1OupJP8ckY1hARpJLc1cprAGpBO1eSsJ+2gkIN2WVyp4+sLtcxAyDB
cZyNgFhIPRSwGfQ2RVsxmhO46tRk5ndCM8za2rdtqiVh6tbYCG0Or4Nvf97ip1SK
XHp5RtjJl7wv5+bJoTxnOmJbGO6qIdyZKzCHjE1g7LfU3Bt5N/rDsxB+1SC8YfDs
A7yuQD3oyIUVSh8a8wJHRsZ6BSjd/ez+yBC9eftPLWH8nu8XWRk6kZTMSS5hSmkT
piaxzOA9qE7RBAe3j0djs2/3UlzLJKCJMx68QL+yuPvAhcedH92cr+fT2sELT6tT
O3l/qoNNO6Q14ZoUvBjDTVcyDdfdhXB5ysoUhYXuYHe0NzZSrYzHH47G2LhpF2Ty
t5HxJJQ7MADuklWY/xaKVwttCSI4um1Pg997asb7Bbxrg61Y28A7jKRsOMVhxmrb
bDei64BOK5WECWAg33W2R/9y1Ag7VAhuEYf5bj6A4VW8rDzkAS0AcUa6BeF+MNsc
RG/smJKx502pa0i+LN/n2LGAzUbGThZKWrI6l9+7lIDT80ZvTyBq7vYSjzWi7uWN
6YBCQ+mwiFeSiFrxLT8+LfoL5PiuqJujFQvuEen1QO91RzRHjW2Nvan7d9l3iXuL
GXOB1nKq0MJwvoLKam0NILoMVVdkDDzO4339lJngsNeVgYnjZCYbZISvySfXO+5f
RWMzYl92e9HZc6fA4rJ81V92URLEmg2cS3mOJZ6NE+6q7a6UULVBStsFoIAplw6a
ooQnmSoOCu9FMTOKTzuHknpi6fOr65kal7TIBlaXgkJDp1Rnbfe+LX94T5C2flqw
RXL4HXVN66UO8yLV7q0R/44FYveZ5Hb7K6UQSKg8JqU6xY5AG5SfPkYInhwMKnDR
+8WYC2mSAAxHYV6mJhzV7ipPVK6gHGj7apaoRpl7z6bVUFugZm0MhHtDOKGH17kb
KQ/J9sTNQWkwaob8bOqxdodsoxaSMfd6reJbyr0JsSjpX0z816eeb3Do6gUjtfMw
amHitEXSE/uJ7xZCwnwyuQh7hSQSEEgByLPx55z7gYUCMTp+IscJxEw++xJryLWB
KKbuTHzzqadfZuLMojwH/WKqXqg6dIlhWZDm8PYHb99VM74yUAREbHNbOfK7IYwk
CxDE3IxcrBIxVYYSt9EfFoj7SBR1qrFgruSZHN5qjKLpgdHOml7LgKGZuclslntE
U3lu/eKOlUHU/eO4EuiMldQD8MRVToiCdkeeYzitG+YXJt9VXcKs2zZf2zvYX+r6
AEjFtELp5pnQDd68On5XNoa+DzwFBiccnroxagMUreB3pdRVfmjjU2FBhQN1RbFW
daUoO5a7PXbTVUN7jNV6+oXUMyvMKHr1sjWs5cFDGRFLMpjIFBHYUvveG9qRmgNr
ZOYGlF9WPldWgrPlf5YVFVRkFD1675/rDEcIR9eZHLVkKcpBeT+a7Bu67qNVgw2C
MtIYU+Z7lmqpE9VKlQ1ngbnArzNolqQem7hg5Awcc/iHxyt93uuWDcQ+bjF+S+mu
woMmQdcjfTO8tpX1Fc2AOAvEOHBKM2smNg5sALku6TswHTS3KofVB0qH7vqH7EgV
TiRS5w81SPra2YQ9ccPgPLWV5wBdPU3DgKDvg3ypRFveyuD4CZbbCB0b1TVF1pU+
dr4oSRBifDTv8Fl3wvIvEeowNYnr55fis05uBU4CPjbj4t/fYvsYZIPhQn4+SJzj
LxlprwyGViGEP41dGRBRdARnTrbu9m2JZwHuXYIs16bk1nShfq3OL7z56mQMco4g
0HZxISVGtkY8qgta0S4FAeyEWYXz0gVkHJue1Av5HV7wbuRCOY8hvtY2VHasTkp5
7laMg9SqIedQa+5AwwrOFOOo2K/YpWME2zAE4YT3XddU9sy2/GyIooACXwmzWy01
kZtgGi6s+rxZrahvSBDl9M0vA5zjpmlq7B97l198wiBv4je48rwXtSXRfrZHaoM8
RFif0q4EXuEzf7gOIwI4eVs67OpZJQOH1d3RsB6FiiINR34OGc5Jc/2NVonAO6gZ
1w+E23YNXMVnJqnF/dJsN++pT5kLlY537k4/b/3hfSUXF7yJKyofhlXaEnffpK9R
Ln+yXF1b7MUvwBUA+oLKksgSzKBsSsNK1Z5TeRVFEvWyP4SXzK3Exm4aDvNvo1uc
XXISWRjpAZFSKGcc49N0F4nSxrCxLqluCYwwvLUQKqQUlWS/T3pGrz2BLjfjALSe
i0kr2aI3sngL+iPIDA+KdhJPNfm3g27LmpJNFZUfwA1GqP0JXoK+RfHGIOX5QKLO
ZsjTlynoPk+KiINg5J7NFpcv9nkA9T8ZqiyxeeVG56qiwcNSKsWjvIr4gPmpRq27
iUx7ytGiUqvKumMDiJQMxufUDnvlVGB6Erx0IhZiZ6inHaZUz8/eWEcN04LTopiO
5GC4g2lRzTL8qRhBhUMiVvc4YmNvNR5IuFxZ1zF5FDXc9XamtH+SrVEf+HcxmIpt
ZrnLUGJK4j6YYsd4/KO2zw1JiRzlDp3kookrRk7CkDbDxCUbRidJwMqOmmMsEGmd
CyHJsp2iCzSsMDDv5CWpmA4fRV5Rdjhiq76iFfaXzf0NwGSpsJvJpGgs9hkwh5vB
HICsZX2CU69/2IY8guzbmj/mwISjkpnEf78ze3eolm4zzaNYliqYRJr0K/AaH4Ue
LbsB/YF4zsvnTR3ZpaxbbYHS+peY8yGatnibB1EM8t9suiHcuMZKhs5MtTt66vQQ
LvLxq4qGvcAS4aiAj5bRE/vR6XRcVMwNqIu7uBn8CmW8AxndHr9CxiB/KZrn/1Xw
vKzOzcO816T8IkEWzKIFGPnl3cBlfUOmzFOOTps0dGPyTUtM9xONhmPnY0zfi1b0
RnFXtni5BNQXIaiKbvVtmCM1jpHfvbWob+O/NEHs0utGSpPzL/IWgih50h/JmO81
8cDA7WXYlrl70B6UsJ5OUxMSmRfaWnrHGcPpHvSep/FT0G/MGJFZMfR3jNj5wIIw
NIUjY/1EhggbYbRXFJLg1AHoCFIMnOr1ZaKzWTh3JFL+m6pVmaWQA9WZZRcxWN91
+VN/F2U049bliT/N4r1r58D/F4FqCpYtlFPhl0L3UPcZfRQTPvz/IIG/iOXBOvtw
siriUCa/nePX2qg5Rkpv34uoWEaKlhz36sa38IXmSySsN3DA1U6r9ev/cKDOng5Z
Rrei1jOybkkKKYIzAEf4O0bJHfoJ6IZNDmxT1DA6PMvUkIXqzxHZCo+RcxLL50Yh
QrVMEXEA9YzoOxQphnRIoxQ+sWuC9GRJw3Q3dxx2ypyWdLTXAA4UHm5zgAb5ZmEL
1dw5NIqy8he4s829b+sF53357yMPAlg/J7Vx8O8UHAcC9PNDyToVlkHAZ+ziREkk
AHeuIMjo8+L7W5yhnxZEEYpssYAo+rYbXgDx7Z5OD+VAbCSD/YQt/hCs4eeEPkg1
paxXsyzPnr1gAYlPMordm/jAdbauPen1wKH5XaAei52yDDzluCjbJzprT8PAdC62
+IRtCimXYzoEgmVhk7GAX5QagxFsk2Xffe5GUpmRZI4uf0r/GtRz9pTy8Pl6Mfwe
MPUGVmXeV0lNnjES6ltQXJTZ3r9nr1zu+1vhFIiEEYGx10kWF4RRG5S3/9XXuc4F
44gMqGWYZQCGcmzPNKLN9+L7f33qeAcR1vlMqcXf7etTtdUskwC9FEsfvtSCrt4s
dUHIg6iwoZNN9hV4XXno0iR8Z9UBDJtX0ot9yupNQsj/DjZaG2usLvWQbg82IeEr
l3hfZzgZp9YFrJs2qMRM7nOCBIBa7cTqsxNKu+pSZ6pOGXQmSKkN0GRUx4x4UkXg
hdLWTsI12BKjFoq2UYIK5QJJAqp+nuxKDUQj7A9z2nIUNzBwFxciHNsGe8Tl+z9C
hAuwoViTIHhHiYBIzr8DLTFoBqsB6DQJ2+oo0ZtUDxvALpJZ2Ysq9yzS/4vJS0Oq
gxghT0lnohWG1OApFl5RHefqx7kftR3FcUPZGINSs884DY9EuMVbE3KTxx7BgqXV
0y7o7BHTouqOGwi1ID7LuH79m/BGnCkkcm0Y25sAi8zGTCMer0bux2M4jijZp0yM
7U6tFIBVXAdj6LhAl+Frl0IIDJ9oPX3GsG9nv59j7Z0uCueQJBXREtQJSposjQQy
7XjmPFHWyXxVLvHyxzidLoOS8siRen/T2ujlMaU0rvj+4K85mkxwNFGsa6zEXO0b
fmMfibITkCwyf1EYgrhf23OcP3ZlaBNJh5zbCxCcfWeg0r9aLArkwgI9XvSAVFTE
9fE1fxJV0Fpvux5aoAyZXd+qFHpk3qwO5+42IhBtCAjJVdNv//idKgvKtm38IHmG
9BNWsrdU4qDg7qesYnkz229FoI0pG3dlUqxRqJxQte6J70H6fpRxMoOrcQUxBsnX
RetHjCF2EtWlgPiy1LXKyN3TwJxgpYoX89iaJmVC8byZbFcdWrdEqg4PpY67lBTw
vrD8l5lBHJbaxZKagXow2c+O3jA0W7eu8U3zeXJUMFyYqJITXCy21zb4yipSdMx5
SUM3XDT+H55nZl52Fdr7P8JGaC3rva7dlUU861D3Mi8SDRmPr7Aw+pp0s5CgeSzO
W4pqkHp7EkmQxHLFmo7SVnG53B7eb1n5IsrC5s/KE7MhT6MUg7ScxJBaAPzq31VO
sncaV+7F51FFDvQffHTpwMMLddWU61D82SsHeRvr/ywC9ah2+8HZdw730lmivKwu
j2Qxa9bqMV6UJV/uM6fuwvuUQWcmOhIx2AIEpo7W/Byx9adDieZ+iPl/VGQr4nNd
mjPUAw7OjSG9G9OyPLsqj0eYNnFZ5wKFInN0UOOWiVC5Se9lG8pVQwp07d6VyFI1
8/Vt64k9IiZKRE11AuMbNFcJooUgz9j9XXPyQ8RGes03d3IuzEMbDpDXOPFYLMdS
5nLSU/h/CIpo17pWLKr9T3uPOoX1EEzYCWP9XNkXZ42HdOe18Lh1hOcc2MqdynsA
NdCWmPNep6WCrgs9wGWklnB9pbBfBTohsH9mAvZdDc9USRYp5MElhRLSXruAeOU5
0ZOLF+0o4xB1XAxSHlopK8ijd2cf+1F6ZXTZ4IPRetXDqMIP1Z/Et4ZEJYvwn/Gx
ccKKbfFdtK9PWQiqlG/LqEv/RUKwsHPNH3vWdJpxo4BMpeW4VQO8wzo8XblOf41d
cuaufPhfBretIfYwFNTEowIfpyFRMhbXo3nj3chpTNmHe5oRQUKx4veFyLOUmBLq
taLV1D847r+ALCj1Y6bd57HoE+1ajfElx4GZ9fWvduBtxt19I9v9US/fs4aXFgFP
6fNkSlv+Hr45w1ITzMJuc1cj7XWOvZMMUWVDMOImXuY+PcfP1BYElyoLsiIg81PS
8ZhRjnUuuo6jJxG94TskwksNqVazT30PMuYiiWPn99hjv7W9Mnec2rXJX4IoL/S7
upljlh1do/kKgNv78Bla3BlIxB/c0K1kagl3cInETcg4tEHVjWzT4r+azcQpfH7W
irWt0K3ZMVvAJS3PRIYNMZbQ9xBeG+ucnb1K2QnxZmNf3z/5GcOSwouFHa6HXbPY
ZqMyC4laawekt3Tstk9zCFIgdF6RMP5UWnL6B8VNnG5bnaNX6mlm4oAdIOHTs/2C
Njup6mbELNbgP+RruV0jF761Iaeyg9gLPWptB8gWbFAkdqqLtSeXE8dJniof4WDE
KQn6FS01xv2nSU9o3/qUo7zjpCms52JAF9auKqA1wi2ODK/ygnn9bSHTVLzKhlVG
RrwVNYc/Q2Tq8aOFiDm1pt0QAeQz5sCdit8z+1h/6tP4+XGzViRHJNtYRS6WsRgI
6dJfqtd+xAisZ1z4D0uqkXZx+2jaQMUIqei6JpWSXpbn7fLbDL/Kq4Kk7FznDGXz
7R5MOler3qjA/br2ooutTLr0niAj8hfdYooTFbiC6ddBRNBFZKFanw3tXTVuDYsU
eseABRvGJFY1PCNF+2jB6PZeMusUNbbNpjsMV8hD1y92HKubI79lOw6EB2NGkWL8
3zy2gMSyw5b6NYSOPrcBBwqSc9dDA18kGBEMoNPa7Ps0o4jjjKZfLFmxK3JuZP41
K3VsQiI0uP9+D64pw/aYVw4kpCRbvvj0q4e/9N5sAZ4Ct+j2ong6MvGYqfx99RQC
lYruA7K/DtS1XEKVHvN45h+vz15YLuanjZCbUU33XhAZK3Kj70eRO2U3Cqc22W7T
UgKREiktrP86z3l/pgjzkKgHX1HAlARR17lbgSEWgUmJ2VsGAgLIWEG3Qx1dinYd
9Kc5DLB34fViyh/trKTz7yA+h7I3jFTdG4R+ZPlRY4i5Pk1+CVmmz7X8klI1hm7w
UXtCcROkcI3GgyAi4NME+iOqRcbNzGR0xi47z3geGUP+WsPJCGJhTTfpvxRGuwsl
/knrHQ8wJeQgf9/d85tUNLkCc8CaHrCpGFTT7IGTvPj6jiS/2WPEaIuHE+wh1Drn
mEsDhRHJ/5pH6PO8nnN26cVqGD4bU16CtdR41BULJD1GVWIaF3DmDXiCghk1QP+H
/5+w4zqfBLopEH7yIJi0iWwCnjg6x8UN8FtWAkLo6RupPDbdPJyKL/JssriVDJGb
Xuf91RKKu2wqGxVC+isuNFAMMURzIDmcMI8oDzaWzPhOPfz7AtCwx3Fp9U5rENsc
hLrC5EkiI1eIQkRLcFijEJzcEuKja/idAyGsj9QogcwonEnoX5XOq7MLUSUSIJ/M
G0Tl9GpFGjqKZTx4jpEV6oEMjKEZ61ykNyBS5JS2uUEqUD/ww7BdD7sC2qFZlTEM
QQZrrCd9wQbU3xTcYt9669Y9mCP7SbRCR4+bQOUwaa0pSfwSviKHr80PUQfYMLBa
OG7W89Ble4Y/jhgc6Ni2OMYwhJVKhE8Pj+rqAyQzK7bcqWknYZql89A/sohlzndF
bvb4OA+NxQkuG1fphbgl7kdgKx4Phb4R1iZ0CiJy4nwXWmfP08HHYm+JnImcDgwG
iffUhyIqiFgO1DhjzXOSv8s2OoHR8/vOfukBrDATriHZOMJJQBkxoG6gG22hFMvG
8QXksRUaIPQAoH2E9Bp/OYKooeXJ2QNBdaQ2pXEoAiwSO2XBMwXExKpNU/+VcxZs
4s+8OK3q5Ro0/LB8B3oF9wIrcx/mK+cmH8Fq3PeT21YZdt2IB+XOIARhgX0xCo7r
G5pAkYDh5dHVDRgdOTVlya5Wp1hWJoeTRX1yRaK9xgwfc5wSJ2arOZU0n5GIAtSA
iyEQxarft7ZbdReiradK2SQ7uNx6bRT9PCUy+YlGaWrbCq0T71B7c0cp+OBs5LUn
5p9sG4LIZgK9qY0pyoK0Ryh0JNjXVHYad7wHJpgc1AymgkVD7tv07Fj0QgzkleXw
ZZWsciBYKGctJ5g88bCjoRLSqIyICCS/tBqek6lmqJbrmhguWECRr4EcJvyxN6xa
dIwt5bfa830ZGhqft2SMbA/xtd+iiyFARIRwyy18JQJHmcGisxuzk8oM+m7/I+4V
2pXhznf7p++GqMUov9G7FcXc4YI/lrgJHX/ndBSkjyn6EPmGvX+EnPr6gGgtIfuX
VOMVqOEvgwdmzuzH8jvVdj/NME9IImqd2Jh2bCZZ0mdWkrifXNOvuif6EjT9NEOB
0jKlzBZRU7K1o4GyVbvtL5wA3uDQ49BzchLxb/IMvaM+/lm7kam2K3XhLIjcWwJl
/Z45Nqj6TqF/WYn0qJa33fxA+vb6rqaXYP2cHxvSdjspqLNT42HIdjuJXOHvQTy8
bAW83+5AuZ0f/3BIUrboycjHot6giCOdP/kUb9zfb7yH67YRaWNq1yLU5UgZt/za
lKFYaMdRudDQkwmWKc3B1bWuEKZVSyxn92BdvuuaCjkR2cq6aGMeKt0aC8JuKlRF
35qMdKJ/yxs/2JvPHdgkKoAldugqhnkpDVDi61yzM8GWbtCwFUQ1ApoW2ExwPg6I
im4A8fM14bjSiNllJyYg7UfVx4nvQjsP+bl+TPGT3dNHjIgUp+g7fhaUqwdmH/yT
8uK/2pi2m8AWiKHiNrbLMBKBYMTYK1cunR7Z8PIYcfFfPa22F9T75vj/U/7Q0QM7
KKFg8o0OXIQuY+qsKvuyR8v5ctPhUF5TjaKWHL6tbxwfb0n07kNPz/rwxx87DWbt
6HiddctMQv2/x6mLZWBqeolrsgBOxo66EwNLv1I3iXTRecIZk7UXiQDZrzLl6e5F
umuIFokAXGREWbcFJQDJSF4cVd38p53eI8SyQqCA7ykWqy7MPgs+kSf8vOqrxCfe
pBAH6ib4KrXks5DbgvtfVc7rgKsWUyVUOAogs0+won5/5yxIGBOT0BpzL8BeYOqr
1kWgj3JraN1jTZwJkozFCW3QkLvkY7A4g+jTDBYqOESH+h2ifUArISbm5Kzd6TpU
ucerk6g9iCkv7Lhxl9IMcc1SucIgP14wXq3PLJn2mGEWfrs5FMScjIeUI91mHeYv
CFYO5YFUSNvjvRsFuvlibtLD9vI4M8//Dqm+9Yp6B8qMhtZgyQuYbD0F85IQ4hfF
KZADoTj/7FZUPLswDz41Hbne0+P8bXQRvHdIHUICAZqAh03EqFQDzvvOHK0GoUsx
95YFZ6zXu9rx69i3p1Ex9zx4jkazho7fwnxhB2VvqEYuTCx3Lqc/1APkm/XRXWg5
AUP2pMLC2eOxOyReBvUYQhH2UlS3U+MHmDhBEXwJWUkscPM7sH9aoGZDF0O0H+Tc
NReFXHqJ8YNjYouZLZwwr7X8Y06YosZJqbNDr02Z3LRakPTYM3/IYVvwsxgiJ5S1
Z6tTcqG0hhule/cjKVvPW8ncGNRtVq4+4+YK96Nc+hd2Rce3avR359XnfEQK8LD/
/naNobMH0aq3pTCOagj9Li3ztbrBxEp6h18MT15DG7zof/tnOMRkHJWnP2U1ir6H
HVPsf2MnE4cEYM8zaavTQFmTShcty4WEfLMFC+14niJVs18IqpXdxCdaZUM2uQhg
1NSBM31mM3ZpGl7tAq9R1vsVIQX4nENJN5W/YgOtt9gGLxEpFpcgB7vEiNCttw1D
CgiSnmh1E3VZfzDvlF3C1ZhNfVaOTMFqDWTjLkuZ0VoIkl/8A8cQ5lsla+k3f7cu
I62fobKb8UH613JO1wIuDjIZTHwQKiEZjvesQ1KaDQfdOFCT338pLRtN+mSugRR1
RHY3ATGPdqrLqE8ASY34LF+voHgTqkfowFk64HvSuMdNorKV9nQmcK50GVlF1QCo
eCQjyxWFZxt3++j2G1UrGX4LQMOYotzdUSlu9W5yNOe3SsXPw1N20suahBJqxG+k
wCTT8G1oJQ3+qhTebcPkDLOX/Qmft2rixArxbMtew9RFsdDJz0sp4Tqj8FnHjGMd
EHUuqx8jK9KIKcSDJ8cwZ18xKY/rPhZtTt498Td1w2K8TX3KF9LXnzcqRgd6GSMn
xd6+PDC/rB3qe33vGLt7jbxuYDbclNYPogH/OflK4s+oM/AiHzWU7AZ51oMA4EgN
pTEcQiMSPhBU3YFAw5PSfUAtjCrnUI59n6kqrAYYBNmB9ESBauK80/1V63Yq61Yc
MVlr9y85JxhUqRtTLhdLYL5K0Sm14oOGU4Tk+Xkk3/T7u0vO5h/TowV/bhKugxA4
Kf2PXLTzbXxp1orzX+DngXziHxIkJ7RjK1JISyvXX2DxJLBW/o5MufKyMp4eFe8+
7OBg2Drmr5c75DM6gV64rR41EwGt3JLcfpE8jXlclMCu7RIks/vafpm+pzNUuno6
dRIVlowhM4me8Qr3WmLxOM+t3xYf0OwCX39FLpERDe/2EOWWxCVoSy0Z7AWzt+j8
W3iY2FnbCSPmT8F9YcrBX3LHrP41ak0vx3FbO9QistzzgL73U1+vMbYq21TYsVMV
fvMYo0mbd+LiHIv2U/JqlaUmts1f8FgPvA8ZQGxMJOhGU/ePwU5HjGtExjxy1B0t
PbEqI1oiC4e9Yt8zpECsYNxnU2zcXqpf3K/sWSrpk0sObcE/NfA6m6NqNF2dCQ0p
my2tjq5ghRfbdOWmN/5JE/cTM5FHRRgsi/kM6TDL0HGjzW1NpUoTnxWUbpYh5P+X
iUlXE2YfJulQCRkFzDLNqp//N0zgBhsEVcGrNFsiYPUMAMEBoPhvoojuVIJHO6Qh
ZRXHRHRjpsppSRpkzVJr/E+HGy4JEhaSNI6pfgm19HuOgPtAtzJvGoUfdCXkACY+
yOQJ3fwgmfEq2sdTR8v2x2qRRe+Q8tZSCteqQdDCRXJCvxcd8T7zO8LhM2GvxdnC
5+lh7iK6trsvt7vpLz/KwcTjsMdVxubmjTDrZiAHY5I9PHHV/tDp05klW7Z1sf3+
7DkBAlb07O59UAQG/C+qVnBeUyKkHgv4iIpW+yq6AVgnpWaOANOdtkeEECdZZP2g
sFbhR1Tl0vKX6q2HnYtnvIsZfQp5vrPGElEVzuGbkZHQDBgtgeFddkWmSq7jZprB
W44CWQHlYSDy/NC0590L3y4BTor2A8QZ879pIO/kTitWlTSAqb1mvFShMeDJv39t
NjdtSg/CORsiOHZ5J47aeSgnY1JOrhy7Kcv6hpC3IYNT1pBFZAhkNy8nHgpoBdYa
zT0wdUlo/Tw2qwsc+FvbZ0S+8gkB0e0rhlC7A2Oa97+tOaACETlZ15h5IYbaVBMs
VWPiPr0hiB/BIk598r6ZNXH5u4TA/clPtm+Gm5YmC5/bgM6NRmGAGazVD1AxbR8T
SDhAssWN/oq6x2elH0xIJKDMHjT8uCFSnXEKreP+c4e93Xet9yfjVRhKkxxXOE3+
fod0nfHhA/IING4sz5Ly3z82V3VGUbNFla/7SP4zQXOS/XMb9BdwKrxHdt6fKP1x
6RXpDIG4SQu8aeT4i7U5/pB7RuadIfx7RxHmqK37A1GlpJCJ6Hmt3VT9B6GNNr8R
HZJegNv0zGSKYDqlRF5n4Am6X57zO+mya5q1MdXyzsk6TqDnQxUJGHTSoSBJzlbU
XEGadP/e/4Ah3rOt1U8HQqac81Zcea2aNMOncio9FKsx3yCXRFEHNzYPplcVT477
oRTkLi5NYbhoRI9kKF3dUctZRleGTwvATHPKNz4NmxD3jhrOEktCXjzzfaVezdjZ
LQeO86UEl5Jl+N3fviQzO99ULbg5Q8lQ3AzTCiZuaUGxDXPN12gM6wMEOlxYpj9Y
X1zsOAk08iHQqaGddL/xj3iuI4syp/gPbG9Idm2QuoEuT+Lk0jxwehOfCbuh6LPd
2C/WujtbwN+P662JXur6ylP0Jz3eSQvlbk42WcrZJWdkYh4a6HFftlMly5TImFsV
aaiSYdsGNdasG5GB30Hvh4XtMoi2PEbCMTrAspZfhZ4epiG0Dm3XcqwWrxsMo81K
DYDu7lYGwR3F9k63Hra60pRkbuQTG39/xHOJFrwCxVvfWgHATzM7q3qVz6WDDilb
yPJeXWja5mFviGZkyh9k5Q6H7O7ozZCTzqP6tA/xpaYJTJ1Ed2jXT/6UkNMypawB
qOo5QUTibOytdupDLW2gSMGOBN2lsLacB8yoPNhGnS0HExEjtSLWs9Uohq3c/nDd
pvIGBQ+sYaASGVN12pk7lyNoZOCfB1AgU6YfaNY5KAwjlTtkflfapQVvz4xpaRR9
eUFP7GN31nvUc+Jhp4UFZ3WSDK4Ph6M3CZWtlFREHeD/0S9N0Z2eW0R21bxHKfNU
kZy/FEw8S33VQp/BJCrex3PmJLoZO84VbsZnVuuBXaaJzE+gPiefGyihFcnRAFsL
N8N3Kk9hlp2x8yhUIke+eJiNSrwMfx2Bk1WJm1QaM66JEFCqDtUTj6SMEbS/dqYZ
ttKsYoHznX3hmkGqiZyO9VE0cycoN5tU98tHMOPiFunpaz1bQrNPco7uEZbYOblj
QNEuXKIfr4ZVKR0XVTPY1i/4f56B61L9dZwD0SruMJzC3rVNCLJVebiOZW6+xgkF
2uwAIDDYiTi3zOb39puj6k9LV6FzjKdUE7XrQZzCFdeHdV5KliCRhZpORAnLc9mh
SlwTB5ahiPzWSBd3fi9e+R6CTqJzI7/59TokEJKH0H6YILZ/bze3u2RlZdYy8w7n
IMnmT6LZKoY1VuAV6MfHYQF2tKwsmFsIE3t06pXs2InjPkE/8hDijDgiudPdFUwk
1+EHU3sfpooWishoCLFV3987byNZ3VxRIDMZhRsSvmvh9NusqCuDgsRwGsXkPNUX
59hgzmhnloYNEfZkltwcAPbExBjEKug3rOZwJR5IZ1I+ItRpAsY7yjrV/DMprgCm
eRk5nyfILihYFQegURnYm4g6wd0qviFUgwou/k/6BionLaDBzlslpMcFEWJhWkyA
78M8J8uZCmtz7abslYrL8AgGcJ4waZ4EVcshcWX+wQ4WVcPIhR9waa9Zj8H2LH7O
V8t5luDu8z7xfHHWBeN0MW0a4dxIzAj9lnuXwEidp766hxCa3vmm5+CapTPihy0p
lP+RodUJmm6n4haM0yepUGQeUxmUku5g/XYgJGstpxKbswqvtaMzE3EQ5iJ0K8V4
FHwHrRD/SLN9gT1pxYczl1xcFd2PsFAqC2AvusRtDQARPeavUgpjvM2Z4L0Foj9R
HLBTo9uKdi3Vm+6LCNAi/ESa+JT35AnLFgHRyWPhJvVqU4+YirqdfBIkBi64/6P6
Eev1kt9y43hk8M3zIJc3rLdYG6G3w5pQDNL/PKP32TJ55AUEUSW2QPgP2F003nzQ
EjsF4MKiA1FsHQUC1f21TJMmjrPRQSTJsP53WnDDeMcPUKBNUIdn7JXthbTCCqGh
YbCd/cg+AGa0KM7nvxSvqBhNCmU9wHgahf3g/E6RXyciqWU71GFkqW62P7aqyp3T
8alSf0YsB2rbNk+8QY6zXrXVx2ro00ijBNl7X2XTxW4J2r8Mdb2mvkv/zU5/MWiF
cAW0rV2bPh6R+G9e6BW82HvhJkE7J2J1oYN3TU7zbMzURcdiI2VOKDEldVR7VnN6
8CK6BzMEQltYB/e/LW1/pbP2YJnSxhWS4kaPzPe7rw0nyQfz7CiVo9fAmsbX+2mt
vZjfENgHuZXbgYLF65fEF2MEERghOLJvkAoMqCTq/fdqvVsOjlTeagyEurpuqzr3
KWbRWlJVRZfvvNEz4IU9hz2cdWchsPICI0IMB3klMrSHYjkABWAZYkfZJWbvmx+K
uK6eCHbcLJDxLjXMf/IsH1ElMe+Lx2GluJG8KUIGsMkWE0Noimpkjik49gtop9HV
9gb3sjE0gNvN54BDxdNf+BIygngNaQwUQw0mj+WiaiEwxVbCChdVIzXds8yVvQhi
g7m12vp/GFMv6jqTk9zbqrnC9Fbd+6CDojD3I3mbECaANAu7xYvrexgYhX4HzfMB
eNSM2dy2+pb50bM+OM/CrlVOE5hz0CLG3S/6kAhCr6ha51RzQGDaKVZR19oVproj
2nNqv8BHj2F3Imf5ODVnKP0/9BsqwC3oqp7qbPgJ1EJwEIx7W7KZXkcVZ4p/qnqY
bS1LWbaeQ34z378OhhGGyEAwFCdJkyotyE0/hrUQOrff56BAZseYjLM/JtWbnozJ
Pm9yze5cQm1e561ZVi17PiXou1GQ6u2aLuLfrc6XICjKPd7flRUtB6pAEcfv+J+7
UdkZgYrRmZQfsp+hYhT4UWRnIpMy33vPVfrZZ6HyNV3+Z4ptuYcBqcXDot9mNAuw
MOr3g6soqvaDMjFgAEuGRp5U7gZize2atpaU6nEN6NMsKKmu+fPJc80+T/61BqsH
017iW9z7tYOw3dVqPmpNod8ElLx6ydVhJqW3G1bmJkXvH0bgrg3OgyIfhyZM9ZrZ
j69dIP3XpJD+zZ3xfwjEWew7+vCkLTQQyLMpNmlwTkXAXznLaeGdwkAn4TJ3a4Rn
vuTGNxajhwuDOKxcBN4Qj4rHG5sD1EQPjp2gS3pTdAr0TBZj9Nce2mGocp6IItwR
7CBcIFiDYhnRP947SwTT527qpiYQDkf+GOmhuLcSJPdoy9ODRPaVBP/YsBXedYyv
zhqsW98NNydCZ0tOrDFyBnWh2rp/Vs9QDp+7gI14PC+mDR4etlOP9NMr2Jl/bxjb
RO5dFpeWwwzglcpWczTAFdlDcqoUyrLImZ1FjBy0W11PP1R8ohclHjnelmb84LUU
dSR261d6O3CumLZW8zDYub9/6/x0Evyr0qR+woZkMHlgZONugjp+b5Yl16Ir6Mpo
1hFo+G7slvwkp56tFIsb7ViQdpyPXsI3JZSmLpKiBMuZUBZaj4EsqUsL2x6g63jV
8s0OwTF1flaEMcc1q8sOiNjjBdTZ58sCXxhLlaKFHwn8pp8aHB9c9e0nGs7vmTrd
AQ+TSSCyrh4E56cwXMJyGYw3/z+2ydncNimoByIPjMs93muyRKKSaBaObKfQBqI0
Xk3Ao+LjRD+vt2VFLYK6iVgUYHzbrMwBHpAvy6sZnh452FaSif3FM7/kAs4rHW+4
HWIKV5O3hxdd3tecq7ByLQ/7Jms3S3yTenjJ+VRW4onaZ/5OApN+McLhd1wljMyi
/ZGRN0McJI1fG1UW+6jNzkr8C1kh+UmPF9ICc17beeQodGSOrKb2o5pxyIpPJrsA
DF2vyKQIzR9GsaSIXDZE1AgKbc6Mkbqy1xmj11DXLWHTFK5lsr61XIytb7+x63n2
5SCJwDX2wmI50md5hheL0GeDwGrgvm4re0U3FbwaanwbRlsNSZxahu0OUDOJSn8J
XNUQZC8U4fOlKd/XLMDyr7HujPJLg/EFBdgb4BtJuR6BhIOTXVmIHgnzX/trjaVA
8VOmb6Zi7kh/IymWuv57W/2G+S5YrRCD4BUUZ7MnK5Je0vdfxW20ZeSNc2HlSwWh
n0umcV7OtM6vLHyE1NdV+wRNN85dLjV1MysBiOGbIzOarA20TdNTG843el2HtKBN
LfPdNp8YipxhXvTGv2M1UAEXnQ4N6ERNwpbV7dgrUR461HlsxQox97vmKkey7QSN
l8UWG4R3ozELtwsEeX5S5lgKvFUHunAaR4k4YMlfJSsl7ceYOSKUgEVFheNgjAec
ww46Jb6uf872SQlinkZ4bOYp47BuBqExpwQ6HkPwHAMVyXyLzlhu9bg2PRlQulUw
JzBPyEe9DjR0tgslX9/hMJGP8KAZuUuJh1K7np3qjEy4m8XAlUTPtXlVAbm+xwg7
9D6yPflQWkDL5vvvwNz6342SeD8eir58D+psCRHJuuV6o5Wwb6JURXuJTqyRDg5i
u0ncJYe79gY5CpiJZNCT7Agwf1fQ1BD+wz/5lWxpN+oUlNC7sT7LV6JTaN4dpLNX
2Xhm00qySLpXmR4mj92oHHbtD+yUsRGq1BLa0ohMTJBg0aBaRlTruXI6OM4SLosW
+SMs7XLyMkXLZudmmrRxGcvShWh75g5opHgJMHJ6jGGTGACbyKdonF847KXJGDfh
PypsJT1jCPPTovUqDG6Qqnxwf0ra0zA3DB54NnMU20X3YQPcnjFiHVIA0sMBYZtb
zKwO9aKsNAQYByB2hL8qw0HGbmbcP1qqsfclaqWoN3XHcFJTT8rfBfZk2QNZTj1O
HwTA8ZifumdFcav6vGr23EEif1HoKrYWpmSNCiKJx4m3ZkBoatkqslVbRWSq7eTB
oZCHtzdX4Ud61a1fKRWHBO8p8S05OJk3gmJqMCjYGn+eSxxaJpMvakGT3mf+4bGn
3VE4+AAuSZe/hLTXXHCS7aIELDjHnAlZ3eVWlaX7zdElW8pHeOz2NWAB48BiA6tJ
briw84Lm4CJR9EkwAVt1ru2r1t22wegeVP8L4C5NU/0zeFlYfnFU8E+lsA2H4jth
DooeOp9IauWxgBAs54N/G/G3CuhO/YgxP71HMD0Uk8E4HWoiDL1GJP6Nw+kLIsje
ZsLeK4OPgFVPJE1uiDAR2ZpKxyO2V0x6kO/zXCjlpPfKfiBlyOTHGHOWNwECNiqE
3MW4FzZ1DN/AoIaKbHAklhxwuQp9LdSjNga13U57e1XyNMdRypIUmtKhGl7IkXok
3qAEgSIYLQ5NQg/lNvy0xZe4YbXLHKQuOVcTczfmjU1kzV1EPSzNbaEE+2OwhpYi
Ty1QqEJbHWKILycUpDCWNBlmxkkSxdLtUOu4NIdh5PE6U5+0rtiezQseofOOsVw6
QkVuOM8/69+a3q6pMLaSJmWDTdSlw79RU2V4daD7XXuCW2W/oCKTjtETfDnJ7E89
+EYh/cv8sadK9LZko5Teq+kLsIk7YboCvJhS77M9blK/cW8h4n1hqJfRlUBv4gQf
XWZnhllBZcLFYkUr/z43jolDJg1/Yg3xAw1xYxUOF6PYl0WRQFlDntSfhBumt+/c
0P/Vehn89lHcnAPg8+L1HPdpSipPFCiBTb1kw1gQ+e3StTvIorfJw5CJcf8Z0IJF
urbpdhj9rB1XPTWDUSGWENMkC2EyPvXTcDwQwz4Wpma/5nv8pH+QuzOCuJjeEljT
7YN9eAJOnzHFE4fnwz1jhMAesBjurbtFHfN9P7XYJotVAiOe7Z29E+EgRXzebLcr
Se7emrlD90XveEDlVZ/9IBSVelOaaQEzBg6GQ0jReDIPQQYm2REBNFuCFzdN37Lp
LZSzUjNEhHUwcPwop0uKAYanBsVTty8mUxnPFhUM9nxi+p8rkV8/iYtGg3GR24GF
VGhW38BeBYLKbuCcbKe9PG4kijHAB75/rQPasEMZRv3Tim/Ss+amG2NAoA+8bnOP
wQL4/3WSCL/9zBnW2i1S8L+6rpxkBGNpkAvXYLAFLqX2+Y55kKtCnCpGQA4XXQec
1EhPAm2ZJ8IrtjF792P0RZDlkH8SU9tsK4qvEL1QlXahe1tdtxQOYs/bZBfeOjOw
UDuo2z7svOhPAcol4kuU55B6TfZhzuTyygAONjdC7BUR5aaJJdBumiuJJE++4V/G
jT/WmInzkCfTcHx7AxZkFL01aDJb/aGsKP+0qROMhsjFCU+xbfmmNNGZRzSziba4
LHIGn1Fmog0Qmp4TTGvYAFk7tDRO/s/+cP45vrk2m1/WkjJyMANJJNq4zuUCP5hu
AelECvxIbzniVgvmMkUfShNSXfxncunabyvYTYliGMHTJCG2bAveRwkKjptSMdIx
REGUeH9HNwV76XsUgtHpzf4EjspvBA4Chc1o7oDqfn6oy4VH8g2YYu5VR8NvJjI5
Ugkgo2QiLh8jYvoqJzqrIatAOPjsZ6U4fOQU4FY4Vc2CQR3VjeRhe2pOHNNyAJzY
smDBIN/ZEhlmb7ZjlCWAocifxhAOHoaA+3VbX/nzwztCuAyyzACC0CjgyF7YI6mf
8rEhbtnkCG3cyghpxsDbqaMhMHnF+pqxCQQZyIbC/+3xJ68AdQAL7+s4CdJpuo4l
yv+Rb4sEItUT6npSHe+gSTN3RcBIGl1incLk63jaQOBKDqf9Dq5lzssjLYOS0Io9
AUukxtqsc9kb1RvRS+A3sLBC8c4S5SYQSQXSJGFZ/25fmezrCQMzIoKLF7Tgsmky
KhUPZCcsi1t86cGaYkY2RMLQCLKqC6zttLm0yHNDCghDXcJCW5mQekUTcB6bjyYm
TbQaw3u2VjWheZok/xBljEKoa37ZSOUTIDXiLg8BT1l30PNUD+zi3sQ+LkNCYASh
OTiSpZgBXRwv/cScPDK1BL1d35xH3ytw/b1Bs7W5nncHUBOw5DCugjI+culWCs2R
xe8lV9LOt+Nuf8KQzRvQyIf39gdjZuDhGuVBwwrC11oEZx/d4UMNhOy0LYdh5WZS
wgq59jtnFytZNE7O1JG1B/APV46cO37H7wIkNnZe5025ObXpytPCDNR9UlMTlWo0
lv5eB0E4LVlmNp40VoZ+XsPrmaDBGsnI2GcNnFg3vuMeFcQ2cvePLUex66oo4Fc0
8IJlWradvn+Go2D01952esPKDmCYsReIODP7gFo932y6a7v4+XFG1Kw+BQIIhZ+X
xMLOQTNJ8ukN/x+6PagmL+zPb5ywVb+7hlfCC1h29cJVJLFvJLAqx05k8G0Zly/o
E0rE20SJbfFljM24srZl/3raWbkwxyKHT4hkG/KFBMa+NNF6FkSJRPLkHLDRiMV4
kKeY6yDONDda46NAJk2K2luV+6re6Lx52NOz72sTss0D1Tq8icWMmvSnfvyynj+i
+SrJ0H7nmcJfg4j/zvgTtj72RS7Q4kqGNMH2jTePLKUyppQeMOEdtp9HZgJozkUn
REadNHh452Zwal+3QAU2g+fmP39iNlMVv2sbzIWjQjs/NGuGR5n6jwxU82krXR9P
dBfhRXWQ0wVsI1jHHpkDBSmMndUlNGzGkBOG6yQQanGXMUDNI/WEtx1zQRVJ8gd2
SINOayeQ/5aNnFmMwc5WnwGAVUsmAdjUH8HoPJ2bDMULHit0q1CdVHOvau7nM+CM
dBaXQxtDz+36GZi4m0TACHyWHLqjdoKz+HrKBkXfBJsaLeVU0bJpU1sfJxm+PO49
eUEQmS8GZuh78BhMrOqeMkAFQFz16n7/FPSj8QgSRF+wXTh4lKu9chlz8jnTzmxY
CnSFASFscCRnZ+9IhT+jHmrHBFeoMZ+GGJWQ0cAvLVQO/oYL03ZdmmS5UyQdsAIO
ZOYAhd/9WpFXXdZO1brguwUU2k5zJXSGhFxg2Rd+o4Gr0s7g77sIU7e97hUwGKSR
XymOfPpCbElc1WZ6/Ct6KJyqmCuIvMriP0tESB1pt3MuBcVyvsf+kvngWkiqm6ce
8cnpVX6N4vcpf7qCTZPL/sZZZ4g8LluWZoGS9VRgkYsYvASSEiUpubXzKuk8gSna
hK72giqPqMIytLNbUFlbSrgVn0J2gk6zV7xaQueR0EonNuGHoW104YCSuekQuv8Z
vsFZ2r0BvaMaefd+RuCLTncgfdCwDE6epeAwYqV2lBoqpT2EbBrj+pT4coMGrB70
G8GoCAOsrh3betfj6i4s14TTFQ+LS6HTja0p3SKFASZ9kuuCGBWJA6WuH4fbcOzi
YpUwsmuBLpthZm0j00YvNfrGKMUgELgFvHAkVbQoGf5LlmVHdmMlzykuM+yRVOep
P3+gyUry9P1Axebgtv1yXbQxw1cDuS8OrxpxmUP153SQkSdCY/b6eTMgR61QixIx
ajdYV2yadfjOCrLYWrWNxTSr7M8HOBwxnres2XIp3HWH5bDGQRuCs1JEXJWi8/TR
Q45oigN80CU/cPyNHSgxYHRuPHfL1Q23QIOsEi/P8SjY8IzPQDZBYco6qlsdaiYg
414mj6L0/pylqJxjETpX0ZUa+WDpq0M9hgRuDXrRQ0rpTl4IS/HyrTDA3OMykVCC
TyqAV9rrrPwHXniuv6NQHBFLQ3WYL33bAbr19CLeCQM7u/CanKdHjdQxGxwdBpwj
pHLa5zVDgU7y28m0PA+6CgIiesqJaZmw4DT8qbZKEzzhMFdAZ3VQRbDvnIKXBXUU
vwH33VNppxQS/jUaaAeo43VvJdHYwjvFhy0HQnI27C7Gc6Yu7hSbtVx1Y8b+wxOS
dd+lVWd5560ZwjXnajTMT6aMWfUoJ+JocwVkBAZmdcKNucxP+9Y3skBYlHuQJ1nK
mQkz/SbPa3WNvtKCy41b3kveAXu7eoCJw0VjwUfdnFC3Guav+lrKM21IXh816lpr
xuOos/WDaqA7sSfZGYXcNggK0RDf5qaMzmA643tqdX/lAGejdhJdY5D2EMSebss7
eSpDkL+1J0Ik8GrCn+sR7/vzY/5C1LZf089+DI+V+ex2I3Q7yRO7tm+kbssI26Cm
3ILlktLriT1sUP6AsQISX/2h6F9a5pPzf/wOxrwD1Ywl0YtYrwshHUBZ18F9Lxr0
Bkg/5NbfeJRwNyqjZGtD27pTgclZPsSI3kjiEizumLsc1gcqwLcLpHch1Ix8jh+F
8GFre/6h5DNxrt0kG3hN8E9yLzsPaMQ9s3zHhMnSbfdO2k3aKBW7zhxUa3wow3C7
BSyLVr/rpF63g4dqGIaRDyxuYDAZ4uxQnZrdd6iTtin3uVG+JRzySr0RuN8kCfvo
2e4wxZEivc5LOzXZvWkQ4wv0FIBqxgGWyGnyoFBtBwQx18glwXgVDzvjikrTq2Xv
iZYzAwhM3wvB08lNtM+MgASW2Q7hngnz53EXfMXyGaxOq6SBm01i7rg7oFi930tT
hT/LUoFEzmgoWHFvorDWmG1Slr/0++g7YcoSOHTR19RojMFzINDHBLZW0D89pFu8
rcqRj97SSeqCtjCV7KewwCJJHPEWQagU5qH+3Y3w6pBgJKWz5zzI6oW7FCiwjZF1
ZK+B+UKm/vmHcOiW+1AYdmansPtvlVA+JrgJ+JxjZ3sCRScLFQgugN+dq5WAl2P2
PIJEK0e789bYgpxSH7Xnz0Suu6WY7x19ZFVG8GIyGbZCIcmaXdtlht1JCHMw5fUf
VauuBxufB+RzjoqGbHGeJriPTLy+cpcfQandVzOR6wDiO7tn+PdnZTvMXxuPS6f5
LnOFVExl/3cIUBXw2C3G46wN3SVmMbZSFndCNE32whj9pdxNbwXwm2Mcg7rORNlv
Ii8JnmSqwnvT/3Xp5dTPXMm8l9W3797kYpe9znWsZV2N2X3nC/gmf8SD0cIarV6t
82qEaNbYXnE6SiXtM6HhDEgT2KXH3vZqh4flzAqiZaARJ3Aa0G0iKHgwh7SXsyFV
AcHaBdM0wOOPjl3MKK+TvWuEJXT5G3iik10T1EMa95jnRJPCl/NHmmV1ZTa0hpb6
X5vZQvcgHP0+u37eqpCweDvUWVdBXRSbMjSFQF9TSyTYiiSFGoH4cb9+HBHKcKwz
AfphiSwqdEzWcz7XnevTJrCs06SC3pGHRuosf2hHmFyv3PIcEKsJY6inVIRY6N1Y
7YeWVHR0Vgq6OlGMFa7Ztm0Ltkxz15mFuSe8LA8bczEx46CLKrrcFb08Ug4907l5
T6Zz0kiKSXJ8yQX+LgoA/8KBpDmylKSETx1Jh8Y5qTtNclKWQieV5eqlEAR0FnQ9
taJAvRGSXFKEPFBshOEc/SY8jGJ5ok8nZ/Vkegxgw9DJQWzszuA6ihwZIYtiZeBH
5KrhZn64Gfattgg+wyVFUmkY2y6eSSXr0Yr7spW4PQVvNpsWkiB98EX4JB6g5x5o
9SWu8VDzHQ9fl6gzSLvTbLgmhlC+HbqscKNpbVeYn7wVa3CB6O/PC2axtgEGc82z
H9Sj2fE3ogeRzJopUVGm3viCPld53KX05LtUg7BP1N2T6w230rIlCVUwUTPX+XjQ
yG4fQ+GCjRTT3G/ebAq3mx6/JpJbsVhLKl7QcwI/4YN6YOOm35JLl016QeJ/jNhl
+F0sCRImaakNjswiCk89rh84WRDnwwgQgYwFaKNAOhyOnnFBiP86FANMU7h7Nmax
2BP8HBs9hNPat7ECa3+9YOv/1+uffVP7o5cqREiB6Kw0rcEBAhv+3PYq7VT4MBEA
z3lv+R3mPjpf7GQJirPILejAL0kLeUWHAxlh/D7CoqzlPnI0io+HVbg2vRBk32dX
93fINrELPdLDLRU05kLfYaX749qxdHrlJgoIqtkArmDeFAWJJJdpba/wVy7pyRee
ttAvBetEBL+y+oZhKAVRs1lqAM2ucd3bLGoo2/0elrxp1jdWSCMoR1da7avs9q8V
cGWRgN9JzrveMtBeOLkA1X5t66kpfZf60mGC//YFFu2Kz+1xMc0dDI8GDnFiIBxV
CfszMKsbCxWX2LMn1snIXLJZP1UHlf+3/a69m4tyP1SH7BmMpn8HrUHHhB1Bwdbi
DdgkmVhR8sKemscpASh/acm6i+VZkFDPqW4FJzFZECBRsKonfBmGfOFBBsz+GjI6
YS3+Krng2KyUsNsOjr4rShcofqErYgLJPf9wfPIFqRf7g4xh2VWSITBPrVNNKmMr
aYYUzdM8I+d35mFrpam7e73sKVKw8C1yJcRBxgRYqxqfsbjIjmTlhikQO8Q2Zadx
kzeAHrn2keKm4q55FNBaZEHCUnmrL6fexzczZnuiaddr5XeeTsD+n4gl60as+bb+
0cY4gUyLD3NExceBUoYiD5ZgvE7z94W60OmIjqk4OL2QDQroQLC3p+d2OCkFhD/L
u7G9/wSBTPq+AM7HErzNKUegxBgL8iWllhlmMTHpivj6kDwLEbRFuFioWg9lzZzr
itaf6/PuLJ5V7l7huN9O2K7mcnu4HRKUTGMVvnQ/I8/eChpTxJTgkWmJhTes44BI
ZWsiswrMDsl3s6ZSe5mAHJTQZhpKlCtM9QQVcdpUFXNWT0LHqDt+C+acv082vR2p
m2S9qVeOhf5PS9xm8rqs5NSaHYSQSXK7CDXwH0ZipC/79fdihhr4ZqGswSWSXPuR
VdMFDBo/Jn8irEF/cWoixcqmaaIRmlyT5r9+RYTTfIJXC3imGXSM6az7TJJMUsY5
/uG0pp6SOz/p0q5CSM/3sd76kg/Qv1XFWcgQW5hFTgSblJTlr2okytY3jkJEmW7K
pKd6KijOboH5PGcJblbHTFIsZO3kirtSkZWcf2r0wKrOJAWhvjoTVaxx05T14wLe
Ja+EUvJ9S2fjjj5GXsxAfv2QkVZjpg5QvwFzppRJcb3nxB6Lc8yLjhn1vGwVUAjN
/0zTCYrrGFQPKkJJKNozXyH+3Ss1/ZXinyITdRiE/RQ3INUQAzp+TJzzLyZ8jHAv
XRV16x5JSQEJH3z1TMoNRfNruPXrdvdPwam3hl9CC/ZekwyPMidXsill09q6vyPM
Z697/Hvwf19ZqtJyfZn2VljonQgMIhMTUgCpU13LJ2sPX4gSqp3DD+wc376Fbgf7
/2wdrsV59hGKkSeqW8pg2THuwskUyVyCg1Pv2DZgpusvC7YRU+jLPrIdu8iwMHmj
hgaYig8YkAPW7+9q/LYL8PZfsouF7TkWxihptkp0F9DZdStLLqETMdZp06nhJOsM
ofz9sh3BrQkfiQniBRwqYFLdA87Ed1sdW8XhtWPAcLkHkU6ewWLPDFSa9CD1Jxe/
GiEiowkffo0qbFD5lbcvnMmNeuUDtW66j16d124oSJlR+k31/h4ZR0Xymm9kUVYe
2VS+F8hcPwkTI7fmKOSmFaGnhD0bgZRE44DOIzqwKFqK1ywR/qV2/lCqnLpByysN
rftmY2UzqS4lqQ3f+BHYvI3ZyLzkAWdLZqADo7lZ9jjKUbdzWVrrElpB6GyUEt6a
pvhNFPk0WwSPu1ayULxP7IMBoUiylrWX85wtDSfXBHK5lD5PuN8vArWXbGyk/pL2
w0kz2pSRu8m28xbQMqafcW+1iOQ7GqBRLZry2QZWzj6XR7VyjdjhJ7TieJSBoiu0
ikBd4+emB/tlnw9p6hxq7jG0cC+E+TDZRqEnzaBAHL/qMckecSPSXiKN94odngeW
Laxs7+Hx8PYKI3b9uMghxryHyAcCybFCPzbhFocv9sD041dWWeOM7Q3DfV3DPWIx
wjx7HbX2+i3MA80KPocnSNf8I8+m2utEJywjn79tGyoGzBzPiNpZmsoqIBNo7zFW
72f3Sl4f8KnsXS2rKY3BY16+vk8bUxadAjkuVIvw4vuLZd2H+V74bR5dAbod0h1N
6n9jezAX66qr61S+M4Tr68JsKa8Fj5CRnHNpKFohQhm/i1WsPAMy4x9FpDIVZx6m
oVFiJIc8ioUZdjAwAZ1wx6zyAjtWqKN2bKq0RtOwkc8lOha4Ny5Xc7GpSzJlSkBW
sX66y9TUYpmRc3S2Bw16SsxbXziqFEihBMEeQSVJUDkaTjkzTl5Z2Ba4JJ5BUy2U
upOsKrcIOkrBAJOtgg/wB2rfR9L87CTV3VNU7cR0x7SfQtyFk2YIXQdTBjZ4h1Cv
jYWxhpxGS6BNVPMOI5k+ttohgFkMgQHjLnTGO1bFByr3lhxUcVdD9FhCGp6ndKoO
cEeN53IUNeOfJx29VuMFTh3neMJJ58k0zdtBHjXpnzl/w7mZB418So2H2iRNE46g
3AVOKaHJpJPl7Pakf90TIMFUPsRgx3gZP80G+fkIZoQIF6f6dIWS9xPrPdrqF8S8
2GcdBYILsG5bh96lA94Ntnw1vsIsIY3+hKeAYVYeq9rLUxOC2duiTyE2E7cfynCu
At2xed5DT6+gjiSP5wq33S4ZfvzLjQsIEsPLhcZJYZe8F7TwZiQK1jV0WIWamLAT
9mp31cjvXBxB6HhzlDggiM7PzpU1spP+AsfdmNWdtS8pfkVD+jjQf+QhExnKbEy0
XmUY4Yh9Bgz52IsJXms8z6xf+FKuV+DnPTxRebQKsxZOySBO5Ym2F1rdAdD3192J
mTLNL8egDMdnUe4xgTeNAqHp6tlsfLhDtK6aGkXnUoBOprK9Qxn9Pq3axskxQpvD
7WFWO/STeOgzAbyIWC8BfT9iEp2tzmAmBIriSrqPO+3PNn7jTNzgORy9CHHD491L
+znMLcBfQ4zpm24TGaJdyNMVHLdNEy5hhOtGPrva5anLWhCSeDsfCk5MZIky+IVB
dPvDR6hkrBRXkwLa4Zn2oVYcUViF76ztbdyUbJXhBFqBeszvTjyi6DdjfG64uRRD
9D7Ou5DKCefElYUrCm3K0zsHEr7pwVDEvZ3AXdnDZ0EsUF2FHaF+uEecZIR1Jp3z
oMk62fSqeW36Cd/nl80MWBNdt5AO3o4+QQkRj41NrX5kojx28N67A8bNGuLbWdu8
1mv3Kfg/gvJ+8XU0QaWmqW/xV2jSLdgXmfJvwPEtzVZjiFHFOfopON8EUONNpqYr
8QZPEtfg6dfIfW5V59WOxsrPbctqDHBF1JzBCAw4zKjfRkytf7m6xmrlyHl6rLTZ
aVJYZfrBejg2pKVsDkpiaFc+OnCL65pcda/YSwKz1HevclSSgqtke7z41sc9ySuy
SoNHMUHyJHoThKmwdGKGZGqDoJsfKUcXx+S1uGj5hDUWHU2JjhTSm49eiZl8oUup
ysIdDD4zieclR9gtKJtGylfdE7Q59FUnDtRrVtfgjT8u7HlsuKVpdTCylTWDSJXf
lKrigcxFD3F/XiLHq66Ht+/g4Rt68FhS5YOIXz+NlKqBf9PiZ6jar5hLCqhycY3w
TTi82keBdV44LI4xbHqSTxK9ZoOO6uKJJfSkN7ehAFMglMfUl4Gx/9AAajzMKfvg
FBc2BGU861YbkM7au7IC+AzAo1TKGv1oXSElgjKFwoeuyzgXfX9Dgf41ayLrnlUq
9tt738lrxgS8p/a/IDnP4/kTNk5/r4MH1zxWKviV7FqTKKz7xZDW+qZDVMDROhw2
QufKSGDWzbxNywQrJzdHTYfOip9CKqpSbVmfd0pcocpD/mG2A81OiUJjEsNmFr6t
SszXZRRTAmjzsyFKhGWeXjVwTK6yz5UjBpBh/ZPLNBc5hfwR+bQH/DnU8KIDGzFi
/vJutkNP+qac0bqilC4oegkmpojsc3cdteHamQOeB5Uro1KzEuH7h6zChof7slTj
E8yT3AVV6EQJrH3KcSYzJiqyMsG6kHKIOG7G90mQh8+owT5Wv/O0aw9XoPdVQ7AM
EQ28O+oDf9FeUaAOiAcnWdPHGfrL5NJASxYAi9sxfDuTVXzUywXym5LvTxe8E3Ko
oBoREwys14GiyGLYgn5CYpHwO0hZVb/FwoiDRgl9M772l73NjqdFIJgIo+rsXIf6
5tkOJ96N2IfJhbFazBpAf0rO6qMRjmP5XsrshJpFSIkLrUpEfGT7F6fBxgTO+pMO
gRRyU4MyEjl0Vll2gqXbs/tZdIMbh/TNXNT8Ofvp6pkpGPaz/HctLG8uxWEWTarc
I8jmqWdy8bVhFfcXA8MBWUUvIEZ+STGTfI7pFXJ9wrO8iUiWHTPZ+DyuxVOc/byS
CLNaB3CFvzaEKgtuJ07NLn76/1FSQYasC16WZj991IOK3m2OkQRZB0/JAlXREyIR
fAd3ordm8XkXkliSw8bgzSnVoAxPnvWLXy+lyDf9ZLCtZ1+Hv2DKRzfA1y2SA+6+
HGcOarKKw6fB5701kCO44MJ8ji2LlITzET1JBRvz+WrhB4ttXmbjfl7IX6BZL1Lg
YOcSCtFrDeaHbBefVc3KU2kaG8jPI7AxKka8poDI4s2ZqYtTZkni5JoDLsf/NvO+
rZLgtsP4qfvsbpLXNXrCeFuAL+hT58S9AOZMHDVMwqkcVZqen5oWK5KTVvMglIDQ
aTeGGjqlAF5ATmOqsZE0G8rnwaeh0A2au4w08Hrra2nQNlsqQ9/SzEJYq2l7O0gI
zTs9zu7SNumK8CwvMkXOxynK9bSYG0Swog0KApaAwz1ROoA4HeDgg2pQWzmj0IlA
nTJRRDoFVIfm7KxKjKrkIz8x4z/og/5P16322muRmF9OBJZ7eJgJ5mQzX/GiO4n7
6Vizdj0urtuzwzQ46tienIxbsIj2Km6FjkJT5Q6SDBBrfCWDJ/gytL5eiT8qqzlU
AH2xFNFxnscYl+1gMYDBUkfCaLybVs+PlQAuZHKU1zCiC68cvHw5Q2C9g+vbzx6F
92xkNcJV7Rh/U2JsQPRAc2u4aFbEQVSkkSPhHt+G4ivAA9supbgZGz9MwY9RW/KY
ZrMOoYc2BJmjYg2/1Y7/m9aS+G42jZciu4AB4UcdnYuZKpetjSWUbLiiZ1FlximP
ZSGr094I02GqTgU3NFGJPuZyBmqiEJq6/dQYlBOoDwmrkYW6ptApEBATPhOl6u8H
koLybTcPnfCd6AbqjdoiVzyGZMejmbxqaZAv3fRpzxukmat7CPgZQIH3qXMrJW7Q
vgjePDZG1+URtryC//XOeY9bqk/x3lnZosph7KQQgtCA6y6hkCXbDEkb9YUGcq4g
TcbaT/HfdA5MwxPtLrKKZ6UoZq/oF8BVOk2gybFsK00Ro6PDYGOby5R8vp1jPuoO
44uLvknPmzy5rNwhsMN4tBsFkxy37LQr8fScjIJvAI0eqAaBdIdZMJB46pADTIwG
Dljx+3yzCZscorMbKnb05QOujvey7Soa1kZMDHJc0EmEq3lTWqQMgXMuiFikMwaI
skRcKSuJv/DUPcA2AhUsWWyR4URz5hfQXUSdWCQNt3DsufgSoRtaciGBCFcX6LTM
ASxG00fwBd3o8MXBr1SWDNeyBvhyMJU9Klya83gzzFWDMKijX4Z5jkATfInaIFeV
jQOTKj8rVeX3B+o+5tpYj8n0esFiibVk9n9y/ezFFrrazjSGGigplHK9j07GKe3Y
6yD5K7sUyIqOAqs0NEHC+hmS2vaRdgbfIQDz9d/9k59T9NxML4fAx6LHVu27AEvF
Lxqg2r5FClKLVckbyDCOuJ2mXvTfHWvGDjBAlBzeCclCnnssLMBJ5baBDom21tr3
v1oP36eLf+4AD4dpyrHsqzikmqiDS3q40nUFMgOW+e8x0RZRfAL4GfC+Zp6nhqb7
+PcMNRKpZOUHHHZrvnsrQZq7vwdkSLqQn6uS+lxd8JqsdzrnYxc7JhXVWTc2RxPt
/8T5h2yjBQphMoYEn5oY5er9xtZwE25hulbnGPAcdiW4JrFGOqzd1xeZxsanisQ6
LnoVpqpgPFTC6oRlr4fwgiYJeoxaonTDY0MyUrQE6PM7h0mwftetSbmqTVGnAOde
DWVm7RrvdXSDwGoztLIM+KbgEVRw1Z5G618NLARHahg8ybtYHrYix8KCDu7wIX9k
hyUmn8XwDXLGnnHN3sD+gMccU8G+3J0vJKrA7v0AjmHKTD8DcMdpEHr6tmSsDC51
1nxad4Eh3PQkvPiE1L/Dqwdt5j2/GJM+W3RmSsuu7IE2oBAfVjDA6+qL7qEHQ7by
reStacCEB+ze7V6xv+Iak6CKFPH1JOsPZi7JBBHseNc/9LJXeCEbB+LWWD3mbUXa
RJWbCS9w+b/xYmT3K0YMIeXFl8on/aMWHLwwVz8GV50vkJY9FSIAuWLFDEfRvGMU
sOQ68KsqrRLrOAJNV3TZb7HgDbS4v6T1BgTO4OOshSLNhOeC6AjupsrjPLVa173H
X1xp7UW8Bt/r0zZGKynMze8D/6woidumTPouLLW8VcLUdJbGV6YqkbclD/8D813G
9zTs7Ymh5/+3rNFiHYFjQqDuQYoY8j9pdbPrdDOSSzT5Mxx2SM9PJlgnODc8kalQ
emTISnIEWmU93r5Zp6l104eKnWaeQ/uKv+Q2Lv0XEKNwUJs89nKbZhhpc1a67S5h
e1fNWVv1Zip+Cxd79KVdZxG1X1/3Je7r/wVNsaNRLij9uWliLJ1biKmd+6/0oI2P
MkFqaQkRvcOnpM7UxULkK+p2/jYWFW993D6LKVpmPoI7qNaJHQAGP3j3qBwCa7kO
hIpLyyaxGlyOtHFWlwgUSrJMJinz3uNfbCzOb3KOKSOhKJU9zh1+vdqgJFYXTJ39
u9fyRwTlyYsRW4cUr7Mu0rt4i+hToTc55kPjpotbnDKaa7PPI1RpiyIxwuocOlbi
IP1w4bY0H6546jDyPMz30WN1uFMAPUaitCJHFxfLU7Kx++NPlDoST/utnoNagWxX
0Tce/mk/R7KxGnNwyyMHceHuE1NVh/LCEVhtUWZ6GxEzBhjBW4/t9HOQuOdsFYAf
zt9GtWFFVwOzw392VHfiY0Q5ZtRbwg1Zo07gakM5Mc4hWQJWuPHmFAH1+Bkm+5S9
qsblLRxFtyCediJiQONfNsMSDl78DqRuKnSKWNUijKjbFThhfJCmKrSk0byIkNC/
wgs3P/LT22wPekOGz6xhWdRzoDHxMUy/WFuv+vekETol9fbguos8yP+K+4VZSHDX
n4ZV/3Kt8/vmx2rl/jI91u/vi0k6N9aXtYTrAIHY26AM2KYuAX8FYS6867DsDqyD
KOaQQf9Wb1CsiR0Dy7OwLrTUiXN7arWzc6sqoJ5qeHsi0sKDQSz5nknezVixzFWe
uX0zSurx4R7tJG9Ld5alJpvoIROQLeOgrC3ajR+IlBkQ6cROj+o83r2DtDQJ6L+K
JRAxdGPs1r1jxqx/3UKhjigeK8cLvCS+3cnpDQTJ9sMVUlEqaHpcUX3k/0EaTfmS
dGnJfBtydZVNA7Zqxf6u5s99uQW6l/1ro8GQ4OU3g1DpJ37ky+3sJ/az0MNxkdiL
lRWb0yeCTJVT2zepTrSU2c53N816qJ3UXYGmoD7K1lY/STAYgGodHh1oXOS9aRWI
JZ80CUzDdrSlZJ4Bv80bgATcUPHWTiDOXp/IIpxSU9T8o3hBhuC0wrnnlok+jdYn
TZDh9FEG6jo5cGJRGIGe83+buFexedIO3mL78Egq7jvLAIHJcAw25E3RU7sVZp9T
K1eILT841TW3GaggLUaU/dP3fhjXtynCob/E0i+a1NcXO+D44smL0o3zhzo10ZgI
Hodyu0Xg9xnCo7eHsm7jzgBvTBjOTcuP2kC56nSYXLIu6j3uX7G2yrVu5QWgq7/F
RS8/M8/8rk5POcpWfhx7ZcBRFX/WYUN5KxeJ3aT1SUN6Gr25OM/nMzdLQYj6WSvK
I1WAE1R978jQ90Q9ttrFrjwvOiiJWL9gE+jo90CTnWIjnpB49TtCzlDPI3LjUDt8
vVS51jtO87cPQsMR6VUNx517ueKznBV2Aid1Dg+litn1c6NM97XxaGrsV+JplrLg
MoURGwtWkKHxzQ0LGJhZUA/2ITArLVTp46Wd8KWmtczfW7y2o+matkbpF93gSuR8
/pkIOHUVCOsXCFuzV0JC27sd5H/zGqgRiPVOYWnbWSdRsTh/Q3fCFgBOgj9+7fpk
IfUYap2U/4wD3HH4epE8uYygtN9zPQfC/bnW3l9XNaP8gS5P7yu5HFhxb5eGMwjN
whtci9IcvOvWPT3i69JhY3d8bl/8NVPvziw06G+fuQX180KuQT4ZhTUdkKqB2tLN
D3M8eL7PvrTp7nXhRP4kM8udJTvj9o+pFn4C7xO+Rgi4hmjT9Iuqsm8X9CWQGRds
I95yD9VHqXdqvxbAJumuNtosHoTzYfEIAS4VJqVylhzUiEgKyuJPVFUvIPqfyZ++
kHmh8kOQ2zk/L4AqoR1BZXbzy5UDwRkXSjbdYKAgsz8vQVEJ7t6osgpHbp45xJuT
9wlFk6pL3xBn8XdXPxEPbeg2sfzYyC/9NuKrVVVkEkrDprGJSIofhfCxi/QPcMHa
LfekjVmY10utBI9AJJHdLWX8Pkx0ufiTCZKv5D2hcY/C4utA8kKsx+bZZ4ObL02v
Ke/wIPNKdM3QnKb4Y1of7/hLoc9D5xrfBoxbVPip0KtcpstVPdvxatoN6x3ADIC5
UsEKBtmxXPJ78pacxmKjPsGdLSiKRqXNYPl8uSRk7rOvp5hAv6M90Rbv+YJXMPKZ
Wu9IvFt+RqtDo4msxE6nm5wYdU4L4s4prEJl+am5C1PMTfkgEklyMx0nnUQ4/W73
juq6i4sxuk9iYvg9+w7xQUgzkQhsgKlEZByIxzbXmTsLNFb9x+8aRvCJh99sjtm9
OTM1tTCFWP7par66Au+/5CfSZwwl5qeAymob3Gnnbpr4owErlgB9y/hPTPtBKghi
mOMJXG0Ai8A8fzIfERAn0oK6BlxVgjdpK09t5s3avHDBcpNtsec118NGxAf/LfPD
NtwnOJZ+K/o8BlC87bhbT7rubBqxOubQ6sM3rU5fBG65IpPTP1Ch9XJYn7anyIlu
mJefCRENFO++9xV15Hf7LK+zOfqT4j4aaxKXi3j9XUOlzmEdJFWvqqHOSMJqgMbq
+w8dk06XlcDOkQOdwI1MWKKtYOx1nnG9LCua4TWNGFzrjND43WCplJfpFgadTvHp
GYDl7XNa0puLtiKmtwahJ9yKQ/m5N/Vw8k6O03zCi7puC/p9+tmwuo/guZUeu1F8
lhuwDI+2v4JY94RC4sH+Z5AZ1+HluGODlO3ueAxXYWT41p8kP+OMSvm6347pHNmj
ws04YdaPKCbcpQO4h5dl1M+yTfKnqb7ir4XA9PThf+NvIGPhIdOsahdlcN0eylc7
dDMLAOu1aBzDAinFyefvMJeX+QuiLGffXW/LF62fFmJx0bQXREcPykkf/eoyILTc
BCe4T0kuSXIdosgH4S9W0+0ZykHLT5BezChsiSVL/yziZfHE2ATuTYgO+zpzaxZl
QyHi5DQFlVHmbrTEoxqPUtQrVgCllt21/VJlGRohOXV9VXF1/SrEXqAanErdna+C
8DJlN9yjWAJP39pbWaxfbnDoAyQwesxvuFX0C4HErGZByZU9+5O/3wsdOZGiykz+
9b6gRHPbOUrii400F5YuIPc4O3YlLqckXGTUMM8FK2xK5JJb/uv5MU6I9Ql14XWm
5C527OziTDFhNJFV5ntbBkijxssf2oAfb7L/yfel4ILzH89vdsMZxEMCiNdecPKy
s0sop4ByOWUchbQy3WHtwEuNp4HaE+dJGKjnXBOIJGObBgj7y9bHO4dqRW8VQDeD
52Ua5dUon2l2wItRXEWa4hklP76f05XProwhmLkzeES37I5XMi2HsreCt2+b2IKj
3Jestw5NsczDa62jRJq2LN6B21DPAXnxXdABT8RCvCq2H0O6CpqCJoZj7PaqvTU6
gOUfZ+QWB/tOEYwgHeOKo0b9ElGo52ckeiYH9HdHNpyZofiGsm4hTQw7ddXBBlK2
wvpiPlpVAAxOehoUqZqnKu9+NAcCkM84xARY5mQZRIUeRie9oMoO2fjjPJJFZrMZ
MeIQwWCKCz4DGJyJplH2oUgFgsmS/rgu+pdi0MM+Q1WqOn8TpeRGItvvUsetj/Ve
I/Q//7Axqr3GmCq8wGci5i0AD/3OmzihQ/SmRYUnFphnuQgbcuTev+dYOCrz3boV
7lyMGajhF6xAgCkiQDyEeFxoyS8Ms+VZVLjx3Ept1hN52bQXm1KFUaBiiyv3o5iT
J+83Hu7sLZ0wmfKYZ4X4PQmg8ST/3N1yUQ5k9EmCYfYdwJStRp/eT3PedXZuLrE8
bCoHHG+/XvKuYnGUhf6EtKzlNhV22AxYuBGcZ4lsoZ20YjLwEAeDa7UW3vwn6QUz
xI9U311Nev/zSDKia7YeYtQkKXALDziPZs9vIZ1A6XxP91QrdWTEpVYss8dKMCfZ
UXhaCdjiP/3mUxq6s/T8fHJsuTY57jcUNcgSZE3LiNtAnZ2BFYHcbP3wTdC2CXer
M/TjvVwpJbyGOUVa9n6p0sBYXCRXv8O/J+I6/bzfeDwlCDUgbZ3UDBhX1WicStNa
sc73/zOx0uHwd2LxTRpvRBzi13PsGF9KK1FYr0zyuvjtPCoeCNZK28anVtegVxcM
E8+hPYafMu+IsF6HFfNHMaV4MrSGYYTx8hnH/2MSsyXGrZE71KIKCZ0CrLLiJSA4
FJDbDgqyuMRtTysLkzcXqBGLo0DEvTnFUQ+xGA5YJIUSD+C8Zsl4F02KrG151uEW
s4No+32KZVf50KzqlzF7cubMUOer04+CdY7u3hgpNqUNoh+XlaLD088lqaUmvhx6
EUI2pPeop+6g6wqi6QURDZqzanxEdsUYzRLJmrYLxRlYn7ifuqix36oF5+6a46dU
lJEFywRiEsw+xIDVZIFCCPxuJtwlZHUtQGDL4BcaR2bzvQpyXpjI/PNs64Yl41fu
fFOJslHcD2sV96LLKUudM804VlzG5mKipRhfI67KnaYlHF6P1hN9BiHYx7i8z0kC
fJi3ggN6FhqvptiXWeQ5sgeRSEiFLhOz5u0ARzCM7HZzsaZRLl4OhFrK4gav2IMv
fd9yUzni9Awu1iCEdGTJ420L5OjBREZ9GWIUN4RPRAs52swFzqPAggC/NocxQnz3
wdrY+ODoMj/PJKjmuzOST/9Dbv9d4RMpsEnAPXEN8VVRlhrsjw2GwXoDgBJx5cEm
5+zak7q7kUytv4vx/G6gVQRg2whUoJtQvcSZKhIFrpyKLDztbKEHYYC8a9UW6z7b
2E7XlVQ2NpdSRrWEdMQ5CFuCBT0WgyZkRnmimOhSoMp6b+H1VHr8lmN3MVqJ4JZn
c8O16kw0zIS8fPcMH2FHlUTNuuiNHkcYYmhL8bO/AJecgqTN6esJZhTrrs6oozwf
5oC/Sv+ZfS04SHwYSDZWjo1aBtKDnLfHW58tAaBHFJouev19H+xHBr/yRmRKRyE3
vmVHGOv392KDgwrsd9b+ENE/v4lDljPcdt/UWlcxudjxdiunN9gEETYr6zMVslWr
nLkngNhuhc8n2R2Y2epgc23nkFddwK4meVaYTeDdOy3DY3DTcDmwcDgpXds9Wzna
4yR9anlyAisRR/zcME0+jGbIgMxaTxS/EuA5FlsmADDdS4xJ2ML7c+qOSIZLRI//
DTCcMdgAI0tKukiq7eOVPjkEOQ3fA9AulLpr7ZohZO799xCSnPcmbD9X9rb5uCYI
JDt38M3wXmvaxojeGiI2KIfmJrIRfcjERJcnH0pEtJQ0MEjtHsLpD0xZfeRbKwzg
MXsOz7fzDrekinp1qZrXb1Y8n/6CTNwYvlc31G11WnCvJpn0dnYOQwph2G0FTpqW
Bw/iF6CA0c7kiXOh75gECOFYSmmJ+00e5FySJMDs/Db1Hlmbns66ztLrVUO4fSEG
vGOliGfOuCrxcVX6z/BVyFwUm2BI3EMNIAWSAkVgHYX6+w5m0Q0pck5zW/ZNsBY1
WaY4zPUilLqGDx+RasxrU5I+yYlXYgoWuhAXj98wApkhevEvnlcZy02jRz0f2Yj2
MJUsFls+FID5fmhaGkp6/CyIZun2bsDyGdutfHVVqIpYOVH04zcDdBFNXebRiwzW
5yp7duCjgbUJsXbD7ZNJURoVjdog3z19s85WiJAQhCQgBcDNuCPLA+rJD7MBv/GW
CymFlQHYghGWsmI6BnEUB2IA9dHXN/FcIzV2ddmbD9PtIKU8FfJv82IQuU6voUrn
aZ0cseehca1SSExrsw7x2clk6+iTzEQ05C2cgWsc87IyojYtuiY+coCuuqcdQ7Et
kzGH6QTArtY06hRo2+Np5ygBORPQr1o4caRBxrfTHYVEkdQnmwUidP2Brh8POBLk
TUrZAZSzJ8GwY6SMeX72EZf6p53WWeWxQP0QM0W/GEKYG6sM9S6ZJu7Ysh2hp3qY
qXVxzBp3c8Rg5I+xzH0UG0O0ysA3fQ9bv7tYiBXeHBRFvmDd0eDm98kVmt+i9R7D
HOzrRLDt1E6xNDwAgbelDSa8qIz9pNG/2IJFsXPUYzZHKL1VxU7lxiWyKMwxSZB3
L8aAAzvM8P/sQLEdUQfLOPTqsG2f/2cPovWAxJKNqxc2c0yDCzCY8pMDcGgvdfZY
6RdXTwcYZbwx7UTq6B+on96aSAcvPykhqKT0f130jdNHKsEQtpOWxwH7//vVHSS9
RosykExvFp6UXR5T9PVSgwUp/YPe+nr6aER8z2g1gkYJS+fjpsrrNBRPGcBaihpc
mea8S1EVhgx4jSyozrBD3rRqdnKq/C5LuwtJc6xbALrftcn7bvesm5vn7nLTvY0l
PmqM+a5M7O/bwcOhArXXOcNZricEG0BiCQGelHfb0nKARWNF9s3UwuwnPwDkjweK
tBNJUTDu0o7Wvjmq/ga46SpxbfI25JhhjpUvs2ndJrmINfrm/uEWW9mWx5CGnhHK
uxf1KczVddcyP6x0OeBfI1TNIfv1QkRR/mbZC9gf3AI+Kc1MCTK4I1ixVgQe3hKI
cwF7aeRHIhKXp0yOzbX6KO3e+3mleuANiVxfCAvPs3jg9DIFJnrxhw5xA+BTsysL
cJ2q1E3Smjao+ctXak9Wc9GOxUAJZPnV6u5+dDN1f1IlU/QIX+ioXZTovWkGbmea
bOB0v+Uiibrc/7t4gBVaOGm/CIglxRxV8J5syhDcrWaJlsRMSVz94Gwuk3GaeYND
jgp0RrDfoaozNBLtIsLYVFFddQ/ap/2qELBgyUsYWutaAtwXGKY9Zgk+wAgBRB9Z
IV5QOAvI9ZWloKucILUN751+LLkdr1r0Aqa7dbWgXgCo/nNZuMgbOGehf1D3fmXA
gp53FBPrLXndCPXGO8KkztUGrsv6h2oq0I5o0Cl21vgrf1zBY1ip0QNfCEVSNkAg
iNE8ziSegqacoZutqawG9o6IEV6ORKN57f4BNw+E6dVCusx/wceVHGO5DXXJHyhL
SBstVCCB3QggJgX1gQuo/K+T9zyMQcomyqSfRptMpvTW3rrz6deZTS+qEJDLR8Rf
tXYXhH1zcxTekLnuyB3RKumUYhC+V6HWBGiXrDQAW+rbRYqZCfxmH1tGLo5ZbNPY
Hn6FHfz549PErHMoxRwq/cmMUO8LqHBHzfA8r6Ah4k008XKrYXnv1dFMRI2EO1Kb
BPm7CRw9Akh50hNKs8CPQf77a/H2WX6HBtTzDFIGhyGjLkai7WZTUwvVYREto17g
XmcshaNX6n+A1HX7mlUo/RLmRwTGcgQeeHHGLlW6yuUT4w43KWdF0dXTP/2A36K5
0oaxtfdtRoNTGm+ego7VH02Lctf9J9BbptwZpBCAY09ogDdibKgM9HxdzX4W6Xdu
cOIHvUXRvgXtbZ6A9tAdhgO3odW4XZ+q5XvrIcoIQJobJFwarGDn5KbGnfuGQOvm
6+mGYBvtUg8DDSZPDsLESw/oujrKWsPRSKFd5zSvndAUsJHlle8ltpNG0jc2uqs4
C4R7dW5K+uUewsVqH5pi9ben1s+YEBcox5zqnxs88faVxAsVUs5Zd/kMRYG2QhDk
LwDw22+43NOJTc/QJDkO+Xx518p1HJUvJFOLNzGsW9OGhC33EIzqk98REP4vqot2
mHlRQJ6v44mxUh1d4yLKOaAvzr+tkrf8fmkZO+8nPJae55IZ9RQmr7xfsDS51QVm
1jrXZaAMbgTp8gbilaQYZNee7HF5+v97/YPH9CBpztc0vlw1LxWpiqwWnejExaES
eflpLAXTjlxPQtd4IMCc0OlbrJUvjyiC3WfAXmp3rq7Q0n3yR7h1FXFY4kX7TfFP
U2qv8V5BkurXREA3qyn8EyrdDV4/0YUNQ5eL6FImRK1/AEmFaH3p6N3w5YOT3B4w
Op83h+5SNXqs2pSb+6XGhIPY9o4DA4sRvb2jjaVDlOZVyv/YgDIarcfcFNMaguYQ
K+L3ErLBYrNgMsv/xL7H0EIWvKAA9HnI1PB5Jlj0TTuMAY8BSPjbz457/cbRCYWu
gyqP8oLQN4xiFOMpvSiBJzwTaIQkItQOgnrB3oslq0lWWOqM5U3ZL4GNt4RBOaNR
zNU5M59FqYsSMl+2SKsRj6advHBaeafClRreUc3TTmuASAlV1jRB/Hk9uGdFe8Bu
fSvjexdBp0A8u0YEuHGRvmWy0miVhhLR73nVoqEztJ26BCg6W7zRgXIw1uEfT0Lk
MC69T8ZqnbiMiD5MVt1BpQxRfrYfUhSMsujyu+uW2NAgKuWIuJxULVc3yuk/OhLs
+ftI7EXgoBIis69fcxPlVxuq3vKyyeDOpGxIWgBUYwNNZf70yUMXUHcGpPuGfF7e
C7rSkF6Mz9D3EOSCmsifa6CZE7QwuvEtEVUTVRFtVQ8Fg5OSU3CehFprESoSxE80
lckF3BiMaf1dovdS8slE37xyGxgMZaMgXfPyIs6v9ZG9USo5k6rRfTncTYpkXgft
bNgexeOGfgztjdVJwZGu9lGsa2kgvoTgqCtKG7ifSiI35FPzVJldrX3ajEMQ5lF2
h/U1vSadZwuNURzgIPitDNwUJ0aGvGhxbFn1lTPJLOtEhkbf1byBoYVk+fFKcAwZ
QG4+znKfq6Ya+i6+bp+faWSe3Be3INPgsaE4QIIPWjlRxXcHlg8+W5Z/Udjms1dq
lZvis2SJM/RAq+tIdr7AmvZoWHSwg8KWRcGOHm47OrzI9+cLr3m1q9tJsg2FTchB
w1vlIoRhGtbfkfOrqZui4r8hpNyd7Urnrp/DnM1KLcmOwyD4l8vhfvi7Ipu7CT4/
4ggUJXHXMy206GGndM75+fyruKxUA0Ha0Wex9JiIxv7rm0b3Izqedphmh7qfpeOx
3EP8t+suozxnWBsrbJTpgdimnJuEm2rQFapA5hv0vzXrE+kPaJqmc/qioxw2jFI7
8rxKukmDcZ0COXbbQl91PVw3k6Kd1MVm9MN6DqgMjZyz2RkElJdeEpmA0pMFWWmF
mPAIL41b1wWrXuogT0fqZ1Uhgk+0z5QK9jK9un7NGJzNca5L0AhG5ns//QOCASFW
xmwXIj3z0sxpGQ7T4zm8/tDlOkp3gzSft9hhA3inzzbBaiJD6irE7icMUbtNGJFc
n+p7k2Np+6TQWt9QhNmm3fj5CxiBI1V2RaI3LMD9kXKlfIigZxQzX2kN327cqPtw
0n9azv/O8NnbCMv154jyNVKAWlflI3RMKWo9Nw0v9lT5DgL9l2BNpAI7N7m55mMJ
lHs4mkJv567oJGFsN+GUdnTKq41tH8J4XslXICa3JOdt9PUbW0q73JzBt1lHDU7d
iDabRCKNp+f2Qbs/S2O7u+tM/WvLQKaTxtSCcrcfCo5w6XmxMKBmEHT2llAM2wPr
6uR8CUBKxMIky54se/xViqYEIeMV8IVQdcctv8zUxW1HPxnz38UTkdob1/aqAPeN
oMoLii4YAE+TlSF7JZzXPu7yjGVlAwUcijQ83XcmXWxKMu7+mRexoGEA7mNGLIM6
kAJmjtov/hM+lzLxPJjj2vigAn9vviDbJFCGa5bwVLJZaHvcl0XZwv3R4ehvcrpZ
KFYSXpj92k/WLCaGVg6vKJtrj34/VB3mJV/5OwtICN4B0Z80MBb50rl/dJ1mKtIe
uMiXBUEv9OqMniDBh6cQOOFIR28uHMYe4eE2gFs5RWicZ71GHas3Qxd2KESnPCkT
5iu7wE79zOJ2JTN2pqnFZo4tqyD4SfS+g8xQV6oVU8ERMjN/mV7pOKVzWsp9Jb8w
q1BrsSlyUAG7x/KaBoD33V/Jl5HhyJlldMT2B0AqJZWKRo3hvjmWG1y/xdLecWQB
PVN4tE/AHiZZh05KtFodpdkK3SrEn7luqqgDZzLdOgsowft65j7XGl8NOjlTJf6Y
fFQcnDVmH4Fp9Mgux/oH574PKDdMQF3x+IGcOSdLEEL64QoDvUOm5o132yqXJBxZ
lvg1nkrnsvMamsMlvqKgCJdgUdQ21V5gymrwDBcTpkdD5UZt5+hE1ef5VEMtQEeV
ttmh8DCgt8ul89IK2jEkp2t1j3ATrvgo9LtFHTu5tT7VcuMqTMCEyaRqnB9pPvU+
XULQaGpgy6e7qu6Pa7dg69qut/85wIpbFjcAV3ud1mLpg5vBTUdvaboUdCr1iIol
bwr/+5TrszV0P2ORUgKrfIr2Y1zmeOeRN/W59C01vt8lWuLohbStAo0JVBhhe8x7
AWbo3v/+6qnV9jARgsLFAuNNkYzGto4ptHf01qwH7uhAxmf5ypGt0apC4eASNKLJ
h/TsqV0wUjhO/vhSwjcwIHLhvgpLmPVOjWr0mcJyCytPVHkngzReeq6a5mlmMmsB
XYL2o75mTElody430YbuT98bBTyETXorUX272Mfkmdrneh6RvlBsTjbFBsDPwyHU
8KHyd+L18whmTD9SJnH0PcN90wvcCAVBza4bwvYBH6/EQXvq5Ka6EF3nu/SQb2ha
e/p5FHsQMLwCuMniZ4WQqr8VEExvHRrOP7wxCIA4ZUA5Qvhx/K5AL1bCDjrbU5To
StNbXI+OY7T3WALzOu1dKgTsRgLhOTHk/hvNrAse4YXhbiXfkhzdP5Nb7t8my7Rc
mmSs5d9qBf7A5FaOAipR2CXw/Nw92YgFP3pYsfINJ0fXHRIC2cgik+N0szAgQUJL
5W5YixlAUtd3iX19jYROfNFD3BE9GXxtQT4pDZaviC4HJ7g+IY6tuVOxXHRYRAMT
RjeRtz48MgpUOnrZhnzcv81V5nQiucvwg23Lti5mv4rj9g5g9riwumHVBzBdO0Wr
yY57QjJJ81kiCc5rW4HzZYs4BADDtNlUk5aeABHW3cWXNhGGFf/AdblZMk/zi43O
iH/k/N9iIECdQmYr3FcXoyopEkqG5SjeUKhBYF+unjso4nFphrhCJFIcl+8MI+Pf
FMutQfAo8sEaXBUmAGpcPoWi3xH9ubZylFlUTbUOcBNX5guFb/YSMVJt0jWzFJhc
UTBWF32B0/wY2QPWsge9vVesUpEC8a4ZGSEACGnCUESD2PO42hwGzXWZuIbPSa3o
suF9hvZCH5kw7eJ9Cx2YtfzX1DkkHvFi58b/1c2g5qjxIU3Ksj7WtVeLjes6q7tN
/Iuph+ktwlAbuET03ucHaAWcSGertJuze2REcksYvKAzkVl5xfsusLvpTEfDD3pY
PLry1oW8wJyuEFANk/EjKBiZlsUfdNeflFSGHSLEYn5VVv/jhoSSjTx+Cq2u5kr1
GalowscjyoddfROF9LG4oxtPXG61KMj5jm8p6yvM6cy5I6+aWHZfVuwWloXtw6t6
ge7xen4sZJNpsaGyJDlKb8b1L7gTSsi40J7bZG9GaeBciUV8dl1Gh+Xp8I90aHkF
8bpuH6oZW7Im8p9vAQnwkl1HtlYDixwiz1sVySf7nVid0I8fmUzlR1SSALiCCy+B
y1Ilu124NreilDwvTvK1k8ldFVQuPLWXPT+sfFshGQ27HQW9YWaCArlH7tAMKfow
OPpw5JZZ0Bd54KccpJrnzkHPk6A4mk7DvkvHM32lbKsoXEA2xcKbSdxG49qXk1RE
Si9KryHCtRzsjizGkoKm72raehN5BNEgVGPm0saww93bP84nTCQpkiP8R5dgIToU
rn/Nm4MXPp+PaqPygOBq6ACwGPNfmiiXvIyASrSo1BKT6NEc4L2dAMcvTOgsAyoh
4CvPVzOu9xxTlMHW6dCU5cwZTgj1FDRb4iFYjIR16nzf/VfyawubBR9nS2nTmMpX
zTVQ2fKMJ+83ujAY6suo32xJHv8DKz16HKpoYgJ0uCbCrMtXbg0WWh3JPyrXMOZe
sIkJkplzQgf96NwJG3p3RSnGBW9hjZVdAq9oaDFD1cwX99bduyfQjojWBIWydKjs
/v4g5CUuaMoTaHQ+ZsamX3/g1dyMa6Sshd+d+l6nObJb9tRbZu+LIj41UQtZUYeA
5VyEtS5Ascz8QuIl2GV6yvJv2tNzbYksOvjlmxGvpkWmICZNVrChzoR4srE3dF1Q
h+GvCRodkBAppw4nNmqQWVLgyNYBiVxn5hcdGbq0aFTj13aELlhVqVn6DDEycmRN
zLNsTfSQaeOsdcxOxtWZ8NxR577D07Nry8msbF1KhVPEXBoCZtgj01t3cPY3CIjt
+6kb1daY++Vne1pem1ONns5sZJ4k8ddMF2Tkp7ZNhbf5JtS93FFery+XTrM/XDhO
Ba0JxRzd67D3KyQOTyUIiOqNkPrL3lCrwPjjCaatTxlG/JGMSdrKj+6P56C2/RAl
3KV3w/5j1JqN0vMfBbTofiT/P2GUrEeKEpa+MNxpDjUjnwyPxXKzsrmiqmxU/vOA
rX1IohUTGAL1FgP5dahqw5HkNXo0yDUUZpnEzphgEmOYvlGj30rN2FLri1H30ZBu
Uew4R1ccij3HdktQoYXUsBN7o8qVP2ak2TaCBu7kH6RPVUtg1RVRBlJDYCg/BtxK
xtBroxtccwT8B6U27B9SKwTkXSU9tAfNVQ34K+9hGM19KZbVivl49XLXtN2/UNAU
4q0RDIpgAQfRySkIbZrz2nknQdPpLl9jSSutAFXgLIC+X5KKTU6SIcC8pQwj090S
PPj1XOXETLXy+1jAZik7oFb+YMMcG/mJIzbQfSUGi7736UDys2AbcmO95ldpTt/+
KgcS2/UTuCQTvTW5i2tl+UtVfdtaZnyW7bMiQaXIleuTNt0UVJvkmElDYUOrYoIN
pAMCz69xPuYtGhjMXtW+6RBHEcGsa3FLet9Lf+7oL1PYs6NkWj1/mzmQE4c/pErd
sSmC0r7giobUh3TAfHCvQ5nuAm3IAuwSt7/n/GSJswGwQEv62LDpyi2LWpTsEcag
LQ9YhhhLXcbeCHsovYxBhJFyiaKW5WQ/Nmo8JYLiiOEe34/BDKJrzkc2xbM1KmJ1
QhyrdxZaLy/1HpmjWwIxEAFrKSMyQVeiki8rW8Qeekv1+NLnQE45sIRkTtbaoiRd
4P6LyzUCLHkPgkzjQDdwU/Z4QFaS4C/dp9R0NoO8wMHE/8/DbF2x1/PBhSxEvvZ7
4gyJJtUkoREEpszlKqL8m8MmVrEFOVs+Y92LvsUSR3B5VoEL6KLj/qEgGX/Jy26o
x+lx1LHZCD6TXdYnvdg76roT8o78yvbEp0HbpgriVA6yYUyLqOgkwLetNpch+x1d
5rBcOOMZ0mzBv5ybqEYfv1VO/rZn7/d+JwfAQ6JvwznWGZx2SJ06w6mjU8R1/bOb
F0sXkd9RN+wSxbOLtO0CBiihg794Vfh2AckE+5Tq6au+ZHaDFa5AqLAb0l7BH36q
Mu7xuS9kOr3RxTMwOeHs/7edcN21bI9Lncqe2Kc+RyK2CcCRgdWDWivZU/yr9arI
WxPJ1xv7HZpXGDvJ1HeLOYs14cC7Ik22KyRBg+dNzXUOODd6g+DLLbhCN+Yjkn7j
nSQjgWGxsxkndRuXE4oyLNxvhWc9DNtdP+uJrLo4G496o1G53EhZSd1BE+vDGKwS
EvhelLKMrLXn51N0/F2jH9Bl0OQ3AG81/gUThEeDLGIPfmmacOaGDUpzHmeNr2qB
jguZBoymbxzlVenyZUdWdArxv6ZF2QDqZnuCOeixEY61g+dzQtH+K4RE03Luimny
1MH4LhIfLagmHq5Ff0pMIn+xEZrH/uYHe5In7Ci/16rnH+wflViUOz0hs79bOAzz
ZHPs7BnYJk29cgbK2uYIwJphAnQ+3/b9OEHzvr0aG4qFarHjq3dI0xbN0OT3Ax3H
KAWzE1+DXhw4zkx8OfJr3ciaHP6jfjkHkYBXaTDDFl2EK7bkut1xdDbP8rW+G9l/
uoPNh08XJkVDECJ+37SusHHOnH6TQzKdPxZhYxqYekjEkTiZgqAKNnmM2dYxJhP2
g+f0c2RbG6FMl7Nq9lZ3OQ2t/Hga3FfR2RVANQZuHLDeVaS3Y/Cp++0XanSZlIGD
Vym35k4dKEOsofCTeLS+hYwtTHAGSmI9g/N1Jno8JAFhIHoSnimmnqv6cgKGSdyn
gPmTE3xabHtaePrQ5FWmVCCWLj2eR4Gtcgqh+1eKXNGTQok5T6vJwL2wbJpjXUB+
OQCGKcUtnPe3iwCJ3DzfoIqyLaCR2yCq/Lw9cFWhUBiMhXA91Fe50PFLeHMcaRSm
OS6CQbbHQUCCv2OzzyY+p7BIplqswUEkKRkkJSVnOokeIGtlfmSX7Mzo07jrC4ZX
7aj1rzUc0dMDVuajcOaCz4t70bi484lhuF3zEwZjzvYHtRS55Ljp3wpkABxt0Kpb
sQYji4enYNBumKtOycvrGlinxUuV/3OPVU+cCMlLWzUk+uMrpbcowSy58XNbs+AW
pur5uVAcshLAUepVQe9o8MGzCW0OavFwfyh9NBqJiqTjnsfTTQum5qu/S2iK2tUh
Ey1F4YorPU2JzjRedX87s/Smpd/wQ44qXcxqno9Ko/Q3DaS/tT4Yf5d9ClCfsKSx
85SZRVX7fcHZhsJVtGbRPismQ8qLl9D41eqnQOnd9G0hv7rYXPM7vpjC24LLIvE/
9JbebSgdxSgREbkgf4zJq1IJDySz2w5T6B1WiOtEEmK1SUGpIpSTcJTLOl12wJXt
eIHqULlPuUY6C9gra6BM88oeRPc2hL0+Vp1aMpjs/nG3oju21K2pGCRS2VNTCcYR
YZdXQKy3bHUyz1bJx4NsCY11k4dbkg92r6NF9ZEYvOCkIgWt6tF5abjLDEzdB+vs
ZQzIdMlpG1WE1oRoQvUk1THe4YM+AXxqGQ+Z243GWieaBr4UEP702VTgmc6K8TZ9
0E21eL73pNLu4t3OQ5hn/Xrj87Y7DEP4/GwiiFnVAYaLMbK4YIeoKefYnqCUDm/P
SBMADxOeEfFOf+WmwD3HXG9EnTX8dGsL5qj9GiuGf2QYphgrBWLyNvRlFwR875pJ
tyhQl5gqCzwHJ4dG+4tJS9gHEE8rcvTlwlHdLbX6ZqT0uefw6fDRhl6dk/9dRrjC
AgWZu4p2DuDmJLJENLsn+b1u42DoHkGIEhQ5ZaH8/Vp8cVUDdg161HN0QnmEozRy
oIJakyK2aXVlgYUGwuCfmQCjHxxmIDSS8hWKpV3Fs+GAfhHOWYMpGdt/W6RaO4rQ
+YUagZjuDBxFp+OPQw1sJLLTqg2oeWM8wgKNyE7QffJQkeyHWWO/VpqSz+bRduE0
9VowAYd8QLgNc+o52zR3/zbpjPEKt79Xe4YjelG4FLB5EI+5KVKh222YNM1tK2g8
hD/YvxrRxr7jAs9WA6M9TJ2jEyDp423GfDWS2qQb2+4feS3cVa2VeZjVl7Pnp9Pc
sUpASG80gW+RrRMw3xU3dTVOOZw1YnPdkBf0p6C+S4JmQI43ifH3PdfkaJB0EiDO
g5LYb75l7y91aG2rHQrQKbDYF6dnjYjK34+HF3w9t3J3OhmevXo/zMndIYefYXJ5
kvvQx4OxIaQ6NCoBZ5EUW837sGzMGlt2lBz91TnFM9dJ80W9FGY2NcwEKUYe+MWR
uc2YzTqnNMQI4U9bdEP6SiSMWwNhz/HwsMPipc7MsOvWIihPS2HY/bCIhaUJC0Cx
HMPvyeGd6owBaoHXrQsb6+98eD76whAaC6UkppFqK1z9IY/1yv963EpDCjlszkVD
LEhY50LLeJkvlel8V5cOjcHIc9f4oeyUWjW4bp9lnTzkwuJayd8LWPvN16WMHsIX
rcQBctsiWIR75WToPegfQE/ODhHtS3VTp+n+G3DMQnDb/VoZFtPWh/xG9a98BxL9
kujCWo0pt1T8xXGodWmeGbRXhGBrzparuEEqn6BhxnvxqjaIw6cFt4WxLsOIA2xq
uMCUaFPHzr8vyJtG+398uh3meLr1f5eUrQADIrF1mVeGCMHDJilfY66ZTL7M74uW
TJmhAWXUMA3fxNkAylhiIYIm3M7YuXxyFo0L6uxJkKg63ThR42Ah98+jzh/55QdH
SFv+9EqaShehbQHVhmVx4j4f6l6cifpiXlax1j3I1qCFIUGbl5SVR5mUAV4pn9TE
JDmGm13f1fnhJ2dK84EiN2Tdl+Aa0ewgaehQVYg0iWEXXsvvQocrkIH41gu5jTzY
JckfqQl1UWh7LQG5QQMns1d61BswqotX/jwV75tMF/85iF39yoGjhYJxG0c9pM/G
NhmmMv8I1K6fUq4jPYlTqSDK9jEpqP96rLzGw78b9JtdvatTMbh44n9oj8oJYNah
RTDPzeeaDo7pAshcM6QTk5sMMKLWOeCRwJYT1emcYXx6yz381GJR0aoBenj8H86B
AAku1RioOu8Vd/NZL/35tEKyUbz8YKSSDYqtwlJb3/KEGrdA1yI/Knel1XxTbCD3
C/ECdncFqLwTJ6qmXPPS92D/v1sF/Aqd0gyEYVgq9tASOXC3fM2nhr3utQKuP8t8
1CrzobuzjH73sNfB5UesHUoHOvAKoucd4m9ZywwnZfTbPnjK7fJCMgqtloDenT2j
h9/yyzfVsWdMoy7dWLt1buBIEb+Bt3cSKHS6iwvfxQAjFRt7SOmSbS+lm80O7Ssn
0jjPqLOFAu9sxtiHeM1SFHYE2XhLwWLDvqAnEJW7XaghOAt12YNuWLGk/tIBqX6D
X9X134LOxxjVHjLiXLaR1IUz1pyyj7xTgJdt+RCyehahIqB0p4D5QlujwLNB9ORB
wM9pKu2qMP4Ij3srHeA5LxgdPdungvNuI+4bykuritT4j2xBiew2lgSxQ6V/ML4L
jMLvmnEVAmw5QtaUAHs2IqrWFkmWxD1M9z00sAFKqIzik2aIuN2BtF7nIusOihxd
iBmZ/2AYKxTbmmXwFHrVPrcBnsPAF0E03hq9gtnAccVrvYmAHA2wdg1U9UKNYHwz
x2d8+fOQB5KqXVwfmDvZkEh5twlTGlQIwMjjIR2E6C1xR65RchkOWfJ2iMxQV7o9
zrcWlMlEd8NHxhbJuyofjoBKfuNCKGBwagbsM0Bnih21clnFhD3ssNLQWGeAxPko
HyLo32P+MO525zFQHk+8NgYiHrOqkV8zifo2J4ToAT2AsvlFctrqsNXfWtk3lN5p
fafaknG9Jjjyx/DgTaRYWWa0qsktrc5Y9fqdxLYZioZL+cBnUanZr3ToEcLDjR1g
LRiJ+F19rysLvThSiOxvtmuS7xCi9p/TYVTsArMptZ9Hpz/UjJ9ucQM7fxnDkUV2
V4u1bTZItxB9amlu0jKMGhvH/wlFAHqrXy5V+IN5sI+fRlHYl5/mhrsv3pOvVVVj
IYBwiiu61dzNzYtHlqRzHb+qTTi5Wvr7waK1CNaJbAHlD9H6yLJ3NgSstFufFY8b
mvCWOJ7jVL4Uro+IY4Qvwzu25mj1VgBgUY2b928WeyrhJ/+KRSXBeYMCprviUCk+
q97ZiLN/iRGIXrR4y5f2xQydqS+aDioZaHJ4FOEiX1NfEO6HiZJKE2w7sY+FSOkR
irAZjrbM7NVH/9RQbl1LSgBxJhp7wJcse9mlD7bI2cOMC8gwzE13Vdd35CfHf96c
MjMemlpfcibAhQESKcj4PLfdUR/gsXjZab1pFC4yqkkdv8fumEfnSZilDu+LcMlT
y90muLbtbShJ46jTXkPpwxYmWyHEhIMFDZRvPKPptfq+z+n7hfyF1HsS3cnKUELM
7fRRIv/8EjFfWDK1S9lGxSlIZ8BHEFlVt/NbxOHHOrz7gOdW4bAsqpbf03MpbE1H
OQOaDJ5dJhYSVAX/2wpO1njuyzoBoAPtUjTJGQZ67MtQtEz2uS8X9lmVTlxq8+AZ
NSK7bVCZ59chf4yWTkx0SiQ9tahXabHQSKZPm1uVxInNRIBWtUL4A5ve4z3HTzpJ
zZq3B8zKqEnGKyNgYTCNeJBx6EAjkTE8DCLJlOxouP6QjBf4X9eYIVQmJyOZxDbm
mRiRf4UD9ixy7TTsBrV0RGoxkfcNP945PSWwsJ0SqUuub0PHLQ2HnRauOyCU/sda
i2RjijoErFZ2c+F/e70dflkmdSa8iICwFZc6SoVxQsCMGut2JdLl4XZk0kLgYa93
fwVYH/3yMPQbR+k32OQnClF2g5x+9/oC8/cn99MNGXffpeW7ssh9MFB4C3NhA/0z
LWq7m5J4jyOHv85oqjPQeIEtJbKa7qJo6dVHhUYGLIfXnC41vP8GTmqQUgLtx8dy
F17fiOvCL+BeTtbRWDgAXoupdja3c3o8D3XAxMV9Hx2oZRIDsfTJklpK7GEQfWO9
4txD31Lpf2jt03yLiCUwfd9QHHgw47gCIJROP6zxgrILRx8+pTdgIzDbEhomS025
tvbtXZuoECiPbNNNNRyGdjj5scGNNVGIidJJD+wzGsSffuI6BQEBnXzPRefsK67T
F4w7JYguiea+KnBEGSek5voUKw21pLkIxZjSW9F+pH4g2ll+CkAmAQUwvJIhxpAR
I67H38uVuKw9VinuyBKT287V9PjCYYAnsjT7SZhvz2477/Y9a2FGQ3gRmaan4ZSN
rCq3DBCMFfUmrK3Ydcjod+qQINEOhBR9fgGt2AEBeyXlFMZzmX9CSyjqFbPQfoh5
F5NAoOFQq9G7ARCBcwL2Tyo4gLZwlInoPgYOHV0L6RKIGbORAEQBNWre0kt3ibc0
vrX+HahTZuss3+KT64gppeNcVexfgpnMpOt88pg/UJLBnCod0xdGuOHtUZq6L2Yr
/rXlE8PbM+hrKpPAGAoEO+r/d1Rh2e+sZEFyc2F77xFn7DTOyrU7NjcsIo+j2zIb
xGq6YyBvf5WhqTBSOCEreGG2JUd8Fj4By8MgEd0ASUolppoIzzPojQVmvWUywlzb
GJ8/9+wuWOtYS+oKnEDTkdVWsZFm/rhLtIBLGfzjdxTjnVF62jwPtZ3QzplEp8yg
SFnkhOiPPBiWbv6TGUgNOYP9kZbqJwkb0LBlCvYG2F8NYlsc8tVM6bxnP/ag4cbV
VKDsa/YOUIt7cI7JbbpNJ9JgHQVXQBQUC4lOd+fExP8n4GYmmLgNrwOx3TznLgv3
s09VXYShrTAjVJ0IXBegSIUAoYUaaomoaEOiS5w9l+4AGn87aooA3jMFY7k5ySiz
C9O4U0wQXCPethDXPXwLhbct7XrGPAefeVFm5v84OIN8WJbH3UI50KIER4UGlHPy
bJKDixPj/bPIFq0cdPtu0BAi8vEv/OALBIxeIEh0pQwRL8f19A6pzSVD7thLWedu
yY8bNDW84utAmKUnz02RncKc239/kPBOmXpdBP+xd7+ZVaBCRpHVJBnTeVkjMADW
KWaQ6034xQQeD9u/OEw1ZYwJ3VZyiPFdzkTAA7sqS8IwXCujSKv7o2dfMR7P/rER
nQ9dgkTp0A3QtJ5+2Y/R0M6M/jBRtxvqDq3Hcms2POxiDF2ZoUAE6wnDOxel2yRv
mdCZPc3lneZ3sBTg8UlIt1Pa75/Xaupx3DTcnbwOt0EO0iHiBqElBJozaN+Fjt+g
xf1DdmfZcwFhi1knBJxZ6LGCre+v1QQhYvvzrDGFaFAEIWzVTD2inUyw+QcF2gMA
QgdUPWYnaC6m9kwuWl6rX093Pkl5HnTz70oZ2lleUMFGV2vj8y26GgCrh2FCcCzQ
8b+x6qjQYlI1FosepeHoyLvj94XGg4CttPSdzyc+ixjT8R2oABE1ww+Vikhp9pUS
quzw9xBwGKbrNqucrvyWj+TYzlP2Qa2lbMwtvveEXc+/KlFZ5eLiz28E02uRBorj
XFaHgu4fbrgLhy4e2DJipJPokIM0vGMvhFPieLXvPUiNTq4vH1hk4/9PzsEYUipU
brDyf6+4B81/ZL/b4wA5unDTl4zh7wpLdcVBSxvNVHxvjn6Xw3gWKCUjpi5MeM2s
8icKW9JSeMSbXzNrKUnaITuvpoSTE49zqp8xDGcOKr+uZpsH0qONexrDY5CGHbau
AMV1mg0IQaTEylObSrmiwh/N8F/PAPp43ZbIKxqNpnX6Vpbb4vs+YQEpbITZjLM4
DREaxZIlUyPeZEmGsOivhzKf+TppytSftK6m/wsIYYT0FkwqZnyvlsmdl+MQBU0i
DSUHErPj61FLglfwD6pU9f4Mcdj2gnrhbrmchS79I5E7ZcFEbZLfN/e4QVdJ9gil
st7GLNaTGSAAxfXqNad3bIfnUxdJqvqpyyt260Zp46hlaed3x0xLsuTNSMyFaKB6
mOJnNlrcCahCAdWSN2LlSZ+6gnAH0pIlI+DkZvtfKGntABIKRicXOaeaG+qqozIe
Z4YqheCnfDdBq7qBwjaLvIexDMe8QFczfXw6SKI2zF4C/nuL9FAzHjoLMvHCmC8L
YP0/AbVi0EYEJFToA5hFlmy1x4XFdyxCb1tvizCP6XkiFdqffXtn0NzSBL1C3eM/
neG5lSyyae25aRImr7or/eAaV1P8Tf59QMq2eudZd9SD+D72CzTKn7AXMYh6x7XB
vyatHRodZ9atXPDYWJICdHXEEJ7JlmgUNU8wMTZHp+jywu6d2vqn030oPBEWIXy4
wJexGcWHTQ4dhiviCQ+G8o8ohhMxSNC8cfW15PBMQ2PFxeWfGU+2KpvL+aXeI81q
zyuLkeGWw96Hw8+CcmM2XxChujmG7Mg+GyheeDmNvo+x3atZT+noeG7P3Fu8l7Oa
Igm6wyvBCA2q/9ncrMHk/cpoS30MdzMOrRNcsPE2P9s8gIwCpm9HWbEX3v5FLOx8
bIhDgzE8De3yjx3FUYPKdx4EqEzppzxEYax6BFA1nVQKkRAMUpGSPojtmaJHROZd
2tJj0jcHm0cFuRIYzmZZkA3E8mtXOphaI+9MtG/ssNCVAznxD0U4nBNu8CQgD2GQ
T/GR9WqytqBWMZvOlM6qGSXtL8tN6DasexYTD9wZtccUaSx/jOSzmaPBLlaI2tw/
EmE51nt17Em74FWtResrlo8OBNgmdKcXaetUXyqeDWKbMu3xAulV1oMp2wWolxRe
TF5ocHGVqhBcni69cC//8SoJ6WgXRujloA9e/khbyWj42qCs/0x2aQA9tl3rJ6Tv
5/6VJdGTBQHZu44nc1gxbCxaLSRHsZ0nSt8rHcFPKm3RNMb4gnogfJttbmElYQYk
WLhnZAy9NyilYQGkUV9EzRtxPAe1rsdPbVHKsHC5gmfvyZAtFBibwVHKZN4wgpRO
gB5eeoLtLFGXdlAIPLeDkboMDRzggtwdHihV7+NfYNPWt3jGHEkojzlnvE2onh3V
2e1jLwZGyN8FKs9RLhn9m0vFeYThD+IMmZUJNLBlBY2P4VHXjMVzGgI3I/Y9Dm8a
hxv8XxBHboB6k/jjl25RcqGu0HzbzvXcZye8eyxtmkLQW/99eThBYLsvxV3KtC9C
uDpeBbBet0ngToN/WzQExroBPl8zri8zPU4twJG3r8Lt0pY4jE9yxgSZ2FqCHqen
xcXYMHQPaCLQ87ChpFaWD6iAXBdPVzwmVrIURojvI+GeA1jvtvQPwqPx5g6MgXE/
GY46es4eO/Kkr2gAfWy1qq2g7mNhBrEzq2K6BQ7macCrM1ACb+tJYQamqH/M1zk5
ib7r4AvRjOrSmjTqhWvzgCrSkuJ4A6mWdXltN1DbOJB9h+mmZIKVaeJA1WsztVd6
UCr1gtL7MWfi3phZ8RIghrCOnKjN40rjf6hzW15/jUKa7K1wNTykxCGQ8N1Dl9Sd
j6ptZ2WKcP2zjFQbCB9yWzzQrcjew03vJIpmv9KSDiR6gy0Mij4U2//H1/MrmPjl
S/IWiN7S90WnNT5vnmIBjLEzZ0MS2EODpUsw7DopYRtZ2hs4AXAWFylJ91LHMbSD
4DJVYR9VkRPunZB4ucbWe1/254WKOcZKBl1Ny3RdnpwAGpqLGgMzkMUNpGKbLx4q
qDXdLunMqkJIYMLxmILKMXhuJRgkH288UawX5PFPeIWlZkxyiXu92W5BSEU9UWXy
6ZeYE0L0an46IiFVQRqITWQR39Ir0UYSq9R5ExrP8W0PWmp9cdagrbMsHWmnDx03
87TYYBXzmWUoNR/7g79rkjFknJARc+RVIyGpK9tXKpL4Rkg2zk1eBU4RaavcGB6R
qA+YMZ/59jtcUu2/SiKD1P46bhV5vQ3vnC1kEfK6HIfYVhO1H85YLLn1sZlpdBHc
5ztLODxFDS5Vnu0swhjciQ9tGirzfEknMbN+xiThZDMKjQ4u6I4r8Z5IN3bATpog
bbtxn52MLBnk+jt8cc+SOrMt6zcdaoarUb7VsdRz2DEOFyzI4l4Km1AGvWWE+Wb3
Ub1XsbiNeQd3ZLTt6j4hCxsp5CWyf2YUntAuYYRLISQcjyqLSecQW2pSEit933jB
AQwR3ZKowPY210T/Az0aDAVwIiKjgYfDJn29Bwx2Z9L6N/59vz4dw7ZdlnauTl7q
S89vMG3+7ErmucY15+z+p6IiImUAtTN16mTX/u1A1svL9vIJaXLJJeJbdlLW+vaK
061ELd/zoYiC5TxiNsZt7/gzu3RcJ1CHMQsHrYyuNaNuYzCOuqLPAsk8lMDL56g6
B4j9JT/icIYQCpesF4JJZxdh06ua8pENoHmjObKbLLOcxdb3nSPpoXU/OZrT9FJb
SQd0KfzEAx+hDu5dbPyAJw8mBDOGfY7+0umkHyR4vi3kwtX3xzcgaNbXbojLSbDN
a9Eh6REIAF/7K1+FsCRaGAuYgsDiR145XeiCz/YKYe79pkTgsQikWRppHpMejl8g
iGsS4mx7+Cngz7uSNZtcOOb3SbA0xMB/EAb7JEKeohU9YLdu+VCd50FIDvUSlDBE
AijQgKOGsepwig7iyD/UIf54vBS9pfHQfrCzl7os0w61to27GD8Qeb1NY8eU8ElG
5+XmgRO475TVoDp8VNSjuCJTj9tJ1TWvul1s1ppBvpkzo4yaMm07uvK28nXJcaQp
dt/UjPx0U748xR0eUj0seTsNc6ISQ/uWQ4/D0nL9RtoAxvM4SNDhhahU0XuBn47K
BRN526+vUDvpMVGK8n9ImQ5nb7AL3j+6XPyVUvwqxHHHdePbg6kFu81UtVIZQa8w
QuREoDjmAI92AuAyYygo963NxtqOZeFDQzGNtxt4MG8+yGrPsJrTjASJ42imeo9m
RgmVOXC/7bPKcqgs2F5fIBRW2kXybZZiXR2tN6fyrQwv4UGb7wyru2vOhmxs1N+n
kg0CHFgoEuHFIqtBSN1MsZzKJ583AIVFXZDCb5cRBsSPlRhwWfv+UT1PQZZWF1jO
+PsAR4JOAh+Tjo2utAH979uROQnSrgJAbMMEP8IBu3hEfAlJmsKvsmx8tnC+gs1x
EziWEkeqREQV+70MFFpi7oR2+roJI4digPNxICqTlWJvA+8Vkp6+iIrBhK6e6vdt
DG9QAKlOL+zW3e4eigX8xTxiWorUFEBKLoOJTc73zJgzQuqXYPWVziaxlq/JD6vh
6re1Gak4jP5PQkf9oJZmqOfQbuSoeNeSQua/md6afCIhGeJDUDGVRlaKuXz0iJ6J
0vZSUg0DXed5dPB9LkjENCxUfNoow8tiIIq9+azLBjNDkFenFxxSgEncnp1CJRo2
59dHgAsDHuMCiCEC1gd9GP234N+gLqgWACz2bBB1lgocdz5gKI+qjiQwhGVRDrMw
EtLTYmzwhSKXDo4UgfIE0Zdn9wLlijv2j+0cY+6kpnLBcRhFsW2cokliWNnFAW/Z
Mr/VqpTIGlE6ZjUACIlkSIrMWrRQaFC8/cPX3fTPbmf5lhz6gH6BoEwdAxLXJCs0
GwHuaHRG2V97VyqRF0rfmX62zaBsioNpyuf6HJJihtbBbOGYq7duzEjKJxJVVFm4
jAL2/V7Yc1W0XNLWUtE6EwY3M9hM6pZ4P1C79LQ5lebLlNiiC67g9huZ3/MRf7aw
Sk4LRrgXLlyNl3EtzIZu/LybmJ/64wKZeWsyB11onRt1h25hOYU21C3BZfuC5iLZ
K4OJSr2Vzr2NQpY+nYCBRxwPT1eKZ3K6Kt90Vg/sar6rZ3REk33qx4pGEwbdUpgt
/e4RMAA8NIv/SJ6GTIuvdeJluy+tXE7PD4oGib9qRspTH9fkiJN4vrM8XvQNT+Ok
KrRw5lJO+mRITNit68hi/rUd+XchJDW0A1LlNO4RJMXXaDiLfGeoo9eRp2qprZ+O
mzHu4sc1Wd8Qj5bvA6v/HwcP98Ql775YnnqEnMY4/Dy9LBk4vjSkxVbliavodMMg
Jww7q7e8ky5gMjsRsf7fJBFy8DNDPP41Kyf+SGPDjTQbr6/oI69zf/RwqhYRRH98
FlBNKF+XTbs13qkvfbXoHl5coov8G0osBsiKXlUUbsottC8T2S5UWEf6VVwB0FeI
4iqFEE33R5r4MyHM5Bk2jSgcXqRzoAh4H0Q0kYP6jHka1C4LdEQ8NEsFmVsfvvhn
EQOSK4XsKAzvBbUB9P8rImj9T2DjlmSI1I8ge8uczYcqx4tsKptlkSK99XZV355p
33n94A4ra6efgauA7FFnepf158sXusZj6ngtgkYl8vnQtAv5x1nIvQG8p0neiY1g
Gg9pUU+zm/XMZKABvVVK+C/fJ1DnWmyjuV9MqZmfW7E/9SqHiAJFJCtwBAHBU5jT
jR1tImkl3BSGJVNVpE8X5f1GcgJiZ2ierf8kRC7CGmeXKZwwRAZ88Iu9STeY483A
LW3qu0fCrORMWf8cYKpfxp3kcZGLXdcB2uXz7rWOGB+Mr5y09YEUM+48niHZOPXl
wmCVoiu0hOfpU2iT+y+HmS08tvI7qxVnkdbiCS2LyJM3EtVJLqsoo41chmtkta52
P3A6+8yb2YYZYvxvvzqEIiEkR9YDFAw9J+EblceP0XqfKLqqKstfNV7/16gq+GW1
WLQMa0q9eIk6FkqjQs9NHTn7089+stkYLoDEYsiceNTfCtJP8H4SQ1z29wpvw/v+
1mdEjL9t5tdrUXaT/vw0ZselgGDc0pAMF/R8WEOmLb/1RUwSekWaf34aFmOG7EF6
YC99ODIiDJENhfpkL1oroRirhK/TaTgpUUmSd1W6D4zMNpXrHqUSSsGhKTqmF/Ut
+7Q2+uTY/KNjlDQ7BI5F4/R68/BZiW097aq2QcmJQBBaJ9qCil6MwpODcJBYpoct
NrHcfTRQtfrX4FupBsx018hn1VombiYXo+RcgBSFVYqDUkvrwRSPELEK1QDZypZw
3UQ/bt6Oqge4VpdZ1vEEBVHPg59NKMN0oZ0HEezFGe/B8KD7WLrNE85+aVVkYZZC
n9ackp0t4fwijCRwy3HgUgrtuWn5AvDzPrGMS/nrWV/hh1VV02WwvLZvSC3PGde5
IJsndRP2bPX0gQVZHUIoSTqBxRVTkQovmJbCzuahSn0kmH021z+VPB3vaxl/ERlc
WSppsDJD3jvUG7ZSZybtAyuM1Br7e5uqEZWgegUQLhIaxW+rJ0BMuXQV7ylwyxXv
jJ4IEGiE2xwKWlqOT7uCdVYHvipemNX24Fd5TJ5nE8l83dqd+mMawlETCfLC0Hrz
pQcubsab3yTY+T61K+y8GqzYW43Fm5Bgg2Wnh9dr13A25jgkCIZa27/tfgHQ7ox3
dEOL0hcg3CvSZfPsfNjPtaUtuRaY0t0JmC4pcpxvAmF/wRuvFPGPOiNm/LdCnJVn
cu43XXuEYnJx4T5+ZIIpN89zagPgt2bsWiEAk0Rho8Oy+uDJPK1fQYR3NqTLYG5W
36sXc+IA5S52cAnv9VaXvsewn85wxROcWUhOKeiTufFyZxd4W40Dk3X+bZOTWIIy
LPEHspU1Oj8/TRk2uzz4v9XvyzyPaIEErhDL0APnRfaA/zPJCuJQ67l2kevvphFn
oNkIBeeu8RTzFWShe+2oT8teFYYqyVQX2o+Gtl81zqQFVl8/7N1varOVx/JQev72
8fXmRURWqyQkNQNfK1fPNXMVcecGgiHSj/HrcQBnIp+LU1QEyDCfqPcSUJJxwwCL
jYO4fa5pxsWmKTIRdoVmbESCGiXbITf++I3jgSTADH0RHsaNRyvjyLJf+RC1fwbI
lI9Ykp/XCK0WJxJMhFr+o37KUFaZ76ptYLtXVVRzxidP/4sVO0QAxbpTJipqEdtj
BTH3GtTzqTqNa9hHydpub6J/qfgPFB0IZ1L7DbEesR2ZhYK+wHX5MXma53ouT4GO
aI5sBmkqlFvWjhuq/RXWzHPJOnR4Ee8WWWfnUV5grqOycstWu42TW2GI/5G0J1Rq
UXvFYdA5Qv8iFg4ITrJAXIF/BkxZf/v/p+OAjHHqNIflu65/gcm5RC+itMkvPcX5
Z9WwrtWSYCmaiu1gLoJl6ycF0zP5dqqOL7jyO65jf7bQrVVSpGIlpyuRM0ng9lko
MSTVDYCSn729Jx5K9P5d3SYkgFzcZ95rhmszyVykqGP1irJKesKW2MyCgxAEGIGb
qK1fpj1nprUfwil/miW29iNRTa+QPcpbeYjvXJUnvBcEYZDrYseQWbJrHBOaS+up
kJl3/OeHYXxDdsASE9R5d6Ys3CYfTxbInMD0d7v4FLe8XcvUm4g7p/XhhopfgWtP
VuWD1xsJJuS26RkXGPU+oIU2OCeXnsMNSlXIEXmIydCvFSP6hmg+EVPZFmN1tU/O
hAd85gN+Y28fDP1LrX+DCLoUEW1pNKzMPrWkrF+611tOv2reuLqtabjCMWyJgmJO
BuMA8305sZuC8UQdBlp2gDA3Cos9Vkx65F8/W822SKYHgBX9x/QmJJ+R0ZRQ8C3Y
5T73ps+XIMCQOAhWF/XHBK6PyZ9lBMtHGORPnQJJ2TQ3BahPQWfp8ag88dRdaWdG
6NjZEd0ZEZM6mUmdk5UmovEpwxy+giewcWzNH+4aMV6wwfEW4xyvaL8DWB5mfW7J
/PNHk8RXPxe/AvGBN7jKKdtIDAsfceW8xBWYFFByClpDTSo44I25gDIImgdDrtDx
38s4cviCMvZ7Is7ozNAbII8z8dW5W0qVmsrVlmGIRpqm7zAOBepc1Whr5xfzi5jZ
n5u3NRXDV+cyCBNOr7vbH4DWKDRZ/7dxQfjaZo5zQ1fb79A4j7eMC52mxLKgQ4EG
OPCOOeJR9Ki8ZlXg9lJ8ocK3x7Lbhnqqx9YZyq8A2Nx18sgWGt5D+gkXXEHfcYVI
F7hTLhCkb3krVHEGfxPurq+3hgt1cU682JFgiXEjOl6G51gmhpssC6IvvjHrVGFV
vCSWg9N5OI0IEQQifXYqXF/Slf4grWG/Kk0xZQ1owNfkeW58R2UHP4hWC8hkH+/O
vTCubmp95XzUAPo7TWDglNZFxcXJ+nVlybUklN3YWryhr2R9wLiBDdEgIbtMKZ/p
rubxYNczSyXesEyt2mPHGHrvdGlkv9z6fUzz656tK5PdGIJFXC5zY9BfkfHES8rL
18EkSd6fEMjK6sVMbNNm7XQfV7UH8yaxSvTE5uWOEVHgl7qgXAfhnpsuIceL5Zbb
0RYOX1Xqpz5eaD7q+fENWQQf5bytIzg02F0IfYhbYw6+Nd8qkbmKjbURXqpnMDQn
Yih6Lf0/eycAy0GO4W7ASt1Vl0n/y6IhUHFofLMDIB7q707ro6wmwraiiAvpyE4W
739/4/y4rzijOtJNIf2QvLVZAI2BFMw9iciEETrPUltOdF8xyXlRhYiUg0oxoKsR
uoxQUIapNjNBRnVTsvvavh9JEDNizCaB+/uDNfUIPsoL/QK/BdMlx+ui1h+ZqCww
nRdw9BlZJFbL+6iG5eaYAFpU4SThDFD58yEOgQ72pWqD7mkSCnh44g7cM6TQMG5Y
6awJKoLW0bzr5zOy39/oPaILdCuKIt+QDT8NmonvobQ/acRxulVQ4g3dE/D4lvND
IyRXFVTBfw8UEHs4LjT9NmsBUKHzjLvkC8FHYV7lhLrrOXurt6mGijBQnlZlqZX6
ulKJggr548IGuxB3fVbOypIyJv6BFyIByo/E6kVrq5qTNnMzNp3tomCYM1LtyGLz
QoePUh5qVOm3OfWCXsupWyKfBnSrosJg9HPKSIDeI1tEp8Vxhlg2HLdc0CMUg3dS
YKBbO4Bs9PKkH9Bj+vj3nKm7y4dUazRHCwOvG7n4LKYz8XdRuxSEs97EGDSk4O5a
a2T+pTyj2oqpK5t4+uXlQNugeK2OG7NWWpC1BXfhJck5RzqY3zH1R88e+t9m7BIs
oPJVqO6ganMUf0B8jdtlFuvFrL/5ByA+e1CHzk7hOP0CzDyMM5Vup96s2alf3BKA
ywTkq0nzoMF9J3GLsdOM1/IXWG3i6iPdQ05b8t2n42tBvt+QicOwAnRl5ObGfvv4
EFzciPf6CApoBuZq+7VlIWVNE/VPNCJ7T4zROkTmw0EssceKNVXMOQt30bhz7ci8
XsJ78h+OpJfPgjLXYo8oBbI6gREqtP30Q9wyqtxNVDlyc+zJsFBQe2WMYfYKfqbq
aFaZAP0Iu/UXwuIqM3U/JOdySHqlqu2kbLxDYlRK45Mnl01xIw5M6ymO7gwMojto
cegsHYUJzwfOwnDpVPMo44AFKu5MedFpY1ilrpLRmxEtGdxQRYYtIfbH8u3ZQU2D
6tnH7Bfx2lNGKDe0/uRh5ikUhsGkwpGHY04YEl5BDHv92iBdo5g3d3AWDF8uTpqQ
jlQIbHH1MWcJ1fqPsqhOcD3D/QyItHMrjA9FqP9FhZ9mKLjyiiB2KY5hPCm5iskV
GNbOradz9EPWfC4b90ubn4s138G0Axd+TaPfJXccuZPEqsbwbLfokPA0HFuu99Ut
XLdel5LC9aiAuehr09r/uQDPE/kkU/cBvU0dxOU5N1A5nldGa2I1djT2fj3vpzz1
8nHEx4Ge1HH9J7++pYLp3KsrhL6VFUTUlnIzfU3lIOdl9Bbzhq0oFbZZebduiQP9
o7DN/iVVwevyQgVH8VbiBD7RkmtvVa2oVBws5CC2fxg/YcM6ByYWoyoF/xRQ2dod
H4ryk8dIYcbC1Wwk4aijyJhXr2AFMuPJcRyXghfTPvdfdB5P0kPOlbGa4L+Rq5pT
R1Ag7extZ1QyzZjP+OdeIfmedXJHy1Bna96EphlXi4EFn/WK4Gk9Upm/dQUs90oq
gLUVaA6ToGy02TfIMokwYKr6B4pnQuixq/jgGxUfqR7xfEQAldAwOs+sdhsIJ3Nj
RqJ36bxnjrYU4bCgh+HKcoSVgB5snJpM0fUceRPzBwkTDV4DD84TUw53f0WIbthI
35iLNLnh5yCtSKIzUWUsG2lmfXNvWwSxD+24QKzx+Ber2IbYs5FqpZDJJUIu0dyf
RFxhlJ3NEuAaUo5ob0H/7QfgiWe+1U2qNoZf+N0PvvH6SYVHBsGtvTdsa/qiI1aS
GkM1KoEKwEaxz+zxSNag7qvyIdv5xYRTc6KSCjAoCCzsOCaV2++SGvztjVMtMW25
WiAK0sp5G5UkdUS+uujDH09FsuyyZYngtwq82ugSoL95tlkar47tNIeHVO3pXxbD
F8dwbQgRl7MMuIDKoY5lzCuiH8TKZ2BbRlJtrMmNLlkqcZn1i6C6923Potpvi36l
pzej3t+vTOIDYADHnnEr97N/EfdXsgiSZgZ7XqT6LWVLJGo0M24W8oGTiUOnFGbY
vPmCv5mtRJT2yG9LAjLu/BFkd2zt0b6ngkcmu4UMvWx4/8z/LgAA+688VazRobuT
CygflQWp6U511zT1yvF7IdOFIhIKtt5Oj7TQnvLXcJSjfBjnwQwd8W/tlzntQgqY
H+quE97Y13E530v+3fwTiM3x5bOVecjzAsKhwJTTQ60WuZ4wWlafHqn06blrLnM2
8w16nmZiubBW9A1bgPYkVwLT04MqJJ2lOJp1FHC9AYOz7f5fvzzbtrheAv6LeNyc
xaWpN7eBSZj6c+rWA8gAkciJR3tKd8LH+nEtFXilJRuxTatgZ0u1y6depXAeUjkd
n8PjvYPZPY737uMLNAfghsKxSeM1jofgYdIMgh4RhkEQYegyqUiOSH6cwFS1QqAk
kV8I1f7Sjv9lopNIAulpP8RRCESpUDcGjzXgGRXFYaOR9zHE2MKrLk4cS7Nv4m6W
ksY93Qn28uupWB+ueAq2IITpJyibceSfS2CTz1NkoKCWb2Mk+p3q16phfPPxl+zb
ybVlAmWQyWfdTdJ2erBRmqOYngf0tUybgC4VGncS3Qh/dKcpyzFfIXJ5ciNEyReE
VGXCAj3qT4KTLaaEQbuPjw0V55gS3E024B1Tr6HxPYa+x6Y43YpINFLMXkEgbTlc
ZzcS3LPOnhFbvJ2M+tc3DEe7U4kB0yspQHVSZNHwVXMOqy4tm3XmWQUQyy7qpvFl
WYm556dI2tuOvv22QpCTpdrpchHa3oYPkE0Td7u/ViqobkQRKTXr3Xnltq6Pijy5
qYH5cCbtGn8ObJejPSRjWSL5Pb0jUjRFyY0FJXlb7o1aNIsiG471cNEj9qIDwG/7
FatsM03yCpuQhLIGzAnzeGT6RGdPIrTcy0dg8zyvfvLsFdWpO/6gekSdeW7Mr55y
T/FxClVRoHztKsiRTcCA2HGXEwQQxLNVl0/EqRij6I9unjN8/ePwgPYe5bQHsZWy
3hHLkqcbZjm6Zr36L01aHkjVX2HdF5wVBsxMLwJr7g2FDVVVzUl1l0c44gJ5C/5s
g4Yo4K27aZU5mlBFpc/FvQsEU4R253XPBy+JbDpBBHWVCyblsNOAjsn6joesr6mQ
woSntOHvE243d8JiHNMg4cZI7dVukYigaR5cXvwIgDlB6dQ7Qsx7bHC1VUVPGIwV
tW2CFWpuomhJ2afLk0yWKS1LSPyDCBB4zU9w1yaeD3emqtTMkhVfWb40MFZ2m7Zu
wOizHJCEZ9MzfcQkBA/E45a0noMTkpxZsfdoFOXzkffOatluqufWIxPoCY9poMd6
PMCxNVxSfB3wdQmFnOyV4bw4LoVvFKb/Nixuju1RYZhPK7qFSOIqvbSd7klGGdCp
r9roKSoHLANqmSh9KKLmR9rAXPDy/HL/FwW2a9LNdvSN+q1YJRS95rENfhGGZWUp
GhUxSCnmAuSdj8HaEYk+Qc/YCOdS5IwTfCWTl8WMPbhH/Q/JJ1LzNxUhYruXcnDM
34JBkH97wOnm8bGF9JEVRsOr8oSeikZ6IPNsJnA08ODSnaitZF7HaLhsjCHZWJHE
gBdtVT+mfFK0B3i4kAOeXxoqmIPPbRg/O/Y9D5LJOqk3x/UKzoyzDeAbsZQZZUqD
bQY3IcuG4E1FC9iJoNcezFCls0t4f2/26o/OT7YjUrtq1Q6ctgLwy4bvHlC5moZp
AaFSF9fWy3zYZeSnmrJ2QVwzzMhX9YZgGpZ8BwAGNEVmEd/hnAzdZ6qxa87yI8s3
TB8xRw5TOLLVLxNK9EE0TohBr2qMLDCRa4mwM5ASR+2B0XEaWk2yumdGfrmypf54
cl6NndhqHuX1yLl61gGWI9Lzl/8i1wz/qYzbw7vhA0kxQn1/clxJdSsgLsJwcmFW
52lFY85LZR/8LmNheWM29OYxiuHPuCkP1Vh/ZIrrL3ZAzW45SZEyrNO7r9TJoGFD
wqzy6aVYl9t6jILEZ9Sn5rC5r+tU24TxDznv2lL5aC7iDYjU3oRwNsFX2KFlBQGa
usWBMCgaMB0SlbR3imaFDN5IwKsTUETPrE3gKhf/94qHrNScs6/y9XnN2dpaqDec
g0upkrTEwN99bVj4ZVTOuRt28PvYHkQXqVsOv9wKBpl9ZN9vsQIzJQUlfNROsCQ/
qjWwvMuxUgYh2tcLP6D277n5g597v+b3ENyWmU1nZtMd6CKz5nKLn/2YiLLc6WjR
rbHGbwlHWe70Yb4lV/W4JP3Mz8WylrPEtsW0XUmwkGCGk58EDwt7fjD3YO/zy+eT
BgCgDHhW7N4sx1WvJlHemCzkfEmvBoniLU7gxYas625mqF2rm2BJemAimzfSftXJ
Y52W1dM0eZWjl95L1RlYFCvZgt8Vm0c2pTDKpDeu94Rn7aP6Cq6HQ64LPSzHtVF4
JWAbn2BOTVJtASKxc3PJXd/6VMJtHPqeS239+4PbKzuPdd2+JVKCu5tu2sOt5yke
G43rW+IghTuBrmY4C5Iu/2XIscswy+DGu1p+bMIhOBXAR7UBbbEJCgpDtGboDQQy
whtx2KCoOjttflNVaoexpPMGsIoL6kNJl/GYdwVXtFZdficfYD4pciXkil7tP1mn
iXvtBHxvlC25zUNz78ytSBDAXugKlPivuk2Rt9MM2k4SONhSLERZneDq4CsB2vN+
fT5FXi/4S7gAaykSeuhxrfX/YNrRGtc+r5fEmacUlfeKhgN3pw4TN89kfhX5M78l
WKLhk1Z23V0MJrTBbMAjh5hvxKT24kg2TEFqv0elfnvq4xX8gwcQq2oqtfoa7RpB
YLmYfbQVwdvJHcLppImyB/11RZq4DrptiojhDPWp8jHfguhKZQYkIw6brvTRbzBf
6KkgjDwU9HEzRaQyGwCLg0C4vBfG1VZrF074XvYbNQodDM7XU21haDMp/ut4cGZb
T+PpTaHhhauw6PpLVGAhzD7Q1M+g3wqPGFwI1QrqSUGH54h/kGCl3Lf7/C3IgiEY
Y3zUt7IQAh9UUZf51vrnYQZ771yx+OenxY/FpHuqr3percUSZtcsV798eQvfYfSH
zhuMZLfQIMLlJ1sGW+ZhhAuhk7d5shbKkE15RNJex69Blm1CKrRzheVsJYrYQgir
5cQNNnG8kGZ5S9YY0yPNrLXTidQRFULDwBSf/uttO6tpr4jiz5cYFn0mAqbH1Kt8
SJlYPjRZCrOFGBmRT47FC/PHt9KtOeB7Qwpe028Qla4W71ymesLa5ORwF4VCTyXn
GLubDCDBSnMffaeOGuBkNQsJUj3LJaPd3e1G2tAKFEc06JAlr8TC2pzsIi8KCTw6
xcXy0xZKmrNF/0PQb6HJvncXn4HDr43Wq2VcJKRz4ty196uIsOZ9jDqMIN+vA1XL
a2TD4TXozegJLdll5XgY3vHPoSN1nVQfgwulXuy4Ed+/ObD1Qess8L0tPV+iUmF3
BnzaKWwTVDvi5RCVM+dQ2c7yHRI7TwVgUjx0/pU3xcWi0ght/lj4+BBKROIiU7uq
mcjo7YqtoXCycvVXcA4mjxG17QGps8Aeysi4XH1s6Mgp85lwU9qu0r3IA99sEZ/a
2YvcCgIs1kW/p10ScgmUZ8WoJCjqDhQV8/ONC3z8rK9xoham74zOb4LQ+77TTPAt
KjnsveGSYdSv+g7l0gLFeTu1B3cfJZJCrLAJzJMuVoL8eNxJjxZA5qziDxx8nO5Z
Oa2zzd7yGX1MYX54CukmWbLiIBKt4Nt0MGHv6ni3hQ3+k0lfojx4913/Q3D0460V
23ThbSvTG5Y3fW3YZGc9/YG0/OJikB6Rv/6Vdrxs6p4Hug/rQUH0HKLs5rLN9Xgx
li0CrYLvRINnyJT2F6hKOvN0zXF81/daf18fQF20l1ca2Xf8NCUXaOB7W7jr3Npo
GAXfbTEMwlCygVYpylJgex5AnOEBFQIv4pP9/gmveemGPTgb3Nl75G5uuioKyNfw
SNDcvc1baMeSIM22rtYUXrJ0nwEUbLBFvgZogIQwgVAsgmB5whVnBYOMEmsAeEVR
I0GssPMlflIlAtaZl0Z2XyIqV/dK5izeofh6rVJm3gDCeu3cXw84suhdfWQeYu66
XPy/0n1Z4tFzeOhZ1roY74PaJKZEP4rE1FWMgTfUU5MgGck+QsOmsv/akf5GgsPI
59yvBZznBnyvH4xVzI0iiY866QALbQ1pTrpYMatWGeFNv9Pbp3c83AQMkFs20GYr
MiOq7lNKy8NQ4ksNxG3MLiTvvHex79YBs7YybPWspmrwulKEiOq1lt+4XiZwNVhP
WF/dTBwoUAogTcAe0bZlpn0kCkDCB4HHdPb6x0ygM1L7NaaP+OyBD9kFOnKftnTO
WhHKElgiFW0M82a/fAK874gU12el96KzbCxRcy1rB+qq2SVBP7H2sdQuM39PFaJN
g9Vv+70AsAs9wT+rhRoCINYINJFWqovw4Z4XiMK7qWBbJKoLxQjuFSOhVydTns97
wPCagfAyyqohufstBzN8tFu9z0hshO2aEhH41M7p200EKlm47+cBDOmOzBRIw4OG
zTRn8JX6X0Oe0+P+5epJBp0d2wIgIltclQKrMJuM6i1RaTK5D8oryYBnDaYuKnvy
cgL9yYVfvF2DuaESyb4xk4Ue+T7mwEKQnHq+t4D+nyzZouZet5OiKHxuxN4O+jxQ
JsRs8S0F12z77yzixPmv9+uEUvPy6L0J5K8f+aDwZuJlwByft6x7qKj7FK1VD8Au
a4q7WwK9YAbCjQ0EK9VoHlVwQ8/GutyUjRieAW+4bB/+Q/Zp36unL1gC36Wh1W0j
I2eYPmtwxjzPcP8rvlYjM3mnR35hmWdWwD+vcIczAspS2+TT0VAdatIYPZcE6k1x
JTj3PFlDywNZx1kS0EUSV+klR3lM6anWtGe+6gCuwKfYEHXrg4lpfy238HKKSNx0
HWZBKFjB7x6vO0RyKbz1KpoDfPQ2scS62iiHx2pum1gQ0hi28LRWOCk8sz1mLyKI
KAmxs+qwFgxTChqmNO5MhY1gD0/g2lms7h78wBXdLP0EofQWf+IM4ShLlxwNa4Ro
BwDRlLeekGl4kQlryLvtIEF43i5yAufzyY4T0kt1xdwv3QvK5BefWc+HxWkk3NIL
1gy3DgowHUeSXL0eCWhZHQlab4GKrrghufKHSdsfywzsU8U0/MewJKsEaUKpda07
4Oc6e7vwLLiYvf/TLMBfiGxnMISCpyICAVJNVuXqxyrIOk/N/LhnE/NA3kDrhYgQ
6r/FiwzSi+sjS4W6vH942x9GXzXDuEh5umLz1sU+dC72Xq/NA/o7Sg+QAN77dhl1
w2mzqQWFiNxKXuX27rNY0fwLRvkVfoHFQn1ZCB/O9GfekQgzLgUf7wHtVcYDieIj
uDx9CmOaqDQERP4dG5d7kCya3k5xUn2TTX6qnfxkpNsNDhxHWmqj7bpaQJI/9qeR
5VVYZn3/C6Z7DOOLIg6KBAIoaetov8VFmKuyJtT2zDYycbUT/sbRDQ8vOPGil4Gs
Bt+iLWb1qtAI2tfVjhonUq3knbHHWIyZoVZu14/vROfWMZqLroKAFSLy/oYYYlrA
mV2iGXDlTDbX/TOwl3tBn5h5DwpuLu8BAGd5oNjJN5bQvIxfNOzS0eF3eQKDI/Fj
kS86ZNmsdS3B17uhBbiI5HviTyLCUtABsyqJlDOTt6nGNKry5KsX+K/3fXx5nycA
HrYGcCw2yBzWHD2blA/sRMZnvFDIBrXq9CVIOhQiIQ8lq0PlERlDwyGUG7m3kNkH
aSX1JTsZl1WDgjnzJrEtt8gHg5gJrsiM7fUMIXlcOH7ibOYCVEr36zNQe7Sszt0R
wMmqbZutlfBsQ2K4JWjM+RZ7Rq2WeQwQotusT+cQaLIgET/HuzPV2bhm8zKesZg7
NtfQNk1rK354RY6o+wBW0CDnnfK5ze/J5Ey1FvRUXXdLPjkYV9eA/Lj1bA9QTR2c
DBulxBvLVx0cglpeDzXVme5cQhLuctNwNFJE8RD7JNxqQntPBx/ddvwtRUwZSMO+
p4XLjxaoAPOK/yz7dATX4FZepxmmMMKwHx0rP1j2mtv2M8sVn50COQJ0A6IiIZ0F
xYZpefsryV03scO3WgITwOvueUkY9NDR+PUhwL8GppPXi6Vg7D6qLnZQiiFwFWj5
HKSqMIuxTenzoQh5lh2FFHcdVL3auDnpKgp1b40phDWpDb6k9ogMHGZvulLUWMCj
EmHaEoDyUq0PdEPGc+ThaYIL9WlB8AvU4gC+gysBb+k2XvxtjyNAYWrr0Qu2N7wb
yjUTBP6SICm0M/zFBiJ1DMujfBWyt7ZpbKnv/HXgCxYv4GaoPuqad3TZt/TmamFn
FkZcsfvtIscglfnGXaHAjSlTnk18dolNU8a/ECOZf//QF5+6LSqhBQTWQWs7Zy2w
biNdemXJAQn5ThhtPMhZ7SZhMV7S5NH2ngYCQu+TU27O4ArRbuF/rQSJTyA4r/jl
ms7dsD0Mv5QI/WIjRPafx8TWht+eLfpwXFKkXMXdc7C1NVDjlkV21BzACPHaXHd1
GmDpnKoL21QHkW2JePz2iqE4iqGKpdQE5m0T2SWrXx9z4UMowHRJuUF2RjwamRCB
WZl+7QwteKcaAHdURlk1LfWAwwY46MtAiVvHskbJWocBPvQFgasij0pc8cQzqONM
kOqfvjPf7Vy5L8UNqqigufFP0K5qRxMLBN62ub4qHkBVQriD75rmp05G/Is0XFI7
FvkuA3rVXd6oTnwUepKnbnBY9MCkPJOsBVdBMm4FlFRD9MmbldPt57lmzTssrTks
p4S8GhGFWeogZyUa/E2gUUHqWEjLQRG1V9jl8os2zAlRihwq9F8pKnvZYrgm60Y7
H2jh1VFzN0SjgM1NPiZ8CpNhA6emSAgzfOjgIenaPAWvYs2LHXaMkWTwXGqFaLgz
xM4YQraLl68mKe1LogHAuf8jASfpEl5czOlVx3q7dTVe3eQmIpKZ4uKeIcnCvI4c
a1pGm8n+s4e/ZMrHTfUI4FcRn0veJHAAuolEPbhUnrBctgVIZXiDJuHRgkMm8I8p
qvlyUbV+OwxO0M08u9LzenGN5nKm5eccFzZTvSM0KyBhrfjI3MwcUuFvm3IlUvvW
WxVLDLHaVrzONtBR07pYZpME0OBN0i9/5KtIwCzdkukhUNygt4RcTzcAiNgiNSXc
MQaL0o8pSslCDJJISi9kOf+hW6FqgIXpSZNXwaL5IIGehDCF3KOnUk0VZoDfdm+5
B55RWwBWPBrpVQQXxfHFLylcQ9A94/McZ9sxNt+o61Em99a6uLELPgTKqCzl7/j8
8jgYnm8KPTwT9S4B0/QyDz5zu1VDeHXOWiOsVfJFofcIdN7EI5fNYobUJ0xrgoUy
drcWPDmnxWelPAS/y+y3RXjcHffraRKBJPxsFzs58GPminuCcyRATP1jAGX/5+K5
1Uj4NBY7X54k2uEsCJAw2yfWRGa3Ws//+aYvSs91HvTZxRsNorWk2egU9qzWw8Pr
c5bNquMFNLcXAYluaV8k6pcNdxs3zkjQmwZFg/G2sDoIdJkRoQFoGJiq/yFu0ZRu
pGySlCLMSYV3Rii5UkdnDeO+3IVZPQlePKEup7UTIYnL8vZVZbHaW3z/CbImQH5H
OLfo8qlsrorC4GzdyQorZo0sdSsYkH72X41vveXyPck8jGNPaCoPXCWCQbEssFZd
FlXkK4frj19FfmpM7Y2Fh+wCWhBOhbQGXfdaBx4RgBkAxh13RKqcvb+JJGa0nbF6
pQvrI6pXaj+b9lXkYiLG9h+LfvjS5Qsc+bdhU5evY2nqvhfkYB1RK5ZyQeSOuCbx
R8Fgz6JkNy/oxULqr67nyCWjLRUul9tao9/29zZs8+wNCoAxsKuswf/DxthDNdNA
5vF8C8CEmWcB1TzNFqX20pU9skSEXbaeioOVNaETEGw6UCN2T+HmoSYd44eSUbl9
TVQyNzFhCMLkIcWtDtoTSyoGXfCZmVKDenLu5Z+j/ypNip8ie6qNfal4eSeJa9jl
Q5xoudtNqfhs6QtsVd5YrxbEIXERLc+95eY8VrtPUwXMDhfdrkxwAxFKVByp01xK
Bh90Fzevj8lx4fj8LKOzDRsycP9nXZkYcYVPMY5S4JpDTHJndqzA2wfk/i1VYZKF
otz4HkHWCXu0InEnD+puTV05zfeCWs20qFMJsOYQ04z2UaBxk9VPsgxAPYkv+iIr
zVpIkqjljq8M4N+SIDZum0tZ6BOwvX7xxrq65zv8+j7DceviF5WFkC2VZnD69AK5
rL8Gpy+/siJxZQuf+1m/GjO00AVEcOrOB+sicS8AJpqUwePAg8xWerXLlB/Tk5mF
580lWIwl2hc4tsVlZdXPVUyf+Arvf4GV7hKSy3Qr4SYfKKpDhtfcu2UXEQX9axP2
t4MBzINz9FxWwbijyRUhfhurx0RhkdWeqAPB/wvxvYQuek+W8cxJkyKIbT3o679K
TJy7uEen4Gz/sAdfOaBHIpGvEVjOxhIqlId4x4f+IKZ1Gw34jBk5ldQspoTu773r
19L3+RRyazBNtKSM2ZSEPmJ6bvOt14Zh+tjSk0XvVemnxniTLnMzuzwbWp0wSXJE
grWVoMbd5tomQVnK6IERBVZI1AI/jt1csfFOJyrodAp9P79VGXOCWCpHVJlnkUHV
DRvLBgU2n5HhEwfPphtWwCj2I3knAAnzxxhHDZti0mD18q1e+zfv2ogcaQyVHlo4
kVUpoD50kQRBMQ3qg60icCwdWzo/85yVUWNF+1Q/+T1BEt9eNVsb9o7ZnEoa2fct
Yl25ucRBS4k9fE1ZtuNJk3jHI4COGaKQaqdeZPorJcjNQTMlgGPQdAKuyOKEdemJ
GCS/cxN8OI9EcIc1cojk+dHjutiGIQWQBDSIcaHzz+VYSeC48O7EnjlWTh3R5AMl
ecF6jYqLUjM3ucwlMpNEEL4cZ/gIWqJOm9nyDTOitcGlaxTQQwbR2EXswDVchwWJ
pFOHO4ZHVe2FTFa9KTemMDlRtWcj0Rpu8AqtjwMBcPEhVj1JhdJp5SfKHAJw/WxA
kI0opDoQ1EwPdQ8ThTuLE1tn4i0PqlV6kjPJiGNjmP2SREqirqxPZi4Bbu68R9Of
HfcXUQHnh4OFLku0kBghgd0JPbvHmkD/2Xmm4TL5hewOsOk+Z9jW7uJSqn15oG43
CuY+kGUTQZrcGCfdhxQP60FskWmPFnd09eQ0TPRo8BY3zRcxR+K10zAmIk+fNsrz
UzgM41G7sVu98gD3iA08Z6NFRcza3JVQP7oll2mJJlqfGgaBvDvUx9JezNfW9SIR
pub7zhNr4ERFKO0i0fDWgDX3R3ArHhU8ByKxlG6YPqa6NSar/bsBJuCH0fDDJRh1
SZC/FddOKKTgl6rTTbNoXplQBS/1QRCojuPVtJwjbV2KfD1tayf3CTZo3qdrY+Zq
itrx3cmCt45h8YVwC0EPqV/FrArIZ0sLWn9WVqnn3geK4UeBANt6Cpx4hKPLFo4d
JJdualcuBgb28jnUtpx/2wD/1lIjDiDDdSpzimhd4cw2Vc4d+YaKR3QN6RlBXQag
ojPk1I5+PjNsPHokwy4YEX6byehdKwSVkX9XOReo75ytGDNT9pnGxEpX1scY0ooX
JqCQp8bic0hgJkg4ZDNDNv+ewuzIbjCDPHhxvr0orDcb9AQgJKqQxluSEQObB1C2
vvENl0SrPXEbC6zmeO2GDuRuevW8bkhQeGsrY28h2zD3Xvl1ezQaYcMCgVbjKbv3
hm5YdZk24KMaYlOuzC99AWSC/N2Zx4Y4bSHMZQpIOtlFNEYBKHg7DMcY8P7cqwng
PZRz4gjH4ptxFCu02V3Ob9MB10vzMean/yGJYCC+U9h57Vb6Ju6ev0aSGuNtBc07
7kLuLY2i2S89ESE8QO7IlWHjKqfR4yTRu7remOmM4ejIIiyhZfLp9UgC1MAw0+Ae
+vTrf4sfR8rr85jkQqzONEwSXANPl/OgPuYgMRjyIs9AKUNvook10yUoaagBgncw
k2P6fn3WVMRzlrOKzwhxQtvRqin20PMtIe4QvQXu4fE3l9T8gbaNFEe5Q+bDfJmk
6wjSmkJ+In2R/nuGTViQ5ZINhCNpIJl790mVHN3zl2Lxezt6vGKwS3zEqGAvBdUJ
2USXe6WWoSRY6CBMyzix5I7C5gI2fIah08MWZ8wpl3FCkvROSD3zrMXkQp1mWu9K
G7PNYJmycvh9ifo3I5SXoo3o9cOvRAs4/znx/q7EE7iNreY88FQADYwwxDNePOYC
KujigxqdIM4N7VKn4Zn72/vWx2kBy9ka9iOmTCp09KMADtMKODmNK1FlQcxRiFns
VkB6aSSP2rkFp8rNzLEWFmHaJSHScGHt9nKUfJ4cjlhoUS4s+00ezwCEmniE8Onu
qWLPPNTkkBscb2Sajxx2rM/y9nndo2boJCOnLbFPWomdXqXqzBd6JPdtqzGRhdCd
Fu7KRPzodIbuD0U4BDLWbkAEZW/vmRKPtbsTCZIzBY5UyB3Ks3gSs+c16g1A3Iuh
UQwDg7emQIMYp26ckG937vDAeGbAWrqQWrNHGFy8PrlCfWTbLiQXAnWerD0zU4Dc
ZSa81ZrwvZ2ed/1MsdLZlkEQCnrmmDfQp4UGzJLJi0Svk1qsLCWx23N1ckrr7MIY
C5dixbpGi8MKcXFJBLKVuJGd5FPYWRjN3sHHqU7j5JwOwd+WhzDZqyPeyj9yrbOY
sVHd75cQqN53ibLI4SaHnLz/KiX7KL1qHh/Sx1wTq+o0b216V6NMtx7VMhV/f2g/
h2dj1D73jmekfU24uFoRNVJxOp+H3jmFx+gE1WMaknhaJfX6Rw5CVsa8pVL+X4d5
SM7mtL2T0S8D3DNfgIj+cDWa/sxOZLTLcxNgugvup6Hw1xOUH/pcDWHEfWXQSNyo
E7sBQHwPrAymRdbE7Va1KT+KtdBS+1bGbtVDFa6VEj2s/6nBBWV4tYVkzriZb0HU
/dg4eePJg7K6+S8i/cgJnUbqAjoUS6PcVzkI3EqA5laVHHKgjsiLMhVDn2jhbpG2
d6owSRgkvYb6TXMrHAwaQ8ofUrHc6OlVMNJaQesFxOgoEk5ZFWsAMm58kgPyW8cj
BCYqyS2kQ0b80B2Kt2Yq0uHhRr36nf56XntLaR6Ymi9xzdMfIdDw8GBFE0C+gsq/
7JHCXN9imm99yDwKbadBzhFiiXCx/ZV/RHeNGoHJ13+4rLfj7Vbf+Ls3uBscrCVD
krUCr3GefZwYCscZH1caXFD8WnrW0gEd0ttWzQsaGaDj6DOh7B20fr1LiIvlPYiK
RZaxlNNu0dEaXKq0gDmbmFzssQw2gzRJ+pKW6YVZTJLJwMcMkDqjlMIl0RgbGRIs
8rnWKbUNG/VTsFcrtLj08sknTW6lRqHUac6aygTRJNDhCpcZjbAaX+hmHaGoK0zF
7uC4HyEpudzac1D0079u8BTzDg31HY0csrDmpzuuMuw0nJwPw1I8SUi1qw+nctSh
7lbcLbaD4aYSm/veM4MRm3eFti1ihA8xLeAWzg/ODzMawMQ8EQ9/lqI/Dgtg0qd0
Xv34Nh0GzXq5LMQBoVuRaPH98wkwWKuZ342mzE0w+5SMvUP3ANdrfCuml/5ebVX3
Tt/QPuRhfKoomZrl4NAImJGsZijCgovLFq4ReE0Fqo8BwWaXU7mAUTIhY0g/jq84
ZXCMvYC2PVSe2/zPbHD6imEJ5TD8eS0myetaWgYBtxZgWWwuImIaT6pmcVFWrQJU
/Ojx4n92SMnnnwxCC6GWe0La9nb6ijbTJb9CHkzGxZ2FL6m/JzaaCTxEOzFqOXIj
lK8nfyR6ePumi1aXZaNokAHKcvNGPUL6Y44LEnN1t4ZpyaZ0SmNb/7tncfT49rK+
AZmeEs94kHrz0QfuYIGO/7JnbwIH5qwnsBNXxf0KG9niHz3lr48sgt9BEJE2nFVh
/8I8iZu/69KgIVa9aCdDa59OqbH8nlFoRl4qrsNCFE6Mv25BPs0S6R9t1l4/SBgd
vmyw0X1sT1113Bp0PNH/Y4MQI2uPPLXRXhVKIrkeCWNd75FpVfVVzViRxxQNotkb
/QuNRykl9m7/IPmTeWaINQFJzVKJZ9v7oLAvNb4JiWMxDXNgR9gOhp6h94QfCj9P
E71Z1mZYJTSgIrJE+S/5YryTY2xSwDbo2DPIbXpF7l4INEMqG+JzS39ucwCWjv0E
cjVE9I60zDOt9SqJpKIT8HoBywN/yByp8VtQHrpwT1l4IyQzTlrp1zv58ZcdbQW5
K1kaDFnWCPp0oZQVWzc/oXWuhJ43ArG5oCRayLU2eQNMjH4FG6oH/Z2NcZVk1JFY
t9ipce5duf0s5hBx0oJ4NYavjv/XzPzz5lL/ildkX0fi0Zqu3llu/Iz9ihIIHVFn
NsXxBH0Hic3p2wqXtn/qGBk2y9tPb0TIgGGDryVByKjBEeSzT2qyQaOXOjck0PPg
9mhNNy9lqH6b3pLenmDL2JHafPcGBWrC7+tLgj9atFhkN0OuXbe7IPwerVM8xzfq
gnR6pyn2EdWYoaAmBcLpWmXWiajgTKx+ELDUV1criEUCILT0ALLl/Th5+lGc0/uN
SIgByUCY6zpQLdSDLe/FufbfsIPpEjtuEju04EHkY2syjbBjnsSEMYF5vniyupwq
Qc/RDfC3Br/JZR+5ajGgiQ2xpiLsnY0vjKyTntaas7Ida1n43rHO/cuvo6oIlKG2
E9eR86IE3qINDHcKVnAfpS+dQBQu4ZBXe80twVs/Fhwt7uPldqTCwbtJvvIlv1X7
sNr1LxzYjavFpNvJLs0SS8GGLdiAwtdAXpI+sNpnsc3nBnIZ7Tt32NyTf+BYs3j8
AcYytgbnACceS89AqQacUN10IVA7bHzyeKX6RD87swIpPeinwQ+Pp5upphts4yPt
CMhBHwTjpOBKmbb9Z4XhtFjJyjjnj3xwQOthvV8YVZdS3QCHrFlql5PieJK7bW5j
B3NfbK3t5I7Rt+vs9Ild1zLggQcNy1KSRJ/Fl5FTD5hyJebHp3QC9EQ8qhwFa7fS
95GDQXGCmWBmr8hyqrqjvespLEcgvQx9DN5/UYZdeRklHPnrgTF5k0jwHrHZGSMN
FtijCBbLMcrrRrt1c55iMMFcKCDbAXXmQe03klV4k1rprbgSfxEfmpFlQLRW4Lw7
WUAMDE7cH2GFOfDf/63xMyGQsr6EGL8cujYk4qkwXxa5YuTbMZJN6dAiZ/RgmvkF
KA9ALTz756b1oBWylZKZLWG7tihx5vx9wUcqfu7M78DiPh33UL0QnPooz7nCk8c2
lknIxtqH68koQiJmnZDJIx9b+/4is9hah4XjKC1cP3ryEX2ecBJSi+vFzJ9wXxxB
/dGMdfbVpEEerSj7/5NOQTIxjdZzVhW3zQ/T1jdh1FsCMxP8p6gvIotFYjugpmfa
KjRqvYD5L9uzL9eJCvIoSiz9cPU7Dp0cN2kxs2KXfkXDeA98SHeF3sbUb8CuLDfm
BTn7+hODhIPOPmF1ReSi9V6jKwfJhzGr8EPK51LJzoYX5+rviLNri2oCHi1v7Sb6
j1FhRJOGA1ANniYOfb2Kf+1YnLowk1ZSGup9tMJnJLYjCefibXTPesB9Ia3xV6mI
kjukMwHBVmhuQs5TA2THapEN6FeufOP08SPpBNKQEyJ91+17/jzvndiAULz5t6rW
LrasMtbvG6dBsNF4n1DqyeR2Rshv6Mth2PM0TDwUw+9SsaUsTQjEEz56fQ9SDxin
8XEaC/UsytL0scsUri7hU8ucBrUaIpje+027ZWYeE7XIdSsJr5FnBt+bZElBwNPE
HSOyEP8aVDSZXv2vInAaRB/LqBqDYTbPs2xzlUr3dcQBrmNUNFAMK0J8DInBD8Cd
K5vjjdsBpepQK8bpBhRsUMXKweNB0HVu1ULgfvXwXzPgaZK/P9xJw+tGjLHhW5CU
grZHsmbi6IWTvlCyjUM6q73X5BA0T6ApRbeCokx+5a0+yxuOkjVteafCmH0rVNXB
ikm3/LJDGnLvVC6NiT5IMzUTD4twCd9h1gIstFlL1TA3Q66hkAiK+SCI4oZ+TK1M
HjHK73zTaxJsd9uS3SSLn/IYpRoyfEluLGKGwxAFargte+gd2++8BwnxQhgAT7xO
qWwh+2U2iXDRsDeQZoFBKToxyjrITi+aYbFyJ9Y20ZdMRyCbgs2Hxv3w7Bjvl6Gp
666B4jCiCY5cLVyMlxXho0zZcHGPHRP/JrN1vfAlq1kxT65HgL4ZalCJlZwYX9AV
7PNdUKk13c4E5xipNj/SVcrSEWIu1+w+feZQ+FbB5naR1kLBMlzbqaqka1wEtwRe
EOYfUF12n4VH5hVTTE6MYE8IFsXGThGfuwNOtrM3tk/UFyiv2T5C/YSCsf5aMogh
1P9Lc1NduosuDs22cfOocszqoSlhv+2zXcj//o9rHgZRHHmxc53qRCZ0L5+2NZIo
0fU5a4wjjs1LMnVmROap4VflYnrQr3IfIUFvUCvHcZvG7Es5focdSca/mha4ws9G
M2LZm7EuCC01AfUofIhv3A7ho5iJtGvqtnFlu91xP3WtR6xNSduP+Fwj9E/mPpQt
tf3dypsJUEW72Gk/9ro799Pw1gSbWy4uREJR0F9LGM5smdb2zJOM9BhCe8YM6AGt
o67z3xvKDBg5a3cWOVQs2XgHRFCSMA/04AufYt5ABbe/y5J7H/tFWkcEVy+E1DVM
PaWAJfVGZWj5pY7d3gkfQpF3CX3OJngtXELnqo/B881A1hzbLiCf6BcGVKGMGL8Q
vDpt+AyUY9537jDHEd26QML4i1YqRvOLhogVpoLBfeTk9jXhbL5gHRWr0lkWhv7C
HyOr+Oym4pm3dGqTvFWQYTHlQhi3hOsV92oDIIe4TOyWAkTJ0LVGiUjd4pQ04muK
2GDocTgLq/Izy/fW4npnPBnhObmmOJ+1VrUaXxksQjv1bCIGXtkBozWMTP4JKMkP
VwHB+84LIA4COqbOdLWvWLtSCpTCjVhH/J2FsT+mh/SGxbIYe4sePmC8QQ64WI+d
/nONrV03EQuyBS9gOJquF8p/KYkTLgLrSZ0O9JJrA8Bl8IFnABpFGqOzh/RDQ+qN
HHzgBgfct05YGrenmDgtO/g3W1mc//57i9LSn88JwISvcp1bWiwU6Su3OvMr7uZ5
lZiu4o+B9mu7btsWiLXhme/xzXbzU0M31IO3Gr4XX8BXs49oaxgTzIERVyYnN9A6
c9EmwtPlQK3VenDbmrggJxWvgJZbq6iY+8oi1t3X5h8yqA2qYEbIp5Afl1pFSWzV
pJAgX5ybZIpFNW2Csk/05Pe/qiWaJISmXGOyyiVPwS/jMoLuyBNr4Pl1jhGThlt5
ipZv/cySjXj8DYFQFIuMqfQiBOlUKS+n9cGAXBD+nGOcZTFVVw+OAfw6vT+/wRNI
u6r5GJ9rA9juM0NoMG6TP+4iocm5UoLj9e96M0VngDnXvbP/usLdCcxJOYWj/z2j
dhg/oGya00vNUZ8qqkb2QM3obaS5wFBdkONL2luCWIkuicfVpp7Dc3zx9Ao43WG0
uyBlC+rQYPTOtDS/IximzihbSRHH6SZeFZ2X9jPL6NRJdcljIpp2hCjra4BLUq2x
tH/Knc9wXxur3UBW9eX2Dut4FlAaX7m4Qq699WqydUIkDrRh/Fairwg1H6wya2NT
T11qpn5BUCIMERKSh0MqEA5Nd3FNxPnk5jwcvF9+TKCE9GKF/ehpYQ+Tmh5Fh6hR
6sIzuOOP0FhGkc0mBcp6iA4yEQ0jKFokYG/k9F/VGly1AzmSut2JHpMlfvJqQDqq
Mi3G/mkLXRsEK0WrlAB2EWlXHxslo4tIfGJw9edef4zpG9GODlHJaEJ4O3dauST1
ubdcTE/4UVGzFRfnAqo/pqa+OHTPj8kP1gHj7lKNAnMz5+qXek7l+8B3SEDjzC3b
WxGrx+bL6oPgs7aDQe7RhpmusgVRowK2QRTst0H0zm/S4hsh7kWFJqYtoTkgHrRl
qfJ2dXhszBokko+Hm/qiKN86uPqWlk6EhSvozz1zOkyZjZZCYXKxxlNKVgGHZ//x
BM19C74it0pMl2S760564n2He0IjdveelFQhZWNZhF4vsZ2CZdOboAqBBGNf1XUE
tlaeZ9vlXJH2iuzBcL3fjxQlxHcNSZHhSJ3o2h6bL5nEdY5CqVk/p2/0/wtzXWb5
8elL83bQSFtGIgsJOh64rCZH8T1pWdqX0bZk/Jv/GMhNFv5/Sos6uXbZPZbsoOC7
jbcYWOhhFN29KX3RhBAVbzZ6VpOQ2p26vEgrV5rVNLNNaWCw/q0IkwY+d1bIqT9T
Va9mH5LlhsZ23p3pzErbqgFmsqjKrA8K5vD7nWZMCouq9qpHWu5WJ1NwZINEqwcg
glSefhAZQ1KuY8wjV0w1T8YE7enl+KWlfOoxwD5YoV5POHuuoyX+pm6blb0z82IU
QuJ1YtPxrTCbsCJjE9Ynaq8ySTqDjHfhglrcmVKDhUO2AdrpzZsZuVPo2drhp2L6
wMVgRY90DPWu8h+xbnmc/h7TyU1vQeT8foEU5sGzZXdSx0lxRDitto81+obNpqc7
LnE0LTMPmtS/LKeDNEBYiaQnNv/MOboVrsEWat/XSsnfu2wXd1bIXtXin2A/0hMg
NwWP9kAZGdUuv4s1vQTF1EvQmSXr2Bd+m9yCng9Pn4B9QrMB+C/CH1EIpK4K+VMC
ZkK8FraHm6MpXZIgaL0u3xx1nv0Ga3R5QQAsEwAPiB4Jcy1nRAex1w+HHBzi83d0
mIe30k/n0pu7vWJ/atqm2PT+LbnX0VCRXzbjG6KgFGgMlG42zJilyKi8IWUNv/S3
9I+WreNCl7jcpmvfhRjiipm5pa2oDUB+3mq8S/o5xHp4aKSh7Cn6bjYyV3grFbeM
t08ZnxpaVPqGecLflEpWZow0JDHcDeRbNNE3SnMWjzIgjXnU2gWeCM0SbvT4AZ7H
A+b4e4ldI1NESkJ5Bxll8wz0+or7S0HUaGpUVs2oYeyyDGlfkcYtA1nbcAMm9QhQ
tpo2d1Z99RGolO6LP0K0HXrgPK70mCFiffOa8ju9RHn5dZ48iZ3skxz1TCSa12fe
TgnCAKqzRffJp9ar60U3pVG/8BZvLkKiHwgjUHXkpHZ+eM7WBJR6+2V4/nrt2CUr
ZNwLUbgqESBbBes6ZLqDyego6xPkUm2phA6w+JNkeDNvyCIckthcj78i8u/FZDiz
/7K9By5A89r0SJhcip7GxKl+nunNcGS8phTj2ztnkpPZSru9pjJDdjGZfTBwNK9u
zgn17bdvxx992J/+K8urM3GfNR90xGINoXOymaI02AeTS4rvsQHYzgw4R4WN1mFy
UbSYGvyiRjOgd6VpLe8FVdcUfWemVYk6yxpNphP8AHfkLcbujM6Drx99G33Hflu8
VJ9w1zT0NzdQHgJx5lrm+OyIlQxYei5M3mykLTtK9z3Zl5YLaSiH9+EaT+kpSTnU
97Q9YIn8MBbdfTt4ocQMhYqxmnUIZv7yq3aHxddnZmyO5bXTjRL6dFu+ZqJJMlX0
F9tYTeCUjMIHMK+FTrZdtxa7FqtyJ1hkNWrGrYtTSdxr7FgMo/svz22KYTqxq9Ec
9QB9L4+EgXo670+oS0nZ7MVIthKcrtYMx/JGXyvMSJFvTiYd7EbsqGo9xKL0rOZX
+PmAj3WFnN3HweXoqi8nK5e6gt1UK5aoZlbSLc+e502vhHSDBdffQl+O9txWWTeh
4+nzpnDf2g1/AVD3l9opT3bT+uAJDe0uyj1RRGueaMLvCMx3dzqgWq2fmWMOJhJe
KoTYSsXaPT2VAT8VVlhlOI48GOzQ/NqIDf4PA8IL2+EnXYdIPtJzM/QVctdIOYEp
immzgWHTybM88xAQmnIZoQ3G1woREQybah4P3ndr9HPZ4D7scr0vwSC33BlM9Zf+
grtM4gOCs2qTHn6xWmfamZbAVxKAk3QhC0NSC4KC7LQTBV2MUw7rrFWpkhVeO1YI
qav1LYVepMhbliUk/XtgBCYYWALzr97NoE3pCi61Woi8zixD+kTq/h4r/N1RaPzC
ZURDW0bZDavwFiP+676OYj6qo3+wuWS+Jxa9LsEtdb6YV+2WNIKyAG8tOdB7NTC0
koOFvoIea0DwnxTTseFY7zFRH/s3323AZ3difciDFB/p8Bo4qYY/uiUasrwTqIND
ykaeFBDE5lZWatKMBCFkII2beHDnvxsL3NweFisUP4ez7Hkp7nyZgcplbsSMOErc
cdIWA1Y6ntErhD/WNk1S34v8Kllbi2/gn2eVByGqlHQg8AsNff1J08j/0cblheOG
3M1lV/cwd5XQt6AlU/xGwQcRlMhBwT/YPJoc1frvAwJhONwmXqij00gLu6pjKOYV
jK/7dh36fhsKgUNuA2sCmQ5KRZnC7FiYlo/8MIj8XggdX+5891R/RbOv5uklydNQ
XgFMMIIdR1zjSPS/11d4tcYxvLOihqbRO0B4L/G1rTC0/BL4ViOI2clmOaRSYf9K
cJdfKJLxYIWcNUgD9VJjIUiG7gc5X2FJlPz9CT/Iz4CeIGJkl+FhbUPV/YN+oaJW
J5676IZ7+WTKu+hSVkvUJzkEQ6Jxj+aqz/IKts60y1jGtVG2rJJrpeFhot1H51KS
luhBieuT9rIH7SphjVsBIo1IUW1csGb0ZbXbpa+C8Qujkqq4mQtVK/NXb+tTGFE1
LtUgHpna/B4lOA6j3B7P15uEABeCWViPLA/79MX7QGXVLzHorC/95vHjgVHCXuhk
sN/LKbmBK0GUMn2JjGe4gOrrxFw71tGj+VDrfQ9WyRNUcimxpySo8Djaw8tzqd9Y
l2RQqqVzL3rRnetSymN23OYMKzSR+1Mztt3q4Gxt/bszWx0QkPXkGXbsnuAPJwLj
QqjCw9l/G58yWf4jNboaJkKAhXpwRjBmJ9Vl8DLhOelXCrSMcxMkogn4Qf1Lq8l2
UZoiqqW0s7afl/ju+S5MvzDlx3k/4q1cbTr0uJ9f2oQMh8cU3uPJNd4NuAyeIji8
5sOzB8JsL+D/pFtyBeY55cTSbN/Q+qo9lOzj3mifx8pVo74Aftv7VO0AeTajPpVw
goOPgjKr/woHUcjm50Ie4O/5i2TdS+JGVhq1DokkNjdySdIFA1tWy+pfjQLLNkPa
DlGh85zEuZDlLYWGxmWpTsqrkpkcMZoDEKLtV6drSUvDb4kB4StKIWDB3ufaVf08
7V9k4Gkz0AVu/e4pqgfsXgaEQM7DcGKjSz/S+yCINXGsMnDzE8EbHBLaQch4RTK6
wTqHOpgltmAWHpvy5k4qcwtJyBmkCI5I5JFhREQScApbERHyi4RICUBjRz/mB6y7
x6dA2ySFEV2MnUST8FlXtYkIewffx5yPVylW11k9qB8PeZTC+82rAEQ3oF62qAUv
VqS2ODcbOnpeEeGP0dwkbQMH6+cVI70r+q+CK/+z8hJi8qmTG56odDpdw99baLlP
dikmw47j+ovOuI4TI1UQyzUF8bFwQzuWkLlsigYgUrilNRN+MUO7VcoxwhkeNeM/
SSaHzpg/GBhlLAdB9BFNVG7/KRmLwS1MfaoPImtxmYump5dKszs0t8dDBS2loT5S
WW1XPYIScid+cFlSi3OPoHq7rq4CmAZ8u66t1Kj0Hz3KbKVeAbXjQeat+i26GVKc
0KDvLoDqs72myUe7OoZKp7XVRi5GhAdr1TXwyXNP3IKDrJnK82bz22D2a1wQLFUq
VXarNvcDObK5+RWWSFIlAb+wTDlgVFXUqCWQeB4ghZvtCxUcdCXHhX8/vDSoB6cP
aEWaTimMGJlqcCpq25TjYPNgMwzZQ+TNdmEoJEhN4QWgXnOzjWubd7lvl1gedsRr
M+jyLceNo9HtZSFFTKOsGYyGHMNKL/sBc0y6Eq9PEBuRuc+Qm1tpBRBLxXo3KZfg
YtKFwwdkHoYitBuoNehwQqZw2tw/jbYy1TjfDfCaE7C15imX5Ur+x7rtxmi5PF7/
jM+4LM7eII10iiohd9cObh1LcCadZAU65FpdLIzrS8RpkflKg1T5UbtP4lXLOA+t
MnNjW6lHYe1IchRb6TnepvrgdzhJqnyafli1QY+RawfZKDbkC6x3OjF444D9QyAl
AGYV9JJMGEY9J3MqMhw491GiZ2YQfL+70etWFNnIlvMQMii2JwrlpLZMpqqICkcV
EsEA4Jto2gJatesnFCLRU0ger8i6bq5qzeV0J4kbGGgG1W3A+nPp521nVm1klAbn
0K4KrTfMnuQW8FCGaDPHkgNku9Y2VonAvqEbg8E7VYvmNcUoESZ5F3ukaM/iIHXg
hBoujYUya2coXhq3tqsFo5zux0LQjbHTSz7AQXIjU4Kd2ZDfKlo7Plx5xz1qSSWX
3+cjeBhN3NDKnGa8OaIljaCZTlAaWM5GTClXVJ+HfVcyOPd7J+RYMBfsopW7FLuT
2/OD8kjtKXoZnqsOj5filo+L09nUV69GmquGWi4fvDU0rsW2yVjpUAsNWV7QjB7x
nZNZYYj5z9LEY7AgxwLVb8jWYStT1Ic0aDQSDJxXqmLXqcpB041+EVbMVXsMlRwr
ofU15nZKq23Bt2S81Ka2Kq2EAsIwpLze6EAk4n7T3IwSnTXA4YEGyRJ4f6CMwL0K
0Rzr128/8MfWTwbLV1dXMU4tdxR8mLyS88cQX+UgA717Xx8CwLdTNvJvSkIW9Jns
BxYfPz18nvqKGqC+avVyir3Nxd6htHie9YKdodAPhdzkGvnr0HmQr9RSw+3FbiLe
K/wK4pk4CmAC+IHFnJ6mYm14rWNlmlEgnhegpTe6JZ9vzI+84n22t6Zqv9PjRB0z
0Dmf04759V8JQCLQWr2vKfKxlZgb3dpENpnMHXOtQB7Fx5V/4F2gK6i+fjn8u17K
mQx35Z0S4WkiuOtDcvAxqX/Q2G9WujZnvYxfiAtYXnByP79KCZ1UgQXjPCzbSLxf
jF1fPwndqBbfhtwoiwT86IzSAO1EfEAEblckbOqZkXSQKsTpc4M4kBhiWf9DNU/b
mq2lAyG44WpufZ40l3AIwlzwdbx4I0iUBFODtwqvMetVcKbJBfO7SwrRTThPnia+
PKqYgBW18zaORM4BJUu8w4kfTwEl1j5msnKh3qciObNqswEfwZr77/qpwhxB3aGI
XHrUYLt154URcWJpbDkwsLLbAmHppIBuT9GYtU+5mzSZAJLE8+gLg5L1WrC8vvJJ
qJ4IY6cx38iclmOWkUaOYRwsKAu93nuokkSpb8HRW0yu5ApnqMMNwPmWgeQcn+3f
a8BR6qEgwZsDMwGYjS00HivErnU5cTbInkfCSabf1JB7X6sr+iuZfURHKa+QV0wB
Rk17HO28UDeumg3VfZ+SGQQ6imIQtQbkgYMHDQWrIYpAcUvjag1G/qJnrOdyR20h
OiJaS6I+dxy8++LTCY5aqAdtCL1t1KMzokN182Dqffhctk+NEBHxlDQUwzPeSnlP
QFIwHZ5Et+8GAWy+ANOJkKF/jt9M9y6HKhGuL2FsEOu7oLzQ8wSdGadw/PD2MhT1
XDlbFFFnsN+7u61/rYETtNcP54pr2B5QAkBA068D16h17MTbAYuhYsEVuMbQQQoh
/hiSgeLXVnduS3bKQ+ZEGOi0s4yOrCNKcF7JRo5JzRIl8ZJ46ndLwhlMyL4XwJ/q
WUL+xBPO0YRgJVvnU8XvgATVFHvGOgjPF6jU4eAzo+cZ30nH38RZc7tpEuvbH5dY
UK2QhoVJDCJv5aFrFXtzeEXepBW4KG3gckKsfNYlACs2v+JYPb8gkaKJ/0RZ0ZbF
2mMmHjeWwxj7BhP0puoW+huMPfCdAe6oLFeTvTwoTpyYalAGuTx10HxVLhTswu3P
DALao9nQMP/EKQSfiVwRB972VvpuX62Ef4XqAa46+KkwKP2oJYv5WvjYE535k+SG
XoJXaXJlA/Qmdy/ogoBld1u6kq1vYAC8b9olUjHucYAzTfwOQKQAuA2Jl7mG0Yk9
CTQecdsF/SPkgZuKqSEiZp7RpQt4blbesoZ+zKZm+LiomYEXEiZ0U8jm6U9oEhQW
0TacKhwGFo3MzjTYlnMpW/KZQwHVmUxcAtDQXMCsJO8/AEEn8TV1ycG6Kh5ponEL
m/iomgds0tDBMFWOYbDQ8cVMJ2T+DeQdc+M80ILxGcs7H5BC1TviinNWCtZiQQqZ
KVMWOgZ3N9MZAYJ80nATaobXAATEfoev6mLMLJLMLJ9kcK6+u/ivcF5apmVFY3uP
oTYq66rX/+tDvzfTgRPCCO44zzMoNUrnhfTajKTwwLowouT2kJqI5N0RhkPap6v4
oKXkd3h3BPjcROGD5q0bg1mn52X6pbq46fzmsxQ3Qd1zz9p04u1VN3vocYKox5lL
i9jPDUj3N2qiQQ6IR7h/5u2ALs2C5ETrCniGLGQZ0muDS7ZClqFX9vIDn9NM6tlX
HQWn6vuHet3Oq3qSizJUFF/LZrpQkyjUhYxx/xzfysjSs9A7omlWjlEQ3EA3jwyX
lmCq5uY2sFLEyf7Cnq2xEFy95imEq7Gu0cW1mu4QTbpYAZ1kbiW/eofM+GgDRqIr
+eRYNGdVhXt7URUxe4+XDdW8JzSwJqfZaKXzCL8CRXW93qmgfDwEHxHiviJ4pknu
CEnl1fzBLtEExudFMe5SzLS1vI9Yn/p7C0PCZx0rmNwiWgXWWG64Jgcu0BDNxhfo
GBJgk0t2+ZHbkag7YxLkT+g3Fc/hhCgOxjrXgmGkv0yxGm7j6TjQr9/lTtDDTAy6
jnhrmfhIA7i7nIY3gb5SFauCFT9gATrp3CkUp/nPn4wNx62qED51K/GtnSjkwwqS
4ChWzjYdfB8CkiUnh6gxWlMHLrH6B7viHjWtae1RczDtEWjDNo/9Knb3ICO0do1/
DRhcNZhBCowaym4vtB0qnQz96DEq1RHGPXEJefNgFDJoMIWBYQ9GdMmDwC//i3Nm
KDv+2xpCzCMVEwGQOe1XTB3YGV/fNzn4rCmC+m12Qk247Mth6JxJmcbwZPI15NN2
qYK68LZlMxM6Z8+lcf0nIKCo6B8UdjOQFTTTVCmXCBmYfm03oJBu7qtvzwXnC7bA
pHB9ilFPLHNbjVu8pBZMC1xUv9Y5QPW7Gr1JAAtwLPmoRRjfy1u7rtTmx3FN+J+8
fBwtV8Bi92650biRbRubLISW8VzwCbaZbIo5YkVXScJn1tSM5s5Yu5dSe6DhnnzQ
utajUUTjhq3lc1KpIWr92AKR2Z4tNHkWKxIyoUcxw+AADAKMYgmVEZ+HEWbgCNbZ
Z1mhJ3EokVvMgmpszF/fMtBh0zqM3WXzRn28tDyZAn5DngxU2Fx4dx2l7zyd63Ub
NviiymnUT03cLq2aAbbtTk4UxlpsEhYIsTEZF4/7evz/hHyc/82DeByqJd0wcXsA
GL0P+OWhDs8oaUBOdzPLrtCo1xjp5hMrDCg+0/KPF4SwSeyuFNl4CrB2oAEflNoi
3jBtbmoFGAL03Hfin0eIhc6PpDSG8PFPBxCPWu6lTnMXNU8wwqelenu7J+Gz4otE
RusWtDrz8fS3xThnUSihlMdavqFQ5cTJkxWve4drYXDhDe3uzyQKN0kHbQC70KnV
OOQRFbv5oYuQsu6SNwOQRZQ1SSYt4qauNu6LGhz1/HSxZrP8uMOriq+1BVn5T1ML
+2AuLSGOVvhlwRKGrHzeZ38nNowymqXaBnmzJqTGhG41rmHRtZYT/X5UECuG4uWu
h3TB0SQrKWlIWeZZsGopJlONZTXqcQpgY3GRzWoNAAaHoxEx8wU4+7jrqS+mUXzN
yaZeXJBSZL+qWVemoA+KIhWJL+fV2QyuPb5DqzzDUBhm7C4nlGoxJj3yVE+THBeK
WBHFHLGW+Mqwsra8xF7K87SqQoFfZchYT44Tq4SPyOBYbH8cehRgeB2rMgfwHgLO
IGTVrqAtB4bF44+LMBOTy5MtJNwrMbnIQWi1NnLJZTcYNODQUcgVrl1Galgko6NU
kXjHUkHeTzu2rTi4I0rvGVTQB4Q4K1iXC9mhf+LfwQwkpbqse1YvJpOuHXYNYEF+
84ThL0TrhxjROhzs0Fu9t02MmhDZVrcipVkPgOos3Mn+tTSm4DV1/kHyg4/WtWV5
m9E2QVBCqa7aD2HZrtD/LO8d5Oc+b/4UKK06M+UPcoetU0+ryTxJn5mdoBydl9wR
M50WPWKr5rcl1v92rDOl1p28L2gxBoalyf9AglwGI6cRj/A2yE8ylXXyX5u0jA9Q
jhoxUZZY9b9PZczopzA+UpNUcp2uUUbnrMnLQ5x4gt0XNqc3M0fSRFVueoZKV2oZ
wYSbLdof9GR6cvttvcLbiTsUVrjNfpq8pzjtY0LvUUfxiBDPZTVWURzv8etJQQmB
jZ05oQg15Abdh1L+nw+EMvoXtw9eE8wJSW+CitfbXkRRZLqsjFGQvzCXRuwcriRC
nh7Xj8zlgqIiSAj1SZKVM1ka4CVyRO5tgdHTmTeXD5y7MXaXOj9mCIlKX2Jpb94I
FjwESIJQ0kdnIeq8oAMq4BOOzmVmURAULZ5S3BZBaErxwyXFPEUgmiDc2D6I6Txo
WzemTJj+ajcAhgS+DMP3m4uT6cOhFKMAA9VEJw/o3FuhbSpF3QdiMu/pvJ5+URUv
/RPv4HkSRNH0v7MJPtaFBfNAZPAQRmkytwwSX/5qzopnV28hzs1Jet4txvkz3R3p
XNab8ampO7xVqbp2Gnzs/8Kq/MwdYYQ9jlOfG9oJvP6B3i19BXaeiHfplJwfSw/E
497OGRV7XPx+4XbcWY6O3vZbcFkG7rcq0xpNp1cLOK+hayPxQEvP9YZYp+sG09t7
IU3coFqrRtfYcfrv+imJiqaVhExn6KZ7rAYL0Wa+0wIqG+IwS/N4a6DzUwb4TQog
lMUDiu89LyJQN44SCQEpBcGHDzQuM3nkKtlqFZ2ipyKX5UC5e26hSn7Vj45ckWPJ
nOmhB+Jy3RqDBD+13mF50caT9bu6vAAWWrowDmayp2yZQ9tZGvhRcpYOtyGTtAnW
KUr/4jqCtxz5os5Xjlv7HeIaIE453CwWjzsTx8hlcbzLXDU7wgeiQb89OHVyd2No
UKSE7E6z7elK76MCNN2IoYkEUZy6Z2hKaho6IrjxFhgwOo1h3BOX4Hi/xQgLusAy
yLJQ7pGZ6fmkDDodFKqmlHHpVtTkM86CX8OIKEzT916J31JModkUYgVaN/9DfDuS
mf/frcmUIU2GpKNiXWkGqNYkKYOg9tLyXiTKIX/M0ScGxq3x0WYh8APFzL6opPln
v++XtXTYisB6GYZLxM69UH8UN5e3ooyiA4cx90uvUsSDHvCFDcAYwoGkuZp/SZGb
y7clBMFNzVch0xHIp5pqv7Pvy3UC7NXiYPjNF2p3PJrdXRUukmnf4WRmrtJzNXnJ
OpnAQu5+ndanDh26IO5Pxax6A5RkClOE7ixDToO4ERak2ROhNUQd2HY9bDLPS8FT
TYbfCAIuFgr/KKdYaP6EOSWke6XG2s/n4wNUSnqDc5z1r9IX1YQKmCbMQeOZU9Dh
135dYNOsrl20ZWDyRkXZ1AFRVsAlWD99VwEug4jVs0qsiOfgzwLa8OlRhoeJkxRa
awP7RMxiaD53mpM6q3Ah24GsDvuFQbA4n3R+HINsCXCK47AGsgkGXR3sjmTbnjfZ
+n6tuMtQzq5ykNEEdpMQdk87ZU5UfrN4wkCAlUrz3Dq2HDGXZwQXu632PtEbfy+x
UFG1TcTA4H2Bd5NwUBMM/aT23NsIKHfOxd6YMh2XnQpFR3k/k1ImJ8r7twQqG5Eq
Fy1Jl1krlCDogQ2xQ14w4/M2vxZcfUyxU4GcKKiPIXuDiDIN62vfWvpGuKZo0IBk
e80cKl3c/o2d2Vo1npOTwpcZUMv8geegEAiKn0fDOCyAEn4WdzrFT45SCESrnXe9
TuIDv0rKJhEmrv6llXyj50tL4aPyt7/yVnBcVHr3gHLUTE/mj+UU5tMygMaqUbUB
n1tvMdaA24d+1ZET8CVi9EwvArQ01zQaMMsB8POkrW70GXKHMBdiRq2L1T/Vrrqv
t+hMAJZ0eWxA/YRsi8ZNpwBVlt9Hu/q9h4VJjF2USPHJ63EkaieTjxhp7w84YcLe
FSs2X1G4zYGYk3Zb7ghiPzVbYaU7httsNoJqUDnvv30naGbPEDHZ4A03vwqivpYh
V/yTPNpL+VhIJ3p5XXAIgB6zW8ImqA9MUs3GGsJ5MO90XDEsd+9FqqrjfvnHKqLp
4RNlV4BlPtfSB9u59tKBXmcVr1WnG3vFMLzcRQYTcZPqv5xZ8la7FDA8EFZRC9Us
pdrROP6xEGDIbe+ykC+Ln4msSwdKIa20VTaNlANVRKeR2DAVCwPij40o8t1fU1rm
hkHyLLpBJZQRwlaE3OLkmF1cBdlQ/TkpOs3i0OGqsL0yE75EH7B/Vu0hKRh9u/aR
nzD3ipaclmgpQaQYTaByOUfrvO+e5mB5WR6NeOQNVoR844jNASjLjnF76gioBkpu
knKZGXVcPQttYtgzFNTNUIX6ZSU0R/mX9OsMCMdFfXNYtxqHQ08FvNmJ7jRtvL/7
vF2fhASzGKCQ0oiIDOtS7SDWFoM0r/H1v5CuAZzpQP8xRUJ2cXf27YkwTSYbscQM
6dHzzoaneAvoHO8317Eale2z9f7bi3w/PfnlioRYkGK3Y9w5G5jSLSfCqW6dn99I
ysS6RvJ4neFRThPSJiMWUvF8fKOYt6aqCGzdYmVenM+ZleSt/8rHH8d5UUpkbL9Z
CnnoX2X3ra5DIWMNcDjAK/VgPY8/HKq3KUM3RjT4EAqRANiwnlB+/IhYQeXTFPnR
XQNQEjzfB/4Ghd4qsSIUXEsYUhbISHTm8X2KedLDyt+JTQfB07BT64Itt9yZKePf
SV2/KyV+QtznjZ8vyYReZ8rq1qt1xIGxxSFccXYUH/+6f6HzBeUs08f+i7IJI4K4
omSrWHQi8tRmN7oeMtBXiFPAUMTElpbXDVDDJAZ645YgXFf5CYbhhBxD95wezKcg
igkFTlt4zObxVqIdDB8Zu1Opx3V+aaoDl1HwI+sW+EsnNKhkR+NNzIK+/WPMJ6Yg
R21B1fs546pXe2JcWSKCJ9mvXM1mgabBXfw7G9by7ZV1W8hjLCraxrRPCt2aFdi+
F26AGexX2YCllZR1yf1aYgvAu927UFydbmSaAMFdwnOeAKlyN+SsSM1iJOmZvSgf
iNL2ZHEhs966XxT+sJwM7I5WQUZ2V87busDRGEFHvqcYzA+9iDSZwDhBoPR6mw9+
ubkP3YY+VCHjqiCdbAMyeQak9q38rR/4A9RRIG04z7GadNX1M/WStVsN6Kw84z22
TngWzr3Fjf+39KmaqnE6zOZzcdhyJu9Cti90w4TjxuaWoPrgiA9c0/ExCjUxmLw7
dvGa6YOSivdTpsA5/RSAvg7gcnTS7ig9Adm5TKc7nCmy3wyFq2c/KOuJ5qaY1Rco
iisl9m93Ltbi7y3aKn0261Es6cuvl7xs2i8d0SkXxHoVzwhO/R3vTNhR64Lzagq5
Tp0HOECKNVhUBjlvzNTSu678XpC+RMtdiPkJBG2CVvF1SdxE9PolGhXp2vSF5XbL
AFssw12Nrp51JP2ZLdhMupbF1JsAImEzj2hSx+sjiQ5UjG22rqLcGfB+XJbEgx9J
JiQhLZYmrVx6T3rmnM8B1JSD7EKDKho8bgBDM91LJfXhm2PY1T7beP3TgXLI/WDl
Rj25e9fERun72PlczkaSAxf00YF+T53+Mn8Kn3mfkL3YaU5PDEdbvmPd8C/eT3DW
8/y9yf8T+ZBTHq30LnUiAQ/JRki50F9KF9abBHwKT1Lq0QOKtPpthV8AM6Lty4AC
WmPUgD7nBz/UJCFsuwzP5U6w+3OY5cXL9Fx5J6m5aavxuynsIUQ7XyTUY2RDnR+t
mMiYQpTpTUhxfpPVD7ON0K/nE36ytHfzQpX6GTu3DERIC7UnBY+/lVMvhNbf3XZX
Z1LuXSggTHd5HfT4OT0YsUl/v2LrSl2mAYH7QCsQeIf74WHWb93BG8reBLtCJFtx
QKHrn3UAv2lIkwbgpkgH3Gam/sEF6KIeEJ623wEQFNAhQ5ii9ApEzAkZvDh+svAh
ugLH2f8HLz0amoIRQ3ER/eYfZ/OsKYm80QTN0r7Exha9r2OubTp+rigMcnKzbJTr
0FOylyqTHVkPSVaTl6Z4koZFlOst1+QL/areLcmfaePnp9jNj9P6rLhtPT18Pne6
5sDafdVCaVIdmr9ERLmqHMFr58wQRvb7hP+3vdbnDQD21sacnvdH60QGpLijc3HE
Ze6Iu5Wtd3cOKmURVBr4P8wui+XeeKN8Tx/oXquWRSiCz5NmgkEZbIWykmxBgkK5
/8WONcDV/0Utq0QmLvT1mPf2I4tUzPab/8XD0ZFMVmZma7nMhmrxYLeqJyGtSNVf
KO9xZEsSC1JWVjAQd5KY+Ve/ctxe07kr7OjtpmTm1CHNUQ6hMRXDwGTTlFzUaPQj
4BhBGF+AKHLHt1s230cGR+BS5QKVbtyxd3ZT+uotIbyFXB54Htjlv48tl8gz2EGV
KWmqrDZQAqlYanetaUmJZBwdDVacJiV0tA8J5EeTcaIIMmkDgLXzK8jcSOqNBPyK
cdyJKudCJl2giQrzkHfGQThSwx5PD7iPUswM7NBKakKL8030wfrx03iCXUD895Gi
RvdO+NrvScOc0WZrUP80iHbyr9KoBZsfXdmtJFoXWHB6Ejh3joK58RsdMM6fyOOM
r4DlNMOHDUOD4whdHPhHavXPJjSxDWlHQwYU4vW3czOazQsQEiyqJbCO1tdRmnSP
SoWITCK41ZTuFyJg4uSPlqHDm35Mx0cy5+qu6slV/QFYONKgEZo1yid39F3cAq2j
ZSOSEkfJ6ldt0nPEL3HhIYtA9Z/okL9ayCCChyafi2r7hnbXTls1vUH0PufVTh59
YXYDM1Z5rqqMK7rAIPKsDGbh1UOvubMbkCT1tvQAz6etztdr65xLp6D1eE/fOLzc
gztefWQnKPTohKuRF/TyDNu2Wq8MoPLu3rpf2SalQwstORuW6sBv98u4J3V4BAju
iviJGjSi0NPz+p4gAA74GxrlXSfWv+xec8gSgP1MUrdrpPjBpvcbeqzvk0EGDlPc
Ss6KGWQVrwXIgkgNS0r7XGqmIXZhbxhXbqpQ7kywJUo43KhUwS5vpy2l+NZeN6kA
YWLwVk09J+q0mV7EMQP1ZgxGMThaIZB0PQASSxhGSE8shWIuS47sgnAD94mkXvd7
lgRZSIvQvHm8qeHXurlT/+O5Z/Z++91aIF9wYmFYwqzSv7cVHJq2Komf3oAZBtEW
kGTNZ+gtxedfszAv/im8c2IeudQqzPbbtg3OoZFRYlckZN4KZLHVY93TRBIc0dXy
NTR5/wm25YRkn+T3ORRuPTTFuXwfrytM5wpoFeLu/HUAlmcR0MoGMR/a/mFSojja
uj8/UHa2Kil8JO1KVfO7LW89cMG4KkcFmiVdHNOjMra6iVQaK29R++lAcaArc5wC
AgSgxT9QiPKWp2MvOl+vgTl56pqIcYn+qpTuFqaHWNfp5fQ+0ufx5OXWb72/ViQW
4QowvOg6VlQgnoJ+fv9V+Ulz/Tjq5NbHtYLNVkQU4Hf9mWUbUES06dIa0LvwpFay
ErXuOxsC0JsiRgQNLeofTghR38qZbVjK4UBP/qU5tmeDDv0wV+v/Wd6/PWB00QdF
mkFpZ3s75eJoQ+HmdKPJoBTbQSW+ZAm8hir2APhMJsAAgL30fURJUU/PzvxTkOJl
ZpWqyMZyVV2yN1YXJXMTlQ1pjEqw07INbnJqF/mQhJnG4znlWs7A4422p/ehBoga
oESrZXMaPP47qYCUICBn2hTpxzPeS6wwN14XjT6sJNJR5oxDmTTBHl5DHdn/IPZM
3Ym6CpRqn9cxtzlCSZ024mRdi7r8jpqJzRke6tvGAnB5VX6BzihvETYsd4LePFVB
IYqSGIWekERtncSz+IpewYePEtGKqFwN6hVQuHgrNYObBGdg5dPLawVJp09dY1xO
17uPmTbbb4Bt1s0uj9G1sSxir/UlcHZ0mB9htjbfZbgi4V6djE1BX1e8ZoGVJfq6
clGN2L3xq1E61qoeyiu78qiSFt65kAKBg6edYDlfOFqkvpuvXaLf2QobQK+NVaCs
IO6J9tNxA5OYS11DtC2ZDQGz2/kUs6T9Yo2zfavjwIv4CluXN6tBw8UWcy0XcEYf
g++ydG+F4hTo0yeTkQ5Y6/0ts0CXur1wICuBzfXuDjsB6eni+g1CPT0FMbN6IB8N
mshDBt5knpR7HbEkMhNPDM+73vxJTmqKYhYHA5ijvKkepMuUN4ZlZgpBNJWHwKF7
Vk5mVuGrdYzVWttSl4JJgz8qFhUNb2ZDDMj98+dNQEtA274XMVBNmrjlQeg+6pg/
MgtPbrapgb8Xs8OtqDHxxqLkGXtUP34wBSFIegNA163lst3FihoOvyaTVEklproA
oLxguhIfMtTJ7XaFJsFfiPL2KKfPAsjDc80QG5v2DeqOV5loHsf/+GJC7YnhBZpV
rsvsbNzYQ73Q/EmOLbrQzcI4GNX680CTkRE6YrcesXh64WNZzr037NAE8Jm/9mKb
ziUnFRZlXUYEAZA3Jxp1Aj7TDIVcxMLROkCpkEFEv4GUXrLSOl54/Bbqxg9vqzYw
ptDiiqHqUK+NaIuI3xDngdLY4SQFvVD0rcwrS6Y15DWSeVQjvXkK5FK/Q3RS2NdO
804vblQra3O4O3QnkR2v/kMBpb6+k49b3V/LrVO3eFyRIDVWPsOFClqKswtC3M+i
E+IRqCpkcOaq+R4RQ2ntL7Xy95MIGCOaxbmhQdNOcULs2fuQPLC7FYR0IpCgf+gX
NgVnuMzWmUCZcTaViS7oAEuk6tByK7r36fbOJ5Nwp0cAuP+iDwUPA/vpul+Vn5Zx
pBYoxREXbOF5DW6a/04ZMptaMf6C3OpzlB0jIQlc4HcSzp9btdAOMPeHX8sf5pAc
S6jlVC8I+1RC67fjQV9D8J7jb3xLz4YcBHDvzidugatZ8jBHTumElY+FLmvNM8bx
ZWch4f/QV3SrGfpdySWNBbjKHLT9UbKD6Tsss8FEONvQXkuui/LprhyQ9KlPTE7I
XNf7SMNwp0lM9B+i1VMs6U1HcJgYNrmKKMai8rXVY8ocKKzOn4gmqzrq9Qx8CEj6
5zru1ivp7S0Kv7OE2TjBNIdi6aPhuOFISDGPZqBJEIFkZHKabRE53xpVbm4ugvn5
3EH6OUHXytNjapYxolUIBYX7O2yY72qhNLvuGJ7iFr1FmXsiLumoH9Mhub4Fv/ut
mnRxVwws+maJOEpKnapYxCeHb2BfDfXUhhn1k0gWUEQPEMxhYlyLjP3DZYkj8/Pz
7Js3blZMnicyrkiktuN6h4tWYq+uRqOX/IQCXkDDaM56uvSygdxKUNdf6PEjCpvf
RmB0raDOc2xYw1PFhnscpvsETob6f3VC4HaB4q+Na71JeJ9DUL28TKmkpG5LLvfq
uczgBqXr25MNOaDlgGqzJ4+9WJ2WvKILd1xC4fBSSw2faPEMUoZd7YLSz9iE+/Wu
zlVF/fznG88jo/cLWll/EbYZbS2WwFb3dvnMvfLEs/26Q2mdo3yC4FwRO4v8PElL
GaOfQGGCSGkQPT24sEYy3H1hABxagam1K6rVFP4oomc05qLHq3x843CXly+JCdmO
rv5gNaslGBVgnQ4kmpIdv11n+extSihbWOp2cO+nmkUvAjGR9FxAPZTXx10dZHl0
2Lw2jopI4Pl5+0gni9tgtbSng4180I8xSI/s8GhXfD6f+Xkf9G32BpQWcivdenQx
YJ8TERSK5blMHkoaFnW8HhoEe6I3oBJNe0lU4rQ7DB1Uk+lLgInRdVe5S0pKYOgr
uFyV5KvGepFrpbcKCdn4+XjDXsqWfqlXv11nYKTX7JqXk4ozIpn204DhNoy6Hvby
shRIdM2NMKjCud6SbOUB43JM8RnCK3BLGwRSNhZEWtxc1HdXPElN+Tiv1wnrlkwh
vBuyizwU/VVHj/I9ERf8RKF8Jr6knCR7FOmOIVzE6tsYizK5d5MXWzDUlBfu4MIU
NsF4Cmbux5KrjrwRyD2QbPw42OokR8F6Eb5oRCA5KjNNOPlxOCmw9sAbke8VsKIe
gPBJh1eabB3izbNtMjI0vUMsjdg6I3S6P6nAxOVglVYaYeZ+k0X20Ed6lvjHz+QM
oXY70AGIIOHp9x3M31s5+mp4SyTRrHozgOL4IzgSJ6z6ly5FrBExn2mXvuZarmAu
SPiwXHF/uXgtBzD2U6L9VnO/tBlnJMfnmggM7uIc4P3uOFxiZvGMEzktzkWPwW7b
tx+CEqP/SdqaMQ0VtT8u4CLsuk1aoK90XvBYglzj3xmihFPTgBJLb6K35PZyNi85
4X2g6fQksFU55rqpVFNAUJCI2/xA31Bxpu6uERQyvoW8U22ZmC7ngFgD/679FMuE
LFupOfYpHJpIrMcactGVf6Lscg9dLB2RHGvfCGSTAWD7h+bLX0PKE0mPjt7fe2HX
YlOgHVm4Fs3ceYfSVkmN9c4K1EO+8QPo6eK0iohYnEvNYXQ1JVResLRlr9jUbCJ8
woI2jsHfcj/JYKzUubO05+D4zv8Eu6cF5vRlXXx3lTtSSmzUjd0A8zwBUiqwL952
fgFQn3WsIxH0kIArqWq73/ee56sbnqLZOHNdtLS0unk00+JoFkDuaJSVJXePoM35
d5GzHO00N5PYpgzlUek8b8RZPdaZWLJCaolHmFYNGIfZ6egiqazx8MgNjBtfCnDO
KocSMqkBUzwoCr0GDglFvo5fNcUARi/kK6w/TAOYYopKxpEow7FU9Mp7VykYpcye
qc0R3q5KEr+dDMl+Ze/L5QOO9wRYwNxot/MdnUkGP5ICKhz9IiWz1jbCJhbroB5u
lOMBlMGAq7hI2cB12oP87QYLi4WdKNrh4DUiRjqUdZ4JzGIBGd5/oqqCo6cnXelv
t+Nuz9XUG3tpoN4leMOuOPgxqMrtw0uooW9LpmztVfRcZqdc4l2bwpcYjqalDsIY
xfYM6FgHNO1n3D0qq9/R3vyqF2KJurEcdH2qj4Zy5LdGNOHfbGDfolHk4OuQVUK2
4bler1VT/tr+vmUkpdF9fhl7fbvf7bSGolExwD1s/SZnm7kXrUbQhNutBQCEZhsb
An0z9OU+616E9/w3au/HjVpgifvYYVW4SLRhgjLgUAlMxhvZmeypCIXO0Si28IuL
Cu46BYOm8RE1LTCJGDEveStoY1r+NAJ69dOfp/L0o8T200gtJgI7vTimtQRcumvn
YA05X9XnpW8DrBJaXrTTn2ZHwHGtnk7+ILSqo0/SP1lvg4Qas5U3yTEWUdkgl0Y5
lLSebaKq85Hjv4sXyOmNdV/30JX5ZJwD6h1qgkaegZ/IP6LLkxkTtPNZnN7swmNM
PGTcjj2Jy6jizqLHss2LfBHFyETML07slIuPyFjbVAJtU9jdcxPqmnpH5BrqoKqq
wlQ/A9TfV+4skR5CippcKCBykIC1arf52H75+ePZhX42PKSDd/VT6ti+pikn7JNp
tZyb1N2BhAuvBXSvODYPdLLVL03zbzSlVFsRaa/PEwS0Ib936TbyP/kcyttyu0+m
iTFDXjRXday1fIVXoziX+MaQD6cjY1PMcWRdrkGiL3To3V6UOTff4OXkkG4U+vzG
94+CVsUVKn34quGhF1CYOHxiy8wAMQ7kR4x0AYPBQM3ORx6NoeVDEFdjTn25Y4oa
/nC4kWN/rLBXnZ2517N0A1jlUrYcIZZ84Yuphn38FfyZ575+oq/6F6DjHUowNEr/
5w72sKoirLDFyqGXu58evtO91BqpdpHYg5P7OCdhk9M9loSkFsj5kV2MGZmLMaSS
VZH32RZnmqlv+2SwvyY9GzOguLYiF6gUcMtnoptN20prkq8kYCj3FBZcEoGmQAtE
fyNmbRlQ7dbJGggB1B9N89mNkqnZ5vItWV/iHLkHNLC1qTjVNANdtylc4o2ff0Qx
FYaPaF6Fj7yKycdMhh9liD98KqnIGHE/oYPSlwI830b5edvLzcgqBUzKMm3Cnns1
1gBoD2dhVL1XR5AJF6ytiWv5D5uOYpz0TKHeQRIzq3VVW2mu91CFPdAZyjQNIoD2
7O80RIiIuxeDFLeEMtRX9s43Ws3tLp0JLxho4w3+PqLQenX4cKORwte4BZZ6Gu94
SZOEt6CBUwn3XhwCjJ/c3vAXGvxqeKZVeHd5UTlLHEZZVlQw0l38OPEHBDmEsbMq
79L/VlwmoYZOfmb/513565jaTh1Dey4Lc14TULllfHaU/6gFvAl8q7M66Rl7/4bd
ChxDMvhEUCjrcFrPrqrmuHst9Fv+PmB8E+lcvTQt0XmUM/D+yX0fE1yZTK6agbtG
z9jWJF9JnX2OHAmrgi+oX2+fPn6auA19wi/3ccXo/giIewAOHbrFNQhJD4PxIaCq
v8sgINfvFBypLU0fdN64IF8/NHzUGZRrBZtiEr9BJk92MlncfwXe+CbLm8jq3BLq
oTDfTHOxYPSk1eyXJYiS5AImMkicKtkc58dIGed60NoT4m+N5+32llpVSts00MlZ
vGZcT4h1NXCKE90B1UZhE9KBrLMwrSFcE/sPrJ2Jtf7/cj1FW4Yl1locacQP2EYG
ifQQZ2t1EotejB16nr+Sj47kkjHzoOq3m6usXxuU9Eh6xDkQaLEfLYF/8a88ydeO
WyobCV/XMMII4sBYr9idKKY7QtHaNN8H2qugtspjq5dd+ZP9r0rBEO7TNcPBoMBQ
Jt5KSb/v8jspj3xmgSm1Wj5Mik7U4ukUT0lrwyDgMNhO8U81QZVc4tVWnSU6nDq6
F43hJcxwLbUCLGo6YYZf8t6kbgAjCLsvuH+b/ESOV1LEXaSFgagyO9TIT8aqYt0w
uMwl8lcTEbMGtzPLacREOAG6w+StISSqGyBltGyT7naBUvkFPlSkfgpLihksKiWR
2+PNZmOIOVS/yptWWoVc/umAj29phUbC+A9mMtFtfANlC3OC7XUiL4PFs4sr2rm/
Qji/8kOGoVVJtmLw+7DofGQPw2bmJdK8Ud2ZX5iFK0C+rAIb4nXmvu/Mr42kem7/
0rYPaCUR2y+17jnijNbzsuj+cwu7cKr0GdVLCKpeXNIr+NackMBjEold4R4ncfem
d/r6J5CTFOVukjp8LqJX4lgkfcLxw2vvWS9pP2v9E4IY+YuGxYnYRJgRjvHZAHMn
NsCi2lUrWBvm8Nty8tZkAuTxi++8AR7G3Cq1/iAer4bj0BYAWlQPnLchE0zwhWjH
9FbHGoFihEVxj00fTAXzRawYxCpWS2+wZIyuGB7ySFWF3+W1g6VoIqdTkFwNR9d6
/WooKMOcVNs9ek9T6QyAEy2++xcz1lL3CrxEQRogtvMXkiHHz/9k4zfzAkJrgSTY
zOvSRtKdg6Isl6DCNTQFLYuzHjAjrBW3HR8yQa7cNglFLtu14nJN+Gl5km/DTaFs
NIRx/Py0EHX/yAtngsgIknHpMT6f9sMR9h4a2VpKaTPyVKAyp+58wdXuRX6HUwGI
3QVQ0/45k3Lo0a9ImZtdcLkvOSKUpptGruW+J3eMeMUPT3tEC8oOfel8BChnidpJ
1WD7WWBf4VeaIsICRbhx7uXfbXEtT3YZzKfsND9hAfOpdZQ2VOKrssJaTs7kJipx
cCNgQl81qw3PbQ6xA5OeFErwE1w4csI24ABGCrx0nURR9SqW/d8na1teV0YpOsZn
gLASRDv+znAJU156dBGmwMVIS7B52C2JEHttrasDHwu89iFz9MHXw9lVvQexufQx
Paw+Bo9kRY40bc2dBGWilBf2RYS5SoyAPNhLuFCc14KFDurEUc50E5GEkZaQKAr3
UZ9EznBfecsYBECJSzswhbd1m+/pNcskNgByLOnNeK1/YoCXQ9BIRoA/VU2e1R0B
Qv+b6vyWIVlBZjEoX7xODenYOUoNlAN/9Oxb+Cp9SHKGd4QICKyUZdEtUdLNvjhi
n/bbhg+LmKjcCVd9JMYU0pO8HvxiXGWhT09Fi6pmeX4lkBrBPsiGiD7e7FYyUldH
3bOwbf3SaNF8jPHDRWZWrUW0a19WfVQOOvvMCTGNi4ItEcZOeeqcklEM+Hqmk9h7
yVDKg+1CQPSQgW4Zt3lkvDoJUU841T1jqE6hIDjis2EZgm+61qWhh+JcwPks1dhz
Ii6apL/iWu07TN1CLG8JF5iY0f53+/i8vvQqIS5WRYrV7g9WhpH7jVF6fJ2Vbh2U
IWCpkWnfuXnpWKmt94ItLtjELiiqOMdb/6eLf7D7a7EmpoBljRavj9zNOX0+/kZW
KRVehVqwvAeCjZqxSNW4fSap97aAZYG4CeibTMg9w/WlNzYFOJ2OVMskso8COpHW
2UJjZ7pkgCqVZw8ViKC9EXKDGjrR1ZrHUcBGn14bC8IS9xGCdlHq7TBip9ye/Kfh
xWwttVXYM79K4DCAmaKYoSi0kVxvqI49ylZbPFFob+pv7BR1ijBJ9U7eUDq6EC0f
LGS5D5NstXNYmXtHS08NsKdKrzwzSoagGdarNl2h36xd8ywCJSLoutqAw0W03Ntt
GjoqcTvMFdDr/SQ5QQklMIXtsMq4JzZjSq87/+uiT0UaZaU6rYIXDvNRDM1VHiaI
wgF4sH0Arrd8xoG2g+QXw7AjL1NVGe+PrUP6GdKrS2A/UKrlL0aM5+OqW2UMr1kD
hkLl0D4coJpsXkyNnDMxVVK9GtosOB9PGfrDAn6WR/ROK6PtDJUbDQQegFE8YHrH
DHyemNQqtiM9CQjrXJ7/szdygug9tvQHGALszZ9YChPG+J5tRwTRlpWZmS6Itb1t
MOo+2zerMbw2fF05fCn0kOPCJh5PQWetBiHsuG4/evb0r4f9HSBg8CkDuosKzGfI
kg/Ut7XnI0bpQzBBpfdzuwZyl0JIDwi2JKNVY4F+IhuyrLdNH/7dAWeOIHOe9dxO
ICLOsKF7gSYx67CNwGdjzWwyyPzZ5n6Sy+N/Zw1xpduygbohB807/Glgyhsq4JwW
bwBIxysczEgh/bvWjndBe6rW1ioOpA54OWIOKOFQ8qY2IlPDLQTnjCFpNwIoujNy
zLazlwqf7TxNmyx8iZ1X9NgdYC6v1Hj/BRdjJaVaY5M9V/EoO2lfN+dZH7HqWK01
OCX02l99HfUlOEQA5dfyQP6jSgnHsQnsHVknN+V1WDrYaxoqwez6ZQaEg0sMIpna
9D68Z9b8f0+PDR+OIxo6FAX1/Wb4FAwVdMpb4ptxF9B07wT+u70HQ8RYDobbPZV5
QTacAKR8dbJMC7res8WpD+xWp/VXzRB0ZcGx9KOBWcOKdHkEZ9Wyis5ignL4fR2b
XVmQLlqa3gwo+itnp4mkPh5qHwK1mSt9dVGEqZbrBUTQVkS9BQGX/B1ZqlJf8uGK
JSfx+g5PzFg5pSt1hbtcQFGUD201RIysceCZbeRd0SvVCXJyAtXA9RVmMsutBIb8
JxLuWVfx04h7kvjAkw9jnRX82I4Fm15X6F3NSEeQQ5Mn7dqcBFeF5ebSrUaGpUUO
r3xkix6SihOpI9MeNgHcJab6C2hCd6GHyjpzSBv95Z7pAPeDdsuLwMUCxa+qctVM
c/eMBK6brTEdwYrGUXxTPQ6zxJkQepkkKclfaq1ZhQ5XFqPUF7eNK1OQ95uk7S9E
oTerKwSSdX88TjECCACwbBl7siiWlYmgtQKAwyDXz2rzlg3v4IKi/KFUjJsMFdeJ
7s3ehqXQ8FNFw+j719Be6oSrHvi58ueiIt/w8YbFyps7UOoY/kmwJVudjL/xemr2
6vPcmitmP9h3n13z6kS4ngovjEvSfH/GBVO+6ZAObak9d1gypAsAo8svGW2kMTqt
8VzoTT7Hpga16LfmQde15r47gAw0vlvaBJyeA2xiwgxu5AkRA20JzBBkly7Nk4DM
8s/OU924lXg0e4RDV1mBfABS1Pe7PnqiMlDZWoFFgkSby6NmctBL/PThQsaf3mth
jXMw5W1yZRuLNgky9QINK8KLxDam3IqYWBGI8fXHZdgWZDkiN0Qg4NBVMWQ9wAM7
z3SqjnumvfyOyBR5wrPAHWHUMhYfoqfS3u2K0NChMInlJC68vSNClS2t69aEdBu0
JXkk7LEZXXGAnk4xJCVJRKzRprTE+pR4AdurYpWKuPRJk+bjrxlPiEB3LpfpaX4e
/3VqEOP0rdXvvTrzTie0ZGqa5K0BoW8fpymzauOPUfBxUs1MKyGV+e31KKkBcBHO
Sjz7V6Kz4sdLpFXEIQkigHD3lq3mJY/KfSGePxAxldeJYuBfVU/6na4pu4tqe70u
EetvVJ5o3GSZU2vvq7XZJuZw1VxrEjX0PTD6AH3ja3+gQ4ezQMAJpRp9oR2dYlIF
GLq+IWTeFTVsFYJ9Umc9E07oCnTv0KeH2zhhjSytrtVhMNSU5Btl92/E8Tu9k5Yj
VLleJWUcW3YTGLhOtAVMwSCZX1XCQPq2m2jZZ2uRRW5LwyJlhyEhzTBt02PxS5JG
nBc4lZiwKrp+b59DhDYEwoJO4wQQZb+PrSogDb6S3WejPlIMdbxXwCcmOCg3NFLg
HocjDXLgZUiXSYOFfecI81SfLpkdZMvTFAEsrIv4jhAcn5CyopNbfZz8RnRAXFBH
LGSqz49NH92ZzlgLYO2HNt+4R+XFHsBfR9u+k1PI/B4fUwf7MAT1UJLACYrh31KN
dO0oK34zE0HeemCJUt8uRNF3bT5A9W7V5lA1AVN8/Wl84teWamd3fS7z6iI8sPZG
m1lkSm70NSiUhrAu6j/4AIIXrgNEKG4OJ4Cl0x4xQJvVTft16KJdEHei4Al7nH2u
9SGklCAPcC9v0X3DopcQ+Nf4W88WoNM9z1qf5KGR5SWHurSUkqA2rgIkTtQa/UKY
8bFlzEhyKFyz5ca7KPpKrF33Om2FRNMI2DdykDh3pe6FRFDRhOv466kP+F/QJx5u
BvItq2LZm8y2KoukLYWMz+rfDTs2VuAs5TyppLG4yZwjqQhvKjqQmUbc6lN7neCL
l33GNAbQJ3XYL2Yj8KgwqjxAOnKdRTDTd6qBNyOt76Kuvr7B6I2Ms0uHX7LkE0Uf
ggWaV0pbOk7faUtR1pWGqB9NUv1x8H1H0yC/445hR7ZJF1x6LPJMSEpgnPGpslAw
1jTcG5Lek1+DlgqPl96wiVBPiNuiLTztGZKpT3fk5wOS0zS+O3E64us3tAMKxgw7
lnzOjPFr05KcTJPbpeOjqGMIhBLugV/QxwcXCk9QFTUNoqrCc2zKvPnwrTTL2uJh
daF78UZsOStj1DxCs/W0x95kLWGRBRl4UZ3oGya5riP6N06DLw/PwgDMIQqQ47nx
s1W1Z0RBajD0q/NcecmKqWROwnfGYzFnHMKWx4CLuoUyZVctOjN1CC6VzvuIjt9b
jU51vS2Y1z8BFBpXAeRRo87De1LJTbJl1AqwA1HTuOWoMCVAIlJHCwZTWuh0vrDq
pM9HRiXq0b58NntwHmPTOec4xp1ZovHtOg7xHRvGO4345qyAXVjokJQUWVUn0PPG
RNopJzhJ4Zq5vvg99BPrLeLAjhYjFphWcXa7O9rBlCDp+4EB3Pew4CfQr1qSNDDI
Vun3YBtmQ2EWovkRj26EZuOCu/wXERKQS8YLeRHVvF5hsHEmclfnU+nhXof2joOa
oluKjqGVDd+gang5OpInxEwAZSheF+c+qW1+NMQNA+zYn0H0CpfSyeUt1kFBFcaV
/8Zois1Kp6H1dItVtPQhwRjo6v7CGH+Zb2ldyVeMUMXOV2p3FKbTZNbS8R4sYo8T
N5uD+H+PZ2V+ZvCc/eA+PCBbC7HXQdjlPUMorLTOEUwzH9ndejkGEEvVRt9+IoL3
vGpVjzsn5hYV35szaYQzws0COQbqXwLhSq51cF+oIBzDzJB6cMGt39sXOQWB7u+i
g2e1Kj837tIZuuKUL2xI+A558oyBfO92JGu46vYnkKbWfBmLitUfaXRRUL6c7PT3
ESUz30QTpvFK8sT7G71zxU5uOTr4XelTU8CcYNpR/LxMk74riD3dDVg0b6SJyqlx
3TcnHK3eO1CqLSMeWlOCHitK2eAcRjQ28buezVBN0LZajJDNKloPD22sykkGewzl
jzjbmQ9PpyKrh26bfg2hpfYHNogC5BIFjdp9LqXOSmuBHO8s++YSt/8lOd67L5hs
CsBHKmIlNv0xKMX7eHWa8eTVKcp+PW6ZzV9Yh3K43I/9GnnEyD7o6B+Vp8LGVYDh
NgppaHxWd+re/iP/NCzKuI5RgEvipJ20wxyllGzHsIe4QLEd+aq/ScJFESG+n5im
84z9o0dWEGuKuUodKIKkKO0XKQhaRA274MqW+zefzIfQN7q5FtecSRu+MWi1jC6p
dy0OAKPsI0Oxhlnp4RH7f5zXfI8jrqwxn+LRf6uG/pbgcHqcMYuzpLh+QiKizbQ5
PeDoXZeZd8HW9AVCoQOVc8YAp8Nf8lPt9Ae5Rr9bChpTjtoOdZaFwlrYS9vhQ5CD
l1v3CTJbwWEKHa7ph3Igv85hNqb18R8F7GHu/bPNIv0mwSAhsUUa7QRcjk74+SNQ
3OJsv/f2gSXm5djbrczEE3lyYw1smuVQPbNlTEvSUgPiGt9fOnOxcIiPKyOIwt/a
yePqEvCrClBqp40BJyK+RjWm3oQJMOH0/terfhKUCifXVqOZrbZLPiUr9WnNe8jo
6BMCvXUcYRqHUVT+hzVINHJi27LxZ4UNs8sEjtiXWMPSQgGsRfKJ1B/I4tKNdt+B
aOr5Oho5x9IZZt7BVboQA4k/vkzVopuN6/Un/iWYAbGBz9c7w8+0+xYGAhYu0ER2
pyZLXO3rQQnkM7ydgHCy2w/il2kJ9qfCSHl6ONSxv0Gf0RvOs8hWh1tb1yXXh5Wi
/AUjTGqCOhjdeq5StfuUbVOagrsQnkLiRWpc5rr4DmgStXsVBRBQeraNoRyO7zOh
kikZ1DyWgyUDnpcNyjc0m1f8zxXntAK5p7bG3N6m3ah3q0WkHWCHPLICsNyD4ptE
BKeJk3/FpP9wvKHXruMiRVmtc9z4DylZgisbLbpWZdNNcHU2//SZQbbcj+BF+lCI
8mzSZB6l2QBzQ8EnZyKPdDkSG1/8m2grp2Umq86x6h/2TDoISs1r3xG4MP8EVuUK
EiBHvEYUzHz0Q3TNneQmZWpEoL2ggmDauSy2VtU0aKB9Ujth6dOnpUKMvq1bw3jy
0E1ArXzB/jA9hJCihRCuJKQ7D+rMnJJ2XxhPOWz/k6RyhG7s+fRO2KiuyWnr1Eob
r6PMEu5JujLZPEp0j5N5nYc9C9sTu85b22h4EBkZElX8BwTuxqE2BV2kV+UAVNck
JKSg6LUgZqgmrpv2AwURdp5RfOWx+Y2nWaJXlBeC1Xg8m618kp9wavHTjttkkjMx
0pwucWtbB665MJ+pqwDjuIepeu0fdOvQHCVRbnBTKW/CKhFw1ej/I2Tx3ELkK/L1
qcK8d4wHURs55slYcUgtMWazeKPEJvcq+SJFX5PIr4nhiGHEY4zPuHonu363m1Bb
fmJcoEDjErAXxraBjxPS/fElAK7HTk1BOFMFaL5YbGT/k5B0D2WE3kz0tZolJ1CS
nL/D3JeeF8uH7flPrhvBUPfzGIJ5x/09Tgk1OitoWFTcvcUBOWECynX0NpcQFm/7
gj0/glyUN5FkwiNXBOzmlqEw/k5o8rKnooT4VSMGAR9ToFCDs8YJlaK4FE8uCVy2
otJkaLPLnj23zgHCOWOJo+PRMYqWCCiYtGIISb/UfGH9cBIC9oqjoPEshtZaX3Nq
GTT7B43pg3yx8XnQqbfcj92ETmkDGwd7IbgAPryBFzpT/UaJjGcYVqJ40tQko6MY
9QnOwPxPgwO8Uz69EUKkveJYr1t5QGdxZDNuIcFcNrxRxuP/21x0wVu+ZjSxy14H
bIBTztLN+HThUu2TClwk5SFfMMKb06En5g5MXdXtSO+eOQKt+amM1uJj1UmCWHfF
JizMVSzhWeTmLA1Sk60wNACWe7pZv38YM1vrnKCmAk4eUZJdA1Yv9oFuX6KhY6Z7
TRZhmnPD27/xi6OusZVNivO1wZhQM8+lOJ2UXzY/063yVp1Qgy0+y2fih22XCrcE
hyhU+GHE/pxg7zxKrKBrPr9jRQtYSl4Sc6SF6DTMGfq6Pe1i5wIAev9FXvVeKbnW
2L9RvdjtWMnFspxTv1XcoacgMmnsoMh8Hni0m4ryi+qRoQXA/NxPdmCP/vrm8/HX
kKn/BB6HFdWnUZSlKhar29YhhMsH54WGZm5Qhn8EBDJg6E0sg0jy6cZurMoK6/J6
sZ/QsEukOGsvvD2e5/EmFdlp7TLh70PEh2gYudPD04SA0xFRtVgD/RoPkv1kBGW3
6hS/8jSnS4iRytLyx72HN4UZQMKb6HujT2vDI56YRwj/ZAmm/S7GDfw5AcvKHHZE
xv3ZJw2cyoNs9H1oInhxjTN2fEH8XVvBy/nqr0XO/cNfwu1W+o/pzDx4A3nj8OJA
dc76kficgckhkQPTDEzFezEP/6+Zyvv9DiV72gcWC1PusicXibu/m/qcsVsWqVyZ
MwXN82Bv3ia5x6RlrawoWKG8wreyMQo6dfgcq42QrsNxDhgR9bL6/rkhnEwwteMG
/WmLMBW70F/Q5oOyjtjmzoHMButI4beSuwworZH4b4zMF+5a92rMRRusKCP2HMRA
bYjI0PsmmDm48nI7+NLqDtoxHiIRuiDpjdxFnyGWgo+L/w8Q4IlLvimD+jdzbHOE
0unEBcjmRIHl0e4D11GY1pdBHdibVTay8AXm2MFAV9HHY/Q9dlJO959ODEXhoCas
mc+hDOCzq+Z5uxGQRQiAgrigcY+uzMNXd4A3yHLhPlo+bCAwRhU3r+ypvcNct+bd
29Qr2MtXYxQG6uyIXTrbSdJlXgtyR6ZEnjlH0NxyXZlRNNY6cz0ouCAO+TvWHRf9
1M1TGmJc0lg6IRjt68+sW9+JFALBGE5RJUQq+0TqPvE4nSIX/iE2tKfLnMwNxL0B
6NgaF28hKl4jVXkjCtlcilcaOtQ1Eid7DMOFHXnSGjy2EwO08Le9H3QR8o0yVVkx
CJdbV76UyXt+f5sVFQiwEfIkqclHkRq8e0B6y3gxEEcjDEeHcp9+GC6WVSjsN69B
rkjsJRd7yzx3zkRYb91qNMPJocZjaRwoghahtBd7bT5kQ2Sr0AfBk0oE+x+AV6FY
EIudxxrHMkm74/wkzI/vJlPsbjiuWJ4LHryD4K6QYrat6E82RnKu5ESs247k0JMu
lCLCV0GC1MKxGDAck0NeDDGLA9tIs1TTiQyoVIJrfsaU9rKFITqMLgnvshyLhqQv
FUmIVM7WapibALqcR52+xNCRDT6n/kRz2WlMcleIwo3mPGaWYQE5cKCpYrE1yKjw
NI5RuGNuN3dEZgVukpfM7wxIOyzcUn8mM0knK22d4UY8hdesM7T5bYnDm4kjKNPn
DhArDWGi7JYiXzMEE2qQZoOmZ2zTyAJ2jbIBxHQP43r4jOfTo6284NfffbUFF/nt
CeEQyZ+evK1Ulj021WGKnWjHhSFnidklneA+IcXZf0n8fLxNOoZzrRAXuudrDAXK
BzRyBk5mlf3mET04SCbcnD20vaBLvPVz8MDqNVHtEfOxNkA5QbelknQCBlMT2XjR
6yc4FPxqGk31w3PGy/zqXYlM7iVAY1IL9yCopvH0N1nAHKpj3+en3UfHM7RL6JmF
R8LUNsivb9xD/u0q7MsPUMePENmkWxssIa9Y7Rxtp15Gj+hzsPTRX+dKTz1kESsi
PBkXMQyiUUl/VHRPsYqm74CtGSIShFA3HNLvI12/IaWjNPLvJC79HQpwOsney01H
J1fylNwAvDDi71chbu4Jza5k7ANi6id/uHOCFvforkNsLlDlYHfdgjf98HBz04/u
GG5reer22nusv48B2njczKC2HO6vjQkUOiOtU7y9lCe7vRiqkra8Yy7I4UKyvGmd
1W/SNN2iXbV/7EfMS/UZPwdhzPy/W0Yv3YZG2BW1n7gqrvBYCIX394rxso/Ra2+n
0zlLE3+37cOoTMmgrEfVkVVk7cfeFhASyXpdT47siwtYnf5eUPOBB3JvwiUilEuh
U6ei6hr0PgOJDaHPNCfhBP+RTC+wiqSc/o0NMGGKz88U2jZO41P5zyfxLSgjls4+
jEqyqeOqQMFaaTjpddnXZXJ4cZyhD/nBLjOrh2yPR+nP7vnOCG7+vezdqWF7IbgI
05u3a2jNl7MnYH6Rhyn+Kg/MZs4mwLmWbYEAeVEAjlrQXPyfCrHWWEuVYv148VoQ
4z9FR5wXRB7EfNiCytbx7MCYCV+RaMKhyL7jmI/BUayKUTQ10o2BjnkeYKj27JoF
eiULdD/xCBWISXyXp5bIpb82b49G51k77SU3f1gbAHYSzY9TBM4N0jmA+5Zm5C5r
FPjl9LZVaiirEb4xq7ftf4LCvvNiR7bKy+FEjVrcp4OubWI7ymFM01AJmK23ppDF
VnZUQoJixTNC+pJeswUnFHu31eRbDSUjO48t967XyqC9cXg2FNJwx7iJaVBZjM0q
3/hevFg8XmC9DBq341A1Wf8Y6ZS9wTLJ1QQ4+jcl0IFwBD3EzZ1LzlhsbSNAf8w5
e/lAmFJoLtZna7v0AkO3VcpMGDAlS0nSAUjYbkZ628oBfw0Om6k55u61UwKzX8IA
DW8aehCcMd0l6stdULTg3wbEVTIiH4mpO2syxF/HoKLrdavH8Ch1ecWq7OlF35i3
aD7mXlZPSVk3n1ccRRl5XGw2M/mROwdltUKaqr86++SA82qjZG9Quuo7J6G4U1wY
dhz92Fy8imE8TYqBXHqG5mVOJyjb3ES32OLVU9YuaiNgrB45xUkme+Ci9C7qeIjL
VR+NY5BqNBh9RG9P2cgVwMT2QdG/qcNwrct857WH7H0CsSsCxr08bCoxf1a+aMZT
Pi5bD+AZqcw1gIIJqsHznRVcRvy52O23rNcvafO+4zbcB0J1zLy0aVsru9JgLdKm
EB4CuIq2gvSjpG20awzNbZxwOfNVM2R8JewWJ6nhTTyLZyEgZDtIk9h3u4puHkTm
UfiCpBb32L57UmYUzmUQfXNWbj5RIPvdvYgCUnHNCsL1NtH4hd4bQ0YqgxrqlXKP
YbFpeBIIMYy8jEqgqxJxguWY0pbhJDle4caMlrbmBFnrm6b76zzSjvVM7G3UpU1B
YwDfqWptL4GMqnMf+jw3dym0w0OZmv3DHTI6qcZpFyx8OgAXFpx7ezq+aYMOzH1+
LesViyAM7/eBYp0t/4aDlGbLO5uQ63tSMvxiaf+Jp3hID71zuv+ULA4qRBn8oZWk
nWwz2oVmRAhxvuYRXckWRyJT/0h01eBTU/qt8cxMehCDilsmIBaU/76tiBM5FAis
kZgL+Mp85NwcKn4MalwpeBttIDeRzaIP/NljRszfRCNxKf02tZVxk1GC29+6hFIN
MEsBlFOw6Cwi+3Y2ifrIuEwBF6bVO8FnVybnFmXyb482XqFm3buySldSkN9qUKC6
rg8poBDPG6oWWRNh+QxxSACucMV8MisHFCHnDTEZnlDxjOVTEW4z2SpxXqYxW5lo
yJvxGF0xRMP+bn0h2pavs22l7b3zfretZg12aQ/iC203apFrw3jOteX/yLvkdYDI
FSUT38+2EhgcfZV0w+2fZhK8c9TVk7CorbKVzKEFjOstfpuPjoaSVOYAHtHjNZeN
s2vgMAXfLBmpPBfp+Xf2uJ25nvQ0Wm9eC091VuWnUuhr46s2pmFzmuu5t+R3iJwK
J3DduFxUdo3gdqwlC8Hg5kdapUWRgimIMAEu8TYmIM90jFEzByg8DE4iI3n5r575
ry7V635u3eFHFq9d2iOFYm+99pp80z61ISCaVZbqTGFVtuqbTvsXrfK1wsiGrNLJ
z0TwPta3ekPZEBACVetM5CCBWjLOCQ9/ss2dSoSlRzl2KwcTXTUDNiYfFBsfF5Vr
tlvedEnR1Gs85xSWMp2jYud/wdxEElM9kx46wUfoP6TvOU5dipEaT6HDqy2aH5Im
G0BM0/Z8/cdw3xnUxjskUs7AQ8FrBqFQukHkdkULh259ihVI5rMxg4tZb6jLneT1
9zo0bLCftDP4d6vp+eKf5UFh4Smb9uipMQWtRQpsLp5P1GQQyNurv/TLfAwqDi1w
rfOCINuu/nqbXgyTenrh4rWhl4PNLSaA72x3DB31RHgM+PUI3XyUFctk0z3OJr56
z8lWF8sIH4Igmt38TQHLw1MHbOxPUg/MtxKoxNrw6fet3219mqrgM5xfBC1HjQhC
2XWlumdDqskZUwXTeWVRgf25BGZITKLSBh+Zf/J1B5gIaXb0QgmGOg5OKdloeq6c
RMaPhlBAqSq+AVSU2XPrT6h+CnrsQzo78adJW1IHLYYzNI3taSwBDkBlTUuvVy7C
W2ZzZCL5M6uo4RMrmvp6foLtrNQer9nmvPBqCSE8qgetqyf9VFU6yAFs4coBau/d
qTeh9D7yc0UBB63WSdxy/gaJcPc1Ydz1vYgKvMVSLqn9uvW5HeQyFHJfK5IUtQhc
ZD5Puxt2SIUACl7y/D638Lt19NF5xtk5tW/milqbB0C6aY+8itPDQAgxY+d5D8nd
6V1p26TDTJfKQC1O4OGKhRfmxJ5Ysq4w6Hcaz0kaiug4BfspwU4FXZcuzk7P7MQX
wxP8vZGkGzqwd5NMxD8sxKf8HVW9DWn/dTRQnYyHRo6Ybtz6X+VeXaRGoXxLtOVz
TuGBavgP73y9Sc/uy8COb6rhoLb+9aeQB7/88z4SzW0Iirg8+dkvEnHwInOUYcFt
Hx314DaZgqR4DCnqmLSvHRhTcPyw03Kv6fin8tG+1+xeNPwBAiZ6eJHha6O6pMr5
U0Yv4gKo9E3IzEg34HaJurQDX8kuf/clZ2zRLcIQlk0eRtFNQISlpIlmMf5fY+iA
WzKSmr4YAVhzDODgw4R30SJQ1bnaNziP/HBlKiyj5JpIocqo+PoYGVRjbqe0SxJv
6goetA0PAeS68OlWhr9mY8GPyk7vlHPKeXFwQ5fZNwMVle4iXucw+ARfqhrqUC0P
OBUn/dSYeG2InYl2a2hzF9JCs8BJK2gLA808beceKNe9plHC9khSnSCu0sdoAvFJ
bm2DqfNf0RW/ixcAz4XJjq8JnZt5LAGU7xc+lKPdc2kfLg+Q9N0eImZpekEVsJgS
PeYBZNizQoEtR06gdv1mHE+JoX3RLiK5DHeL8dx1V3yCr42ENOEg/X1F6YOfTfti
ZQtcDfzDCr8RHT7sQ10ZQKrwpA9Ts8GqhlamXn+Oe7w8G2JNefG5Q+SkcNU0TFc1
IWiAeRL6rifpaCiRfMr/joMP7sSjKWN5HrItx+t5GN3andnKDFgCaB9bLncFEGN4
5ISESAvyZJTLw4iv7o3OtCgphwoVL0ruW9PTiCyJPifUrGadBMLm5NP/ag1Ajp55
lu8fe0x8wzaUZIz+95+3k43PBqPQTJk4fJ1DC0YbNShVToy68gnqTKaI62xf0zyC
Urdmn+Huu/jlWaMM45RsXl7kfGWCcLDJc9UAfnyV+/8KcqK8ZalIRMAYbGBIpJg8
goH0EljnqWk2k1VPzPKszX0FyqOmskASCIq99+VRCUw2wHDWeBHLu6Fj6ATCMLE+
dJMW0hmQaNi9mzaZvTpUn30HviLWcblLE5rNAYOstUcL945HvwM/efxvF2LY7DRG
g7KheYJfUgYYxaCavxepDfMdzN+bPRrllVWuXXl58iQV8NuxPokFM+QR+APifUdU
KXAadxLLdQNh/lW2YtMmlJBELmS3Vzkat1Wry/gzNIncbP+KMj+CZWk2mH8axIsN
3n/ORWJ2sQ2XfTH6kOSK+L5nW9b1wXSa2V4iMiIQkjTKQMRbUt9LEQhro+QofiSz
9UI3BB3EDHhLis4syL78Q7AIfJiXz+aCCoFpviJycyBPvOe0/c7snlCSrIUXGTEq
qqTAuXCBWveEb+D0B0v9fOWRSBj4Vq2GwXv6CdLrcL1gQUtgxr9yi31mJiEdaraX
LNJ721YryhyNcZO0RPyYClGucTcsm4dkZ/DnNXy+Ahd/EqE3pg0NCZH9Hy6kyJKZ
Zpdy9ICCqWvfPrOp/wGw2tVOKjPuGZBSgqMpFGtbcM1IN2Wp2Torn6HyhJmj4VQ5
LOUnEsdRHOgp+qufkqalEy978H4ixjopMQE6PqLcwYNUtMfJ6BCFiZcExyY7Kkna
hN9+TJqZEpdpKxVK0OjvYL80hZBjxU+G/DTQVY4y5gfd6U5OFEkwi+G98ZU+ANzc
ZngCWDCL4PkeTVk6nE+80QhGFqtQwnchfj83FSuVZzz2i+BPCTL+slVwk/aYJkeR
0lqQm9OVJw5xAEw0nt4ilpLTrwcE3fbOf3Ihwu3noR7ZRN2xnmZo121I0RFL196V
NmVmClPrpsT61bLr81zni4ts1c4X2fE+w5DvIlWuQMdwgfso1+bUcflYexBVvdLb
Guq/giE85HpzqZFZ+QOP7krpuSbkzOAlDYQJrwYKAAWnO1qAgpeAPzS0qwN7ZuOj
iY0kxOScJhXEFdxYNRqVt+LZXOPO/OYqIFRbMQqNAHBYWR2rIkS9Hpqki/x6Oc7N
In3xhPaluWwjKaT/E3RxeVbTSJNHRhzpcWJoDMvG8Xe9VdngpO5HBMhwFyJVBab8
n9LBN9+lc7I8B18Xdj1awoIzo6XY7RcvS0UpnRT0j9cpnhOG/ikTQlJ2Ced5iFm/
M/HnhSVBGbIzTAnEf4aPXPG4f4uXANslWyWVcaKuQYMG/WdxjJUCbSRPRdJkVk65
98a6ynM5JEaV/DvZsylkSDieVHzDOkAErLwbnEtiZNW/qEEfR3nN/NssnpDrL8tp
7owSRCBVv8gRfxXOSvZgKa+b0D8smwIdW0TH/8DEUH+VLp3cq4sfMDWdT28hyBtD
N4csD9lq8d9isLAVDhGE2V2eEFBl5ZkrRVhPkhb4HLfZXuGhTtLLJmnC2z+8yeom
1E+AoX1p/r0QBQBdbxJjnhPjX0z4VYykrxQv3abaq5VVJKXJhY/ZtZP+QyyAf4Dw
c/EWDPJTnOprP0HdLYyfGfyEHUWkhSLlQsxHrWkItdsCqeoBbPYBjzsXaRe+WEV4
9k+Fb1O8iJLLC8xaI6Kg7ufuaIaNfFC8umcOl82Huul+uUkaPXI776jTxVsHMtxe
1zJf71SXZqjQiRfAsejjZ6z1vbrF3zsBhQzlPp7mh2hx+DENSC6aWaCGewrM9Wbl
tkiSpPg7SuH5UHQaEbt/ZC7tiT50s3PLGfq8pGOHoRgAm8dMNfbitAT8QTs+W9jT
CfbERzQ7eQRp/DTOjUHNu3Hztmk4uS/IwEPai4+jmtIglI5Z69nvoTXeTBEH+QX2
xAqrtcKglOBVWjAmNt5vCjAQSD40GGWmDucvYxtq0luAEXBdkBBCMIdgPdbsaY7Q
juaXzn/+kSPRpKsUkM53pr3BwzJpkjDAABuKS2yXl+vlJ1oOGRDiJ84OL21MTxGr
UmaEE6bRmt2u40B2EIFOF69j212gWlxPLEH9ewirTXSDTPcoUQ+xSuT1K/ARYUCw
o7WqAFGP+SOhzQhllycuEhmUjV3UC4a6Q4T+lXsiI7OcQr9jWS0pruYEN/cCET/B
G5sOS5/FVyxrFFA0usAu4MEtLhAMClELxwYpsQ8PRQErDT5/H1rjCTvCh2IvyiI/
nXC+hoAsxVzF5wmqGMr9PCpWAFpDxgsPkqKJRwnJBFYX+fgA4EDUiTnlTIgdPDko
H7glm2P0HziQkPTzYN5fWIqg9RCbWfwjLKQTKXMS4TZxgrlKqNsuVY1gtRYFvQED
EbCSvIMu8PCOSZrqhaerCRBCVyJP79eUpB3fzQr2MribniSGYQmtYBn/QqADG/kR
yDayQpu4cxxzTb4ZSPzVNZua+ceCioLYzV35cGVXVMAGI69NDB1LfT++/Ilkml5P
FDKQgRvLG86SooFVAClQ389r0JR3hDMwtaq7mMPC7kyO1z5t6J7cw0N1uutOCqhc
RoP+Gnap5XUkYBsuyPvMcF8OGzh9WaVq1uuoILZCMYmJA3DLHEI0bX0+iaphRUDV
3atrLqGvf8JAk7TnnGg98FQnqFa8vcbbaDqZOb1QSlfOevYoAWfE8xI9gvz0d3b/
TDHMX0pRZ6Z+dOhtlhAf67m6TwyLh4FK1tqApS94a8dKZKNp1xugOfXqBw9s4vyb
tEt8rLfd4I9ynBTgjt2GJ8hWXkZWISsLlSYdQTT7gxjlHT18ScT8FrVRMwPoYp1q
v4Bc+0GlOuhXRbxPPzSJm//65IWBDdXyjMUZLFDEdl9jzirQXrnWhRlbKpTEdhxu
ZMFhSmlC7j51mNVidFf+GVc5yC30a9w1ZBqWLOWOh3/i3RSvi3nkzrdW4/vmeF91
eYNuhg2+JzLbtttCWYNlGwe8557xVfblRqcW/KQUiuHY6uyNOcS56JM8YkhlUYsY
ZuyjHeOatJ9NvoE/9wdTuVTB20Hi1ElMOnD11wxR/iBl+MDoWwqQ5Ll0vJ7kXVdt
pfqxBDhsOImLYn/mM51fplUxNvzTb0ciU4gN1yT9TrJ5yivpGJDmzY8S4uFBWu0I
IIW2XYrAAULpZ2RXAgZXltoiDmQMlG1OoTJHO6KOVEZI4Y/3YBsqd18sRu8yIU58
s6nethTpMD2gFU+Qz401zQ6hhbH9YXpBfc4D4WTzADfaAPMnY+TOXMdGocCX+6dC
o4hpXlt60KmjMPLn4pcQIubJbI84g8WZ2kn30xrmW+Wq8gWPYPNbYyR8GsjTPNcT
dg9elLdVtx2wBaaJhl5+PRCkMhidCpYGyz6/A4995EOnpr9i5koNTILYYKWRBRAQ
P9bUwgFuVcFczgOfOoQiI2YhiLbaX2h9YuVgTFkViOihQHm/aLs8SXcPOEbbGfST
yncHCSETtYcg2Sw/xpGMawWVcYYYUutMA1ARjhQPKPspka0U4yYnMzGM82lh5hf+
xHY2Yw4PpVfLR0kxVA7wxUYng8ihAyuctS5MkoLc4xm3OknjPxEsim95t9JuVT7h
sKC8AdrKRW71KPqjBhy7oAnfVC7NSpT7/l1zO2JP0Y6Q5qOpCnEAXaZ+4dKODCP6
v3BaMpgZWcyRg9xAKbYJD4P3lvcZIYZZ5E0AgYXsSLzneE/sajTTUcnhs0TUsmKZ
e+eiJwiWp3N2X0t4Pe7ImRuvW7cGA1Rd04R4MXl6HxKNTcZp7Oy8P7FCJqxJZ6iE
du+FkIdpNnC57ggwl8ISH7F+PYq5kEp7rPneSFE7tAY+fO6NZLAoIqCD1MrGMGxZ
VBzSkxrwJ4p88r1kMt4xYKoIADmGsShu+vR0U7hu6oXXUODIz0MxOV5SCBTEal7s
RZ7Wr0H/RV1ZBB0uRTOVkAtOQ8GHWe+6ZKfzMYsZpujjKN8eyobDFmMFMmYNNYby
r0LTUj4V/CES0/JaJNeSS022AUvciala7tr+wjOfn35ATn/HCf/xrFIRONP/1HBP
Rro1hrYhDjbK7THX2hDkZgPagJA7Dd9r9nrsBE6HRyhpoq+AgbqwSRCRqMbrPrQI
klrpTsgiPoZr+BJl9Y/9GbSXte6YvHmh73suW6XR6OJG1O/GPtOHI9n1JmXCsnOk
f8Fj+p+law1XCa+jIVvOSzWWlc6ovTQK/RwGPvsDY8VOgI8cL9DOde7fdyVlN1pV
oTA16ID+5HstxnmDtLNPxc5Uy6leoxKcVM4+vebpet/KYLE6nAMBNbjJRsza8kdd
zQTz3vpTcByqcw7ko/oy0JvFDoySJ7E0OIY94NMUeTLLcIr/HzW0z0Yx8bQ+wk10
0NT2jJ0/7MzpbLYQOfB4wdHbIcinoD/LC23823IPDZ15Bdmxk3u5aawoTCxvLRdK
yuXl4aLS5hSVSyKkJ9SDhwZ5A9t6pdb8XKJrtPU12/0lgq8ArJ/lIw7mLncQkACu
NtTWDcCz5LNZByrRlszOEdi5YBIwSrl3Dh9TNLbadSNKP9vU2yOxUVNuUe83Eu9O
cnNeJGpbXiuGtZImAgEPWMI16wmKpi047tLn0IWLA5IEcU0FivgVGO0MFSkD06b4
Tj35pD/3J95N6F35O6AKQabf54DchMUiuvV/TUSe2S+P8p/CWLDyd8DVnMtM0nN+
6mwUUzed/THYzRi0D1OOKNIrnnKuDarKsTYNCxvW8xdSAcnW5+LtwAQbiP0vOLPX
d78PbZhdE2Xaj2fqF5gOuL6m6P9ap/QMB4YXPt1VXxVcVEGsoZhvlv5b3aZfc0fR
lMZ06/8mOPvBwyLZ2GT08Wyj+jr2hIwBy6aAx1N64mutqjVhmcQrdhfPT5j2lh5R
BZJp6KS5etnN7lJgj7bBFWnHroGikDpcDMw1atZD4dqYx1lKlG+JEUvbIUlAAoYb
Gq+TgoD8ZIgUlkj/CPck09C1EV19YBZmJXm2cR9/28ij3B6hpy3zE4oTdekhykdI
dhBljSJbeVy/kb9MylnHcmNmfMCA3D56l2K75+39UgC12HztroB/Dz1So6eseUSm
wRAgiyQGxEbqoTLiAr7vU5kWqh3bQb3WxUiHquqrRvq3JQhcwqSyKh/5viAWpCzK
Zmy99FCqTRnKvzK4GMivmfEwb4n0zwY+07xj+0ttiWmzydDmn38X0p1ZzGRz6TYi
3sgzNHBKfVJYtvJoqnSLXr/b/MsXOLh7yZWYt4gwEuNt82HS/18/5j0lJwPVk/RR
mndm/k2U2Q2hnyip+1f6IQE1VziFsQ40A9RNnQ6NA2V1vdMtvz33ADeG069U+nej
oQMFo0iAVbeCMDFxw/Zaknr80wPCGZIa74yrpXQO82QhYHOAXUgmYk+//Ht3ZzvK
17iUbU2+2xHreVe2RVEA80+xeER0pUGjLshIxEzX80VMAoxSslcc+gxNM1krTwwM
JzwfNCa0fxgfgcQhF+M94WdVvG9IIAjnxcGXpvrpciHjOZExtIRTFQyeIhBLgfk8
jmbUWJLpC/n63vOpfmINo044e9H/+l1HY+VnmBeoO9/EPIoXo2u5oa1BOHrn5XkF
2euN8dJ5Rghi2UJnCILVGlkFwub9We030cka0GARDAIWBMMrTn4fR5Z8Hx2pKqDI
7WyDRN8D4r7C4renLMf98kZ6MyyYPaLWt4XXbi4ymjpmNwF25CRXw95SjnIAbe5O
14sJ9tsWB9MWOkj64m29rPOqp6Njws7LvnoXCRw3FrTrNvtS1me/4bLVqgAxSXaG
afd/XvfC/xSsdBK2Q44kn8UhbaHCQ2A8hPuTVQjvY2QCblYa12C7MYbvhnPy51O7
RnHEje9lMBlzM6+SNMhpiv3AO317Xzdswde0ZDeij9ymp7OfjGwEX96o0b0VlHj/
mg4Js11rpaE39vVMK19O6rEzCM63Jod1gE1MQrq5n/Up26WuuWJEOQMFtj9vaFnU
3czPcaCgLbcX/m9IUCy5UeIPOSFMwRy6OqwTI3O3UjWqehVU+34dpbhhb1XhFW06
cK6ln6UssNGZ9/bJ/+Izv20yKDgjuS5R7aR4UbkkYxjth4usCefJ1AIUl6c5B+1/
E3Fs4vrUqbqDyA0kY0lXjREfAmnn2K0gLYUflGLsGzYWiUF5b6x22POsZBDIkDTs
kQLRf35VuxIhiOnKmWjOkjcLbMTSdMB350fD8saqy1drHZw03JNnrcP9Z2TWIVzp
w0isO/GBWJZsviCSHw5kKnNKKb0k6KGRUUDQIcqOUvv5eJPz5x+6WHuvun7MrEVU
Y/6mbu//WPo1+sDddIziEITgCPXoD7GAFyprKmtUof/GaPzwVHY1OrwK+cfApVKz
jmv9Vh/RKj5Ww6NACnAFbPTxSV1fTcJBZJ+yqM8p9SIHfXTp7QwagRLDJLNhkQ23
eVrMAHd5sWH88kWC7DfqWvaTEx2kV4+UXNrT9KHI30yWs8xysBH4Vvpcm189hZzT
P/OOysHk8AOIYgbcWoYriQr0UKntBBlZbT2pr/RCumwTU96pygcOc75gIhAaJ+Uz
m7kFaTwtVyZrE4tl8KbPqIsLoAmYUn8xTuLaqfdRDxwWyA2sfSKqb/qzOaTq0wzv
wt36FvsFil9VZADn/fsh8Fg77ec0P1YhT1TTFjH2+ltEGP8LYlu+QN7zV5y+jx1u
MHOxEpJr+gv4dpb6W8TgeMwC+RF6BulnNEXaIpM9exKrlreq9dDhyfcsfmBhM/6Q
Y0rj8vKtZvWQtKEgsy9N/ZPtbBzuJULnlLEiJs0NqNK5khgX9nWCQFxrowf3nM9P
8tySHDAcINTPh8Z29UMRKjNBHlZWrMzdnAjpGVCdEqGvfsAOaq8xHhICdiJEM39h
8mgw/btvQTWgVVYiz9HDe2pLvDyVkvQV7qFmcmlBWLpm2yIx+58GgsDWWUGtWLl1
PDqvWVJ2LI8nzmV5nhPdsj/eV8KPECatiDPHRKgF/pAYKBej897fw7AtMfYkXfrd
EdY88DIlNgef2TEyLPN026C7mf6X8AGvf67UfWf2Kek14u2UjMKsqlmzRf4raGIU
UCTKQVcK14mn9QFW+X+FKAQT3RQDI8eOEPw3ctGxh/vB8ir5cktKO9m93CHRpx8W
yhuWYHaGEbt/DDLl51JuY/T58mPETEKdC6QB0bxHfc3ODT2YQoqoTyMgFpxe5+//
fseDG3NkzUu2sIZXp1KCoD8e2vnpH/XRGPp2tK2NrGfBtrGFNykUW1p4TstZqZ9t
fR2KlzJejUIn9AGiGPMWNs2/xNUF/2HgpAW6D0kdXzJdWWWJvn5uDSX8WJzVZX1g
/JiDwCOfi9YvIY2NqJvHwAL/1JEZ3iKAz3zPL8jjtIafM+inUrEfveBmP6I8VWpy
mofyfL7OKnthmFPQiOTFTrHV2SvQhs6YfknIQQu5TKi2XMiW+D3X+xj3KqQRN2Tf
ECD+55yLZKWEvdZIoQJTQmHEmyNlKTsDgL0SrHiKkU7TiFfRTgJXOHicd4ku4LSP
JiNO4haY9edSFp2FZVIjooOwejgCSXcq4MNlanaHg/4y+diFhCQPBxs+XEbXJBWs
yNfuNYgow+sFQ9wszUwUG84gX7vue4xpiU8gR6Vs1ate48a9VdyVsseJRCQrDaF6
JLEGLCadhSEwCeAdwlCTt1TE24fvsBPT9iIZaGOZYdQIKkCo4MI6U0mwDhKR2aj8
i4mm9f+SZsGE101sPhK/QqiBlzerqA3Ux5ZjOJQCn+9IV926nUP4vQT7c/zHWvye
XVv6RdHw+lSFENNSyMZqzC3urZCd56+rxaZzvRo5l2K1/KNeM3Z+tckyfce4XdP8
qyt7Q8UALHtmu4SrbcDrsMfWzQWmj2mM+daJy15saPpu69rDKktbvdCdTYXhqBBz
YUQoiqoIhUTh2Di+O8J/rmTdcKQSd+KMEcXtBIJDR7bpwEp3EmQXYTO3272YPiFe
IwTpGozB5H0Qa5RyfVcVgXpsaWiwQfHLIorxauA30vaex75IDBW+uw780mCbTvCa
z5RntbLT+myLm2PEp5KUdQcdUDvdnkUI/ftWbg0aJTRU5yf0AkV2ykO2/nJdcYpK
nDKVv/jNB3rrOD39d0/LA23m0Fu127ZHreMn+C6aHuPwiN60OppLkUXok+Nt4ppi
5NhzBDrOo8vAIumB4Kjm49XpDq3MZdi0tPfA1cBsEi8fHVPV2bMNM9fQXz69lbbE
M08quy6IfhqNOow2VRCHAgxBzlZ/F/6D803Sw24ntyfiZvjGCmh38wCLOWhUjDy3
KRpSVhLYlcI/gepQjkqaa5boNPeT+OtooFnjlXf4SZOD4PLSyGr63ExCbTove/kQ
dz9Trv/qZrlzZvMjMOCQfJc+6oq/Vrkqqrxav1AXe4+AeMSE9/+wQG97J+agTZHC
j6wqzY2wdDenhyFi2bVGcITKBiy5oI7Vt1//l2+Wk63S4BpnG7JGP3sZNb4ddv4h
q3PCuI3WjSVjcB7lzdUvBv7tLCewITftoJKznY0aNkQw6XOOVoN4uNYQIfMxMONp
0k4JkUlHisFY0YxZpXR+su2EXAuN15Y4lUBmYU2KDCbGcRTbB0eo/u+o9ZtJXVWk
Lq7/Wq7G5nq9lAqoyOgg3eExxrTK/O5Gpwbu3NJh3KH33uV27ItkQ0Cw+hSbautR
o+kxIcPjBZ5dSJOPLpdpal4XfLAV3nC2sSQoXVafFsw2YTRzjrog4j+J2J5paaHI
ojpsg+cEnn2Nyxj+cJD4Mwnql9NQG+49UvFiStpS466SR2egeMyWHpJl5PB8+KdV
4YtgjXEnXgKvy6hHr8o2cOCEMMPoDYyuBS0h41DFdh6W6vDkynwufd57/+u4CV36
lXQMRl7FDTA9D6JMmJq7v3uKcN1NU81CgQKv7L+/6/TKOrA7SxWBLKq9SuiDwMOr
30s2rptQDm6+75quGbuw7KDU1to1nie4ATtqAUCVky1dE3AO5fjtplbWl/tDlVjh
rG3JxBrTvuvOR7kwVKPDXq3u06YtRgCsHgpOGtjdcHT9hkTYP7wis0/8Byj1cq3v
E5ScOC8cehDygkMdvBcRoVg5yorQZfoXpYgpm/bDkRlMJqizEWZfYFiE7AjJE2B5
evoJNQnwm/BBNO/EqVj7RFjigqcMOyX6A9h4BMdm22d3NL5dUmLSShVY9/yeUy0f
nC0YCSOo7JawN2zqiXVVZ7iGLJXB3ZRSV0oqPtx6A771FwpC5DeYBASOOI4l/w2R
7+zacd1F6UnwJoSN2quytL40g6fnlXuWgn/RASpOdrEkLGPyDdTN9XhvxwkiY+WS
OlWjYvEKzvTY/sS3/YOLn8LV6UG7c9DAluOBmEMpQCH/e9hAwTTRmh/Hwh9zuKCc
uaMQZLEPVku8DTXlB6L9YJLq04xTn7DZ7Fc8nPRFgl8WeG7AcRW3WxQKAV/xlCA9
hN145aKYJZbyGDmCUlwqqR8chZs+ZAFAQxvNr6T/0fVWeS1YJlHMd7sSo7n2ogzP
u/3cBeD9kJUiTt7ZOZh6W0iGwP0u+jrdVUahiNQQwEOdoA4/ptiryUQqmCpy4+mg
Cf/8aN0c545bjAU/SCx1Qdy1BZDpi+CK+IDiTXy77IZgUuXGlYKqTuYP4jRDmra3
f8zy+2Xm4b357yZrr/C0aelSCd05fgttyHl3XwKNECzKsddC8AoOY0+/674jhR9v
159hn+jhhqQ2V4KHPIV+fJO+B3uzoSxR4O0TWGAm9+ad6HDJgiadXFkCgru9KC2f
AqwqBT6BbjWpz7T5F7V9oRk5g+xtR+zHfOKgDL5yk82cLAWg7qIBtSXEZ3XwsqOG
pMZkdfpDy5z98G/eRg1a+KRPJDAiao+c6oP+Rv9mXP6iRkjJ/rZjOx6qfVOe3Jrt
CJ1+FMbjRC+q/K9EJO4IYdCPzXRmpmlHJgRh7JRo9sxp5X/siwG+xAhv1w02GmP1
hTjdtGI9JY9fhdDItjAkJvGAKLmUlJfmphsyVfbLKIQSQnPaoorO9mBQJ3FQH9r+
jQSF8EZA8/bvLS8RMcENQhD1ZIxBkZ5bbsWCKyBEIfDmTbWgYkh8Di2LX5esPjlw
pbdAOJJn87PPWnn/DWatJc3j+ZqqqncZljS24D5H3OQr0z1l36r0+gZOPUblbhFS
5PNAO2ElFZ05hzXopFajJ4UQXjsf1+614oWRhk5ugTrons8en4iC0VooZAvuFqI8
pZnWBdKSA0G4zSIk1u70pKC2nCU4u3A/cxhLv21/+tt+jCv+RlTzN8PjHIjC4m97
+eoSvi6AM4cWlKb/EGo4ZXKHl8rQd6PiBQyz1ZwXQmc0yqJsLZ9ioIRohyZKN9Tt
X8tHBfzGkq1XdfTAkKqpENBIU1AgO6ePU/BvKPDNCg7XFIBzhG3Q68vaSZMmgBbS
734nkFboJVqYHesb66568yXNny5kuhovrCquhrSr0jr9wYVTMWJFyhd8Vg2Zadfi
fD8IvtD6LYpkJedRcTVdAeKxInkY14F+6cXcyc8RSWRG4oCWm623mPWjxzroALer
S3tnL1ih4dO2GMxsnNiZurBgNTGehB9GKtAO84nfdxY/RlcGfelKZxDrPm0EZw1b
9lfzRnHbbMUg3NoaYld3vKOvTYQ34Z+LHYEhiVslbLpORWxeLwYNZ2jrHs7BEb/C
M+Frq28l378eLf3Ljx9AxWxkprFcdqfVlpQvJCjxERWI0x+6lq5rG0cEhz8p1noA
OTmbZrRdfqFeOXFl4BqdLId0mdHPqcVtOaLjmn2c6+CAQtzEbn066A3I/+gRZDtj
J6bHJV1oGceHT05R+KtNMMDhjl3P/9/9aJ34iKWNW3W/9YncYtte2ce1k8sVOEBj
LOssNJH1Os3DUDEHNwXOVep5M5/qAyVznPT4glDDKiP0JJ1m2FcqGZtXnT+AQsmL
B5IIs6umBuNEsGZa3nah5KXBS+O7eatriOGDhKaU5JJe2OcmT0EBlohuW8i9EWUp
szI6Up7VLmXzJuUdywp8XrTASn0wJl91iJmYp/vb3KWie/HJCwbfnoGO91eoVf5m
C8lTtPO8Ihs5IA9dTnw7ZcVSvlW/KRLmIiRpgfIn0uDtxZ4Rv2bDSUS5gdaUpM82
iVl7dZVS0W3hnRWX4Kr89AKJSDE+fUkK3o85oGqTwkCIMUT/Gf3dY3XDoBZf4eYP
mlqviNynvKdGlfsEBGeGBQzkjJfIfgk7n074KCkSAWQwtebDXZCXdLcG9aJ9atiH
GObfNILvQTTS6JdJBfROcr9O0J/P0kaijHcuib5HhcPm8WBSHi5ZMCsMdLiVoQp5
IcIxQwoGs/QeRkmNUy/xvIFi1GVtAODSaFSw8XROCL6ZNiyqrn+3EnUvdTgCeCbP
j4neYDU2CRLrvi+kxHS1JlfR1inDpePFjoWYjXaEcN0M0glDRMLuH5DxvTT0GJ5m
eILcqRV7qS+QyKowwQQmRFtJUuGzbqhY0YEmEGttG/S0z+XRJWXITIsA3vclOMIe
8kdWJSv8Atv0GcLYjqp0s6Fw3QCamaEFo0djL2CVDneDWhpt/RS6oMesnnTcs3Oc
cBh//9tiU9KiQYXE8X+7/qiICTu/wKuqo0ptADXV9r0h6l9Vy7k6RYA7QKlha5db
21LghwZrQqnxq+s2fCTuPb5vGX8tKftJyRAgJ9Z+6HdBfddC3siiZkqKNjK3fJQN
U+vE30pf1W7mmxilVbfcQJUx3QxZIp64tX6HXwmjgDcARVTyYuqmPBl/wxUgz/Q1
pncEipKeLDTPo5n2IUP3JsoyZuJJ4a4gQ8YXHEXSbRcIlodc8xIT/SbM1Mh6iEEk
rn/4IjTFwoXmVYUFqG6UX+mo3ydbZXD8RvOC/5xIobG0pQaYoe+/j76crtEjvFAN
NO9DlvOdFGJ4M/KowW8oRb9Z0T4GfTQ/2ZxPY8T3blQIYR3iFfVqSIve2gsZuh07
2fj7fubjJdU6wm9cJZ4P1g7hbFvixGXDFfmPlOf1myRkRvbQ7Lok1EAsXPoGlU8Z
5fyZgkUdzvXX6GS14NBIYOGZuU/2z8eIqnJrHuChvK4yM8XbJoVouXsYKf5WUOVW
grKBC4Dq/eBR3m+/QxJEAA7y7luIZx3lrnnEri3X3w79LKAqxiYzjRSLtopZOVp4
5FSWKtng5wLJskeSVzIIqLyHWAZdMnilevBg36mlQ6oInDuP4r01m8F6htFfLjsu
6IKKAozhvsVhu2jRCk/5DpvbRSWDEvu2vN90PiEojqcbh4k2gC8Dkrw346i7XLDX
RUeJREpwp9RHdGLYUXcb4mQbenRohAuuF4X9vG0HFEBmV8pNuMlotA+vKYwEDmEV
uzDnhh4iO/oVXTiYOr6PxwPHhbaAgs7mkrZ4bpH6ajzkmoHOTp2SpG0LJUxz3AKQ
f5/tSRVv15vV6mbHdHjw850DeLx+DFNDJrfCjh0wQw6e6EApO+Bh+odUy7/SFnXc
Ep6UIanL3Zmhw70sXFjaAJ2zfyNgKtN/BEcdhZK5+9tSdqFNMrNvWX3Ob0kD6kf/
jFhR+uXcdRTUfoQevQ5WtwBQUU7Lt6tWU0TK8dGqVdsxm9GlySVxN/IqRFr6A67j
ijwPCtdV36aHudfZbLJJOREFsiSmT9/p/ioArlcYi47SvvyJMOrDjYCymgXt2mDp
X1P29eQjHjBfKtME1FMJoFtPCymi/bWtyUQ9E4qR29jPqYrPLFDiDSpBYtBCtWdk
DUIBMPXTm+mioTQHv6zk0USi/2pRXH/1qS/e/WdDJdZTD12wnDrpGJl9fvVEboHS
x7ZLzoPucmaVPSvTKnLwk9pJYFQUmrSsPsIHIZR7JPKOABnipY3OIno0UPSzv4E5
L22SiKboNuzGx3cMK1YEXmUHtf5ETAIBKFtFNMqvmRNNyng1H1O+iZ9c6nOqLjfK
qq/u9Ih6m7uhMfYzM2XM8lUAgI9SCjaeYItQMpzUcwNMM7Lz+cMtgzBXzCjNOztI
3gRqb4p3J5nJEzCm//ubE++4lDUN/K+0TeD7eO7xUrQis4OKohi4dVjIDg3Qw+BR
fTSYV+qV967Q8HvDAIcHulYZYD5YcfNxUDkLqT4cXbO2u/3JQKhby5DLS+h71Xqn
OThrRCyAjjW7FUclayYnY38Cn8Eujc5vuGL/Zi2AO+JxwGju+izkzNmpazmfE58J
EOw71NCJQsNKs3P/NNhDi9sb96bCcxMpbbdFgbXFMitzj5QNgUcubtq/kZD4L6oW
WW9cvLnNg282mEdg/a7009SwTbFy56gMxY11XsVVnD3RWnh2JdUvM6FFeuXqZSl3
nOLMS+vD/tyjI8euAG1V/o4HnOu3lY7ahuS03dYpPNGNkEhtFDm7qdDd8N4JVOfT
3cUHRblzVRs8hULQfWdS6IwezP6+XFJakWnoC44HgHrr4jNNRXtKdz2Jle0/yxpV
iJ0sbLKJAtN4fhL34+9l0kn60vxMOPLWKsd7GoKYFfspRZhAGCdYBsnrSgzuAfBY
lW4RVTcLT4T8NdKF1+dtPjuAXy5QEO7mrTD3LxcEOyaaOm5rR/8ADYkIe1lL7ZMu
pc/G5pnTbj9wH3hOy8hWmzHvIO1mcWbKVAG9MLWVlydT4t5E32I8QuUu78zpD9q1
RiE3ZDR6PCBh/borZ7F6kQfK81uMk1YKYadOBoJeQ076ZH9y/vYY6tS3XKr0kznn
tI5VS1yUEytjxXO9DVuozneTpqK4hzg40dhuD2ahr9wUB5VIYNaKvXHCf5RXkqqT
X34IjOFBnf3ZLLrQBzJQAU+u36p+lEWx7ZMEaZeMB4Ort8P2O+SLe4H7TndzSggX
POXgqF+9wTfywU/zyKcKZlx4bkpNsyg0MizrahyX/gv4sncmmm1GUXI8r7h0zZdX
IOY4KrIUcssKCWWicHgsTQBkZ43+jsupXFGLL2JMZHiN2jmi6bFI+oA/c3niczup
z9weHkSkwtqgErNYv2NOg84502ZuOB6KmP9xxN16dnqBTIcU26yHZZ/Z2lxULhJV
JgkfhErzyYqPOYvog7mth1JN+O2ApJ4rq6DfoU477ohRARKQZEjPFOqU9iCkiOxC
B6L4bpfJvyyg83ucHWrnsQvqlnTWP+1hDbSYN2bx4uzJ6xX3HCtd1a6FMcE32cd1
xQe5AoInpEmOYToucCssI8l5I56DivoisbyWo5rQGWUZn4w4Q4AZZc2/C64+bkcM
WCIatlvpF6kOJ7eRh1mupCvtFoOWlcPEoihynkHpb4CWjE0xG71Kv1cnjvyeKmBh
1Ls0lMn8uXkUaq0IiOTNsDVuVZLj/6C8YpUij0CQ/kbh1ShOjbyxQSCjdrT1ME/6
kUDnf0UqQG3huXqA622sdcjcGSBB4cfvVH1UDB+kGj+76pj9/DYWRAGVMeorEtmO
jxbBcYDwFZnqBr9M0SdjBa3i/Evwk00gdvES63EY3Mg0d+ZksrS82GLIZHD8t185
OnlKONFs+q3ubi4aHkpuq6xJBCfPp5+qiT+m/IHdc2qQ6Q3y/ooB2NEeO5Km8YwB
cA2c6uCqTPEA/c5r9Onb98YPkn93MOIDAvnZ7jxo3Xmf2gKN3+WeXDJyHH72l+ul
yHMmhKgLfCINjTopCQZKiFF9kcROtdPD8GZUGt1/4gHVkUzNGzZ3FO3ZZGPOKvTN
B6A2t4Dk6ExC6m8oZ3fHyMGMeKjlkGeExoDgbo0RbTCYAIEkTrNHbkFdf8+/FxNm
o54IM6V7dOhLY6T6UQRuR5zq3Mb51VrQTo4D3HqqcWOggcNlUp1kVtRf9zx/BDfu
68TnzyYzmmAkAIYMmqP/88hMfFaiqPF5AqMyKqPIpHe2oAcOAsoydzuksblBCyl9
fshQKA4B54PpfX+IdKzg7u+vWa335zUQMmN5Dbpp2+YMcsb8lNgGRzY4UX/Jcr5Y
TWYho2hKMheFrS6rotfHMYQyi+jFX1Sygm85eMjAmmW2/2EitNJB9Y+2nzF5BJbp
b4g2IlFSSyfTavvdw+PUpgMK1TqGTKglsZs/X3CrcA8CHa6nvdMBYNpy4O7ODA4E
iH+XUsshnSVl4318SP9OmvQvzWfQYx4CYw4WSeJra/0rnd7pmtSl29kXpMAdQl1L
gcM2YcLRGcwQ3Cu+6M8QW/TmPHaeIQsUAl2A4YK+cuK4ztW6mlFO0yOG3hL/0Kll
x8cyevlrPB+fyjp8MAgu0X7rOPSjZ2e9Blky2pwPWlbEanfEYKi3iNd7JseTK7ee
xNUGgVAviun5tk9ZYRKi0+SH5Il6H3FhPTvZUDzjWPo4R2wufeLRzmfBTTF0AMMl
w8BxKIlxA3xFz9ALTNKLQWfZwBtBDbyeDBgZ09ZUWZ1oSvjIonkv5O3SwCX1d/nc
aORm2mqJaCfCEEUwqsJ7dKwD85KzR33tHOaXcPKfvAMvp02r0EWs/ihaqT25TCtK
+2RmIscrwLpsKFTvxPjH9YvjxbDZojZ5yEWZTTpwhbiKXBBnG/EYfuYeuZIvbpec
dy7Z66gwzZUwKBtecVtp1TPOfcdIpaiUYikdgqe51BdNaFM3ZVm+roQ0ZpMHORfI
zI35RV975U8r4vMsk0l0NoQugkOJq9nK3qyh6PnVjidghqyToiN5mCg5iwYO+4uE
wpDA5q3VErM2C0xDrsokpjZhwKw/wZB8Q9K4KBaASLphvLasKaKD3BWs5pGLvLZO
gkAE1/hz4Y6QCvhnf9FzeBwQEQAyj6cld6O1Y3vVNaChGne93TH5g9YzdHLcEq6v
dX135mL5T+v7DyJ5ijs8KVX3/X7ox9z/eqeDUPvaQSzbCGviCN3RTGpR0lCJ2QqF
HSy7Z4CTApcQbMeBmUtQUV6Ydp5yZLL+sTmgdX93EjlTqYPoGRDvqERHmqYyfFz9
vw3DPnVGkQ3d6Jrc8JAipDEUAMC1Xe22sp8co9ZOBqSleOqwpzhvBW7Am4jNp/gv
rHTCE8RuyQ3J2+Y5okpjA2jDFMwmtt3ZppY+v/h7PBwoGnZMHkWtgNl08/gkzuQX
pBv+HmH0uoSdLqaQbnR/8Rk+1e/dHrBpmJOW340DVEs8BC7G4pdI2zEQ9KNPxgik
29b/916C+hNC3yDEZt/clGIxMsFNbrUlAUy8ucBG2K/u3L3ht2N4hWXiMEi5J+0g
HM8RpSylZsJNm8WUAlW9oJhGPZhLR35yw3lzVhCA9TY2u0UTTPR+S9/Ntrzm2PwO
tkTVKLZC3DhW0uQxMLegCu7qkLwE/Wp+XYCEBpeqJmSiXCsyBApyrPvkM+vxAWt5
navNnQVC9rKHl6Dg5p3cR+idbF3CyoreX+iauB3n8csYXCHfznpGS4bkHA2gg9PW
X390i4169IIXiVceKqS3m864BYXAocWbM2g8tEfn/yehF/QpOHyZJJFovAGHcdTO
3EvKkrTvkDNQme+JWfJnx0DOw3N3iIanXPr3uQke2fPNakvnD58IqDlvoW/DmKRS
gh5ZfZB9IooEoKkdSYDIdynYr6unhfhmNsXlIExdUBemeoDCx8A5gzDRt6YYWtCD
DTk52oO4tfUPNPdJ0XNDPE+VOZhcy944D5eG2qmaqORqVZubGjC0+XyECX2pBFbm
STKjn/9jxQBDVloTE5OEObIDhk28Cw+8QVHBo9Dci0N4VV5/P/ap+dfY6YQZMYJQ
DFCpNHnJx8YB/ukAU7s/pRNGib1zjdaDAGVgCmSgWNs7O2+7BoL8AerG6yLfsYUp
P9lafj5NEn9sXbC7+FV3fXOADzIX5hmg1xQIScrEwCKg9wq/e18GbBWJEiy1In1y
UTDKWeppgwU402O6dvTBxegABlxGsNTeGzF8scdCGNypULYi3VbCMd4XWe21gWPz
mqZ6D/H1LBy9aJq3V/lL3ZeVd6fxAt8aL71YS2ljNP4BjwbhzrFtnq1dILKt1pt7
BAIHFv+EjIMt+v+Od6Qqz28NiH9SZW05iwye6/dSa5iJ98vUj+ECgOo1R/PIPoVW
qkeiiSCTa3dfc44DlywaBwowDWrlpWkPamyXJMK6pzfAi6a+Dsh0+nygJjMvTZ5e
FxpJGMtM2pgHCa+X/hQdfqJ8/tjbJ+jYw44wZxEiIr7wjk08WzJXGB/P0pJxYiak
BwdFFNEa//6TuQ1+1WR9IHtZEZg1aHgNRlSkeVXJNRGtBel82soLudllPK/+XY7H
RVKhBvQzrUQNuZnriHfQsNpEcKoU8Vf6wATwGjMg3vNNCGVACD8V076UlmooaqgN
3s0SODDP8lhcZbINXqgIiGFuxeuNaP9vFT66hBRqsXzh7p3FVGJRQqq11pkD2y5j
csAq0amQpdjoBGBPct6SWJOP0GkMtfLwxN2L2yBW8ppCskDQuII5Ag2Cy3YXAzCz
8RAEUabnlRIvlc+dm8e8TS4VZenvx4Vxr69tOQ4ZL+6dyexZw7YWCVDLmufPo4IH
A+VOzO8+YBHEPHT47XuwQWT1rBM+OjNa4rGccrx82KYva/vRxeJfX5sM7pmQBRvq
ZLaq196FKITEIswKOtegZ/b3N3SXSNB+5ndv4ZIeSsAeACiHyvFEfd17KcUZKhS4
7+KaL9s0LIDN6hSTXDJuiHWyatmXCm7YVPGnQbmnAbduhr5cbt6e+XrXLIjeO3Q/
vSQaPu59J4xBq0J8FMgkm2ubH5lvRH6oP1vcKTMevVYID0QGRZq2KLxZ+5cSBi+W
U4Q13jf2atDCyF9QUnKgJFRUteOkEo3u07uJGgb7D8q3X5xzG0ZYEbSaUvR1UzOE
Jqu7nryZWL5tNE5eRryEeF9wO8ZNy8mryD5OqlNAeNPAJGsmGA1g4Z2X2ZPTyBLj
ufgtUQ+ImsC+L7Pjb6rYf/jF26BbMXvt3/XxGtUmRymdp6IUGEQnv6mb1H3k/eRK
9bsK++1g68dmrQtfNcLB1C8+AK4dfmj3zxBD9uso3KuDnp9HGM8pckEUXXqQHYJG
AVXG+wY98Y0twTpqx19SMBeVXQueNDdc2u7kEuaOaC6jrXEdy7AM87BVGtzguyED
D041rW8dQb14OAiDQxGBk49seCMQmSIgdwEJtrQWNH6iamnbgDUxMaXq0kz9cGip
yE02IQRorBpQsbodv6yYai/mqcYVPwBdcGN0wzM8+SeTom5VN/G8Lxiz02f4vCRO
L1PXkO33f/8CfZh8+hyni0EQyq5w4uPboV5xpJ60lZr6GB4X+xn+SZ4hEGp70oXz
2e935lFxE/bxGq6uoaoKK9LSmJr7vckpQA5kqcJsNKYOoYyr7xPMiroogIg8iCnL
lxMxaJtBodBBPupokWqNLFPi9jbyuaS7jN6UaMna++IeWLv6F1hm3rBNUqSKb1dC
XvRZ8v7yvVAolpiPLMaCeB1jMBwot0iWqU1phvLo8tHwWV76ZVEG9JaPCY+Hurbm
Gij7xgymvQvCMu8F20pLTa95CgDy4XyNgxoBgw5979zhXk8T+dGDp/UnDopTlW0M
qjZqP+94JvgfR5HFHbyS4m4pCtSYkmqWVBts4V5FH1dFF5M26vzDcpUv7E8CZ4QH
wIjYpJbzba96kdMt7z1wJyQ0s9LKCOZ59uQg11ND285y8HgdUJUyrDlSC1aX7LP5
1cWcAbzGawDXrfx/rotTlEwHo6PscFFLLHJQC6F+S3bbqXo83F75lyb2qSlTZUxy
2BHGdE5H8jGPi2yRAsEgPefBm77rqFnZYZRFxZjpfMg8WsRPtMTe8tdo8GWvQEKd
qkDaqJFnI57WX6fqgAXKO2EDkrz9oyoLsCtNe7vXhzKdbqY9u1XPc0GsJbOFSy0W
g2ZCg7Kzau7LTwdtyoZAw9fm7bciOwj2kYOIhj0f1OL7nmNxQ8uLLeapS0dVOdUY
sITHT56Ngyn+8Ces/I/8BO4mLIwQoWMeMmO0rehng4F/LfZRum/PtI2j2t9LqegA
ahy/3c0qz71YyFyz/10Ih/i1WiIwUDTT78kMbdOP2CVnTpVwtmYhQocjbROmJIlr
6dLWlLFA7TN+h7dh7hx/mlwxMPdZK1BvGz2bKBu8vOOsqmz+b9cw/Jf0OwWhGC8E
j6dWxMAEFQnhlp17AWSyFEZWjSGwdQoylmpNg2beT97rT1HNoamDeUyvuA5UWAXj
FpFtA8aNchSIDhZXPo3sMPSXBGNwlghj8hMH0ohlgT8Xji6JnbW7B7buMTk0VL2X
eImRL7Rb2fe34CIy+jApnbKhbzNtD/VSq64kGyXRDpxgtT2uy523/O+CZ9Lcaigw
IoAahetlJG/ATVEbAwju6azB9pEZhLnsK96q+HdRJYz0PwGvi/0qzBDwfjYMuhol
ej74K/5unisZAf5k8fOUX/7MVEInO+XzfCL2SPVwbfzLWHFYU3/ONtEPWqXAbrsR
E4OLZLt1EImZLRqFFSQ5txnb8PHRMIK09IIZz80EOiwXjuVXpWKA7nAD7LjHdQNL
No4VH/AcbeNjFw4ZKW2JOLo6LSKgNAKPBLuU0UuOa16u1Tkk5Ug9GjImIsOitgzZ
mDYuAi/PEAg6ZbfoktmopOlfVqUt08N1P1M0+GOkMwnb9aFwLTA+SY36e9/+qts1
qLw3gs9azgLdvUlpFu1oTwOvvEREjgV1CSumqf/g12xjOjaqOrUHtAD8zYtBm5fR
KLZFbKJuyDgskVOul8ZiEv/jg0+dQsqEikb8S68g3F4zp0ZzHDYsPTjPIXv1g09X
omvSP8Nndf69ojibHDfYiB9cN3ipbgxR1U0Dx94kxLni511xj+61LhALR/bEVlu7
fWdATMWz2slaCCOtaRit5cAwSEbF7WsomYgfCJazCidQXS7gKEVhtwVdTFbOcnUE
+eUgyWSTL65LwtkDzmo3NQhq/rzAX2iyV3NSZKhnFVlT4fTFJz5kpiqWIzZ6BgHG
ohkLLa87TueKohWUuVtcR45jdfxmasG9ugrXvztG3PjZwDXuuMOTNfIvQcZePOKG
0PYZ99mDLbOCo5yXzIjjKpBGLLm2wd9WG/ZGPR8x8igRASJo6u6+bVhpM3JAVHZE
71T3lXKj6bQHO5V+PDvtSdi7R9pf7wskCX0/xUutZxyKCnOk7Ncbhn/ZR5ZXcAkH
rolszJRvFw6BjE3f0Ev3VqLXObFiH1APlJhu3UdEGvp6xVHCryxODz1OL3LUygKs
LkEqsCkxGDMyH7EIjdRSdy4i4qb+kx7L8jdsQjXaN0efpA6WjzRX6pgUqErJHr2T
DetPxBlQUkFbKNfwWtMhKBSUJgoNnm4EKWE9dE15np0gsWtVGXECcDkEmlaHNuwV
MzBo0jtCMYxfyvpkUPT4SmlkUE4zgSc8z27qSShFVNBGuxHwp0Ev6dyqEzFsW63a
hjc19ZVK1UyLDw1Z2vhpTyu3adfivL2slhgKbNG/lTIfrelwI3fe/P+cEZKcjv1/
tY7G4ALc/k4QvkqgC0O3k/y+jiMsoQbJ/3VcsaKQuYuBI2c8BARdVodsmhpe63pI
GQJqPIHFvuj4RqCjPwgZ52LFHVnfjnJnSHrDWum8/B91LmAhN0MBXNUSSeZiE5/s
yTHGFPe+/O490qkcHq8uNpWa5SJYXjdCVer3hd3l6uIJJ+SY1KmHPd/ZZZGWBn9r
TDC/dRC/Qo395bFd5T0GD7FfRRrBnBdxk/lPqpw8kMlMF6Bepj8MHr8ebcpDwE7k
7Wtu0e/48SnsLW7w/q/G4+A1wNhhxqAMquMO/bw8U2uhTGSn13qQWUH3DFL4jLPq
Y98H9frj07pkmrfrXgnffj2WxmWG7Y8LMk29Qxd+BAfvqOjDfZpZNJEiN+qqX6FM
CJZEiq17KrwXnxiwJLExRyYcqNF54AvacuulKdg5EcGNk9jjW7m/R6NtrelZwwyQ
YMk+G2NNl64dLYX/x8F6rrOAwV/aE2PrRBwkpju6ea1QKfJqOYxteA5PEHtLpalh
50aCCdTcN5Hn9+dznZzMYkf1w+mEOpZUbr7SWWgcuNAS4nEzX1DCJ0G6kiDX2Xpa
JB521btTTr8FZZEIo+5KUxqngIOde866AKomz+Zaf4QYN76cZKgGI8TK1miX/6/K
W6Pew10CFC4o+/8Hv9ILaPmVY6oRnr7UXeOCuEy0aKkGNstuqCRK1MrNZ3VvFzT4
gArklBM53nNzDKFO5/udFYzzcltZTGLF3mbI0cTvwKuwtJQuI+NJJHGKKUE+aQOR
ZzSCf6SOUVSftPIBl+S8ED7N0EVC3zyi3YgoPqIY7Wg3IwN+FOPAgQTpnqURJmQW
LREIeVWzlZ0+k7TeOfP5UoQ0XekrYioQ4Qb19/e1gMRmQE/zDpcRDlV2a7bv1Ov6
/gH464z1mFxuTLRiEDQXt56i9nNldCOH9Ovxpl+xnravXpbWSpsE+KySF/x00cFG
f2/ME7geT17TNPdWBQSxV4RN1WeMc/tKS8O2P1i57kMOe9bJgEpKeBBhluUbVx9Z
YbyH4WGEwSQsvR+aTTwkHlRlgtK0eBhWwqD1YaxBhauczB9QNsebVDLOjj+2jdBJ
tUYU87DKsFKDlFQB2G4aDfkfsyxat+qJ+AiQh3Ms1CjtNSH+GspBSUtBQg8T4hih
jQ/WuM2n9AnDcGZRXbDDSZpQh2RBNbJqSaTbVrrJBtWQ+/3jIT1Ac8U+jCkNbAJg
05gQkBNZvj2e9TDWZubvzVJBIn/ADx/PsVTJHE8IUAhGIPtgrLYwfr8gL4T5lsan
oTeUyxs9Snobyq1XwQxumqY6FoqFQcGn2QNr3hL5OIhyXS6JO/ZkXKXstXfwCXAP
E70Lf8Jpm/IxFLmt7tke/sgeMsosvYfBoXLVERZLbec9owdIEUGHBLRtau4vJmzu
uiMQSaufqQ4aFhAzXBHn57JB7msyCa16G7/ae83JH7HjvG0IhJz6jStkvmdHgEnD
MBvK+uVvW64/9WJjAcXurZ08TrGIlZ1rzO95mzHwqqelEtwzidyRvRmpu/lB6tlZ
ocVhyhnuUikJR3Gi6JzQ29PcZJHF6N+Y2pe8DTZAZP6qZcyJJ36JupG89UbWDkl9
DCvhUlmWiLho1gEY/qtIvQqiPEvf3rz8q2kyGgPOiipRTGgz6vlJ6HEz1juAWqmg
K/dMNnZXhJ3skr8008/KFVFYF4u+v1TzndckhBoHeACpRQ1yT4FvFiUI+VSf/4F2
Mi+DzKAE4metPdnvRNzkYW+GbnHtKnhWuk+JgpQmXu+0Oivg139WMavq3sPmmeF/
f1SL9obA/rUJ3MZgEi8P9duRcu0hMoqpjG7wdokwjphGcXuTJGV/q+3od43QCC1j
7J9qRldt302ean7cdHroVqwpiV7R5AlPD6DSiGdZHKgj75f8Zrtq/ccEBE7P6gXU
mZXQvFARKoBfo17UdmdMMCdqK6P9CO2O0FGKOBj0XNWuugUNi+2Dk5d4qKA4UZ3v
6m3PrtIFGw63qovUM4dPWajia4FtLmEh5wn9itZG95EO3PxvItmIWphtd75qZQyB
lwhmNs4SJWTF6rhv9HAwJclICKgGyTXD37RPUuAoeJ07vU3L6wVNHEyAAgQ1PKHr
8WtvVapCi3Z0apD83XIvVYQWqPPdp9wACW2Y+dodeFMBmiN2mEnXger0VkOySvMV
6xWmniaEHr3oY2jluXSB4f3z5JYIcn1j+e+KvX4MW8yeG05tpI8v4s2jauO2GgAL
gRu6bLQhvunrnRZ95S6Bg58MPs4YtasU5HfhH5gDW4bJWgso4nXncNWKf67ThU2U
hVVnUaRez0tGIXUPfgMgG5xF357jPA7+g4pWdrb2BCEc4g/fIKKehzaO6BuLjZty
fNM19Ij59a0MfpHp6mRTGNb670MFsa+Xz1MmMTMCf4P4s7s3+jvNS7MHt8mkiuwV
XpQaqN2bboKoq3/OZ44l8KA22cD2aWpSco2Jv1v/lTR96TU0rgx+h2Ip7rFthYW6
0Dc4CYRt74VKdV6sDXhLZ07i7lC84nNWbsYGPsk0vvtVqxG5YILiUo9aQNdrArRS
vcEVHHCR8C2Ax93PFc7TnaHyEx6rV8aEEHn5fnebfcQBc1W3O7xY4wG+ATSyKO2C
tZ+n/oB/fgs0isJHNHwbEG2wqnnshI4Hb1OKEO6xSOQBQr6ZUzsXIWWfwn093tnF
0hrdX9ID3sPQUmeslQVFg2MUmxy63xeeBX7B9HFMq3lSEuS8xrVEAKIRmf+1Mi6B
OySIWdnUV452q99kgGeZCxUwimOVNm7HyJHtgmv79CS2Cyqk0mtnrl7C5EVXgSbp
0tNssCd+YqWO89Z4tw4e1gm9346//Nz2GhXw4ngxim0wmMJ+0wWCZIpdxLvxQQ2Z
/Rj3GEfo0hzJ5Mxr8MzOoXTtDuOL/1Ml3+y4XICL6Si6h2mQrP3tPKmFtv9mnu2q
aP7qeAnxB7CADb91j5UkOt1ZSjhJvZwEqgShFCtJ1wKQsyNcGBDzf3icX06VTok5
uHZKtlm4A0ldRpKOFiEq9+KbV7MH8fBa1YtW5rehrTk2sflsmSHeaWJQlGR2DGPx
duQy+h0GdkPyr/Sdpf8e/B7iCfNbOWQEcO0B6OXWMdO0M65CvJtdF24HZyCKyAUl
hcaSgnN7VxtKwZpg8q1BxzH2U3P8QOYrXQq7Qqw33tX2yeYCCXayjt3ZAVdCCOKc
RTNgfEbMTvR7cSvjkj4YlNfWzLI0ueDmH+TcWsaHpn/ZhusSNGfWgsHovwwPZewk
xl6KYpG9kFhoHTR0u5sAgBK8uhZHne9KrwlGTPuDOp25P8zfgmqBQKFtpnbUsL8C
NETss1qTu9XfwQSyo5cgpYCt5C4p3OYA6FNMR19uTp4cEYw7sTKYlhKe3NK3c0w0
f83TOF2l0fLesvbfij3CXhOG100JDRUSxdDPkykwv9sjdIHYP0wxL/qTOWmDdYhk
5fjb40LXhFNxfrM4H36yBgzQdcra2VbubCpQjefaL6yriF2aiOH8K8SQ7298p5lj
N3OkRo/+p6uRXjssKbGXgyDQybORBbFxw8whjHKDPdwc+mrBC0/033Gk+7SF8Gpx
N4zp4cfXtVcRZQ2Rm/B5SMWQ5JR7xcQTeJD8UFGkekp1AoZW79Himgj8q23VBeYM
aA0J5AlJ3rWxUfBeI5VH/n11txy0R5t4bNCDZlEGDyoqEztvt6YILyAB/KyocZAj
lEWVGMpkWaIy4g1sr1u7+DdNOlFvlU7wOSeY3xcDjOiwo4vfnaNgzgT1qpAg0aze
f5Ps4zZPE3dNccDpL7FG5FuO6v3SjGPAOosN/st7CybJFPVk4A8ny+JjRDw6XGeO
V2VNHQSWYxYMkTQisTsBsyyvxZU4nDYcQV1iJKeFpWwQ//9N9vRE+Y8ZgXbKHbAr
eobq1pp1hdzcJf/Zo1xtzXcWxs0d9+sqhPXkD4rPJUk2fcgRB9MJ2EFlAnLXXQtx
MG7qqwES2YVLKCUqcsgzmtMfryQE2HC+wJC2f595HNJpZiwEucT03J1PB3lGP/m0
zGlnvaNsr/2l7Qaqj5ZSZv/GgwGASNNFIQI2Ld5eFeVrSQzVPWbP82nkvfrccEO9
LzKMN5a3gKyx7ww2U7OOv1qvPAaS3+1waUpc0ndH0QhY9KUsQFtSPC6rXeXwVmUh
sG6nCXfpJ7YgZwDwGmvCt6XfWKnFrGWlgjyGJ49ytb/ONk2ZFgKeWvPyDnYc+tf8
M89EPLKQnH0vF2sQLzbPI72ANGOB4wBM7VdLz5IFyzLzc8XlApror6B7hiLesOoS
mbfFWZgCD85M9+FFZUlC143VbtbtQjxn4sGZXfaLXq7m2bO4niVMnpfghvVB49xW
QrSuR1lKfpGfs2gBuDjZ3XPHdig2RmkAbYW5VXxd1WqEIkzYsI5Ik4aeicGEys0z
2QhviCaaNLhAyfDNvWp6os92oLxzOHRVJcM0nOTTzPaOna0Zpk/4k/Td/RlleF7Y
0v6ayWx9WpF2B4ovG5863+CyePcl1kx2VPhc+c94I2I9Z39eK8TsovGlCHIU0Cb/
HpI7ZEY50tu4AuOi7l5v0dCx5UPCuEExovQcWq/+JeIMlOkIlM40z6x8CCBgOT3+
QheQi4bxwJrSqBv3bRS0rIE+71uJ/zLLjzEcYxBBLMgb7Us984YSFc/o0XwvYkgd
Jf7VwkYWr3Sti4nKqXjnSLu/0utFM4XOXDVDsDXgxoOTIGblbStXqRpwgIr3R4hl
uyvBwZApvZiH/7Soh8Ixxi3vKbHIJy/duxQj1THYQfX8z3lMdHEdQyU0yZ2i9Z5j
weBBflyCHd/EdFnPmB5pOjbIS/TjQR7PfbW7CRCv3XHYTWaPyr7GKlmoJMSuP4S1
HbGAkTYQgrBsJsgZmSlVlJSTReRlmM1LNBGr5+8wPaZP812Fa6UGMCd3VSrWDi5d
jEKsSfJsbKK4ambXylh/hfMbXqrvSZLc+tQsiUwOyRyPVMFqp/CVZfteqcbZhUW4
F3s6sJvJAb9H7XnG1WiQqg8bex8d/xQpTK6iWczbQtD3uHDtoYhxxhOY008JTGeA
rjjJrqDqa+XiINZ4ZTp0kP85KPZerod9cOgyXrKQy6U+G6eitgtr04MsJm7BByrK
ONKoxmkj6tp47xo4Y1jHUxEhkAl+uP8fl0FaO/raLNb0LfUHXjFLUMW17YuOi8Ib
vQZUAE/iM/NnP7NXrIBW1nBodAAXy7oSUDHT3kxybmRfdphkJM72Zz19qF6pcyxh
ZLt/YCM1NsqlI+zH6Z+tFWojLCDdREXKPDGr7uPU2x9EGpWqnyejmFZTD/gr3448
TRimj4J5pgmKozn1oPxjzJlyJlIQlqmFUdPPRbYUxe7pUIupqjm3c/Gc8G8QBFq5
ZRLEjBab3soUfn9A1OylEX8uear4pVYvfOqNrqLlVWHXWERiWWcEq/jjNCLrkROs
0/UMj3QXDASmTg3XS8uKQFzwBYOqJUDQ8Q1CnkktcAYZ9SnyDrO1C1wVs4qopgFW
I8e7IsYNV1Ao9gGqiS4MiTgvXvyoP0+x4nfYMymZGdxBLmmKvBx9UiRgMFQpySs6
3JNOU7DyEiETQmMpBMCZDRQYap8ie3drmDx2KI2K22ayrDVluaXL96XLolBkAjVB
ji9NukTKursDLud/hqeg7rgQTTtll4fFYnj0PBYEKtn8kD5IPwpEtveiuAUnqAeF
1+jPgit+PLSJF05UwBriu0bECk4p3rNGtQAfw6UMfxZqCnW0heHKTc7Unb67vDlP
HrbCuUVJvsHWXNkjslAJrodY7RkKKiRg6O2FMjlsuUCIXlmetggQe+Fy0csxy3J2
bv4J5Kl5QQHyx6EVhWTlow5g1YBi9gvcZ0EpN9sJQksA6zNOKwNpJx0yT6mZAPRu
rZimaaETnKUEh1Zhqcj+WeILpja0+7AO73D8dU5XkmmCgapZhRtLCHB0H7EKp8r+
DOZYo1lueKLYPYyuz/Y5L59tY6q7kVOUQ/8rog7Ymum7ARWhU87bH12vtEa+9kG4
BzDITSitWdw9d1iGmAs/i+iGOiDU16+MowzPmBSClq6i/P5Pk111aJ3S9Pf7ul4c
NTdRCllVv/Tuk9ok6TWBpt9uldeV8updO7DvDmIuDLZ6WKHDN4bvCIBIXI+bdL9o
b9hVEPXFN38LDsmA35aJ1tegUQZutT9o7ZHpg1ev3CDIbCtjtE0u9/3vFcoVjqvj
Tlnj3tNw+owJB9nJf5GwiMj6yLQRfSY03vyuc+xDuuOe4TSM1ACgI/0ohgZWyZwl
a9fE9QyZ0T66pyqvascuBydtcxKAe1jHgpOulo6oi3wYYgLoyu2JZ2XI2dxzntjW
mEaU5It90UUnyUfJywZxlvTZmmPwoXXUI9Bi0AcAohRXY8ppN6S/r2sVu0o+iKH/
MS+E6ew67Pq4XCQmVUV1t3yqZKbIQXYwaJpNjT2EdsIlaUct4HMejD7qxwam9XLY
SkMb/jQkff0s9NUV6jISfC3US+YyTEbYEvOkDCdiIQQtNgGXuwN4mgl2ZY2zuhno
M/zZGtLTTknhp9v5Z0VF8Ygl3gcNWB5L4QF0XZ1ewZ2L/Qwl4Pvdy9atFnwewK+D
TMnqi8LfXGMguny3rFuv627H1rWJJWbUIsEpSW8Z6vnNoSsaV05cKeSVvMM49oNy
LuKD7YKmhCVv8YgLF2nww60+TkjGbc4VQd/7FG4pVQxkNUN8dOK0NrpGkotXXXJ9
EWKzrX24jJiJhiFCvzNQiggpPUamWjdUhJxkJh7r8fQ+QY0JmyEK67s7jyEMjdUn
LEO2S5diGY+odwfd1g5TEtvKq00YyPZHanp6mL6c5fpLayu/AEL/ON0/47r3vKP9
p/rC0zpisRA7ZiS/T7ZbWEmYrgE3V20R+mWqtFPPeZhEramwUl0SnKfLt2kW2lQr
hxnPzqUrQRIj04/8kPlRLpd/29UxipuT3+KZlvQ0MnSvZRiSguOhC5PDVizHDdco
tkMoh0O2th6idei93JErAKqB2/JrLdu/Amg32oI10a+MiylUXpSagaE0bHDHr8z2
QFhyUkIVtcYixN83d8V+0zJ39Q+I/sNK4pW2gjg3X05s5yL5daOHcddJDJxNQOau
CJbhd8QP6CiRrBKlrgrft7AszQHBHij9EGZ6gcPDVIO4K5OB/MOrvZ21jVV04djP
fyUB2/WyiwifaN1bzubxdfj2BFkHpSrVyH9y247t6kJ4GnUIdaWinlh4gFUh7Oci
f/xgAw5dkJBq8J2AVYI6Dg5HLzVhxAWkthdjPGjTSKuB5QUe7CkglpPKunX6wa+n
R2i0yqqFD7XVTKf5xFuWHhs3r7BgGthlKIPpQnvbGJGB5s1nmu0gb7aZGyRHhLaJ
zjZaa9K5Vg/DWNpybGsukkwlt9cxdFB6aBAVckvold/7yTYWmWjXK+KgDG9RBmX9
wLk/Ph+ZLtjFrdqgsVHl+jIy/0CdetknMkgWmT2vmcKTln+M2FZC4o5wFuPgIFIR
3K4RKSQbaqSgYOM0IOcjZMZ4stS8GFlzjBWPFQ9FLGFIYJgk2uZPfaiCXTuDpxEk
rDZ76hhwFHPQXucD3MvoU0jAblGjL7+Vi6BW9eQQ1XFszYz6F1iklrjssLeqikoz
JsJKfzbiBL8HO+9umuRTkuNJCJagaPwmtambYkogJdDMOzShAR9ueHsLVFGTIUOf
eWHmaqRGSS8r8ZI9KqDzpHyrPvlKmS5bQDVwaNBeHkpMNM2RFiTcH7ndYZWY9sGa
DnCOiXIwAt0qL3+dOh5DxZ6zaSFwV/Pfi3hSda6QB1xtZ+Jk2+A6eV8oOOwi3d8y
zA7GBNkAduyJ71HEtRR731Z4E23O1l+pUN493cnyijwU719D/Tg8jL8fvs6ySBWT
G/DFa0ktfQ4PmqwprC9Ta8oKUkaz9ACacl5EZM8DJlpnnmZiKAeEdQNTuo95srMJ
GR2g8Q5RIaKGEOYj5lWs5slCWDnt55K9IoImnzCG0ZibL0ZNmWW25AddJJtJw1Yf
6rO9RDjrimxbxWc0WlgOR1PAy0thxwE6uhTqwl1sKvYJFxoVGEHOO1Hk7GTBPSoW
hPCD+wirsN3ONMmgD02u1qNx7wGZb/0WOvEBUgPPcWaJ2fzmPcuQtMIruPgd8nox
Ne/JkAOVMceIEKnBHMnZ/Pjp8Nkvi0s7eWu/ifO2laKLd8p1yA/tqpEfXQqpWbh+
BtK73SS3vClgjKqz8tzZUszhrsFUUKNu12/7j3wQwwUslS8Z3LXl0xqb9nVxMC6K
4tEjXyXc3zyyYm9tzmc/LqdCrlhlMjMiGkRav8LmyvIx7PFPR8aGK8sQJNLQQbWY
GUWrOYkjXlBIcZ6o0ToyJbw/w8B+t/8S/A259WY4bEQFpFTKjxjYh4RH3yYjOrZA
RgU4OXV6/hr3mIXAJUFQditvKVFHpIiDc3X5LIJyajNa4wL0Ae6Rcke6rMsJLdng
w2Q0hdt4lYHLbvSdH0FKDV4O0wg+kRlyiLD02i3X4YB4DMSVOk2lvzcWKTO9+1GY
ZFiuFEM3SW1KNtDNHn8bONjPsnMNJhWyaB/gQECs0B9STlHnX38EjHhHzfRuTRbD
HHBpoXqpiN+AM/SLph5UEzcwi5PWPG24MvqWFbAOTRwtjykhVfCPlAd2B5ItMNCD
un1hI23r5akzyA6+0ytS0zBBSfyz8iVqpwNmc0FuLYEYEz0csiU+kSQUpx1m5xHk
CV3bCAlStycaF8UH+hh+/3CnoMRbq9OXijSkle0cFPbk7ThL2d/QOm9OIVMt97+i
ythYMfR6TjL+ZTy+i4cKEUQx1SMRzne1GHh/Sm9NHqbmVjiDhsmzWIsaJkAlBb3g
VCuOFmN0DbkDhMO/w63Nv9RacZZBmNKu/it8hXK//Y5GB1jsFWXQF5mnNW50B6u8
Ox2qlXx44mDa575wQXEhmHF8Np96YM9JODSJU7iCcq7yLL5LdvnfOVg+/zjRJt9/
VJUecKsfSlKB4bBRPGg9FOw2eTql3ES50Tges7LYm5cHl+POyKan6b30otwtEbCX
e34TTl3OiSQbP5TqBpq4aBkw2nxc+Z1zRa4C8kVheofIbf3RJvI6s0Bj6W2ocOfi
hEfYLAO9IFBn7r67oCXN9IxoJo2HytkYjW0bjAsNnjz/GdbI+Azj/dIbn2V6Z/jH
3apzS6nL1+S+ErKf5TQghNrGK21t0jrcnrmNiP8BrQYWCqvCKM0RMuVMwIn2sReD
3c1m3jzm1BSQATCTnIZ5yMhS56pfALg2X1Zl97F+YXSmJWPDNMcgpRTQd/xFht8K
yXBFDve+QjRWXuRpXcL1Z51t9IMLFaVgn1lUmmof7+eGxGcqXddf99ICiYnGYMZb
BpHcOOUlB4NqsYHDLnWjGLLMvuUtSFk3QiR6KD4aqn/pgCm2vJqrT1R2sxaqhwLc
V6cL0fAudcuohSIg6Ux8kinY2xKFoPdurQ/TFszxU90O+C6M0DHDnJ2PtvKiK5aM
UBQMFPaWbHIVH87u/qXQpKSOmfhVbazOP7sSCHov/Qpl6EMx7eIEFpEcxrzFMT+U
uffvZjzYjnQfhJn+t2r7kOdqsxhgu2iP+8bGOMhsYlb2dP0A2kQWHD+0CIF8rtKk
rIKKWJ39YCBl4M0La98Jo+sYk56o25TyA94ctIk7VqAe6dgcfB4jEh5xOzz/SHs1
N0Kwd8lGX+uPCme33Hp5Y83Zz94vAXkphYLNAp5Iy0RuZQQ/JDTYY60y4hw9TZKV
hiTV0HzJB8TGeZvoMHNyXiq7dsw7be26wRBdZO/R3xcCVtIrwpbXniQv/zCt7YMy
jFImG6TKs7Um9nE/JakD/OjzEsqNUudaS1utr8oVu4FNvGoCwT82FZfOpu2TB5BL
qGZv4n8Aed8P0vmt45+wm1lnXq42b4MXMO08qwjeqa8kz00HfMEt21J5QrkBJwq2
J5JHFSQITspIC90WZxd5krKkJngFnzPh7D+pp383ZMtR+KqzK6u97Qasez+CzCB/
YC1oiDDpXNU5wPvMv0+WfqQQ7836sTiG3U/QQA2zxIYZZatCuxgHv/s2/JrJIFS1
ZMf9LOqGNVky5IzVqZD10UJEzEW4odVV9vFLFRE+W+kvs0bbLfey49hSIJjj3XVF
hFmbd4oXX6jHJB+GIz2lGXQtis9FcBTdjDS+EnBIdNZ7ACsdh7rsoJ+2sTtOaJDi
7TmGdL3PZSPn5b/7cMK5CEaens8zwWMAJ6F2g9/hgcSIm/QetUITstZEGvBKtphT
LX4xkaQWNknEfc6v8nd0RNP4mFDkOXKkAjiy4goGLTodhgPBtQe+lQBUHq/k1nsn
cIt8vGoY/c7wPUBYptA32pt4Vq6VWpYMT4QVlMF2O5UCyE4XgTfOZzYl9l5A0bPm
/gzf+nFOefOTGjOYqn6tT9uA4UksLzCz1isyhjcrYaCN6lR9IbxOyMI0XK9bfxex
nLYxOAP9GjfPzHjEptbQCn62VbzYowWJak0rws8BJY215+YiF9GIL2pS8vz72G+x
redoMUy3sdIbignwnyuC44R/UjYG05caThnSo8T/sIQJEtpzqTzY8+j4KiV5JwDR
zOc25Tj0FkLLxPVPMoez+tXg/JK+lOvNA8FwH8WhF+nVny6afbDfxToOIhfD3MGF
Zd85d7h5c1w6UJd8Dy+dmj+a2kYIkmbSkmIOk1uzIjVkuVyEQNjBq+dNWDaXa2J7
M+RP2PoKYo3AuG9ukkvwuqMC82yh3Gakh3mm4NcXNLvrqlP1oVeGDCHDk+k0+fr5
0L/Tu+FJQ/73L2eQh/jEd8UJ0tLeCc98zi0LgiapPjXHDQX17OkiZGJ+YHgZemvn
uCL2myq0QuxZTv7gSYKnH96ussu4wwRFj+lLvSIUXRIFyvqARbnJe+acFZyJMbdq
k66f2vwAzSrZEF9azfPtyztf3ZBs2txJUFmeS7ou5V6L+OayxjdVTUMOjVRXoWur
HiCzo872v2oPu0S35haD2t2P65KATy+BZ9lQUAjaL3RVLgzwfITl2y5hYHLj/s9o
2GXjci6a/hCEMsAVJYEZQdt86cgMsBXpneMGwgzdbJdsnL3QyA5mpubBUSPZUJik
39OZdOonVN2bwFPiOnF2ooJH5ex/O7w7Nw4hBD+ae8lCCJWQrWjBmKApr/eVG55a
6lSnUF1tyArRBNCiS2W7olVsk1NMfsLOANMdWUEW7fglCGdieGOis8KFTn/TCu1p
XtFfSOQqirQlx1xQilv1cnnAU2JkXU8FC+PAdrcnI92uSEvwfmxZNfwezhWC+n+6
U/9n3b2fMryl/G0V2TWb+OI4PAki4qOARRjuHoEGwXN/uprtcs8g90hbd5ds7OMv
cVAJsGI7v+xbluGNS5Ce8EMXj8XDe1SfLXdBZco3g+ea2QhYx34J04E9Bx3Pr3op
0oHUZvpBRBpvyPIx7LkuMkx/3fj1VhTiIl6Z8iu+eyTgQ9tXQUqGZKxPTp5vf4R9
Y/ASkvIwpCKLPiPWWTKLfD5sWjxOMKdCsm9EGxwjNbZmmql9nDvDFUliWstRiJ1k
RfcP+mB8dcJF7NBr9bit8a8pyCDh/8xNfuK1Z182nFYByIWUoGh4ESOSC4M05umh
4Ag3ua25BocT64deyH122v3tD2lf6SCwJLbamyC6aKtazBBqtC8Yo+6VeP9vZMAc
L6VSD6HiLSVkpTV3E3eMS8V2xr4J2QFn8VjUED4ETSH+iAQ1kZpEG6SzOlWh7oAy
+vJjADz+n6GO+oxBuyuKR9KVf1gLi+SfqZMS6ZqYIFS0XWHQ3FkOCmduNG/rZsNh
LN0o/iZ5a3AqKbtOXly9k9zVUoFipU6N9dOTvN8aSNMta0rjOWV/K6Xd0ywtqoab
8GcnNi+qiTT1xugLozY2GUCzCsVaJfHOGXlS91HxCzolKROhjgu2Y2aIQuavaMuE
7fAz/FM1/ikyq2xNgQCchbTew9sy9x92WVHgv7wEbJqY08/Yig1hMLY5QrxHcUXs
jwIt/n9qg+zwufFi0YhRviQoVtJoL2tyuZd+KQrBFdE1bqAw/U+7ILiCXZdWJJBk
xDBAkOU2twqhraegESd+HRdNc+i7g6+X3gnjybCWsWT0h17v9hqFpqqxGxMfLSRH
Nfq9EdHisqwi+061sdnjMAQLMHzgdqNi9v+ylnCSesi68E3mMpRWxesXZMQlHqz6
2lPM9a17irESrkKXDeGV7LIyVRKRuZcjsM5JDnlCcdbQnbrNLPTphE70HVi0gs3H
NQNgpSUw7fcmH8tgJZvqGr+AR2hmJ+164XuHNTZm0EpMDL1IygAkc/xPF2mmzofQ
7M/znt4mAOCOcRHEe3wNGiAuwCxRpSqN3wFqPOvXHWVJ2Eq6oKVZXv8OogQLjSvn
nurzQ8t/DrRqtLZOfvZjE3XvOGRjtsmihJRap4hcO1LGK795eBwsrSkK8Bocvj2v
lJpHVUTbNW0mQank0K8Z9DEBWcaSAxcBNh7LWdLgmKfJ0n0C2DVOyMjd/HPmosU2
6hHvH3Sz6bZGdKoi3QW08Htqf5RNavv4gICr0L/SkxWg2KFO+LDJWMJ2i0xnDuy/
3S5sr7OXZ0+rvsnTfMLu4gxcJtdPATouPoPF7fsHSVgph3z+65LERRL9b1uGO9ys
n69DoTJYZROyPBJrggs1PlsU7lfr68ohPqc3HBhgVa69z2u2ko+gUF5fpCSrfZWt
Ze4yFyIHN3yAidRtCtn4DrwkdMvI7EfgDlE3QwqkoK+Fx4VI0s8u76EWnpbnoZ4O
GXeKtGJ3qY2QIPxkeR3TSNBckX+uX9I+NoviMrtWz6QG9XjC8QQgTWhOH6phN8ZC
G5k7UmNdgIU2pld7V9GpEl8hr28fCqvw4VcjXX72FJ6ZCac41VYf2qwK4Ut8i+4T
Xk4uhi/G1511yaLEDApb5VKLJ6TG8mZzZHLGjAtFOB0X5nFx+JvjVr8PUQaJzH3x
PpDzxyXnCQ8iAoNq8D/7YnvS0NOxSe8PQtkmAdNO7EQgg9wq6goMIa/DSMkb7LdR
u4bm4MlTyXLYuDKGC0GPzaW7FhavlyKCUZz5Ud6X64grXD4Jk+0p9bmeJc44KXBp
lUA3ZYMe3ODFKLjo4EPn/XMXDd+1TyeXMx/fvPKOtM6sXf3aEqtFv5I1igobCJY8
1DYf22zSdARNjeHY38Qfv6u6szryF/0WO7sQgYkJiMJl8dENp0nginS9ssjv7/ek
/nJi0Kx9PL8LtnXNh2fZaT7I2Z2bJGC+JS6cj0aYGoeO1hYcRSDXtPjN2+bwT6eG
jferoKkp9kXzieOn7rqx0D2Rgc43g4zexRHVtyfvqueKlyLh/xqRCrX4lz4k+8Fd
rNzF96zrXCa/ODf/iABntkNuzsE2Z1ShYURf1mlIi4OXlBejz5DdKncUqOYknnKe
DPcXWX1183RtLD7xCIGpRJXXJX4c9GAWpqQO1AQYG/zZRr9Csr56ai708ke456Qt
QnPVswIQPzHsGMfuUj9qwRiZ+6lY1R2DHrYbo+x70LW7UFYBwn52MS8OG8ZMvpyj
IoIbkFOwzilUTXR3wiVp0So6JYy06JQKpmp3zPMGRjvuCbT/rzyfgFf7tjNcPUxA
sYHWlsjOIMok8zgzB81iHUA5UZ4Fjzm2GK7s5oLKylO63mUMiz/3UmcfEddJMJUJ
syiPruocqV7ex/IZaQM8wbrGy1ffT6CC3eWZh886S14TeJhreThqK48RfmSkOWpX
nG40GPf78ixVRa5wWOSoKMRHAP8ECoKRIfszIvy5jkXVWYdHBJM8/32OAaw7T0ym
mc5tKWj56GqayaBpQbvU38mzCTmtUNS99q2HGWc8nXyhtFCGXpmeNE0ZX+v85Adx
U/qgo/UB23TByN3akk0fWK3N8trgQHyI4Y3Sas+V4TEF96RyM0w1UvGIdsgUDnlI
IjRRITDOzQSR/fDUaMoTEfyfWdPWwuYih43Qsai8VvKpDDf/CAyYdpMcO4N41TCU
FU9oxHiZ/U4LD30kAGyozoteeLk5fiWRYunjKIoEqfXz31Y2mujpZTAf/XG5HvFN
eQeQEPwwcO99rozTCBpFBpv0SsHCzGZw0AQ06xrpeSw7dYp3rtbXIaXGsuajk3K+
V6yxaB5Vc+ey8I1GaTwV8ChC8ZaXDhnoQSI/cIMX470/mdHrwimnNqyl6ftuReWJ
zXZawQEDdQl0l6blfOIa0sQRZYmwQBqZDhQHpD1Q9FWubt3UkFXplhCu5rUEuvLj
fp59nESGOCpYBJzsvLDIInJRsFr/BTvz5ByPRfZmyQmYM6fUJhsgRMfjqay6WF7N
EfHtLL9gJEFHDaRtftC2Ue6kTzbvoNVfQdMlYPvi8DMrGmf8unnnVQhksUT0FZHm
440RnCmS9rVaE7QqrEG4+mGrxL8I2aD12B+wXIMA9f3aGF0RYGbijJ6oMmdd932C
y8W+iXQnrzhgSi/hY1Q38eDXGgSvgwW+O4awKf8XkydLP6yJ9Y7Lnjl2L/rbHEpG
qRsNpeFUxUUG/mAttbIcdvx9bf876dCZ4NETFMZAZWC7vh9Zpe1zV4cI+msqtL8N
WennS35Dib5z+ec4vT2M4Agm+JHAb3vcjJv8wnbQ0m/ou+1rYr/9KKZnhnfFp77p
91I0LZm2z/x7MrBYiLjdyRqYNrGyfNNbHG6rmV4RMvwTvMF3d+r3Z6LkY/MR7BBo
rJ+h0Xmyn6Jwpv9Q1N2H5yhlUbuolzdxmQYxwK+TPvaFBHpQeGGFW6t38DMFVoci
d6JKtWx7cq6JamfD2NaGl2fzqJ+xI1fyd6qxbnu78C6oEw//R3xBKX/3tp92BTfP
5TLW929i29Iho5BtrOQ+fHPupP4URl8Ozo8owX3E80fj4BRkZobnfClhb5aAGpvh
DaH+vkOYZa/FUUHUj5+nRr9WN9L4v2P0eLD6uKsWmg329w+kpG2s1XaH3tCx7111
KIpXXdc5IsMPTZTxfOBhmBO9gLOYZcLQrUJ+Io8RLtuh4YhcUstH5gYrBpA2bgb/
FKOJadBRdkjGQsk/OGBnQqYXbBPOi9DMzrPt3yjkTV9EyKYDJjtBz6uz/pPh59sW
A776sFle0agARsMP4Hlsn07PS8a6cwzjLjzCdb4T+6XiOdKy4Hjs1bY+6DiWECeE
AnBV4o29iinml1dpeyJ8cFjFLLd9zE4KWmO0weW/Kz+rZ+JSKLFicLWinIhIusni
EPtWrk20uRT9xuee1R5wcMJ+CGahJyBiVUPfN885Nfw7//NrI/UiJV1Y4OM4u4SN
7s+Dm7Hx/FtvceBZAEIwYyqiIeyqO/Ol+hBHTM/1kNRK8DpPGIFNX+ApxP5uW5k0
wUxYTcY0WXS6HcDV8pbwT+zKLslXj7k3ht5JTfPDQF+1HdM8yDzXZlv1gJUYRHNB
mdFSeFLjxC/RDtBChXn6yHeo8vpwQCWp8a4wvnvcZaxeaCoSRo7prJ4jlhnRFk+p
b6zoOrYagrJO6rEYdDhfQv4LCMNINhtAsdXiVK15NzRP083h8nfN5rlOJIaP1K5r
zTRtff/P1slGmPpLu2WRH7BBnMotOe8UuokLvBHS7QIKlkVJYEapLWowQcel+hDL
Fjcbz78Hm9WIFEl2R3dsufKQQy6DHH2D4u2rRRPQepA+lodS0VTulm8bY6doLqT5
Gf1xtRgntzRjq3anqQWTmeA3uIWXWYQ6sWEJZPOv84wU4uvg6K9h0sVHZatpFOYn
tAmlM+LYqatuj+CY+95FM6d/fHz+22Eu2LNaqrQjhXpgwk+jYEKe8JISwavWweuc
RCWbRgYqywwlcJ5ACioE2h1b+kFnJZNtGYdq/qKNEWKMI0g5uedChPhHqY6SHMxz
BnjHY1xiX3svQ4J0q/IOvEojb4HiQ7e9lmzmWD80pVHsFMNlNQWkK7UfHVWYaX13
/lkDXw4joiaLpH0AdflbcNI1tT7iXOVY7clToigEPIP2bxqytUOZctI/2HQ9DpfX
r8aP6sOZd8zShq1UYcikjQEvgokEYQ1d8vxdZbarVJOqoHfaSMgci0LdMjrgYjjB
LzdttipSaVM6omgLFgHLO9FxmFMJ/wPo0jnwGMUK4WOdNygkQzA+CVS2uwxxDYM7
TsxsIBREmvgE5hvElIkIzjQs+ZKTyIojxgt6rsa3cdNrHM4SbMZrnGNoGqYVGdEO
imyrEhz//VumK8aD43fFgYWRjudRlmLCQht4My0SJidXQd9hrK0485yD1FJEOYal
Nw6vqeaK16i0T8ouQxf5fHaNL+ShQ7r23gFlr9py/9KrkxiuJ9j5Quyq2rPchtLU
bh75M2NKsWWL5Z0PpEgTHROlo4PBqAQKCJuPveDU6k7JbVne4lXxBwhRYI+WRbD7
51HeizGFEkvNbtIxf3PVNY2XlttcoGUBsOo/fOFGU2EDsC/nKPHlOnc4Dzg6RcFX
s1PunucNUjKNomgnQrutOcgg75R/UwksurLVuq36CBQDu6nmG0Ztk1qbc/6rvYTT
yonx887V+M7vvT1o8OnTcdjknHQtgZAy2WdYttSDfC7janLk1a2mgzVkM7iCo1Uk
ArhETl4TopYrsiQd/rrUri0Yf+4xmsES7aN4eGfFjzm+IBRkfQg75vSrAExWlBzn
3bf91IApdYmmnXLCBXAHxvqhUaU91Zgg7ATPgWoWSMtd7bShf8fCW81O9zKUbGpD
yPlwaA0+8STF9xCO0O5lEXBQKc4SqogZnlPGqwAzLrdgzjk9ehO5W+CRjgqv3Fg3
dHVdfO7ssm84jkljJrNRxX8Q7iTUe6e4Mb5nUw2/Ye2uQLI5Xm/kFYwW8d4B/q5z
e1iIxoELCJKGyz7GaZOsVGOsfAsVv2t16D3EMd4KfjlIxDMaj2NVDnvPnax2L8Lx
6F4dxPzDT15FPPGPGWA2dVtXUeq0NY6M1yEkoran5HZtiN+SjrVySfmDzcfAj0nV
t6wRn/HdxCbrnsczMuc/cWEP/g80vAd8RBRSeBGn/vVDA/abAKCZZqgc7FsvJbs1
c42UXqXHcQTRuGw8m6rghd18WF3+B8br+ADWmFyLAm/Qt0qBi/MbDmrtW3JQcdsF
PFhqZCFQxwv03buxNNBmaJnuP3bZU9q8R8wqimMXO6P36dxOidUqXiRZtkcUJ22s
JDzrrV7SC7bfqRtQ5uc35Y5CXKGN0rlglXPuZfhpOX6EzQc5U0ihZqUxggYlmlfx
h1Dbx200R19ZXPe1UyDS5ERAbUP5CVdY2MqHhItZF5v6x6eaWKOk4rvD8vHg+Wqc
3Sun+DMPVWGZLWA8EqfLMbQAWyPMi6kDe4R17L+BZxwPGDhewqINIsO1pnTWwNo3
MgXifrQ1MWI+VUPvKJDMBwYF09RPUkOc/BxcBLcR8a2So1nMSGxoKrkd4+ddFL+b
svzDAYHMrT0/mpeWoaeMinGMV9wuEIN10bfM99KUvxLM/pDym656nj+S6Pvl85/B
SvNTsb5NJFIHS/EyCT5ew81a2VVhhZJTfT/xzCZq+okztGl1GISwKj+Qg6EgEs2u
sL74/yYPhlL/IM9cKe0E4OScS4khpNZaxcGWlG/gPe/pbSjpFcbkKY+e+hOGJfij
6WW8bCdZ2yZWtgTP0i7/bBcvqhvBk5J3nL/+uubIqVoKX9tGgj+k7rZqL5bbRoeD
FHYnGQu/hNsh3UsWBymJDNvF2psQh7LgOP6cAs14OrmmP1jM0IL0+wZV40HxDxIn
xz8COv5vO85FrUrpbG9L3rnFGJkxSSM0zM0UmEEsKhd6iju8F/R2EBLZlMlYXhcU
o4Ot2hxcUfLrV2IN0uKrEnrvG1HpKuIsiIvLuf/s0cWZlRJiXdubNPktf1HKAZw4
VYWmNKciyXZA5JFkvdzZtGPp5+T9dcJTjHTHsT9tJJWpSvZ+IsmLu0/mzkK/ifWa
rM6HvHU2nBvC2G6RKAZr9wx3k7bUuIu4FETUyHKKr0QJSRKc0xEAhBqKiGErcN8o
h2X350jsq3VO7zLOX79ugFW0CA68v6my2wNxKx+hcId/ykWQMJhNEF0nwfzRoek9
Gi9WUT9Ie3xDe9UblQ53P/NeKkikWFZ/b6XrRRwSuQIBWbrNMLX1SNtUmzA7OGg/
g4bXkZ/B31U8Hqw5oGNOYwBQgTDWFr1HqXqdpb3NLRj/fZSVpGDVDmvK4J10Oxyx
ysPC2scCLV4zc6OEBa2jpvm0xI2A7mP1tcO7rN+m/2F3fUxxZwsJVdX7IJP8de+O
5LkuKV1DNOziMEKHLpr+tKZl7mXfk86eHOeSJC4w4ypmP2u0Slw2RBwJT7V8WMie
9AHMQJCKyvIjs3SfHkA+N8yZOwDBinCIiL1AyDfRH+t2z3Y5Ei1oVV7ZEbnFIG4z
/+hmw1TVh/Cfs2NWj2CGRMKTZezg+KVKqA0RUlTp5Hov3l8gjhjQY/tcIbTcL4zK
BUhH3bimdFPjwiHBcWJd+LpHeJoilPxJCs3qRsIvaL7fUb0IrMBfbSzOH4JlU8pV
AWtDc0C90YJZUOMKOS2J/DvASDFl+JRiz0UbMj+ljro1uzrwkb3uDeHIFnqyCJE+
u/4wUxJYhs6LJpQO1y/mfzNngesV7RS5fF69t75Bct/b/1IXmIhD4+pc9wrAkiMR
R006+zDDSZpcmGvrLfFEGTQPjA9mX798pDBqHFwRVnyKGZ+NgYjj5OaIzfAhWilt
20MI3nRBYvnMV098QMfVqOrInbqUJGghzR5joneXSnzOqHR1AV6BAIwB/TeqSWsI
ATpmwnmucT2eU5WyfLlmmBOb2gYj+ub6iu0WtNhenITbk/LRa70pxLewCpcgCgnB
gebzvKG0pDaoOiMi/cR9vDtnrbnvmVevRbjPiLfGzMDivQvTDBDXBGLzf/IMJzIL
m46/X51Y5iP4oXiaQXleP9hsZzHbxpwcL6qNxR5zlRvTV9mLRSH7Re9O4SFFp3LL
x06S90TkWzj/P3nsQKkM94w9pw4KFe4rlxO+DZKvM5IqzJfHOwub2AlNzuWjLq2F
efbt3LfKsVsaychglKp4UCkATsJuzuIEWqIMLalDyy16luXGvFFJ2mo+jEcyUDaf
kSDIH4e8+M5oBAPSkNRlJQ1quRRXEa1u4Rh56Ba5SxEc1sNAtkDTK5Z4huZFWjFr
Im9KZkio+c1FFBrZv1lameZsEW3ghkVB1r6Sbl2cR3J5btU80W0hl4m7nymLlNvs
H/b8zNubI0eKMBXF8CqOCCHDkgbpZkQ8SchIAwfMgeM5jqP3fXtEeQh4hn3S4kZD
jqk7xBRec+PUedM3vnv8j+9PixWkA+VYIMTTba+90qbKcjMLf2VRafOnKYWw3c+x
DuT9fTxgTd9sZea74okXFuBFXzg7h1whSNFI+bmCC/N13pxFxs2SIpn5E4H7oqZy
BvzN9+aiLZI4qoAtupgacgHcqlWtUo/03khDsKc4uRdhY0l57ARrzqCYOSAJxb/+
JrbOvChMsbhnc31wG7UiwIS/knCIg5R5qQqREMGwjKvpFZB0q3W1yueXLuN49cPp
0kxzEScXschjTnooaNFDO9uvmj7Hsn0YyVbNdb+jU5spzCC82hoZ/3oDjFQYEMqH
SG1vaV13H+Qsr4ujvB8Qln/ia/TFaE20hDJDWdwHvPQxuZ4seZ45L5DjWsreTDbR
zuaQ62r5VVjUbvX9IoJ/McX9ZZ3gw6X/aGEQ95ZaKgeGBouCSxyz3RF5QXsXcQw+
Uqh8gLQwJS5QH6qO2pOIJDuymRHIpFt95cWv7Lmp5fjNG9nGAIcHgttTgh1vwS+k
yLyyrmTCMZQ330XO5DZYqudK+XTsvecCFCrithzvLdT1uyvEPy+ac2hSA0m+3sJM
36v/YQ1eDdMfpxMZROMl10ruGFF9ydhDRxoJtQ4a/+OD41Kqmiv8IiaStTkqdtta
L7C5pRubgbh2Zmio33vLjtY2ohrL+HQyDMU+2KQCboqXeAKetbE3CWewlPkadYpU
aRoKxg3HSJyEfRd++ltW6d+jWm8R67MBNKVABPU/75TomWeE9YI84zgnDDuQ57P7
iW6qCnH/O3L7ilVcxRpKKdyRtZ7BtJz08CZbemkSKG8CQvzWOK3clPV6OPDnBl5g
7NVYi993C5xWVJjLJQ0KJDqdEUfjNGjr60Yk/vR32BAWMr+F2IphUo/S4b5h09Im
hu5xtZKxTsap+W8ghDh64DVuLkghT836yH/5mpM80Z73/oDajZJpUQMFAxDcP9Ln
vtbgYIdRWl9rtB2ecvFhz/nWw5k7o0WkT2LkzhwQSEZsDL0iNMy/4HgL3aEIaZEm
R9J/N+ewjNIJz63jyF4DI2c/1GAYsj+9S54O8FS5219F1K9FulPTjX/PbG2s2Sw4
ugm6murx9kaWFL/rQL4NKoAJoQqDdenr7YzpoQ1GrkuylIDMhMXIxiDKFK2C3ABa
7dlxveV/iGjOuuRUY3taTyqUaGE62hnYV9M5aoQXrINxXNF/XvUca2FE8slysp1R
wtKxXTnf9cHsO6h4ROaNLXOn7ljf1S70hW3JcRHp3W3WJhhkAzymJ2PQUM5Tg0ke
O3yGWUIgx43G5S1TWoJRCRDt9cm52keOreOL3Tjxis0c6TfbOxhthi+WcKduUA8T
CnyIWpJBZye8oquAwHAXMj5bucu0VvOTB6xiIBOtiy7l7k5ThEAOuWYmblwhn00X
agffq40I0bS1djfn5DoS5v8ri0sHAC5kd73/xRgsm40u0T8EDxGoNoQF+MA0Udxs
hScumJlmTkoidJO2Frt3nCFepCnkAIptjTAALQc9/Af5YYLGLOC9bcqls43d8Qlr
8vHF3VMMCJsFEUS0ZRaiROtqOfPzolgnrcMhvl6PRXTFp0MddcpxjFpbU/iT4nrx
RKGLIPb8w9g9ez1rnmj+B5ZHVtZjhz8TbtXsrsmHX+9JVz/pxdmqxNxMQRmpIVqg
LflYd3iZqmvv7Nl3ZYfYR9bijtQe61N1MYsgBO8dcgIpGzZBnha9nGmX3zEEwtvc
Dh5XcGrMVQoyzkNCp6+INS4z4wJwpIR87NIUa2XFngF8jdEcBodKybaJzPw1cAZ5
rOtxLbmP7zBFbYa/WeIgzSe4qsNL7BxPGbJ0wdBJah8j9ywkWbwZrKQ0RmXPo0Xm
7mhbbiDJcvTqImnpYRJdg5boKbQQmcOQShS3l3dZaMCrwBmVbujvRHJI0CuPUq18
IhI1z2NTAKTnWacIbDFwjzHbj99KFSv8iX7U5Xgyis4EhTrFoZJRO/Y7s4x4IZD1
3R8vXN6Ow9lLPQblXi/Ka+jxXKZhvM6P9zJxnwm95njyeRWqhF6QgmGogtqaxxF6
NnmpinmgFXW5MRWfhWeJub+CIJ92rIjh7/og6bdeUQJhXTfHAeyELykp4I7vHCd5
NhVXE9ah5oFllDuLnbKgT0m01PIcqahMUL0/x0FO7s5hbHeW2NxU1VWoIvkV9Hqd
eQe0eW12z8UABp8MfolgeuJHiMg0bpSzXprIVp1+qS/OH31wQgza3DwrvvEigRoX
n9j4p/eA1Zelq2QGKXzBEQ4LreTSkSIemOHL5DdYCFGWckd9UpsGj7pYCk+SX1eu
4cZ4nJF54JFPqzYcDeuIGOUg/u8xCazJ622siFFnnJOxMvQwn4t4b2hX83PDINfg
/eummMyi7+uLY0eVKfUqfnT8PPlcTwQBSxGdaVsEbyHOYiUSsCg+pWIvhMjkNH65
L3x8Hs5wJg+zmAjlMckdfbLUcgr/Bs9/JlKUXuSy007i1+PY8rXwWm5xMbmu/evC
u3664QoiIjF/IFYtsGCq3oLe4WpJrtKlwFjTZ46mNaYgqOWHHt6jAOMlRzV38KXe
LfT3EFmtJLwQFhRwjagPgOuwPuzb/6R55ZfSz3nXoWjHU9SSBzzJ26GxfcDyc13j
hmVm9oAH5XZpwGk93jos6EcGQfqpiebz16ydfcY/sr4O0Ju+W9SiSetQrS344w/Y
HFE6iH+9lchInpeHs4M59e5Y4edFlzZ6RbvnJZPSLzRjCXFbtgHmWW5aBqwAqYCs
iWUHbdySSTY38fAQrkH1NQDOqVlo0/LezUO3+u+6svhk0/41NooaI5kwKzdhOBbC
n3/H58y6lmkW6imgS2osp7wCy+UhO8EnPNz6r59rm6Ab1HuXHHhVoAKft+SAUPpb
Z2nH7oOuq9Ij3Qsu4PX6Pz9AdS8xBOPxP3hWUJOAos7ZA6XFlfXeEotSWsr5AJ67
Xn9WZvtUlLtKH7yQ5z1bGVRZbp9SowdIRd76JhuKv5QapaRX7DBY/wGjaCrtuTNe
G61Q4+Hae5PtN6s393LAdEkp/6piUtkSULW3MZvT9XUybzcOlTyeZoxq3tG2bOJB
gLGnSxyINwMf14TR+SZR+BJ31o++WGqJR3XnEcvnm0yKJIqci2oQznSd7bQBmq+Z
pon8j90KLkh1HyfpMxjhT8gpxxnIC65F4cEyoh9iV8EeVi0AEiAeKcY0DpEiuGFs
uYChtXTgfjkvmSEFkONWwJatHK9uIgDUD/4PQu4CaBDNvc5KdSD8K+TT/UaCOa+n
+ILLGfT9PUiB+ikTLoWx8R/h3RapQWwFGKBMtNlGRdnbXuZV6T5ABgZ3RdMfTima
sRYQhEFYSiaI22pTRHEJ7oGsuNmTnbgIAst43Lpgo/GFX8nJ8QyC/S4vsI+63Vf7
XE/MWS4qTMiAc/MXnT3Q92k7ZswWdJa7D3wOe+F1GdYgYANODTuU3+taWGjkKWV5
VIay2ZsmsHbpW+3xQobSwKFGFOaI4U+NE3g5QVsnsupaF56zaD9TTKZCngxWjXo9
z2LztLuHtdLAnQRDiqKNCL4BYGgt8IHu70MRmdsATXezRdV4YGExg06BzJxQTKVZ
K8T1K/PgVGzhMA6o+dcndZtzIQQcTf6yjM7X5Q8BII+Qny+2roQoUdELZuCz09m8
Ujio6fw0e5F+8vWO5deX9jJfpD9GePOrphJJXcJKTmkY+awGnjhxuWq86+NjkzOJ
K7Sl7BRMwsixfR//zmzRChEajUQsNHrCBVz3zoGBXx78w3EtZBi0BmEfASssPccx
3xjDlW4yJ0qk2hM+VSeuugoz76Z7Wvvrc+mE6d7RLMm7TrsAfFZ25q9uk7k5+dwU
AwcAS9lfYuniv6u/946LBhYs9B7qWA0y3w5EvBfMR0neuPofH6pmOehC4u5KFX+/
tnS04s7XZLv51b9WeJa2zcKfI8ppekoHktcsfccn7LQpJpD7jBz3Nb04jVpB7uJD
78/hHwsrzP//bNis6jpYXe+gwcvTtjL3VXW/evHgpcQEDMh1TponZx0OZYApsOKW
YFoSrHsqHEcTHyIlhO1nYgxzSqeccEHfU9SeaSUToCxILJbfCQSdm+vpKDrPb0g4
1IVX2/LBKtsast4pE1LgpYUI+9Lee5dbcumNlMI3xul6Xjfi6FtYC7P6XnSjP63A
NlnbhCtRVFR5SX9B0K+qRV1CoLMjc7JgCIv/GTvd+Sc4ive6YjvIQ+4d2jQtjQfJ
/zHMuY6v2GL8TkkGyajPOxMw4vC10+AotTY8EXyeoEoEEKqMl6ODuJ1qZeF17iEx
zgFbYCCt5Y5kK00nOmFK/kmDYucJOYWphNvBkf9c+a84k94h5eWhv/54YdyJ+3Pt
1R/XM8WZoDpUoREK5x4SaI5bJacpRlp1xAATt/zqHRiRpWUlbyiQZGM8FKTji/Dz
z/ESwVRtrmDC6pTU1wLZ7Vc+iX0Ub0QVjHMOBJL37UrVlk/t/19KVQZIZVipIaNP
b63wuMZfEttfmWUbdsJwyWHPSGunWd/H3R76fBUcrWJOr6x8F9/FIlxCL9Wf0JeP
SjSU2X0ib9vK1u/dcPTPjUw7QLgL75kzsBs2TRBnNMT3NlmQg3Af+IGZydczRJch
G6JU8OyBltC83a5TK3GWrBB1po5pPVK3YpJNi5hNZSe0Fpnis25bMLfL/n5ghLm0
Gha8fdwVyIS44AXw2m16tNiPnrLt9W3AprVkcVvI+JlOa8ReIM8AwEJ1QUqgOX5h
LniIbb/1QqAhJKqMs86JRweCQCclg4eDpy7xQtX8DZ1YJmlB5g1nMhF4iTkS+CRB
KIs66IQGPa3o2lHY+ZBwW2ZSoyG/ztvEag11W1hki5XynxNO1e4ELmtG4OKbCaDt
QwyadoBc1Y5timWTTPFDdDBZWtKnWkIHyumoQSjhrQPgRAJVceeJvGmEq9K0d/NI
B263votZxB3on/bWPZbr/RtusTxgziJB5ifYFh4d7pcFRIIel+XgtbfyOKfbN8Jg
yqePaPB6gdOMpz/xJmM5DXKgf8cOHUcwLgnyDYJzdmz2hupKrM4kFAQwB9rD0QD2
QzWaK3WylfPFN0g+a3J0cwaCvHGXyO8ww5QeoTjerMcduGjnLNiH3HSZfCJuCNcL
B82MT3mp6BmuWF916UmyKeTof8+mRRWY5LISYJ0E22rF/tVyzIsjVEqRF4o1SvtG
eUOQHsppwtVclsKhIq970RjFsnUlTt4qa14B2VMzp/nff51m+A9Ry/xDAWtiqRg7
P9XY5T0SZVNkpimDGUWLJeNpblrjlPP24mEys9QK4TC/LGaPZKLjeulfhuiZbiu8
EtUCL72v7RBWOcqjrwKMk2pCUZT0K+I23flMZhV6wFoK2WYQWgdjei6mBw4uqkha
z0KrplCrbV1c3NitRdzR7rovbkB136uMZfSgWRom7tXtrfx7SpRxT5eiom9FJJHi
PljsD/VbNfkU8v0txri6uCXT2Ci7QGewdFVd5kRTAUS+sZgv+Xru+Aur4LZfI7m+
IbU0BEhsMKW4QP94XyYsFvG2xhxtQF5frwfTl2xiFFM6zz+qItU40CJWtIPnbcRy
2UfiGmJnimVnS/LTRWGSmaFlSJmPBaO9nE2xpvWr6KTXiJslXUOLmLAlhzV48o5v
WPfzI/Lt3L0Q/wq3V19vs5lRSvvM8JSSVRrZE47hHk42L0PLLQOYURzZz18bwy5N
6+g57sfd+6GSMgc+DNvj9pz3e+p4CDClts5h5ZhxnKiAe5dX1fNlJzUYA2XHSdlT
CpOYQ5FsjwsyzHNqwElg26Cvk9/dunQGBNekOTOtTpiFWYwsIxyEJ+df4JfXVdaM
bLwFMPdHTomIxwkRgUHElyIV+JjqyiZZQLgQWawUfe73Wjjyj+R0f9NVNLCcbKt0
9JHHlYk85qilT8fbm3I7HwW0nxr8mjdatb730E9uFku8FCS9vvQKK5n86pQlhEY3
MGuFO2BRfmlSTbECDDkeUMrif6mxB3AioOJdMmucRY1L+N/s/xj5Icle4i3DSyO7
bHA1Jkm6lFHltEl8mZycSg0tRGK0/oBBVuHuK4yEk6Kt5LJoD+bw+Ti5h7zPnE4T
GuKEPmu/qeKke7CS6koopVivG98gD5cYbvD+JTnAz0V13xjSHDJVVBivT2N/CrN/
Xu7+p9efIwu0oAHBLKDwlaqe7vjklfUJfqnFHC0GWs2k0hEfUCPJg66SBKd7+v+O
4VyOkZ1dpmt2J4HWeEwudiBVZHackgMDp5gZOQ5W2TcPlDPLjCj42HPbSp0imcfU
bhEE3GUYdnflScOF4mj0uOKHHeucTX6tpC4c9VyuKCZiLQnijPT8RMczog4YwfnN
dzdJ6uM6BcDV05xtUo4WiI0SHDx6tjxaUHd6kxP515gC9TSD5PcdyhcefGrqNk7w
pjjOu7+V6Hbg70gNM8T0nCS5PYaEls1u9O1x+jf6k0RZvMK86JV7QxbstIepaCCF
qsbRi39cZjOZUSHEdpe0DoeR4HZm7b60t5nFm7WU7Lckhlat3n+04gznsDPOtvbo
i6gGN4ai1FmKbpnn6oUajiaEIKSCU0iDDy6y3WBPWFjTsdmsPlBnKbq4DfCZPq6Q
LozjS5cPfTbGNyWWDmPEbEDV1Ky7HbHEk1ifn24+emhZzCiFk1LhmUSSMwJkyLNS
F+ymEX8WGsKh7qKAycRghTtP3tSN6YSaPNtFxLwrjZXLk2Q9s6gP8ngL4CW6NKhY
4QRa2PnXnuZhBWgb2h7KBOQ/ZG4JAoPLYNFwC5omS/3EnLm7F9tIYJUP8ThbrjRU
lM09cF7MLMyMuaGgASG5EKh+fJclpLQOExhvp5s1LW9FJunulz3E9vM7fsuS6DXY
16vFYpMFoaEuAxu197GHj9LT8NYn8jhu6eKQTHPA+mDdpc3Ple0D9W66Wtu6bU+6
hMU6YrTdZtuMrFxgERU8rhcQ1m8K0OTyiXrYEw3F+JvpftHIxLVmsBYBBZcKMoFK
4QgifNpzvx3nNLcoCQCO5C5UhN7U5VtIuewy1cZta3Ux2GygG6l+pV/Rd41oLgAh
0mlJOwOnQkMPNC8ZvdCunmujqjFYHuzbRaK+pYUKsZ+fsBtSEYG2YB1pWpxVQGEI
0LZ34evPKjDhslhRZRL1B9GKI4ZwAASSN/4alElscebvSol6NV7uiVw/hGq7x4Un
QzwveyU9Y8KxZTr9Rzu+tTwUDs90ZQ/sDvO3Q7mhb1P49O2P1icLB7vl+ynkYePU
J2DvgLY6bEi/7LpzUtzWJY2+3dBOuWwsFGr5na+ipWbZQ9sD2XGJTU5zgOInq6st
L1bswqdy+rrZYbac1n1id7FP9gkc5l3L2nn9pSBrZEtauUYUO5W+MgIgKk7EVwrX
BCEqadM6TsgZ/N2fohmidesF5agKk57g7HJaOl3EUWu7iT/kPXAjDMvnYI9DmZrW
GEWGcaPp789kQtY5c/h1q9T660KXPEAcxwekE6GSP6raknXqYeJy3P5cqpO8u6vg
ea4sGAEK1yGqsUBQU3PG8x2HLFUbUEg1fyKOdJq64TfoPBGYcOaoSLqIJfBmFi1l
jIKPYuLyHRIMquxDLhPy2F6qp8hR9gec8aXjBtHD9qni21B16qkVgK0gN33cmt7H
gJ7Gi34C1L+snz3Pri6cjlfyl8wR06cXMho4ZY28NUfi4ocuROsIs7m0rBpht5SO
h9q2zo0fQ3Q5R4OC41bAynrexHOCDPWcgideRIvdtn+5M6i6Au25t7Ja9gdzqbdo
ESnqN+IVlE0wzmi7WvAIHcrNnLHfD27wE86xglYCGiZTmBpM1Z7Ti3TQVbKXjv0e
yFCEC0a4qbc8sXkrFJJX2riMqkIxsczE5pdhtLyk6NZFRgAvdjszIwYxc/YmppXM
ujxUenwRq1pX4sLwT5dyRoOkfbFcoQfLjx/15YmE0VL++SMmNp3q2+Lb/L9BqNHV
v1QNtcD0uYEO63L6oTus2SZUXQBS2FXAd5OQAqT+WNeJzMXoTTHaTDgro8YN3vWJ
dCsD5wHaxK/wxS+3NnHEpikXGUahzC1x3Ntzudf+aAQTCc8E6iLjep6L8MCZoZWU
DkDO818y0TpL0krT8CUVKAsOgMFUAnRovdYvzf9NS5JN7vhL0TW0ANqlniFQmQj2
kI22MCRO/hMyYgkvo5XkEM2m847UjL4ZkFzztBhPtcDdapOuobqoarCgSzpfqLrE
aUwClx47R2HIk46i9gqfstY1qwlARr/zeVsggX+qH6F+QpB9gKP9QmAYN2kuIOy2
nLs3/H4atumGr+4ntwi8jLvtS462Fe5dopRqYm62cZLlKCLGSiNnj9BXR/R6eI5s
yuNI+AxgLc5rKEOI2YQmBBJAcxACbPvp7u//rKOKQ9Sw3cqFxDCY4dWuAsY8Qibz
QWLv9qfZ1lgjXGF6ylk0PGTeUjI6AYj3k7hoyRUtuVQ1TqlkF7ouT17ntWfH7Xh5
nuFCrGPpKHUbNXoz0m/83XDku4HrALeiMDxwoGsbw7h0LEba2JlXbpKdbFZkoGqr
EM0KMdrcZJnzdqXnky4JtgE4cbvXnJwWv0b+KZy0kYUmFE2BgybkoUH2XG3lWIva
LsFXSWwMmSaYtlDZIrVkBSB90qowZPyfTh8xI46FwOM784Nzg/13MxDmdJTY0G4L
YozcPJZLq6Y58mtVWaYE+FPGWf/9mDcbf/Luml5OG1ZlzfySuyzAtupmY2lU9Wxj
PCdmFHDhUV07qtRzaFZEocGekICZccK5Bjc36r1CW/egkQVGpJpjkEKN7ROs95pR
CUHn/0RJxMOySLktfRHxsN812ECo1MNEanYpNEugnsxc9su53uQ65iw2HKj0V0g7
vPu7bG9kQySSsdnsOnA3bfx4Y+F0RJNzJTtMKf/PM2TpFnNifvAysCseGzekJIUb
tKU3SmmTK/l2cx0bYHjj4zNw2OKOO3lusDhgzCrv1mvfj+p4PgL3BfQrmBih6Vxm
a8O4lvIoiyofXwnPWdNLmEY2x2HuB36bjDXfoQZa8+FQFNuCB51/dvUyhJ3Jfwww
knJsYmV6v0pg7GP8xnJ2ls4Z65o5tJ1Yvg+Np4GwoRRBXxDQM/vfKPfhUpLlY1E5
Wjj9gymWER1frC8JpVGutThDfxWS70mnbMeKWddw9JlYe6Q/QgUFo9aJqayECsEn
ij1xarpUHyYPPtr6wOl+UsVqvkwD5CcIcxA5yjfNaYHe2eo9EQyQP5z+qHNnbXY7
wXSE7AUcW/qXrA1D3Q1q0hwENTufGIRjysUjOumRqXoFidl5hPHBkhJrLk4n9rEj
X/VZCCLwqPcyJSYg6apmxCUJy0Em2ls67XJC+19I8DV3MCfBsqqS9Qs00wDz2GCq
uzCE7AxcKN9ATF+WORh5dLaaORtBNqyY4nh/J7pwAa5UkOYziQsRfqL4Iy8Smwrp
uzHyYdLlDLZYqBScNV+0lSRVkG1BbYeYEfbrSqkcSEF7KdC+GzTq7dXf4vrsF+aG
dTxinxjRW2VxkNIl2UiTn1OIJWxamlmB8ksjBNWf0OX5qxLlDm9a7iJWU/oRgcXx
m6F1LC4iM7wJ1NY6CUkCgyGy+SHJtVJxQXOIvA0cZbIk/axcruzJZoTbX1rf13CD
UuxhrTKZFR71CCQOOCro7ZwfNCOsz8hhaxuidZlt6tf8S9qjRVxWfOV6k95gY1xL
eoiyHvmSS0ASs1OXoGqzA/oC18+6P6VHyjAaZGl0Jdqb17ahSY/AqPvSBbb3HEXA
Y9aQK2wC8ZUjbxJj/F4RVANet0My3LfTljbpVBgnBeaQUCFGwaeWUW8W/g7eJtCA
JmbZ9kGiTx2GUj4cFYfrEguu3hbb0Z0e1UAsJzHNzp44lFLEs5lTcuGVdUWqPJMk
cR1XZ5UKyjA60OVJyLDZVRwp5+I51kV8nVkkUsUXu0gMoTa4KhDsIlOMWgqJ2SeV
ujoyAWQu5Ak0hEPiBOcX+y2J2xGbfYD+yXFvB2uqam13cCwg6LRV/gPq8ujGQHh+
Yprt47UNjjbQAdZVha8BVQkBTIGD4LHezJKCs0dPTxx0hSIzlHW2crR/Mq52Qg66
qxprC/x0Rkgpt6+6I2EqwJk2J6ogiF9GrTjLNCipQG7vNqVNMf+vjAkmdUcqfHYd
DdPHBPM93oxw9jBqjWCfAHTSD+eWgDcJ2mSBARKx71kAi8T6l+ehtFJi3VIjQLAF
pXEhaEtwuslAOdDKtV9uircvCO4wN+hu8EwteTUXheUtq0pU1s7wA/LDYlOmKLNe
Q7vKKKzH0rklxj4QFZ4K0dYe2m3RmtoHY310tyznFKo6MLvXp83XOazThwtEinKm
sTYfxUVlv2Ru4REqdd+PUxADr7HudwSWB3L4PF8Ow3LoiIR83pzEzEHzCrjz0gIy
byfccTUK1ugh4tnfb8hrEov31iC75yR7CiuVuyXrTC/bDVxqTA+abe95aG9e4F+x
QP/sunMez6rknfnCAu8onk2FpVH7vJ4YijHnVwF8psuKTxEVz1OL/tbmskrS97HL
jdGIJ8w+5aHPl2hLVt3TT+XQ2TAqkqzLKKqWuY06/lGqVn6Il3pqDRvx1+ZU+Hz1
WIhRGGCEtFXyIyDwRHdYhDE1UJRJUb2EhNRUmeHWMKvTsbIzcnAQDWQy4Qbt3Q98
eIU1XigDw2bQXQHpAPA9l7+HkjkCK89qR/5Zz27lMmKIkzbpn8K6m/8MM0C+qmWU
pxNwLdJ9Q+urpmKqszaeTKGp3zqrNHOBppGOt/yYwfaL45nPoCvaY8DHDo+RDFb0
4lJpS/agID2d6H75nEMyOkh0d/eOPInOgOKGIotbGaM7lswbQlPubtElfyNCwF+I
EUTdKOPjzNwLv6VDotjFSAyvEi2jQ8VjhKersH0gfrgkGeRkEhZFEQr8FJPQgA8m
DdPOPFi7EEmG21++KvpfRKiAx3CgoQlEEWxwa4f92Pgllkdiqn/7qMU+1UlSZxUp
kx3uSaOztDHhcxczd1mJPArsiPobaCt5pZyVxdNicYR5b3HbiTw7novrfl+N9+NZ
yOrU6uV2LBV5hK/UipEdQBoSMUpeUw3C6XgXSHGW77M6Ev/KRYZbw6QtKMuWTOhm
AbbM9AvWv6kfv+4stp1dPVed+lmyuYCtAwepnPIU8x5MXKkC2VoY2zzhHmd5xlAh
7b9UonokFuqW6FSptc4DQZEaaHgfJ25OY0ZjO3CnJM85bD1j3gw3iu+wiy02eaWm
fvkyCoGr3JcTLbq6pKEpGPjIErv7nITlkeUSQh42Xd/+WvI6tLMlCKLoZ/FsF//J
QzmZFqLUxj4SztgJpLE/SccdUGV8VacbLp9/Nfg6GZgnV6lAAp6CE7sjC4dARYTa
9eNUWUAgrbhf6SVRLHn9plydOAsot62jesELDKPjfHcBYHqfoSc33/WNEapeYccI
9PasbzEP1rEJ4rnl+7SARkAQwsnd9xMDcpYqOY8SBGlfVD075lWR2gOdITaZNtZe
KZYLKiXAqSTJH+uFRsIb5fKT1cV2pGO9dWNOxWbvzYctakb1OiDoExf5yazJO7Ab
mOo19I9YkG+p7twtXKl3OoA1QK4cQDtZg8rJ7C7ZJQoX8eWWdufOBtpDcYnnFwtc
748rvXo0wrkTbJ1YWyQ01JLg86IiAuMkiFKrJ4mk5/3G6GdrgzxGc1LLgzQVJxsu
Kq5XXd4/QtpXHn0EfyGujf6sl5lReIiEQKEP3+V+aB+FRaiNoo1HvkPtCDQSeg9J
zWU3vqE23MXxPlN4AbRowVprR1HeiB7TGYS4jdtXK/4ghdC7SAiE7PhizYbbm09z
3kcdeYqe2f1GYRkJArxmXkH3LT10Gz4QD5rA6PciWyB7Wn45jGwX3WO0wOxorY8h
5FPkPKh5IlZBVpfXQCQ66u3aE5MsU/rL6+WcFuWRzwtyY5fU3rdmouTsMfNuQ+ZS
BQtRgff32C/10iejLfrTbRiJc/ybTBW1t72H4lO1G4X9xz14irGpmBszX3FedAc6
dORCcwuZ1OBUQnje3rUGDyyR114AmJRgLpeP47gkfIy4CaNziutoj3948niVITW9
tvuh8Rz8ldeCSzR+EE+Ld34d/JcskKSKYNrL4w1uROSe/BJkjsbwetCnrClk0odT
sKgGQnTijpLQOZIdrZCeWzBjxSuSR75ivS/TdM1rIIoP+SlToVOE9THhddPiAUB+
9bAxUZhEHDVZyuYwwbQLAsiFF7eZIEmScg4GCCcZmGWKRs2HHpz5p8JxuijppMZa
qYij945bDyBfNzP5chdSLXzviS6cR6uJzN+TUkxzAmkVP3ioZSF450Vr+ETrFe4P
nmXw0uF1SUFNC00L+g0WPzVIC6YO8NtFdlnJ+LxMXu6ZNpvFGt4GBMokZLKBu2T+
uchPd8qf9z134ohsTSe9RNzEuKlHJp+61V5Codvofese+xOqayIc12GzjNrQJ4jd
hzYwI/lC5zEvLIfwooBu1LEBS+lraNkQ2FJAA19hkQXW56XcpRJmNJWAG9ygWx8s
ynp3yJVXaSyd4NEFNUWgu4LvOuxfYUp6EvTmxDgY7k7rWbTseDYywuMPdzGw7x03
OlISrE19ibY7d6BzXJw12T1nnUr5YCWlfUZ40UrjV+Q2o/QthrS3/XVW2bL23Ppy
4L241fH5qN/3ZZmY1KLa8xSmD0IdmamzNCVMkGbwTSqyZd3tqdPNODEkezkcAsdL
83OVsPKcrTk2sfS1L/wOJY4spiCGJGo5fhxYJPR61P0VEUBidXjz8QFfxAAdIRVI
BE2pBHUxqG1w9rCOexR01doEPwAwf8sifwNCHaus2V7sOjrQKBwqS3AEfry191Fs
IX4YlRACXPi4Knfs84Yqub+nmmSn2iPBybstPfcGr2NYNriMolBju4wS2DXQt3QL
e/CS2pO6O457uDtG9GC1guV76qaRDnnttyzyYbXqKgjaAAnrbPvLFknHYUYC9O+1
5LKuMHFkI3Ds+FXyLJzUaFHb8Zu/XYQWVvgx7cm6lCwWQNV3hLiGCWOe4pCQ6U4Y
sma20brcWJCKdzI+1yP61SVaGnPameojgSM0Kdp8xDsFJ/+9JwHP4j39cJv8sN7j
fUIm61SI2TeOVMFnfGbq8R1lrMeYQoaiXFZLCVp8N3AQSckNAzYGErFoGakr7sHS
0P2TX1jsOXZMG6updEuOUla951siFYoyELs2I/HRm1nO7ceQMHo1DZOLv3dl5xsG
X7jXhg1uVoNf5QM9iWvqTI8gKpOoE9q6Sa/gdxqtYZp5r+7oLTubT6tX3u6QtHq6
9EJUkipUqCPggyXyS0MD6iNE5rIYMU1I2UmtMDX1OI/U3yTqqcrS7JKypxWFwM7g
JKLoa/6/7j5Fp7qmDjvcT7oWstgawcze89xDMv3wQGIybElXTstTp5E9sPxw2XTI
gK/TNOMamJNaBoQJMJGj97jrlboifWYFseRtZuE+vIWmzWJmRGcq6zfvK+ZR+FEt
rw1DdweZ8i1FfH/TyRKyaoAiiDI4IzyxkV2wjjR1ctPrhNZ8448ZxIIDtNMRb5EW
f5/6O90bQLUvsPgoH/x/DyR5JyCYUfsaaED8d1CXAytAMZXQ2bFCOrXMe+jcssbL
4sqj0OmfZTrgTIIsOQYj0UFx1AOxecWfZGVGxHCeCu1nwTfKM8ZLVoIf82lFFfB2
bAEgURAKW85q9n8Zzhl0++9DzOMc3wNxzva90TJ24GeRmjLDevU2NbzEYq/I50TS
rBqeev1+lbtolJgoJewS65xvQTXm4SWQ3KUuf6yVeeO+KIa0Q+DBxawKCob3uR0p
W51hv+GONgHpDezXRfbRzL+C9ZI7ltQoU4qp34pAFlYuTQFNs4K1elqFqU7xIBw3
FDAR+62gMbdGkJbRcB48rDEiYOG8tEQZGdBRAT/ZHGzYvwDJ4B58i+ufLZQD1oSg
4fByzijocn+Ex9k9XcurHrhzVLMwTNuIAUj2d+CrrUBUKTC4Y7tt9x2TOVcAlbRa
E2dwtwfnmJBUeAfGrcn94PAfZkYPzK2jkbdpCQuJ9qaEW6P0vagQU1AprI7L1lTT
QeZPsUXiU4e/DxWmG3JxfG1BN9FoVU3cW2VTw3GvlqJB4WhILgTT+IwPT7vyzRq3
rpowCZzcHnbLDe1IDxs639i6KGSzNGsyLXS+wUfFUdm3J6Q6y+wFwgzdFZSteBeh
HzS+CqUxUmKHxA6rNkutwaQlyYm3HVyjUat7sWs163qCwY8o73PS5HEqeeCS9xvL
N0S2a3op0QhWELThk4DBTtVZHPEzM/VzjGA8p+hZKavK/UnwncGuGjwbJwLmcanz
YYv0lmKobpLewW1apbPe2Si1r3iCeTv0K/5M0ON4fCKC/8eRWnuiHC9GbW1GZyMS
QpObkzwwA2AC5y/Wtegk+88FxcBsod3KVs3Mw+5cyvtb7q7GcNXMwJlQ+8EoVFGp
glTWaggO4g3jzVd6h3NwlOuR/Rwxyd0rQReJe3j3Ef3u+W6GbarKal4AFXs6JE/+
u/FIKkMVvHY3xVng7NqAebHvK3alLzkomIDKUwGTHmOJdvDBQ12NLebc+Va1Gs2c
gXSP1Sh0NIKKODjwIWkL1rvcFKsFfTD4/9qGOUgg4wvdINVCPg4uWBRhX648wrH7
tSHN/HsTNHSCI4AwuaWOyqBJzU8ZjbqsjaTNWj8ZKUf4r6SX40rNLnkvdSNJ1lxV
v05KSyTaBuq4dvxDecYI5nUVMqS2dt6osBXtE9BLwjNEs1vsXIvN2Z7VeuihvT6q
fEJc+qNiBLR73ERz/9d/7LTMHXCbDfe7IxRjCYp6dtB/tPYlV3hTqavN4Gg5X9UN
KXVLcCmntEvutwD5K39NcIjzDVHAYZEXbaRFNGYUFbcjnigP3VCuss4+t5V7wjXj
coGpkAG6+6czE6JHh3wYTlANJXp56gHKvBN9DFC0atzjoNIds/xT5sMAxcsMg8q1
FlB6bvjoMu6KrLpz4lZhGCHIp20ocDhnOx1tvXOa4ZpkatN61vUsEHTbZljpAxu4
BKNhcLjhZWJ1Ggv765iQLFoYZwNRjH9rCci0wLiVPAhWZe5VZhyF6p7XukIYQMee
TjKy5NHr0Wn8hS+gwhp4Lz3Daioipz1AgBcLer65Zb1rlQ+5XLex3QL1GGU0UNX9
doUeyJ/sm0rgykPBCNzkaiqHh0qt25YR6IBUSOyvNSgHEoPpWIqPcHyUNiHAR4Ip
6huzXr/7zMDhikx17e6EfC4h53KrB/wbIGtrPqDGdSsrlrDB61FTSsQ3LgMWkj5h
MN7a2nW4sFjZeaqG0GHRE6d9cXHv3eVxgTdZDk04ZfRyoOb1PI/ega5GXX16O0la
FoGaFhMo7hjBiiZzVtSmw0KJl65XNtskDvApulXz95lSSNuA5CFxqvz6QkJfptob
Lxu5vH07NJXfHNjv37a7l0FEFFIiMdLomLZi4CYrvIO6gIutT58I8kjse2Wj5ctN
JStnSDjb1DPtsuGe8+R93DOUR1B/kFC5W0S2Bf4ewCsJvtxZkreKfmzRoAqX/9Xu
TarvQDBvvBLCiZktp//PfHW19mv9QxNDZGxcffuny2jJCWcTB1A9Kbx18/+ZnwNN
ccXCodjK63v9AnjQUMx85jWt4ioC3q4wl4iXoOs3iM8J0TOsl5caEKKn4GtOa9NS
QxlwMTv+tDdVM7UC73bcEm+z01+g8PCmFDZwhpnUT6GNf2T9WA1JguyWgK6RMxHv
FJMYOHBePBXjn/2cG1tc9oM7dyy0ywdCflDYURFuCIWcQoW3HjHZ2OJIuYToitoJ
I/6CGEhq2c2Bn62af0RISKL3UtP1t3fX3gU+Na2hJPc2uk+DCbvAXewRUrbF/VM3
SKToQmDxIyep0RrfR0Zsb4NnnwqfhVcnffSsPDveqkrI8hSDHoCEWmWZulcSvOie
xc7UlU8jt2FGV3QeEfX9sBfKQeEh1q1U4FQPPSoOhct8w5q6SRalnLLNmBK9oo22
OKvq+gAM1uVMrYXKkR+W3NdDJ8FxbJ9e/wyaUsLEPs8hOn7UTgP2ASRzaUcctPTJ
ZTUd8kKFYAVjxr/Pyj7hPjIs4mFiD0iafuQCNisQpJZkvrOcLpDOBtenPpqNR8Vn
BPHPFUcTK4pgSSP1P7f5gTtYId4NQiicovTJUpd1NhxS/CBdtcThlvLD5loSOki9
AC25/Kbm7SWX9yDAyQ4FaKVsFC262GVqD3EKrVN0IEWAuH9g9UJDY2ZWIUZ9kbWf
tQ6EIj2ZCZecRzf3OV9kvYQkq4WPSBhM3boxB1vK7EsADqzIDDha/XXzhQQWd3dT
6D7Jfw/SAiIEBB9h8qh36PBtJDk4sp3qzKA4U9mjLvzfVK04gfN3hvEZpVhGo+F0
rh5CzHUMF9yERJsDCy6VaII5tqTpcxSeqrr569NeRWRJM7IPuSrmci5DI8R+qso6
MOwBqEqn8tOS1mS8YYSnkJ+HMvPcB3L7CNYpdqZMh96OenaOc4tBJOTiLFp9nvvt
CZgrOxd3K6u95xvmuW8deSJm6ulNV+ps0d45fhW0ENjfzPEAXXuw6MAWFOIYTNp0
IohJDBPMC6mWVzeo3KE+VtAHJsdtzP9KgGJAgu7xaOk7mhuxex11CEW7lGhVnQpk
8u7YCdDjkv0S4jF8jYJMpyCSSB+FWaz/qPR/4YP08zPrxa3CKlZvdqh7jPs8PTY4
KLJxDgbtaI2w3oGH4zDxFQnE2U9RUMnswsL1fwi3p9uI+yHSiyzuP1RnfK/cCGyy
OhdOy9SEq8NAClxD2T4YCuY9eVF8/qbNSnO30BpQGbuSHp4JfL8UlUVkl3A0WZAm
9p4YYaeWCZzMjwMUJl89v2gQTV6p4AONTeQRt9TEn41XmnNXRYsKZl/RAtKl9eeR
+2xlZ/DThSD9g1DRPEX0yD9XYfZOpI/GmS+90ChaSjutKEok8kzOKx7B7h1Xxwlp
pUzO7n8jJ4A3x+3Vi25ZaNut8XwXkbC6ob2TW5NE04qmuFBbCyN6rEzNTCKeAHAw
I3uID6qawvetmi1d1xruSuwKwNxTwuX0EMvCVr1hr+eUdK87wGlRTPptHZBreAU9
zEOGn27BwJz0205EfxwxyUzmP2J3NQrNsX+FaJe2zXTD3iwz37WSErNzch3sX4NL
l+Ba515dTTD6d4376bNRqpCQEsOyEaodJlpcXZJzZoFWLHUrdQEHK7ZgdtnshVte
O75rUSKApsMqvM11WMqJaavkj90PROVDCB8XwoQhVCdgk5Fc973OG9zpKzk1l/Om
xzjjpmTtQ/OGeauZ8d7IpWyN6V3+Qf9qSIwxV3uEMn60D6jPHtPlJRjWliVLupdK
7O+kZKlG0vekTl095jIgn8VH775JmCpn2Tb8FdmqC2DUQVRPY4RRYGUVMKdleEJe
3hCDvAB+d5BXCTptTPRC2Mn6szp4EC6AYcMGsD0Yxxlnx5SSifAhQ+X0zxA2/vrg
+tBpOOJn6YJxOHoWzGVjeQeJA73fu+2IhjdjDRAbgyvN1D8t3VGq8Wcx0CGWEtit
PVjM9ecnF5HXzQu/IUj7jdevLrSBtGXhLU+E5FgLfGcwI20QAcncxBPQd55wbgm2
fmUxEtxbkRJgqLHoBeDKyDn/H+KYhwd3tXntM4HxsW0q6UHzffGXxaDY/EnEa7iW
066suotW9xgC/sTyUfoUV2cgMh/5W4p6QmbngJF6RxXR1noDVL16xmIvwuXj1PA1
aGIVkdojJe/XAaoW5sir9KEoXi6C8XNzXgdFsg8w1ZJeJFWt7ly/xXQCJw3n8r00
zhyUPMv7McYbB0yjXYjbp/o0aqfcNPacmu9T1J8OhLARsiqU6x7S9YOV4Yf8sizz
bZBzq0MdFikPXEpHUtTTfuK1Cv2D3yv+gXGQj2kcaYsmB98nw72vcRP6p8ke5G1i
ug8c17uDBVr5KEolJ96P48x+bf61SAAxJqYSYmslVqk5mlwL2n4nmCa8Zp4s0PsF
AcaMR90XVztvExOmRW/UvD1UAN7cLhrOiOdmjuq4RxQAXuvhTOM+GRO5rhgx1oY2
9oE2i5HIZt9WO9MB5v0+U/ad7nvmT1/0eETPSFnAtBHeIZClRY3+6yJeXh4Dw9Nt
FvZdqGCP0spwww5rTVQu843SyjjC3QqYIURjh/g2/kLhfRBkqDjo91eA76mqoVFE
UEoJNGKzIK+vXGDijsqsUImu61447IG5rmuKf8naU75E0XRH5BZ5sJVWjMjpXG+E
cOAxIddB89IF1hIiPi7Pt2R1ZmHEbfIfXLLKzG9DIvreoszz6kzzYzWRo29MoNvW
nu6lVqy1kTvL6zBfUjwgLbtq/Yi1mxJrZoYLbbVJT+LfVktEdPvGxi1gQB3gd16A
jQmz1xw8BVPsqBe5cVxWXQ5QIMA3P8pq6XNS4bHWExnteEtjQGiLhsQgoJtMee6L
+rb1c4uDIFgOWkBMdmYT+8NLUjneSyjZr14SuBKXIiujuW42EH0WSn5Cw/dK9YRS
uVef3F7+CKlFwHB4nD2IjT2sPbDmkDEtH0/PxcSFzOF12pjMJ2EKZMSpkOr3orxy
FEevG07q4XuVDoNnCYlsrzHCOkNwJ6Hzk+hmZ8pNf+FdtJQp1D5/WymBb7/qm4n6
SMwdQXE3enZQCZGlLnPAXVca/vAF0y5zl3Tjtdgx4pjda5MYj0Bi5z/CL+T0Y9p9
kzaGrm/EKQ4klfskBL4yU/KezOFIODyzUsO2IYmcuh+SyBTgZm2cPliZJ9GtXO7n
57peXaebGFFWjHHnJx5Z46IHrwlLIDDBVc4uRShK/bOpe8cV3ydXRsBLPYRG26bL
1H3nK3+c/jlverPz52XcSadJQYTeuMx48G/TnAKvuc+bk0v30TRJm792CxFFRUWx
GJRmRdjLc0WKoF4k6fM6McVsUcccM8bqUWHBO/R/13C6kTY/8NV/6hVC8N/WVUqI
WzsOIGMuzD5nwM92sJJcpO3ZexuV+fJT/Hs6LXxLRVXNxYFPRPamd9Pz1jzJrsAj
5E5AK1ZFmjB6OUP3utmPvhCgoHIDFFO08ouZLXjEFDw6iVHeSwYTRiokovszgbzX
47CvWJIR/b03QIjCUlRIyKLc/wEp1P81c9Wll8eWIjA85qHH8uLDHylLnUgbT9h/
VbQcXNlGKRgdtjyudBif3kx+hnNZR5fwXbSuYVY9Qt09hyalnzeHUn5v2eu7d9Gl
/4UutTy+KVFtGHakX/lWqnh2K1phY6zk5GRB71UtxkcRVSDNrqXQnz2WFsoqmeC0
oK7Bu0/XjkMm99qDC/ZuZLGJF21Ij2KfVgUFnaoTFGgXDhblEEei39BAOQ1A2CrO
zThqqi5hEOSRu/bngfuQEIZ6Abf1O9WVCZpnwgYXqbRQUgjcjs+flNzcrdNdFHfd
m70vo2JCpt4UhXiACMqvTd+GRTicPmK+HNz3lyWcU01jZ+H2WeV/x8aFGnPMMVGk
et+l2pnAElLpEH+bctxPkQasst0fqI6rREbGOvZ1nO3yKZi4U4pXNrz7Dr5SeG26
8gyK5sRQFSidjLpln0i3XsBg2XvCnlazxC1u8l644RbDuYcLIOEVDyib7aH0xd96
IURgBBzL91SOVt/3FLE9uClqt/MiF/erGdXg+5+BZ0CupZP2lKv/Q/dSHSILEyzd
pPXTfP0QeTFw0Ro4DXOklcUfi8ptFYFcVSJWVfHBbqeYoy/zesumKT9mSwhHlnRF
9izp2rCpOaFGtbRIfx6oiWfN0ve5pO/09wS3idbWDSuFPoU1wE+CEkz1i7j9igXa
39Vip8U9rP1Rr4L3dMoUFa+nX96Ph3eoU6Feq2g3Sq7RnvUorhe/7cThMoVn8IB4
pef3QDm1TLRu1Ti9BByd/QegNfEs01PPLslzx4wAIsSpQxMeLpA3G1vOosXutfKu
ABz1/8SHIwBde9VmnFlwrU0qsIcALA284K7sWA3xPpiz61DnHMSZt/Bn1HRmdgRs
h80I0k9L6ObZ3j5aPhcvvsXyOkLcvY0VFVT3e6z22OD3fDlo69SELbz/Uxx8G99S
VdJcB6HfD7Bqw+t8xY0eqQI95TChSnWVEkXzkSdUxHkKwx01T2m3cufH7nxGsTBp
zlZ/6QnORNOwUPxsv06JzDTWhKv6wP/1x91grh+oEAdF+8pFpGPWhM8zV6/VC9hK
cZq6SQNl3QikOxU/avyMw5ueBoZSY1JwPktpvZLrzlPrgOUhkTzX9j/m8Jxo//ir
VLJpTQi1ZcJPxetGJNoxtwed9uCTlp5RSThFgq9QPV4Bgb2HB9wtEcZJ6CQ/5N73
WK/Pff048F0OM62cEV8SpeKNk1ACDKN3QhzKPtmh9bbCwxpKHDrtFVnh61Fs0wQ+
k/WvJzaKJGbwebYzvu/Cp5+XtagLfhKgP1cD45Sp203xwWDo11BcStazZIo1XKTl
NOkAPJMGv27BmBP/4vQ3CPA+9tCR7L4ifPuv2DmTEzLd9N+Z1IdM1f4DlmugfGDm
fLYp4WhyWSPutitt1U31stQ3DsoQMhaNo2wRcJNB6WGTq9HuEreB1MWXV8CPrcnB
9Rh2U6LYE5BZ9tcSQsgS2WNbf376YSJaMEyKFXCEQZydSeFZ3bXiKC90c0n6pPsx
Ewc5rcmEx+NNo6utdOWJUuAp9ERk2jO9d9zM1Ed6ACgez3goL+Vd8q7WybRiCqT+
v5whf1bsCL+U2OH0FZI9Ft5WoYx6GhaH9Jfh9ujgedDy9jBT7n6V8COldmPfpLwc
RmffFY8SrB5S+M6uQ6MBXT8clKJpVM6kNHfbfqXWlr9MzZqsyrr5Wh/Kr6uqd6mS
yv6HkE/+CliBb8PU/Pj08T8TNV4X/f296zCFkqUZOI7YvayIjz4Rn//9gsOp0Y5x
BhDy6+xN4hO83JY1c7jHpiWu3aOncRNf1hcuY1eNJ/aLP9iVKGS23ironKZ0CAx9
E1IeMlRKDhPDfr+YouPLwBnCU03D39TL62lasv7MxggHM8ajXARG44opQ3ycjLkZ
qhN1doXBOoQouBVJU79PPALljc/4OJ5P8TFU4ZoumEO/2yrpPaITdhjtlPLmD2zR
Iw1NCyLpWWVQwIREP7cHh6jpgza/RpEUQmYmxFSb2T/3dk0vyIea0YNDHJmrb8z/
LWio88MW/LteGKPl8xVHzX9ZuX68ajWKswBhFj3fDnR6TL0HxwI8/rWgGOI6QKx3
tSzf3RA1evs5fe7kCSeQp4cjSv5SNG49P6yHXsmGHx1UQ+8V8w9fh5+oUgklGR86
A8l9liZyMsr/e+tD8xuc3h5tDZ6rXLQQx7Xw82PwG8zd/ZWAPt4lptC7/yVOUsZp
9iUIRn2M0FrMvezKJsCitvSjhJqFsfJOIWIJ5Y+povwI9GFmaXTQQy3OaMGcMph0
/D0w8jv6HJR+Cavjimmal8pSvt8+ZocGvu/dwl60gker6oTo61CtELStbpZIO3C8
GMekd5OE+vIIf3U6uvqTAllzYh7EFCHxbDRkiE9g3HUvsLOImh3Kc6hGvgeEoinj
0boBZXl5g8jBFaVy8G5p/D2I8EP6jqlQ6aT9r5aAD3+9ejtnbLb8nb+bQdHoYlRu
1WH2tB1ptdHJYdTJbKIirN6kExgOfQDwWpQmXTEjRURee2xKIoWUtxti0ymdjl0g
kKyLC5loZ1WU0gtjNmkqtAcqmeS26o8cRCI0h1X0/X5wASt7fMf1XGtV8kx9jvgD
kqA5wDJLumWWgN2AQu2UY2Z2V6hrOZb7dEOcJf64vdYiOOpcD71t774qjb5pwwXX
KRjeAskk9g34GYSoeKzkDEnOzspSSs1a/Zeq2sCH577fY0tugZvI53O2jbtORhzX
6ZcUzsnsi8aeG5WvEXr4uz5pwWcNod8id5NTqWX/U9H/RLW6n+fs5Ln77JTncgJv
qacpQaiLwXx5F2gGdg08ca8wTEIE2XLomroh3WQB5A9oLbUcApppNRNOJ58gR/6R
ZHbtzhp5x0bMujt9AVSj/FPe/nPdx4dZL+SO00WKuGXrVxQUTndwID53Gs8voqeT
oLT/TgDaOh72EXXEjIzXfYIsWIkSAQQnx9zM0Q3iJEVA/xbmqGQrQEozufOeJJcs
u+l8zQNVXbbqbIZzzGUedaHkwA2IyVAN0LJTZTzpk/T3y4xv11+4flJbntVDRyFx
UUepc6nONuxApZs/pCWWJ5op/vZ4PDVPrfISkXs8Yn30kg5JJeEvAtR00abWpNfm
9UOMPQWwvegZ5Dinlc0WFHDQel/Ny+Xl1474jEInogQoGCImm+RrVNGrhWrVIk6t
3jhRUzObD/0ubGhNWJ4wyl15NWwsGJstSxzw/TcPkqIOYU5ljMKOBVzVANfA/gZ2
KR5S9eDNxIsHIQXMYgLFAmwZE0mpcmAurnoyFOO5GBje/x0R22N/cOVPaqtEboG2
uyhZnMjzQk56L4aKxCsIQWv3oe9JXlGRuJhjrGtglhUpoSePAfs2sK6G/rUa6xgL
5X3xzNHYKMsgcqpoGKdbtq4zbmhiZO1x/q2LiFuZ328PYmx0Qg5qYS4rDhtP/xCv
aPU/oUlrQPI3GXFesm5lzUoEGzKYxzGs67e7pafxJIwATGpifZRgVUvpj2Dod1lZ
SQjCtUA5qDopXpfZXCFGkLPkD0T7TNMDkfjt4BLbTMAEi5V57qP4ZpI1Cs1D+pWq
3gbf61OGJEO4K/r2pI91tQ/5ZAZV1IXBqxxBzLJUO1VbHIaw2W0vqM1bAVN/3fYh
+sv50ON10HsBsttNmelR/8l4mmi77k9XjkvuzoYCo1r7lu1taFUROuqfHV8fBxv2
wa0zkf6qp6lzy4aJj4AY3TTkKArujx3XpehBHjxSJy/F+r0WnCsqx45LkmtzDMe6
wJ+nOvXZwuqjKcKQj4S+D8FORYXksHEkGeGWvUafsBU8IBPL5rn1gf2XcED9FRzZ
rsS6PGUgnVOmoTn2GTmJ5pUBjnVDKN2lWfRC4OARyb7CPUbHFwmkP24e5w0qPejr
7PDWNKeP3K9O45CNj3OvRvSZTMfhwoN6UMuz/mU80kuZ+7zVsp8R6a5c7YzK3nXN
0gZZpejwvvQ88qctAzON3rIbCsNgvfDSfx2VF3Uxmc6jKNrW5/jS0suHlO6tgaEy
djI403cKjlkhpirSmYXGJDhX6tw3kDxTuvqMuDxT10MReoQyvRCjXKyj4Frd/ADb
P3rwKS6RoXlFnJbfwi16dz+NPSM9DG9z948WQVRnZbXnDxsUHS89StenRfNXBf8a
/jXhSNdN/PJ7J8PHFcN+KJC7ao0lvnQwu3V1Ed956HpD9TnB50puJtkUz9qPiaQD
HV62Cv5FSRRc1hAdDp1iowaDJ3kR+Nkk53+axEUDMRLInq7dYXK1OGbU39HbciZP
cV34KXZtQbdgR18mp1TLKzQ2kpeUZUy3bAJv3E+48ZZk7Ud051K7S6RcUP2VSvMI
Q6pDfUD+3fUVuyYoFYpueXWEvr1Ze5/Cx0O0BTp7z70t22gfm9flAHSb+ekqiyFu
gWUGVbCjInPeZS+5w44oL2LF4LcChHEi7aZyC9AJVni4GP/ZMWRm2F57DcahpRya
Fdy/vBuexqK8EHMsxNAwKAIMCPQ+3MmsE7deObQP4kYPvSMOrI4cehpZKjD5QaOT
/oyyRzjZhZth+hWOOIiyYhkj+NII0qKnOYPZSaCjR7GjPeGH68jGnE++cwPpfSlr
LIdBpr/CRxcGHUK2M3uzoQr50DWBd96IcXkkW22fVaBMwJllj1ObR2CIdBn7IsN1
BnEXaN9ywHSXix+/IpZsU0OJ3Jr/Tq8GaKZ0HxfO7uJ3uBupD958354nv15QMczt
a2QkscMYLzoPyeQz4o/meSMObRAzHBraT9ypYlfBAxuPvGK3oStdRBwKjnWlarln
NZtN/+Qq4RiX2/muTXe8dr+i3Whzl9QFWg6/OCryrg3ap4wyj3CVjxKk+7Lcg80p
bNdE6YS5Tpp+/+9RFZ0nnQJesU9OM4gTnzUqk6itKhS6ob6W5a3RE4VLE/TwAwkp
TCtRkwFyznFerPR7Gou2Ps89IuKFKB+Uype7/EFh1U+WBx3LikWTzk0E5rlMGcgB
37Uoez+sh735ALT94NXTBfOH6c6goJTNCun14wWSmDUHlcPtvTTclPqjoALYfq2v
9hNrsI1b2pG8ohRUivOGG24L5W2Ca6jzg8lH8T1Hd67DzJmNGLxkhuHwgtol64BJ
DKfUy+WNDtZj+5AQYn6O27iSPEPPqNrs2rhS3iTndI8izv5LMJW3D0Tmh2PjdznY
VGPFs48aNzjGiSnHU9xoAydFNAf4oOuHPCyXxDfKnmvkv23jmSC7KF09rO0D+o1I
EjonLi/afs1l6+efj5jRcyzyzCEuvfP9jpVlZPmXuJ8Cxp6x21FCDk+dtCzaOdIv
pJcYVJCOYQLa2qSA63EPXKNcC/1ImAKvw1yD0FgKtfpBpgKz0ZrBMiDkuTLNasjE
8fUyeQf4YqsqoqJM35tpSYjaQMKRu5dkkq7hg++uj6h+Sdd+ZlThS3hSMNW2fB2Q
Doeh+IpMRuuckfNngkyyOPnTfXzsy7gdupu+Rr/E8560EU4ve589d7IZcIgGaA1I
cJhpXSq1Cd76RBO2/4UQwbFzkuJXTE59lC6EA8IlLguJG19V8V7snb+s5+/lkNNu
zFHTbKn6j708gknNUt8sK/9LId9HBKyBhN0bbIr8tR7atdz9KclTyPVQZ5+dq0um
ljCh2y+sf+HgYiH3QYRXrEWNztoew5wvuSQ6yRbxRlIJNhh450EGvL+TBhp/+N3Z
XKowhk2Yo1iby0WYYsEr3IfzlPzyeDHI7tEmbDhQZZg577Eex5BDhRNKa4OJ9Re1
KII0BqO7fZJNJwCRZ0UPCiIOY4yv4GD/EcEth78b0piaQ9PgRK8ex0MWPNo4PBz2
EFSCop0SVvP7yF7QvGDj6jE7LlRhMQiW7W+s9KD231HIaVD3Hm7pIYxCDopOgCfi
TdQ6r76qrcin84r6my+nXUSXGFECSi5bjwvpuaiS8zztHbpdzLapTVYbLGdr/yJj
WuAO+AqYoiWhgRqMXIhH66DZCjXbtdbrsu6YmBRbPWq+TClLeh6EUUAIxMDbisU+
7Wqe5irPxxysLT7pywioNQKhxxlh2gIWZgdb3kWJjjOqBA+6qL7IFH31ltvpmYZJ
VT6geOMGz0QZR3Btib38zbSOdGWzy+p3CMp29OSDZwy/Tt3IAq2g4XjJkikP5H17
Tlb1aGa/ihVXO24PzwrIEL8QXqd+OirJqSmqwL1wnIJcHRB2hCfkJ4yZc3v9w/ZH
PJQvrpWIwp4xvO0ZdQH+dewDzYQZl8ZYiA0tYx4ctslHPIM4gT/mf+if2sZP5zyn
TV8XXsgDisYQk8/oPhDcekAWI34Vhaa71q5v81VKleZ4oz0yTAcxgCl+t8nLyMtX
u3op+BkFeOXVfAPz8WhFzL+1YCxHoL9DpvZ4w8jqqqwrVWEX/LETlZd6TPClU6Xn
bHfc38TspoX9iVTjts//uHfumDoA2mLQeyGIVKPD6wBzzR8WrRWT1YE4OkWLxqEL
VOLZ2biGSHecXQNjun3Qa8sbafxkd9+Kr/QcsJA1061j/RR7CJE2uXVFZQMvwgf1
WeQp8ozBDmr6bZesdpXyNjsHizyiWDz+X5vvigMU00nLiGnJsBQYMz4so3A9DZWd
ZyS2KXTaEPK5oAppwEpw9XdLPZxKvPbaM1WGNqpykgFb3UB9RWhdrdYgm2G03M+R
3STrZCg7bgjcNL7u4BqKLL/Ds/s74ztMZunK5+Rl2CDLsZX+Wc/s8ujkmtN2PATq
dKVKWEtr+JP+MCNR/C3Ns1XXSNiyJrZcsQ2xhFuXXtmQUepzSuCOuy1Cui0lVjxV
vv3extGgP6C40Hu/jOpu3ADLe2M/0VUVr/I0kKPndFS7nF3pqkX3aoAoMQ09lK9l
Zzp9akpZYx/ERc0KrJFW+fX5wriXPnjHsKPA10NyA0rSTXQwjejpkeCOw+1xbhG7
HI/cbbk80YrfPPf/AK9Q49Dc68C2TfXHUSddeocMhLHioP+4AvtLm6/57Ea/yiZK
2TMj+n3dWSf0xWPEUmqQkMYfJb/1+CvwcHe5KnLPhlqZCuFdnDHh/fXrMPWODrh/
4lxdzsvPfbMcExtvzQw/RGZ1YXtkcaAmTcnwC0BZC76VWiFe9xjkjbASTDBrJaTE
bUPCEULdFmOqocLuKl6VLDjDdndd3VsxuTa0KMeZ9to/VnFYQT/6i8YAzQHYxQ8M
H5YaWJus+ojIyznK9oEriy5477usGA874ZXQsBJcC9gZkZXv1YXqXYzdmYwqFpI+
ByMhjpdiGS4mQqvVP3dom3xFD7LY/NWzIRJ7f/i6pt4ON7G8GOPPDrD8ZV6GgBjf
NZEAKNUVMzEV5ulDJSq2+hrl2i1TzVMLP7aGcUe5w4HQMt/JcSmjRDo1rXc1g0xM
mLl5ugFRW0JHOTaCwyetERNRKfR5OAt16uRo1GhlPYiqbtxwKk0bZ6N3ZiyGZZiz
WzJGMuSliUnDNQC7G/4WHSrQT0MaB5pvLe7/cC7J7a7i1mTGphS/9nl/esJq6kxi
iUBJO3er/fArfJEF1iJKalJhSQUxWkMm5Hg4+cRJ+9irv4mgBm0WyiOX1KaAKwCk
stsz+j+x+kor6jWZly/Fe05efwaeOXKQBDJEzvsYvGx5ODEKOQOZUzxP5O4AH2Nf
nrqtuY+W3hmrV/Sr2nA49E5K/cj/kZ8ZDRGQIDr4h1Cy4sAnZfAxc+qEWWEbNaoV
Q2uQJ/Vx3ZoojIcJErfEmxhHkAakny385hc0P9UYUQEJzRdZFi4p33trCyAxiGKz
BR4cI0vsoXCwVHJeC1luH6zs/oqAdvaGlanFYAmsi8rjwA9KMeir0ASSuZhmXgAS
lAvrJlobEldpzxGzk43T8hfhZecHFaRD4OiS4hCVksKKEmZZNZ9G+aVrOp5DlMih
qu2dZfOZiYgoq5rIolPGb7BKJ/aicwO/aDh7LcobM4NLEls3M9COP1kJwNj7s1ME
53BBv0IfbIvSA0PxeSTcfi5PnArQz1+jIPxV3WiMkeQUnoEBMyvlWAbHsr2gWxNd
UQJYyi6eIe43yEgCgoCHrzP3kS7BuNdp17tZP5TebMMKZcEJ1jYlasMtsSFzaSgU
cqACy7u5/mVDNhrLcAaMkbZOBYXDnS1N/xKR6kGS4EFdr6WzkiqIJK92yQJLkm8y
3xT8qNPjp/37VvGVUZE8CckdQ/Cy5kTuxHKvGvlQbU053n6ZygXZjbaDuaG9J8CD
VPL+xa/5ku3edN0mHuM9zPZU8tuaUdJrikwanXliZeULo1R0yT5xURrxXO8jiwoT
u7SEPPfF1oXdLy/ZK01dd+NI4TMDlkzJL1UVjntfTHg02xAvTeoBRB1jK81Gi/19
LQVAmKQfyk2+NjNhvF3+6NIhMfu4Mx344LpqcbCxLUA9hOMsAa91+MCjKnzUXP/t
qzTocF5v3TUaXjrTStSlfyGSO2/DBKwGoaA/Nwl1fX7AzC860YEgpkjNrixB8SPz
TPLsEjpx7vU7GysQFRM52VZETOBpoh1ka9cEeDen7t/d6ZBvzA0Vuph2qharjZGR
QjqMhopZOLqMHzk4JKy/+dNj140flvcf/SkxiYnuA6669PpDs/WcRrPgBhkWRqsr
ibCBEQ22D+CFUnpd3PgYnuNwRIzlTqsLiGranxutYuxxXjRTZOatmObzM/zhulY4
ifSUL0AJemTOSV6Z8Es4VIj7bjTGCCEEBEes1wVZRc5jLT+UgMztucjq3k2kALvF
UVVbxauJ7jLILNB6ZAiSgi4O6D45O1CK773GlxmkHxqmenzyNN0TrJZxsrbMBr7y
fedm+27FpaaufX/gyDBhJJtNv4dRwk7o1ZD4Ymm7/rj5OYmxRym+uwANJZjmS0M4
+8KR+c/yjY9H2IgOsu5Y64yr4fsQoEkDmMCyDbUW/EY7UChwLGV8qvBJeOGMAWca
zmEzDKB5W6dAYYxHW1Xiom2Nd9GrFl/sHUPTWZ96oQFCOe8KS9sCI6W9nIws6A4E
3H/cwua2rX0jR0VDUGyrfB6Wtz01ly2AHBd21FQ/Ua37F+Iz5F/+hwarJ2TtIaGD
uuYdN7vwuxYRD54lGWJzWBMUuN+O9qT+uJd/UgsKqgpV+la7H9kZiUAhECxLpbLi
Ft8nJCZKl5vm1eBllji2uLJImL7q4SITa8gejRBC3NMZNzGn9DQqrpgSeYP70a7s
yJxv7rBHyPcWVTJiEJBxMvrJZfNYo0ZiAx8tgJUI8WQ39eSSJWYMa89pechgIqTo
blx8t6gNjRlY2cmunmcBrW1vS7I341ZuvBkPWa4iSwXxxULHMy3gbXiE5hMplapR
fP+VdA2BuSY69Jth00LSPkO3cUywd0mmMk59GyRqSuBeJpII1frRug0cJaQfNZV5
vGyRz66QeMUi4WMp2PUFuNg0rC93vRFvguvQBNxIlgETNL17sWJIvdzXIcEjqfkH
14xTKF/4qZcsvbsgqLzv/4l1VMHre2A2kVofVdaRaYjrIFvLOecMpM9GiT2Y7R37
1tDYpwZamTvxhMJ6wlKuOLHV6I9g1KuRsIWW3UQ40BiSA1Ww9lAG8Fcmo/K4JAOE
wKdLgBAEXbZl51bbTmtY4G3RPt0gxu3zVBn/aAE1gIQJzLFxz/a6EtmmEVf08MR5
DSFya8V4x46/86YmaWWMecaT2G7eMKnwyoWCL2KfchqKWf44ygliruJoXOkD83qU
f2ASfuvbKunFyiczt2+6dzsiWHRY9Km7YahMcPkjxfN4q3E1ClN5q0xWkiEcG54Z
SLhWtnw1Oo43NYSRqDbPaJC9IlDPxw8Xvkt0pGD4lhdrM1gLqNIdDuoE1KxGu19q
ATw86xv/kWB2QE2IQT++lVAgfAf5OgSKTnyRW2+mAdTBdO0XTGR7ZpLcCD/dha0v
PcKvgimFpkm2WDxfUVvgtg6GlCeVPijphqzOGfLWoisXGFjrzn6yCaYC7Wf4CWhu
SCulBuGgRcytZBrgU6N7TIjsBymjH+mOIFEHyCaluVoxrVrVLgJN/xgnqmug3QaZ
Jel4TF/i4rSLRzyrdZZYXmwW9U+niTAi+NVH6HBfZOyIfhiRs9ddNZarTp6tQgth
oLoRBAcb/K80b1i8c2FJZNigrOdkA87ga+u1rB34STnEcxVStGDa9Azx5gZL32CD
BE2e+Hr+XllPaiRwKzXnhJ5H/O049gFkK86A89YeTK1FFCx1ABoL8N+Gaic6GArs
tHsb4iyEmgl/1vkl0yIuXR9+q3hNy3Ng9yH/Rs6zer07TNRrzR/9cCd5Sf1xLQPY
7fihbKv30kHUF1T6O/KYb9qPefnMnnLMEhSB5YB4ADnP+AjgWrKjqlSRX9vpYVDC
A3MoU5DyX41eGSX4aPs5kSWGCauvO1mFNe0N4Af0VuFr+1t/W2+ficcR+YtIO0ok
gSvl8OcSlwDpVGgilTBSWJ1yWZ+DWEQrth8daZhVINTN8PjcsKCOeUpjxz0R644Z
e3n8OUTI2cFo1HWteLMw6gxNSQHMDSemtNYe7kbPPDO7ioA1U6upQSWK9tzxPFxD
/7qhrTzdEI1qu4okK9z/mXVTTNMEO7YjhQbja+ncVB9eGvvClgIPvEU3hZb4POLA
ZbcCC9q79ftilwBl/n2C2WkWx+7pEAaAQVqwJDpPQDbiAo7LuI5Cl78ZvRtcVVoQ
p463K1Vv+QW4zC+nLLiLoQiqbe+nEdycJpPk//v8eXGYZVsn1mUCf8Am1Wr+CSNN
iis8bXFRpMffD70Sa2q8fNiForYZ0ikgqnmevfNGmu3dJJQVsN6oYq4d0fAS1t8g
GRtxXQBZ/byoBfvE+mzxVZsznpB2bhnUl0dvNyPj3w8MgtqqdzY1bY2rgUzxw+Hx
uOpHmoGvPkYOq0hWSTc8rk1D3S3YkkxUCjxpzCtARHx8YnnN81UCfAFC4mOUSa/D
KaZrk0DgToJHegnUNXaosPuwHzQeLWEca+3dfDplBdRA5lb4X7tWxKFwFL/S4TRP
cLge3kFeHURxljJr9MZvp++QFP1wc3Avkh/deCftcMbjmRXahiRE3hyHqVK/Sx4f
eN01XRMrYvXWtCTDf4lUP574qor4JJ9MCAx/vypsujYMuiXvLwsEt2JwXku2xLoU
jUkL5IUFMYAf4oGukrH32vJGZIXv5lTGUaBONhP9hLNRvEEk21r02Ud61OySRMtd
roBDfyM6ygb/yek+WBsX5u7OvmFfalQK+tX+poUEGWGGrjlW5PF3414VXK5WS4JI
Kz0MqOESBVk+vlGXSE9kJ/XjMS1ZaPoMCJQK3M2U3K/QEPw9Jk0rMV0t4TB1wXNN
kR+1URo9vtDggfiiF4Ys6S3hI0nLKywPBGz6TzqXL+STHxg0l/VUPBoI4Pe5tLjf
bL6wTTgijzl16jC+cDNgEZPdgjC7hch3ENpZSJxKAmYLvj34Qoq/SwLQnn8dFB3F
ubsmIOiCyc11IvWMiehlzMdCrQBj0PNuM70m2E8hK0U8fZfCY7KGDqNf5z+g+ha5
w4JCvUiKrtb4Tjxi1vLGnVUm2WtTx6t2omWV8vrA2CEZiHqSHz5ZdZmgcTnnjxNb
lSNx3tZzUkRgjMLpvHAzTm/kkthLDyepjbXn7vWbNHs1Q85cVBZsDO576BAppz8l
ASUsbKSRxDXLmqM0Xb7jxuMUwGMJFlKmQai5p6HR00xKzKE69OtIqExNpDwXzVI6
QD3p1sXhGXaJ9ceHCJBBQR+3hhA4ujKCvQYFq0beHvrVSMjqDRcaUhMQM3NzrapU
a/I3mweomGW8Fy0ezZrX/Mk+UEbhg3o3qAmArwjhBVivLYXz+gU7l/bV+RFgjV3t
mbeevZWrv+9InFVJfpTwS0BnoO4p5ssYbdVj1H/gJX7Koc0Fp+4Jq6kcrFxMuGiY
Y3Op3H6/njFs2GxG88z8zVWoGmy8uQg9O81fKtsn4m1lN7Zuy+Uigk2hp2RgYH2+
KS3z2fq7NPjcLfzs040ZUpN5cL4QrnO8WLne3pOLUDvk9iKN+D9ZHkdswS0uowzh
ETERt+N7LDqDY2ig7w2DJSdRAy7PNzdSU/dKY/8z3MDjePCdrqoBlJT75L6k341x
qnnToTV0/QLQlWZcXW8bZKJtyIEphswMv+RZ9Eoyt6lOlQYMkF6ViaKIj5LOr6nk
XHIJFiI3cjDJsKkSVI5TPirVLC4M3rPgMf+rCyhsWBsUQHfEJWJEVTIOTZhbbGxw
sWSmgj52tZgCFmiVUKRhXZZPJeDDvYgsaIRn4CJ4+XUXYftSdzwqjPyt9ZIHj1wj
a7mrfjc6unUnPJIhVkLefX9W7YL92+BrDbJfszEx1A/kzUsHosKsr02PLXzKdfrk
vTPxkUjTBSHvFyeaEFQ9CEHgkdmlAkZFd1XNN4ZyXYEBYdEZRA5OcKpbB2jNRdDh
PRHdggZFny/Ejyyzufhqf3epVivv93BfAs2fQBbdtnFjQjPvUElhKrkZdDSlvKrE
q93rwMDKP0hN7sKXp+1n5KIh0kl7EWk9ADMRjCpd0k6nrFDWe99slP0fdrOYGFCn
1INkERUjwRNHSAxi1g8+OdpRwmSbMlHJzFIBANnbrGjfGSbrkDGKIUyOQWEu02km
wzEN5HJi/QO9Fp9KV1Fodc5vhmAo4ezYazKMCRuEL2vwifaYrD2LXTXluTbpaCit
770DkrpEhWgoFyW7yxtWaFlcezfl41rS176BtSxUseufX5AoC/VyJ52tabKlQ1g4
J2BIDQyJt4ebntV0+3VIJOqTmO1kmFM5yplv5GPA7wa96o6E5g2y/uTsZyOtbYhH
+5QCcS8P4oBMM1VU3xnWeNNNVkgLiasPfsbKny6Fqq5c+M/mdBHa/mHfsWQkSiOM
uGHst+Bt4ihHrC96frTAtrYy/9efUNr0IngQaKiCNRv/Y/bxaqslfCRbP09gZnn0
+yUJv9QWg1k4a4FchGiJupHZIrMVgnK6zFoxYsKdPGlvtv85qkH43lnotO7ca5os
4J9u4EmYiaWmi0padg8qhz9rjHaY9qi9JrN6CqKvZ4G+5AR6rNv4RVP+WfT81bqN
SkKC3HpLL40dXsE1PyAKSezgeZ8uJOtmxVLek7YtiIaPlgpqgiQsmAz0gvzHfZZ3
j2TfzlOUwkT8FUb3ieAPAMvzOGV5kXLrStz+Ja3tbdZyIQYoflZcub7icreJDpFN
+WDK+GcJZ1YbTtRkO9C7C6dlhskgVldiw/ookHOFaF2tb8Grf3M0LGCabTclXbBp
zrMaPU91O1OLLf0BNKyMRi2yUqnwgPm/F2d8SOx/glD5rnCsx6FR8TrZtST0SkeE
CfcUpdSgdLC6X+6ldLjQ6uymtO2jPO4a+cacRjeqCAqRs+XurpC8J0eFFs6gIa0p
kBcons7UtHa08vreUHjWiWap+8+ECTSIcTyJnAPqDBPJy2eA2qK5Msf5gyxOrEvC
5QxnS68/7Dmxccyc6fIh8zDbIvZwGAP1xOs1/fPtz9sBXOhTD1o7Sz9QDSE6nrGx
OnRJm9qS1iElsJO8QlemvaLUDDK4mPqf+EOV/FLmnYt9/cBjGC3l0b+fuQQaGgyV
zvhIp0Mf0xhLH1gmbhHIslVQ/51fZ9v+RhdT3CS9ltatLIillQ0pziT+a+LOWX6B
ABjqBZXlA/EF9VVgqDB1SY4R4p1H7FvGlXHRPLZQAeF4q8SfXYBIemJ8wEhQa/qm
4UCmCgTlQftG9zlMaYxpH6Zmw0CTTrjKjxKC3OzguM4XXdENTXxeFBs6uaUbEjJk
I5eUOv2706smPMF+AqQeBAEWxk3vkUIlfDGg1PmWTIByRfYdZGYPzRTHeb9nzp8N
kfL2UwPNlAfgDXrP3E79u3GE588z4m0hW+2/GTfEZu+jv+e7o7Q2F1NvqnKcMAcT
nYdgP2Txlgj8FetAmv+JGKQegQlsduNQKIFpd34KwdyMxrRvEHgepSuLEn5CdZeA
NfoI3F0NdOTSRTA9k6X86PggnLxu6OEhAaYAtCn8MqQfiRmYXTvTi/tmPmRCPL9i
LTx/WVqkANND7f812z9klU/1fPFtr1i3F5O37/76aGBjIkKm7UvpiMX1xhTc5dsR
COQZqSxNlLj9VHu0f3EvEvU94dR3bjzCp1Kd6AdLS/7ntQRFD4Z1ic9PAJR7WuOf
u3sgqyZAaXIH6FGxFwd7leKM5CA62zz60AoXsO1FrFI10G0XjFrShFGDvXYrZRdk
j1ZvsbPRNKSI+T8uJFOtjoSrpTzWKajpEHHnHYs1s3mBOXiFDSMCBQzeqdbqPsyd
BtWVhj/+dShzgUi7P2QRFhSKepHxBMZy2htuc0tBsdKe2/SA3//jHtimATZvcTZq
L003TOKvYOQB4aYcuiFAR4dN6rx4ydcopOzWH2OJ5W9ZOuOcYo0AcdMxYOAIQS6u
eq7qVwWTUD0iUnQ1WqV5jHES/iygYM/moxNMn7s3y96RD69jioVnfaVa7sYIh1w6
ZpniuvqslG0BWbk8BBqqYsJnd4FnMELd6nBInHqGPznILrZxgM6iWh9b1HK5q/Ae
NiX8qUIK0aMoNn1AMTF02ZUvasCUpLDQJLCdsodTi/0tPjti9aX5RajJ9mpn3jE5
ACE2cHKxvQP4ijubwZfRqujI9gBC8X2C+DSoUSX+c47XVqpviSZcF9am3QJ8iCx8
4S/bbDQCnIbMuCDcV/eHQZniEJMmT+UpoF2vW4LxS4iUrKEhfpymeO0BFx6shXxj
6EGVqNJSgdsE942wRdVgIF34Fe0c4X5Iyj/d2y3sKEGuLANBMoeY0mfeJm249FIK
Oz5DrXZLanQ6spodBceBMsAXIQw5q9OJsk5z9qNhzDiF6VmRE84dzP/Dg9gm6Gt4
Gsvf3Yy4pwbD2f9pdeGPchy+Zl0RL2Y/wlehIGsh61xJtPPm8Mx+/TKJo2v24QQR
qfZkMGIBdHU+b3pDDAwruPqDZfNWr7ogC5vTAHv4iUoaAzCtSdtlYM/JPPKH14I6
DLnXZP3TvCoxQIx0Ljm0Eg5NqItHt7d5yr/4MPhCMbpuM9emyM//yaaow4DOjSM4
oWK3ZUacSYNT3OCRbDC1AC2KEyzdLXutFZx6PpzykDzmWKUW17tJp52w5Ll/LzJ1
kbxqyR47vGA48Boenmy54ap5vVmlc/H0nWL3Z+yo1lQD7SsZlC++Gtd3lgVfwn8d
n7qHf8IcHZ44xgf1peSIKO88rMPrWqUAYo/hhhIMxtcluuQ3NlAqSCAIgEZatWpG
0b8tkGZF2koR4cICAqHAQr16hlICz8XcTRctE+LPyRd4NRJWvxaeaJrHOjJ3Y9gD
v9Pc3NWlCSDNlX2iOBP56UVZGee8CAQ/ySOvEk3w/cWRkwOOr7blCW309403Cc4u
sdcwnLzucVRulYfXana4jeZhEHVZNuLRPHaBkG7eVycXeFzl32iH+PpuS+Ksw3qE
7dwoGDBiW6Kq5rJPjujNk3rTj1vmAweI4gpbahfqFdiTBTQIwBFWgQRUPJvYLGxb
Tc/WHuIemt0i4b7dbfRHJHtps0VZ7c9fmsuKqOY7xu/K+dX8vfxDSd+zoxoH5pPH
zZ3NeQmFhrqGOYziW9hUimoNmsdUbk9VXcAueZD0fbBjtyzqiOgONmFy9ClP8+an
pEMT/NlxP8ppGZJJpZCclybPyxlPd9+63f8va33feLrSCxRqNR04lvvqLgIWPsfn
2q6IgC8DQhG+53LfWJqbjUPzxbUxwW/Msyn5WJr1jsftY6ajetoGGwKygO70jvGD
/INHKKqcIs01dqlApDu44QH/aNpgRQ2WZuVeW27+3Z0rB12+qs7tPisCPXl3mJer
1P7zb48vLQ1Rz4RrGgO8Vu9lxHkPl4tMsog6e7G5kJJ5bW+rVzcELrC2/hQRB3tD
ldWwQQwHxz5INGUuQLor60P8Q93b0S5rwQ5DZESkGWgcOsHnL3oCnbPE3+LbU0xs
7pNJt4pDItgi/n7lii6F6dyOwzGlWATGp39idvrXkWJvVxB3mJuZ5rmyOJNzRTXv
23bgS01h8JGxrspiKFEbnU+d1sRKQPZcBkFMj8z3sMNHFdno4pSAAmPh9Ud06/KF
VuWNO/6GUgSFFIoQEPlNC2mhbfbYTFiLqJCtk74DzpDe8KlM0oiIdigYFG6jxIqt
85ep2qaOQyL7SZbeZ4CqKOZ4Jio5lbSxXNl/Sl19qPnSXaoeHNCQz2vY37NcGKfJ
s4uKht2C2VnBwHdpDmoDxMamidawWhDAd9J4aiVjwbld7Vg25N0N2A/RDuc4PuKS
cSG/KQBIlYjc984xvOCR6pRx3iMPzIi4+caPIqoHBR6zzAct370E0abdvGVvd8Pv
9UNwrnRuzHfc2YF9hT03gMh0KEwhUq3/LH4eh/M6RTrX+0qQphZJxr3WHe3kSHzI
cLEvTenZuZwfjUYj77JY+BnILEEJrSD7lT/sEFdFpCDbexuSyvjsLcgxYYBsGKfn
QyVC7IKnvc5c1L7QOM7kE93KFiSrS2axDA41XNOYy5Tcy0f5RGW2Qn3bwDQVMw5E
mPu3sH2T+qCag7+e5qvPscApvSOI4FFsN88XA8MIUYHBDYo7O19xkvsk7imNo9Um
oMcDIc/yLrvkYabcy06poJIC2aRwUuTatyXF8QsZCIEagNxJrXIZUA642KeTpUnc
24RLGkaV2SWZg5gm/Q5n5bKFjH5bbNLOtamswNmBeCO6kpJXB2xLXjXU0/IrAiKr
jWknFyUr4r6lzcuRMd6HMX1pglHaZ7X4uF4aUlddPs2Bkp5n7glerMXN9M0meBBJ
gEwhoq/wA5DR5iuSet4dDR9Vu5JjOwVuNI/zTQucc11JHFKhnsYDpSKcbIhj7ePF
lX5NG0Wh6gNKHALqTRK6c5tnkPtyVe/Lr7n6cvA5fg9/p8HNQtZkr5UikE2Avc9b
o1j8XeeUjcWGV9visMGSt3HU7SDdLdSJRbCNDECstTh7fc4NlN2Uxm70MVq7x9/I
0NaMDlsLCNXWPknGQAMqjyg/VDBPTduBDS5cfV7Lsbe3UDYaCNZrZhusN/bb8Pos
pGubblUIBnoQlav5OdGMvDKiZimrKljQumz+0wIOE4w8rp/OeT3Q2lRscTBLcd7f
NvG+nA+9JOBo5QySH4JMtYplNX6dxi5i83kcO0JVts2riA6tjmOY2tECj1d5S4Ek
Z+MPD9tO/tIpB/q2dbzoF4Ai5ljfyVPZpPe6q24tUFqmfv7cEubF2T50cdPOJ/Go
OisjCFy1Qrn13MKGudgRrpEhqkJm0gVTsn5a4WeMGAbD1wBS/StB1kzv3YWZDNZJ
f1bjHDtciCoxSc/vZ08Ep7djqcoCFwgbs4jbr0EwL2ahJwOay73ODu8YL2XkL2BP
wwt9kyku9WHBpc1zTYIjd8/1HBmABquVcPG2UVIZG4Q3buRO7dK9Pl+O4u5LlS15
82hQS+BTiaHY5wc7Vgo7D9Kye638GI/bPV914u9ROVNWFWUZDIqtjxyLVyT3GEjG
kLTBeDXT47SZYFDSpaGqrWIoTx9jPGes9OHB5lfj1GZxOO02LKO2Rr7Uhs1qGRMj
7vGioEbLhiWdKc8RXkvghZpK0K5A6fqO60fwVxw+iVMgJNOIssvV0PhlgyAzQuxi
i4TFyiLc9130ClBtyqNPXQOWI8YhJttu0HddXe2fzYUY0A5SiEnjkXcbo04pmvQo
10/flDyY84vqJjB2OBuIDmAv6f7WUahW1VlRQ5T0E2przUL6LOwvizFU1CjKfHKK
pLwVjVPC5/ffVEqD98IwkkDQgl9JC/4XsHfz5fCjxt+P7ugkyWo3sJwVWYj6qEhu
su6Pc+Ji/VQMy8cpgVmaCIG8ZpqTqV+UUseeaH9YcsngHbQTqUZ7EDk4Bkvn+r+A
84YpbGMgJziKHqiX14ZM0q8IOmpqfgyJfSInS2LvoWE7ft/7kmtS2qPls8hn/R2e
tO6te/NTt8XIzjQ4GWRpu5ZRPqonFE2Qo03gBKbzDp3+AcOpe6YezAZKUJHLaICS
uggJPVcX+NhTTqUyPmhnFJjrvEMP+8Y5hAmqwekSJSEAZRqdFptJSzHk38uy22XM
Udpnj6BMXmkMNcfKN+6/BgXNDsfgSefhtit+ZhF+WKuIMy7ZK8FpQKAdBsEh8cY7
zTh/Ol2/lKejJgrrBxN7XS9jPcRUF3IZ0g6HU/6ZOb0QDI6k2ssniO/IyofUcc9b
h3/SLLJDj6xkAQ7cNVbME9Wk2no6ZHrxXlfED6aaGJNGZOjLxYQOboVRFTa7R7+W
XF+Kx6JoCmB9Mk/NiY7mwtIdItMFpXGYBu3l9D3m+uj20ncO77MBjAi9Ig9eRzvd
x42dlRzhKmnYydddYVTm2UxkALseVbnhqiE2EUmKGvuOfS03aFOuLNGgQgLSpsf4
hYq7lrI6e8DcGfwMNGbG/eIvVmncW+WaLSUcoLsNHaZj+X/D5dCQ+XJPRNRthbBb
HHLuDhWyOVI4yE7wrQ21jRrFgozvgm+Bc6CtquyzMMuFQLKvNoDeM5OQgpR3/I6W
yFfpDhjyJUeXmdWGJOn9Wz+Blt/4XHve7/R/K/iCMKEZjPb1Iqef5Zi/KF+boEWG
JASmY+chizJVzpm+twZa59rQRUAVfBj9nepYw7dFwRWtxVJ1CELw8uOy/kzOK90S
PeWZdgkH8pFd9A7J7IpcV+z4HAE4mXKNX8bNA7hHUR/t00nNZ/CSK3u7XZZtTHcn
JOJUaZM2pmwPtT7OCJnmWzfqtMzHwjiJHtcTjGOlWjLAJy5LgVlTr9BhejhCxolo
KlXpqma/i7MwpgFuHAzhSyXLGoY4Xf0nNOtILE69dbW3RydyewMKI0XauBVXkcnx
H8ehe8HMLri3uZxJPTVllNVJwjAZ9ioOkFm1ZndlbtgPHYHhh6uscGED8rsJ1Xxk
FHyheYHSGq2rusfJVO5dihFTvV71UFMppWPbUadZ+L4x4YQdnYhqcdeQxCWKiDPZ
YRHGQDJMLPwTYILZhAjuAiB/YJJI2hr6IqlGvIAn4cVNedbKJMfacfN0yDBqgKpJ
t6oKqB+L6iXMFKNQSaCTILeduAS3cbwLRe6RRHFcHfAkU+fP0B5GyF3luGcVfi8I
KFGeZ/Z52Xc1vuLTORi1IjVH21esRxNBzNls46it0Bc24J+4376B4/rJEUL8zyIf
rHmfpXog7+cV1nU3+eiCqrR2XTBvLJEaPlpB2gzkGfLUXvnCTP9oHi/7sF8p0lPF
F2cNff7IzYKvss3jJGhF5V2Y/zEwU9uDbwxqC3TZ84Zbg1p2TQmCJT6P2oZHR8+5
Om4chwu9TnwtUwDFj3+tAtENB403xNMpFFRSHNU6vJ+c74FIzi/FNUtqCwbCfOJ5
hfh/IDgDrh+xWAHFNnMJaJKE0KzniwW8FHhj5svNHh2/Rzg6PhzOwCOxqv4Jaa3b
wAqJuLIprYj/Oe7c1PkCYRiAZQg/oUoxyTuA2Ai+Fx7FGowjHtQWuQtzwb0UjczT
ZG/+kn0NVt5ydDD1aIKG2JK8VDBl4cvYcYQAFQ0KwoFwK8I89hQaeTsiK/9CD2xW
WhlMyyg4ZxoxKK0WHtktr98A3RewYiuspvnwgB86AsPTjozvPtIgNphiIWRmgGVg
39MnwAd5ghyqVIuZ8I1pwi5V68PLdNogxTjxAfF5dOtrfT2dMAH1+V20EPafP7rj
+N5PjIW9Cjt/rqK+D8w10nCpxl6wvTpITMVE6lY1+pPDkceFxCMhPp+aXJCU1OK3
FT5942efHCfM9gEZbVI2aqKt2l+LiWqhRA3Ak27OVCItPgGJTArecQMIFA5PAF5u
QvlpX6ETyldR4teLS3CHZKPJ0FY5K8WPIyYip5f11q16bKXkK4rI7YvudnanNmQT
rU215dOs/xILUmQ4v2SscrA6dS0Gc4S4XgEOBFDq7ytlbrbcu3x95RjyZK66b79n
7waR4FVnx1gfeA3Z6u1Tm11SlVHgkxYFN3IdoKPZRySWPnmjMVzWwkhua2DiEEOI
eQD5SbTtqgApih/F0sIKR5GAxMDPmglv+R1OCh7Bpp2dMoxA5XO7Sw5+3L59gpl6
eqvDV8YV6dAH0pLlvpQYKfDVoqLcMlr0bx9L8AbWlFWa+Jmrwwy7PZ3YqzgW6eMB
rFV22Wfb2si9BImpJeDx3TTuKisjXiUe6W1vz9PygjSZ7Lyj6aG8o+Mp0azPHFnC
DsSKbwjBHYPgGsOt0hovneEQsMA+2Mu09LjeShgh21N2UXmN73061vYtK3wPr+UW
4YZDvjeyDU0Q3OyLxH/ZoRZ/fpbx6l8SGvjeon/MlRdVzawdxp7gJslwm6ZBpkeZ
c6NUFD+3y9JNrSx1TaylLwVs1mLAjByL5crv7s3MArEPdct1HjirAQSfJBhqNB5Q
XFF0uf9/ld9C7Rx8xs23saj/vqeqPXL4n7YIqvqQ+ydJklUBPhgzN+4DjKIPnmCD
Z1Qt1w7Nhv3qpnWZ9ledUnRcQvMDbhRbbk3YlV60bwEr0IJ4r4+ATTMzwRNHd6kN
M8tHg+QjlN8DJpKZdXu9UWz55r6Ze17M64v6eS0kiZI9EFwVDnQqwjjddYC9843+
zu9QJZXSHxqSIuRX5JRKVRlTL9QHzpfHz6mLytki6M3h4ZXmE38tJgRcLv1r8YJn
x1fsdLXUVhTMlGzVvNsCaq/imuaCGGkUd36bg5p54EFwBzKDaLtlmZajaCVldymb
n5u5Ks8yRd7xfT7rh/XkDW7Ixy4a/sqTWxDv3P/KVrGNR3hcdmfudbzo+2hqJPcC
qG7M7hRkGQzuxTw6Arol+o0UwmkXfY3nksKhNeVNqadh52I0n484xWB2uGqkZhs+
Ed6zwvmSEAnEVuV3IsLYHjAX5eRq84NbemduQ2ZO8vvTT3W0lYHH+v+Bvm/9gqfR
b6RlsLpPLY3sU1X/psP36LJC5gZg5H/IU8X033ce+IPeB9lzCl+7DAnsJzxfHKkL
TPBfSN8WN6tDLHBZx9ghvcERxLqJx2x4bjPVJnlcLQ1H/0Nrq+7K5OA1FYOHSvyw
aEJbXK+waRxDjeuwLiJJR7DTA5M9QjaFmWO/4fpV8iS1QmXLmF9XecY6llqRngzL
4uHeHDvvVGFLEkYNmFly6RUhDE4ZMWUIjd0Rm8Sfzek2P716nA1iKeqp2d6Qav5J
JeX7iavgeZ9UUd9IBUOkZ1q5pwOtBAo+c/X89vuW3S/2YDDlyBbnH5oXxQho8kf7
jWBb5OZv1FNE8tFxMUgD/oc4SV9P6KZ6z2Xvlme9o/KpXpivhWWiNwv9Y48iKT1E
lF5zQ67XYgdaEpuAOeKkKU7BiReqSMTIlNuARECErJBccUNHGox6zxQ5Z8p8IU2G
M1fKpAmTORlQwH2ih7bIkqtdZk2EDxjIe1//xOw/AejVA41RiPGex7DUOXDJDIiv
raep8Q5Uc0gF2liaXWnEchue6REClS2Wk5MkjmtoExkUHYCOq1pCo5l/y40X4gFN
szcoCI/DhVyQEqtbYO2FmKYqjPYXxflDdBRIkZfek0q28MViJHDByVa2WW+31Gx9
qzPkyvmwYosyO04GCb8K5vJcEaadKed5gml5zKooG08uVkCsy+qCsTwsxmeZpqnv
F4geGNXuqdjRg96SUFNfYQO1aHMW2V5moH3DFJFXYBHwUseBMumff+Ku/yGYvTuM
CksMuuRN2biYVra3sWnINd2llOeSLsPPl61znfugoobQv3kGo1bSOUGPTTR+jLjN
FTcbI4yav17Ep4759+CaqL2M7+heNMdX3Qq7Ib3IW6QdpDNhrZ1OQ4uqFGrpJP4a
pA8+H6Ml/hCWm8QFVb52hUvnp/mSj7G8dfSqtPAjcwzkVwzca9d8SktnPJfrPw6U
5j3BA0hg3dEMjEkM7/7oxfYpRJOBGfwLS/Cnl48jRYzk6Vye2axJF1oql/oyen/h
/RcMkRPR0w3pSJnAE9E5rLpbxi1Evz2IGAXa7+dGILJNxgILs/0ard+4KSTbuabg
wX43h4d0T1y2WJ8r5gROE9mbkeG3hEwO9QkxEj96LpWqgBDlAvtLqLv1rMEkFJCj
fxySB37hbPcikRrwTOJGdQcowhxLZCW4vazBu1QTKy7kGBNxnXTBbQeCkqpetnFs
zPCVNPY8VwmlprMnu2c0YO0bhw1E0Bzym+ecWBnJYG5xv0UbEBAIgRZ38Ac26mHa
Fihp7EX4T8dH7G2uPBVuJfSpH6lsWyd1AeT0ONGUxkO2L6Nf81OnJG0H5JcilO/7
GGRihYlNPlezQSCZSNju+VWfdV3pWyx+gpnCEbwbuCaKjfY9p5UO0P6cNP2LWH7Q
I4oa1gmfcgTtMCPxaeqw12N3nyu/rj8vKGf0t4LWdqyE6UiIgFcVTZjf+Zy5bATb
me+s0X25O2eqYnlxkHYFA5if+1cZGf7YzMCv8XsY23DMCVZyFnYKL5rMtifv+Eps
j57hsaXearsYfnljyGjN5V/W+NZIws+8onknoKJVN1jpxUGbcyl3KTq1qIJYVsnp
phd41mraw/IeQi7Jhqy49SFBHVPdkkrs7eY4SKCH3XesG5k0SbtWAl3gSsfrpdgw
7PYGEmk4GD1PdeZDK1BejRfCvBx6xx16siA32a+I2mIGSE9+8FSS0bKdPagAMJPy
dkz/Rp953iT0mu6Jjdol3XVpvEr6i8YiMtDtMIGbBEl3dNMfVFgeU26pwhEPKCy2
3yy6JPjvOvXziYiy113MS9b+6hvRoI7DFsybDF7Iip7Z+AtFRvt74FMwD9yQidA6
CuFqqVgDMnsOd7FZ8eKL1dzA8Em06T52u/R2u60baB7Fmg9dSIgvx5fLVZPK2Ydz
4v09x7KkpnD0KReOImy+F4hRIoZr1vs8OcJLLm3jW3uVSm0tXbIc2cn0bzpd/zKQ
zlRIJOwy6OSf7GXtM5+41amMINGecCeNRSRlJQBldCv4OM90vCzSTlz1ovUQ+6uq
lWPaV4GGfRmSYvjtOND+NhaMKzP1XVrN99/sKhm2/tHEvAgSlDautyuYBQa303Jq
plPNPM8oBfYlOv/m17JxnESlIYqeM9VEtBTgN1X+GLZSTv/l94x4Vzy+croZeEFR
fKdr5yYpBU/YqSYZP+BcdcuikW4caF0lXh9aBabN0W5Z2+nFRACRJ7XeN3qdHz2v
kNr5nVNW4zbpufmDkbyd61u+9LChWG0CLr9+mMcASIaEYKo8M1Ob8Lfynx4zN+Xa
S0gse4dt3ryZvk9jNCa+ECb4QwVDHOA7ySrSbuD0pCjMclUIiufbinaezb0oQtik
ErItwqDvOgFDNwmsBZF1SxXU/TcSFkrabMBjy5UT8+PodHaGIiEQxphkk2SxltBN
CvOgy3q8Qc1+HikouLRI9QdbqpLqjIsRNfBiyWv/2ZsaO5YaT2PGnmRKnQQDjqej
vumWGCU0pYRJxErICqFdBz+iENbSRYwA1+aAUvaSjwJtbPtmKJiBpwFUpiFMXHi8
kLyH7i+EkTvrMtACAFN1IZYho05bRhv9udQ0DaNEPxwulRFZtlGW6DVKhNCG79uk
GKODP23I3beHdSyfb8t/C/50uewPOq/oJ6MDWvE7HwssTiFj6aoNpV9ydcCBnq1O
qJQ3WNT1qmjkTVOmSxAdavGMYuq15IEZzcCbRaKOGs1rtlaQPPXUJN5+yHgRdqco
DyuQjJvHqlzIw0jdTOOima1WsqcS/gycbi140Ec8HawATCQJQWBcS9AqfnwMqKYw
t3lOZiqv63+OMzzKtVkqsJ7ju2KZCOHfhOT6Jg4ccYKqFGpWkm52hsCKoQ8Fq3a5
lDI0w3NqoGBDXOS+00NoBSyusq9SyAIMuHJwuBdWYu0RvIj9FJfnx1KyjTh08enR
aT005mv2+Hsle5MQCcG5ZTglnVEi4zryLVMDzQyFIceGGcOl/VRTJZqfB4wgJTWJ
jCeIa9YObf/J6gPpbUAbWAkAB8EIBbGeyYU8w7mAgDQOwSftW2s4GYRMjvICCMcT
wMvgR5T+m3XXgD/EZVpUtc4GcO+UpF1qgwV2G1n3PJCYBzbn+4TIkR1dkV6hJMdV
JRO0dJ1mWWma2Z8v5GVC4ag8u+hObfEK5cmEjsbEjWbw1ElB/4ExrnVaZj6elUDZ
cF96236f9OE/NEs/5OwGP9pspe1Bv6S7WhRPvUUi/uBxRrzq72Y2dTNo++z6xZEb
YEzHO0LS+/K1un4CGEsFM8pmFEttFiZtbb7bSA+E4kzTzr2NQ8veph/OhxMF085B
O/crHYxk1niV0KQKqAehgeYEdqqBrAJW2xUVkMOcO1ZPJ8Qm+CozJMXoCQx5opWD
mfEfAQ2Xqkjbt3qGoNPLT5pHkh6quSxYq0Q9ctao7gXPOgRLLFSPja7JmkyoK7ZI
JG8w/AD1Qp5UI1aZ/gkvYioW/oiiyv1iayEqujLJnOqjv+XOxe2JbfmDJgfRLK67
Q1nhoqjNSl/7tDMz7KP2hN94BqSbbmH+OHN/x3hZaWzCP6U54BxUoI4onsREe4le
L1DDymMFtQqWf/QiCB376lTvsRwPq83o+VwJligh0oJ8uu3wjU1EFsCqfW/MVxmz
Iuo1OYW9v+TLtz702VBwiuqxA3DZ5rqgDtwqKHBLrppf9+UdwKdRqvQppqfrGRug
5THBk8fQinWeenROBtuMITGwQQjZY7uaAks6o6b1wwGNhZ/SuWxohSU0uHvB7mXO
0x/P8YgU4kIhWBrHmXuc1n6CIatjera/p08/QTY6LP2saeMjrzrNfwVll+fTCeWv
uJwNYIz3DEy9PyTR36EqJlX+KZ5VWVusHDdSGdGAQKarOSq4k4d4MHZLqJZPZg4e
kz+rP3XXtcP/S7QvuuAszpOtj6Ip/0O8entN1ZZddIcMTa/ADb60Q7tjQRBA5e6/
KfQmmJ4CKAr2WC+xvRoBpmEyuWVtFQKPBj2G5f+CGFRA7H7+IdHwPm1O9qgOaFrZ
4mLmfiiXXqEg/OQGNdF6U7GIDR/aZVIdkzmM88jTvE3o/oEfQnxoXWU95AwovHRR
wKfjUaSwvrkN9Rlv58cKjHS8QB7CQGn8EFh1pC5ZWOh2z3IM2SjFJSMTtO88AUEb
m4Q+BZYSY/5WIfA8tFxP4MBhItqX9dPhdnethpBoTFa/iM/ndHPk5k0OqTDvFYiW
6Khl/P2EMAoB8hynSb2suMFxYe6JY8TyoI1kEBZ9McRl+ZnUau02u7QdvhY3/E6D
L9L+dnwk7/8EB46XuuqTzqp/4hlEhNrLAVfQsyoBLg9ZPeqB8dx64wWK1pnISsS0
OtgCWpQ/RFdbk1p83j1fEW3CxB8uofQ39BL6PstW73UjY0ucUxJ3Ltl+GlaYFRdk
oHIxe/dTDqyXirgBtXZusYiea84UwUUfMN/hh37Xft9rWz4uvsUte+V3Svj0jpSC
VmWevKMZct4Q+y8+g2FlRnA3bpKGzFuZ+1Xtcvxt4tQtg4yrj5YttRSfwiGiH3qe
AnoQemiAKUxC2Xx0pwbGv8ypyxjvAUS/0a96HjnuHj5T8Lekjy3X9d0TpMcJcnVK
YElxDLBhEpsYBM6fCQXKvYbKhCDxRkIfYck7MOL/W7HYgycMMInHn/ZnW4DmcL7E
Dg7kL1ThwF2QHSit53mvZ6AWvXyHwY18pD3TK/z70bS7Ls7JCNfX3bIKxB2LNkLP
3XVfplLbUAHh7+D7l6Ct5JdW5T+4UefjsPvytTM3cvrRR7C8790KVHBTyU/06+uq
QXpFjJSu3dUzUNyKwzpvLtmvECiTErc09RXa6R3ggIABtJ8r8KYKW4lu0M+Hcy+h
/KU/JtxwGi8bp42/XiUV5M8hOXHU+OFxFiGmGjWZ2M1cUmdFJg8g0yPq2EqJxdvz
5L+jU3Qim6bTuov+HFuKdqiDEciVX7H9NH5NjDaZMgO1id0ZQAAKP9xE30d4nDWz
gw/uV+gTInUO1VAtaxamd1/kGtGkCULvgDt45kzgyQqN4C/oFLGl3unOPJUo9vwv
E0kmVu8hrsudcnk01W+i9cO1cXE6a/OMh/uLqQfyPtY65jZKVJkKPDX9AXCf8oWV
4vvVEfh0vQ5kIw5hg8XKyWIqSo2ndQ+gd2nRHm0itTTpZPnpSZ/xcPVj63uCBq2M
32PnFSV/YsEAyKbJKAuZR6/556kn7kVrsrQ60G+4Ycn9lxRUPKTjaYWVSRhkh91z
uJELpGQFTgpqGDjWpk2wKYqE2cdF/VUampIqZczD2jWD+uAODutmKDT8KTQx9KXm
/wKe+Dp5OiST30fKQF6/Q8fRfzsnyEE0CyxxlWEGFT929uFnMCY43c+PBXz8Li6d
1TCy8cJM48AC1xLrjxcwzlRhBtrZboNJcpT1ho8A+PdHtX7CD35QQdnJ/8rx3MfI
ywnV8RAk2CrH1bfax/RoKylzI59MxzvA1MKR3pkQxNG10Xf2VZdafhAUcuayKTru
FYvri3Tg3Z8yaxD2HzfWQpc/Xz3+BBlm9aEYnyd2OY928c9trUeXNriqtepjl+DM
f+/qfyudumkUhef+u6CNv6PT+fJuP1ADqng4MFtMx8QTL6TWFnJgLTtDsCs49S2K
Vm9Ios5OoibkhIyctekAvNqP75FSnZMAGZT45o8LNzrWT2OdMXn8QPwu5Dt6TVv9
OTuDFck3+ib3g3ziglT2j/EoahjIiQdX3r5aNtluB8q1JbyX4VdW9utWiBk/B6pP
OUGXDKIm397rAfL+0zVsSXFjL/UbuYwwG77HGVpJho/s0Zlreik2GVUym+ph2kFR
UiTFOcTamYhRGpQa2WJaSHijmW8yF4ua7IcWa8y7Lrit4ltP4fh4vHx6U3LWtke5
/89JUiNip3ekkOE8EB018SmaD8jU4+uiQSncsLrRrC5VWsOkxmfXyq2zC1gduIfl
7xZGoXjhcVaWzfA7J0GNmzFNI6UpgF/zbK8P9lr38JBtZYHjK/PB/U7KcKW6UGkt
UGaQtFFhMuoDJylzxmv0KcnDaHLYoS7FwvQuogG/IJahLOfvbbxOmL4zaSqGR4vc
05UnwlXIqKGICKM4P4WnvNZC4LfibdSZN9y1HOv5/+sHGB0JlmgD8RQQAclkjZyp
IUB3fm+fKs8+a2JZWmRRXhGTj9dnDYP8F2jLvYRuQtPG287GuqOey/rBX60yjpnu
D9SpCjY+WsTSiJfNkHVWvgjaP7Lx3afF/AMSlyP8tPADkRTgG+X1kOsndFZzwBnX
2WzsAYARBd5kAAoS4H+x1Ck48c+IdsAYlIx6gIVTSn3M4kc8495BCyxfnZlJvCSh
ovV0Kj6eaJrt+6Mpgx+EcjPk8rAjmQRZhBCCRnl9RJmT/18ir6FcaSwjv+uVk4a1
Q61s7sEC1OFjGyBvjLddLHHJyP0i9N28FLYHwbDg69FCIMy+CpMBugGfrdCgs00A
bwSVgVbECOYHCs4oKYSq/EPDMoK/UmrXuiL39MbLLL727QazHMYoceUPNjCs3oht
mk+Xgw2b/S55grNZUYZuBzhfVlUa9LxXH62WLyRjg6QJpPHWszCWZGDxHogwXnKK
tl+nJPz3Oo0GmPoW+ZrYwerXJZztsDhPQ27ERuS5MOfEdVpP1L8FwXoTUfNRhWUk
YzBsurVpv7dXSNbQWmF70K8lL4bbGlb5G8JxLYPThSLaI3zTqFDwCEJfsEmKKZfE
DvLWBe489fo97oiEeSkWZxl1sVhU2g+vh4bVfNl4Kf61nxPAqmAeIkr9zYyed8Yj
uzABZJGMwBfVHRcT8Nq33KMmJwzHGMPWOaZP10bKQGhWpFnCfJBP7rfAlXgC2Ast
f7NkKupghKQ+8OzCFdDTTUCgMbDKYfxQrrnDjfuCOfBSzhcN32qbxpW3blaTuyAc
bQMVUuhui+NqKYOdp+VzyA1+NVbqx2zNmVCE0dDi05uErM4omc9o0v8u59HTSICt
g07Xd5DJ8GjpgNh3CL/jYcJfi1knCbCCqMJx94WGV8h5YSVifiCaDwMefdX2olWm
1mmswX7I9ENamn79IRrSeaxcr+JrHFw/8Sdxp2nSCKAkBNtlZilGVwg8u4wfQUz2
ZWU2BHQjzihwzTGhFcfM7/DleDn0mBO5DjU8POiaabnE4sm3hjlw4vm2mEn70Tt4
ZbnZ0OAa2LfleB5GQc6QcJ5HoUHfmv941HYYjj0F+uPgYJfzbddgJykao4mDPckN
65otarABG0jWdvO+1sY3TRWwhdGE/y5Sf52m+6kLuVt5dvpuYQJ4SH+JEkedGmu4
zC/I2kJyD9bKOXlxiq8eKv2g4CdZjfmhWbuBxH0G5ERw/D2WYlfevehN8Sfs+DlY
USXwrpO1yxpQuMWdxat075yzuQJhV4wN4UyKrSWR1vwdaMdzABWCOpCyCRf9Bc1J
C2rivPEG93ndR8brCG4Y2BkPgnqS6uZUWiCJOMBVWr10oHwDwwekn/hWzSMdLgv0
SkqiqsmIad1AcyRZqygCVYkFx4/7feWMlonHdz90+/0Z6TjcY9wZvODHIiAoF23y
OjqWB5fEBaUgY0qf+5za4Vqf6Jq9XkKt+TeC36eQFwNtbw3Qnne1yaFVNzDU1ipT
MRGgS2wWfnO6192f9HFaMo21ziQNWZkqUSBZqS8ofY148Vyh9T+K6uAwk6ncKT2J
PnEcmEtELj838wLGCNxJCLFkCilDvUmCgVdBm1k8Okp7L2TXDAhFp/iXEfka54nz
lL7/qkewRBbaPavpiqxDwuTMpPYIBtgdtAX//I3zgsMHBf4kFvIc7A8ArxxOZLSZ
wccUKCeeInBWcR3/uLsapFnTjuM6A8Oig0u8z8zP2V7MqLZF5b1reMhkcqjvx3R0
dgG1sVCUrifjGERsK+KVLxFLqxuSB2/RiwcNj8q/DQHXbR5U01hviAYpRqGzb9m3
lsjNMJAC+CClLDXsbGJGcEenaVDM/Iv5x5f4pfKpMpQVRJRzzuYXnxYGO6xESY1G
QKqruuWOHv+4l2ZsmALW6Uw2X4JYneQKWjz7fCTKO/QNr+ES9W1TaXavoyAfkXDO
ncBa8w0G3wJ8a/esv1aQm6xYDc7KFeEnoJCKNPXb+Hv/JeV6Po23Ji6G66Pvejki
Rx1doNklsrEZ96SRmq6f5bjKiLLxU1HhA48eIsY4FUiDjByKyqnPNn5UtjBz2S2q
fNHUcKwIbYqWh9DIDjLX2n+weyu3aGEacwQLxOCFKrAg+RfLKjV2n4rgI5zqVEOG
ibAWAs0UMKCI9h5RUcCPuH3WwBMV4upxsIIp252l7SoXLQe9XvYIVKLfzfvhlKvw
JG8wIWLm8s4gYL3tS8sXtezhU5Jbad9ALr4K7+5l9RA26vIDWAtZOuDsCnTwq50b
o4oO06TEZcuUkepqhAJwT3RnXf5EEncrS135wm6ZCmZRb7Rm0vn8ruNz+H96PAaw
5WuyV4ABPgdV5fJ0Vax1ziwCbsr1dHqbAqGUk7saRlWRLwclOxOngG4NvVu5Y3Hw
XVaXEwNmwZiGLMSdm8ReEX8S8Wzl4ZsTFUN030UNCG1EN0HTAwG3eN50ODOSb9E6
E4ndUWob2DRAllNk10BsKy/mkknMhmGax8oMtRE4bCcDha+ZmztTkjYAM0Icab61
bzDWlahbFpHJogW3Gn1A2bHLheAd5uCq0W0PQ9h+e/RGGnqzdn9laVKBYB5QHNir
kjyoADgYF4DZT21Z7NaYv551q12O6wJ2QKV1QBhyozrW5QIOVkfTJAK6kfahdrKh
C35QT2dxLdDTr7p27YDqaZGJAP+7XUT+UjRga5NXpBB+ZOpu8sRZmT7zZglt41BY
WXjZbFMJQL7NrtGenuGpSoc3Uinc6vTfDij5EjTLccGtEK11EJuTWXSK9QrdhwTk
OGshc17+wrch8F9hCz3ceiSw20fIunVf+NLZZg0XNKu7BneUumLlYoFXahgoFqqP
FIwPtcl/yp2jeDa4xyVnN4UKiu6vzR9swm63/OOcdOwv7LZKC+GARpf2x3A7fcCA
tjDWPN2RGYV4+CZSLP2US5I3nicEtD//X41zdJ2bR0jusu+JYBmGtdg4JhO64SOS
QOb+5ymhewGGhvF+mkTziJJtUzV/0aoIvbKY/MEHcQr8TeTr2mTkrF+2ZKxhTy2g
1eb81bTffW3Cc0VkwYstKZoGcm9KvUqXYI8S0bbgOafahVtcqrqUCxpCjBodr6lz
/7QJxX/rLgmIMJSSxySW5wJgDHer2Vny4lZDLo1tZjcF9Em01Wb03XQjJAHKwqUy
fSFr3yzWMnKeL3HFqPAyEX49F35pw7gXiw7EdQzoFYYJ3trhhLwv9+AQqc9P5j5a
hiv9n/4M77FX/J+qj89VX2rv8dMin9rQdhWXzDZWY1vDY+NtE7UQnVKfI81TjYXL
AATZ6kIoYwSVrb3LlGtuq6a3qCsgWkiX8DwEXA2BQQTzu+2NMAzuvmDwzKoJv1ai
7nGww0oxtlkrZDk5yoieKICNpw3xusdd9iG+Xk/5PPfw+VK2HUbdOt7j/5TVOMxq
uYxcC5Cqbx6T0IWai6DtZwe2S1NXdHHbej8qnqSOab5AdANuQit6kezzDBv/P3uY
hxqSEIFiPgDT39UNOUxw4n3+aCNR8WUtmf2C63t9DXL+T+sB7V0HzHf5SLhaRadp
ShZmm3TOYXMNb4dScqQjpn8g2GZnh7UNcbJrjBoNu681V7spYB7+/kEekl9KCmg5
fLh6Ep6Jrj2pS/ASUsBAz6DwXEGCe8NLGxwsKC+YgavkMWhFflLA9fkdalqiqyR0
DpZjC5Q8VQDxW6DXovr8B8h2iQTgVBP0Fu0fzkn0BLWJzvSK85fbufPLJDfb6UdQ
wbEDTWnp4d/PyNroB1Y4tGEsDYoDaha0vWzFHEdvrTK/Rf7GwyoNOIkkl/ZXWVaF
sI15dOWRk15aPsI6Yi9XV/o+H1Gkc6PdoEOcOnA38CsE/FhfC1IGcLbq61OXHjKI
bTPxbX5M6c7LXUZ5c2wmif0KwOpouURhbXhIISPX6kbC4JCH3OE8dP5TPiFbiO8P
sReC8YMWF1IsgOuVeDC5hFCpbWpYiyc3a1fNb62ySG46ncLa/CAZeLhZuYzwa3aH
ejzahhO1f7BSZmS2mjFERaX501WcWC+69Cl4+06+nmY91kXwUPqhRzs6PFGEZSDx
q15bCmauCbrHuvoZbtZY8MdQtyKXcdD/KMYYxDqkIuuvIuaL38N0M5yksPAHi/OV
qg3MNt/z8v8i0kkgkF8AmhP3eJwhsBwTngxfovMC7pWFMccYDq05zSEV5XcYmsZ7
GcVSX1IzJZDCh5WRVqgG6ESYtsthohuaZBNj+fKGKuSDk8+EDCeSb9ijEfE/ei/n
I7mNngkJt2xXM+3/xNgReJ5Wmi3xXAaa6yJAoAyCGWT3YP6bwFFeMGwGH5/7SLK0
FDbMYxbdHshx9snVQzt+Nv7SSchpbJ/k2rR/OjyM+pYVvkKHs9F6A4+J9U+iZmPb
AupUgYdxMpMbdM7s52+0NJIln2B44QCA4GGyZwUYZwB21Mlve8WCFV3ukz2d7B7r
xwuDL02FciE+jyrz16a+3R+cYwAv61bEFmAor5GvOwiCivO0E9/3ZKLIcjzw3uOL
ARu+pNqREzG4Gza81ADPteobiRu5bA0Tyskv62vv9PN6+M6/sXqbTK56DFd7VG3/
H80jwc17BIMoJkUqf/TERg38O3mCDw+/guqMVdBt/xPGQxBlQ8JFUS2LfwK7yW5u
iDA3ylyhCWGEeyZmsR+43xbki1gu9G2L8TU2KkxcbS+oPX/9zwiPXKsQFh3SjRgM
7UuTIi+7TVm7WUkbsQcIo44aLzFUl5x+1l5kgyODj9v17ejQbSPBlaRpfw51p7Cp
67uGInBYtEE9jL+lme6lGwXdWfCqFdTBTb3La1/6gurVjZEY8whqNxP9B8zPyfJd
2AU6SLWWDb3TR8w7GE545stdaYatia4UZ6sxzKWWFpwLUR8W1QrhwvEGkDqbnl6f
Bzqd1pPRUPovWf73ss844P2mN4+pXNUUzZjHx0XSMGW+9YQGqNbrwgzuhRB5dyEm
l4DkKn8PcKHcVJVALqXH/D0ajQspm5RghJLygthmMKU7AYLF85NA2LsROcrcmrUf
/ZExE9f/yPPtNuhV9WsPAiXH2aG3AY3b2cZlMgfZf8A1oG2LpmHMbK2DNvOtB8pO
5T3GR280iLLbJtDeNvEKAzgn79ahfYet3vafwum/vh/4UDPGo/1V5vF2Xt8qAp+H
NBc+lqNEKwjpEME3Ghlr/NY2kC9LxR5IgS0m+7vS8C5BAONixm1el2XX8Tq0N0qG
tbIvWUcBBWOH4cHjfbWaZCUh7rM2qwYu4OdmfSMzSXk/uc/YIZ5cH6HrkQW6vuKX
hjNcegzPbLUwERX+3cdC+kBo8r3aJeAsmFsg+tV4G/PNERetz9WyF32tjfQI94kn
No4i0KmmCafxBStt2yhylxO4nAvBX6IHTGRg8khb3RQpyNeOF7mYm/nPICfEJYIm
V7Ta29QGHlqFc8BoA9GG8PHHkW3ycX3IVWnhIjvfcz/HEWhZfCgekxnle3tte4zL
q5WIYN86Iglbz5nDmf79LL9DH9Q9PHlNxHd9yL98gXmvUTYzdCJzw5E+lCcGsbcp
P4zwAMWDGIohUfomACXhnJO7kU35GZe1TWsSD6JBmm17F6CAhc9zWoP62KeNPsgD
utJHmCHiYAPrB/B0HyMW7XXeg258iSsRXdfcUq4NHWCEJUSP6MB5Ym0qLfBMlG7L
+yJrvnI6lXb9jgNzaai61gdoe3DbBuJGR0V8nFpsepxgF4LnP41HJXMJe3A3ozpk
ReOfzppwIDYUcYVgbwzHl6yYHiEb/OiQ5nrIvRYS6/modzZqMbeWe7EQMDsA1+f3
3eHxQdJWQCfF9/+EypOaN6w0ZCszpebTpsiGW5CMqs79H3tz6tQ9VgAmPNQlgARJ
IAqmiKaBX58sgO1b4Z2ZGvYt7LXzzHT/IjY9VbrZvUzrXLCv3fwKqqyKVGrkY/2X
htWxr8YSFMLdyx3nOgEy29gwXIs2P5gNexlcfirlDMEsUADojRmA7Z0A3di5LBtb
QEwjyvJXrR84WQKZBprV8uKGJc6qyM8m2qzKyoa1uuNMbnDC2IM1+alzOinLtwQ8
RZYRChFRUvX+EIg1Wp5MbDxPsAQcK518bjgXelkjhd+p64pVsp5yeG8o6K6O2rHu
XAnbJe+G926L3ekBCIlrP82XRSZ2qxEKG6kd1nGKJs3uy+Ax0iPo55PmnGf/63+X
BDWUmZa0u7raJt8c/Xwov5dSz29pliEZH7w6jeupCYoX4SePdPwXf4IGfd8iezKy
gF/SD4EERs/zR4TQI+ILqzCrUnJ6r6+4LmjJ5AyIi8Qf3rljsLB4BDm1TeHUl3gL
7EmKRFidXPBc6PP3M+vtKimIINIOI1l1Ai2lJEOtnQcn8YuAHbQg/N1c6RwXfB6x
EcI0LG2+xjlI5C4rE5GLSMj181OONN7JV49rndkPmS4LHmNA6psomW25wqgmGPJ1
NCiIidWlpzvnVtrnu/PXjyRPW8sc8UsG8GyCk97vKiMHsR19X13ZJSp/SL7NwtSO
XHxCJ4mV+IJvz9J+HJIpduw7g158doafqiKxI2rsskZEey6c8M2C5+HdV8q2xfP7
2HmJEcVqvGG7hYWfwo98RcZmMsVWyFPviB0ZY8bG1wKFUrnca4DI78dhanM7kLy6
9WraySRPh0ME3D7HY4O6824PvB4LWp0NchjMXwtaNySQrvM0qrqZFGGlLEBEPDNt
v1rbcvMISaAWT1zGvNl/rp27j/7I/8ZdIkBrF2QLcd0XhXsczhTcdLhUk3Xf2Zoe
c9Kf0wZ9gBoCUHsv6KHvKWiUtdNn+BNJ2joFavjj/p0kHkZ4hem27ply8cNBelHC
DCQf+WAKZ+f86ZAPSR8Bp/0fFjihCfvkwEYgWcB6d3EmsY+lM6JPBsmyXxM+BzxC
DGmD//kGBsCRxT8O+S42IP3scgydlwJ5MyXFCm6D5GUrjHOHPQ+CQSu/A8jC4SS9
RKc0OOO/3fEwQyCBLWFd/Wlx4au64HTUFONMao4CG7uF4h0osFT4IT1ZFdfvG1xW
J5FBlE8502ELVECzXGasiLol2L5mV/dDaK/Z4zJX3YIrDwrHoLSrU6cwCc/TaRar
b53aeWxBc+k3bmf8QJ+NEKULF5JpDDGMu1p7pMYwJxy+VZ2DZfmeFlOXgIcwAAza
cjEGeRuFL+De8MA/JZyuZEHshgUCNlITuTQO2o6bucc1Bhr5CV2zvesCCK1M+jN1
oVU7IaEM+G3M2hcmhaTf7PeoYVeSxXKysqNLVNHFlAVoM2ArU3aD2o7MEXk234TY
AA0kIgwoppXHUo3QoqXZWG//LzVYPwttEz4ztFozLPzvx9FD+eOzYqp53dQJwGoB
sqXSlya1HBUKYllthbG9H76PomtsTS0KlAUs0Vm0S3INlkoWGZQY9NnMSTM+v1Jd
jSKXvsmVJ6QRL91zhSAWSMh/eeiTD6Ha4VxuZH1f9mQxgV4LW5jlF4IutbCHcb5Z
DWwrRgkdLtWSDLSLXuhEGYtFzyOXivhF1INKBIyGs486o0ZL+UETYao6hQ74M0pN
gpL/1NxZimo0O1cj4DIrBo4609YTsd/7nKuNeUokBMlYgzTzzrCF0vwPBaoFTc/c
iTiqFSkwDXhD0buofALmh9pam2SF6UMlPcSJfmU2g8rOVdZ2bU+j4S2X7haAUDb9
XvYLfJKsTE2IADp8kAi5vkcfeOTk5AlmEQmJKz3e5t1fILghBFkigSpz7DaxHr2f
mSobsHqZSa0VJS4ZdaqqQ4BPQmCbVmpcNdeaNNrOmO5NS8qlQv02fFRey4a6cwLe
sLo63FXBij6NXvvsjhNzsVu9/a0GfHc6JfbP0s4W/9fr8/wGUHR1pr+0d+aY/1sD
SaZ4LnK5xCAp5koJm9yMfQrBMnvYHYCbNKjQOg9u373XJnN2gYdAqS7XOnY7V8D5
zku3m/LdHroVqqf7aMQDOqC/ZmXr63XmmNwTNZYlGIXTCE8pHZwrMfwX6+ED/sql
R3wQIh0ZvT/kwY+Ap466AHY6jmNMPk0JRSwpxH5LXZyRDhp4V11XEbSLhMAhLCzV
SEjhJVYlV9ZxvkvpluFU8VZHY+8tOd8gE0qhjKzsST8FZ4o5tAGG1Bb3bJPweP16
9snN6sCs4zyVAWsIyETM/5PuqtDiaGDkUWf5wG5joDACdgGq4sC9Rs9EIVNN2hJg
Kw9dd+MINQqxkZp2Nm8DuPkEH8DkKuwKRBUEz+L6dPly4GEBq4uJ6X2U9bH9DmzP
5Ia6Xj6plKTm9w+wUZs1XQNEKAIKbzj+rQkW/J610qAVmopU5+M0E2oedseyxHtM
UE85RsdqMsZPDTBXeN6PEgmCSsty1IRwy0phEGBiPnf02n45WTkkRxStuweDPUV/
Uv69ueHUezXW+xVhzrO+hOD9sEAmngq5+wKG7oZrM45ShzVgTovGJg4UwCJHjrMt
Teey/S904K4rAh9fzJpaTirIvGQ1rbmDPR5zZ97bDJtZCvqv65k0fvTWQOfFWiEB
wfXz9ck0g7DtSPU9G931BH2WdPrQlMy9r/HeDCdg/a5RUlvMHutYq+PSTKSfKVIv
9dOoB2oieIPuKglsEf0aWJv6cNHpaFXpFGA93jMLgzxE4sn4QyzQx6ZTEz8EvMYT
wK6veFFj4GGvBHzu9WQ7taeObCbtngoMcApm/lW97zcFRJVh0pNPsAEh7oOnT8Rj
hiUUs1zR1g+ArDVgms7kxBaWPR9U1gA7ZMmCjYJW4NZ6BSlcgT3YBNLbqn234LDj
xTbMIBnezkd2K23UrRkFOZx+5to77S+9xllVOa401h2wUje7clJ/dYpx6riZQKQR
xdDHX8PuUul+aQoPP5sySTU3NZR1BQxHn9PyMp/w+FhIjQbA6lUVvIilsK0W+DF8
QA4+BM+z5MYCRkCV0RsOLMwfDFv3VCFQYo8KCSr4c+OsoqZh7n1QSb4RysuS9oZK
nRYifMQXCugSYwtMD6XaZ8RPKar7+zZgGcxz26n9hHKJH3L9ZXELEmJSZHMJzRDV
FgnlXfXdDVazk5j/YMMH6b028ZZCqr2+vZA6zzkdqdIj6ZDSKAVYahw0aM2St6fN
X+jVUrXFNhjOvxaMeIMOTQXjToMWMv67DP7hdoczfwBjyOB2b7EZN0QJUfkMYvSk
qBddLLBThS8x/Wpnryl5wcB5tBUtYYYa1jMkf3Bu7R5UAW/jkfLVEBT4VDqm22cV
b8ubGrgu6bkOUyCzMe2LeZvME0LGT1fGcalZ+2Issi5wRQ65EwWCA17fxYb/6rHY
4UbZhV0x/7GcN9/T45/eGmEbbdLJM+20CvKmdsvInLpaQ+tMtKc7xd2+qrTalQLX
tSAXiK5O1KgZwk0wZgGXTlphpkobwSuLmF0mA1qDOFS+sgEW12drum4dDtT9r8cr
gEtAx5ckCZmJFo02yh1vzhCthTMwVzGNUQ77Q3A1J0ylpG3qQrGz3KoQ7ixkQO5g
cDhb6W/Y7ADQqLmCTWBLkidZk6x/UTq7M8pVkCmhNsihhrsxL2KDMj8IgeYzBMHG
l1GxuRXeVFqVK8Z0Om02zOIJ33K8hu32D8d2KNPtASTEemYhtDb6+ZaM6Iju22ml
mxhU0RFGdG98rpzSTlVj8yNiNRoblulftb3cQnYm4Tdz+2CVLe40dsPj87Ag5rWR
U9eVumVSZRFsQqs6iyLrKgDIJYsIvKHVAKP2OZE6Yt0R8UKEwflpmIYqOBEilEIj
WaecIGXUMOp80E45zAPq6eNduLMZOVbHEWYslC5254Opd1sgdPjnPyx+3tfJI/P2
2aEMv5AEL4/vZkcaaGcId5ecyIrqmsDsXIRKdytethaxknL1KArAd6V3IMRVxRle
aPOb2w8+c2AVNnuFGpHKuozoF6DHfap3de3kCamoHLmLMxV5JKx2SNqAoMuOlEyC
C3ddjtzEXL+yAg4w7gfdquCUcOJYfth5HLWWZ4hISeScGUVEewvUtb7olpSAmEaC
vY4m4fQmzkt4jNC9/yXpFLTGsmn8VdqkIdkKEg+ImQ2xe0RkovspZorbjYr54Bfv
1JStKnZC32ILo6Ugg6U3GGPvXhSHHqDiUkTKxKxiO9UQtTplFTCwc+tXIXrh2K4L
CaRLfj7ehSpIZzic5JrQQdFwdOn8v3tfeuSYVRplVH7KIFjsKuHTg6fNAv+n+xUs
Hsw5CNa2yiXNRtRbPqm8zaMnHmzwQXXDrYJ2z+/Hz/m0mjeDRPFwWn2EU/UP384H
9WujJwNakXCjI0UaJQMhwGm3eyP3kKkVboxIL2QIlq6hfWfhDvgXt5I9sAObla53
WlL8unn7BFSvP+SCW1Ki3qUEHa671icv6MC3zjE7F6J22gWPQnrgJ0iahsgJbgqz
nVhcNZuQx1+xhEtac7SxD/M+liqUSls6CK1ma5YQwl3N525dwMTX3S5pjFJnecc7
HcZACzGQTmpSzw/N94dqRcUcmVgvHQjedvO2ljc7UedO0fx8kByFI7M7YvkjAbgl
KfFf1Wiv4x9i+ZjEn13HTxZyl6oryHKkOf8UzZIfOdvrK6SUy8BdqeNRS3WByhrZ
Nmv+mEz9ibC1RbniAtwepw0RQOVvCZHCRpDKcZVjn+c7Xpkq4qOu7cxo8t32G/tS
sxRy38M8BURYDb4tmONoVKRLrujTD4CajRVBiY6n+6A5fDxx9ZBOTNZsTxifYi5I
GFKvAwhBfiJaCMsDA5U6sszodsVStaeR0VQTk4b5P1quvJRdr+mxdmvsMGPiJt/H
obEm6/4vVAS7nyOeXNHoTufKEeZlrkVG5o6ePDETkL/Ckf3Yn8YnJhBDXMbLvRZM
kv4cKzz6WGQ1b8YJGe3cNnBnVkNidNC6U20uDlNJCDuxn3o0wZR+23fFUaaE2YkL
mTkiyS7al37cBZALKglOfarY3rfPyoVLx2GyagcOFQGp50s7821t/glPxS79sN0b
w837rtJOUrjoXyFS5uPPM7vmvENpbQsnoWZc2Qks1T5NWei0Y89g9WFLVdhtT4pI
3CgfrC5L1h61GqvxoGFnFu1eu5aYJpkrd85Wvm8g0yN+DQn1BPoR99QQTVoZX3+B
f5w6Ih3HyUEQjFgGvPLMypJDKoYjnmEqIjd1RQbgfsx7W9r0aOkc+ujSuzPuHGlv
xRQMuD2fbgxYdugvAOnEzyWmZoj8LrcM8BqKIXmvcvtiN6SoL5NbMY5oddlg2xpC
eK1RLmbboS/Z41PG1xD2j+4dMh5fnB8DbtAimR0iZGMWJCaRxBC8nlY/ZPjnLp2x
wjBeTsoLIsV4MmshKYzMbxfgeTDGlXn+FUpYzZ4m8s9QYs4SpHAAm5ISK/2gMZ/X
8yZKnevgC7g4dU62PEKyBV5NBL0VeJFMgdyBhl98CNyU4r+YLXp/RiYOE+wkJ8rd
vw4kYOVRaETDtTV8G/9e7ZhAcVt+Pvp/YEIQHBZsJeCZiRc1CcfEtw+sAwjGZ/pO
y81CX15l74L5Ytg1UhJ0Cb6A1n+V5c6EMCuhJ6eBvxXlWWt2eQjrB9spdNcxZ0M4
KsafFuGC6b6BW4/aekRELZo/5qOJftPXvVBg8016JJTt1ViBptMb/rC2hHFSvJ4E
MAeiLuJNadnOovGr1lkR4EkHZYO98qE9l19qk4Qo8B+GovzXEN076+Yj6VmTzrte
4u5BpUS/vUPKrXQFqrBwhJ6i71pKIiCVKVEJvpqeGlzcs18LL0Z0/TiGMW2dk/QP
H9X3+MXcwM+esEraYk4HS0h+8CeCyf8NJTt7XzZfpv+xNErVTSZAP7HqBRfV+iJr
6i+jLISNTmolhnioB0nkbjZceRWjgrd62ZswG4CNhflmbwa4YlkXsb53QctRn7K0
dkjXZhLtHX1PmVh4fkt6CfZ+4Ki+ivpFLgZ2GcFP9X7Qfd9l/KiEOpRJISCazi+s
Edjb0v4fZjSmEuUOR71tpSRoVwlqtWKkVOpiTOndJhGBSRauvtr8DxQ+l4W/tbaJ
wMZCsdTZsV8/9jmtUokGmFqJAO58E1EYKKsRutfLAX1R6l4dbe4E6y8CCcmzMa+9
p5AxlIs4flGetY1FNdDCYqDSlZfODZWv9upfw1iSkkSr3X3mm70H7dcLqkH8Y8/a
bmVtXDmJh1vSODlOWTk0lm6PiptftBCsJZntjUJeXzgSf/pE1nmhSEm4pdrdretH
GZCeFrbOYr0Wjkto3agj3dKV91qTar8tGyfFl0WuHGX2YWZLOEH6PERH/UHo3lKU
Wg+F3V1+23nPOBY4Y1+NK4X6V8v72Ur8u7cmxj94eOIKdb1JBQ2Omry/6ebGYN61
EJpvqMY1NBDnyT2vr1Lf4d44qNNc8cd2SJ/x2Ti8iTOq2tDaBvsjDJ2Dxnou0QNA
rIt2Ha9JlC5MwfVPPepix9FX3sLAyZNw6deNh7vSe/jE6RT7oP6jw7R8IPmvDmau
emvE3jT4YTMJ4Rtk1WVAohoOf+zB/Woaj0BmFq6rW1OF/pCRvAt2g6De+OLH7Udn
hkJUr/8M/29sZnd+Wg8VdZ7iV6JyUUAS2a0DljfYxSIQwO+BDPZKe1ZboKUnN4NE
mxzTrYLedApSzd4bd1ZPHbSOsM6VI2loIRwUEsc3eFksy2M5fBndtJlA0ga90srZ
VwtcPrMy3BXako+/EBNOjX1kWpBcfTtDKyAhPtsuzBfKb+wQJ1rIdqduipc9uzl1
iW0LugRkwE8Zo+eTg64DaKxJ3iClKWmtBP+7ec/NeAXSZg9C9oD6ihxPWPVtztNe
w5xTOWJSU1gHXrtGWmZncLUHQ23bIk8PkMZIyTUZF1IEuroPvfKmgEJwANL8b+n0
DO6SWF+g2JD1OdSr28/P6aohReTn1Qa6TiayZllGyQwWqebd147lLWPiOsQ5VW/T
IAWjGAMloyZNugAAYR6d/UvTGmItmgraGAiGfYg4Sph4UrPUtfHU7L6IX72e6FZm
0/69m/MmrR41Z/miv62ei+bTEw5x/Y7HXcKp9V0PkrU6rWT21BAdJP+pd5Ld2T8u
tdLJW5v5xc6inMd1o5K86t5kEbj4pPwQGjikHYGS5JGo3iVltyTp2nVGYYipwLyB
zUEl1ynozkN/Cr5fMzC/Zr94E8itUUc6OJqmIjARQTOhnbI5+SWOtSH0vbzgWndm
JtnQcsrks5b4aY6QzvKf09dJhPsst2Nhk4+Ktf6xWWxqqlFIOAfN4npPatnAf28X
KyNxIHN0RkW7oHSOj4pPAJq3zv063hCvwvREudTZDMmDqoNu3ppJuqAtJDJzKHz2
Y+HrzHY3PgbFrQSHDCEIyjr0co0vwuo90LwFRn4pBrWu4mdX0sK36pfJXtYOdKrl
uWpSRpkN1NmqVN2Eal7ztZLfo5OkDvDjd3cE9L73bGL5dH17nBVlHAJDlHp2837I
nhaUjUZbfNhfDg6HG71FpZxQfjHrO91Uns73i91KdvdvWiNJ5yvnoVMkhowxpKZy
StNQPUYx9uNOzt/edHcJpq5xmXp1kfME62MeNukLDllVRDykCJywIKMr36JaktER
Gx47/0lSaUWj2J8UVRuydjmrpILW8kafeyQ17aw5Ty20igNEGeqn+TADHUOAtb8b
27QM+xSDJk9sTQuZd+9swbhhLcEILRx1eRIFBmiO1sJpRgOmhZ8zIBZ/yHhmbOCM
3VMPUW+b6kgtzISYEYeacLNMS6nQNWRVwubMYqUKvKuIK0127axYlf5CeWrutCI+
JxKfVRILovATC8xa1loMVoC4U68IzUZvP4Tya+5AxUuxEeEJ86F8/mWCG8Tb4c1+
ta0PpqjSzxyx9l8+OAIZA07WIKIQRGFWHBR9rRDaMTnJ7Jdl2GFZ5422OipkZBn2
QWVsgZ8r4Zs3xCWbTymbudDYq6sqrQphiQaODaJym294BYsz3QstZywDh/pyL7V8
OMXNjRB8YHWPejvX0AxlBgh3DcnVfAMU8y7QH8AAYJMCP1YkZR7YoMJO3XSx0iol
TzYTa+m4ITy/MGIQwebUk5HnBA80Yv0S9ho4zLsHvsfLAHlgV0qSiR7csgAei/7w
+UJ8+swFHf1mChW6FR1GeQ3n3fj/ntkOp42DnOTYpVWvVQSrL82PimUmId+JsOcx
zIzJxfCXOc0PE57GCJx41wJNP305eDBlmV25wGQgv0z2pnBwi2/FCejJSbjeziOO
kMqR61KlHzWKEFkem51YShaMTMEshKIeICivlZbYTOVfRotoRfE5Pwy40x9cmitM
sT1eVAlYnLSTdd0wVFmkwu26CYSmsX0wm4ISjQVB2ENN+v1IpOWgGGfzTYBnWbhf
NUsskV0/hLh/FXJ/FPn0hRQYuxtnZt2chYqmGDfF/9oYOEl2It6FqFDAHz5igS7H
YJazmOf5vn4WK/+YLCoXWAYa9UjBgKp/9TbZLmK9dv1cpBi3n0PNDEgBJPjXCKz7
xrPLri//RPtDtNDF7IucE+9uGJxuKekbSoI6DputQLbSFGPKMUutxbm6MA1gLxNQ
TFQsCjPSzS93CjvQiZhBkGq1ffgWVcNfJT+On/blhpU9CWvIpbH0Q0gqYaguBTjZ
X0yzK1k3qmmhZscrHK9VHxxtmJyZ2fK6lt5IqeebB9iEvxnX9rHpjtc2M8YE9kPY
G7167ZuouNZDPue0ceMdNPKl07FQ84d6LFFy4DO3MY9nka/F0KSXkWEmqbcpF7wq
q+dK7JQX+neqf+l3HNlrfUQSS9IwKqvs3gEmzWSbAuQUgrH6Klf0GyiP+B+Sa4TT
D9v1bAXBg4w3VT5qHiMhSdfvK5pfRh/SR7/1uR8R8eg7rlPDuYF7eYqhDVUNvIZ1
oSJkYh1uhHvh/jRs+uc4vGIMaimrfUKVHgzD34wY56yDDncQpgPM2whkCIChJMi9
iHbImDjT3JsB/lwMuzTggtgr5ICIi61nqSMBFAe94WS5gyzKrh/s5dRPods99pAs
/w4mterlETq2pvw72ZFL3SV0y1Pd0kaZXjCkP1c7y+GL0p7dWFac9mpxG7bXZOfu
uM2qLkIvQ1Ye5t5kFRTP6BrJHYvuDVZD+dQtFaqZdQMW6+C1zt0eYVpuMPHN+iIR
kRnxPx/g5Ox42JvOL8dp7e07kNS/0DkbgZ4YsGIY/Q0Xefyt6RarkeoDUKyTIUZb
ydDXUd4zEwafY2d5FNCok2A7HSRXIUFN4LyXUZ/kATeDg4pFWasgEz1E8XnPtOWn
SXEIMIbawvgIINnzmLaDye+Zi3vpLxhfLifn4G5Bqaun+0n1emUE67cnUMWQ/ZMo
3t15y67M4LNq76yeG9mPLcsd2h7mwjHPKugm/9MJFaVlfl2iyd1Jj6ZvmohIgxxV
c9F285PKDh2J+X8hIX+BxRXNeZmwjijSJuOHGD8R+jdTc0S4uuJfzWi3gw7rR4J+
c+e1Acvd2CRK6SYT1Z28oFNyjKDPgObJf/9dp28AwPpUrOkbKCx1oKUWCTDdVjs+
dNYhI0HO+ic87yRVrxichsLLDBhL946B2CgKQzuStrDF/hP9MKji5nBZEbs04mJg
d0rt7SC+riXohaEN0TCLb4KT40zoYSPSHnHMDZBCpknOZbBrXRmQyZv2Jv/6TaN/
03ENZfndYrZ6kJ8HiLPsuaWolLJ3nEFJPZhSY59+2X1Mz5y90TvBQ9pRvkRSGgtx
OuMZPNBtnzFkSVTRs/mOLq4nCLr/il38/payoBNthEQAWf70+o1YpK4SuXEFYC0e
B+SIu+ZbanmAlP+Y5K9HBP10U2IIgLLp2FJ0MlSGjhH9EK2nXh81On017HbAWBGo
A74ymS9Gf8xOBRCZsd6+e1QWXhXkOxWHZFAq2pPdwF8vaB8uYj7E6NylYzG+R7iX
y6dZctdwF97x6gsDQr7f8O0GKcYkecewqeRE57wtMCoFA7e204DfOtV4W4H0ogZh
hH9DyY+aQHRT8Vp52dPyiVZ4Wx0WoQkT7MWTZhmEHC7pYIR4/aIcvpSF20Hb+Qve
URO7elnpP/MDisObyeTr1eFSLH+EdLvY0vZQAzaYC3yQ8p97WsTO+xkucsXGEvft
5MbtABT3AyyZl3zQLXshXI7Q9q+k5efU5dyvJQHZQRkqCsTZYKhlwKG0wYzIewRp
yDpLrZtiE3SIPVKLf1unAmb4vjhoF57yLn7LMicYt4If/RYGKj4CvJwHrOxHh1yo
uTyhxAl/fJH0XZyo4lLRKlBhjpQ1tlW5hqJLa0f2T+iMm/e8NrowLoLDOiPGrQJh
QxGL/fv0RJcAKzxMQ9A6RoAOWqWL2lS+oQH6euyEkBF2TEK7s6ZWPi3v2IQubsAx
CNRxDXPOX2SXvRU4ePaXj0Alakgj8ObQbY6Gh5gQD5g4EW8Kyru8ZACRMamFpp3t
gPCd/PSLWKLxRbRWripzPunB/4CfwBGQMoiIC0bi+PgxkkIht+jmHnErFbKleazj
Hpm/7nYWQIFqx8ITNw5Oru/TzsTG0DVFc4UoNrk7jVUIkqgYVRYWQBB+HJ2SXxiW
+A7rwQnm6rFs5kxg5d7fxiPmBsiVsKLhhrpSuGsfX87KUBq7rpp+rbPYSuPHwLYV
vHNYfBOL2D9d8+QYmc7ZV02IceDLpAi/YFmcE3Skun1EOpILoapfLaklEdkzqJxp
1pEcRunV73AXGecYnhfMGp0auXlWB0rGKfqq4afBSNotsFu1n2NNaBOwEgczeF0U
iVnYCCLYUUc9lb9pxK+lb6dTtxh4EhfyjHXozEXKFFg6gdt3mQTGXpgqOnzqAuO4
8wD7Q98Vb+GBAuRUTMc+Uxmi9HdBpMaxt8N25rCmqvao6VOmMnNhz35U91uC+yCX
4HROtyZSGz0SEXEx3qfodnAOaHIlPO3Pg11wpSJwcL5bxrG9T6BjEd9/unzYYCfD
k+CFIY2foS93KBho5I/VdF0+Y/LqGZBtbt+JHgc7LWy22HOrUmjbe8I7uv3hn0qC
6ZXlJ9cSRsocbvA1TkqgcoaqoQXi7SZr7EbmBBQi/ApHGACU7Fa/hJAsbma7dt6F
C/9uj+/ibQxPG+WvG3K6SnFqR5csTDPS7Wh0JOV7LQ//YdGxU2xGADe470+iFBQ/
diX6cduJTU++lrBkMJmp4ag7BVNinkeWSoZiXtVPyQx14mmu/kL/x4U3EyKxUGmw
eXbDtwFNZl75pzXgPiiScScOhzk0SCU7AeFHanj6Qs2BcrcKHMkUrffN1OAayM6L
/9/V5GQkGirKk63feC7uQcdKWcuWoTq+CJqTqmt25fkfN/+oYCABfbWJIOd78nu3
VSOhDgoSM1rdNZQ0aCC6Wj73p4IEANxHj4WwKu18nuUMZ/dgzvx87T/ssFaOVyxb
Fma/4orwcT8ftbhiM/KSaMi9JfLyKDzKQBqy2w6pSDBN6nMhQtjMtbTc2xH98b1j
RFGdgTzzRnMOkxj79XM9dDJtE2soIZZrecGXziSzoHQNtRkSkZHJS8D72jkyjdX9
0np/ByPCqMAdMJpMLvZFTGBA+JhxL52Q/7onPRlfZT9CinXTkEfQ1RwxNTcqTwOq
G/v53mJS8deFqzrXC2Hadv3xfbOqM2mAlUUY6RT2ZSOgOnDNRvZAn5+fLGpkgqy5
VzCBiuAt19QqHRuyY4J+EiAnf5YX9gguyfSDzGhumHncyw5tdQgFhU+P9s0YyQZD
KXdItpoBL6zhbsz4yFtJLQY1DtjcJz6e/+2BAzvJg01SLV9gZBl4rujQuwMyLJHO
72LkEnTKTUCAJF3y6dKHWgoyNLZZXqlbMPMt56JrEla6EWj8ctdrcv1kd8quP39P
Jy4KkHGYarSHTliOW2lv2CRlayY3VZ//QE+f3w9B5PbmSw3cccTw5VywgJzjwLCG
oR3n8COxzopQzfnxIEpyCf3qp0WETjxY5z0djLBDCitYJhSA3VG1tScIN1u5M1kZ
FJ8GqSehEsBPaPOXp6aqUFrhTwWo/Q84xXTryVnsuUqg2uWutwHePGQ2DSkm/HuP
fueLzRAliBPkU0E8m/edPoMZQ03yJnwyr61jit2U7n/uHBI5cITp1w1PGE/PivZl
J/0i80eBW1U75pa3+j1jhzZDK5q/2y8NYLI8Avgb1V1rkHHd9PpAz3zTJupFTeGd
xCpaVFsiAZpI8133Im/M3ZTaIeiJ/g7ti/EYpuV9XRNSgIm5YoFdZpE2zxrxRdYk
vVRVCZle8GSp3IjDcBxyABKl8Adi6d1po/tSIP4hIcYh9q9gjReSwKT1ucL4cT+Q
Df8MPtlK50D/2pa1T2xrjqebH1lje8mgYEONpXBfM16J7+90wyhqIgiTJmNXnm/2
2vGrrKCeY9DbSB4YQa0cYf7NLVs5yVQ2dOXTq2tlfPWrQwRntlMVUIFrQXcccvvE
sBBhokaI5hsinPmyZt03LwiuHqjruKgdUwwNKP24GTz0IX3j1MC67h+AQuMtpr1x
6mXzdEyKnDJIkUTKeBDNxLuGFGuga2xcJaoqAPsaRthcE5UyHighdoOYBF8IaB4L
LNTg5iziXeGQKFMKJBXZPiO9WpQCdLxX2P45SlBxi49mUumK/CqEWEwXEL/Bm/RT
NqgBkqZZ0F2D5/2Vd3b8LbxPUD3GaGiBEoXnIJe8XrHpmbPLx3YeCWg5vF1jyV11
fYVA6p4ayD2WHDPItjWbF4zHUSZRvnkPG2qtYanMtXFvXybYMpbeiO7aK1lCvYwp
vhavUBE9Wy+hKWpQN40OchuVAqMGUuLIFbZ3R3GzcO/2Ba3WLSctrn9u6SX1HSGd
aZ+Q9YE2mpV1T0VeO1MY0LU8a4fIRH7Jn05CNzJsIGxVlLK5LDduM6h5BVNmmT/A
8sZL/264OYhE8jifmdnfe8RgAkm6ZTGbCi0BH9SPfIj1rSkfm27qzljhHK9iweFA
Pw5ddq96mKn9dBGptMm1eO+20AnnhN/nTkN1fIZve2huJlNb8Rg3uwEPws1UKm9L
wqmuyNIk6H5EZ2hO6On913+O3O2xhXaYIoTny4+di+fvDVfrrlLuOMJ3vy6XrA6V
CzZMvzz3Y0vX9MlltSR/FeE8y3MRgjQyqD6bud+mcie9bXk9DlJhiq+7l0334YG5
h3eAt7OOnJ5gxbe4HS250cVDG2/LHWieu8L+6LUkkP55rX5gUexftF7jvYk4bOEw
6oGfgRArNRCG9LM8zz2giO/XTAd8Rf9atF2s2XTqHwtNzEIeFLsFn0GusJFmay1l
u+uF6Q/H27fuGv7GnJ1cs2+WObD1v5WayBI5NWcznvmX14V1C8AmD1eAeDh51xCv
mOvWcatLCEHxDjH77RRjS3y7IhDMHFZhyK6FHNpfUi7m2JYhJyaE0e+mFQYoSyid
WiwWT8HrDftTHHxjohr0F5aYDBcwb8KLueLvcWOt9HmEBFD3MTkbT1VrP2r4+O6i
xerdV5YlC/LAJLXBUL32/r8WqoMPZL15s6v/0C56Q9At9sC+QeZzvv4LxyiCBw9S
dkuEo3BeUX8RXaGs3IK5LfNkKhenBbTuczWQTeTWgwX2/diVl7llUR8TRQw0DuC6
6jiOTpZSeWNn25PsBBm7Bz4BqZWrGmmO+Wb2CKg2MBoavDIepFQ6/Vbfs/VcC9Gv
04unYwyGcozYDPNV6Ya/R1AmjpmLvmgNMTAQx0B8OHh9MVF1Fz7HuUdrjr3XxMWj
OaHV+zDWl96tDvS6Ov6Kjdf15Nb4SdSxdIyERDuAsu3KZdqj1W0VcUgXToEnKKqr
+WROSn9ly18tcw1x+3qZSaPx5W++Rr4qG24U2vJGLwt0fhIeet/XHxm+8hS5AWtu
rMK/fHljCCQ4WKzGL4nWftwd5GIGC5+3nsrltp7a8R3TNsjw81oqY75CtJY/p9x9
n83Ze23BrSMf9E7U5oVXiCJup8u8jv7G4zivPzn4rkw83yWUYxHpkJsvziYBrdxZ
gicTLwwXAO7AXPmKX1TeAjKR5fYUGi+YRw5VSNED1jKiJIY1ABJbUbjeApg379Uq
uCCnaJ59Lxno/mDXOGUIMXii8vJ+jECOQHO+nvv19M37sUD4F5UOGtMQffeaAg7n
aDXeZWqoLfUuCp67NR/6Hl1DjGkNrHeTEhbzVWWhknIHvc+l7hF3zpuvh7bva1lW
GWIhyFOkDdHL727N56qbvjpXvT/oxrWMcq3439tbF+NQsb5/RAMzSzOraYk6E0HI
RxZQGB9TirJP2wNvGx4RQpCcbv8Q8JKQka4G+R6+OI4XR9y8ni+JNjSvrJI0Ait6
7Db+KMokS0JBuJy+MXO6MgmJas1drKnnlEJaAbArCWBlD5XZx/NETxRnLvl6xzln
fOalUEdvgLoVw+I4bQBb6efncAHoWwVyrB0AVqmUzULF8bb1qqlFIZ1401gJxs7J
so+76phNwExG50zyJxmtmUZOKqZqfBAJPNlqrqxGBw5UmlShGCUkfE5PjBMhwGYY
VbqsSyCNfVJQ0cWPb+j1v/3BnTPlKJFNqPWQZP0XjJ0LyXm2wmYju3fVQltUqdlm
ZoJ1RCZPveWVSdQD4BegegTNdTVCBAol3g2pbwcxVZhlfQpW9VgpbA1R+LoBUgF8
tsYPPueWc0mGwJOiBBTQ9ia5JtgjI2BYwlAzd025cfv/UWLHi/4cYyRF/8ZmkTRs
ujhQeK9Ml+4enx5BPga4/LnSlzrfcmz5JaIcY/ZIheRSePo8xnOaQ4mrDqd4Wvn6
aRv6ITbsG9kd/5eLChfbFTtMifngp3nh0U5RoTPRBxNwZpNi0HVP0BMy1HvrvEdO
U/b+wLUWndUnqYvK/XS8TwXCoYRkdFtzf4skVoabwym6GJVd0nqAC6pWXCBi2qha
Ivcw8IelITM6yaGGKmqKegcw0gqoCMBY1HMun2Akuq+xO+8TjLoTxAxQZbQGzcUm
KbmIrjX0E5sr/UMQtQ2yXrYw/3iEI6d5FTlpT45HWzOwL9yXWKq+e2/fNx8s8KhB
T6H5dDVFg0pO0ZJXfTffBYXhzfczvZRR7r2ojBMwjV7Cvby2jQ/SF7GZCt7vr0QL
9NXydMkIULBmKPHxP38BajcKmFT+U9LvIAbKezcOteVCaG/DT5f+rEZqbCvHflFX
CccegbfVk8jZxgWZzYfmAc9nXm3XybCTw7k+6CBi+mSqdF8LzsqsR1X6cFov7F2c
gGcy68DF2lISDRzVSf8faN+HjoSApP4wFBGaiFFMhmYZhOeykpsv9gbJIEYnTIfs
OztAeOVYgyD2AgqjWN1s++YMUYADic8Z7H0Bbr9+0U7zRq2OFKWmJ7EEgARPpVAZ
8mfIDtQOo9taRCd5nSiCV197Hxo+qOO/RH3uUe0W5uWMpwxcFkuYmOqtDev/o5Rx
WLXgpA4PA63Y65yzNay3CqmP8YhNBmgJFmq8I4MJxSgwjxRhE1ThPRpPQK2GJynC
rvJrCA6AbxOS/oslq3TaZZkAoHcDAoHCjmxG2A4zJwypHe3QIdU4VMGWitUY4tA4
jkwkjRCBr1dRHynjQsj5+bVlVbIWGYWq1FJ8PzCdebDxBk+lBrk1u7WUPX3HxdYT
Y7zULW3y71NwnEn1jwv6EbjNe0mFL/vwPuPx85BPBWMRrc+wFN/mIoaA0TkztmsQ
7SumqjN7NoadcQW5ZQBlh9w5OvZP93vqtJNT3BK/cFdOLKPGud0D+6CJHp3JDWVc
fNcYoGgSBwuVUfiZlEaEtqVokrGpPg0NGCFve3Dg6TskHCArx5my3VRDttnjdRqe
r93Gx8mr5A42meu6VdeV/h8bcIasYx7MPM2/Yh4iYrNIs06P6l1/VvFS8E5FzXji
DqHFoFXElkCiUTJEl9g3DkQbMRHI/D0OAuvJoBS5k2LKqybpEjyzUcy2BTs00d7S
hvNH5LbsT4bFS4gsRNhe+HDZQwZ+7ppLjE00gDDQYCjd4+z1X7IykGJ17P2xW0xO
bzqOxk54u5S5SaWydK8ILVVGI+soSU/nXbnO8/S6arfdS9uzDSQtSd62wfWXFgAZ
Jt1dyBSUS9fwhQm1HoqdleZDhRvwKcyWDq5s+qV4xhRU0qs+iCkElVVX4KmC1OYg
Ot8ysQ/o1wmErfnWNOdM9mp24E/andrC6aQOS6FD/kcRSH7tlqrV2emikaOU2BEe
NCw6Vo9WHFWwH0T2TbpgSaQENDoQdkLMITwYHCE55JZmOH++JgyWsmXSEy1MitgE
45jt+2jhioKunw9jQAygdFdG4L+MU0VCbfAl1qFgEoJr4x6v1GmTTO5jP5Jxv3G0
35ACpRRHgI7cnnhs4c2Kva+hHSrBEJeWV0aqvgD66qcQhg832M4ahLzOnw2YPTAy
DrHjLR61NiCkSH7aRE7V3I90G1xbqchBUWuMJSWSU1pwZGHMrneDdavVzVZ6/vwm
zAqNtcYyLABFZBpfby9/ODnvxVmUn5mH+eEup5hbt/ol5Il7fa1XDLNW83Ki5qTv
1rs/JcYi4ueEsojv/bj46L6O6nI40ovRhbPxYRelvgV4cz4F860FfMG/Q+E/IqhM
V6vpzXFqLZofRk4hqgYuWhTFi4qu2xPp1X9jyu5+aPKh5Rf/vy1ywFT4tFcJbVYi
cR51NFBsP3CWTI46usXbfHZAuqiYePhSf3lBFf0Csa0dg1A3OS3SlJZO9BuOhTeu
phPk6CbIS8TQgz0l/D50yM1zfIue5pLYd+Uy3tP5MQSVi9TPTK0/E3uQEg2DS7B9
CSZkYp5ryfZSUCfvWPEM5/LjUjXEVSZUlvZmkgx8/WVyjP/FR6xkrb/IyF6QmOEr
BfliJtvePTvrOWolFNa6qMe099Jx4masR8DBugagj283mJoSGxk9UMqe9dNZ9nQ5
Lw8Z9IJOyQsYY574WCuzeT+tj6bOP4nnhmx9lrcePpy239lzJnZ84OleHVb6F2zC
5IpsJrMTZIizADnz7H6uQne/v1hTKYHRODe9HVsDD2i9yXOkXi9mENyZxKdLMZCm
7C3n6viy7B6yM3bNjw6Qohlp3oWGVKm8ublt6Y2idVxpNx0sCO6lPO1pOCW9BTMX
ET6+x6pR9il0WYC5F4W879N4UnpdqFJX1uxrYai2+eX8yQn/wMrpkp48EUw5NTac
XfdHopMsNmkpBdbGYLBZInUxTUEfANL1bpzvBOBq6EbrsyZt6urxsPDI5VLDTPMi
k28w/u7yJAKzcDzJGO3OYI3wr3WDc49fVJ7lsJub5ew/TBI2pH+5n6RUBrTYh/9b
J0tjIwtGSMATLzz/XmBo40C/7zuJGMGwvAEJXmORLCMKooZwmeYc0NBUPT/Nf1XK
JYM9MoAkTmhmsZo64mmZjddmHq4jZ75/qIkWXqnMHGgOxHgfSFmhutRsLwOE3XIb
NiHwYp8SldzIHGE5TIYJCmAnYH3bDKb+fmDbA+s2CqEf2yORxoYIddDRGWJbFygy
fvzpm3oDDwEXqZWdir5IahFStEMF4VPta6vQ6SJbj0/2g9t6T7Dy5KEGaN9F01yd
4hWxZLyCVkUFjXb7IdGkin72HXydRr+5KyQeiR60H9ebD5VgfiU/34KOvIUPe9C+
c7tkbul51QwsYgO3uDmw9KjP2uwRjQWRbEVI2IHoVzJ+qM7O8v2ULbjLEd7qH+Qt
3y75O8TsNk0l0Y39TnbhyGXOiI4Ghy0DM0C+M1BlHN5NZYMncMRr4sHomZlN1B0R
9geuyUNwXgOdXeDC+C51UQTFVVzM2X1+rTEOQk7PqMhAFdL1o+zmd14qPqdyZHsH
05kFAjRCwZxjDPK7LNm7k7ZwbMY7J7MfPa5nyn107LAe4p7dBKqbrK87UPStPJxc
ELthAUQz4YOJKpbTRm7xAPj8U3W088zMKsnWs17IXWudfwAlDhT5P6Y9JweZIGEt
EwQven4sQRH2rTnq5+XF1Rw9fx2lkKnm+2+A32PTNxNBxBnwVh/uUScJ9RUJCQHk
33haQJfBhi2dXxu7OwVlJmHBLd9w45//1NEzSkh8Ft437XARGkyqdspXk9P0e8Bk
wTQwwFugH+wYTwy4cd2ojvW6yRx0ynavbEr+/AVKDrbSvxNILC/6JmnuWGWdt57R
FahK0R/93AFFWCozk5Bodwuq9lvCO+m5/p7GnFbiDUs1uGZfBG2fWXdSDuogvPii
umbKzoIO7iOFaiSwC9nCOJ0hvBls2VuLMyFxWqYcZ2F3BRQh087WRyK1uJRISTqj
amA3nzu5LmqhPVDaQ3bJdQcCXZ1Rl+t+NlDYnZoQnLGjFActwUnRHJC4sj9ZQPF6
8ClGCO0nhDdsrqckOGgyDKBvk7kSJe51OZCRHKp8Uq5tizfxvCEwhwvtCUU0E/fw
VPIU+PjCTtg+eWIsxVQThX2wMkBLgYNDaybrd7W1KQLTK4Zh2BvM8JCVwnZLAtua
S5DQsc0jiWlTRPyNc/TDc38sW3619F8gMYvqcfYI3Y+8q2U2+qMu4iYdzQqic8ie
yI6H5xkDTA5yZzTthWT6dhpYfXk/8OmbGReEpFE0uIuQAASAvxVg87+t3W8yb+7o
gCTs74c2fARrrHVE8qWhQHoNbCUvB/0No9TTINS1UkLJViSEiRU5wsvs5rY0hjQD
5JCMuRYF4gFuCyiWvQQNbBA2Cwd1sxnO588FWw9M0CCnEawq5DbOJmatE92K+Mvv
PY2VNCaBCtP7a2gydTnKmhgt0+XlG9kvUjhWSU2QcDJaS3s6Pq3PQGWsfu8si8Zp
8/oqxgyxUxIlXi3jsRXosd5uSlhT0hrol+6F8oaJBDW4R3fihiUnxbcAcWhg5Gwp
QM8LrmPpyA29w+0KjPBNSbrxFIfBN9oJbL0sdigLS0+N8Qdc5WeegozdJBF/faRi
xLlb5fraqP45Gp5GThY0FMzBWvOPB7vNU89rygaaYprdkH/P2tejS2kOIFScIfvN
HQ7qmaoDkuusRHJ7/liHxQE8yW32+jXHHbBox6DL71ADA8LhDZkieUPkWvF82MgD
D8PWPp+uGfXdhf9szkAJr6nEM3nA3FqctYEVH/kC2sZ7UeVQv6lcHRj3EPVjni7/
nNkyQBQvYOAizK5gCRC/zDTaDKusZc5y2wyrnY9XjTLfRIjviU3l3J3iWOEFIm35
d6lxa5AUxEks7IO9doxnITwoWDhZCCtHM1UkPfzxNQ0I4dCsPgjRttvMVx0oBbwe
ELcnr9PYiZzNsOOZRPF0zZrVkR6CVM675FL10coK4pxnI/y360AvFkLWwRNAxX/n
0WH/1tcGBF4Jokh4hGic7aCVWZQdDBwxkLPjcBzhF5luu8OvlaHq50wzJuXwO3GA
wpUWoX3XHF7GKVx205Yvu9H3Q8by/1Px+3d/wvVkZ4m0hoYgjn+7E72EqVYqiIsV
oXsZQLoiEVNeQjREfGOvbXW9aUvLsCohLNTsSwzbkbXNyiFgnAW0SFsCP+FE9+Rp
PhIwTu+0d47m2h7gIQhB+e6fPqszgWuiwSVmpgDVbgCW52zLvMzoL1QykIb2yRZu
k7ilLfzjUY1dmCgJT2FwvAVL3hYpzZ2IdsSRyaDEKeuqLtZy8WKMKHbv/tEa0tp7
WrlSd9BCiF4mKyWkmDHHFuBaniPZcQ0xT4mbxcSFU004XpxcB2ua1LXW5fTF+rYZ
6MEpc2EmmV3oxdeAAsT34KyLIqLZRGH8mGaZrX6RhZYuKRHdYmT7sejnhVyuxyFd
HBOhdKaQvti3A2teGeV8HfvA/JoO8PHru+cN2K/4IoVwgasir4x/nLmcAX6bFzE0
eIAtEi9rOnX9Xn1RSJxyJ0J3tJWlW+M/1BzC9VciBOknLUhnTXeR623HYqv5GhQR
eabL+udsGZ8NNJs26WrCtYnu97V/rIyotgZUk/ErBq6G6jP0r0eFu3rtzUcdkayk
I1ykPO2ngCWmr5AVBIfelBNS5H1Ti2jGgElJdAU2H+jiDMQ25VCabBDIZPMWPx+a
+6O2VvHxUFknVX/yzc8DB+CI/Bmh0w9w4ZKMCNfIJy5YfqmzMRLkjIPTBKR+TQGL
1XF5pu/k+1lW3ps56RDRUFU1qzAcEDR58VsxF1fURcbyorTBfIY8WpGqk8tPWbVr
UAGzMm6lD+Y5hzN/z1jzRrFL3Q6dZWS1duqiGso08eqFLfUbA/FMTrK9SJhIoiAr
hfxMVlR/btykQ0cITwj498JRa1U/wPiVSv+aFDasfKGouWXenJ6CZFXcm2U/WJFH
yEobve76yBLPA6pBUn2fL7MjjVbTbYX1jUwcG3bWfHEeQX+apyrbuplt/1xcJPl9
XW1NPPc8uClHu6iuUuFPOaM6uFEfdHia5j+rG/9dAdEudVZbpHd0SN3TlWiRREd2
Zd5sXnbFGfGOdXh1vdZjhH+ZsHdH94hXpHjNod3gHdi67WdI6xQMHsQCsAdlyElP
JO1UaQ/b+YC9UKWhaAXC4e8Q4iF7jfxE5zVNAeIxgHShwt+4ZkbW5fyKeLENj+XL
/XrJTxnBtLhYkPqpIBnJ/CVGovqivv8jze3Q0vWxTZb/hFNgYrBNQITC834+QbMV
ycVuSzCZYdf0EQVJqPOtC9yiAmWQRnPh2UWnqxC/t/plyfBZ3h2IonA5I4I0qxCt
dn3M7RT9ON+EsqxNPZeWMF2K/l7Ow6L9GCAOgxRrFlHBxddG981EJDHknxmRAXO3
reNfQTtHriOvRmwgJg7wtwqaKeuRjePqW8zGL4o1izKJejPvJxssxnKQMknO3nP7
t8vktYn+z0YXwrLHNXi0eJOZMnvdBbCzJtBPHUo1ySU4fcLLyEa97TWjgUE3QSOE
WNdIitQQ7m8nGTulykutW2shtt43AWed+R1uy5Jyao8BYqaSKVue2lOLcAPgL7cZ
Xr3aNhQRSeEoemWp7cp4zuccRIoxChbMNURO7mZLfV3xtR2+jGqiVK5aOlDITU7v
tBvzOst6jpc8wGmL9TcS8zuo9LFtP7VlF403WTm2cFy6QVEw0ota6CnaWO4kvq5/
qMphMRU3usa2SzBfFrlq8E+p/9x+QAFjfpeVTX6OWU7ImfUQ7tC+WZc7fNArYgBk
VIwSr93yjkA4RcVShq2Jt9sZBMuymaOg0fE1XMetvvEs/HNeAfZhkKsKN3M/kdXb
nJ2aaNFiJDoVB9Zo5DAOKzGK/7zA8IL5SZz8KHEYBg8UXdDYn2Qi3qv0wbEORqHp
W3Mi/poEwlgJ8zWmaZhBQpIQVn3rr/Hs+DoKCMPqMHpDn2sTgodkjd7Jc+ETvpDT
OeYlo5hQJixHte7z+Wtziu3fhQbePfih7U9rwcu/UlQ9yiCIlzIGStMM/gOBh9y6
PU9IaYmrNZGZMM+Pq/HgEb1iqJvnQgt4WlFuy646oCiRax8CvbY7qzmk6bUL55xn
TO+o9aaQihJ0GFhEptndsBp76uMeQomllta+aA3Izu2J3Yp6x/FDJDCG3dpWLZ9/
dj2W4mkopHPMZLZBUVOi9b331asGljtyJ1tGPoyNCXiMXeVEYUWuoj5AKRtpQe+2
9j2qG7qCmbxXfcw3M1MLsD9RLloNBpGAx2iNczSqlqbiN1Nk3zTIctuA1XUYk0nT
57sgRny2Yq+oKWAKEsdUhY16R9GbAouceEA36sBr0RtMU5Fx8iushNC+auD4w1cT
oKNHtVk6Oz4Nxlc0ONGIyh5WrlbasXhsN1dsZpA5U29IzIKeiNeE/lRhAfM0InAG
v0O1hs1fIywZ83ateDrU5HMja5J2tY0YwI9mntiZbo3yTokMCcgAb8ivvMNAGU2C
E1SFTlpiYyxKpQuIlZdm4TTSQrtLz/vYnXbMjNRGRnwRc28hcn2gkOOtonZTjLu6
65YUNru8c2b5F9Ise24fr3RUzRKVe7VDh8I0Iy4TG4MARDTEqW12FqTKuKrIQ705
koU8JA5j/fWfkBzJ2yL2VxL8qY/obwSt5y5gsscK3JE4V8ZueDEUtfwQgESz0o+O
Pe9sw0OR+gNh1tTxSmSFBT0Now3XTgHi9m8J0JazGp0Tjf1L7H6MsQ+P53EI0Jgf
30RBTAVJCoa1glTiQxGkzpBxTDVEjWzNm6AGinVkvKkf/TmGzWjwRzLcRkBnu8H+
d3rxksj2X04kD4JNt3GHsD+rCiqXAdcNB9or0xP+i3FtsVZdwfvO0wzp6rLJppnO
JCCbCxRPBtdjU1MbqajRZwZDIFLHeXHDmw6FuWNCyHLR8I+vu2BJawMxugJuhnUt
4HirA78IpyOa8+kcRpqriVeXo6uXs3ye8ZSgTltBcDFr1txFRO2FJncn8T87fmx3
GUUjqYC4Bkk2PqPAEMqB9fHZNHI4NbtIYz/Ocn3cjbrh13kfa71ekkKUEXXhlEw2
2TtlBF6Io6QwsdOFRCvBw6RIRjIDiyFCWe6MEEk1cOS8cYZpLRZOoaDqz+eOGYDR
wVx5K1jvkueSBDOhZswvpFI4JihdtQYIzO9aCAdkXMWaOZKWdOgqKk7YXvUFUf3z
LL5WFSLcmu3aaMdncdvNDo+yWfTP8gyLqPBWl+Q+3sHT6CaXrMwcempwS3J5Ihka
99qhTbu+t4qxdGJxquAguA6lrh2flHEHhFGt5UiLREA7tPIepqmAfCSi//9Huqjm
tysiLJfKc0J3hJarxbIWMfQOHg9B642llaIxq61jY+pmpjpQoWaRU6uQ4YNYkCUO
u3J5bIqjVJjUbR/E9R3WBZTx8zH+JfAf+9WLe1le04sq9V7LGSz5MslWccjv2FVO
gkS3P7yAGtdTH5fBfC4wYu9bcED4OV2aG8dfM1NANxTZqKnst9X+4P31pAjdNbO7
6nqpdcbV+hHLrEopaSlbOIYc1G8IF0isyjA4jJfgGEQn8zbyIx0iW7RwqrRCr6Ry
a7k/OWzuBbAmELQSDYx/ao/UVPqlh1e0EphvQ6/5/quBBQqqTj7qMRQn7nC2A5pv
cXCmSpsb7K+FWK4PNVQHvuC/SJGODeCZyCC7drm4QXG+TLUX3ZFLHlOTGZ5/vksT
GEKM/IHvi2uEyP4o596+tlnfannLt6TaS8rXT3lzBkfYMCuO/9qptN7ecwC8Rp69
oZh58i+OuzI59qtc9vtHY7kygE0Px4dpk6WIe3pDXUPP61qV47xkk8AmGE303pb5
cwmSeXFhzys8RPlS6SO7s7FTTELXp11rSS5Qm/iUBI4iDxD04B8bkxaTssYiqoDa
56URWIKggfXs1IL9aVO8uaGC/dEoxNZOzo+V8j6iUcLub1f6taOxAF5DEcyJzlJH
x/2db+YA2bMHWRqCE9mgLrfW8ZiwZXcUc2pccUthBXJnpkrd3hR9NXenvxA08Lho
O073qpjIy6Mo+CrZDgcqAeo5AiIi/9HIPUyOSN6EHMVmOXdUGU8QT6tCRs+9nElC
/4nxXJkvzptlzKDEdWQBnFdkmbsbayMPPTOJegdM9gJ3w/N+Q0Xas5fRYyIbtV6z
M46BrFYtkP+7aND3dSXj0JZugrn82wN7VIui0HlAHzgivEuA32axn92F83w/TLLA
jHtTFi4wGkzEvLU40AygzSgEa6LPeL0POcjpG1B8+lpjb3ekg3qYuluhdXLDg+dv
UMi0f8ZZl0LXROmubOZlJtxchbAVSgKH770kKO2Gn/rLI6GbWpMVlUZmzGZQysk3
bMuuHeFg+yAbzaIr5wMM2LShyeAuc49b2rcwglNLjM92OCDrcZZ/zj2nNkGnfkmv
ht49hpgIif38/xnesZtpixGa9B2OmEVSLiAizefimxpxB8ikW6dqEG/olSZ2j+kC
/oRSkC1/FZ9owHs2MOVLFd4IfoM0UjXqHT/psxL1n7FuKGE5bGU+0hFd1GDd0Ex8
+nSxZYbxw/T59zsbisGq49vg8BUguM2cFu/YSQBYqhdCixNqi00m8z8ld6bKRhnx
1uVEFSJKFnH56K61wStnowViZNHAyNkisGYa+nyz3Br02Iab5c/SHE+Py6XpJwXv
qXerb4t8I7IkMQexqd+Ol/1gN/XhCHgTFDSO4pNelUskxSd5F4jxnaY2OrkVSdZ6
ecGIiF0mehaf8+b9yUrgax3mHZyfeGZnYBD7GsO1mnvIKq6oYj1ZHMOA/kIxz22e
q/GJItezG90tDVnYJ0979mQr/5jeyHq6LiO7lBIsMAnFQHB4py8yn/yBmFbrIkv4
Ghoh/85YgCSLsKmcw5m3SGaiLnNP2sQZvpqOAkejePIRdgSaSHu9PX3KmKGsWb/J
c8Pd8KUGLuKsbFLMIqvG9irNt59TkMUsb7NQ1uPeE3q9Su0HdmaGcoMT1hoHrCbU
Xs+flB/Cir/cw2WPkjGm8VsnfLouW6sBJ2oZisjaJf7no/SBJ/5uVlp1/HgNVGpN
r5qBupy3Omwo+/EeTy4Qd/ic+wKn/ZqaMzlqqMxR+OmBYh068GSUyrclpgtYroMr
G6Di+y3NYe4w7wZgxMSXRgTR+idTcu09GumAcKyWmZVVDNcqqDqoullho9x6PDWh
HrePjYpBTNOpUJ31Q3OeSpUGHB1BoGGhD50iwyEa5Xz0We7GNrCwToQ6T8kYyY8X
UvPrhmtMGBYTUYnmFe3u2zNRRxJDN8p0WeBUDQ2jQurC+scMJiQWs5VSJj3QxvEh
tOEbgXpqq3tgqZ90YL/VRsH4OartmLNFCecZ8PTFmXtViA8IaWDaHSz3h2YVHtdE
3iC3urEiB4TEbySyzGYzW0Y3QyYzOSqWe2zkvPQGCZytURzRX/cxPMPObYM1rr3P
tF4NVXkFU/PEOy8p5ofkUmjo0Dq7+ytEjzKvucB9bY+LghVH3ZmuPKTzdrNM+9Ro
AMG3+eAbyT0BoC8o0jdt7TY0Ln+tAxugtFsNxT3lmMIGlFPqGlYpKawKbpYpfz9O
EEMPGo3x4bJY/6iL+zIObMZILTsQrU5OcPT8DqGEWR9lWWqSQdBLu9n5jZIFGSA9
6IIYR+Whrdp5uVoAcop+ICCAp494qMtWzyu7VNi9Kl9aH26VHTCGmzGKgfPdbp6l
nqhgyMTtCKtkM3YNoEEKkyiEBR79ZsP9QqjWN5EVKJoyeB0R+2VegeO8kt7RqbgL
VZke8aya3xoO492d+DS53/lwbcrBUeRNatnzEFzgjLVLqwVpJ5rAk4dbxhkw23wR
w0DH2zzyQVvEJISirCF5Dbj7n5JcWAl4pokTiC/JMFNUvvnH6xMDQTBaZJczsf6n
esNPvYmf6pV74kNFU1WKY7kk7hdQwJa+oFNGtpvcoeOJrfJBvX5VUtVCPAtQ11+9
wiShblVh4hsw/NMno7pWep1+wMxBCPLJdrmZ0vx8JtgOk8KPFbgvyoB86SahT3tw
0w021yncOXPE+dzUbpMB8ZtaDSZzv5nhoLGJIBuhdMCMgczLCb+ZfpCA7Naro4DP
kUlNSkHSaKbDzbz56GF4Jm6AKmb8eF8Mo2WbEDEw7bHNB4+Mg/kU3+G+QwsAw3Q8
MFlJXxrHEq4OJTJ2J4/2t7j03vzA63EFbwXALbeMvTRcJnepP4UoSLDc+zSwUNRL
1b/rXQE1PkjUj7+CcHCceB2OPrSh1UqIu4yrVIkcCQ+NXYYEEYulnLHPU6J7yQCk
/sRJD4+6M/oPPHW805GhGiN3G25GJ5+Ko0VZ+U3fxFA8bYGtCGZzr7fYHeIiG9od
CbIN2c+u/NtKY6vMDGiretDTlOE3RXrJ3xrZLUjKJzX13sgtX1Q4nMjbOStUVM2Z
2+LLzG1omCEDViNWeO9k/4Xgz8dSZhneE2EEVxQZCRyRlH02zxa+TaF3JkAfAbt5
HX8iWSYfK5OBsLVyRGwnrknEuZFmHKmPnSlBEnWX1/QZOUuxPzXT21er6vKyTWdZ
Z5c79d6LVCRafwLKz0JnNlZgttaVNPNUShFJL7QcjOueJrIMks5Ab2c/j8fC2gdN
h5CkSLjh0OGZ8KrhMnmnT92pyxAB6ztVLpCP3hXz74LYwQCCFYsRPXe3ka92ELN8
26lcCo6Ldse2OelqGIiKu9n49MhYpaiNCFVM67GJu7nyOzHjSItdk0nfuRv5nvWz
JnpVpu9KF43QoWXh0PVEX2mcr67q18Rysj9Ku7joRGBVZeB7BkXw9h0THpk01NX2
t0UqGJOk/wGfOJ0vOfMxlQHw+PZMXNn6XkQ5II7uaFW6dUWoUOzjpGJ711Ptx0S/
fbt2Zc9uvjA17Nsd16esw1jT40uhl2HmTD7G3lsuD12iQ98DmJMaRnyOBi0PN77L
pThmjpGl6eXPFYIbxG37QUC/Lree19/XEhJCQW2bwMEkUTabOMNSXCQrRN2PkRs9
7oOtL4B9ZauNZkyNOVHK7wzjdDTsja8dY+MZlum91lA4nJQuoASveC4xZNRHBN3E
NdxZ/xwDc6wejc6h3VPFTjl+kZRyL/20VR7RV0f5yK2S2tRTDWL2O34ZTCJSeoM1
bER5pPnjeFaH2s6Wss42pVHEJp4EHtwCTp0THaaIQZ/6CTbitT124GLLBlopZBRO
On77fHjjFoEHqy9+2BLUQpyFa8ShXWnKvWIYlLxGzfiZsMEEoWZT8kpQN/uwaJzu
HH/Hs112Q+wQUbZE4J1V3KtBIFyam0rch/a3TJxHje2w/vUP+8lXfMjDw4877jME
angCbU9CKbNSZFHaMUmMJt1YAKRadHMSDkoCkk835KxHoAYivmL/itzk3QNwqRUN
oNC04INxQxnoNzKxcSeqacX3xOz6e2fw7Tg8WGdB+sqxCLelLTJkrF1+3rO0cEP3
0rvcF0VvFuNa+xwj4LEqkuUUjCQ9nYFx8d1vKLJv0hcKXiGmuhcyWMnAHEpr3D5T
q0R39n39Zl+69rH/1pODA4fXyrqKxu+4s/YBqfI1Y1DBx+LjU+ZC7j+G67945AuN
1GNYxXIR1WduLAMA3BR7gDvBkkuJm281WY/7ENnpbs7zOWlM/Zh1g7yOGjXgL1e1
K9wTJ2cFoWQhi/wCSBfiOhzXMLokAWjqSjUN2FkSMbLuIjpXaZO0Y4VfR4BAox8N
o2OqKbKKJuj/tekn0qIUYrx9RUXAUhNh5r5Zv42H9DxzmQ1NB/tIXuXVfJeb/ir0
GID7993ZyNbKqCJpF7Sw/qET2e9T6VoNPEcZ7HZMe5PzNlzztT3cYgEV7YKQLqc6
Tgmhga7rKTiRAg+mnUUhL/qlksDXK0iSZMyjgNu0w+y06Q9DmA10hn5JkJvHe+NQ
/IIVaxLJ7L2g65uML1jOeE9umJ/n2u3ViDI1hwhvmk2L+NW8BZQxZOQg+ho44EnO
CVNzbLciFQCm9yjAiJbo7wcYx+GOAJCRuM+IJOVI9tMrwCYKs32b6ZowO4CEgOmr
+yLZ+lD+VKz0sDmPuG9XmIbqa4S9Rs9iZ5m1805oNJRw8EWdRRB/6njyXJoFNJYB
0xnq4lslHlWoZgcAy5whKnJoMRwyqvyUWXvulELML883x03x4C1Wx3y4nzrAOvYb
jfT+GyoU9Ggj0vZJJKlEuG/ci8koggbh/KfpAEsRcxamnpo1sC3bfzyJxjdFWfpa
lZEie0loFLRgDRW02WaseXPkoN6Ku4cMf2hWEqwhzikU7quIwbQIW/uiMEVfKhMe
X3ptyfxtguPrVjjdceKOhUxx6bzo88ina/GMrTaNEkZ8s8Axo93+RBj8K1vnSEYk
9iwEfYOHYGb1velwFJKZcLnuM7rXWz0u8jOfYf5kEFa6DfDnQBruPfC7TZZ6s/+r
3Rr7hnXS1uvGVCBqfTOh/lsa9InoH4xH/LKgVB5lk0P0BpeFLyS8fczLDcOMP3Ko
whd4pGvdtNkbgdQ2RwdqJyfMY+JC7PriChzdDA/9umEDaDX6Ff/WuMYHkynVcdfq
KF6ESsPCR8IyerCE4j2VwVoGIiHe5eMs5PYFgE8S/P+dgHqI9762iLPcoi7qWOqp
SAqDadcnV4zPKTMHIPyFiHGjSmiZnNImbwTy93oPE/TlYxFtazvy2uXdot3BqXeR
lCFWDSJwaXmDGGaVz03ELcjfTE9zlR7fup602KFF4KUpJ6QVzWprKDfyEUAhgo0A
I+620k/dV8qlNKSSr2RhRJ70oCDZkOT4TIeXnjbt0i19+GMBDp7fPa5vrtyF+CIn
iIOrR3AQjzxXl7B89icWFHRVH30qaJzUHesrLQKqVF6+iI2tihBvuB/2BAq5jwo+
cjRZ653XPR13ysPLcgiV2Hi46uSaPxK0pDJhgvdbLpPL3rUsAZ6X5Q1wnHLsTSOV
C6pG6FKDx5ABTxCQ7dANrEaSCL+4tvnq7Ze9RBxC9+bvYcKEOrk7HF92/UGE904p
h628Ruu4Sr+Nfpf+ofqNaNMgkDHUC/sKazJINrmQaxBcXTK/7jpFEjOReggM3KJ0
l0nwhCadO1GOVPr+hmZsjscCGmiV8JUPTIG1AiDBtSex6NBXfnRIDjS6r81unfpt
HKQyqT7AsORfsSUWbbO5ZKFYj3j9e0s88wOVYFmQELx+01DlDE7qluBO+EYDuFxF
620VlBH/wCVLGMYXi+8ulgbABf5bfhJyoTQXAKGL8fbLMvFBw8vTNIbuAdq71oaZ
23I0kel9a3J20PfhCAonp5uV/JBtNPMpjszlo2Fd23ktUuPat1i1KYBRIHYHpCGG
kSKdY/UMCEq+2y+oW3W1JzGi+gyv2ZEtjhNs8dgkuvN36gQ/OaumTNdV1I9LJG5W
vThKZZp46G+omHjS4UeOBAJw1mMdNnYDWOL5a6u0bHLhcRpHUc0VBAmL73ytz1Na
d9RVLV8DFs9KaxPy9m5hxYJt1COT5xQsuwPJz3Ws1HnYhMhAzk9tcfYi7hu3xdZc
DGHyBePUpIZv1MGtoGjGPictL8dHTa96xwT3RN36m1yPM8qSfZJeQlGtxAxOLmiq
j8CscZ0zgN5EvlYM92NnVA72dbKa5vqo188+v436lcdl3h8eOE8vLjxxHlF3O/mv
WpWOJzFMubFr77MYPRjk9WORCstS7PAbe7w+zE/c8sF7FzGYgtWpaLByzAC8wcz/
Rl2w/tZrAyvqbvg6T5FFaJEp0ZPaChn7bBPXyT7i9tCqG1hdo/PnHW7VCXKwJNWm
DP1Th15Bqn1ZNAADvvVoKPZX/hTv5YZPmaXt9mYNe9HN7Fm4FHssUj6gbewUnPqr
nnJTjSjFpSc+JHI1vjyC6gpgqxHwqoTWW/7A5wx/o4itptIQrzDMWkfzQ3w0PVqI
rUQ/ac/xoCK/He9R9TRIx4kwQ4ZWDWE4jegl2AquCK+bOuaEPhMe7d2iR2RnRGtr
cxtCXpVuGRe/g5/VwTKx1biyFX9FtzjRmD85+Rb6lCiPQteW8PWJIPX3JPz1JXGW
iiu+KT5k78KDmb5vbgr0SVnLpOWBS157UhXuImdJpxg2nPaJVlq3zbWfrLQDLJ6j
qb017Agi7s8CVyFyLNPGtjMJ65Bre2K33qDdnbA5szncwPHqx6hmM3qz0F2ermDb
95pyUPSWmCZmXcnS8h8ZToPurFtpnPUgFzs421+jdSENx+dX8HmkPJOHuZ56dPQ3
F2t8nGPphPB94Geas/3JJfJF4TjU5lKEgDTA3aHVqgCADwX/qqVb3KokiFks1uNF
NDtiBTrF/quqtMN7+ZreX+mM0YM6aqyjgAAUl3lwuHujCKBT7oBtwNlv9wnISvc6
CXS7NJMrtqWlbGee3fCmTOGzNQ5wAvKY2tq+AwjKyBOF7Ipq7P9hw80chCwLUuAP
ROsMh0Q31DffWs+8uptBQ4Xo10oWMsW1R25RlUDBtNKzz9zevuKwI6sFy6ZwHdXP
PX2RxwNzqDKjPQ6dSc79yfdemj7Zyat6BiUFC/IrZmQZoJPio0av8hcQRs4AgFa3
2tlmImZPkUeTlXmw1xKjmQvWtZmuYje9I7gxuynzEgGftwChkU0X9/Q+GMX2frJ7
zitFQ22wrALRu7TN97Lw7Ff/a0VkzXj+rWbq0X/o/ik+vS2crwJIJ15zzRy+d9rM
TdUXIGsj3tID0DnO7YuFqkoAEGjkh/xKydU8P6VU3IRAPJ+6GU0H5r97PHuSrFcw
2BOQRtAA9Kxb0FwF+ICDzsEyFEFnmpCnThFYDunG9Mj2ylSvXMDBvXIwpJg0BAZH
UtL5E7ylCNiuq6zzQ9/OaQMAbRMjXNI7xIH4kaOXD02Hioamg5rPxnZ5fsamSzyl
SPuCpKJpUncQBePYriRtay94hXQUMpI+9GL3rV2Mf42SfM3q0L5kPSrq4D49MA3n
uOi/YIChRw5bSiKj1/0F00vWigPoi4x3oGBLjLJz+l/itTdxcvXvC4vbZML1iwrC
Wt+PKgUpUnxmaR6+cLvQYVgaYYBEBlDppUe+wN4dhMjv9aVAns8jz5gYTYg4V9Hg
e9C7huNyoGq+wKvABdfyaPawZzd3eLArCFRvbyo4+KrLeyaCMBE2WCgFqvqd3A3g
BG5swGA4ThXCCGtMT+QaDfXj/gV91hg+nUAGZpN3A+3ZYecnZubT5L7j+n0zYBko
pxTrohYVHNT+urpsaH9He8pLCmI3adtmFH8BUTqrzFgvINSUMsBjSFaxuh0xcbQR
G7lDn74aCkaWeO/NKILkCoHBsbYJi/FiFAHavsBWLMqPZoupuACjY0Qtj5BCdErt
ZctMWrTy2oZjKsdvDEDR3lDf5HYEX/JvC4I9dAAQMot++UOkib/ArplQ/4aUnXhY
N4qdCy6wtQHWEyPFS2p8ZDQ4gPyzexX/pXlIwoiZ7xt4ASWC4+KemZEvljBGeMnT
+iMe4ZiBlmYyWO/OrQwlRLSd/CCyCbqwNvGwyI3jhqClG9WqgKTbOWz3/2Bpy//I
A/TE5nJJY0SIihjTPZTCAlnnnmiEtA51ZA8fq/QmV8YoBOhTkwCoBDJymk0s7ndA
yh1G8FN04RI4tv9P7+Yhdex0T+0t/m2vXpPAuiXzJlTvyR8ZEYf8apU05L4koTxG
P5oA/zUJmVv/ERwXk3cfteQbsFqwLRlBgJHJGW0WXPRSbjDuZ1Z5i0XerXH7bPe+
s22UVpPCPwkwTHwDIomS5klBHEUwnXodj1aSXsyWwWKpmqCEZO5/RsCWxOm8Qmui
y2QESeM897mtoghY528wrlSM7D/0ifDBjyvhZGA+fcchI5yUPuhvmtuz4CHpH7Fj
EKJUl5IzI0jHjw13mUWj6/t+Z+eBDcVJoj5/0rStFjaISxHS1YROxSO1/AOu972c
Ga5idjvB5pYMmF6TOQ4O7/HNyoEKAKygZk60ROlIimq6OgwmgFx1W9nbXa625R60
rW2jToMW7T0KYdQ8U9wH+kdnihZuH8DuTnU3Cn8tib3fHyQrl9r3WZYlABAHHoYC
GmJwIFPC5skqBrGcb1EocVogZLZYq9BXP0pW3Q4Eit6ypoW0FPflBu6YjE80aJqT
HvViyibx4pJMx8o25mOELvL4w5MirIDwwE6FZA4Uyy9praiVW77TwUmVBLYGH1q5
dQ2isyrWl6v5X3AV0ZtZ/iCih/Wl5Myy0wvX4M6AHcrKhwxMDYrp3kEgoqSpcNI5
w0PzXRsbLsaZORyK9y6AvE5gwE4wy+ujqoAfDkFNwbo9eHjtt/q5rWhnjGc1txWr
hV+47HsXmggW439gdODe/JO/Y9KLqvMP9EuASCkL484FdZ30RO1DBU7TIPoOZ+hP
rCFUZVqMQ5WG+wym8Ppnm4QB4O1Qzj4u/yzC8ytFBiMP+YnUFL7v4CLU4V9V5z78
xuwDpD/40/K6sXXMD9y/J8M5jzrbRBGuMoeGkf1akD1QJYgjDlN0dLCA0xLha6L/
DmoDM/qI1XohiYsmCfpxTUTp4k8E0G6eC1dr2lN0lJebY5AKBy8FpcIP5UgPLUJU
zT+rtv6WcKp3fELK8SG5R43kRH2CZlif9/+1IXWaeVlx40MoHaq7VFpb4Njtmda6
f1deXZn0QZhvPo8zT91zqmP6yiylLr03sQc5Z1YJpnjoquNlmIkC6eHFNV8ejvpN
QHaMvRoVG3u1Vcm4J68A2JlcKUhwbJLkLQ81UJ3YOsF0QbMEu6UUebMjUnoNhZwS
ettWMYYN9TJi8NVd0ILTy3jBuZbSYy8V4SKRSdad+ehmDm1K8BWRbbPL2n4qUFR4
ztnIab6owAwMEGPRv/j+hzrifOqb/gfTtJeB/B20SCwEWGV3eaUm5e33ddpUvxE1
pCg2HR+qgqIgN+mIArYSepC8YUzi6TgxI897PIUd/GtC/ZaCqNzyrdnDdQ0eSffL
KjKUGzvKwjXLv6vmBCSNxPAJtIFs6Y05W7L9ITMlLv3UwGpJEVK36YHs+9XQyHUC
oIMPBPDfHbbTzseEkMHW2Nc/vfxIEI5/k+FqpeZqnyikDo8N3eSd+2uavNKi9aBz
WmJhiWhXNEh2mHtVyfAbQXov2PX82qTctoShcbubFJM9sigmUQSOM723CD9AvBqM
zp5122LWbW7AVi4VxIum79f/zckI5ZymXWwoLtdz0ACdgXAzhJFjhRIInksgV8A1
m824BkzHjxIzrw1+2KPdtmqVFKtT8atrEYYp1u0zteiMKIVIP2aWvbrU/Kn4mWOJ
b7c87caaqApAQ8lULAMcqYKGQinf9qyJhei1vVmje5hvnA08Wo9PjGd7FfPyRUYW
BxYJu4xaHg+5amXjvlt9OngmsRUXQoKq3Ih0WjbUP4zZ/i76dPLxEHLdpkaUiXmJ
hDF0auaiWfTZwrpWeWxbMhx4lxtD/l9phL42EvlFMr2f1txMzvpm3k3p0CTUL7T9
tFNh5+3rpFW/lJ5XbJmQeQ78hs9kZsY+cN1+GGx63P5t+vzpPk/gUBRmRGNgYvLw
1JscMBAGK2ZnfUPBGbC8Ax3eRKtz19lx9wjiQoOjRB5WAfhoRZIfj0rxz87C5ifw
Eux7Y0ra1VC+IR2k0rjGC6XW++hV8vyDLAetuP/9rpadYNEKfveqtguc7RBanAQ5
YcksEcrDXNs+8rYJSZdlwfu0K8S9QTifUZQxF3lnuwzCyO/pzH4ysLuQDesOiONY
no+7hTzOW5SdFG5aqdnZXutf/gPrHle/2d1wrCR48eoQqGTCDUksJJXOfXphAwyH
xriKRsYg87WsDhPIZOqJORoZpCM5QjmjWCdh+DhTyDCEfJTddILdgFb+V4r01CTq
+ZkFSBAN4uRdF+lKwU9G2nONxUd17wWo/43hvP4wbSboSt01WZ2uLFWdeJsk8nDe
RBOTkD0eH96f2vhPtP2UXtWBQ0OyF8fAMANyOBUVw8HzFFiNJbz8TsQuUwf6AA5r
2dsdSExGWunWkSjHOvs69l7eNKjw2AZyFYJN4Cms9qgVsjigoDScc9KIkO/nkTes
u+mkdGjl3csKoWQPbwXBIEHCVLCML3k49Uh8KduPrdT3pS7kfYyuJnWBsLuiJeC6
qLTDWKuoqyg0VtqmO9j8/VMHjdk9+Y76ByPyreQ3QdcaSBF7IAsMzVkFsW0zJJiM
LwboYBrdAWtEam27+GCE4BCmZ5DJ1/gKRv98c2jhetWVR8J6xXKcyWZfQfImvl+L
9vdhUqZ4YlciLQ73T8uqOLDahSGD2LnA6xb6KuOOlN2iB+IFbUdCKxbccVjYH9hx
Zo138bHuyrUX13U4E+k4WN1tgpVv6sjs4VEVk2QnQMZGUsYQ4lz2oh5qHiQ99G3F
TK5rU2CKwhY/iAHfzTKzqZPkvdfKrr1PSW89ky/8qXMtQREN80rN6S+y2Js8gNWL
Oe5xene876L9PiEJwsDVmgv4ISO7KyqGS5BNSq1/zZqOvoThIujLRmhiLWTLNNQ9
NvWs5JQQtBeG4FPEyKZcLjZCX5mYEapQKWG38Od3EjBUggmYEkv4XTcOUhubL8xa
JJN6SwDkGa832UqKidjCcm6c0yPcW+pFLqlKBC8FRvK3BMwtYYmN4lCfhEtukCI3
cmfyBTuswNPX/yp0vSWA6tU4XuESG6MwWWhH7g0LYex9MOSjXe3yomd7jl9VJzi3
EF9Cz4Ehka2AaOF+gDfMpmA4Q7Lbpnq5C/FMBLgQBaMqpGD8UteJX7WzfpClhJrf
QvLUSpce2oLPWZWns8NacyiueRwho+i61u6Oi3zQBSXFALXBVgnN+oDme+fckB7+
1nKf/nw7MYJgAlIQU6zNaoqhFBo4nF2ysnMEfGufNoouR3DhYFBVFWB3fPDV5jb/
cFjpWqol444JeNCr25i3s7nIn919FiF5Y/ZkXgzP92MbVR9DaB3b/eQjLD4Y+X+C
J3ou+Kz40Ef1DqQDAdOF0GLDQljt1fWZ2bf105VsRD8NXwmn8Ftz1cyWrUS9/cff
hpBkfcPjJjZLPnyVbKJWZAyP0+HNctsYUiaKG8PwBT+1drIMLNqxvUT/KLZtDk2C
Wj76smR7nOOrVe22EyIwxMM7bKWDaFDCY/eKVVFxHDv4lXSQMm8sFc0ECWqBKYj8
Y0Fr6LFLPa7hDit5jNFqDPXsu/Wwbou13Q0q1bCZlgeZcpxHiO6CPv6F0qXTX1T1
FtgIEz5Yi56e6kptnKdNrcmoEQpibDBoSzzwGfLSCCFxZ9jzGa4tKf7SarpZOKVr
8rZzKMES5P12qzTc4nx02TmfvuGEJBwGjZetYag0X+4HbNaofxFCM3eFATtVBZIl
gjwWcDBKYncetLL71ZuYlkhGp2qz/HylsCeNP+jFnq1DJVajskVIx/Z2CIbdC95h
kf9k5kRaKMg58Lj02iurMS6q/mdRjdeE0JwkN22yActBPGtelxj2fF+Ceqg+rxfi
HOKv9XrlNIDrsrneeoP9a17tnoDGvRdso9nt+fHzJA9bji44IuRqinj9bb2IbGSb
dLQ3DCwgPd5yqdo1tilRlbtBn4OGAz+Rxo206akWsygyuNrRB55tu0NP8/CmgGjv
CmqoTMtzbTJ01rUyIBmM63ZA/n8U+Px/ihlrlktbE18aTKTvR43uE6O/WJwYvDCh
BD4ro9yh1lQGM4OE2krb6C8/Iqz7bTsaGaLDoB/RoL+yi89dgW2lgeVoDHMAxBDu
Jr3uZU5gpKvO4JuOShPt++Fphz+19fFCXaTsNd42qvK47cXePi0wKQuLoj6hIsl0
yAPVvttVO5IifkXZnhGMHGzypvnQ0q35kqFq8Gr+Vj+CvOYqrQCh6USKbjAUOSsv
iCwZ7EJSFDBxm746pbhhy39mij2Naw6m/5zLN0DPXoqfl9WwstuKpKYhfu0UBwGv
0/y6e9gXjhGKsq4tOA0Ajb+cEJL1fnrB6eP/bBI8FPDomT0nZ0zrQuGEM/H1qv2I
ydCZimXFEfDGpM2ftjvloN4i+m5BOXuACOMMx4tmLxZhZ7xY1bLAB9RQXVbh1LzD
AQlNWRY3CkS6iPF3IaVsCwEpM+MGHEtrrBaziCjVTixVAEGkSnzDpP8CKJ1/iO+G
MtT/maHmBztaBA3LR1jj06TXA+2oh+IznheJmDQrvYQFNnNXosDPoD74gbBAvP5p
hc5xcxG5GOayTniMWb+kK5WwpcVKEjFXJEJRcrNUlDf1NiHbjSq6Mo+P1fVlx7gq
c/EPy/31LjK5Osoi0a/TnmsbPP94X9a9BnjRbSQpKKBlgkwR0dTjTlCCrVw0Tl3b
pyRfUwyQlA5HpL644HhQs4Hwpg4odEKd6OPcelGBAPql/AQVP5JV0HPUQFisWEQN
CsD5qt30zsLDscsMOu80mFgwgMTOURWGxUV+Z/rqKpmI8UjhbpvHODgVOLEiBZmA
fzaRnobUjfSDx61o1IOnFqPT0I2v61qyiUL+7nWjqUPrIQiSCq1sRv4iPOqf/5BN
xs0hsOcrQ2x6Do8UN0+r9QXTbZ3vsX4fMPad2xwrvkE4M+ETMbVrRQHCQlfCGKFM
wcma6LGj3NzteU021QT90prOI93OBF34iNJdGaJoi+HYkVZJLY/oa8FXu5wUCPXv
1GBcV5uv1U2qw1iAzkRWOo2w3JV8Mbjzyed9TrXH9fBxX+mKfPNGAXbO3euqnKE5
xpD5DwDFC2D8YqY+cQVks8FBZRLxnz68oOp7z5VAPtIzqn09EPrCyk4vVYBzpEnL
BRJOluhEhJhb6tKnB2KrbihxiwV/x1ZmpJQzfAkKHCj5CBtqFV48xOdH8OkhtyaW
mRePXT/mH9KW2L1Nb9UKaZ7QWBTXJ5yCib5ZtD5E3N0qh3YtIajuBJrRAO8Io8uY
XpxuwL76YzXW82OAuOQUNcAdSMqCr8F4xJvtth5h0qeiYQYinuRfDkp+5ty5nSDr
BeygNRlUxJiHwAd+yxkgH0zM7gwL3ARhT17Zun3kjgLsDHp83Ed8sDpbQDOjTXxv
t+lNQAoRvXkTXDORUfTk+xm7fN4OwRvz101s3Aa2feYD9iKQJnFdWc7cGx9dWLtL
ZQDkQuvDTGI8zAjRRZm2k5XQt+tjm8xoXcVUt8XklQIyDZyFGuPCucAUUBL0TYp3
Yiz2XW/JFMA2MxyjybpE7cKa93/952+ertzXLOq0hkDAPAPCluM/lGm+4uf400j7
fwfUqK3GPiRSCoPXVLB1qn0q3eBF25qZFcdl6JXV12mpzg9Q9+n2b1ZVrgoWMDF2
jw+1a0DZkPjDeIRMZwXkiim5S0iDphqjncFelIRXuC71yeq10rDNqKbdjwXa79Kd
VH32mTZud24eFInrrHty/eCNXMltJf3CPhoW4cFLMRC+KTqkwFp1cBlxPahG/wrx
KFMoiJ41MTCS69WnZ6VqXl4ZYLxkBv3dd6iZcdDhwttcNdTpv2euK+deBPeW4g4q
vGRllyJKZaLqVPycYDIqDvi9+LgRBs3rZzqGdYrI7Klc0fNi241H/Fpl91TabntB
o2QjWhq1wxfykQ4qgqgZq/hO/3JUOS/Ek+eSpi8z5sQ+4PzATtDId8QtJL+6sZXH
F6gjN0qMljCcr3VaXHH9lNGWXru4HGOT0wKtH2xVg3qedniX3adjyISJBcBV7w6g
ojF/R8NMlBeG7lrc+Zp+kkk5IL6aVIHpL/LXyimFlTzyRmIrnMuflKWrDH5THIO6
0Eb1nn0wW//Ma+12zN9yCbLqQS/KWMOz9VkeiJltBrqQaV1bHNbxjvq/GUeQBdqL
aeI9inYO0D4uQvlfYKl2mAuAKqMS3F/Q6sxYyzQSkWZan2DS+SL0M+OQPd1onghq
P5PC4ZHiewsq45X2I0dQFZyAxb0G41dgf2YMh0T6wN890wp6i/x6MPaZy1GapSTp
p7191rq2rKZVmCOo9cJbMcmVPTzCjZTmPIV/vH29WMaG9+aGCF9pdagA6owvsbuh
kcY9fsO7pP/sJ9mlP1pl63EVpYasOExdqVzpb2+LM07nHMBIqGeBoXrKuSf47oO9
l3YaxOOf/VdeUm2UOaNadsXDD6hKXExdeS8FfPLc1qOQDnVaqXHQfuNe4kHSiJla
E5dom2t+3JF0f2I8k3ZOFhpJ7yZm7G9hGXhOvaukl7uQfnHojzt/OlJsaGjwuXwY
JJx/KlvdJw6flYzpFaj67lJZajl4AoSV7hJvuJCFbk2linC370AoK9UCbkuGzZXf
spMCABnmDh30WDMjWeQEl1ZYFdgH349z9Kamd93ivMQtNRfZgFGtYJTbfNdBFwNi
Q/DsvPrnlCCEpjXJGnF5pQUGmv58wLIZsEvoZ0UZ5NDhAn+uftwX19ZhBG9YoRWF
G66kMLAqmIed2y0TRgHyo3HayuKWFUKgIqDJrZ7p8SAZJTsd+PFlDKfzGevioYst
3MariAaesyT/Cf8uCKJUSwfzOH2BtOnM2wHUZlNFkmlMw/bWjxEF8JhJGHLgpJ84
UyRDtQIInViVvyNQYUw5r4T4WjGxmVXONrAv7uq+pOBJz492VS793uNXTv4HPObv
G8DT/1PjQwx2A3Yv+j9Chwm6UpuUU6OUWKbyTcXulDF2WOUv+dpfvWPGdLqTqflI
CkhqNYvefnAkjlhwB6LBT7ytCkqLow2MSjgXlFHYAxOy7XiQGCxFCjCnoEcIMl3i
vNLVd1FMj4NZeJg7ViDlcjxvoEr6Mj18aMlqVJGGmiIPQA1T56jEo/8nVwE7kIbl
3/ieRCX13sSz5RFPuRVWiTrmwS6I3O6WntyFf4igsOxN2G/+TctbvRqnbkCrDWDn
iA2T2fMzCWtQ/jOi7+CPdvhIxP1fIZICabOzmfXDuvToxFqdAnOjO6SIG6HcGab3
2jL65gqwsWJl6FCU2/yoUuPH7om5OHwiyscynvx5yIQximCz/TlW8PDSBlQCTpt1
bjV5ZioOaklEkXN8sOZ0BDExTD+/yN0Y1DDuXFkwOJ8psoOezC4JlMwT5WfJ3F01
RZnw4JBsonu0zQXofqqkNqtBnzcGwjZwc5ogmsNp/BRTZqnBDqpoulPZs91u2cEN
pq/LwPRnzwdGtMk+2v0LcSpSLrOrm+yBl+Wuk6mEgRHJPQRiRGq/u876btoJk8O0
2YQAttCdPVSBwUT/xXh1/wxVsnEw0CPyk6dWY9tuOZH1iKgBFy5Io4AKCQhENJw2
VtLLkJyzIHuLug1nuL52ObDT1ISW7bhP0Gxgknb0s44O9miAqR+3EWt3yyRKh65s
qIsUY7PZdAI+lCK+0s+RWTSWhPfTeWMZthOO7T/fjDFSWaC8L8Wl553coHHEJWEU
4Khz8MIoVcX+NSWLvwQY775xumgpm5PLQrkv0pM0nq/nJtX6FmZEBabm22MaM30A
Zw3byvNFqQqzdRQSVDRZboDDse59I0QBWvMMuTC5xP3AEm+ubaRjClZejdmAS1L/
1TtPOHOre24IcEB1RiUOnZpxoqjDbYeOGGYaS4X+lMa76yUQUSnCEUgp9K5bEiij
lGY/P7FFtVGvVIWqsM91lHjsMufGr9MnbNUSnGnz1ROFj60i4ZU2CY1fF74Hw4CZ
OjfMrZH2RFJM7wHXyT/79u4fRzHvFsZwSt5Ue2QVQu+TGDBDFUyx68yB853rmpOw
SCiSv4U+7mSy0VcACXB6J7udXKEFZNcqEbqKr79c2RLRrHsYty/r9WP/fVE/8gbH
PDWrngdFS9vgr3T2bl+QkKA2ueqXObmb7Xl905Rv6prSgya8VV2O09tiUvsqlDTz
zOKJ70VFa6d3dhvX8PvkBeQIV3Q3xHscffjS7rlmOcnCnck7nVqpGRYII81sj8IK
qZEFixT9vZEYm+Zy23sVXX4yjvoHZwZ+U+L2S+JEn4VDdS4qmbaou0N4jZsoa2ED
DAA6IpIWOTbL+C5pQQSqq+DISS+j9PxEKFCRURzkxi2Ib6ujU+RX1jPwPKF2ntSr
CC+moqNgmIw0DeYBS2hA78T6ZlFRVNHywqQChBEQsiqJbIiHOH5Xt2SEQl8g1pYv
xYt4GtbpDC1OJF1Phgdn+IIYMPQhKchHl02D8F4qLaXoFoT6trIguDgkTUZmgiBs
NXcIWPpjVg0FBnpK09e7jlYmlaEEjaOFItiE0FKduOQ3SOMGXk8Ayl3+0SS5M+H2
N5ehYSO6vqm2Bg2B12GgmC9tB+sEH8WynRtebRuLWbeua/GnPClvVCeuJ0rGPpYO
ot8hh1YsxFCB/E9z+KvwZk4YOwAGXoz0KZg90mbyzfI9nGRcAEEqm1ErV1vMCSiM
dbINsPx7zZXyP1S9k0NiOvyi/JNBR5L+rlEIKQL6c5PYENFdAOLFv7bhpTtcbNVa
GrI5VfdtsLWOpvDOCYUrt2G+SfGXeCBki9n9BRZfXXAK2kzHYaMebqlJVKDSALcy
C5+0RosOvY2U6HHYm/DjRNT/l20/YTtTfw6OGnHVoDmmlFbwE/wCj2gNLccbxOFE
1Nj96/JIXQ4X72HVwo+3cGNgRKPv9au913tuCFjvCZi8fjxENkBRvT8fJOSVKcE7
L17CoIddZ1hHeEaFbqdHtiafsrZX8h17ZkEdRWCPBgBvh1K8ovbsJH6oW1G/XzvO
2qHfUUlUiiz9Lguutoy9WE5xjIDYobXDH68lEt9zcYqPE9mzQCl+uVgNM9TQd1zk
4au/H/zPaiOX4N2xaYZ7CAfdJ4hDZ8Yi+3lWL/vtWtqPsAQWXVn5Qk+GsJLuHdIb
Hm828L5ZfzjTEsR+rautzj/LaBG9n1/eTn+fPcC0w+V2J+O76nvN+aBpFLOGi/WJ
lvvex7FIX83fp1du57HbbqXCgj88AwRat8k5BaNmMVZ8H63Msw1QIQfjfm88HLGd
gSB4P1Y6J61xon/G0jByf8fQZS/3/A/1Q5w3rp7SOBiLj6UbwyZenyvmLT1n1oR2
1DJvB676ndz0+7EjJqR6scSDtLb4YsZDGZwg3Cgt/KUpUWqmyzd1mGdX1SkNB6d9
wm05ZBRoNaDE3EJVwIZ9ZA6Heh+Zs/S2A0uwcbD3I6Z8XIoLMaWKWx18jOoqQj8a
4P05pav16n16Sa2khZB8akLO8jvMU4rvutf2OiVyfECbbKqrejCURFfBosB/y8JZ
akh4zMMUngPYlDzcQk/LT3kTz+gGY0VeV3seBX1jhb8IESLSha8ACaZRZljPa/tW
Z2JhBtuAA4N8mTYWfELi5/8QRTMOcZlINnboRqw+zN1yqS7+z+34XUqHiNaP/4gq
j7OvHja6A/ltSkrL4V926XW/XgldZz5LhdzbVyl1xk1qRij9me3a54/jy9Mc5Jm5
FD9LDFKHRsa34Fd+Va0VANsfsnnfg4G6V0aMz9Fi5fGU36T2okypKO9e46vRKa3j
9pyc5ojkGfufp+3jDoiykcJRstabcPogQP3H30CVQn1DZfRf/QsQPzoCHGaBl/Hr
358KoKgwrdLYYgYi8aZXI3hGcd4g4JkeYhpg2BiOlcuZelu4a+peSXufa25eP0Z8
aJRyXs0DX5ZtmksSXBafI4XI5EmBpwgnoBM27k/jB24EPMyU1Eaxy8LuOHzS9jtJ
/2kAIKcL1Eahs0R8ty/k4ohtDIQLuY9/0a9HNf0jZ73UilMvUHKJdkfrHRTLePl2
7kXiS/ezEnf9usge5upbWfYINB+t33iDQJ3SK3AzxmwqH+vihViyEFSavHmH71JF
/L6KykiAaDghTgOiDdjl4vlZGeM84m/HKC6dRapugsazPrLmZQJSuq7f8LD3Hxem
bSCLyO/cIOZ+p4/bXsq6JmyHsczd5Y62R97LRS3O6H8kNvpSs1X9FHSK/HiLL1Zx
b3xbP99Zwc6W5yIEeFilw2a9bpDpB5TmWTQrvqm0E9uoHIOXxQQLyMw0E9rkMlKW
awWb1BY+RMr7V8SDbhA9LRw1CIAv0SstEyLleV4+qzJWcDoiVQgEINnQbuTOpDgE
GwOUAvOAWHKJj/fNZZkA6lwX6qr77dhAJjcf+gEeWq6cTWsDo5V/IKUjHTLL1Coe
AxBdhPzOvuWIzbUzVHCGgYgEw6/Wj3rJEwRlX5U/hhqmu/1AhwF6Ux7F2zFizojw
WmEXxoTu/JmocmBLXi2QgymAFx1HJnEf6VogfhOZ/k74/iV3X0RsO3KWRc1lQ5Cx
5Fz6SFN7nHUQ9pkXqlCo/X2KWlO7i/h0RLZByLDVtMfVEMB5OBRFF2JHgNDjOjWr
HFfQweV4RYxVp8UPmlGmnQyMBl8yM6QTW1AxI5twxvlkHoidLPN217yCpm6zgMK+
EcswhOeeVFCRM+0MxO6rmxAYSfYyn6DXBIMkH/kU99CApfl8/rZAoUs8RqC7tGmX
DfsWE0BvkraLCHr+Cw6Y8zRMsqgioRQX2vxG/HUjpf2fj2Cecr9PCukBKDxN+wvb
5ghDY6poeBgTFb5iL728uzAihXAiIh8lKKaoity2g6X5bTqj5ocWFrYwoDMqgjNT
QWrFKk6lAY2hqbzRWM9cQ5k9Y4OpeZBn0Av5Is7srFnf0dCW2qhfoOl8J7z9I/yD
lyBcN9QJL1FA9WaWIldV7UwKDcfCnKm9Z3/rzU6rLtqvX1EEd3c3/7ar/gV2YZ4a
HYDhXB5/G6JkoD2qoObF2VhafgaMnsqNImtVTp06pnmPeGtl5bJJi9Kz5aeMH7Pp
+PK4YubmgNByJu1s+vwHOm7zSOVIal9VYi8CzvF5EBalxHC6EBv4QcOHOciQOSgZ
neWETP4rur+IBiRKjb7OEid/7SMIOM4YRQKPvIUw10j+kF3kd5eAOJlkn9xtkJNz
T5l7TJtAiFHmZhqSvpsXfpLdUAxjhvAY39F5LVbhHFVZexIiyKahNc3+qjikjBgw
CjjlLcvgr0cHBNJbU6GwjJoPLC716a4eiRQDN+Q2QjxHqn+8VqPe86HNY9N/Mht9
wwTEytDL2sWYuN7fJ39VOxSHxpwliIuwM1Sw8HzODfBI5LGyomdYQEzAEc7nAtk/
kkv/Ncaie2ok8pp7LTP2G78MfVGheTZ5QVZXWvdA7bidxWVAGokTgDEL5BIzTe83
5CQKpzLZAmfnnkRRe0cDBEFGdqiJDEmibEFY1Nf8XgUPYUB8wRbP5FztPARWdWM2
2AHtr9zHbcCJpIHJaoyTS87WFgMi05xnN6tzK8vwn8ee5xSt1jS+SOyoviw45myS
iNU2Uk2vXSmV6pwiCI8MdLYk7JObBxtaAi70wn7SPZKWf+gaNjqPQBaF1iORoTcG
PWY6tACzOBKNnZ2isIDRP4wqa9rgVOf91GyyCznVUk0r0O3YbwZN8jxo7ousHBes
ubErKbfjC8QTBLLLLS0S2i7saZvQ8QX5/n90BdbQZvAGUichjlRjYaCx0dnbhGVP
1iwcRn10e+ZYj+tOvDtTjJ7/6KW9zPCptpagjXoz31u7g/E+ykoQ2Ni48mmcVBxH
oa7v2/qtu6fL2KtGfpwrtoP/fn5y5Nih+Gf0n3gbeVwJxlg9AXWiILjKjJ8VakYx
QeGAW3YJ/RbcsKeQpy57Jf9hE4l04WRuYZijKJ5Z3kVW2sC63DUa3dy1RpH1KM88
MY9+sngl+1Qt7ApN2ym0WUb4Z6lqxBmO0IlUcsqckpBbvqbUvbuiiA/hGKuIAdFb
nP46VV0jP8yZjqts+6sw1SvXwR8qnI8L8oCAyTlQgSrA4PXDgafYYSCfyp5ar4No
pbPz3iJczrBkEAEyQmAwtJ/O2Bvydqyd3Y5uu5zIcxvXXlBKUlD7T38cwj1ZGNY/
xOm16wkVFiGWhcdPIiICvLuTN9T6jXa5cTEnbvQnjJbTI0qc4R5mN6uOO7a/Es3q
H0PwfBsnudK/ynn5r9EBAzR5RfP9M4M4M9ZfnKxjRyfIeqVpdW1tb0e9CCKuFgbm
6gSpDvHvXgwq6ApPQgiKXr/DtwLqffX6KfVOzzjfUUxQezZsP/S0fuKQ2bVMbskg
etnDpA1FaK/Qu4/aJ7Uuq51z0Bs7GPpsMHZXBfxiw3vC3js0YrdCPAErrLQRyNBq
m/rsVA64MKQPdudzLR1l8CCk3M7MD2h6U5W4wiir+FB9qIY7j3csRrUlMNNeM+cK
v2T2PRqHCTithH1OHt7c1Z3p+luHJLtD64bdyw42kgW+Rcku1GCfeUAP6SXgoPY6
JbyuNrf0feS8wVglqYEXd+JJFetc2pE+ZRoM9LiHkHibLSQRA3K7z7AjuCUDHXQT
X3oyxIPUPGNUCdhDAki6h+ePxMPUPjmemk0ies2HlDq2xDm820aFtPYvZEBr5lLT
PLnw6FMctKTK2FjiRfxx0P28gLyXXLiPZB61CXlBu+Qt0Kho5P7N8u2CusWrJrPL
kyj6ncNrAx8fc41iE5J9gAdjvXDLYYde1kfES1nziRW6Y/VhoRt7NgPtAOuVKGWj
WhDFl3Mcha+WRq4u4//BIg0yAXVuuHPADpJAT0OXqpTAB4uByQmhfx9IeeLIHp4B
tywoUgYOk4fguSAaJL5XYuPByPC/YJ8DzFp9cV/w6p8GaKj0TT+mWTyGp1BFZ5TZ
ZQX/IflI4kd5GgrY7PPcFS2+54lbuTovNnFT4AHV7u48CyBu6Jvr7Mwca7ne6LYB
rtioydv/OC9UXII9MVx3IHJv3XC/bCHqYK8OpLmrnq5NvWf1ib8xi9p4N0lEgevD
nnE0RLEQszKKlOcSqym4xEzzRBkzVRr8Rv9GQTTIfrLz04LdDOy64E1rkCgOARt7
J7QS3S49EOR76O1Oi8UstovGVHTKbbszFwygKJfhVO055It5vf/IY9h80sARKBvy
4eKOe2iGqcg1GkJd8t3yXx+lHoFVmJe936Bg65Btarxze62p8ZSaXCquQDpuo0uo
9Qy7LLyHP7HIM+3O1AwryT0YQ9HBPlINYytx1vWL/MsXHvK+jWvDy8YqERyaRoQN
+rhSgHqizYqQK9XT1EtEo/FspXkfIBA3Z8oPQyHeM6nvauXAh59idvaypjbx4bNB
cex4n4B+jBKfv1/Kpo2I2KAot9x6MMsXABtDgM/AGVtm971tA8zsHVXxTdY7pEbR
GN8EO5e90zWS6pKPbroqw9PrvaE9SquqAuIIk+NotqyKk5IioNpewzMltBXrC9dJ
b2elqpzoQ3fA1DcBJSla25lUVpJxmeYWQ9cQ+5gyfeI6TmtfMHecUJFAAZZhOKrQ
1UmciKwXI+I3vWzp35r5b174GzcOKJprhgMdQXWwjpr6eDIJMpWVEhklnNL85pCX
KOYyiOo2kfBAHhL/XlRDKL6sBYStK3FFNTkgngifTbH7b48FIhhOFG8HqaD3Lg0j
hamC432hfmiNyHfXx37ieY/sdr++8RQDavyYiZZiBi+SpXfrFfPH5w6FD2/BRkD7
s5dRZsb6SKXZyQpvB5js69E7eQwNPbGYxNEOygIad9joW9LECf1Vd8jX+8bwPIJh
tPdx11kwuyY0c5lXbOwTXu7FZ+0WSTtAir5VWIXFevLyS3exA+k1Qvv83spPcwqg
GU+TUAGmTCKNIzCzJmbe+mPMJQhJMWKfwvbWILz0rFwCrjGP0XbYj8vSWopjSLaX
bVx48GWNQcdd2K389qJcknLN8U8qzonhJh45aGsuuJVCKk3smkxNxZRZVMy2IQWD
L0hRX9h/5k0Xsr3PszOHRM1fJivmNf/X1/tY1NIJAYe+ER9b2QprgOwqiJ0KJphZ
lLCO3W8J8YdRKxENRShBhoaURyP5KxALsf42oWX4tAwZ+xqYSbpRjVNCYYkEUA5L
B3SAti4pl+k57hW8mZKLS0t8ufSSk1vtEVoqOWtrvmvmT5nZbSQUdhXPfFobdFNJ
GuRJdU7T2Q3LEF4U5r89z7Zoe+jaOkKP4AvHRpU1v11MbYZL5IxIRzPzP8W86wjD
VM0syqQb4NYzS6nTkwBkgcdHzcdGbD1py/176V6604vEP6iOpcCe61es0NUj1VAc
lrwSc1bJYy+kMjuVk+nKJMiNfIxz+wclX7MNSuh6grElPXOZwBnENwMXAgxpSD6B
Zp9/sx+96IIZniMydXkv8jDvTnIkTFiVNpDEp9PkaxmsPb9r5qCac9vwnmSffazy
Uyw5kKqEVYb4K7IZFqpTcLRqKZ8J8Kuz6HUUa2kymRjJpRgo8s9eei6BWpO5rFLg
FoKECj8D6hlcdcpQcnZI+mo9vmU6ZlMAdDAfkp0OpUi1vSjXkl48SjLILloi9SPL
oPjbw9mS2Zf/h3PLwvdWgYx8ztBEP6KN18/lmu8YimzSrZ7IMKZe3xesywE+FhzW
ny5577zbSOp6nOyVxCY5lDx4Ic/XUIy6lrZmoBJbbEMKtHZHZ6JaKcRmgJk8poft
aQkIm9GDqB6luAibx85v5BBcTMIJlzObVju1WvJM4fEOyhah1320YyZV2hfNe586
kYI7DP1YpX6x7B4WG9KzfLZZNUgaOGvs8nmUcBayF7mfHIKc7csR3TFLsc38xxg/
chyF7OoTTMPozSqnonLPVlPe1kbWw0zwOehOlaC9z5gYt+O2qaKK6lb4O3m30BOa
TTWB3zmJETT9TtNayhkIfdhRO74auIxiQG2OWZc4wMW0N3CSeUI2MhUaZPsTqIWB
fK3/V1til617jPsLLlp/R6e9zJHVFE0xuOtzQZkhLySvlta3fUiJf9R/YRsfFhIf
0sB6GrQSTgBHTnWy1/A+KbIOl2zYhzqmMgouvnXnl1qv4YUWFqZ52UCPzU43IRVT
B3lHk88KWlIl2X2EruVFNJj/CVx8/KTbYNOHqCyDuftdbZt+C2TycA8czC1IHHon
8ZVScCEle1rQtGqc9Lb5DlOohrObVnUetPl6TgKSgj4Qx/zUlV0ZNHf3Yl2yeg5n
t7RhPjGDSvPZ3htduDfwDLcgqT1RE2t/4FBgDL10pmMbVGM+znVhRejikeAKk4sl
L0AYaskqTV8nxl3VLdjRYvyFeeiEiLsR4lyycHqAziTA42CfvbkAWYwKhF+lSB3I
zOiur+fkXDNWhLh9F8Ne8Q36GOSufkuBnaX0B5EglTfbAGulxKPY2Fq6Qx/eS6RI
1Subd6BSPeqHGYN7fs5cOpa1Ow8OP3+es0/E3SzPk+5CI+IfD4xVwLXto5PeYKhe
5sUwiac0NS/w34APEIpZb+n3fNQEbzWsOQU/BbTcDI9WkL9CGBhcKcxI8BNtUGXJ
o6l7GfezmfR8JXt5GJUhalOgdoKYGuFN/tkSe+BQDl0obrhb78E0MaC8zstfZBHf
N+wv9D1o5Qg7si+UPrq7/aC1/bcoo0zxCSJRQ+YhH1xNa3gaOrCrIXxzrUehZvT7
djGyUMd6o9eIIoehdIuylNdJSYTiSsRdSe8oFwigvxuI7bkBc4bOH5gcCnOIqLiP
xoV/D9zs8bQ6DFlj8BeZgmk2IuazQpZZW2ZdzNtvoK+rCDtDnvgfXDRP3e8puLaA
rg5FZ1vbQ4DcIr4OGlPWfyvrUxCln5S0CYrczMfB0hSI9gvRi9dN5YkgraD1xZ44
TW8FC/2S5YWeKsG9nSjNfBP52T9rvsmIkKbzDSCfhCR9/m5pC/LI+4Gqngus1cYc
luDXETUiPoRsmhBKp1t4Trtx6GJFq/SGkej1leHPYS9C17kr6N1Ti9HBx9FuRhjX
6MLBlfBEpNvfpwp19MbDiXncQ96oIrbMBFJV+EFDCmr1219tuJjvSknrm5VaSJ0N
hrIWfkMwhb4+XLh0YsJe/O4PNLv9ohB8QqCnOMLr1XviIhl5PWU8AS//DoME94gZ
8p92MS2i4GJzNdqGILF8yqRdsqfpzheIJYXWxhzhFcRwVZLETnPvvquIqchS5gud
FKJGfflaWxloZVtoqrPyzIsLCjkM+w6a7qnZPiSk4aNcNjV8VIlAZUU7HEZ9VZye
qBWYgjOKTVRDMRKdocndXJ74tVTXdlUyVkqlPLX2Tv0j127etXJeScBIXQ0HJ9QZ
kUmHwkf/0LKUgyZrvWq+hQKbcKXALFxxE5wQTFTcxDOSX1jGQqx27crHO789kCuo
vuJVJtjV0fEDyKKoDIIsfc3UmCEoFf13g2C+K1fDUIRa/FlkbhalLT6Q2BK73cvB
VWs9M7A6UMvOfKwsX5uMbbXrbJCrYU1dOoSwEAWBxH5a/3vWayF1aCpRowPeVoLY
88PwSEvbHLjRey4FvizS+ntB+Civ/MkHpNeYNz+/aTrDW8XkUIjAnL28Am9K47y+
maH29MxJn4zxgSzU0tOFnjAfAP4DmWdPhl/1vnm212KFSW4NfHI6syRUnJD83aLu
ztXhPZBdvKOvoWbK5d51GF2Qpx0xgE3t/EuMLtf+zVggbOFHJ971pHu3P27ONKuT
hjPvY4x7DorAyKf24cYRJoAi+gktGzqx30eVnxjT2Gxnc9r9JCz+TJP6rMHzgx21
qqItV3QABl48FU5GDhvDtak3K12mWIBByMTfAgs6qNYJYkeU2tWIXBWCtt2lzIYP
cLOt4pWwU4VwRmkbVzAuQpyjr0DkoYa41TTA25bK3SK8okeGV8IdqhXRPBL7sqGX
onuOwwIl6PFrvnuDikcGvqkFQV526sftBPRpS41SakKrqIdgm5vXU68V1WZwOCBC
6sN+EOsaiDTVNyUt1+xES5QcfOKka6RFyv0efxoMAH09TFjrunLzfbROXbm4Zqly
VzNyAN9p51K6ungtTvI3qFao8uuAdk8cSfm7IGRrPXXJhA+BkqCikEQR8S4H8L7e
u+Z3OGSyWX+ZS272oUhyHe9TFXm+UAAIGmNvT2YYpNvwIXSx3hEFbFSTCg+hNrdE
5i+MN24y/bQL/W9GzYRTqOEeaPkVZ5QDgNAcDPDfGGxJm+dYooST0f2jBiy8if1h
CpoIQ+zxpUUCgoIVIqXwXgbOzJsGMF5Nn8pWwv+1QDESSpXWo2lt5s+2rAA0SDbd
j3ZUlss+2ON783RtuxvrLfJrOhod7Q0jaKjeRCtp/S3J8Dnx0XUUTHXujqRywrBC
OfEsEk1UuS7C2pHC46mCld89xHdB7FFZ5j/9k8b7A4ZZu2tc1Zm6ffNErzNnyZDt
1EUIw2oMs3KMkAq6Vrf+0gyJjBWpyxP45xQ58O0kQFOw3KCFfcZOXRK3M+5GuOUY
+x/PUhEiTEd1owv23wI7YwrlxqJccE3+0EyBGy0zQfIOlP+y78jEC4iHLd3p8Yn2
kczLIkwEwolDGeogB+U6Bv8QjF6UyG5GtvfDmOXG5JEnVFBTkjIAWcwmUipbn0Q9
FtiMAOSWXj4In8HQCvN+uIglvfdsWCgA3xtmk3Aar8i27RdfBg1N0itUD1vF/3lG
zsymoxfqCahYFQfVZxlodd4VJazI6a9baRTxWaXZBP/YpFF95uEu0Of+xFKS6BMK
dwb9RqtCF17ZHKsfqypM++tO3Ja+wo1nGgzKpiB3Tr2HpKuT7c6Yzqr8U6XQpuJO
d2xFl1ARdbk6OErYYRRohNvVWsa1T/tW5fZKtznTe27o40r2id01fmmcmDT9+Y1/
f74dh5LXykfI63byghVTeW44+4HxyiOrjl0DUNLYGO6kjLNULawrZ1WJim2J+dqn
nrVAOJvzMoihjppgAwIaQY4i/TL25kujJZARQs3XJ9ZruVVo4+qEFH8+KJFd68al
9KxqomudoynfhJSsqgWfiRXjAwlA77+1feZq3pzBq/BvYh0w+l3XpbwYSM+dGON3
zem5pI+CWBajFyoar+SQxzk95ifPx27agfWiFWM1UzkfnYpPzXpmKBhcjVVgwXUr
nw9rjfpQLvngi8fZ3XYUOS0R5iueyF8y9Oy/AD2FlrZAyVWpC10FgGSsV4WEG+Sq
Wuf9U0c9TnG3Q6Dn4Lq0psK7u7tDkvh9PjegZxy75f+WQb+X8MCAZzEA9uoENHlX
zWOncFeBu6ZBmVmYcZ1YY5OosBiH3dGwfTH2qeV5pS66bYoKrQg27tk7CqfB39Rm
N77qbR/ip0DnpsF+5UTHpfq1HxzhF9YUzzK2fy2ewprVHYR/LLvTsAzsLDZ8cehw
A+zT4JPs7JI9L3GrJL2XfYIRlNN7FNG/KlhcBZfdypAYcRG8PTSm00nsaXvfh+k9
oCIM7h3ikY4Fl5RimAFTPK52OmVrfQE9Z5hsLKjjc7kJhfQmoOTJqjRNQr5uxWqr
AmuOSQv7N7nvkviQHirO6Jtfp1wbf4FdQpSLbWn9MQq5y1UJw1NY350iEQObl8e5
qmMte1nkWJz1qi7099pu0KjRD6g1S8PnShMv1QGAZBTbQmHRMGUfjkZ5Ku+rvTZ4
5el5Pz8ENg63aXlNvzT84v+KlxPV5GW+VPv+TI/PvsRCzrVxWdYVG+yBBfYWBRY3
wHeEJkh6tkorUb8ns32N6RNJUVVr9G92KCFpu7GZ4vIjdBOTmYGyh9ymPzd1nSYu
g0dMEYOZnxLcpHFWGQNKcplk7c5K28Xp2pl+OvGwU8ozO7qAddpD3rBG7vkjjZOR
r1FWl0ly9C0oe0B9fEKbtAmNcInyfl8JVdFzlBCqO+uyg72Fpr4xccv+QYz7LsJz
lIZ+FiIbeoW71edzhuf9Auervn1U5EGnAhABf0lYfyTcn9knGXHB2lXAbK+/fB4E
ptPvQsg4gTZ+U6uMnqr68lANmGmdGLhUveUFeGQEKUAWuFYuylXLzLdeJ4BCUo3f
ZDt62V5MiYYGOrMZgY+E1Vz8IEYdsfMtnHIjRhgofHU0/Dl5xkj/CaQRa9L54oJt
CwMuLpmmCc/IjrBIAR58NmqZNV52xF2v0ZVtKRs66tknx08efjPrJe+RcQxhlN+2
XkUwSg/a7ZTCIcYvvnLmQdWRcfE5mYAQY0yYBJDDjQ7Jf3N7xq6e62fExv31lu+X
pniPTFkzWS0zGp6kji/edNltKbQyn3ZwUrIMhqRPFOphtPOP8Ovxbg9J28wyf5Nt
qR6V8w+cdL+PwkcGPJy8onD5VUkMggRbsgfk60leh3leC0RUG6I49l6c17mMd1mt
3XFShcKlCnVagMFBVU7WjS3l4i+b8c6gU9ekcikIs+3Rp6BPknxUWaJdMavqGJwG
VWFIFfTdtxk8v5zf0t02yEqGqBW4hTsNm4zgTSOMsPC115gqK9a6Is3Jgw/RR1ry
c7e+1JH80UsLaCEAp6rbjz4sfMOtzsksklliM6TW6bbIHLig0xFgeAFWFTuP0qU1
5RCw4+Yb3/J4yyh3Uu+b0Og8+a0OoWu3roofTO4rV/Y75NJ94gjyB6mVtqyVC5Vp
bR+1Uw7QL9i87teuk9lmardR7NdanzCtZE8/Z0pOzYMafrVirbzlVV1aZlOciVEv
pUhO9/Hc/MjIxtSUyeCj5FDRvVJTfPEHCpx4Cf1gzGhm48bxSBQGxUMc9iQEWtrK
Std64n2QqneL/F8pHGuEP7vtam7QU6wLcuPMuNkiBfvbTbsC13QcL9Y/VdAVOyse
sjeksBOwWhPOmchFaMGNl9JiwC9YmaFB/nKK6IZ1fuNpjpQCpEciZf8hOCSZBK/B
k5+La3XVfgN5zztGx5k7QI5W7oAOIeAPDS3HM+L4oXaH9WwVpUHFP8seXRbNDAYY
PD7+R1X1sZXz+PmWhYpXQAoHd2HkdmEArvdw8SuSLKQWk2Wbkkb82Q5c3z661JvL
GCrosteYMf4B3M1O7kGFpJV4xuy8ra5evITtObk2Ru8gJSQJBvc52olkglYAVNx5
4EwAxYw2+ItrQFVnV64UwSHys0H40VCMhg7IBDhGvcMW1agXqSJB7y7LcqGuXYK6
1hvxl8DLKqKxv52pCRjM2He3VvR9I14F/eZ10+ubCgRLEniI5tuMKuXh/5BfV3ui
wIObaJrXSmONc/r3qpP/7X+NJFfrxpiaGIY5UUP06fkRE4OMF2KKhzHkkneYm6Ys
decHnxvtR8ahWUbcZAc3NAPdxx7lx1pk8F/GQwol56vIGuiyn/SmgC3Na98D3ejt
fBP28nTYReHX7Qxf1XosCo5SPe9npCHFTTKzpzlkXvrMkPZm8N4izVT8WTtjOoKd
fqnb+1HFpPaDazweRSW3Y54oL+q/6WtFxeUOgZw3DR/oBi4DDPMzEqqgrESKqpoc
FgylcdzdSSgD3IHi3ixYvvWJuqFC0L8+3LadlN/QLDWz6btbYEP2bZ7yeBt8vmpS
2zm0MPO8YoGofrYZOvZ1tVsGYg4BnfxITva6uVG6vTVgesMxbW2PWcfEkemj+T2K
vWcYbspBvmACjJZHs/tyqeggYflkO8yL8EYf69cvwSYMnXRX/8HC5mmoB6cuRNzd
YkbqFqNTJwRi7FKlsmkewGc6O5+NMl9cFwn6X39xf5LPscvizHN8QU40JOcgQfI8
VEgDla+OGGDkVfzyZkUAsCrrCQmQp6JU3RNe2GlD5GDRnFiZlUtU48rY43CbDJre
RfpLGNwBaGjIQ/Gh2oCRJXBI6IX5KnoeLlJvrw3jKSk+Mp7eEgFQAGHC0emOe0xx
RfO8XpWYnHSnZgRVejKaOP1QH8ar1oLpCZF01ZzeTWtgOKQh8oJ8S4yRP53S5DOp
LwBWcbL1r8M/KG0NbL2MtXnWTDwq//ioJXR803D9Y0kKbFHiUy9JVBznVPRykz1b
+r8LkyLA8oTmZKAPn7rD+XWrUsPbcgjDYrmlWn1cHWozkVsmQz+XoJFM2xuWEg10
i+Ff/iJJvGXxgpYWXDEHL3xHZ5JNHQMX4mFXzX6HqESYkeFB7BHv8Axli+kXUX+B
VjVBI/D00t0Ycamf+ch0osxmpqWQUm4ePRPdWAtppLXBGZyiaInzFEOYYgz8SNuB
KmPpKEsvuNsY+ocF80Qw1hOZWV5jxANx42NH4sgAqZ+pIK1nvwpSRMLGG3/PzKSy
YmuMk0r1kTOuasZdBO3BFhuSr5a4AhfnWf25wXDaqRFLJHE3hJujFl2n//Tkjr4N
SZFfIwENSXm+Te0eES8Ddh2FQ4cHklBUrWDsqg8BEGIo47bGFf+PPKibVlTeydrK
2AKRlsbcdOr+qpQCocJd6MoMsd63EVYqIjUD5rFVugEKT9WJPXCNB8pAIzb22qtZ
au9iFbgpFmAiSKZK9sFDUuQ7ud+IDwg33fQrrFrG3hBNSTFVGobptVoRXuQZOz62
iR6ao3ip3SnEECNGefZCTySuVGGoswRznelrzUHv//uzfm0C1UB3+x1Fp+zUynMX
etzrdQvjpeICxgj14hwN+ohqbh+rJGpctm43MWPLCjkzxIpl3LcK0/mLHXli0pzL
+SY6qiVKKqYNGRpnXCP7kkMfq3kWrMJr1eLP2flWRmgVSdEVq/fj7HsCjoCuWhPJ
nS39YbDgAYrph5nT/3r/Z3M/dbbFN8Smrzm5M6yzFAFZvtwadlukfyAUzoGthKc/
qIQ/mBEookQGahhSVsFqPoT30okSGm3e8NYNtfvut/qdDZxo+YwdjRQgrS5pXWHA
q82TrLSGylm7YSpGRa7a9CUx0zrGper6flP6B+BYSbeU7bWRDhVIehNiNwTVcmOP
Rb71tmfhPuDzOhQHPsRWatrYSDxApyWU0hgwmPjp+oqYNfM7cvgFUtLIXLkrrzsO
Z18iQZILKfSSz7JLXb/wApIWmdGOMXK9D5nXih/KYSEs14hvFRoMlSCRdJRdDE/i
tCr6yLdrFreCxDFTdYRvTv4ijvGb9ZUMqESZuZv6ohYfZlAVkvu2wUAaUC4Zk9BC
NY2+bkjTgtmGpYB/rxgE3fZ6BzVCXt8UhND4AwVRLtKNYa+0bYeM0sSUY4fn/ns1
DprPyi7U5nzyFQeSe35oQbKvoPycpLiFZn25tiZyn1q3puC1ONKVriNv4LLvE3q+
t5QJVn4EsUvdvKBPjOdq1VsRY1gQG3mUf4vak+QY2Xgq/5kBturXFkTzIdQkT0Fa
wHIJiPoKTxFyOj45iTv5ZlFyIvzrDLck7t+zQytn0B9mVQZ3nekYSOYZT5iEOcD4
rF65fNmBEK7uPBDz31or/JN0nwEUGQM9h85kyf1WEiBphLk6bWn7mZ7R6w9gurI3
8Noy9mX71ckrKeMLk8pWBOIkPUDRljVrlEtLMkk2nwWMmCUNfiLUzOrk4VvRcHEo
tyCmpw/UpHjvNhSWiDYhKrHB3RRx9b8e+7UZPEv8qLoxFPZUdU8UBhyk5+es3Y1i
Kg0FkMmyq+mKVhVtk1AW0asrcqNaWje0R+zNjDC6EvG4a9+tOLvbM9EB1SgYYB2/
3P0XXYBEvO1yzYIuMa/OlX3VPdZTKwEFoGicfJNOyvZiFm2RES4ZPLG9lYXM21Mb
1fPQA8dDh1EBqtLdLhfjrsM/Jf3oIf6+A3zzqHgifh7Wqo2DGhOEQoyqarOQqm0J
G/n+YCvUz1ylhwOGrW4QWQOHHlzZ6sPDDz+mokNMNhLPxAonrFsCO9LBI2ZbtE2e
irvqF20hJuDMynxkLLPqM1zTsXgKrRNP8k74RI87XRjmzkMzBRlUrrkp3l2B6z/+
5eAIzyIigCoUB7+nG45MhepDXa+DfwFEKhUB0Tvzv6E54p5qaV0sfwEwElsDeJiq
LRtdvrxod4no6aevi0vUWM4TdgwbkOX8YNGMfxnKxXBHosLwQKU1IvFHhnQfYQ7+
LVBGs+nLDtmEGbXlQUwNi0PIf2R1dNzhUF4XIFeIpYCKdOB6tUdo8ObQg8NuBMtt
VK5rKkBvSm4HYKjTpWAneunJ3k99Y2kgmb9ckoEkfq26YCdR9BUkTTOPJG/sA39Y
MApaiFtBlTuxUea29GervBHKncEVsnadpE4l2VJ3yPNuD2/gTs+E0dyE9YCw8eN6
ryCu10z8NZMsLPmenU7NWrv9undQ7J5wqZ8csK5hzyJdlwfhtH86uUl64uAS7mc2
1/EgXut4R11asVhx1CRycLtG3SVlhnw6NngX9RxEaNStUmR07IGJmIpOkhBM7jKh
Bgg7sQzxtZkCTXoNaPgGtCoJExOFXkYB0efZ1w4iSIPW2dOu+q2SP8cCBQ8T+aeS
SeIjOJwp7rMiQJkyLv5DCc5w7CCTvR0kN3SF/Is4e12tvrpsBBY14DHelPE25wkp
xCfFG4zAWX9ZWcUpsD403J936fkHdRGIyIE+HkbIZZSC25ByKg6BHmP9CTTVKd/c
V0mCJXveVFRtLuEGFrtjjQaW17qRnWRacbJVkF2e4fjp2sR+6BDBuTKha6dbgWp9
PNWBguJonlQsd+Rcdk7gjgot2EJ+3uvWCoeFQFic503AuO6LmK1TseVA06jgfwiW
pbT1eC4Y+PaAldZsnFa8YkAKnwi35xX48idjFVdQdan8yjJKikGfXFU4xDa4MnqD
xrwmeOQEWN6hKx878t8GHDJzxy6ak1iVMkF6tTVSvSW9/qiaGJVHqcZhY0ox+/yh
J2S3Y/bMvX1jgZLgzc65CyFeeiC0eYbX+EJI1Ajti6npNVQUpHpYvUrWUXAZWQg4
9NwwnJJFkE673xH09x61aZG5D94GR0bx3f0d5A5ZF/5/Ge0I4L7xmIPDE0DqjAnC
tj4+HHXzY8IxxoLVKl578Y1RSR27IzTWZ6Tf1cPuRcLAPAxqvpVNgjisS9WNVk/d
otAmSO7XXmmfXwdbq22LFvbwILUoCFpGDHbbCrTBsZDmRnmNvdocnD2sBUHJ5yxt
sZwVZgcs3UJsTSalJip18mYHR6X2f66bNFY6rVIg+qLxSQHIN/tGjbtA9SedBO4M
1Co3ASTp7BkkYb/HymZmzHQV1PQtq0mW5jD1lzXnof9+TTje3HgmNSdkCH8O8Ora
l4iYvWJUj1W+zkdw/wB6ZNLfZbAI6ah2G30HQy31Q5/7F9CYz1xJpttMer4+N3P/
VG871mtV6wNbtcK3hOjJ0oQqy15pj8Sldb//9SCF0x/rM6vdDYCC8Us+Np5crI2T
MnlQqExCgzeOkPL3j5wz80K7TcmCplwefPwlbryzWMLfnZV1odfcYwzdK1qP2W9R
g/Ihxjl/KYMPnQmp7fwjO7JCv4grUnmG1PXzq7w6U9yOJnpTXT2x0ivDdHZEitEa
irHZrGH92zTE9PPzg9MUZSWotzttencvNPLPmUJVezrVIB4BLSEaWG/QSkjACblq
3BtMU91lN8Wnv4NmtWq80TY6O1x0ymZ2tCs4yilIwjkEyFPXQFK4m/Nn/Jxoizn8
dEHOeJ0Wuxg+u7WS7L+rCUYhSCnbaEpKF1GqckBgThRnfUyyn//3O//ANY+AjGKj
SAQIacn/h1HQMvttDfFaeAUPKubQndjbHm/tyTrOP35z8A0ND2h2LMyEk0wHjhWP
2Ysk4yVvF9HdVfPBIvRpi+w8rcTNzCx4eNOuXqXvQCLQhkAxT+a/XFHccJHTrCbg
susWglIz1fKwpjfgymxk2gv/z1cbQAghjloZKnOz3St4kLV/vW6nyVRKHORICoBs
wA5p0APWlSbBOP20EfOcuOXr6TcP/cpBWa8rBNV5MqL33mqgVwAhuY7cnGA4F1lf
0TojH/t4PSuLp5rXH7OSwVU2T9jtLGTaDYcc1ha8331wenEnbHBIjo7B2mNqyO5k
xVbvnQhqdfs4/MdWVpQD5Viq8av9Jn+ixck7iAZemUVZvKmAfH3f2tQCY3H7WbDR
3sxFQpzZO7rMykjAYQBVaD0s2gKBRHAy/yGofutRb2y7xvZ2rnk2wxO1qRvZRQqj
CDIV7BAcBkEE8xJFaZPSafS4x6oIUJsKaL71UnUDN2GTT9X+unbOFAG6Y1nqHyVr
ebMkP8RguWT+RtyaVfxJ4MXEqekVX+DHEeCTwamfpqQohEXTqbEzHn+5pvP/kOGB
XlKB22EU68R3Yj/4e5uY72Y11kBR+CV/BqY5C/5E9MsSXNclqBRoPHL8dtlFy6kC
e0WsJFkdGSlkMiJ3i/GiQhnn6PQxeOngvB6DOsjoGMCUc/GBe+4giGKMxUjFLlPN
3gsTNxl6CjG1T9WiiVTuc/nWHX/VU1FOevNl/PUbaEXKQadqPoNSChh209+K8fa4
AzFYxYskuQ8tkeLndBm0D0w6sC/vPINNPEfUZ+cD2IibpNL/JaK0swfiZiwmzGPM
+Ehg4hGYBiQxhlgdg05fwVbRT1YPsSfD1hEAUcq/zCK42ogWd2MUuHSyDsFsxA5n
kQ3HZpAzukMK5Kceul9OVY9ismaxhhrDInzOu+QaEkW7BDPLwCv0z5gHBLf0N/uH
zN+0BMiXg4X3g/Zruty+ejCCCrwqlrxmSiOPfsgnzUSaiw+Tl0wvyKDXpaBgJ64j
hp84fqDuWR+oUMJvU9eTIZK1T0DhVD/LHL/p3JJptw1sI4E3FPpB4voiNRc7MMGt
clyqH5fWQDnxgduejCIxfpaoouHqR1I05OEcpnQ9q92HT1I+HqASnU1nqsxabHcu
VZ9sfBMOKkY7ThOusa1DKg4MwE7t8bPOZ/K1nLlV+j6Uv65APMQYwR18+4H+KbvI
Gsq6YPTEk7ZCFbsJi2NrW5DSCwgUglmtbLtJFa4UatgkCMy2Fyu7/tCNRoayEul/
Mw5HED2hPJ3pJuX2Caj36fM00ggOBhF8uhRNmGzs75TG4A86ur4ZJx0UrUlSHGAT
Kcfi0IFk9saa+89J8s51CejCd0DOCC1bKUvGRlt2ShB5/rO5FAHYdSHGx1rY1Kev
I7v3YY7Xbj+ICif5Dl1ofCfxNCUUC2t2OnToSC2LfsEDkiKv3oPey41xmH681ZPS
d1c54CTBQ9KIOn/qCmj0xc6gFzGFGTiz7r2TKiMwwpM2rVIPAvK4YAYmxP3/Bz4e
DpN+dKwe6MMlV5J2qvj/dpPVvJy4JlPECY4GdTMyPvzfhHx6A7Tu/v0Tb21oiMyP
AOH4EykZgfBMkCMk8qmi/rBCJdN8/r182qUqFRg3XUaLnxTq0NgaTL3VaS6YHvGK
t5c7BblGo+yEUJvoVsVThp4Oywbb+enerxDpKjXImWldM92hNACWl+iv1U+ZRMrr
VqVjjKlD1Od8n85t6rjOFhgcd7ICj5QqbL4dKh1cXM9axY3EFBNBs5VVlrumXkHi
4dETzw+wczvoXpK8X8RaErQCqSiG7AIc6jMQA3YAgO+0TrqtqBgQrvrHs65Fyx0u
kRRaK1Vixu+2bWyP99k/V6IXnzJ1Va1yQ6VAgOpQxNE08ZVfbo6gmJBb3SB7/yzU
ZZvDFE+Z3U3xNwxhE3izxu1cs6m5JR6j1AaOdQ7bqV/rBWa0TQR/HSzPQlyks2mt
skC/LpRx3kV0CMdLGEuRFx8T9nXYkZpBxIfowW/cWqCZmz4pIT2UcjN28IvyfK4f
BrkWn8TVbGdJ5fUezheFuZJYoG5zxaSLeN4LQleesvmsbGRT7/wXjTLjnYQXL8SW
elh1yOory81La0DNvKgm7iynPiEqHghHoMtda677IrXXOpoy74KDAwOZz+6TUBdA
w0BCDh9fXw6ds1wcBJv3JihQNAk+/DtOLxm5Fu26RqbO/XUCS1uuSBscw+bjey2+
d4Vbk+tGpPA1nOIvRoU5np/0Ogl9U2HU3+zcufNM5xPXMUPVOvmv2nAzGss2HtU/
RPAVkIQe0OHQF37ipY4w41INOpEKwq7BTkJfjYIFmRkpzmQE8RV/QPRuTSxZUIg4
McjLhL34V/b2gIBZ0LIsXgDkrgxQNiPNBA0b6udXa4IW3Rmf5cBzkRTiQGKOAp0U
6nFBcx9OHYma1wwvZTpkPg1A8EduQGUGw5NR4T2bOQwfKLagA+G6dZrUIL5AscTj
LHIX09qHEWDuAwfaMb2utlmeeVu5WMp8EC1m408IpYtm2tk3JOFRum2X0FxNR2mC
r2Ve0hKUGurbJoFp1xieCYtQjwDSEN+zNQ3UIZhvPZ+OnLqOa4z6kT+kx2HSw5Ck
j5A7tX5rI/OLg4qXFMZOi2upG9XzeCzbAf8rzTMSXocpAgdQhrCDf72FQu3+6Sd4
h7lJKYiUJSdzcmm5btZNuHSbASerkcXkN+rEunBKPqpbqNOIvj133VwMMt1wRCcy
NkeBxPR86M+gGciU1Dfc8om/LoNdBhLs1xWHzbdyVzBlyIJptscO3vsp/ArsSB/s
nsE+OunTF51m74AcmTnR9hQsNW0KCkSBlfgSvfXSxk+Loj0ivkoObwsgwLL3Sk8r
0UnBe571xTViaxr6q7wj60nKeZ/iCXFnjKauZWL/I7eu801uTn1XEPsl2DaPGrot
xOE/LNXOX2NX3Odng8+1nsyeE2YiqUVW66495Hqbp+7B+s0AP0Pj7HCkUv/x0wRM
WeIZOhpGLG5ZN+ulT19Ukduvwc/IvAA3NtJjwlSWc/Rgg8sHzUwBk0o0vMvjD0C2
0b6z5sp1AHvRyIujw2soiec5lf+iSFkJiXCr0uz8Vid4T6oeTcQ2jGa2eK/7SHrs
pS7ELmTJitULI0eDHhrmopvrpBasG8PwIJNxafsmy7ebPt6riYUMMgiXjr/SEzyf
ae35jnokGeYs2daICGSzvl5Vdu/Mr407f0OZv/QH8eP+o/gpGRFRGLwb2u9LnXXB
aVfRHjPvFsN+hHH5n+VUw7Vw0RRhG7Su+4LsMS66pKtxmdUrRIgmcnpjwH/JsHGR
WWvdqZtfBMlVBldcdYftHgPGklqzwiawHZPsWXUhD1OJdsMmQQZGsUmXmLEU6Jg7
Ee29l1UOce3suYZ7wxzQapXChCTCvcWiq6rc2VkYBN16j/bp7obf/fPYgRQzu9i2
SPaADTbQ8rIO2Fy8J2LslA0sIiepWbJvy3wUhL6ZicQpRJcy4OYLod7oYECPwFHV
Nokaw29Ke8EkrJwExRUKPWvaGaX5zYdYCr4NzKEaaBMotDyViUr+C8+SiHpg8lAw
gRZCSzhj/4f936WcAYxsFrutEEjOiK73d1T9ur54TJiofL0yNBdEalSZsRHW1cN1
Dc+wVDe+wjcsXzkdrBOsCDgKtkqk6WnBBgIQ3p9PJZ/N+j1bW7QxeKsSpidSgsqq
6jNeDaqu4mHcPlB0TnBGvOWJrGgOTf4T2vGWEEyPGNPQeKlXX61jgbPn1oLdvX1P
k7PwSeOHJKTi4W1/4Yd7SxvIDRqTNJNItX2uLTb2UsCF5wmNj6d8RkYrmGOG9egC
d7aFY9C3xH4f3zfK4yKEP39Yzzbpl2xSSMPWbIXmqpjhNcn1KFvcJcSi4zZui1BZ
8mXlpq9B5gXwbafVoSUlLsVOOQ0p1m1D/9S8lFusO/+Ni/IAfcqfV9HSeVOL41If
7YYS8syqw5zGburHrDD84f6aM6bVV3EuTXvH/OJL5Hnw7n0n9AB0mWcr4xknF0NO
IIIxjQiiuTTZ5QPmIhWq5sZNCxN3d1GdhiqZhczKJJdIP+dC3zlsIXfSyMGb1HTL
0TK32b9F2YMIxm6atobIT4RFl2/O90/YGvZS190OMr3/KZ5DnHPppFUKuWMzNG7w
ymDZAlA1xxzuTT5zUfI30sqp5f4N0ektKrlsnrcvfCq56VjGPGpEQMtti8kte0TL
UlW9irPfEFErCi4CCXp6RCYlfbkcrzlIkjl4Xaj4STgHXTiuGK/taiZ85SAxve9E
HGW0UgdCso6nE5GuGvAaP/Eg6q7RBCU/sTrZzKNhcm0zAPo95P6L4XDLinjXHLcx
l24zueRwOVbFJFB/Q2UzgMI6GUVjn2KeQzQNlgi7+Ip++WSNp/1SELASj7VHeduk
CBJHG05d2kSqcrOC0yTr4uTQ9600Wa+1rnHTIxgU9yOFuHQoHKBozIPXSX9+gnqw
BZqIl0kcrwOlo/9qgzdl2SjFA37kFfTsk2tr9ENSw/qSj1VxBzMBm4lN4E14wOtb
3AO8GO+lo5bMroLmyyLQLVwJwcsDV/DuQUkvnObmkWDki0LPfJxKQSBb7wDpvkQU
Nianx/cEj/u8euvb3icHIXCnbjv1EU+UkCwbXbrP1380z6G+v7yeyK/5McwxKgq3
f52cOPYkMKn3p4qXhWxBk9Bf2SbjMIYbpr181t3NXuImwhuEsm+gs0MH6XJW8AwL
kveqjCBJj2WjXASX/P6O2W7jMYam2OsEjgXRs9Tl/Ql4i5zrdjYo/IMVrvbNqQk3
qvTTRTpBf3Lchqg4l4T/HKT3+Y81o97wyXskYbaoaob7G5vo1OoB65PYrzLmhjzF
H+W7XI1E86cLdV+kUqlQwBUBn4ExIY1M7+VmVMbKNLSB3SvmFbBu8Wtmm5oPu4gD
X610JyEhfcgZJbNTcae/Lfmd+9rE+9jfOq/UQW9BaHgWffsmPV46OkdCoPYK0gvU
2RPkh0o7oG8pqkzRV7D7aOOeLRHmtj/ONXlLwCYZjeA5CZca2hQxlGIft9wCA4is
1G0iBytE/arfytX+wIcqPXD5y38y2P971vM4AO5DKUUe1UCX+hn+rixJ3X8Cd23o
HT6ajmUe4tXQ7CjEEZj/BtEi0X/rMSBOpYtLQ0/oM9yX4VjY5R8aBW72vgrwQrZ4
DRfiigN9gTGFwebJvZlVPBkP0QX6SKmOtl3MtwHrAs8O4r6WdUFnPICdqyHlme/2
6AgB6895nyjvCo9CKi321EE/Cs89haGy5C3Ate36nAraw0EMpL41H29JF5UCOp/k
aqe2EXxp2opET6WhQ9uLqcyVVAxNDQ1Tn7gtqH4Agb2LZR+k+AKpFPNZCtOWyBXj
ITvfTXktbFEKPIRipPElM2+NvOsm3VH5snE3H6CBpiYKzWtI+1wMpeoa9wfxnQEH
wGrxectIt871sxav/Jex4GR+DIe6oGYVfnyUdPc6nz1ZmQjfNRvJcdyANOwfg7tG
WYfR1+9b4McSqbzMpbG8VvFeSFY39kxHV4x8+z1cMeKSHVrObjOXcyJdE/TuJ7vQ
Hh19LZbxC5S0O2wBdKRoOzW+4VqdCJIGZ4c0qSzKr9vOhPB7Fu6CTaJpYiXZoRFC
28p4UuPUgHNjcCXH5qzQ8ZaA/kPXS8qWIBs2e78Nngn2eJzQREOhdcMpLt++xzBv
l9w7xtkH8aSlyhD7FyS+O0vX1MIB0DOOcg6zkbZnM9Iq+tXib+joYy9b9zRRHbiA
LtBCzZdMon8c2vGEkkAwqTOaced+8l3p7qCgyCcugE1XHc7wjTCWkzQ9PPIy34I9
SyfMP80CjcOX5S97rGEYqdJ3yIEu8yOvk2neN3GHXYSRODOUdOydPi4b1Ve0Xa0K
XLyjmx/+xflCLgc5BpkC3ylBqXekQpXfKXDPcRxQig33cj94iZA1lkZVqzbo6riG
lEsCBOG+udqhfbouA2rafiSvMIzPu04mVaGLBZ7TntKserQ6dHKrkHKNZi45XJMP
M34xeRh1gLw7+JvgMyBt52w8lEcq/i2dIEeFGgfKAjfyTHzZ5lVy67EAI3O1uSi/
iR0qVI3e34PT9mZ/nyjplDLL8jjX7ZeEMyvjyalS35NywIBaUvH6Uo6rHMG0WVzy
btv3MpZvIfrfFOV1w9pqYuoQ1o/OgNJVUiOe0OtbouMstdP6hCiKFECmGmQEwiBj
zpRkSDqbkC0WaSq9y202unhE7i0NamP+kYIGCwOZVUqB6PpXxxoXce3JxhDUfyQH
iGpaKva8vPJNUL1V65Q0sxlIiOye4fxzMDe/dW9IgzYZ63VrqYlJoMh5t91zMyp1
yKGF/In/8ANQMVIlVHNceSSuNNSAnfaG/tZ7J5Qt8FYuy0O9J1pJ3NAkfWkJLQcI
mb4EzDLQ68qiAtWx28vZfxvF9JiUP6GV7Fcr6IcpigqOjf4ISHpIJlvNjIkiITQf
UZl7WPI8haqMy7t409UA+1lqpqV+KCeiy+jPkWvG0PAah+NaHClItg3w+blMTHXB
vtp4ChCvcwLIXGYplXY7ccANQ1wGvpvUGlEZDIPTi5jNphhxrnNzU50xeNawtuPK
GHXle+thpnXNaVB8H31EZO18U0TJUOfor4dVHeN0nPGlN5ysh0KmJU7pnxHWoi+1
RSr/KYGzERZP8JmAPXPoo5n7UjGpktp5NfrGgfbnLcaEJMs1yHnaGKKNkC05/Buk
k6Vt8vBKanwFXG+84AvY9OGzxMlB13u1Rwh2aDb6+LizFHOdnkI4qRYa3hk9zpAl
N1eyZsVFAi5v1b6tlx50GSxfiOLV2HoA1F+ba9gw92XL+89hk8fhQqdTyYE4MqvJ
dhTkQAt2lVm+kUE0n7tGRgFcGVKnWxPpnaWm8MZGEm6GML/hUQyUOAzb89IFTpPO
v4WzCOdtCgwjNyKX3Xvo5lNbtyyzqz00Ekcf0PrZwdwWKBg2OnslW5v+pem63pLa
XkRQcAhf5CYxFCAQELtoGRkfIgLeFoMfE01dDA6mnq3qu9Qh3OAf6OtuILWfP8GZ
m3Mp6kT1sZ2TKW1TBAjDcUDwRZFhLXpoxFvXV7nRtmW3ATWl+gd37xWwS2IFTR5t
KhQ8TYADyCB2Mpd8/pNS3MxSrKTX9iJimsQXcAW5o92IYSZ7JH165my7JpEd+JzM
KDF95PWmNfRTr9iAdZuRgbQROGeoIZO4o6s5S00GxViifcL3AOb8oYFFblHL3NM7
p6whWb7T+tgVx2Q5j6gvnoGeSon/WSzeYm9fnYezplgOnsOQRg1dsGDcV4oy5Qlx
RNe8ZXC6YAfTeepz89TNymvdYKdMIM0l2NmxQ0czC2OAxXonOMEfvvjXe1NNkZKs
yaDq0jlpqyOG3/yHe61l3X84yWamm5YYlOM4T0vqfMpPOG71foaS7lEDLEVps/5e
0ohrQeiYrhF73pPoRn0OieofrOOyefg8Be+tj12Xb5VY9D/gS97jVbWSWXNnCd4I
KcJCYjaVtuqXawaYSt968S68hGLFkvAsF/9U2jWY+177/5XYowP+3R8p1W+rUYtB
kbnibzCavzjbhuMUmmrkCrswLCEa1pCeBqkCRcj0m2XT/HS4QB/omRSwB6WvdhYn
AHoezWHUhxlkZyzsykQxeyYh8Q/eucC1+K0T9Ya9VHLmixKb7HUk49hL6CIduaTy
fuFBxtWGdOB/8R6jlWuTJTSccVxrs1mS7HnKFOYZ5pieWeWrnWl8+Fz32NZslUfd
ExKr/olk+7e374e0aRcpIyGm/Je5wc1eMoArq+eAS2HScNvHN7V0cmXFORpZDphb
rL9t42riw7rq3a6gRjf3dBR5rDhpIL+tUCp+lPrZb6Jvmzzepkd5ZEQbQ9gpjfaW
KFLTDI4Xpuex5XhJVC/KR7lzSpP9FAlDtCyxFqFQ0iNsSVA/ofrStZ1lma6iBCNF
dZ1TSWDZu2QygPBYC1eIAcG4l3FuzXnYFaM+SJjsxyQPuOPYdqvUNNDtoq8NS5+o
/6DWKaEYeGBBrYZ0CqBgAzzX6FIiDoDGG7YxKFWs7tKe9BVyjYu6feyLKslYKnSm
GTe+TMxtaGrwfvwe2aFkTtliKwwaV+3OIpk6qJ1/IjtbRBsaLemnG/e98ZiY2RgX
dzmqdp+8hpYNld6fvfDrmF07TZZzlvS7O+cuRl6lNNzlWEJoOjwIZfE3dDmZ/KDU
dJ0YjUXUOjPEJ3fTC8SxOODzGOJxFlSPtL2KapAQn8U23DaiEe7iYJy8OVE0ZejH
wVuf70+KOPiFwdmrEUkwA2NHW3p/AH+FAtrfh9zaEu96k4wvf7CM7af+GnSoSOLe
U0A94RiBtyLWFpL83J8g6u2CuCxw7SJHWVuEIpF+d6wJO7iQDq79xVPhpekUmOKR
cjnvunJdT1Queff3dSx4MJiNyhljFDi1uO//V/QHgX3FUNrnlNOP2WQSSora35D6
L1Sk2gIFAPvKhyu+xUtWVqJnStf8yWP/AI6M31zAz+qqLp8jRZ8uALznrsBVX+hD
eat85o4KP5Cw4AsLGcrkej/eY5L7Ukg8W0k3Mx3i0OQFiCl35fyr5RxRCUCXGYHW
6MzlnfPtrj5c6TnyogHgKnDpLQe1JlIfvQu9P+i22jx6smeoKyeLmZUn6yLAVMKK
2e7daa1d3js29PbTALk7VsbqAuJE3Kw5uNaluo/OiAulT1GMd96bTCT7SP3DpgqA
10hagK2XiqaS83qofKHaIq6+CW1n3kVVG4xaTeTQ+JD+xIWZ0DApcccldwaGTtpv
w3OCS2VkVzDFDiaAVdkx4BlOw6DcF1WsDYy+tMih5lUqNSkDwZHa7JhvIUdnpC0w
s7cQsA4F/Oue3zVZETNyYqnK1HkCqo3V8Ox+KyB8+XIhU2ZwH+cUgcMrelThKkx3
4G9iPaw6qiEsOIE6g0Dw1Gyfn3EoQC0AR/FT7kjTeJCO5bfNcdnlnt97J33saFLP
crbiYQHro0XmEp2snEz1vYG+gBPy3An/HQJWj0KpeKeddf/kk8fZDgWEs4fH0gnJ
eaGva9u/3WgHlp7LHaf2Hvo/hYzdAXoDroW2Uv9kDrXkgW9iFpz3vWCvFq0mfjZB
6AGedv7c+VIYXb6DSD4lNw6Z7QkHvPYhuXWJxvQqeQUWQ1T+/aEaEYEQeyGy1I4L
q8qnOHWl18cKUvynSpEgppezE2fonRTKUEUly9jDv2bHHyNUI3+UNbZ+7F6Fgl+1
LsziBLrYut8970dX6WmXYmiJykjDFsYl20mOtP8bGR9j20jFEr/mmRdK8LAD/PU+
aNr9EPTOLFT2IrDbW/j+/Fhar3HGktV9PlPWK7nBteGPu9cIRr+THbrqXdzDW/iA
vVl2JhhiSSz38AFCSXj16DtKsQ1dMEBRjZqlT9aJdqfgDtPYleLX2BpUVPpnVmrI
l6mXAu7iscNkBCjlT2+zFhfQyVDBF5uj2Ns4FVesEqx0wVyeAwcrhkQSRojFXEFi
hO4REXTZHPTtquVoRAjrICLazCuhRLXxMZ5p8GnvJNGHzzNcR4JGXDjMSa8Le9kP
ENVo2QI3E35XhKb5V9OpveV6vANTL0QSgB++/j3mIlg4/+QTPjn5ExRJ5Lnkx2JD
S4JOGiQWlu0NT7Kbc4ZSw1qEht5Cn3zisdKv72hDySzML06/nnNEdbNOrn8Bz4Xr
H5P/8sBARFQxLc1tjW9WvhjxPVw7I96BPLY8h421evrJtLDDx4Ziax7vx5XYHJyh
muNFAijbePbv5SXzQQd0pPAjGcZiwA4KNVAR4kEmRYetLNTKjNM056KvzmxJtLHv
7+F7HCZDCY6aRfO/rgJ+Mo4LwdDC/IwaCaXiXszmgRYoEfaydJ8N4VyUn1tkNCje
W/t1elt4eRVaq/D7xCaSRa/uxD571p83DL2zylmBwMuZ+oSrb0jAes6QZonOVuHo
zLbSDNiNgTBj4m0E6twBHOyTeVsx7ZIqgEYX0zQWcZStCS6sjAqqZG0TP9btGfTO
2ZPW74ra0+6Chs97HjrRBhD0iqt0VyYP5mk35UvoE/ZzUfPi59grRwPtRH/wQY67
O7ZEMc9E42qBLULjlRJMeRdoRUM4YaJsgENM3qoaFxOillCGkAHm1ERFm1LuUjU8
BX1tPcYJp37kVR8/PwBufZ5X4NtoUVaGg/2jNNNbqndjGbbNhlNJJ6QWCWHLpvZ4
y5UwaVpVtfrkJuvpgq9GdytkmyXYiNjYMdNRpjwiYhW8SKQ7ZJXE9a6/6Tv0iXAV
lVTijGbhapF/jKEdhxtbUV9RDQdT/GTTgHioBp/LS8aXjOBOTkGLBfTFtmtJ0bbt
jFmGCNWPEIpx94z22ghft18Ge/ekqREyJ7/HPBAliO/ZHvAKZTbruCh30P5Lr/nb
fraCGG6Sk4HQeoqHg7RCIOdGgAVdveFFgJxfsnwJxp9ihG9dyTsWCYBtv2jjyqHN
XgZZEfGBqHz8BbJn4WfeM8e0RTFDKrlUi1NRwRu0p4oA29qTG4Z3ARAFaF6uw/lB
WtSRWqfHwcXI5Xmfkf2w9IMbS9ShccsKaXTF2s63pIXcvCxxbDxSXQJl+i2z5kzC
X6Cn+eLhxNXOFUR6rKntvvFKgwVlwlLcaJgacSdRcK3MIglGva4KROmmxVWKsN5x
EPKssKIbZQ+YzN0R+PD2Sl7n6HN/6gNQZSXA5J2UwkPX/rs2zycNBLjaHyJ00tXy
xI1t1nvzdCDzXDZBPCMu56Maj1sqtQULb+jfrYg3+FGHic3fgH85eEzdYecgtSqg
eY3Et15orlp2HvddNXgDEuP06DyWjW2AaRwGe9GMfMWrodOjdZcOs+MeWMGCBx0r
wyYafa67fpcaS/YqDltWkLk2ubXwGK4gSTMD+tWsg6Uq809/ncivQUk0ufBLOYQQ
s0NWew5tExsLK/qFPGMAcfkeeMOd89JilguAp7EwvZAGlMTHTVDI903zuTFrNP17
jVcGb2FKR+fHxZYvmEeL7HiQTQqiRHZTh6qfLewgHfNXW8NpJBbCK8ScdpxucB8e
oNMvPMpREvR303h5Gj+7Cl/6ClrcntOq+aJQi09eWSDu+Vv080ckl7HEZBEJQTBt
UkzLEFgy9Sc1/RydhPQFG46QPYS1q4m15mkDe0d6Y7RYX0EWsCi5fANXLEewh5nI
zqZZbOUIFnz+UP3+iN6ho3XDE95yNLsg8t+DIqq5xMh43gl40AdIy9abAqRTvD/T
Te2hs9L6dQ6AldWOD0g/lKmFETXGkX+afH4i6k+EIclUH0ewcMeSx6fJFkE/MSrh
EeBIJKG8y6oKTxleYiNwUzSGv10c3A0YnxG+l03c/hjcxX0tQ19wqtyQf3j5QtIl
1XXQKYqCeSt1aed7ky2zQ41g6X8IKeXxfBgsABe3SP+jmtFDWQbtdkmeBhW321t2
vjtWwsPtJ6Ps8t1Qoz2JppLjGzUZYqd/WLewaCXcYbsIuwqeI+e3Os/wirp7j65g
DPeaUHGi3WBHTcHn677w7pvA7ypw8H3k/5P95TwTQeXY07H4JbSQdhnI8nrF2HDV
BXo2FFWa3A6iEUCvD4YmvbTXx4S0OpF1O9eU+lN2yjpqiAjNSoS0QVlmZkmvVsF/
FoI0ZGEZFsIicq1ef1QRgpvTX8r8kAZHzDA/w5I4iMsEE3frMcH3IKViNsVhlEg/
c+b9fvXd9yro0zVlCvy8R81qYGQUpVlG4gZBBrR3aTWNlMXpFgVjIwOPvkdp3Jzd
NEeh3cz/ndJlwCx/arHXdYaYRKrediohCpEv7z4TCVi3C9iP1pgRqW/7LLLTX0cu
2SMbFstmepel4H5ZxhuDbuB0sPpGz19IlAMJYBkB4P69Kzwb7gJj1L96kHYi0oVD
2TVUg0xzNozSWDHS8jPIfvjt4qWgtiHsaSmtNgeHBQ89jrsX/fnWyHl9xdlhTvx3
vUJlOx3cLRsT+tp4jiwoQRBGSssCthv7lMSEKuZg7rRrAm6weCfdhCi3I4etyg83
eZyTZld4XNoCZD0Xw1i0Vuidfc/3/ZPnyvULjSpo8RK24n803ojBZHMWVmlGYBbo
36oCJOrHiQCMDJb9x1UjALwBm9z80I26KvtE7I0BVXcyfrZYypZ7mhmnXRctdl5v
g7VjkRqgiPM3dxnkPFh7jwzjFXOAm2DmQQXgY0IXMaLLrX0twLzv8Rxs+OwOoQZ0
cR2i35xOY/krBQCQqjdkZM6KCLVvniCe+0loYdM6xpkZ/L0aerOZN3RcFXnifNSM
KUZtn5+hEsmXvOZY87XX19PWmE+apbBiBXlQ93vpLqgSj5yiaKcVOe4mlEjJOgrq
P7bvk1Rq1+GWvJR5WgqkzIc5SzHqr38cTkardgNaBeuPqGbwTS2teIdoc2/0BgbJ
o4ZJHu5NC7RvvpM7T4yfCn/+HtNJgTKgUBtdQmAUg7+27FocQsYkQ8YvrCnw6sSq
PP6l5zma0NT0xeiKbpXQ4FSl3ayOwoIbzN8a/N2L86TMznDXHCZuqZELQWof1m/o
eAT8YhFE6u68jYhI65K69uxtjdgkRU9TkK61v02/T5JLk6tzXwkrHAsu9sv4xGDM
j/4+y8XwGNZyGKnbe96V8b5gJg7DwEpThWMFFfcpRTQq0lGYoOmE4RrKJ0CafDV1
RxXrOkSRhtkXau1Q8yJL5kfbAQSSE2Co/KNj11FVmgxsfJlOfiEpNEqUsQfmjLiZ
Bq/zzTp6a1WF5AIoyTb1Le1S+hhtQSa7PdXeSr6eh9HviMUafy7resr5zLXLfyv4
TW6X6Y+Yi3/F/9HmBr90XRrfhSzvd2ksGeBSYqvceTCQWge/1E/79Y7X+iQxHRld
YM0FZm8JzQIa3BOBWboKmVKS66ScOcfveZ96by88PzH8OJ/Q3ali88fZ29nEm3Nd
ofv4pjPzGXB4BrGtDHFyF2nTGcVHzo4Qa4fZqkOawFkrw8ShK2oX3LNZms8VsOnz
cJtXgBCk3YQX/3qfCu1/V/wG6oqiK1wrNWsUWx0TAMK3e7alG68lNbwqtkzW2KFI
xwNe1hlcr5Xs/jqPsn2oNFD+Cp70aMizU75naQ1TmbT+zbuQLkLSAeoBceTMkbvZ
fW4N6evKJXDanrUxYuwRHYtHPyhQP3k14brZtbqCN+sQQkWY5hvKqHD1WbPj+Osb
MtBGuQ39E5UbyvYmV2Fj56mCWvrb0NZuUG5wEYkkY38j+u2riREHcRhOGRPnqm2B
5Ac96kPRhY0CAgczEo0D/gIAMa7ixK1gd3PMzWzUsF1Tn1ggfDGhLq9RBDbjoRDU
Oen9STOjjHO7Yg8llh7Aka4bD1ECLogIx/vPwmFroOQ5jH22mEZ10ADopiX4HufO
IEiDb2aEwKwbhwR+Opa99pmB/u2StFDfspefWOej5TCzEzo8ICQU7hNuD5loojeN
Z5E7VVXAfO46d0HLgGuOdEThS+EBiPg6XkRf6rc6jOFhI1bJ1iyLmAaUTpfdYwld
5gtoNHCWsJZDR74nGtjq5LAQj8jhww2TrwAlwKfgjlYLl6I5Mu8I94jNvJ1T9KtS
ATNMS2YVFaDmV0JsbE48DGFK3/Xk/apm9+dyBXC6+NuN5dlm3DbF81Gt+HTVbkJ5
irSQCW8erFFg37pYt4JJdtiGtlm+mHgC1LfytgWftpDjFIGM+1LZOjNL2PYPlol/
+NLQrfPC2KhjOX68S97cgAgyqzYPLzINCF+5g/O9sDhSnjfbOgATm0Uo82D+5ox+
C6acs35aThHZuvbVKA38tKqLXU5omLFBTRZBtkk3bx09BVTgddaY0dQEaLAEIqJq
H4J3bZZsein3LzZytcGzDez9sH1vzFm9PlXEiNjxWs8uJMej62fogkhTjo6N95Kb
TM5zAvaNoDTQbNloZJbG5A290a2EgMJfcuiRqPsziWkjZ0+AcA5qAc3XRfJi1GFK
P7zLLxwveoEGdK55VrmKMrWMn1xMUvXFK4RAthCOgbL3RTNTihFGgtMb33wmFTXD
zPrDayOInLYfyj3xVfrW32aTQWqiJVOFVf2t8cqXtgW+/4wq5+ohUa9HDgdL/l99
5rax5nh5bhFjYkF2as1xWEgtTXFP/lQJ8YpYhQOrLptq3OtXUkjficVSC140hnV2
ltEo34jjenGHsaXWtKMmEcdbrYgTP4uFEIAK37LYSfbZFJyVvr7+/8X6XIuqQ3Fe
4Foh64l+1A6JeXjJrTkZwhEjouNjAF1yvoLOp3GJSOiYokGjA4vIeO/axHVniol1
IPJsntxUn+3MuR3ZpbNQiet01I+wiwFgGEo7NCPayp6h6LApCamwZ/6u3J00uhSJ
m6MjpL6GansnNRJ633i3DoMDcoFwp0rvevYyZYEKf5Y+CpbiZZ+o0pVqaGtP7YbV
owYafJpGrMDIphNBMAIfxqjm02GZuVmyX0s/J+HPWpbKS3Oes6MX3Ipur/Y7TWQ1
nRV3ryvOckT4DfxNvIDgepAEeKUR6lqr7u0g38LFR3fAyjxDmVGXn68YkiaNK0ne
JXS+yMgfnmgGlgn2+7W7sKXg9jrsRsXxv2bKx1/9gj6hNm4TyVEO4w9pU53ly3Zx
dcDR1cZ/PvGfoYzdMPA9ARYZBwDY9+ldQYguLWdy2vTZmZchrh7O0AQPfwSBCbp9
iMMOwEKMbVr25GayIdJlyr+nFFEKJbCdROFjpVO2+YXrkZN4X1Jbgzj3QI1Pwwkz
zq6w+OhrbCxd2Cp3lDH/Gy6bp9oVHw8ZCxh6YQOQmNm8PwNxAMZHFLoMvYGKACVZ
YKlAIOODsCnu45JrBeesvNVlM5eoWkTaC4vlZMzCYsPwizl/p1Yv4KiItpxm/CCh
je1eM9pRu4XghrjOnpIwJzhqI6yhc2kMzl11O067N5aq20C9xiqXODrvbKP7j2hZ
zF0ONUcBXaQb8cT+iHz+BQPShTVseFOn49N2cbmEknvHGWNvL1PEa8KPh3gNtVjI
Wv8mgy0CAPCTm0nTs5xo9jAWMGJ5as1YJhYsxZHUMhO5TZ3A4Tmi4QH2sTtBFH0y
JAi7qRktlm2x7DXj71dLKTK2GIRuwGIgI7X/2kYuWySeL039hwfBac06kHNueUFY
a9vaVOAR+AJ73XyqCr9kg04NQkXYrdkF5EBI2PCrP1U+sPA8rrzmvKSX5OKVJryC
1giqg6Xt70I5hENxyvkU6EJCZDJAQCw4RHkxskoANQeuRdZyIEnD2kkX3F3j/L27
6YID0iVAjg7o5bEtO/TzyvSDmDc7Hf/wJHf16e5+HjiGiLgtS2CyI5txFMryQnFu
IEs7IKIiDAD55rlmc97boCAez/Ml2DRkFMYhizIQ/Y/GFmeNSYKFml+nTE+iE0j5
NDPiKZ5Heu2pmQxZXVwfa05v+ixT8nKfdFnIvuNLBHS07ZNRKHR8AI5VwnbYMvVk
ODOo4tySjSAEpb+l5d9w95hkVJL9eG+39HeDG807ofIh13muUKfiIO1ZI5m1DyvH
1E5+bppNn5qn7w8y1/iCWR3cn4a5ptR0UZfZA6t3S9uZua+AnZqRrr20B59ZHdqJ
/7BBtyNUdg+9fYPbFWLDf8unM3Uh6F38wFc+tx+1cBlKj92zVlAKnc7pQlFj1ufd
OI89BhWfdwGFFdrTB0/x2VBqKMX7MOB/5AWpZDQ9OK1ZN+3+/h6Jpv1VHjgfzrAf
QsFl/lHuOZGRiiUAWtPn8H9u0esJDbHqjQg5ckvB2zfcNR36yLHEHdFlXqY3IRQw
T+GXCqV2r5x4xcsaCyOc/lg8KYVRZ5k5si/VCl5LzQwlLozfo6vwrlB+S63p0xEt
hou7keGRYgWsIqwPNIRmRQ9J92Cg3WJEIwAHu8i2Rmg7nS/18Ae9ipiifwEOLVjw
KN3fy8D9VKYccDOybBYJiJujTDx79Pfg0QKxL8iqtXs04qNmb2LoIVMbfFGIghGI
O0SIDO/9mVMyJYMdQUScT48uMGV0qrBc5dhmWsKOSAagtu5wI+lLPHov0CqGy5mq
qXO4keLbcL7q9gAwg4mIlkudz6esi2n67+mffeHi9yg986t/JY2WW7zXKYZEt6nJ
Qt5aC+6faNvK7lCroLwI52HA9I9k3ZfHJh+GMqfyC4JBMUC9jDxAumZkcMK0mnsw
ZZevzE/AJdzACTPhS1k35zcxscz7nMADkLoWURcVUGOiYjzYsKqiY3OFRScnpSjV
IpKEgd/Eoihl3oqcsJEZPMaxojt/59mljCfqcFWjtc8qSASlmcAyv0TsjM4qOry4
6MOk0xpEOHGH9ELpkVsqqwm7trYvumgF5/x6nWPorecxUNG0hGysOAuwZalnqqWb
7dYhDeMJ4HvKWmUwiv5JSjf0QTomWORAZy6KVvnFIvEvqRwWxpoqFeWFNOy22hjm
Duu8xzteQ4C9Tcg/BnzuAT0WwAUeCslnnNixIMPdKNJlVzt49DK5jLnqnt4++sgx
EO33mOG304byexGQ/YMaNYF/s+gydSOuADkhFMrNEyz9tX7SE3YH/PTG2YVhN2Bw
EL5MY+V3vLiBk4WJYvAAggYtNy6HDH416Au33i4a3HxzsMIByPihvhytC0YliER0
CV63h3RGNnApnW89Hbkjb6EVRxRpEMNKzqIkFNexwsKMXeawG9rlQ+m0xFmYJ87p
cfYmS2eYs6iHaR2VfYhcyVoogOQ7F1dNyUIxnIDrKthKu8AaXmEiS+4Iy2zer6xS
YfR2KsumPCN/sSa4clK+aP0Nd2RpWG4sNB6F5oa8Unmdq/6BxLunUWKi7lX4BIh3
3gU2SM/HMDRR/lcdVRgv/Mg8vViYAmnH/5DClw0rJSp+vx+jXzPsX/HEL1TCDGDB
HJdePnpV3psPW0EW4qTTcWW+6KHsyM5Vs/ZlXVZ+8+EdXZwdvEnngxsYX4LNruHX
O5xPWmxhXPk7ScMu7d67tgYf54AyfT/n881d6WC7yzK8VBfOoWHLgdqVCIMpzBGX
+8EMJ79uznyCyLEJlc6EBlkhjiE9wEMKDk/Gb1p6Y7WoxkPLmLi5SQPMd9zrGk8Q
GfveF4XXwXsVg8n+cyi6uQ/4/AH9hBuYxDKUP9mMuyWbPWctf+UUam+vzVriQprs
/S9lT2L50TqK5fa9mrbVMbj/XvSqLDgiUMjkozgBaS5wIg6wbDzn1Zy8w7NVI5WM
GSvmLjvtsfNmNAdSE3LBAyW46odMWcojxdMKXQivoi5Zr/WWalp4sEqkVdFXc57j
DONaRUu774PBJkE+TJz5XuwEq6QG6j3qAW7PJeSNSyhk4pCnW17hahq4nsu1DmJ1
+tBde12Z/QV0n8K4J/AqxDnaIp/Iqb/V3ZtacOO0pjHdOQJbNXJfpKmVH8120oAC
8KBL0+xXZadaLJN/+Ps9beXm03KL5fXwUuM/vabhMAmaX1kZ1NLksmByGME4R9d+
JCGmHRsOoy7p1Y61W4T0v0WhURiT0iaI0XAwEf9pgEunQLb6TqTnjxPDSJ04HCaS
dr8yIH2/h8K5ZUeCOt8G2aGex3Ik1HfSA7suniWB2cCdBuGDjnFhfO01cNE43q5c
DV9+6Qeq4MNJZctvTUWCz8SOLzC908QQS3ZNcX7jsAflkuVuEc7o/ma6bdG0uZeQ
XkGuy1DU4mW2K4G8bYOX38yJybxKCDVLF+lG3fHD5i54glXE5wMaRyyLZNRNup4h
dy7zvNcKePnfKIGy7eMsOH4NksTB6xX+gN4W65VinErX875s076HAZDqsvUDiWlY
eioPXIWH+pnC5/9FfOohjnTnYWklgdjwvy3K1T7t5IKHhjjvJd/KhT0m6XDZqBLT
Z99tzYD/hGTcuFdfLGWPF8jaJqQW+pddtT2/qP9EJt5wGQMDY+OY5QmqNwefIm34
/EyNxxEFYl0lUIghcZXllPKIB5dkRaQWm8v3VefRQEvs0guS8FPo9KsmPs7XNA6v
Wx8grCJ+48QogV12G3CiBsVDHEhX4yvh7eFHTG58oDxNpAgPMdvCdYkv8OjFPPtG
+gEZLdB5ZTdM+FwqMlbj2HmMZdUtnZf+G/sZxM29wmbKVSaZ8YgW5QxU80U4XN8m
zYggbI4Xw8GesDnlD0L1p583rOH+Vk+tByUr0AmyttCYrmd3CiH39q8oYXVqdUJr
SZBYlXP9PdS2sFfwz7MCtAfTWm6utPGLwdxzmm/9y2x9zrwSnyfpdzyXlfjVXrpa
fq9DZVa4CsH7KlM4zdSoG5K9Eg3NzpISiulI3AL8UbBdHb3Hza+nsZF6OUydRodr
2kiVcpAXkwOltYMqwSBhRx+iVsMQ8ai2Jw+dktz5zewHJti2FMQvxt636emnbHPj
N79YfEJeSOSPHBz1zjTnfIOx/mTrKMoT8uYxCzeBO+BFTBga0+UCf/7D3hKqdEEI
rloHi6rnVPRK07fxFZaUTJXg7fE1LrvdnWae1M7S25W5L9Bx5MeqDlz5m9CAFzdk
AqWYqQH5dDKdBCcw+pxM6hDm8dOrb2tA759IvYPlsmUjt/VIaAa6CnEGBbQQG8tp
32o3jl8FEFWdNP3Ai50g2fZyUuaqLjNIJvlCJU7NxPtBdUINbC9IhUt8UOpvb2fM
my3ngsiJkE4xXIQPz0NtK8WK2N6Qj42EJSTDEzgj5YBKXFfU4YEf7XQD7sLxCBM9
wrgj/m5m9Xf8rP+b1MiXuk4sVl4HjZOT5vmconwEmIbdOL3UPbc/my8F+wv1bzWV
l76gx5jGGeinsW/iVHeIwn3WUEbk9dunygvfOD8H3pjO42G0iDk9NqPh6KvL6ANE
SpFp0qd+8mDBwusfUH4HY5zzN9JGJxNm6EbdmSN4ONjq5N0SxDu84JQ58mgztaSI
PelnKA3+NbU1YLHLRqcpWZ3qdCL9VD+xQ1mGntl8ZWcoCjx4wxXfcvkXnS9oC9Qi
HcbRmpCHSlTnQtdGoYKd2JhXxkgR6Uowaxw2skE1sN+MdlL15XG/dfcmbKWfLjZE
dK9qAyDULglkkwTeBP4+V6hXg8cGCsbf721dhvOFnffXxalcPhcR4K9rpXvnS7P8
TW6bAfaNFCwgwoj2u0xu5wCYmyvo611OklMZfjogwaQTbEUUgs5pPDIwXe30NrVF
XF52ElzNI7j+1cSUj9be/Pj85iZp+xmM4ixvVpt0qNFzMa5JmKwYxK3d5Wsd+0Wg
r9A7enqRZ8CWr5KDylq9bNy2QTXxBZzVU/+zA2adTlhBacUG9AEzpTFSJqjbcdL7
I3lRrsFEmqMw5VwNOfZiMeqdUs6y1oTADpkkMvIJV0Id+j0VnAMGjYXk2TNp6ibP
UxRIIjUgstXrODuqceVUmFQkmMiGbfdtJDCxv9/daT6x9BrqaZVGQ657q9sjzjES
MWGdpjjDRaxeD9Db9JYGWDNSZ+q9LVynS+Rpkad1Pt6wy5QEurm8+pQZKajKFmd4
dYyifr+VLBNfhfusVRvw8JQ6Q4P/6QrLgzgOIxZ+/V4uFGDEfpk7QdZr1qr3YEmX
XzSfoE0duPM4EoifZn5BtDpVsxzD/7nId8ziYA4lbxrV9o922B+pBSORzapD25ij
O1BV6mB0of+o/lVa9z99UlCakMx9J5FuFWpAEPCv8pzxneH8K8W8bL9n9uiDfC7p
h9oV+UYYtM1PDErfrA7uBhGg9LTnACb6xBdQ5G37nWYyH0fJIwlbwnCyOtnnKz/k
HJKng1xCdjlR16uif9ILpiL/78enslQjs5EdTs7jODvuOQTEKxRJaLBx9hB4Frqp
cVXmtXm6BnDrGeHUainwQ+ap8DlbBNzIKidJd09Fr7cd9TXQ5jHgeR5vFNtBhx5p
zvg7MNnuBxaLsqY/N/Tl8US7DyKWQeRulQ6NUCoArm/crUNhTfi9upaZSZ+dmSGp
vUpqmZ7efgnVTnfPBZLyTejN2vXV/U8BHWDuYJOonaQxTeL1Lr8LSiihwmfptPOY
c/IU0Yn5kpmeHatK4BQ2ah3UEddwlHJPpJIcoGuEZ2bylVDT0fRFDcoYPk4D6e3L
edu4QwffFTXVhN/1O1CL+sAzJct6zyB+wXCn7ad1KqWa/ESI7kl3NTzEOwgCAzBd
AeepXBqBYComzNn4gWlhlE3hkjlq3N69ecX5l5IyxB+cFsr7BmW5R+b9gmEGaPpM
8ffV7J2oSpXuty6uchqsAOP0mguRrT20K2l7uBDF+8TEzF0otG+G/mKmoNehgvwz
U+zxZHR2/YyDe08YfCnSrM70KpsoArmO6YEjyfUBPgZ08JjYl6p+i2lbt1e0RVAC
wF5iWpvqUaleiS8cHL+xqLwQlEwAnvF1nKJbmMYMcbKV0Z3McJmRppbPtugAPhd6
6m67Sqt/aKUaUW7kGhVhG8x9DWVCgzUJtB1xZWkxsk3Imt5+ExJQEdTIzKRswimm
FOvppkQBresImXTmxf3O742FICxhTO+IAj9zG4hcxQklcqE84kqSj9TEuo96X92F
RoUFX8rjBB5xAXHaehTYF9Cn+lPsyeIGz/yDUd0198wRKchU2Vf0gl8TYcNTlKAT
+HfnNvMAGi8W0D7dAN1dtetl+PpD5gNDjQpCOZwcvLnCZRqyfANd3o5nd+k9rFlP
ybInr5TW5/31R4Ju0voLzRoDe3Ziwze7+GttkXV47BzWt2hgzghSCZcRT2h+rAQ+
AafMg6CppWrycn8HMWvUJUSO0Tto9F7lU0rtdpR3hHr+gkTa9wk+GB5K7G3ka0SQ
dsL1Ovwz9XC4qf+DbE43vwtCQXk53UuI5hFk4JS0VA9HY4xHDQz6cNPZwSd4fLpq
fNe31D+fQox+Zr2ByUCuKhKHLUS2nzbb8hmQjjnMdugS3M/DoX5f6bpvjuhSpge5
GiXszi5UriSsCZMa3p0LZ8JEEj8hUHmCY9jBpAWgx64ZlCcehxUCC+6sbTxfJTx6
ZWAV3AQRgf94OD9BglnNTsPG/YRxRVIYaxI9SeE454hChFpSKGe1FI9AGAIR7ZNy
2tpXvZbV/kEeFEnRReKkplaVPfDTxxkmT61eiL+Ws1GdCoTj7Hovfafd63NxVHXE
2pYrcjxj+4IPuDk5BJEdPX5E3b5kLhjkBnEdN26IwbIQFiUb6g/DNxinSc1e0yyz
tQF54HgVtu9YTDJThMJiLAct4xDVWkZ8nq+jbsQzAZ+C5NLLg0nSikw4iBHr2j9y
6VLLdHkVK0elPM1UnGBy+CUO7qBgtOtx01LfGaPYv8k0p20ePyzC/Oozdtkp5NDK
D0Nz+hcyohSEWXfPMgkNOS7gVF5Uc2k3zoPrXfO/dlL6iG+CPXpvHRFxcCEBhBA8
eBWFO0udybOr4yaqLyR52HbK0K4G2GPV+vQ8k3qrdVrbKSYfxYAx8p8hJ8V/QH8q
VTD8F5xlTjvI4qpflkg0IXPBjKLHVa76qtdJB0nwlZqbR71iWSnbu+8U8mg5c7nF
AwS1Ap3vM0CmrR2ZksBWcXcPXa8ddKHtp5F3PqYkFh2smU+A1RNinhWeLYsUZGjt
fN62nGT/kiPgzGuV9eikSzNHKBtTTDfFWhf7IwqJmQfd833fMzmM467oJeKudHol
cwEY0em8iwR9c1BC14CvmyitRLsxnIa6ybZ1si+A6//gH6QHk5i3vSxGdR0iMXch
g3irh8qAzXjkYGiLrCqV6U4FXgOCk0Z4aq8p47xYuoCTlDYWWgrblj8JFD+9CxD9
Cc0kJ8u7EQfcsKgFy4qtnGTdp9Nx493Z4r8KVjDsM8wCYUrQon27XfVI5DLhBvpx
EWN56nNZ5Ow7YhcFEvNC34PvrkJshIZZ7d7vtuJh88JqqRcGFUhCELdFCx/T67Ta
8yK4ghldReK7sgf3rgCPOJPowigVZsbeP3j0C0das7boBVYtJ6MSJaHYWV4SooSW
kS8Fo49fh6dEYiDwGWGmwCmqJyqWpFBie4/AYz/fvtwD14nQFB9axvNNGBnU9C/L
phmCQdWLG2AjZVQRh531BJ+AgCJZt3B3fJ7DwClioKIv3rcVNfbSOikFUGF+e+gc
n7oP78LwHDlJ8QeOxM0uTfNxVp/sPhp4SnDtMv60LWuT1q8F1qL5M98YSyMTJmlH
4UR2GBhdiw35Y39llUcudG6Hq6thT+TrdkEvnQOCbGNWUQ+9h8And8IQWU+VL0V4
slgMAEPZHGXqyvZU7aZf87bJ5/4inUjrPdyuZASc3uCqALSfXjS1dmdqQxlTIORg
7X1+dJA5LBxZnEd8bws3Ssjn3A7PCzCppR+8/riaaJaujbrGo+O8VkdLTS4IoKth
PUb64FdcIOIUWodK/93sSXNnLgIuhdaYutL7K9vReiMx3VpLYGN5uXp/RME5z6ZZ
D69izXb+Mjxf6ejoes9qAMvZCaduob1SIMofQxh+M8Bwqj0hTWXi8pOwcyHxaX7X
GCLPmRiLUgBi9JLZ/pXDTgG2OJtcCjcNnCsxxGJOgkiM9X4PfsxDVUQjIdS+0H8c
UNsiYo1LC4eF0uhLG9RNFxC5eGmXTmAWZ/dWZaOmv6ZXlfUWAzaQysg2ZrxmfEir
FqVHT4RMUKHdEBusb4hT+cTLxgUbMuhqijOUTe1DGBC5IDXzlvJwbL0vyyLnvtoR
CbdTbuJo3otjW+5H+W23bA6KVgElGzS9tYf2xDl63DJAfJo5+vyhsq21oVY7WGKU
Oc/jEyyPY7Tpnzr1zBm6holsODcz7Ayzs+Dy62gsi10bLOuHbnfi/B++S/72FRGD
JZJ/zZRP5jiCV1XG+6cabKECjOYW+Yf0peNUPQ/ExX/PaDtUiA3SF+MsIorKz3/o
IxhGh+yU6QGl7CCbcgppdPvgLXz/tqxYy5LJqs3KdH2Ch4nXRg9J+QJ9G6VRUzFx
rPdPsSqhm3alLVQG4u0a+H2Ejfgg7PMo1j2DzEmJUe+43iU22i3tCkrzRrJsg6zn
vxBKYB0DWMSn0DKqXz7qZrNA82GTVXTFZXwdxQMJWs6p0RCUU1PTx5uYq0DXAgEA
vsRsa986+SOczB6KnP1srfGgyjoH1Vlh9ouj82NuB+1FQjVnJlmFxMoHutKTBaCR
sJCtPXv3FislISmq8+AQaqIH20huj6mSkFFi0/S2M7GGXeQ2IQ/lNahXGtecjzXE
szeR4JBMe+kywnl7BPetHFKAj7D/aGImnUrUT+HJ0k/iAV1fQHLmE7ac/LlLIJ5t
bSqnRiLyMC+ZsjJPNvzPgr8YEZrpTLkG7uLAH3g9As5qpqj+FGpVVoK4PWzB0et0
8VDpVGyv4COLMPWYvC++4foi2x/edUayg79hKwlSYXkBS4l3TpQt7S66WDY61Tlo
XbkcG30JL3p4WB7qqUTurz6Ct/LZ3uTO7qmS4ANWpWTz9g6fCDup9iSwBrWN65cm
lLW/cvsIgcCFPoFYXR/lW8mdXbvtt8rTC7qToE7pBfwX5ADgpxAOHUVKm3Ndh34a
DUVbiEf0TYDeeAEoH11WqeCOsxqFu9cb+oJUE/aW3RJp+d8dKmACyaasH8kaTLrN
I8KcI9ixVMGrytCKI2U6pc1KJv4rRpNxvtLWelGGwcy0vV3mZUwukqDhMgZx+aX6
QQhdGED9q68Kilf4aY/V7xFZT0WtaLOpd912HQS/1atO27L0ndPcZKOXp3TFY6jU
g5lpGXPUDePfR3JfppYQ1u4+M+AofZ306HhPgVambz8DTl4/X5l/t1krqnF7k60M
wmc6vWdB1VXJRFM9sBTNCcysLtLlk4z6q6Xqb1A8QMeGWrO1MfTi8HOrIrMNjb/Z
VGn5clnNbeCyJF3S02yrTvjSCf6nApJokoT5NEC8bozFLOCblWU6ikkG94GLuPTl
otuRUKJZ4encHxToS1VjqirebvYgU9tcjdW3meYqnQxe6A1kd26bFAxyNILSUJcw
p4ZCXp6ynzsLZ3zyGpbRWt7u52oolUDLqPTTXSZ3BpDFtaTILPVND3gAa4idnUV4
GLCKwAfgeGCrWbnJ6CPW1I4CU693MkReRCMBU66fxzI3IiGU0qS4m2JuUdWz+c28
5P5fQitJprz3f9K6loSsY8n0ApqMlg130nrDCeKJPDypI4FWBM1cbrV1voRWFc5P
po5ZlwUDC275x+kU2A7UuZarQAFxXzR9WqU3gHTpq2Rz+Cpq3AWiOXDsvXRl0Hij
N0Ra6P+e5e7emtukq8tLUkV4tL5KBLRWS3kuYwY+cROJF2lyfJdJU5RZOK3Bo4tw
GeFq/s4W8KcgOG791QCw3hmRaanUlJxyM5bMrDRftjs/EJl9Bv40zokN4cId69nl
P63RY6KLNRoCjzy7NcCOpjtfdqSzyAuV4Qy4w04OJTzPqlTje5+2cLhVAk2ypzvN
W/KzVOnmZ7aDtqQzZTHlUNDqA9WvAzyaupo9CgQOtYNzzKunwnK2AL/6qChwFezF
Cguhp0VSDSikdIVQOrgX/LoYYHLA8jW6yJAxaohcIT5oGVUkr3Dnw85sXp5UaPTb
6+9cld8jbVswuUOvZs1jnktZloz9jPeQPXQuvq9whYN7pI58/ytCdygvh5JbKryq
F0+k2+tu+fOA4d7DImGZSw48ZwWx/j/dAvVrmIOuaF9sdGnrEtI9N28Gi2lxQeml
FP95Js3FisPzpPmivuIvDvEbGfIaj2m13rjgFD0pTDz+Idzyv5xIWIkS2h71NdmA
Pm8Hj74k3j7vnIi+LhvDIMdP/2E7cMenWGzm++10jbbmm7Ywiv+A1/Lg1B/l+NIA
oi1gNO1cgVcH5My3nwbNQXLO0gFqRXH5ZTzniVZBV3Zk4jf3bIZ6uIWKPp8UXjtF
giG08kWc2qY5ndV62lYYC1/VC8dIC1zID8slf26Z/3KTd/lGIofSy01ll/b0/7wY
N+/fLA+E675GNnSFZC7HKMoDdVPEGLI0de+jTqLYAaZhM0phpbgW1cdpkj5+M0Vs
vKgFWgsGXsV/jubISzoodrH3Ft260fmFVbkXGnpqscO+m5LfXFKATXKCQkq72cu6
cQTO5Nhpg8sxZAFXMFO/HZMzuRoC3DfAZnCaHyqboUJNDfCyJNdTXREfnJtcOvS1
E0fVH+afCZp5TDr8sAFOYk5J6hKVM+PvPMvH/MQcz+AQia7ctP76mKE7Isg8Ns9s
TFDhpUsLdPv5j835lxU6K3XfJk0oD7YvBfUQ8vipSTbpi0Sc5jkgh52kPHH+pfpN
qyFKOifQjZVW49OlECCFf3eU+ohN4hw3+poXkOeuIBKkxRHmCBurEaAArlOArfRF
1pKbmRWSTPzu9I4kibmSz2ANrpYxT5K4xYhqbushcQR+bdu56QxkGCbkPLpynTxy
8TRNrbXbOXXa7mM4rLomqQU2bJd4eNfJwn8nH7kxdfiXGVlTf9pR29si2UllUY/h
vlm6VswCkk6HRiOX53zTt05g8OyLFltzzNKmaYUnYUsGounNWD5CDIp9VC+nX9qW
w+zmxK8Fxk4L22nDgItrlW7GepUt0qapYu7c4RHBp8nsB4g6FdwlTiFOfoQaWHqW
yF4xBrDpONL/KhEB3hHQCsfIL9Dh4WZZljQZ2Wcr1GN03wSJJrRJyNb5RV/lJxW6
A030s+6LYYt7Y1fFgUdBKQkaNc0v+/rb7RKKYi21TdEEWbT6/qHsSqVKH79qh8cS
296mfHvtUFo5yjoL8hnsBHmTFri22sv3cVTzlI4kvH/OmC2TguEtNkR2s5N6Xace
VFXV+vubK8M8Yt1qZzc9GI6hFSoBfhTrm51sWRwBIzar0BXpX/e1lsquvOJRmtA0
tjV+KBe/QFR2SI2YIowgsITwJj4b13462ta8TdiDt+Mq0nXFmjW3MutPMxBCN3Wv
Xks8t52GiO5AmYzZVq9mOUBfeC2LsDPSoAEPpN3bv6uhO02pZHc7ql+xGsXTZEKB
gfrDLQyDZ8EZ4XsaKfwmSaJZOnJGsE09fwE03VDybMuXzlqEq6lAH6E0To+yBQid
KBDwfU3Asa6lr37BS/mrfbjYVurwhDdaZE1LnN0HAHcJrfL7DqH6whNrvYLkMkTc
WBrOcHPD92NxFu5CJI7RqipW4PucTth6jT96gfXeSosO/181w+AprmGYEd9TIG8b
PKBmr6Q6C+MOKzgCoQCTmKt28iXMQzZPuJFNYag9ysfjYb90ynhfltIuw9th3/bV
41TYrCqVUeTBsQ8CVHzH7dcvp2hHqLQqSOob5tTPm42ajOx7zH5NJTuwLEbOcpcn
pRSwFeD+1BomtyofPkQ/66vNgm4pDhDyPU8xKujFUu8H/f9YKvvJ7VKkhoRFeCwJ
pkXcgbM6Nnkz3f8dkMl8gWWv/hUJhXhxBas0Zmk5xXwtm84JRkEK56+WhA68VKDx
/AjZUaNhqA81PFoFT/DCF2l+Xr/AFYMUCNJbUul6QUkJF4EvEqoi5EzEwo8MTj0i
Hvn1WdXHIzAJpS8bJQ4w6H0j3SCCAb2P89BXfVY+WFHaJCZLWZx2lx0TTMe3eNqW
AJ7xlKIb3uhaUB/irE7an/O3UE5SYh61L5/sxk4ytXdMpcul3XXDJ+w/CtSwDdr1
6BASe5+898SjzKvjDSBaIGPzuv++5F7g+zr3C4oZJL3UvrPF1XMBw1fH62WKnpKi
XbV5ncRSp8fLAYyxp/9bW4b5FYwruJiUxa16d39/3LB9Y1Tli5P0qxF79oNv10FJ
TZAGU02oyV/mCeKokTlWde/s39rG2R4YeUwh5VxuIuwFphP1D7MRIPIrJ4lhx3Mm
o+lsf6PK9mwILr+Ea+h5Y2EkgCxCMPLF8ZdPNBA3ZxyDt+HM8ag+va0SKot5e7o7
W/AChduvFNY5SOBjleWxOToSHAmmVZsLEDU8GEer0pD+bpwvtc/kxiu7fqKgb0Fr
fNBUJZ6QQbpR4kT3bWSHUdOaHLL+H3vECLbNAwuHEAhIEz+33V0p2nCH3zdOmH8G
iQjGaNPHU78LP4owp3N5vkv7F89fw1V5no2f+xUwDgZroEkGg6J8mEldz7cLw8wP
5H0hj1J7m4ZscGNyTb3ek5K+N1UKG0QjItU3M9Jqx0CJ28B+I3NBhpwJdfRwailH
8YGUQyZ1BQ421QV4WQstdrSZKn0DpNTOC0aMlZHsvZd4CXn2rKDyt58kAb6w+fEi
tmNMmJy7KI+kgzDTnM8uBCcD77V+cdtyZRW3pEXNQjhicpCtzKezcmdzGzNKwGvi
0cF0PX+GTvhQafNPcRIZ3pswL4DJNlGkso1PfOJaZjk1uCjAx5Tkz+vOXJa+v3Pv
l/UvAdtlXo5dwUT3In8Hn60WEdkGAP7bHC/EncMSvTqVS1i+WMfwxGzxVVdUQKi1
Q4rQLtAWuXroF27+Y15T/Pj63J7PBKQGrGvQ9QuNY0SjAY38DfoGA8vhcl7tyzql
jPvVFmHQgbXIC9mtOVcupJOj2yn+Mkx4FPpQg+Pfka6PW5BOOGenSt0Rx8QrBaxn
/T43d6UChSYoFQ5ipSO3B7wF6gmUk+57HkGRnZmZskQpAl6Q/xMkS+lW1gFI8m4I
yJ5ydXemOhfe9QObapsF6bYlT44ov1TsxN4Dqkbta1CN40sH5ziTgOUWeq6OA+43
ZS8C25on+P8BJ0SRZ7+N2qnLMGowPeLECtYg3aZlDrK1URlqUYIwn3K6nThqud7f
3ku9t91nGScuaMzHtyvNGXUJncQJYzczSGekmER0xUTz0UYz+nSMrh3FmasKW2oW
T9sZjIke5vD9MxDQ9J+Vp6KnKic722+0lRWeIvAtUnvy/RLVmzXb+7a5B1hWManB
//HYAZee6SeZEzA1qkdckWi+f8fYXStZ8NexB3zwKZ96Jdp+xx2O2DIExl9fDiJ4
QWPg/BfR/4T9+09C2hjmFa1/MZ64jkxPbrQZ5+2obqB9sVppXawocf/w8QA6kHUZ
x+uBeq2Pq39+Q+QN5lsfDi4sK0ZXq3lPk5pzgs6JQ/QTKUvhHW4Kx9AoPa9DIJXo
28pUqO5fBbFfTM8WRRLnWwgH1vUqlIN7ejpaYzBT+RAyV5YiR7S4iCHU2eMTScUu
vKEFQ5cFT6zKHPg42MqJ6tqlTNmDMBDYWRZ/co4ePpJRpLg+Fln210sF7QdaMBVH
SG702R5LVhi1z/DeaTAU65IzXTgY9eUOml+kLA5F8axtCrp2JIV8OMLiKoVT0Xja
/2G2GdvacaxxjvcpbJ8Q1s38SpkxBBr8aciECPcxwrAzjLMF/al/nWgfZOgbq8AF
XEB/P3E+n3+jqiWReA+GP5900p7SFaUMMUFvMPGo2m/B3/TV5DV73DVCthpvHa8+
DN/c4UIZUCRedS8C0CaS1k97nrZZmADOApjrOK2KMFHWUxKWhu8W4EihOiQC9yJT
cnWGetui8EudesQi3309sacqSizTRsSH6eohfWrgTxvLuv0Jiav8Aou5Taaa/naa
qnr490dOWxgxjlywqaXsLYwGOutNiL7YOmJUw/pkBbw2amjVREb2cncl8V39oMMY
LP6vFgq2Ui9C0MK3XxWocSEBe9Omnt+ARJYW1tQmOxxLdgWgsjgrCkjO+Xv34sP0
zEm7/SGNv94qBQuSQTAFaGVJ4dwtlrBKIa07GPIEXc7sWMFf3ajFNGCaJPrOy1G4
VvfgVun1cUu3/019kqcZ59/mGmm1LrvJAiTUoDSYIoA3zlo5TcOTMmVJ+RewAX8U
m+GHHFQk7Gohtq/RLCJJPN4c/nfHv6xTzfXpDWDhPK4tM7tEph6hZs7HPl716lL6
WGxHC2KF+FrFmfn2thDzIUiO1ZikhKm0ayJo52RlSYIc+W8a9tjJ7NlXor4nY1ij
pCmEO5NACzOjNuLobPPYsTr2rD4RM6REGayq9mRVosOoOXXJnuEL/fMi0vdqU+G4
Lpk4rgtgGvW6HIM+Tl+7gsPfe8aC5kix86JCC4IXrttlReKyE2Nqpt84nwO+Xxj+
oJ+8G59BCFaZsKoT4yWGF68jWm7Modcxn2e3ncJjTH9qMghiBTf0Ux8Rc3KIHClu
X9XQ6La/dSmWGKIeXetjLb6ytOFdFP71vKWtHpbc0kCl+jwTbEL+9NgFAHqCfO5q
3u0t8t/I+qlgLUZ+wIYsUmNZPYphfxtvEuoQAAaqvD1u6iHBCyjA9YJz6X+sXhs7
49Qet8yPe8lv6o7tFDgyz2mgIPv0UJD8kooX7xoR670ISVWe+Tmhrjdok5SoZjtU
0FQVDuJ4YSnVohvfcS0V7jdNtdl8DWgWWMq0Ss04eMb/o51GmBqLZW7SEgPtOpHe
6FirYpw1RA49TLco2mvNbKffFNzqPhRmx3Qa7kx5GNO+VDlMrtIVauCvu32TRi0y
+lSNZeDP+FDmUhO3CYsEO3HpF1FM5Yvk6iVQzC4nJw1x/vFneyxfWah67qjnwYRp
/n4suxROYwo9WvHovY8PmxoyGl5nRuhonmS7zpAgJfuPm23itPxBLNlaxqMZGxL8
+KEVxlMYwgv1HlqQTGmCDHmCYdr/tfeqYuXf37vK7cCARtyBjQalMZHPhm1oX/UA
cTodNfLmsg7GkN5aWlALoRHgU1my9KqugWVjE9CXiyTKJShAWBMJcRdoFlYbhvFY
69EzusCvR4cXOiqnZp77i4ILZoyGTKgOJRzM4+pfqQocDmGRoyMGtKMarEw/TumU
NUsYhX0vTTg42oW69BcmsFR2u8ieYW7id7HqnZ7TFV40ltQwaeNPl80MkPYWe1Ym
L1Q4MAvGxa5RMRkdGksjWyqOyugJdX5HHdZ6dr31Mim7+4XcX28NLxSMwK7tkoxO
w+/BMQVlLcCqCc68F2xeGpalTsdD4RKkIZvOPS7CjnbC9CBmSqQsb4/XBF7yr5SD
53jVhKDNvtDRc+R2vjbL+4p9O/mSiKfSFmN3kV3fCxsT/XBIo0yfuoZ6yB5bU9kg
EqCQ9VWwSd3TaOhNbNqiT2LshGf3qxNXhCM3OwiwSL0JvyDlFwC5o8Ljzv4MLETX
1R0WaNcNlzstAcD/2XIGR5r9Ji2y5wQBP1yew1QK5y+x93hpM2pX65Q7K2eErSRE
XI+xkP0gI40JOS5PqIjjkW5LHGkVoS+CbOW8JNj/qHRDF2DZo/8j4D5kcPo8VnkV
wkl8M1T5KQgE1Mc1dHMTW2qX88+G+6GpdLoi0qSQ1jRsH5HNQn38qSo7t+8aFJpF
+Xb/Rf/dkVbgP5CiplmjeTKTLLNZxzFrQnS1d01LoTDjxDfCWxU+rgU7UClqqfHW
A1ZsTkzyXfjF4J0+D1D2oTShu08afBMGVBj9ufZxsDQdWXeG3G7dK/+tsCz0Dj9L
+KDNXWiG8EJWrKFSlKEINGReanY9CM1F4TMXdp7RdyYpfDVugTCCMRuhtbt7JbpH
AAGDRt+RKPWIw6wW3mb4yWNb8vpbFuyP+g3sRvw8Vcg5YcLSoVTNc8NWt87JBQQ4
oU09EkNt83ITBq+0ZS9z6IxRVl5Gy/vBrM/un4Rg6cBO+Px9U6kCu5PnI3+pxyY/
CU1Vv6HETcpXjNhZ1v+AYQOzffnllM92vVZQeHcpiLuz1jQIRzBbcYPkWKdhNElc
W0tY2u7MnfB0m7GpiWGniV4qzkKLAYHSee98UbIdNGl/vjRBokMwhQ1Cm7hNEo21
I7XWOuGqyzgZC5zIf67JBL0Yv/28QNkfSVmlxdQ0UbysH14raoCpWY4hCLv/DR0y
Ps/BEVOKpCJi3CeQsERn3JJFRBI1wuFoBeCL5xq8e3nVzf6oIUIlJjjTt2Ljq+Kx
CgCKBuZjSKWBkjhQQEUtL81IGQ+JVeBizQ/43sO9/rA6W3IG/4ZvzCSBvaIwUZbG
QbcVo5NoVFzjrH0/XIE6Rh5LuwCevzN/CvlnDde0z1imLnp4IqXANrVdSG7IWZZP
8eV9TPNTpJSeY6SHZzEI0q+WUd06/KqEIMeEjjjve0tP5m/LCkYVqznBBtldsfIM
utZHH06VhhiUwoCubkszR/NlusBvQwDhnEgb4iJJ1J774mJbJbzQ3ezyn5KK1Gaj
LbKNHFJMY1nHd1N636irkuvgUIeWYVVylrw8jo77ds/x12Ib6h6gKqeVILfglzqM
utWGI3+xWJPwtZdkUAuEzbBjl2W/OcHqVFIOSkCFmD34ON9V9+I17IR5nJLHmcy3
D7f1qBgP5ba0bQedVxonnYsdjWAzLPAUTxxru5M8rydzBeQSfTHDcWC1paJu3+nd
oUZ4FVUt5hCtwHOzxJNwl22XPxU+hipTPCOlJWXhmS3eKMGniNI1loxH39iinO9x
ojy0B8QwkA4c5/bKVMj3eaZ541RJBLDrg5KFuBieNhCLArfVNdnQ8L3uOimYLPG9
Ht4Ex6fzAB7OArTZ5FPu6HJD3/bZPaYBXQTNOvBmQ8ELdYEVqIOS02g68Aae29Ra
xlEQ1Ru8FaSY+jgu3EhnwvG8sIcS3FV9cyXadxMaCZ30MmQ1uET2G5nnticmRngQ
DqMG3lZpGBGnGAAEu6vFxf173KBVAMHsS6m0Zv9t9hvXTu9/rP+KmtN0IeitD+bN
cQ2gbKMzXfctcGtwFpe943safa/Tmg5Eq8WoPjLf5exzTNH9KiinAPE6hKWic4hb
UxRaQDLwgK+/EyC/avKPjFpnv5FC1yHdgde0awIBo25VeUBWrwu95/HRMm94DUTf
SuV/wR08Z29L26oVWbUm2qEdrtbeOUA+40dmL68bvRGBaQBN7CxSGKiVvuzu/+PB
hDZsF5Q1irHTFcai04orXJNR9TxIEoEUeSbNPMSJyBHXCEowUZ+d4Sx2RDGiAYZx
hAqdS8TKNNZk2Od78VMzpzq32XeaXLq5o1bvRKmWP1aefea3/GzvY2e4b50YDal4
u16KLtHmDYNXrifeXSEe9FmXtbktsR44pLCGPhbAr7DNrqLwtSjWxXK8/9AKvF14
qeanMOpfr6EFMsxFFxltlNeZRyFX+bkWGS6YLhai6nnetkqw+vKPxF11EjRJEYPr
a1E0KVYdJ9dXxzOYeTrt/qPZGoGsiE6O/cX+eCVEt7cTkMq3iQqYsgTqDW2GOD9C
/ooBItnc0Rw+EVDPPme3//GlA32ldPixSDnA+vsW23AYj/GzIx1SdRdkHg/sKHx2
A9FZYOV6lJFw7ZZ7Taaf4XIJViVlH3J3rFfW+DWnw2cCkSdvbaBg5APewjFJ1XAl
TPFAosHQop+M9/NCEBIDG2fiMsbhgSpPB2NaMq6F7PKuiKBP+zTSeL7Jq31Diofv
Vu6aX+UFDVUN+u7SC/5jM89DLtRFDUe133K+16S9sXcsb5wnDfYhc3CnxmFC9URU
r41KnCQZec1yDDR1GGZVr/q4YkHRgFuZtBC/FKjkCQmdUFUD0K/3ItlKdBf7Zgbe
3xiIns1jOZb2hgUxQ9kxuY//N9gdra+rkqgsTh3eFz1+MwTY+0uoDW/0ZLWun5KT
R/Uv8Txwe4UGN60iD42lxa4dhdA+dySSDwasNVmp5ZtHVtGJIup1LDY3F+V8LVhC
YYP6apHk8MtYvM/Tf4BMjcfJzL7dsZTXcAG9teq4E+utNFm5Vcg4BBWchUl9I0qU
89/KHnIpcBNirLLctXCMAt/BjBeATbS2XHs8KuONrhCO82/GFV7+FfsdMHIn/P7f
E53TTj4R+BRq5+EuOdH98FSxEXt5gs8Lzk+ukHWWivdwpfT01UWKI4N0alrI0r0v
uaW7S/11iZq9X9FQei7gaWGTtsdCQgYiSLulzHrsVb67CVpE66PIPz7ZSG0phnT4
qZpdnLQ6I0kV3VITYLgETgpUOCfx8vcf6CQFkacifzeB9ZvWNF4WXqYRYRROMsCs
wfY8DjCp1+OhaLvf9GWOXcuudTVVtLcmoKs7NYOnaciToEo371M9qVa4706qdRoh
1vJ7h7rEYi95LpOhSLyDqi8tYhNyBpMgghvVzP/v/VwZykjVI/bD490OZlCvReFa
cj/6pHcvImyH/g6EQD+rgyj6gi0M9DfB5JuKkYD+vnB5pCdYdlnvyK4KCCVGMU2+
d5maMnuE089ztd1ZCnkmZem5zt9BH7H8S35KqxqxujbybkxkaZ1dOPu9qWGLuff2
vIMx2uIzs/asO7OBIsYsIc0gi8pp7pmfniUq4KCgeEV6iykg4L8Xq1rCcFxcxKwy
iYgMrAKPOyByZJ0lt9dZxmvd9VSWqN94Ckm/X9VzdAZqk9pP25Rps2hVWcTnh1+u
0UTEeniHENIotvpAoSOlRnltQSOgvayvqzKXMHBNl1EkHYNs6g5qdbRR1Tby7FdS
rW/hoc1b/Q3tXEEB0aKZ5GyCUntyHjVqnM+EBB4vBsOcw/tJ5Y7X6dxA/EZn5tNg
HPrax3CS9lXY7Jd77zAw4zN8gDFpOYqpVp8r5yQ0op8o0ITaanrul1B7x/pMmOgD
gD86rlrq7KQm6/6rzeCOUWgx0DfV84QXpaeR3XIdNsRweFdT386+rDw5VE/pmo9d
tcgdvkfUb6eon2WwnRoXC7oyR0Rqgsv4dWHQbcCsaS3g8bUojFxesgMsYvjOb+6j
9eQrV+SFr3b1pJM+rxNqtUJgRxCKbgKiOeNRMKn02AC0hhIvUaly8u1Fz5hofALt
4AY992KjU2VGjA1bDdMZd213JlanZaIYTOTqraNOcGCHbS5L1UIaUPDM3doDFMzF
qGidAisxA/dZVFkwbgVzpRyzmjQBoB4TTf5vcVU4foe/i9bK2GL4ZQuDEZEWK25/
3L6kJWNtA5z3W4CtSDr2O3EcRP+cxhcHuXKBbOVl/Bs8dfWGwWOiPg5rDBmmnA3b
FmN2bXIcoPP3XAKYufK7pmSiS/ZJ6c5mmxS3pwHWm0M5ofG04bRleKkU4/OaS/pN
86mtIUe5qD2QNaMsY2nelrv9XzPksZnTYKSp6BLXj81w7E8CVHzG5MJCDUn0Cj0n
xyD/9bRQFILgi6OQA8KDk5aksfqyF6UKTI25WFQepjj66lEr61RzheosLVfgtjG4
7CUv7PoMj4qqZzhVzE0fSf5ro7l4K4XKPazVMdNBF/9ZpH+KlUydrYjxHEJliYHH
PsDfCocLjyBF/MvvvWUWNj1AWa4+CZ6A9M/9tnMFVXRl9qDvrzuNwipVqCp6G3r/
w/HhKjC9YjxAYdn29GrgyavS05tfWTKyXqKXnn0yc8qpErvSvZxCzKC+n3BalMpg
KkOwgWofnMHKJEYc/1smPRtlWwbx33xIYuzCbldHBylsc9c9vmDXepZr+2l/s/xH
virGqU8hSN7CrhSoIejKlexxllhOR6Nm8YDPxYfZQ2MEOCPlPh034o8fODWKY8GO
kW9oCeUxMLttSlyMR/SzQRi08TyowGyJGzAM06tGI146XT0agcJH1z5PgwKujj5o
XO6m19DfJyuheLpSfA0C6rPi4bTmQfA4Yr0mrohVlxPNuXmgkXZ0QmgXkTS68qEp
Isc+ndsPBJEb4XFiak+658DODdt6jdlOoNbn7/8YeyYapSbg08LFo6pqbT4BL6nz
Tw8GJBoE0bIM515UtV/dMVgRY5wcG7JRIJN6UlTtkLMprGsSK2rpNRn2vPCa94mz
JowIAVQHr5xC0AckRIHvwKWFyEDXjSO31z7pZ09TOdZ5UY0xIq8vyM/fdmk/KI9l
cvotA5LmAY9qCya5oHwFaW3m19wI7II+DVobt373ncl2p6Ce8rkMCPcFWRdtLl0z
HYxzultrZhJOyrQAgftDPVoslKcQz0mfzHPE3iSPTkNUQa1EMpzfbHkM4rfCdPdg
qzdWRvviAx1dwQIbvvUf4QF906/SUnOrPwtYoZTfsldNEwvKUO/kaHi4zud2puo7
TgMvGggBwB+X8fMu1HTR8A4yaeL6WbThaRvYkh3Xg/gsytm5xQZ1xd62ZQrzjCV5
OKEtNX8L+AR2NRr3AiAZVNP/uZ4IIFu+9rtryU6YmFYWQ+97JqKwAjP61UaktXqf
ew0Mhn5YyopLKvOcj/+F3W1XlrxSdE/tgWCw863FCRw0sYFcH8OApy5REHEXgyxu
Cc0Mr3KZzfFUiYHDjTN39rXlB9QlJw08zYAym738+DZcu0VkGQAAfoYSBwQeM2nv
8k5EHYsIiT244S8BvUC3BLcb++bxSULpXcKuxTWnskfcsHK7zcXAkudHYlzw0k2R
K06XD1swNsVLh0P3MUKvdFqBe7LOk51+ttdo/vk0OI7EmefuJmPQqesLIw0Yeott
BE45rZF0mkK1M1zf3Q5AKNN9m+NwmPdjtJTpzn6G94hxY1FFXLcZn7KTTASEyRZC
RWmMI7e5BrdTkPrRuULVak3bx6PrvgOFk4ge+4qSGlfr4sxm56Q67X6ze+sbCSTK
WZ9l/ZwZz6HOf4ojrlZrzOLqetORDa2C79E3dN8x0N0RTwNZx1apmpXUt2frIWHC
OsT8YDzYPrgs1eXxBNV2p2ga1MARm/zbDskqY1crQetouYIypAigcV+wRRkoL2Fw
5ubm6y6OxrnNxdOLCfUgwVo6dD27WfPk/HkNoKmEW8yBkirKtk8YuWERB9XsbcT+
xhZ14x/UMgC0Cuuqu+PtLo9qCMBaBm/bo5AZZ4FLOMhApYqHGyajaJZ7DH9RL026
HMvIFFi5orSYYDLzu5L7AulPGSqRXOIX3CKVDKF0IEWqP+z6mP4KbDACDnKOqmNI
8tNPJbJpH4ss1qdhLSck2dRtU8WU9uKCEv+YuyziIU5TnVuxFvK6CK6lk728F2Ba
6W4D6xnoRznPp3E2yteKy3nd8ulnY150QkNQi90rI4jeD15BmwR9WILS35A3kkH/
CAVtV83g1CWiIthMA2Hh7vHbYvSreMhwpkYf+L5XjBtIpE3g1B6LMwiB7YG1VxGj
u8+gInQQRF/1/cWxbl1kBnj0KLaGxnXlGtnncXg0myLbyZz4ZPCHoEsCMEFXbyAP
0lUxCKVnqoDstkRo9JFw+G59pOcbrOShGvYICOHVIP81xoDt2zaeMPHKGRHbEO1p
rhsieENlDzF6sNIpdG6D3lU1lN/dWOb5iV159bKdCEParkQDczPdjJW1gFTpNMqA
nb6UjUZxBGPZYgrjGbP04PBB0FAJEkj9sUZ30oEB8n1pbOHDW2x9ZgCrVvSA3u22
Hnc1o+YPgfNWT297qJiAQNStzm9TnaYN/mLv2DPVwz/AS2HgIldf8If/k4UXCz0Q
PVXUjOo7YsGgGYlnOGXjO9ZqKZcmT56zC4+QCexdhr/VJj44ZOKZUQfSB4PTMMFl
I1Dt/cDas39d1c6aAdm7hMYw3lenMS5M+53C0ZvqDipLKiEjeGK00R+4xGbpAbhA
NyCI9++bU8D+yWBmbfaWDMA7HBnmuTmR8Fj3jZwL2GaoUcAIICJZAUGOjgZ/4Ga9
ke6pgaiL4hqmg2ebAKb0unaOpIm5nSlI7FqthQxK4NcsyAur+rt/Peg1bdcTACur
vwSlfqa4cocrZTENqcE3lBHDH9/dqrTJ84UOREgOIkn3yXVrey3qGo5hCu9DOVmh
pkewEJExyIRzgMOsA+J80GPzwBzWfAj1W5tLdI8le1J5ROEmsh2DahslAx6HJPdO
4zOJsgowijPuEbIlh3e/ZssUkiMgXX0SOlCxU3B31FIjD2YhHayF9luP+OFMDZwj
hFb5wvdrwzK1mOfeIdFSDM9CZQ1/dshB5dH1s8h0XgwtBYAhij5Pn3fhBw/fAel8
qd7H0DSr2BS0xvUp1zUV2OH2vHtw9CbWeG6iEdNiUAw3wrCGpy4tFxguj3QpHMt8
j4fmry7XmhGR8nv/5RIlqwbYVhALwx0VfxuXypdXBEB11hAXxGOgyFASZRA+N42V
iwlqUQNA7P1yaPAKk55r2oVrV3rIU0h5dVVL4RvysohbNcgrkEVOww+mFLc0s+yu
bHV4dMZhJY0dOsWIt/MHTAcuvwgyDujRv0xcDiVKa3PyI+NWNCp4O3CRVjaNQRUb
7GraTeyT0nnHpU9dnUNf6QWRVvWx26QlwKUg4cPCCU52N4UnhswgT9XD+sSsEcPL
SbqVaOf+LqQf22UfRF9GyKpiph0J4nszn+hiZgh6RRjDC6bfgc75Awt1f1ZJamnC
/uvJSIkd9KQ7TtgyG9j2ouH/iG60FCfDB41TveViOfqnPR4/zK2ZR95RwautqxFD
FrkLnFBSa+W5OBYldoQdbOdQvnPBmoYHRX4o22oSARCEZWi2YC0M36zGdbCagftk
zzsLcUGKuhaIwrtLyCxVc+EQgyjiHPxTW9hrTs49Q/f4j5hUScx2LxzDlHitgdgd
cDI7N3hK91zd3eNTh7ARK/1Swx4g2It4I/TnwqCR2BBF3wMF7llOKtZdcOJeaG20
H3hyZiTBak7PL0E7HmqhJUYAf6HNEuhwj/ehx/uLe2Ov4l1klYUcqLsCm2wcsxg/
QXgyDMwi5Z7XdZLxxtMcMdVe1y9Ozk1p7EQHVqSJy/Ze8jNAQyjXOXu7TKbyuCyT
sqQ60WW7krqw/lQ6g4Rn1lw5quSkgyRuBDhelZkLP/IaoZPV/tGLvyLnH4SSDCbW
IwbnSTTzuW/zPoMXqlqlb/MflSdiggkDtkYoYljtFdYUCHyzSPpke7J3jFlalgni
HTgvxKwdFMgkFgpz26PixE3FXS+A9Q/9rbn7nWKjjURfbKaAPDY0tNib5edah9fQ
fgBhbcbaF+u6HyAghoQsYm43Ti2mXihra83NyfDk+uyfbVhidVGNGvnkYGob3wof
PziRhYIW6M9H/X9L0PzBylnkRt5Ds4nimmC5O2bfA/JtnIhRh61vNBBfT19ssWmI
pweg9/1bR5HKF3V3cOoygAU8qjOsNchnxC6Buwk1JJd33tEGuHkf5ni8+4olUIzi
YiGxEQBIgNHrE2EjQ6siFhfTTQIlH/hTeWWe/WBhS3xdQCxKqsbZT1vAXw+Ntwgk
eMY4OHWMXvhAVtssElbkdr5Tx8JBXL33pysf9kdlz15XUCd/WFj0reLqhNWzjcH2
Q6zf4nRK/CGvwLFj/kS3U0lgRdDTVGZVDzVHUnET41ZVAyhJDO1OXDfxjW7DRdIc
wmadWJqjNf8n98XDGxAXta2V0FQ6xtKHb+D/4FTHMezxg40L2o5XYcmR6wI2AaBN
5hfj15jVltbMpY1rJSvyathGRqV+jBsVjNqj922zgZYwru5Xd2piHFlYMAhN3UvM
XJ4Z6lpp3TPCiIwDZXbinnYCw7elqCVwoBEbOEs8wp93z1zxFTyUDfc6Nb7IEdfD
TAnDjb1oHTszVbqI/WPzZ+yyMRxb4Lxd/MVldXeCIcmapFETgZaMQU2/A7oMEZEn
JWB1c1nplKAr9OyXCB4VYK3Pe4kWLVED9Ff2THqv+tS55leTgbRbb1IsNItNZzA+
nCU55QAnp1Jd/1R7c/mFBqIymXIrVII2b/dlONweEpfp5QgevolP67mhffVXE6sw
PuL4hAG9XrCKpf80UHhVM30OpID6wwiZYYFpq2jqrhp2TzeW7NloKpMhYDHxA8bm
kEs8z4okps8DaXwuA65ek7jywfteGFMNjG1CPJgb95Menvl499q/JU0e+TBOm/q6
jFrexa+8ulZ46Mage5YsggI6F7HDFyaJHSV4/QT5ezN5NgCGLfIukFIzPbdwHQuV
uC9DcTLM+rgQQFfLYvMRgIt0LmoI7+HWPtYT7v9Mn4xqeg8fxTVtIjlHiV71cLe9
EbRfSbPI8bOdDCpz14UH9qq892qhdCe6A/i33ouz+PvnvXYiVoFJO8pg/yl02laV
9XoAHUJPYJwaS+S5Gj291+1rdcSLFdOd4TgN0Sn1D+7YneI/yTRBx3oeofEP06cD
vvcewsFHZA7uLLXWU+ye/xYZvjYwOwzrF5jq4E5ofxVyvDgOGB39ma1JCyLpGMFW
ZCgpVOJJTATBKdGJzsNWT1QQJL0o+Ul+oUzg8PfUs3xZGcThTisDJmVmQqjgp7F3
IZhBgOhJco69ePhinflGZi7L/TqQMaxLq9k+71J0SSVZnQXZFmOOiyxt0RVI9ZqF
OIH9kWSFUWCfVGywLiw3QzpySx9vHAsllFev794R3Uuk5YQS4EHCshH1lRBp9D95
Z2rGfdDAlGH+kQS+W0GnA91IQ2FIg+L+fy5U3rKgeHYgxfSm7O1k67dZ5vTNLXF+
Xw7wS70jjIzoNjLkc8BpQm32dZ7khnR1Cy8yT9aS3PSij+nSOSgh+OhEDs2VJAC1
Q71q/KC4QckjECjR2wPa2rjXPR5b8nQFeZIZpd5JzmA+ZquBxXa6hVwAXxRJnODn
krh5g3pGqB/cjJkJUYwNBW0AyiTB8q5u4g0hj604LY6vcqZcJhVBnC/y8CibJQq/
mtx/GmHNn6C3B4/MNjAdJkG2ZC3XK484dcSWRqNRZxAePhwQ+98T0dGA4o49k+Jp
ieVMCQMi98IZ1QQfOZlkv385T8pIWXVSMbIxSFmm4QTmWNsQEsF6gZRFJ1xrX1mA
kZ4VzYHHhH5poRD4dQh7BiIfVc6Fd/mCSumet9E2Q1L6/m/s3ROA3dwj30KeDVhq
aX2HGQlAYm+OP/qlFbG9rbByYGss6gtKWs/J61D4m1rvmf9qnhNIN8+HbTW7qnUN
l3Ei3stjZ61XBuyW7qWSb8aiN3Z+GgUu2/Y6SuKNf8YBbuPeICdFb6b//eayUiO3
nS8hZL2hr7QetinRXDXmS9stjzbEjgQZKvN9LwgZwYMc2us2MAuCEE/xxvGitDyo
40vQovz9Qb4tmHrIYFktetjRtOpbOTyBuBrRTlApAicMRudznHNCQ0+aXoI/c7oE
q6egp5LpeTOOVF4vYkzM5A71JvrKQDjSWVpG1C0+6ccFTJBnzxCtNid+gjkUcxX8
dImty2Wc99lMuZJ96GHD4rnmaYQIW0WNSC1eK74dlA3u0T0pWSmFVt3nl/LK1ltR
JJj7hCsZRX8bKI94h8tUs9A9MBcRWa5iMRYGN9d5B4Wd+wdcu73yR5Dz81K2omG0
lUAILwLh4gvk/VsDZ1ETv9D9kKKsOn4FYOiI3t2nftufDHrP0H5C3xNj26rGNn8x
wY2lIQ70WqZbZqOj+yElWJTs83AIYfvrWqxE2lDrpaPac08HRxyqMH9cHaeygpo+
g5J/Yn6zoiQfMngdRAkrSfbZu9Z/k+UGgijMuKJj4gb6WNtmwwuVE3VY33qancJo
weX6/BQesTekQ6wQT0szsyshzZ4d25wMhhVONsyrxp4R3KXQWjxouu2jsJVStviT
22+kwIaQngjPKYPZltKPGqTfYpcwXVeWz0xUwx3eiUa3xmxkUlmcA5qcvktP0R0d
PUHB9C6amNRR48ELb2f97hBKJIdMMGCO54ks8XTObmOnjTu7XHwll9hKy84BoTOF
/psvf17SpEORkA+GkidM91nBELKsdIoMafSHlQW0kiM7yVCMeO8eUR7jB/HEpF9Y
Rz70foBxqoRz6V3L6HYdou4m+udWc1tI6MkY8EZAKcGzKh+JSBRNz6Rh2GKfOFqe
ovv3LNjtaB0gY7wt85qBMT+gABs4VQQKiFh51BW/TPrQlvFT/F8Fvy3zgQwXbQTP
gLl6YE8b9CnDlCB7dqFHkZ5jZ8NCotN/sOcx8YowKuGi4Zb0gUyFULYt2L4hgoJ6
81qC037sjDt7Q0uJQV/Ti8yGSkE7rJ0a7ctPI+OR4y0z+mwtTMnupb1ccpTEn6O7
FNS7k6JvapEGw3Kmv5L0lhRemvRxk74R4Qfd3A4L/Bx4vZqqmRN5IrVPQFvf+mlM
85ySYZ8PKG56/Kb8m4VOyaU84zwelXvpgnv+wBPK9eD4vnipnqW6b+SRJs79VGs8
A/9T8VOZow3Gh9e66ZO+ArCAghmn64zb551xZTS5GT8WLIRlDJKKYAWYUM0eGRdt
VQmuoTlJpc813JyPHrZZQ8IkflDuMM5SA+3V/VW8kvwMhcSOIDXz5DuoiAwMfcVA
rJq85SyBYgrskeUp7gbwNLNP1lpBpgbcShIts9Lio37kRggoOIWoWdH0IXbc8ZhK
ioedcCd9KK95iwG3L/qsW42xiWQvsxf1FDmMZHL0B5TPeOwKBvRZOIdaFhfbpROR
MNFvODwChiRDNDfXVOx+TOcw1yMrmiwwRuZivg58dpFZi3ej3pq8JbJEuWEzgSAV
mxqKiZSgBQaUeHhDoqDw+P/7H5FcJMDGd5pfcwJXb/hupr9Qx4utHkuXCJVJG7Qd
mWZNyTCZ1baZIGbdUhFhs7sd2rWdV8TxQvkN8KzrVYuPNr8k5pdceE6CmcFMyAla
FNYOKWW7cjdl2z9XrGnS6gRKrgybNpq1N0pv/UYEatyDmiy3tM9ra4vLl8gatEIx
o9JNVe6ppwHGZ2fg5HC8lEW5gSDLWnvO4KAAj97u3GDjgDW+t4wqY+4afK1V0HfW
JErqxAPXWY2/k8rAjQ9pm1S3uoAsra3BmGolFBFvjaAARsX5u43BOtWoGg4KA43X
BqEv/+v+sHSyr2fYxDrArzEI+a9yP0Krr44wkZANqSn3+1aSTts7/wRa/MveXMZf
zrjd4R/+A8JfZOcM0Uh3DyV4nHjYld7CaJQU9olG9YLnbFlFM02vBFeUEpvF6GKb
rSMzZZRNhKfj7S/7WQLTPoA92ioYFGMd0DqyOP1NY7fMI0chveN6xABTMlQbqWPs
+ruvQKdDSo0EwHubu+RPbYgWO0BdXKTDaFnWhla9H5r+VnEMqkyjySyJJyExNqa8
5FcWQEKOzIQ2Bp+WkS7/YX8le+SimN+GQxjlVMvNeJHqJCOfAIMLIt5RcMDLhj/b
naX9hU2NmTvfPkPL5w8/OGaosL41WL+gYzp5HOwAyiqCAhh3y8SFVmsge9+DpOqP
TZLhp1veGcz2x8i7GqNASg2Y5YVvACVN2qmIdoiQw1N9QQ/Xvq8SVmCL0Jr7Sm9w
kKGt1B9UTUCG44Gau2tCABlr8Fe7Bcsj6kBnJXS9bq8raL5vP+U0XmcenThtWF1Z
5SfM4nG7z6M8XnSZI5GCANce9bKoNE/P30d++FQJpHM7+PXUr4tjGd5pM/ybQ9lI
HAciIa640uT8zdvZthMYCmcaD07KMtCFbdXh4ttY2kKwhm3MFWq6lrhxfNzeerPS
ZG0WHTWFxiRro+EDCi3H+Y5QHUrlzB+o+7Fe5byNNVbGK0aWOfgInbfgu1sMNmVG
i7lIQMYFzcK/cXw4eO1N7zOqi9WgtFWiF+pAeFyeBKAkGzGS4g40sI4xfFi1HbRL
pN97DcSsW4NRGu+x02mVX6OV0bIAdZT/sTMcqQ3lrONqpD+DbeGDpAL5IEvFzHSi
FNflOOYlmRggEWJUfBw/qG3LDzgeLJVnugXnyLxqzFJPfqzvEDB+U+tPVw2XE+M/
hwXTZdlff9DVmeAP/b7CnwHVr17BEN9pxetaSMmymqtr0yU7+26SLrgTkOEhf+OH
+Bd3ARozar96kFSIuw0c84+zGqA3XtWI2f4w2mW0o+EDanIU0xbYDxN5A6dxSknR
Cdwxk8cYq5X8x921JQCOUrghxXT+oekQ1Uk7F7B3RAZRE/eaDt2PUfobdWNcd7pz
mFWmxi2Z6N/Qq+UVmGFH/PoBukjOisNps6KEYW4fwW+hHsFr54iUlU66l/Cv4fB2
KIQ+/d6UJIP4inF2BgMzQigmfCZ7C+FIa9fWuPoJ2/FTq+xVup0P8flEEVqqOuzj
sbMeq6IQS7n8DFEp5sJjv3jwE3AJiNPz1Ajf9hVCxlqbAVIjz4u/VEgnitNAi4IK
qdtCc6v2/rAgncb4/m4VlPZgmFIc38XgCqc8+ZJsbk2LK415G7vFipWc0BUE0zgO
OjHj7SgsPx9bBW0roR3aZNOJjxiXH2JXVeGCSzIgjqwugH1mB/S7NzSFa7W2OK5W
+wWaIEf0XefoRCx439pYuZF4ZHkJFXdzWY0qiXfT7q3R52dJseKxXjW/rlb734ho
8iJdWcPfL5U60CNKsmVQ6oQcLby1lE3MlmUYMeupAaAolpbFIdLa4OnHWT97/CHH
xpI28ebDwhrl3cv+oBU69pVD30z/V5YMIvUr+o53YqLr3Ta1QPJDPA+F0k5iC10m
74I2/kDqzLGky678RSroOvd0rGcBGgvJvyvoXCnEYRNZFODSkJAuwL8zRWEV96A7
DS2uuMHpIgOrIW29LJwNL4Z9jnvj/uDEz68aDD74f3CdkX+099STgXDymUk/n9I6
nF9/Mb+O/vrI6/kXcM3Ps3Qu5jfe4rb1aDxyAIX9q4Ok75jjWkuL3CZkH2yK4EPY
eRpJ8b37B+Kiblgi+IOQ6FlPKhQSnCm7lm5Jjodu66lVm9w4nG8Bx/h9HjxzEnDM
I4wvxNGsTy1umhck/tRVQuRNXPnI6+Qsa8tUX8kpTNQCel5p8vcpwCCcxG/Yk8D2
Y+4Ch5lxIxhlJYNBxFafpyInUDtE3SC47w2BhxvFT5goWH+SkzytR1JaKTRRE1bG
TLaZWbVK5Y071l+jH/Y8RC833/Cc9KBnDErLL7OcBmuiR7CkIdxnK2ZuilSw0Yuq
+LZW+/8DFfNB2KdorIeCw49PyroL4LIO7AE4syMw0uTSvsBJ3Bj70m55wcx02ric
F8XDBisMnukPYPxJqXqU5JJ353tht9XMPzabRxvScoxaVLpm3hwEAADUMpR+Rbnr
ej4fm2sKIT2VgzG0zxrJrvSKSvwwcXzVX7DDShLbf68vTICEGCJJ/Gt4eZrfCTN+
l7An6kcXkxufNQlrcObfqdnBhrk8ZC/y85yPl3HprteVI8qIapXBxmMVgX4lq2PB
qaJKd2q7Zh1ngQOdbqVLXq2U36x61Suzmctc5Q7d5lbliXvEH223oGZ6HbuNmAQ3
PDnEdKsZ8TILlpfGwXzwY5myLGAn+O9/r/SMCkyTZHQQn/oHUKlGUP8TUgqu3wbw
MAcwaVBAo9Vmf8CcjUX6QMG+luY2E85X1RQg171kHgFUurThir41vqAPJqjU62qE
VyRKSG9W6nlrvHNAZNTLk3uuHXW1IgIf9U5Kg8E7SvvKujJJy2V1QJcWTtaDv1QX
T0FZOC/hOYGgDN14IRAFsUcPVWfKeu3bDs4r/3TAJ0+m0SFGSG7Smr1AlxFj4yDI
UjHfiQ3NHr8Fye+tohfxRfLXWxEXwfL9L+60dTzokMPV5stSzVoLlkvsWPl9hPDC
zEo9UbpRkS3Tdmnco/pLdIKpjXgLjffMSwTO9z9ZcPsW3geG8CFf3FA7gsbvzts4
aIbnk/VDaLgoe4TwN4EaOK3FFuF6mn6lGvElVTvYLEFDqKKs2RHuMrnyb7+KV97V
nYHWEUZbuVhVOmU8ABfBO6mEyBxmtVGScpHiqJJoQ15H6K/fLOY8IqBSe//Ay46V
m+7lig4xpANa7T0HakC6BVRNalZqVPsXmhPAWe4n5V5HekA5HvjMDYb2ZiwRTK09
9F8UL78WtH+aMe9EdBquqwaHTfw+it+8Kx6ZgityEnzKjWeJlNlRW5vesC3z365G
IZjAxlTLYfL+rxInVlKOt0tVFhE3afqVL6c3N1wIWCI7Hi4VeYij1AWu7ueMSQvV
UkPN66NEaSNHSv2uugjrMqpRZz8XZ8VTVaRAMCm4OMaiN0ROpn9GyDr1332FowyR
K1yHQZoauFIjS1uhsGtU6LEEyezMV8K75t7y2xVyVl8HDgx9qvvWwYGCaU5tHOKU
o5NsSy3SBLQQMz5ZXz1JITmoUgpLZR12SoP9hHL4LNqSaFtRW0CxIqRNun/bd46B
+f00EClImU5j/GfNDCgewzJBq1DyqE+RiuR9izjTeUhtNf5YSsl8ASWHDvDW1QQW
BQTonKB0bLkXq9vkzb/1bq04QYSbq/O1DM0ObGOzQ500/IbC61MmyWdhEDJz1Ja1
E548753gAPn4SmW5MLNC1zs0t8PxWtL42J53lCVmYUZAUy4aT+lPghLUNfTPMOVX
4DCn2p+1JgTooJ+hRLZoDagzOzPDu0ETpXvMfSjWdz4+abG2rRYn108F0wnvsBh6
PCen0iNhdejdeovAD3Pdbphbq20Truxy+557d2ery4GYxqFNZrrLUfhikxwuPjSl
m5uzhHX6y0atPPHMlaL6paX0ATItGRga3AAJULtLRzNnJ1mmbGEU+JQIemTpJ5sP
7B8YEcziA7zHba+pFct/jG5wMPW0VkVqsDoEWS7wGZsCrvOGEMrJC5Ry82VACstT
0LuORVwoYC3ojef+NkAxaIbEoh96XsCF9UsDHzAePQvbAEBYCii8kgdtb0y+O4Xp
Q1ReJI6TUtEQ9yRXaQSZPrlsrzDs0gvYM8CSR0ACPaOVoy+1Aynd5CE5+Tu7b3By
weLaVaUQMQ+eZtBnca48GKLZ9wb8TtBorjtrnI7mvaHIww1hSq9HyLBl/fN7gaXA
1warDgIYro8/DLq0IZluJ7jSTrh4lHi2myT6df+ipNxvisL6zqapG8sYN7r6hZRb
JRBmG3Q/DxBqJiBt/pjThVRTn6Zo3qu0BZ0AOcxQE8TcYTF+naAkebx5Bkd0xtG1
f9LRq4HNNLcTALSE4R44jZbCtlBveF/oHq/cZ5EbRO4k0p73nabO1zduIMlJyaJf
FD6YdUM6iuXFymTcYa7KmH0HKEnYqo6ECR7H7SO68tFZIEPC5K6+fE/psfg+ZI8F
B3rIR3w0XxBoZfKVS2CeVsT8hIXk5ReiH9hJxaTe7ewp8Dz7BES7AqaE/FkuaS5l
m9vXmEOFP/K+Hptf8z7Z3YsQbUcIZ0tRZGVpzrtGv5ctsN6Yhyv7eEDQA4Zzn5va
myOCuY6SHrDwPPthho74BZKZ0hj76Vinfv6jGDP+Zz72+v5qRKOU9qdqC813BxHO
DxCrEOOyR5Y66JEW1SVhQ2wLybytAecrYWk/ERu4X7oDO0XPQJcQopjGzvl74uAt
iAc3WHY8sPhEsPKE+Q4MQnBABwrfkgPQCFuhq/IzNCYjMdauLyPYRBH7R88IoGC9
MtpTgLQ01ugVXy/foGr9kyq6RONDN9fXv4xX17m6b/QH0QVPVQ4IfBM6hulsO2LI
Hti1jvAfv6XUqFtMt6zriPfVlEEqYm0P/7C/hu50FJWabtuT1IcnvZic1zY2aOCX
JrFkUJ0VfhMVdn/zvYiXTpkjnmV4iLKpJlLm9tD3L9C5PxS7HPZY+4xEvKmzcxr4
Y2Ce5OMH0YxZk03EUG5UNVWL0n8zZzPTvXOjmR2zVLi4URTzSNjPe6GXpC1JeH+Q
OWUwyYlgseImjVjGVXwR5qaOzrbQ8Nu1XaSGJmAOcaYDGOckdtOPcefCqMqfMHR3
/ubS2VU2lAiV4K6U5DLwXeYdOOHEh1Ml6YjxwDuHXkGDQYW+L1n7T6mXzOEyvmKw
qX/3Fm9+EHJj6iAeFfKKi47HE/QX/sLmkDlEpiH/emGYUOv5ZbtWaQIoUey4i/+i
96KF3rFgYGfH121WqIU2t3EhNQb4Usg2LK939EUrhSQ71AjUpRQ3Ow5zro5OQr7p
Wa1P+J9GkiSEdjMAudt4eaenAksskTx5ULXDp0fZSHx10VCrA1tyRKCImMGGZ90M
9K+VChibLEJPXbf+Qr1W1jTfQW2IC5KeZtgErhM36s2iYLar+t4gYfuyO2uCcRsg
X2SWQrTy4VdkTMWeRvWQlx7NbtVTBvDhld202RX3mBD9fQp8rQYY2ZcWCZfvZpt/
LfUJR72GazaZpowQrD+X5N+3gkkBwjS+JJFyv+2PSRY7iq17neRlpzU03RYLIkWC
tT/zl4V0xUVE1knAvRVyK2IO70p+Z2XdUt1wq+Ijmm6uPCZ9IipNxjoiht08F6I4
z4Jh6jDUCeiJ5RQZQ0HACD/igzb8la9GXVVpRRFuE2KGDm0Pz71uyFwVlF4IVHwD
qp66Ped85ip4dtDSUAdU13+eT2RQUn2ucRI58pX8TziKQTrfoak80z4lOYir9sri
khVa9ZBOtozKjLgvPqLCTT8ROWnpmHo8THMZssYs/SDhpkKCAaubWNUY2d1rrgxJ
gds0g67JtVO+FTeRAClVIQW+UwAkmySO7Z2bsWw0ontgHJOMTi4rAXQzp1MMSArH
Ykea8dfLz4GhBGFB/7ECgCK3yz63I4YMruGrA5U7WdWUEyVgcv/Cu+qIROZrL5yH
+7wb4bmZZu1dxHDKeBowJ7dIXm29MNLMA8q9rZ6q1/tNQjWPDiKinSL8KoJKPZRr
2MT1p6cR6dVbidHpBfYfURusWKH0uowxbm7zdIprsqM2MeGfvaenYjQr8zwkta7+
tB8UG0E6MfTX3oeqaQX/lDEZOyDkxskzzgMLPnfblFiBQKWKHLHcxPIPmDM1YzSd
tgN1YQELwK3IsRVi3D4XjEFCMJ6wrkAgDuq9FP04Ta6sMmVPi+RdYZuX57NhPUMh
QCeG4KXiTEkXII2WbOSP/GhMuJkiSOYM9NdynRhF1gJIFt+xwPRHZpbXu+//XBTl
TSJlxKcwf2aMip/Rnl6xBxdiTmIWWxe1vbO75lC0oPmfOaYJa9HzHlwIVsFphEEZ
C+FoovgKqTaZjAHaSlrSaObom0FAx2hlxhuvtpsFwxEA8UFJ7hhpefcCzLPC25T1
ldOFzGjYbrnV35S0ZHLbd3k2jAwugzX+rVZt8aL+pTYyXzFVhB415otJpFcqLVhS
Bx7Rd4nk2IZ1hty5gdMDR8gId6db+vCGbbGzRMU3H4g3HnMcsVDmvsy2PVS226Iv
GQK84nEDrHiVRYd5so5iVKPwL6nQ4Mo40E19vGH23jhUzR5wjLhtnXtvwCJgmOc0
hNwCgEIL7r4mwzeKOWQib14dcFEOIsAcbYfR9h/oZGFn00sjiBlSXhUl4E7c4Rue
74AsClGyCk+ISlBfpLGiviEB7z2tUxxhFm+ZOHCIJtfScP2irWl4nt8iY/hrfz09
2n/Bgki+oYDvi+LPnNd8TFZnp5Wlzylzf1ngWaDZHF32xo5r/pHJy6jBiXr+i5Ws
oLulHMSHjvdQRQqtCUiYjIyB6qqwgnzekn4rIO+UKq2HYF/Mc0yxUG5JlHU+GZkv
xOcyNQY/+4Nodmec0CkJ/HMPz45hmtL52o1Qb88FG6sSxIP72GXMFGpEUR0D3IpL
wm3esQtl/XjbH0jWjF2yvKTSyS3W1qJjEqNzH045dh8T7zD5bWfgHdQiWRX+DhN5
lxmcEDSlHoUjm1Na6nGYioJbdkSYbYCFXfdXYqS20eaLfOXkAN+fhnYJkaH2RYYE
zo1sxOP9RZrLkXvEKNx6ICY/rUUwRAK1Sr0d0SVttwEhKP+TyOQuEwOyv312/0mf
zfhBnyfJzC2oHidBhj9+hyrYVTCG2UpJhDoq9Qynvf1ELaMs1pGoexwUxXNyGZZx
sa50paORteSWxuKluKNKlPL3qr8+k8xVVGpFEawnyXMmNH97P+tzEac5QZKRUQp3
qlr4edLWyc42b7UC4Ab2NSzor9aWN5wpCUwJFK7RR5Awu6x/5dHbUQSvh+sOw2rF
dgM9GRKvOm59lTdsz/png1Pslec2tn7tt3fOp1mm+3VSH+YwtHuvsfqFnajg58SS
8G4bjltfKAMNnLUBULwZk1lDnfUeaqkZG40tVJFMFpNpShbCtFouyHZl81yB6a4q
ijFrNaEiMLpIqT3Cm2V82VB7fGoc+Ta9vl7MUjcF0quSuSznIQ9XZ7Ne86tZsqzE
/npX1V5/U/2CKKK7bhwOSAUzxOIjDybrQ01fP+JtQZBKeGx15SMIWiW8abbxSRHG
PfUTq1zd7ohgFPNHdVhR8++lKqnuAm8j5usiN/tnc0qAIf22G4dAdr+aSCUrx8TP
GV3gPQRRbUNh0WFdTT3tIm3v0dySrqeUcmh0bNFKFQwnZpXJb+mWlbRFK9ByA7if
0hyS3RFm8Mu8UQugwOL5cmYEfmnqgfZhYz1m39Bi5WyrSAg0YragNLPDLRU9cMe2
ZXhgGVsjoRGu8sF6ZlpJboDUfKFse6w7QXtp5iBosVP2v27q0/55i4mNbNXKppWJ
SE/04+tRtQhEtVlpZNylPCnmoXhjC7jfwWZmhhbYz/fHgLo+wit4AfVhy83tI8W5
JL6CHAPemA5AEz08mWUTBPRufH/CWN5LCSEIgxcSS6dJsQMqEgRl/K1ByGoZGwki
vhKPjSqjxlVwtWdMJpXPFV+fxXWgnklLeb0UiAsPVL4A1x9nZxfeEp/j4eVzY0OP
yzpi5TysCYUp4C56rCZYhQOX5cIiNL1WKuKrdyRhnbnNJvIuk54AFLA/c3Me+v8x
pHeMmJUpjTxVBKWmXRwcp3Wx8lwIzGDcq3s0jcBU1ex4qVekP2FwtqWuRbBx5tiH
V9aN+daCnhRFbHM/WN7ickMgtDt+kHartMMPNbxS39ynzjoAGN7YxUVCjD+p2Ifz
2Nd2HfmYnCoF0UlJEDmMFxJxuyAX6pv95S/k7PIY8mu+St9cGXGPeVLHT4VdoRwl
LJ7eQRRh8oytoWpDEfoGHsbDGBygVB2+/GlJiGrqcepyNhBdo4DDmlQ5d5mmWflk
fmJ1pSFXl/SjHlcPwAR/gkYegvkaaaOm6Io6melBgkVq7+XE/CHsDOAeUw1jqM5E
X+VdQeHpC4UIPYlUdkiYJkjd5zsikmMPawxxnD+GOuRU2EM61QLLKSgVO4ObNzY2
+cubaZyXXIGDqF2Y9yyf+4hxpfpdMZepiSJz/J73aAUtahV8gAVzqGj5EIMdSdwT
T+0Ow4YNGBd0fRZuK6jeCGWHk1wB0eqCTe1XoFa8/GxDBWO5tIWBJLBIF2hE5FE5
SbV83I6FbxeJuL78b0WWFSM8hCyixJKMC6Nv8iyPMWyh50g8ogUO0k8UAIAg43dn
xRVzqTQFOyNrzfI0VYLXhnZJ6sTA6GPpyFbvUnMsn3VlMyydxIkw2SLOmrZP+leS
JUMXjjmGbmjgj5IZhIspkWUVMQm1FgyVE/0RdNZG0GQJMZmkDdwouKftE59HgU+6
/rFPOAavJXLYqMBMeEswaQdgJT2m890Q/uFplQVDd7PMQyBQfuqLTiFeV0xI1apM
x/rB/xkGKVy4lGbno3GDsXQDid0pTmf+2nBlidPEL+XAiddkG5+RiQzoyzRn5E1l
sky/3FWf+IwMi69bUWQJ5XeoiinDUNM9e8LG/+522GJrSzeVzA+aDY8Q/TfIYUK8
gDnfaoePs/NGD6atFSy3bU0GMjWttWHatDBg1QntAWMjddLav/VQiH9NT7E3ZMos
SOc+F44K6UpNKn96yHIOCZE9vZCS7r18mcYvG6mXmX2lyKfFzjZPeKpBtEhfj/6B
7RKYgPWoHDQg7yt/rKLBHbu1QfQf/gzatGqb3ya5O8Syy7LKB48ud+TZbA4EGhBE
3GseeR4XefaVq+lYEtQcxBJOZAKTJgJaiM4KUQaIP2o5oUYpt2v2ARQvmucoEY98
oUOEU90XnHOYSggrgmsZ4UuuIjMdfbRhLQ6H2jXoEnsmhyA9NxujmEW9bRWaEwle
25Q2MyfALfrqHrwO5XwadG4cUCsAhpc58ozLUxwIT6edhffhgwOLK8RH4sKN6ZQK
3GB1K+3ez6/vlakJ+mHT9yOrhTsd6EgnX0jchjEmXPGA8NgEf75VyLbu7uu8kdv0
FyPwGFXesKpfIiSn1yW0Ry4+nlkrUw+D+njunB2WhNzljsgdd37FXnREpSmtwqZx
c+3FX9hAGLt9DlI19M1wRnMdJ2lmcRrax5rmSKM1AmIirVMdA5JtHWZUrQZBRv6z
+8bmkYM/v1QS51FRiw9n+UscuDzXSiWSCzTOQjmZA/UtHeqkvKjuRxy5yMET7mqK
jPNpv1JgwyzHk37uB0SI9cNJvvfBBTrWE0t6It2AzDhbWYzvHUwAxub4YCNb0rYq
P1IBVCNIYWI0v8hqIujMUCE202QBFw7EOe6aMjJQT1sJI2S5IpeKyfdOZVYNpLb9
+H+NeOrls4jwchFTfu5Dv04aY57HKAvU+m9xFjE0/VbI+22cg99VfW7YbmNYXiKv
E2Xt+0ec/arTZI0SPfmIBVquJtSORcmZJGVDZeB3VvlephB/vOTOmK3IHgK6V8WP
nzy6iGfYRCTfTLHJ9FchR28TR+UgsUJAOUwN4ySUY3H4td2F4KKEkGuoqMHftMwC
OXLAqrgEwnvds2ngx0qvfIxdEuxLfJqlhP8fcLJ1mHJ5B/lEd/RywenzYXWNNFQ6
A63Js95b9hEqMIwyhrGzc6S/QSp3DivX57LFXCSLNjaPvxyw5Fp3X4y9hhNdupv/
0Fb7IFMyyoOqCOf4xq3Vxo8K8nR+HoVNq6dNu/UYd8RKwJIqugPSMNe6gedOs6C0
lz8T160+Su/tvL/+HO96taI7wrED4+Q0UNwQOyOQ4kPTfRWm0hZwQCx7I+xz/W64
2j9+zXY1z8gPQCACcgxWWMeLQkqR1lmiD83yD35Nmddwx2ZbV0JDmnqwzcCgsqqI
WHj1JnEJg2oCeOk+5HVF1/9NH3ziOHYt654e3loQ8lcdQqN4e0rGscqjVZ4uARaG
iMVWN0plympGGaybLgLMKmsCM+hSfmvuv/fHCxQCx3FULjUo1kdh/Y5qi4kk2jxe
bM14dxNQJwWdKWSXHEq5UePFjHxKq0wOjev9kBkDOzUqK1081vLkgMFHHWdxjE9K
f9fB7AxquEnY1Z+H7L+I6ZP8GpN/JoctCm+OuQ+tICfWES2QIjbvNp3cHzaWw3HE
xxDzVd529JLbMfUcNmZ0R9EWVnRICLNZ7t/85PSpdE6zfGHzO4vJoeOz3AxYqsP+
mT5rXF9DetIj/oCCcnEfulHMt15XXX3Pn2HUvE69L31pKXEsg4pwn9MnfcK2PizI
0WMJ0U1IPUbvj2PPgzhmFuwqhKCKqg5NfFTlY+7eHWifvRTcQH6E2ODTS8K1R93s
xLqD9f4YoeKhiLjDCysM7ngqe4MZUscF0RWJUrpW6ABn7v00HjzybZ+Vj41E8J/w
MELJM1FrypvvSiC4NZa+/CJNws36LAiQttoMyIxsuiZGgFmBqdLcCoxNXNUGbQOO
TvxhTONFiKENFmCkfvrXJ2jyNUCMmFj13iMcc9hiefG3tcNyvRAe1+Qi8x8VIMEI
IN4ZPLkGX2LUEGA2aPd3/llepjXKsc/fcENWTb2jhz/BFIxA0RmNljhJqOTq6CNf
yZ5yY/28NFeq1KFIleXZWpw/GgR3hPDAos9b3a9L5WeXnUxkIktjJQqnfOquKC3Y
Mcsg4FvY8Y74c8AV6kcAcyMR+3OmmEiRLEzYebUeolFjWj4DfWLiZCN3HzaGgSiu
hs+iQ5KHEw54FEC2HtrU7v7Bt5ECHHzzgy+C8r7N5FRETwl/B8Yxj4n2LtOY9W8L
FpcXD132rjwXOhiMFZZWRQL74a/0tHoKxj+DJNf/w3+ifY2XctTCeO+CYZjwqMhy
+0BUkoHDXfhW6SSO0GXHzkVYBMSf2Cn9GKKCGAEtU70Yx8KHWpL4xcVCDsVir/Vp
iVMkKTF1Ct7QtutjN4gwFPlx/MjekJS2uuC7ZQ+D1SnO09SjZI2HDX297ICjOwvX
3ejQXEwuugPM2zE7CWEUtLvo3vIl0W84aMGbTRf1O1RJhLaIXvh8fGI0KK1zgKgw
4OBgAepZvnr8OLFCcqjz9kLHJaGB+CDpGT35jAaoK+taYyDx76Y70HaSL7bO8Cjn
gjqW0/uGLo9hNqKqVdFwCvrCxGKMw0ggVuNPbtVduUd3xmVhqk64UbHkiUYhxNqv
8rmwhW4jPRQb8+0wpiO6PlTIejQdj+54p+rtDCir9+zUUu8IxZ15/gLMeDRlt12F
jZ1ZDXB0vikbBpDQsmJjnXculY1ZP/q7YzxnZGBg4DfihQTZDIM7yabF/mDhAEOd
XiQIfrKB2B2kPLf1O/Q1aUCNi01Ek6V91YBCVt6EcDZ1Cs5HCcIRoTtNS+lag6P8
X11XYypCELDjc9i42QTxWm1SicTAn+6ZvLQQ8DPfF7rFuNaddJgy2aN2IEe6jzTI
d69S3x1y3TZCyTChP0Ln33d33QIfzOyw2D6cstPyZqR9f1Q8Ms8j4JRLCtwq93P2
MQin6TdSiFextRPLC7iozkUS3TtNzZjWaIjQNkubdYvmR3IBBuNi2kfA+gNoj/lo
fyk5kebkANt+Pp65FtkBompEonMy79Fc5t+K5cYHce4fQVR91z/gsa3msSOzwq8+
DMSc2+tSxCKx4FEd9LBOec+2HicQMwT7aecOdgF8vaQxbZhdcujfOrCgjSZe3rda
et5imOmQTIn76dZ8ziBA4G8WlsX46A2z72UNFpZ1lNG6uVsxjA8a/aMicp4K1lRd
VnLY3H/hsKLR3SszFqXJdr8hCcxEt9Xpl8l3s04J/hrVLu/fbkNFgYmv+4h9hd8G
KhyXHSlooFxC7FigkWGpdKc4ufQv9saGziLnhNudN4fGDXUN5VPp97eq5ING5uKF
Ks2krL+nV8cJutDOW7txWo/kRbS4QRmfxrtV8yHZMAvfVYe3n2mJoMTqLZeQ5qnD
R96MY2ZLITsSFSixwmSGjgXn8vn+N3HXTGuSvDrfvX8zTTCKyDM867VJYb1YHK9V
fTc73RH99At1D3DJWg+FVQ/WXHVPPdGP+Bw7IHSlvMGQGk34K3UDuatklBL/qPn4
gO6QQ4GSRDxShtuOz7uqad2klvoEdnfXhnQ6U8XPTvo+Q3J0Ilu4nAYB8+SG96Ml
IfSdzR7LmqbrAS/7SrItuc1IsFkF+tdSspqMhOmQUZJtObsGxQLczaxSI3aQ0E3J
tg7TgvYBizxvSDkqwZTQVrTR4iuYycDBSaoT/0Fkt+NmnlYjEuD8HNleyOHJLMGu
cKRvw5rWJ25m/1FlxZl/CHmo4dyR0qz1Pdkd8BXAUZvw1W5UEUym0T9XxSyobUpH
HHmFX+b5FXpJFmH8mOq/qPt51FyYTfNwOk5iKsT9bQa4ZV1j1Qf6oIQswx11ByB2
CXXNwGUa0jXlsw0WrUJJy7m2+M8YxsRrKrgY+wMmSxa9pdDY6LNoXPnpuCf9I/so
6kp/FmPLzqELz0Z8CJIVv6NoV5PFXIkqlPPmE5UzYgqRcnDy1nb17Nd2MPIFjw9+
4qQrkLYmzsnmw6GHS+IRy4SAr1oZkp+q3TPwq9ZaDgJ7QYb9L3EaqAVHU95YLmh8
v33c50QXZnZGLYVpiMpwT7pCRIGRYHY5m0sDbvw9z488S+SA490ZwFGj+XBsKoKx
H7pOoRSWLgRD6vXyqttN8NFJhOtS222/uX3ZmIzCg7cJEEO4Fg+eqMBXX8bUv+i0
HaJR8g8BDo7LqTI9GiB/3QNEilzx6V4FpAyIR7/BuBAWgfx4ywvyJWDp3rZo5wp+
ZF22y7O/J5XlfVkexFUc2BeYNrAthZdYRfpu9DF/rPM77uV89X2onDvHMlfxHMMJ
bwEohvtpyQhppUVUWK+Cx8wQa1SMod7CL+9B/vPWP8ucgR8QtqX1Jgwhy1fz65cS
4gjTjDVOCV269bHU5tOnpso8WqJiRNkvE44yNdEPmNNu1cBjQ1w5K5OOz1NqvtI2
4DbpVhK75/Xn2tGxJNI29/RFkOCAfgcnNmhUS+yLa6n9cxndHtzCSImcNEtrQNSQ
+1OXqQQnJ2PIafmtR5svdkaZyvc10bPmdUictnqzXw2bSU+5A38Zz9MYYXA0NJX5
zoEeGCEWZ9dEyOOvDwbI6Ua5cSSEyH10ECjq+8jPPJbqkOwgqUvXERQnHbuFUO/u
YgzulTCKV+zTuFKM8yn6wPxDHiI9j81qMrWahETawh03HYTkcGBuG8VwFdnDi+1H
OJDcCrEql4211TBtw58IU3KPJWpuUAvfB/3b0uq3BxbgmBsI0J2hCHTyZygttneT
GKWJQr7FH/K24F7wX93Qc34i9iQ1LNE7fLwwoDWxk5fTSYMBwP2sK33gkgSzM796
7vEohyKuBPPxYiErSalgAe2PwuqFxLESXA9Cy9IOTCcZLbFTa9Cssq+WPC+3W9DG
bmifO/KzWHS5nlLFlWNNvyZMmVheSZGwo7VRt+6lgHUD5bZbrveiYoqt03Z5NJB8
JEw/Fo5wkBAv2yx1BWF0fTlPbKxQao1T82XaU49ekawyc7X5o2QUyuA+MAxqh6/z
/TLgKzi9rK6C2QNqKJo+WF0bFNT4uS2D2TagxO58NXBq8XQftHl0vyljwSuTS5yZ
tnfdasecwyTrdroY5NsJX9XcrT81myYbyP4K1E59D08MeGdVGlLj+rOshtCcS6dN
gOVjYeNzNhoNK4Ym13AxBHERkaVJt16EpMquWiBVE4SszYLhyZwP1103cfy9x20o
nG4eQIdKirmQaD76BbyaPEvp2pM6jY3Yn5FJfG4NAr1yXxETURyk2mop+oqEdP8S
IBUSriDkiScrOhxrOj7kCnwy/89FTaArkT9a4c0reaxJoWocwXCODvow2MOeUnum
WDaPVy0Q4bJtjzMEiY4nYqUjAp6PNo0A2bQwiz1Q5y58ZZNrDeRaE0DXTGbuvKdj
Zssv8glNKjBXIINRK5KGdHK/bR26SCrWQsVJ7WzYFqKkFKAZzGtqGL9gy3CzLJXM
tcMb6d7q7cN7WzsLUdc2VQTDLInIxTHIxVbzJB6bQinW+Mf5f7pWZYCoiGkk0faQ
Cc6DroCu4x6nJVEI5OkYD/CCpayEbkxw4pTGBh8SdCDHw2FUW7TliCUEaCYS0c3y
CDhqIItKIEwDQnvUrCCJFuuHNcMRW3elfPDGU/8yvQPW9HuGMiq7z0RShxe1iPNB
dCVAbB3h+/mhuKP8OnP2vnYVnEq4hJkCsVBWYHYUslo2YyhMLgIYwh9EsH0/XxKD
Iya4NkSYboSmlyTtBs4chnjCQgPr7vS2BDHgytay+AUhIRnfBwFez/oM2NagiHeE
CraQWRt4dKopvcUZ5T476Os/a5x6nNZdr3/JVA1NYPKYV4u1qwOrRwiZ0ONMGG5+
cw1JdrCSgXW/GttTF8lQD+1JXhvBS9QiU7RtiI37v2uvJ9JW4bpRiupKEC23isR2
HhsNQieQo8UmqpcTC4N7+sWl0iPxpuKKcQV2boQ+UruyUSuDQY2oxp59xESQF9Md
gCKdPrVGm2LGtEgi2Pb/fSH3SgTkOK7Yt/y7lvVOHq6VM36cHVQ9ab2QMRKYnj1l
Tv0hchVppdktEHbl+sMtJZhv0Sm5LvK2B/FjrAlwqW8e5WGUMeHEHFv/346S51sI
qoByaUp6NjGiepCKD1Srpo/zEyQ7vayRuHHPnbyRLEzqYfQGgMOZl4fIOtCtZpGY
c9xXb8/HNwoz+YUYz1CWsOQs3UzE6zsTGLkCJqo0JwbBAWzIOS8LMOSsachdZwDF
us69/NDXhzUnCmYtPFaaours5SaicfZ139r6ASSVaEVHhvClCxg0dcX5fZs513Xo
k9S7ugMnda4Y+DqAtQvPWHP3WH+snPY22SYg9KDjYIQF/my1ciJ7CwtB5Gtec85U
mdBYrtCIXiOH+xelzFPZa9aKtAIgZWloioD1e+C9D3EoUcySXoTYWmjzNK0n6srF
vUb4OptRRiuRvLfXAR08R1HNs46ZflZ23XIb5Hm7LtHJqJHLz+a3VNHeh2qSxzJV
MO+9uZwbMfywIG/1uI1BeELPaB/sOfwtq9afeEJ4IUHzfIQxvxyHlGeH3mQpZxfi
gLKLc4L1b/+DHBZpz+QhdHwBVFC1ItqrBRay2Z9rySOHV+ioci9MNtbOhAIVsXW1
c9uqwrxCDa4ukW0wM+2LOoK43495LSJB6NfNgN+3+5arwmMOBkYyVKbhaxKzLJ6y
UXa7NtCkxuC9OPwOFETDskFdp60C9H9778j5rtEyFh/ODAkEQxlayVav51MOHoSZ
lfBg5vhuleIB/1LMZYAcpdJLuuAt4xXl/5z+Wbq2KNDX+sinifJZTpCK564J6TGq
d0NsVLZF97xvfdQmIuqBDq6Ve90vi09xonIGl4JVJ4xVAqHymgvhERkUv7FFEd9E
Clec7zBMfXwsSvUB64+BasLIZCFajoejCAoJjT5HeMEh5qOF7DRHw9DBrvJijgqr
U7UPFrJj7ALCCJzQZ/dS35s4qqGPlrWI0dwFYCvZf5hTL5RVdlb1Q5dxbKa/LiqN
zs5ZDI8M2Zy1iO53pPLnmPbPz/T20GfhUUUqEICpfixc0LrGWHYZcgAxx/hMxYqO
JJbrOpJwTYQ56o8aJur1Fu//OiRwpzEeIuYU8S2+ZmtUOjfYM3bgq5TGQuBFIJpG
0BYRXyPFo6KdwT6+VJ4LdVb2wh1JWJb6bHEksi2/k1+0fOa7yUkR0TouP4d6f1xg
/lhufdpt+yPQx5bIPNDlLeIFs7hc5szANoGtCnwcVXsVDePXTvn+3JFqN+mKAF8G
aa3DLDvSLnREbzEgiI8xm9Ss4m9iH4EeOTxEW02rkQvBq+EM+wKhvP31lvjCshUR
jz7Wnsjj1hU5kkbL6R3xcpB96br+jCnwXIIz5q3TKPtqoFjh+qvwG2zawMEtksJ4
g+P5R/Dv22Z9FG5iee9c5uDO9v8hgE9ZqxJ/f4D0+OokAF6W5zLTRLwT72WTLyLM
LrtA2e8DIUF/5CpQ15Vx/v6oBYkgOaN8DKc7zMlBnv+2X1YHqqgX+8+Iotmmthj7
89sqDJUPzFE+FnxLVJNv41m5fiT09nS8DIVbiGTEzX8+FySUmqMOilFGYIuR+OMA
ed5DXKvRCZ8AOBXJJ8s9mvBqmMtmcWe9BtWJoEwlezlveQvnxdt6jAcR9VOa59Us
kvWv8Iqr7XqYK582nTc75ChqwxXyKQOD9UsmSyY4GltYDmPNXVsPntuuLQIDehF0
NJ+AVEtBtoLUSHu22dJhUgFDwB4wWUObC4lNNGHrsFft5LgWF+z4za/PE670Wir/
wO0c9m9M7Am5fFFVZS5m+pzt638ry1Lecwyt5kMSfjl+T4+WIEZjRBLut3fao5W2
7OU6D4rOqbcV9YkI0cUODSgDR4P5EztVd+CubxORv+DdAAswRSTImlT8mv1l9TM/
I3gPU4u+VWYOGarPCF1Jd2dZd5vYJGrVlEPB7tdGD+23BMXFMzzB2WgnIU35nzdG
tXnNLM1gqJhkEB0MxvLTP1rGEhL4rdQrv3MLFTnpEqg5QoIkeYMjRMw4stGc8TSx
1BTDq8jU35Be1kJEXo6yNlFPq/vc+wnD7ri5V4+Y9fNFuhyprs7QUlif9K8SKmsW
bwr98jPwvVVzIKnDfWef1JF+o+MK8OsrL8sj/eycWGCfvKAZ2asNxIXgdlH3U3uI
kXLN050vi+8/eVUfLwBZYjpXkoemeiMv7hdSXMreFYrovIBjAqXck4BfxZIQpgnQ
rdH6tDF1Waf703kgpLoGF/YFQ+C/V7e9Zd6JZWnpegWuXfOEO2M8RShKKuFrcU+Z
XxdA5aZgpDwDOnDTOGqhuPJ/l++PDKXLklfOi96v2oO/FRksirBp9O1fOKfheRzG
+4bO3ScvXIztsANC3Oo6q3sM0voZwNoAYTJyQLPs7yl7C17kjhF46JFCTCu7V6d2
E7HZcC0aQrWz6qQnnrhnBUOHssJinCqoPsWT2HuqFS17QGxCb9R6diVcG25948WC
4H7RvRYOW3NDMcLm4vC7TGqEHfwjnvvSK0ZJLtQ39bgWuX2B12YT7Y1nz2pfDQgr
6rbYAoTGr2WATPy2GI55gI87EFEVPoexLbiqpF6AH5WAzVZj0wXXQYreBN+OC09v
TuEy3uK89po8rIX3DItE0T+3rQr1KYaG+k+vAdoQmmiiiQkx8wyPdrf3WRMA3ejJ
wh4n9Ag4F+Rk4dxcknC9tPAAn2+6xqdmqCXlWubOLXzh9zaAdIMBN0Fl6ifwuupm
9rCx/RD+9oTYuYjWLAryyNitha8/gUrCnaupu2AlzC0WBoY283ckYF2Edp5ulDTR
GaXm487r3qotoV3S5rr+Ubjp2gh+oqAjxS00GhNNzj1PdSdBfBl/OTDvSipGQepV
uf06UaIkLj/iwUeaVw/AQ+y40PMgxbyybiBGR4GcP+aldB8Jox2voqMUa3qOUZcv
6+T0Q3f9nrQ0b1vhHhydm0Gqtc9iaB0BKkKJ00nELanYapUJ12rNCpaExoXl8i4P
YMSbCTfFGtvygFJ30VP+AKg2oBhX3jwggWG5i89FffSuBRpyG7hN5WzgUs6ntN9E
e5L+229ZmC75asENOzWiKqNkmCIMAq7NZDyeE8cbPkryEk9hx3isTrFTWYatDQkO
RpEWwcAly460UcZqDpvhofz8nv0QyhB2NYsveP4ZnrW3f2MkbLSikJ3Hs0F8xHZx
fHcUC6L5yrDXXZU0mvepOnKY1SjWAYAmKZa+WCm+I03E9rDp4rl3CEx4lz4YoEPn
/blGlGYfp5MYBkaPSHJzBY2JopHC+/GCSa97OBvoIiMqLppISplCpxBCWX/OgSl3
MB0k5VyDxSh3UWNkw1S/bW5fnPbex+E7+l4P8tMU2zzitdXdy3ByDSCeCKl/6ODL
QalHT+lDST+55m8UvgX04LqfARhWgNKU4RJ4FHDGebQztuXyuFj8TWqVP7CpHtz1
WfV5QGt3g940UCP/KdSF/EL3n5fKhPiXG/4XInZZgyIkPwk+74pQ7IayJ74zHQeZ
kinR0SkywTM7yLlUhwVfjJn2Tvh8pEQO2dt4ajPJUXbXd7qgGO5XTn7NYPjfFvDl
vpCz+xAo0+JfCa3UgmfxsdvGTfD3ypanRS4FublWkYThkwgKhZGjXm8G6OKIqk1K
SEQvkONUef1SxEvSQO9GQh5plqPPj/Vy+/haJA4MO/B0A8Ha++2ZYclJ8ljRRdgm
sLElGgAvp6zdl2SECwb+0hZAkrAHWphyYcmLW96FA8IJAObzu3E9I/eFgma8NY3s
91lhuryUCxFuYrYEvzm4ljPosiY4b2IMIN186sZe4Isdx4LmBnA0E9rAdWoSfoqi
dD0FxCiqd6h5gBd6hbp4dFN6wodNCuf83CoPuuaMm1hCHD2XMp1GbjJKG1wytxqU
9dF9LknbgRMqqQpv/pwB9g58GQwknMfKu6i/q3zvq6eZxLXvoYcZVrX42cbnsmip
4ZggUtrWZt/FG/4ZJ5Kwu0rd+2ks6F00KnIEpjcQboN5lX5PgPlzY2l40yDI/Zz+
6WaB85JqbugMFZ9+x1Cmw9mSGG6wi7QYphUVndsJNgepA91jnm2/pqunErC/Diuu
p6BojUJEl0xL2v2lW8apNiZo0lDk11VN2T/UEj3ScgOgOiBCxTWU2EHnr2kdeHbh
g621u765I0E4WGByVfwVb1f407ygz3MKWjlUXFr7kez29zuX+/bVW/2HuaWuXXa3
TAIWrbykRDzYhCYPBEMDDaqIVJ/FywVTw9ErMfhhfVuPWBeTAHuPZgKMYkC0hYfx
rTTNGXZ6zUWw1KcfpVYjUll2pclJMkGllvtjmzXSPlnLi7TVRYL8P6n8SkI/wmI/
wleY+O22kk2I6b1ekcE3lDSlirh+TfEpLJ1vtLVEdaDrPw5kBnrUFmfFrjSZRJ0u
Y+zZ9m7VrWnUqr31SRqbcOuBBwlkEpCoB9ySY/zD+nqCoxRpwz+PvLxaMAP37mHx
OwfjOJRhHzDghQOcUXcNXbZDDeCFe3a66flBTnMDeTQWTOIhkWcwyfNCQihQY+Zm
J0Hg50dQR0IgwDZ23BxelABwOo6+5ezC/lsPfWnPaab//2HLMw3ILud7H2I0CEyI
rEqbH8Tl33RHGn4C9k83d1XAHi1UP5L6cO09DCTBQyfBockSPPdUoDCJ6FjnknN5
oCXtxBzDe+0nJKF+nv2R5SHvzdWUjFWwJc1NWrUuMrIi7n3IKt5MrERmZQ8+q8WG
UT3tAoOOO5K9IUEpIOum0HH0O7/qGtQjVSzWJMemZlZeKtOxiZmpyCgLke/bFDbo
FLEQD/phIqA9uTUybfic1Mpx81RCA3jDqcgpRoEiogOwSYzaMBhvFsxRlaSTjx5B
eKWumpb6oxNAnB5v4ZTPfOrY7AW7bBd6Y7Hmfx3yEtY0WXuhzjAunOzqpSBmDf+o
NZGIaGEY4W4+mQNdooinNtXyPC1GiZ5nO88XrPfcg1bdua8CJ2CEfQVqr76z94n6
DbfNIqU4ABe7zhQNDmI1QuFioYi+2HAeyVESj3bJfT3TddKeRcyy8Dmk/t03lwDz
1pQJCDKM4pPDm0dAGpLZWtqos243dsDeVY8t1LcIEhTgXtlikJJSGs5MyQVsgDYx
UgzLIRlqt/UvxOYubhF7hlMjQ8X/NtZ09KpTb1xRCh53/JUczECgMa2T+v9L0bPZ
cS4Qn74Ol3gEDfliOtmvV6/fcsafIi7ERIuTDSw3gk2pj8AzGJDt4CzlUCAq4/AS
Q1dmkJEYPrXYilEAAjXfTM2Cub0PrgRCL3Eg8DsvRJkFRJ1KFAzeS1OVqFszaTOa
LfZEp0b5M8cXFRxe4YDjbyJsTr/97FZM+5nGGm744iRS4NXzTzy1utCjcYrCmEDq
zO6avxUMB6YeC0aitoh9HA2i5D11bf8RGzc1GME7x5lsBR+5ZV2Qx5OLoiF6TCrx
gXvM389O+C7huleNp7A7V7i3pq3wQq2aYV4PqHcLnyZhC9h/6KQran2VB81ckYbI
YqUl6U47dAjj4i2ocuFgPrkUyob91MQJT0wb4LF56kE6Ddb9zfzFfFrH3B6dmSx2
lJQ4DdhFQpfcscZE8VjJo9nGOBt2phSkr5v77WTefSEY3T8vQNwk/JBQVAOM/ZzS
j8lQCtWFyV9gH7RrXj82yE4B3Xo7PoM1O9dcHqYPPMiOU6LxA6dEzm+C4P/kGy5I
wdh+C/AjSEhcMhFNWYQzmnrXjRqzQQp3Qm0v1Qyrtzzsqx+TbnAIrYRAXQISZd1t
pipVHMtNmCARh3O2WmXeTtj62No47N/7NKEoSlV9qEYRSP8XhUHpLpVNr/lNgwSA
SuF9arECzInGq7RCjMv8PFWD3oW9k3qF6jPJLSdCmiWO7sBJqVixY/1J/sMd4DWd
ICyv6NdvhN39/2NmWfM+ATBgKwqORujffPd7/2AwpTAfJUslZ7ZXtncGzzIJga/Y
m+hXqm0hM4j2zwtNCYkEpZT+QpFkEd0gWh1bVVUW91yep1xqJKeuhnyTRzKh2ejc
ApEdm4yNnViCRxzWTsW2eemyw9Qtq6NJ/mO04sJQ+jw1BZKXKEcOuS/voR2E6lfv
Trf+6QdQbMa2T2jF21eFU90XXH9iVKsujb2uXpVbvrso9RxKFxbmXjJIt9gZZpT2
5JjIWJZKpgAUUAZfKRfjKWj1bHMFYPUOAmCOe/IdUiFhDIQQeGU4auYofv4nhID6
+2GZq/kEQf/u68khHbD864RAOmmD7VDu3O143CsmZufFIfbL0cleL3gLFyZsLTQU
XBNW3Lh+oeFwDdiEtWrFFVrOWWAVqxIsxUmIAkv8GleEpa58x2H5osdLjRi8j1qJ
+o6nXjmeD1hX2BOZZKbo65Ew/+1uWBXRshmM7C5ZH1XBqJyxR9PvHbwGOLTsOpQG
FipKPQz1yHGOBAHNiCflJEaNEUtx1n0MjHXbfjrubpe9letpBCadCaVQzU3a7BZ1
AnQhhHWKXT+H/5dWFN5qPu9pIbsgCXtSk9Jx6Mfpp3yUnemjfBPLTXh4WBn6O1Bl
MpE+7OcF+B/uRBCctqYJCCJ5BRzEwrvxp5rd0cl/oSMDJd7gxFUNmuq4PKrbREza
4b0UFMccEoFZzI1WxsyorpztuFS61bjCRDtBjtYEfrLP8+6cdKDHKafAavsllowq
/7ggnfwxnF8/yQrPVFGh1W/ia5sTYTRJ5qyoJvPyKmxbZGC5f8wVpDIEPZF6mo5k
BXMK1Nj7oiirX9CXLuzxVnmd2s7Gh9oLO4begQ/JH1dUtMsX+8z1xFoeIAVvn7Pj
BZ0GQniRBroh6q7SmijVuQSdwM5W0/CR7QzApSutn+gkN3R79Jll1xIxWgTA4txd
7UF5gyFMToieBr3kXUPTZf16PcBAzOLabY8/JQNOoOsp8dDue/erPXwHd4ooOWx+
SoqkwQwtPWcJGI0mBA6yERgCQyyP1F46LF86fkgesb0lKugB3YAvmA7kghPLLxxD
Ja4dUwOXie15tLlkUYAJDghB7veFhWnzT/5OHtxk5YoA0fz6fcx9fdqVVyGcPAti
b6l8SVTBh3SVt3+O//Ci6VWlpWYLT9fOL493w8NREPEa1irW0g5ztEYn2UQh0tMH
4gW0ZsAxrw5I+4KpyNFElxv1lP8SLJIyaGVHHYvnheB5Gcrsr5ycm1w7eiT6lRgW
Ycz2KPu0+ui/bXQaCL1u3OtblV5tz22Sq86TGBMuMeMYTvm28Ijf7p9/A1uJbNcX
xdu7WyONDDNjXYriCgo4FFr8nHGppoiy13DgnunpFDz7kyIdBfbajDwuyMa8M9er
ng/kQ8LGjOQb9LgDc37bApgPr+gOWYOX3EYqrsGpXjzqIDgMekiyHi/y6KgKEhk0
tr+EpuNahtUDoNcqyS9/VNPd5xgZaIaxNmlQyNVlzsvZfSicYFo5wLUd8pDXNTWC
UVMWP2JnLnxoZFNieF4Tjov++VuSeVDaxFYiDgs08RVBodd0regSC5KLEdEYOUer
TahXLag+bKoZTyqiqfEANvyTNUZsdt9T5krh6zykJR6EV/YEeIl8wMCx7PV7DwF1
cZkR76pG166IxVB8H1Pb8SNW6jfWRF1i69rCEWHsqsE5ivOB56S8pbtSSPkdUBXS
/rEjmLPgrRrA1Ov+9JPeahWFx+uFcSRmOEkiRsjcI7Q4l9bV8OaI4yWdKYILMkIC
5mqq+1troBiKKsjTciWF6aHzvLWQNrkEsZbzd2MS0FWeBY+0vZPHz6gSJv+JNqCs
rmor5I0gmGGfK+XhzRrJ0Uhr1MJ/RMvQYPV9OymIZyyNHRI5RsbyMMqKtBEx44a/
SvNF6Y3+v5JYzZ/dI3WdX6jLwqZdZlOwXvUAQ4WTTsh6WQ7928fG469m5WyfGBgZ
zxlQGUDEIHPTjKcLr/Z4XR6cWEct8VJ7Vjys2e5QDLp+q09Sfded19Mb+Zta83O1
YyNUTlAvGgIurNS08djeSiaWbbNni7USoohvqHx/IfUJtFdYm05iuKDwUT+lq7HQ
zi/iUWhYOAeqHp3NCzpYEZr+PfqKpAbyCB2Pg9TPlfpub53N3uwlIoTkAuXT3u3N
qtzDK4wxml+dW2O8fLSrnfkO05f0BpOiHMfFoyLjBgzBym3Hx3EzW4+6/ZGzs8sn
4Ib1gY72Gr3NB1M/K078ylzEu9vNswVcCL4sncdP2ci7ESFWBlj6kFQLL8pNlppf
Saa0UnCNE1DSblYDnju6DDMqyDWOsIDlHSK2Uh4n1HIIf+arp/U7yCRWTW6Vhf3b
IUW5oyvRMIQezz4q3o54Ebw+j/DRtxN9dFGq+uW1Jbe6+pkDfsRc56fPNYFuG4aA
CgVnZP2OYKWbShJ7JtIhO5gHhcNRAPMqDJirIYiPHaKkxjJKFpehvqnBCCqCIA8P
rTr0BIBxeVu8/rYvoVXHqaLJ3kFcVajptVcW7ifcoDA+VWiaDMfYk4mOGIU8urqI
tW/ZkoBMcwvdhlq4NNKCbcvj/D6DUc0KSODM1hyb96WAx6bDQ8w1oTXVAjov/e4p
fnp5Y9GHJ9SpAnRco92/rduYeQeju0hT9eJ2VL1B6xmxwsQcIHHitCPcPmOl75iu
yYb08B91LVhK5LxqisD0Ub6zhmeRFFr6TUuo8a8EfCkTrff6ePbtsOO7iGZjqBwI
phRIl8JXSKE5hOwwcNR9PE+h1duUxAihfUvOJ/UZ88AxLVDIMPXKO/6n1MsurpqT
VVb56c1DQ/3NHCqgSpFrKzg1xhpHArpjQYrmBQ9yA9FIg1m0D/vuE5RjIROTO4y+
0QYcWlOF9nspNYG4LmlRlTtGy3CASMztVzP4kiNqJDweZBWpiqa5Vwcs6yfLslan
XtyUwkIYSRbBBTwJi94rj5Sf5p3OUXhYPXQRErhSxQEj3kDLSmGb+YCj/cnSVi9z
Bf5HbpsCnMHwSvetcI7lsy5KfB4i1Bpx8VAGyK8qc+EAMGrrx12NCxwzdmIOeRp4
jjC/WUT+GYyrmzZTpUf4JJBRaTcWzH+o5bbVUayxeuIT+K4iml4mvLzv2n5UahFe
ykSlc9kIgFYftXGlA5arQmm9Z6wiE08lJqEIyTx02AQ4USbLxZDyk1IePQYWeHIp
ioFm+L5s9uPCcBt9veVRxgUR5kno50sOaZpdWTx0s9l15cbGqJaHb1go8RU6YNEX
ym92viQFpfJosSvuTc9FevK+VFKawHVrGO66mFBxwjPregT66IlE4AB45rO5DrCc
AirE0dDb38d1MtjF1VefkoxZfDFIfRwjQL9LdznRKesZaw+0ezMjI0H6PWtFVHfr
Fwv+4yMFZfhKmhqyj0a9Wx1i9PGCakAwCdfiSNC3xEsUBfPjUyK8NSRxhkTg37xq
3p+lIXg2egUuh6t4SlFbUFWxpdbOffqZjDYfryU1UorNYWOYNLL4R61oH7+2vNvR
eZ3GsweTJphQ/IPIuKlyIYIGlMQfj8MCMIbgqODussRC3BMt7ew52FRVRegr09g3
NzqTd9NlylezbFg0sdwLVu7TxmPugwUrzkr8Ri24pVDOJYMOpd3R4ui6f0WSAepJ
9n6hWp+KKPdb1jSCr5V6FAOXYGOkkJgPYixBK+cGI3gnR6QAVr5xD6MPubOnzq4m
Fro6FQezEVfHfxctg523giQf45uBqZUgghl4PzRqZaGCr5J9oNsMj2shepKkP1uV
b4bEqb5+P0LULu87BiK83+nZQacLQuzegZvb2aDpHIYxFkoVS0hhn9+E78avXuoO
5NHHQ0cSLT/ilZWPnB1UtwAKJJMap9L1BajBTioOyrFdGrZS0aP4F0zXwQLKcBeM
tVS1XyduHEvSs7htDMo/SggMealgQgznpL84V5GnSCF+FiX5sSZPN6ZVU1dXksDo
tPTmh/alAE03Qu2ZKd3vZlOA/cdO3cHKkYTkNZY8g1YyPtjmSCc95i6uC1JY+6RC
wBARmfo+Fh4IH65nGwSJdQ9V2/7Jbv0LRVbeLt+hyoKkUnqaqTqkZ7NAiVhHf22w
lY699xWxfV95C3nT+miMB/H1QGCOi2vAarm+yTb0neAi1kmsfeBQILKeBe8uTtOA
Tgv6r9dWE6MLdkiNU2uenzep/8rD3gZQILr28jU9t4PaPzD9ONoxHxmBKvHyonDh
9dRtOvCxb0XnaV+MGkuoOwXYH+17USWv2zpmuBflF2fymVR4k753BsbNc7kNna+9
cI0rbQP3IE1lDLYzvbAF2qIGdNsPXjcoegnrSuGvl8WAkcpQGftwPjBjY0+4zgrY
ndbPlQRMLKJt1WjirjqtWpponfn93kNmHlJzFLuGte51TkKHEBOR23M6NleQV4Qc
ZR9ON6F8pF5IC2HjzECuD5AYgjR//iPJObqVMYSrveY6X/ij0tYq3Dcqm/CQqoI+
bNMxd3hAFeQGH8PemNXImv6vbuH4dbmqnodhHT67p8NKzXSuj7MPYbbfvLZiXwju
OBEXgZH0IS42KosbulKk53nITyXIQ89TlTHOGZSqYKabTvxMVnTWZgy43mU72UWs
c0yCVUUDO/w4XPwJQ/BfswvdVCTb63Mov19I9K77rHVC/nhJ8hgMkiI0wzYXU+iS
KGzISYYMdSZzQaBNSIScsWI/PfyvGFfDmVxHjcv4ibpHNuYjgViJuS0VKNMXAVRn
VCcI8KHJD6VKv4ZxAoJsr8ayOtpHrlEctKLNZMVGZFYPHN0VJ33zWa7xabJfmgJZ
Ymq5kQ+yMzsij7GPG0L1XQtqIue1xVV6ixhUIexpvcHBSdlSwtszPn8nuUP0F6/m
vsfs7NbpRU+cXRe1f3OcDiXSJqfgxqNwbTfs4AhcnoT0DWQsHV78ieISe3oImqYF
Rq1TSIMHbCrGKdO4Wi6/i7tbTPQEqVk+FnWsLVS1tHBEHFqeLuu2mbkm6szchCa/
EtBTQb8RWpjrHYnsEPXIfgWTAJM70yKUPNeqNklp/Yd1N311z7E+BetBW76lBiJO
Dr5U1OdNKoJceut6dNrZye/X4CD+Kx6/LIowyrZqaKbfX2Pl8F1dC09HhnnuNElT
Z5ilenuwSk0odqh1vtZvqG8fkviht1DqrQZAmyaicSHhR4HiIh21qZkLRXvMBguM
Au+gEdsySNqghxgnRmhaJ8cWzEQr0wNQYp3zCIEB2FHaIxvdB6sJ1ArJZSJUg8At
j238KgvUKNCj8nz1ZZuRnYbyLgIYPUBpTLC7TG2Dnvs4PGPkZbzJRDglgvP8Cgaj
OqpgwKmyWtBko4ML0phW9WwD1Mrd9brs1tXdDEQtnH8+6h6J3hRFMYL0/AkdvRwH
piwIsPbFULIjSemeCDAPgsym+VhO1AkalXoxERlNyoflf812665c/6x1+CqTAK9H
W2WtRPM3C//Y0X6X5HL5VRTw4iweTI04FAS2z41RV/vncYksjPNcDnQIjS8DCczy
USCo2jfr3xiDH/DEErzcxk8nd2P/WjGtuw05UQOa2CNdGTury+Dp6eCG6vS9aKiC
C0oa+7s8ZujJOCeZynqRdgUuH1LzKNCGPji/20Si9d02EAMkSty/C2ShlBBDpbQd
Dq0YNOSH38kLsbmsjgbpeUJMBRvTQpLPs1W2DssDGKT7ZN3f78VYsD5h7yeVXJ0x
Ye6+pL8trZ+ZzVax7Uex+ribut1GxAr7Y6lTxGyIp+Tz5plh798u44DHBTQ4pZ+o
LrjeIcpzIrvMNHqKiLK+MHz8hGwoKNEDRoqNUY9qIxl+b8wCUWAa0zi3nEDIhxVm
sqrj7dB5nzbHYw5UpkUFFSrSmeJJHEcs1O/7agmXrQfHMH5QT59Eupa4jm5ZWy4M
FE4JPb4AD7aK8cjTKxhpCmmzMXWI3sGrjmqaADGEJoH4it8hycHxnwfzF5XPlAhN
3iktitCpeob/5vglT4svrH/rX3QkBZL1zIruy1Pt9APRm9iuvSDUpz++ViAdqUeO
dVC7TofpELumpQ+BJG1hZgrmyM2/ScDxxqi0+iszf6piarQv7owSmAEii2K3OlyX
hSIPdC67ZmEY3fJRY8lr9HcWLNklZLwN7ZypssrJYpR345S9x1jPGT9BgJEMog5V
pm2pQyn/3Dub2TEeEQDMiLAQDDtSmozbEtMOV5Og1dIF0bz+DG+Vpz/etqmADxKd
+zytYxopX5FbG+UzlbXL7W8SyI6wOqfDgiGwKCilE8xVn1wUu69pH9SATW5G2BEt
FPFe14CpeoWRugeedBsLfxVbgT+LkDdvzL26PsRss6f+t488zFsc6y+Ghzh2kogO
AwQ9GJeOiSrZietVztQG+mLomjLS34yvjHGLuMks/W5jptHa7689gySXnCwSPJx4
SuE495j5zkU+f2OPDThKYP4ctkybz8BIHbGlopMGIMeMu3OhOOPtzZmbVx2JO8J+
McVe53nwB7udh7J4jjcPtc+LZC4XHJhULrk9tNpPyjs1VpMmUs2mVMn7DosvBO0R
xzg4peuO1PASnZU6JLmGuYfNijB52alWc/VVOfuJu8AKe7xToQpLdZJmkrFdY5xa
ElHAszcVOJBKGPHkrzm3z/TIgcBSOw+pTSqgVFHPs44zUbjnfJkg5vncUR9MbX59
JETeyd67E4KodJth8kog8cJ2qBd6610vd+6zgEsYYmVxlB8e5HIOfd3pifPTroUg
wREWcHHOCcVGE7Bq2EgdXv/avgMFUqOIffiRaAazWiZ1AiPC+TJxBSl+iJbbbFu9
Kma7YbTAlqI6GYQ4BKO7g2FMBi1t91n30xfKYO6qisLyRbuVDf5Ly+kEL4kaU28b
GBjgJKrot0UIt8/U/MaCVMuVNd2l1g2GTOsLWPABckJp4mGseZtGHSvs0nqUdyzc
3MNus7cjGEcEgL20QNCtBIQYoMULW1L9HMhrn1xmRRSz5nZQc9cOOFuhInNLIUnj
Bm0/Z3i2+OyUB0hXA3cjwy1E9pvnHLHYvHf4EZNoWOcpDrWKazw1x89muIeNB6R+
2ciSm0J9lMYcSNI2DvcA6zzF635h9hyaJQduVOdG8uLL0z4W3sHoWDsNtQ3g+9YX
x57rtomSrnhvVW/khymv+UeANxu0aaCwQXzoTqUO2kR6zQea9iD12djFe4vku/6b
0gH33S/C96UQAXeYtDbF4eEpuyurwUYEU6N/FxXqhP/tFUgoQejeoSo/KVmTwos/
afx6DlGFM+T9z3NYzTZwHmYd/15E6DTMUpSSJGMmS/pt5fJHWRCnFd+Rntq4PNAR
rW6kXI/oZgSdZ6Co/HLqV3ObLClKAhAy1vso3HIqTHD4AyxDRGMTP+cuBrvPEIfW
BV4++zBHTI5yt4VJJR16hHDJyI7OuEXDzGJp0cXGTVFZaBIcdiN3/asBliM+wU4U
7jXaXtlexs477Xg0f+Hxw714QHXRtQ3GCVfybYIy7lT4RXFPnOTzFaRS8iXCOjvd
X5VvXG2cnQ1S/Nc2yPpYCDsVFqL5+KLYhzECaS0DC74vS715a++rrG8RR8uui+lF
QzR3HxQ1KlyVc22AFc+P/FLPfwhC6q5T3mNnjfTSqC3DAP7q1iTZP1ir2IGw4CnZ
jv+5t/I5imNVKoWh3j/xgNajy1jqQikB/nV5QJLFP4NRi4rchQ9mj0jh4QK268BE
EKywC2J76qGrJihFtE4LXG2vZFTZ5pTvyAxZUVp7y0GOVzPjCrYLNEavohHnjiXM
GCq8akP0dl25idOTlIBsITJnVBi9TEX4CIErPQmkxnepH28zn6VOIRfr70OpuAaL
l6UBDB5JqBnLHYDjOhZexaDpfuNe2ggQWl7srmF+wzV/x8YRrH8ZDgUwd78P0Nf7
V5Umoc+MR3grpOYTMm6SaqcZM+75BRUUPpd5x1bwpGzt7R+gFIN5DozocnrziNAX
lWzZXUBqmskOVOSoYus40QTWw1AUG1lrL86rbozZLH+jK0wPoi8jh3O6jEAksav7
JXFFZEyF+41rE7/Qas5cCUx45t3r2+YZIf1ttltrIVruX++I/zIJeERq227rmZJ+
xemNEVkCtmUoYLxehnZFPQP2vgTu3aN5zLea5YZ7mZi1nhPDvQBFgEUqyCkFqFpZ
PZ1Oc2mOhrOSUvEbABlbT4iw4xNtu6KQkyH4YkVMackWh8e7i0Pw0/SxbawB6V9E
u/Wwbb2IhevO1rxhQvKVPJmac8Hrb3WamSbMHEolmNqJUm3rBKJ7IFsQViZg2Jah
FpZ69SkGOWfmsy5yT05zrCBhD78GxuHptr7xIcyDNb5oLKKKIscKjIn/5AnNY++Z
HcOG1IBkFaTflUVe0tLmS1WUwPHQvvJqGYizqwp9rjgluk2DmWI1oqoyvcu5Km8s
gMzTo9m4IbEKk52SedX1tRBJl3ht3Paoo5trQwch9KILk+EdiRdvh1d/SOue6Z9+
TqiwXooy1jYTGtrx1v28WW1L8ThFOeFZuRcyzXue0ANvTq0YT1fB8Jfh0jmG180g
MXJJuYxbICJ3gOSrhu7ks0q4+4EKoAKp1CjUllc7Yx0K5f+yhmkLm7sDWIBa6gM6
ef9V6Aq1SGD5LAo34WmiLUWXh76iZ7zEr+H8QA4cUAL9G/joNePidQ8OR+SFKRMO
TuQrFGJc+3INqzYZOjhFu5Fbqf9KMjOXFYp+HTL3FauZPLBKz2etX0nbEdaCsOUe
YeBjKoQLMxQs3FYcoT7hDh+geX9KetuuWUNQJO46ZSwsun84iIcEZPp5BfnZklYj
yKQ9Ogu1I1XJOYhVVKBAVmwdVqpyVHGD5VkPbX9gDcbhkdDMTKNj2cBNa5j7Bfcw
LFOphlgTn+cV2f2M7uY0LisByChhUDWxgSh3zYiEaLg6wNlcfzKEcqdCDcnxAn+D
5VB69er6T7QeXsBunMErTXI3Vc4kIDZtdMU+DPWLI4XGfJlWMf2qCPNK6k8qXIHK
v4RxKZtDY8NPCJBAu9TVWIeeH7j+DmMvg0Sbk6VS/4FSgzdXhjyaQGZJwh3HBUtV
kLrL2fls9ses/nQPlJNWtONEU1BAd4wfwOW5HTz0+HhS9LnsYmogOUtUewfLgI8N
RUVvB3VHcMv6T0zPaVQDA9zRfNl8myyv+r05sBZnYIir9Dtn3JthsRG0sb2VzCnD
Y2oDtXQrg8x6xtiY6gJjqQKTfPuRu6LyBYyIf+aM+O+bKe10PEPb0OrnicAwf53v
Wgx0A/OanyokKzpTrNKXn3hHncB4VAOWLn921CBLpuSkHk0rwiPZxRAS8XOJrSJV
xHnz4ostHNn+XdKphTyTKFzwLrW4BoL3exIFhUx87ke6yxX1xAmP/gHj0EKCiP81
zdBNuOwW8Dv37d5fuI6AJ+3uEJ8Rb/hQuDD2d4vuTr1uxWJ15t9hjHj69a0r3scw
BPJY7gezmJ3P7is9xxIaKE0iiZZsz0durV5yjd3vRfjopnoN8FQKmH0Np87Nc8b6
mM0Mrxuc4UjE3xn9zXy4XhCEiXaiwLpPyiN7UlvzgoPsR5Uslfe6+q3qX01H7Mgw
osDdKlnNhfuvtDB8avAkW/3LYQM2BS2JUJblSOD1leP2PK7j3quXc7/KOIzTXSjt
kcg+U53psffUX9mhNbyOJ2NhIJcr9fmMZfzPucvkQL1uFu8xF38QP4i+cTAvTgOu
WTLTnPXo3if6ZxEJKq/N3amgR1ZyKpJ+PJ0x+HM/AduWXr67EX9LpNdfUSyQJkB9
J4S5EkPY9Kec5FxDNAEY6aZEKSRhowR8I31/AuMX2H5gXO46wStl0pu9y555iD+j
gO5VJoGzifiJZUOeyJy+Ug/xqSv4UV/tzpwgdGPT9zzWefW2TgzOxMYFOWFuY+KJ
yRKCKJLeUIhg6KLsS/4xsE32/1yqlKk90aojGGVaq/ARLyKPAdbiTGi4gclutJUc
J1WAK1BbmRoFto7XZNlG7W89zrlg1eyxKsyXn7KoTDnu3cw8/oPDbogmvx5Jk65H
12Yrpb86xIxIw3qSxwSZTvg+MAwjb9HpK2cG3cyhfSvb4xEcJs0aNVzt6odRsNNg
nIo04v7RnbNs8WB6WawnfPBKW+5nTTvdojfUKnMLPAZoKfLIWVwSoLTLC0H6hUgR
iRmbq7DHQLEuAvqtAurDAOprqO/drCbv3xv4R3o0fP+O5KQODGuTpIHT7BL//XS4
mvbab5QanWaOiyRC+p8T863BHzGmRLABRBnFGA7ybTJP578CVbWfRKHCsLGkqM6R
mqRLn3Wf4nJnkQwfnD4YDOdr544ARVKZvlcGmOrjkNyLhmg0nsSakMDCaX3bhS48
Urv+lsli7oXJ9QeiCfqsmRAkKSr9F1WCkDH+1RNveddO0z8BR3TDd6QmVmEMgBu9
InLPLERZ4FfVyjj5awTV8iFiRHmsQj/8jcvMj3Ambn7Kaay+jqvhtpNtoqkkCS8J
IMLCDKLBgFy/1KZpOPFyRmn9eVNtLWbWvf3SFhj7LHTUXXDtZn56HkvTgAHXJYz5
BE0g5OKZ9fG0h+MUZVXtblbFqkg8LElZI0ZLRiirSvreZdDOD1qFhjqYKuVpoV6g
zqnaYRYtPoMnUAwmMBz3A9F2MnqWJNiXHgKX1LTRVm9en9gwJFzqJAK1rLaO/FIz
yfVVmra5gnHLm1zbMPPgPc3XhG/PzXOyj8aq3+k+MmETewvVS8odsdzx94FbPepd
9D188gCfu1Ct8Hfu8lBFGqF0GiiCjAkCGHJVk4MTktmo9MzvRQCP8bVH+6zu0ddP
yhKIdQox1EPi7XxKN50hH5OVb5uG7NR7dZR34qG9t4jZNr6Y0EDIGugUr8/ZcbY/
0jAQD+LOTOZGPrFrNcjctJatWMT6dG07Ly8516NoYzhgPBtxyKGe4RTPpguHmKks
ukLsTgft3C8R1bQmoDgfNm0WzwO8pWaAwEXL4z/9TWYuRvXgxRUAvbXooKXumO6y
KHux39UagOLZuy3p9Q3lfqVS800kyol6yO9NEOIhjMwR/qXSFNvPc/QkfS763TtZ
Nv7snNM5U0WH6LGW4gXfRDMM2ryOoAe1lOIzPmYX6to4AxnekzipBVSl2AiZLe/Y
xFTjypXImMPYY3kr0cF2/MoAG7TyDAmSyBS+sIlpavWaq2BfKcWRTEi+2CKeCmqK
U4yByEBhk4j2j6qLCBAEpKq10GkWHMJpvwEM1bl9jMU+tSnNgz/ocjcfZllBrLpv
4UtKzoQ3hLwXifIGtPUy4vET5Cdg57oIfQkPQ9WGExBpqhN1Otp9gbr008e+I5kR
+pb2WgmJbid+zqGPRDQSv9sJiUkA64RX9cKgcMczJb85xHpJSILZXiVxOwy/vB56
cDCcKoQWnfgtqWrU0VxMJrwaojeqW88ugGExJUAro1pX24WNqtGagrsDqULSBwLF
dktJ1pOVWbhEviItjn5c2mzl0msfFiBgev6mP6yQBVCwb6L07hycXAeuM1qhANvi
IqkPvehcGw2qOpwYw4NmiSavzuMuJ2WqJNDkFeYAcFRPX8fmovOszHPNvLWtjzgi
whmnUWuKsHZYdwoAsFi2SlDYX67aYEFDsmMRM4vOqdP1Q5N2vm0+shJ1cvuxaR1m
iXCZ4GEIEQqFm+HOkFcyuL0c3LXFbvnnC1tcVuoguIzRHESxZcxRnhDpMBb7oK5/
O3IMKWx67nKhYOWVZGTawl9D7OriHc1WDDS5BkSW6p0KrLOgPmRFovFXbRZ01R5x
ax6aKaF2DRvk89/McE0CuYkD/pIN1DWw9KgmH3Vy9Uv5I9lIMKqyvg84zi0moQHC
WrTqmuTJU49uKHW+4hPxmpaPRB+5rjDZjzMdNoqWnVR7c9Jg6Qmc2urv96IU6dNq
azbNPDrxio77NAjWI0HKw4G1E+3gQI67mqvgoJ6LU4a3nO8BPzAGwfwWcDpVO9ic
d1kqSjDJnHWkFLCtR6RFIiM05ePowZWqj/Q9BJ+F0Fk7TNwe1skvZqnUBqLk+aw2
4JZhiSl8OsytJXsk2UVx4PeM8Zc5PgVB2kAwn5LdJTOVWaHWQG7Tgh8e6ZnougIJ
y07lh+jlZ7Iu2mJIXl/ccgFh9fsbkwLscOaAWJBVcix3dMOp7xSaq6k7Nuls2cKe
8WSxLekWR1umFS+Fsx3O+QIm7Ua7Zm7zHAgad/aOGRWFov/gPKXJULQhlSO8UJb6
jNC3gkGFohv1VeRmh/n+rX0NS4zhrFVxiVDSWwlLQOzpNouk7kf0SChEP9ef6Dmf
5XiFDOCoROf9+icN3Bfd0XFxotkmoUuDUTshnBGmKf75c2Goe+9Gj2zmXP5GR/5V
Bkpg8OGQU176KMcLAU4hzVaALnRVpwpXkl1SfmcUifAeiuub1bvlEZLApkEA/Gu9
+vxZtLOMeVUy13SVzhbSDhvKm5d1sH6v909mBYY7W0kKgXIf9hY3uoztQrpsNPUy
J667DGJT9MpKmcEMHThic28RrbA/+ZCQg/pyp/R9nHZJFvhYZqhuGMSpHRp6YGw/
K3IAZOejDOk+moDNRC/BlH0LG/rNPauFSITvH5+0txTmn3frqgKQP1WRU12sSWZN
L+nyAf6I0xiR+XQTD0tysj3nsvqKtVaVjPYehaoMdPIP+V3IBxOjgGMYX7txFWyE
R2Pzb2VRJ/7UwlLJvAABqDa7UJqvw4dXsCpb4DIfsKs7aH6AcE2wqWzOwGAYlbaj
Vcbc90E5wmGk170HqQdv5TaKAk7axcBOU5DMrVaNyvNmNG3rL9iFwkj6Kcscj+V5
+WMTPSQwEbgYsMtGq3ZZQ9teJsFr4iQO4hp8icAaff9Al7dYMM6NdGG/bj4otzeB
31/FZvlFTE4qTSTqp5c2Ku4rVwL6Q/GkPn65+uhhmE+qPUCBQDQxV94qheHqSWzJ
fJ8VoulC7FuUZWsTXApQcseIlHhNkAcJ94a6MnbQQ5Wom7b/r8md9UneIMq0/Y6X
5j0aKup8Z5KOeeuau41UdQMV8FHteD7P3un/ZfwKj+VeFqkpKrx6bhrJGrReomDS
fALiIFV496HM+rzMDuNwin+6RZQdRf/F+voKY8icTz4zivAZ0md7889PIdV4FQN0
aDEB+yvnUd4CnJZkUPZpkYPf1khzkHZD6+9kv5oIHTgGidsLUvnXI7zqPNHwCav8
q2fkMXkQrZ6ApLmT5fJASnNvuUXYqby9OyFLSvfwXsGTcocIdL7ExTW0m4/x/fxa
AH+DP0u2NiZl0Pm19Rfnq8dCTfdoOJt4lTKf3L/Kep9PBoz0pX5wYL0pSulSTSfr
86HQPLFhyAITbEWN44xVVnetX+Q8tegYtKxzci1yDI2hVdiL9QIAJK5gG0x0nZse
Xr9PB5F5YWKQG5YIZ03KOZNoXMmV065Lo99628zkywogDYwFtyyRIVtAX8lr5cVf
hoLEmcQ1SP7yibAkKNMjThglGo1SQveESxeXzlCGQJtH3PjLzM0FrU0uKyQrvq/L
t1UrLBt5gUoNEBTM5s8aPFFNTrFum/usNPX8LMWXHfpIBW4UOYujiagPEo9aIVC7
kSy57Gav67rravU54ufoNavt4N3Gpp3+qBOP/NKhNo4MwtZYdBfaAcgmA4UPlRLr
LXby3LqBmciE76k9psFm5er9IZZsAq5cdQRsNJWrmy3EfFKhNXT5vd/9xmvuu4WS
b4VT/S3S+5V+x4t/uW/ccf0EafqFmYyU+cDtJVb/qH7+r7p0YeblBmc8Rktth612
4+mlE9QhWkvrYUSdjiYcU9VtCmC/f6XovNJ73+0ZbFAPyG/FVuTvMaZhQqUxtX0V
YWn36XLSHzvtPbpVHZZkhJQcRmT6SZGTj9oK9UMtFHcW41x75f0FY3575G4dsbzq
cd6tS9/ytvr4zQhiC8sEhzlJgHyXSnrXp22MigwGD3CFskLTW02zk/OUSMJUNq2k
bwM8h1F14rGoUYYOimf4WL1u9sKaTJulXMQFPNWCvhHAEOQHhHFyjBCQd2Z6bY1h
Wq8GF6PZF9uqmVCokRlJnezsr100dN5LZgfD13fjCNd+sjNAZpUrggeT7vS6qF7y
gmja8M6aqPXmBjwyHe45ejG1W/GQjGV72twCBFgWJS6NtKZqkTn0wJfYel/O+qSB
TYZ2RQaMKnpHlrLapy9TIyewnSORRFOpeWqHV4EkHYUVcmeL2WlgXcLFNtc96Pde
i6ton7Mby+LWxx9OpCMTKxPzebKT1efVjcijZb8Yq9c2DsyY1aJTal6IR5cNbRA7
gL4Uz8ENwlpnMTTErI2COHYtALxtAhDuLUxWzX5ZENwmwWqOKQlhuFZqKbPR6k1c
iKKnGF6fG34Ze5C4qTX69Q1UeJphjoH6st2RnDdSwfzoCKPeIJxo2tzf5v4WVNHq
WUTt3m8O7wsO6pHzh1EPlSWqJiYf47el/5zepK/DaH3LA/2XaV8mRSzExE1XCmbj
4oZwEdEgeektyF17z+wUVNeP7T+m+76QDEGDQMCIvbdzdrwxdTyttW8Rj1ClguW2
RGojdWe2UhtzwE2VTBhbsn3CqWZMZj+8XTcnhm+w8s5k6yyZ4WjLuzBfj6VnH5dv
CXRCKlkPYe3ZvXq6qPTFIAzOTW3zrVJ4W3x7p5saMdEJDOtkMlJweLQ5VMf9wPA4
E7hwPy2dSEVohaVLlsEgGOSCw5IhgI2LUr+NANvHBLSEem2jAOTA0XeVHKZ+z0Dq
5teYatEYLTGYXhGsYAF1kDOA2N0oMO0f0FieGXNglIV9ux64a1FsxGNr478UcPQr
oOo+isZh0BAeeg245znNfvdPjbNgYAQSi1g/7K2LR2g0WFpLu/cOylQzVxQ0tnLv
3bjm1/AeAilv5x/DdLnx5jUaDB5rxbWDCxjI95yTmkXEky/V0KUbkpye7bdFgUJZ
SYo43FuKLGvBBLvIjfRYOqmYCijugUA3a7e3g0lJrldqQQid/3ICChQegZGznm4s
MtQhoQSUtwKw+wP7l5ZWgvZIO8vmA6AIDZQfDFJdoVvlsZOqSEjqYupA+o2J3Gtm
zox12Robwpwk7iaqw6qQDwtSnR73AU865C1olgOswsTXRM+Sj/dxrOllq7HpdUOs
1IsNXH/Oqtogrl45QS5NdF7HLoJ/Rp1K14CnrBmyvOdNN8hpfQLo88qjGAr3M68r
NuJ9cBenHGpc3jTghL+iBZxucob2xMIyNBC167B3RMcc7ma+G1oweU82UbzXKO/S
DZvgPBa7qgnuUHB6qUejph2SlJO5v9yV5Syehj2IL90p5zCi34W4pE0aAFIQnCLl
Ze6rOpy1uQ864tnX/1jh483ZVOAdBrXuv9VrAudM0sJQgEE+LKVkYXC5MYlMsxWw
Xkx7qnEP5RJFhxCdRqGST0O0NYtStjtN5ng8xppfUm5X4TEzM0EeyonLQd5p6fid
9ZNfAh8kM3QhaBV1G1T0maq1SGJSX6MLJSa9kdKng0nRdF3+nGeAd9FfaV0e1WUI
ZaRCl6qecp6ALwahJJWvzoNA217HwkcR8421CDPvfi3f5AFByMzi0fiAAVy6dTjX
3iEOpB6SlYzsithLtOSlRC/jXDoyIvNXhFs5a7m6URBWyy2MObn15NN5Bg1Tp2id
IMzCbsOvZQZ64u7Z/otIGWcYSl+CJu5hzkBPrQ4PIYEys3zffTOjempN4SjwxvgN
9iz6tINHlcAFlBoC9UE0oMF2koVs6qGGPnL8WxhgcmQHnXdU0XpSuGLvsM/qaijA
lTpiVafbXH6+yr+708CVQZpKjfY9JhhXN1jgU7hOT3lXJ6QzQEzy+PFVl8AKa8a4
wqKbf6/xDoV/lYCTJlVJNfXu75FBK4OLfUHTqU3RQU2EZzH6VR4U4uAZrXJ+ecQC
jA2/qpuJUparSJWHCDPauqNYWnSAJsc2HQyvjHtsURAA9VAmtqdIBG0IJjiLbOxH
1p6UX3eTvt+k6C78mHnwpitCLYdlWj5weWLrsp7kwRAId0R1egtGyloeuRlt0Pap
J1JC+9jMRsvHHtuUjWfEEWDBKwgPRkUUgvkPtcbCdBBkemiTXcMNUhGANJgdLS8a
dwf7f3m+mlzzDf5wxw76n/KMiWku876095OxqzvV7Oz8esS+sXEpYfCb1FFjsM2T
wEv3BNBVKyjq8Q/+J9O5MHcjUkCf7vtnGQkZ8RmdZKcbdPLztS4DMQbt3WAYBKA3
wqv+mFZLCARJ0EErzGsQQZdlBBsFxCtJFMjxMWTn2RZmAA+taRtGHRdr68QKxAF+
e7UCpwSTABzIJLmiEC+ZLWyoxoFvX5adn3q34aMMdqSKC4s/yzqr/FoAnzhfi8hc
axkJkMLumMFyTYl/3MV9Su9iGFaDY3c1ufALmxMLJuG/hRdL+kYhaadqQmKZIdNR
8gg2m1zCvzI6WNAfCzz7hihwX4aKjpISgN1nS7n3F4Und6eSeW8MwZdUv/fDz3aP
0QRQ7ek3iYeiUZgpYC9SywpxbC65P71QKLy0NGp8Z96iTIH+Fs2JiXmxKvaVryv3
NPPrqFJf1xB19xqWNXbw+ObiNvjNjUNUzYVWp5jCjiBcsHKntG9RgDq9wQ8BALD2
81fOgl93c68lxEH+lYvasOWokfH5kbcUI31QSVcmIBq4beGoVM+Y/Y+m36BMEUOV
zOVqD1nemksBKGo6gnhrZPpxs/rDKEzYUqk8SqXmWZWdjkvGM1gLC0GH80zjZ945
UEK8u3w6o8u2U1g2Ky7no/gqXobIMOZnGvUxjW4CI7M7L5Vq0DhTKsRuM60r90U8
pE0mSViJhzjluIRu4qMHOIZXAC7/lF+PAZM08SzaP+p3l3j3GYMprGKyLXjC0Rl6
YSc7BBe5bZhiHOhQAzwBxP6Chn5+9EP8+DPUARna+ZCJCXwuapHlsZC0RFMQm7R6
mFeY8CE5ZlgE8736gSEQGH0t+DIYl06CVsceXcbJu6X5tv2eMtxp7I3rrhECBUFm
8Pfre40US+WD16E6znm2o14MjX7NQxrgU/bXcDgLU/SBCPoDg6BkdKUjmNJh6G4L
7UDv0bCB7HEH5bJ5kPtvwSev0oUKHpErWBiK3++5LLna0Mj9rgy+rv/3XStWr6jL
/NuuYMs3Fz00vLnfYvCRK9A2dP4VwvBXe+FOIGqxr4k8gS69ExQoPV9AzG/6vkZU
qrm/8+X6IpEe6On0LqfYjH3dBupcJeB55YmNfhGtmibqdXMT25QSLe93OAQbZGEc
icPVWV0CYxe3Ii//PgOlbv2smSdxz9HaJXu6aitbTPGai7ZYiOioG+1NpsD7Yl9P
WoI+qRdJql1BJvcc1RVpNvxrZ8t3JpbJ+mhmYf+w6+hDQMTRR8BDJteXwXJkUODi
ouyVBmuFwAqK+AXD4aS1DqMRS4wo/+lAjFb9WMvvOHyAPEIYTK7KxqnnmpsMXMkF
wWGZToe2jLJIEBbNsaJPP4a1H/kuZZr5b5Y4bxK3p1SUpJXi3Fz6iwalLmS500Lm
mSPENJLspfCs9mH7pBFetdWSsG2bbJdY9CxBsHxMV+eSjgjspcYQzsGSLJeB9WYm
WacoiuDp6UfU/lEzG6zAxchwDXq5iqy2DkXDGMg5w+eV2M3mQi6vUfvsi+W+PgfW
56v6nNpkYpj3G5zewc4yjLUpMSa5gBVoghocY/U90qixIHkF/GEBC2unAaI68wuv
9vNHOmBS8gzsMfBdItrvYiLWTHQ91WvlUCZ3x1FluBdntCTI1Jr5M+gkXOPbmC+t
7toTO7fCVU1dIEst4N3wKexvPZGscrEC66OSAxdS7VRBQRRVEAfF4enPLSngx+4P
ImGSeG7NpbX6kG+9gvxwiFnfVQIqHXQkYmsfI6fnlj4XaK11cOHLRqdE6IdgDIB1
NMQcFHwS7TC9sdk57moHUbZ3heRRG+p1HLjo3Z++mUEhcU7hLJ8AKzvnD7D3szys
svJd+qV1ct1kCNzl7sO0xa6gzlRhhrZI6F/kU1Ej98hjEHfmOsYBsb+iVq4Pyu9F
mw7SKutM0xdgQZyptFJdLo6Bpq8klBAQIRFM2wmmstf8SnSVPCRbK5SUMsBASqAs
k/ukjwyhX+ma3FkmqSbMTmiYJ0ao7/lduBThjzsDPPqdRPDKzk0gYZpzgyEbXRrA
dPjG0iIqh/WIBwpE+g53AgXk9GCILh/a136xH2+0AjBWvWJVL0exGbOKqWAcNXWq
KoAb+alSSi35CU0dx8/+Qa70785WyXWHbrGX6qAO+dMlGDcAWgjf584IOeOLxQXp
iN7qUO6EAZSBpesl5TOFD+DTs46Z70c+yRiaSHzHdEEKbmjJMgF13DciPIkuZEm9
Vz/1BeIzstzNohoseuvCIDSVoptm9WwQlIxgehbPdefKXgkFETHIkCxDJeR10w0J
r68lFl5UsKgmNeS9PozkoX/Zp93JEc5UkCHyhM7bT+81qnM7/ZedHvhGioq8dtDS
IqQ1j0MlxQI+aagek0KbXFAyOMPSGslN6B0KOh17vj63GrSr6kJ20NPsTaF7Or0Z
26sjaVc3VBy6ir1wAA2qvSwHPRD4n11el56pPNHn/PZY8IPBXSfKb0fOOhA5oq5y
0Mf66ETAURMUqErI6nPNSMpSEfqx9AQGuohaesWIqKKq1XsQT/AHo5i6XXcVcqkt
aSJj72J7sgbY/yf1TLvywcrvErZKNHHFkxdsFCOWzjr/09aE2neBYFn8I4olUUsV
9k7c6pea11wo1zM7hT3xOR3NSyp1fHcSBqiVvrSY4UQbR1diguuu/sreKKCMualo
KRmncxvM0b9gYtTYO8TBhx8mDsuc5t/q220RSZIQszB9BBhHv4ZVZCrN27l2QFD6
Mre9i8RD545wc0YdV9GZTc4/XpjTchJdWMaBNITj1VHQyhuRHJqRavDwnlaaDbX/
jtLDU8gOn9OJ3JhxHr/VfBdjmQxxojplqAw94SMGBqZ6XyFdxsmf8XaWLWZ/5Ze5
mJQn2PMDUbjtH0Yq3by/XK46mtnpfmidfyu4FtOwlU7l2KK+90x6m0W7wFrxG996
mcZs0ohAKbOYZ53LVxwA4Tw+h4PomSDYxMkyAlaK43OxXTWjwyJyKoEEIWhAEG49
KtWcdVk1vhkWwz3Sx1P+SN2by8GiZjstE02pLSejbK0MQykTWx+aYvLeXe7Z0qqB
NEh6tBGr2c299yZDhUBWwbIH1zSbNc0u3irOkOWTH+5BDk4O938H2bDuRUIHILRe
YCFL3D7VVlpNolcCKZIThJNhkEzjO3QND1zcbhasUHxyXhFhfPpWqBAQIE4eqMko
f+lzc6hEOplBZf1tQAsjQhl5ZJiAbN/Irds9E2wN8LqzLCetVlpFaG8MFz8N1HmH
alzwq4PjVCapqa75/UPOFG6vwCGTg6lf7vp6yrtmwLnJNkgJ44BzfB+BMaqGRoiJ
vym/Kkm17RWuC++lzCM0a+zTahu8EqKTyDGrf6w2FBS5m5LpzuuQ6ssfaHEkYiMw
y8vdRaPlpcBXQ/tX0NmOpc3ypC3aG6NAVOBkwFLQPszQaH1JDbQ05kQ5tYyuGSCz
7giQD2ZBT9rbuLvpO7JUUNiGGl8TetgUvdfx9iJi/ukl9c/917MHBBH/unAGFxz7
/orbduEndfSzOIAO8xzXEgL9v9EfZgGZ/+2iWhW8wZQY1HhThIIjU6OfXv69R0TF
7N+vzo6xu35X7OcFiWlsJK6TJA86YDWGZ3YxGJnyFjtTE/XwNQP+7kjhpdj/LNTS
2ioMsJjx+8Vmw6DarlOuomvvMIH1sDaFcBJ9NL9NX3zzre0BC13IeXhN4ZM7ya71
sFiOU5VzZca3xqXJUVNIoYGjdW/3J8h8VodyV+jwKDkujAKdgTkVQvDhGC6W9vsV
KpRDRls1z3xYATizHvHOI+j0QFv5CZxbbeLK8Lw5Jm2X+FfavNgEGmnSSTizRhvb
rVsSfEqQIvvgECvZe49XL1ZWnogwbffWgmu/LQqNY/85E5Mj84dmDvnrMHPtulW0
HLI7anaISuXr/T//xf8y1dtxktWSaaJ3KKdiTjMBtudFeT6czbfHudKOWqIJIO6c
OXH6lrX7Y4FyfXD0iDBb/SA/eUTtvNOhgYYnyMfo35YGEW7mt/Bh/lDxM4SjAK7Q
dtbpSZ4v8N2dgwIM6dmVeWN0gJlUScVqxJaTw54ERmUHu2hOw3apou1JTiJS5Kvn
mWXhBJ5nx6aoAr83HhOGP6+BWdZLgLYRFVIuGJ4663q/cSqpSkW4jxbG+/vDqmFf
XJuTjxiSq/KXQneBppx18BPsFMm6xL/BldirlQHWAna+nFnept7bdJ2p7dDkTiYX
CtVjZMX0DHEz0tvkyRZ1UZYP70ef6MikxYE2CV8Xy9w1QLd5SOAidbpNbZ7oP4oc
qac7sHt0arfFXgFkU1L3v11W1J7/p09FTRe4Z+Ycv9l+lDkUY5Sr5BsjwtheiAw3
reG72bKit9IT3IQwNJW+/zg8CEO2DfjdePBjVWq8pOLYwz5KdCHNimYxzU01u98n
Oxm5FYMkqluZfwOEFKvn9A9kakejZG9rOsJ+FOVP338EQvJS+ptEQQTmMx8NzdAy
3n+Fc18NtgT4QuRHSu8ppnlaPKEWP+sU/Ti8CCpPiyitRJinNLmMUH2vf7kbweUF
vsUvdIDDYe8qa2A3vaIqtImz5qLwCutyJJ2a5LP9URh9bW8680K99syI4TBHohyF
nKwgisGjHH9mLJgNu7B9C/HfrMZlbux4fetZLFgMhilS8bvbSSbf1AY2I62AfUOx
TUkNm3JR7BnAZ1Lc+oR/WKsCUnYNae/JrZpZ1qV8Xs0xpdt4Hdjswt/i02eYLMH4
rH97dos97MDbLH/9qat+GVXsgIWn5h5AxbOpsUm5sZz/zNP7SAIF0E+BK8oU4zuX
eE6t9Yr/xcAF3TMrvAwELReb7aNNvJAeRDCGfn/TZkelL77pCSbcN9bN7cMKmW1G
c68c0QpARqr+CTjW+827XsVERCHqD/9NfEKy7ql1zc/mQO7C0fDbNWK9dM8n3VqL
VNK0rlHMCnLk4Z2kR1aDb5yLmH2uQjexkItao1UBhB+JFf2QpYg5OCb5TDWZTC1y
ezk7q6FEA+7/L+srPiD5lblKB25lMqiJaDMEtXOY/mDLWiVFFtTCmryB5bgd4y+r
cc+EixVKssihdGXDjuaMtIwNqH90jFLKBULkhuxdGkXBhXYFVdkKWyJtGavYCE0B
mdn6Pf52mnp0kyu/SfCi1gnijTrspqRrtAs5RAmAEvjOrBrx0XhwiUzqkVMA4aH+
XrjH0WO9/DRCFexQdXNK3XhZNQad1n5tFqmO1axiMneU+B/Ds2DSjQrmZ6LsHAVF
ngRwoT6kJALii6saH3XI2K1sNKyJcYgTtaJjkqbcOyHKDxvjCjuYx8mhK1GZBswy
08MxMAah8IM7ZhPqpbyK7LPCOnsfC6EeVDRE9YC/4DgiQQws70Kk3VDTO5gw/Hre
+Ah9yfcqLY9xAecmTOwfeAnt4R4f6GTEB23Qe5mSmE2CUM4s9jwU0KBbP6pM3sLu
YE152Hupr6VbmBfaFZ/69Fc9Zk5+oM07LLEoYaHLLtYNPGR13VbsIUSw+RY8NsPO
/7iLbNEL4wiGkLiB5zChtGE0zDrIrMOUXkZ9SIAUGTWn/U1xawYU+uglA+KoQTyy
IHJoxY2oqOVMNQvC5TRT91zASVrnsvQqMXwQ/tBRjNevRYI2rtFuNFT8buTF+g5M
ICyoercwC0sLgeAbbdkrVC4HStzk3XhCVtcWBagIfHq1SIP7WIEnvZkrUZpFIXPR
wi2yPdoMEGUk0VyubtKY7TGc/D+9HNbrWSO8VwEFEV+qMdY4n8NV+sPraT6yHRgq
p1J5ofr3BlwMjW6fvyMyZbjq3PvD7gN0wZG9aE1UeWqg3PpuLW+sEnXnk0Xp0e82
e7NT10pOyErR1HjUQP19OnPkyc1u1bUG2ZXXzc7wKDTfGnnqkCZAx6n443aEOqVp
tdK9X0vrqp/GDhrj/6Dfq1v9gPJApn64fe89pIFLXc0oAxEErB+bAPX755geHph9
1q4rmCDO4DZH9AbEsUtRPbppm7pXnPqtJoYsfzEnM+Av0ox1aYPXS3w+TGLGac7D
u+GW2bibHUYnVVmGxfUgLQm37kE0OcWvmwoQD2JZjYjhLeVAemY4tZufRD83avNY
yO+BnYfOXiCcy2tD7OeW6mGjWGtCZ+NoUCfULWeHX8i/CknSSm/bb4KPRh6oMlt8
c01j5h3gAkTDBIlzkzE3kly7S3uTk02O+a8/FaIM9DxuztMlCwIaAHH/kxWrkNH8
JzK5XQ/azMpaID59yOZVt2SmnHZL3K0QZO2KjSt3gzr1NgcOQtkSMeXtahvxdNqM
nOOgn5KndWEfUkL8KmXbCz6bBrLc0I/l+DL3L8qH5j2bAiIM1OKxEa9RXIMoyLjl
lUp20+hRG0bN/tfmZ+GTjnXZMzx5mwL/IjlyAOY3/7D367dEY95jANjE9t5+kNDG
RADtmXiMppeoPy1v68VB0Ei1i+Q/FOfg7s1CQ+4CfhDrUTLm/Wsb0QgzWPkS20pP
KTxe2xilfN1giAIf36dnYkDdX/14GShghz1G3DNOmvlav3i8YR5BV5wgXBOYZHdm
kwm1Y2FY7O+E9QVimO1gdVgRW9jsc/ab9bt74nq55D06KHnqhB3AMIpqFSMIBDW2
QltAomIK6vfFDRAvAZvv1+TxTas3XPPGwI1YhUt+Pv3CEv9Ylnx4jMqi/oCyuDMG
oj/nOSBLvd5JwLxv3l4GNk7u/SZswTRjeb4SaqiQuBeuAWUFOWITskz4RJkUyLZ3
04gOnLXI/rJ6sj/BXet+oXLM8lZzY1FHq33ZLMHA8l+846B3X/gRNmROeMoICgCc
A9FOGIQfBhpjyXMl3pO+W5BmFJZJyemN1D6agyiY5Lkg28bQ8eflKVj75jZK6F/f
i5+a3GOSmbbZfaVF4jlOEfuPDhr+JQNe726aJfa2b4FpYW4LbsfuYy6tOXb9qXOD
txvv5Xv7OU0yosuCrreVg4uLbL5Hn4JcEsjUetKdCYtr4rh9psqo7tx++ni9r2BG
OEt9ucwjwplGb+imbIDNHb2T7F90GGj7m+wrlDVaWRS+qG6rItmfikkrfi/OjSOF
2OQ+WhpE4QP+Deh/HqX2kLk8w9Csk1FzW6R22hCzdoQeTWsC07PcJ5VphwxvM23q
3H+DpkvaUHDAA0wKOdtI/q9ldH6qT++AVDj+YHDBZ3IW+KISgH0DGfWPq/qaRV8i
3cdET19Vwzkyu1iMkr5/L1Y7lfJEsJXTqw1HXsgXrSDkhNbPOq8flZrDgCz/i1Tl
Jycx5uULOr7boaO9pt9eJbdeMOvgfNQZ+mw+mAd68An/KXWAg8km+BVPMNPDlHGK
L7UyN5+iAHy1Cg5CwiBFZL164kJxEzGLrkRM1yHAHJjXIyQDMO4y4LQY1GV8xBeq
owJBwZ09JpW1PUb9S2gwa88bPMuYhG1Gaa0Lkx8HkpRFgljRHaFbdrpAqF/1+57e
Krv2RhhDtXHI/khzFYPljuR2mzzDeyHuxSzdsiqcpT5QAtO8CjC+HShd2tTwdyLd
4QPBh0Qsalo1y9i5X/IXIROJaI8AlfM1c/tZ7Fxeg1V6hOkI0slNBZMFgF/1LOML
OK+YaDgt/Zhn4hruwfcVMSZGCVJ89CxSQsrHFDCZCFiUHXM7W44AcMaMNuDyXK44
5Hld/MOY6acvoqCIQ6+54arKO9XSG6wsk73/1Yv/ejHkFgKOIugsO2xVC5Yq1QAs
Zly4QrYlAfIXYlmfJM5g87RqACnhxdZ2iNXrEEytmTcyDY8B+2G5zypqv5YvMnwo
ADYwlwoTzGjMOQJOVJEvfUFC7lOxA+gtmQ0ZPBWeSL3/GX/6YfFG1InblfiQXb3d
qGF7+E5GY+xZHDEWQ905tLLD4ScGK731DadhxKCJpmnv/XGBvQDE1xmoTM/YT56R
PE16OVZ8dAh2l+J9fRDaRVzc1pdsiJDKgswQ6L8qMH7CF0s6WazY9tgviuiFXGJL
uv5HmLDgeX9bDEzqRYX/w1dXuNZF2TLMIlJ1peJUlfKCcW4UpsOwnrgScOUL3cL9
ov7YVpCavcXCU7mJMNnuqCqebGfFkUWHE7/b/2ueZcDyqpBWSutsHnnzZFpDmQod
XQwcjbAFZ7vOYUV2j6W7qCn+lBR6JlejN93hpXUYIvsa4wS0scMUeqmeOQtW5hmv
/LkIL/A65jay+699adhomXzZrtBaclK/fZDpKWg3OiJt/5xmwHIMtLwVPONiK2TL
0HAPSw9Uk0IdRAl3th76qMXcm+f32qtV4Od44wS4vnWFel5PVG3ICg0se4HFqq4t
Jiiu9moi6f9AI87u2fAte1VVu5ayhwFql5y6jTiswrGxy74L1bCBCsgZyK4PNT/T
QEHX3u08pH8xVlcaNQm7DHAv3FelOVFtsdM976wE/X6iXyjOFDNsCCFfOsGDZuys
+wCwM5GbtFhWYk4pp9wQS/f+cyUvWuwXnBYSh/r0Jb6354ZjFOvZdTDvPksW4g3e
KPqk5GrjOPP9TnGvDn7P7E0nmTyto+OH6vBRAwlu5hrg+bMzbW7wbRtlhhxALDwL
v2rE21cqBdI+yif8/dyOZXgVHyfzR4ts9Uz8Fg2SuFIPYdgG5KllMkFJPFFTu9Kp
9q2w2PJUOCMdkKQiQ7JIiWGXCAzeus/UB8skSp6m4xjdhXq6qFwxor4MQHeJZS+5
daO8B9I+W13oABSGlBukocvkDNpjfZAK/aMIw4qzTgxNvUoiC6u94h0W5Xv+nE5X
vKn+XwnhiSmVzXmOnw2c/3S9YwFpjwYrbQ1A8AEcl7PTZhpfH7GlJSfOipLD12Db
8YiuVhWKfziT0qkhtynt0nYyKN9uTu2IylAwCPMUzoSShbVXJBf0NOA2FD66jG/4
cwBcUhyJ73+8fTIaU78SnXLKouSWnakgdeAWUsVEzuNoSGtKLHumsuwaHZBeIXyW
GoaDVOkDImnwQG31NMDcAmGd2jF3tpL4FaV7H5BMRkX7DpcARy1MlxVGSUh0tRN3
ffyQrhlLrAdonLbLC53vurToOrge8ssO+iPbGLPrLAMEuBjU2/71nX44Hhc47eU7
Mipr9mMCIahHyiSNn1ZEmYh5vTVWhe2HwpWG2CGiwhcAt04hG6U1qxwAAep38PsJ
+KsOwww06+5Jgn9baG9AFugDNlWbwtPbgzyUGwx0kf9l08ShfPOyXy7ftOUSKQ1G
YvJa042sja37PMcw26nm3+1W9BZvVhF8UbHs3RD88MqhuI5OUrQef2s3kgSuKTKZ
8GbdkK0k58cnc//3y7QTdTXIksvculI87OmTkUqelZ+m8/k2aOTq2Bl7x1mwNr05
Cm+rxqGaZHj6HuIqjiTgOo4tgMv1q5XvooSO/deyb0l77exqY9M/Sj+RqTTlblKC
l2ptgqIBO4/Lg0Ia6qtA/d5V0Bdr263Me3xdwzu7fqvbH/oqHwp4jQylAmStWnig
pF6ImwNv2TsENl/nSRxgiucJbgYKmcdPmPDI3EhByLqq92JZMtvxMJoZ/BZy4gDq
e9wLVy3JcVrkhncTdTwwVH7y3cJZB3SGfU2nnpTj9Kb0F8FSPz9yAO0xaf01l9Bv
oBWBB8K+C0NKH3WLj7dwT/wQLepp1OE9bzERkOSbceA5EnAY/XdBTCBuJYLUczW4
nhAV00gNduiQeKRIwqmTEIRdEl8sCthl/EiNIF513ozm4OA3+xFmzHJ//eIEGw+9
uBAoy3jiJDEf8vFXYxsWoKLmtMrojHkW8TJZNyDsSl9I7fs3vvV7jhrYMN25KV64
cGGfh4OXMVkOvvAgfEn/NI1v6R/fn0ABGsyUElmweQ3N9YpVG8vXxfftWWddet0P
3MxWC3t8E4tC9NgxBNpd3W8JYRC7Ubfsdudb6y+q2WKbZ009D0iMMXFblHA5baAW
7/Jym/glPwfq+fuOW6k+MxTuoJ0zrpPYCbv06uYGo7wkJKJkktRXBxK735o1YMrm
9/mxn1ExFpLTTayTPBI75MOlK9yQ18dMF3I0C2z2OqBtYd4QufmXhHB/frBGGsxs
nl7jBP3V1Zaka76zIbAaiW4fmXotEi41KS3tUkumcfxO0+4ayofQdcjuIcX+yqc/
oh65gaWD8up544WstEFDgnXPEh5npk4DidXqqG1+sjfmbfcIyw63NscyCTldTA5q
AJTnPgIYKguGAVi6ySkkUYS9mLlQbWnPN6vinRjqhFvy9aJIoLQwN6+9/nAw65CG
pab/CFJzTT7qrrdsHnC5Qpz30S6H9r33LWe4u0dVVqLrKGymU7pgMVd5oIed8bSk
z3w9JKhZygPM+NsDTbaU7SKRITQ0vXPeA9RGPq5409/M2HL2Qo+CEWuszo1xQ/0o
xqF2cJxOvrwTDNPWaHi6r9Uotu3kpczPpM+3k5cz1WH8rVYTij+SPBnWIrhZT/AU
Ns1mslGKWfr79hWvUoUcmajJdw3T7GfnY8H0rWnHycmB6sACpuwL8H9HZKQzo6oa
gWS2l7dbqhJVF+QPdFd/+WMughBB846lcQmz5M09L4p/vqj3WaUxYagxZqtIEkA5
Ew9yiL66gpGKwlYIwS51pJHR4HCQjkhXagGAQA7OTBBu+KDdnZ+FQaiRu/LbdtUi
TcIuV3F0ib/fzgam/3mvib6IrithJ91M52yUX7w0XxYB4G5cZrEOQgCIauDvMoqL
ZprHylQL20bnLahrmxv5OmxqNviTj/g9bJKBzJPD9z8qiHfiWBkNLmxXNhYgfsPl
JGXNyC+DGdVAbZ2tNB1BhWt2Mvh6WcsWZXzz1cEZVLTdLW4hR2Ezm3aEenYZQDFY
CrYKfUJJPBB1/DWwwyiY6mSGIAVJ9fhZfz+zBR4J6Vei12xVB1YE2x9GSLcP44Jr
qBoSdPft0gZSagLHLgGKMkUjhicdGYGSSHViKJrwzDT6jF1u2kREJs+0APrNPEEi
s0hH73FT21xh5fYlsDVUH3mDfRPSgnTyzHykdxVN42UHCAOmovHBwlEKxVQg0cIH
WcZjSegEDQ9//IKYWyScRnQhNPeucy9s778OLZPSLt6xovJ5FGT1hFTJGENi+1UF
XxUb0872wa0FlERiGm6hi2NYfbM26/hmSa5Qypx9UV4811afQFk6pKJmH1T/QpXB
IOa0bFGVsmHcus9hv1zqaKAaqCvJXCP6qP7i0ubKg6O7i6N/vZOlA7I3eNz+IcRO
qufpWQoI6rwq87+zM0Y8rdybLBWIg+0qSDgU/0YxHTvSOVxUz1EymnLLKgOnjasq
d6/sy5KoYVk5aU1F+KQQ8khfZwyl0rWPomobX+5z2nI3F24P/zQmiEk/HhZodtCY
u2SkQX2poyUiueEnv59ro0k4vXqnpgI3Pe54L6og6Oar3hDY5czn9CPE6hVpZRt6
naBbMOWFxj98/3x4QsWvOJepmSNlTPet9x9bnyC3/rgmqsmzOeVe+Dgx0NjkJtRY
JawSl2jCKEa7M2NU28DyKAiCis75yuT/yoT6CAkoezgVYIyqplpcU0C5aHe6nfET
yr2+xSKdKe9Eb/IC0FAq/0+VlKnJEdc/7Ok0WVOlQdmF5KJPR6DqYcUfE6H+z7LU
Ur++JdFSBCU+SsyfrRSU3DiP16qeE+gi1BPiiAuomvehV71M/Gu2EQJVaNgy/S6H
yi0kANgnm2WQNhDQviHqlLBNy5HnB389hBIF9QQVQ31otYprgqwHbSubQgr8/FDj
TETfIJFZbcPByrVAfnt9bPPNp0eIyAiOcejp7r/CkZ2BVkdVOnlGsvXr+UBGKsFI
p5+4xrhI+Kp95IoupMu8XbLXYBjsrDM9fXXTbLFO+EGTMNNt9zpA43sZfBOmPWEH
Z7negDv0tMmh6yeyXJHKkio6rfuVmxy3Alv/1MMB4I9LaaWzFUEyPHqRY9KTEP2j
yELdL3vi3JDSyRPG1/xbP1UVYg70ttvVm2xw+w1mhbfqAU6t1aIL4nJIdQKNzT63
LUD1LYUxgwCe9eyMuz2sCgMuQ2B7dcXceEliyKVpcVRr5aI15aX2pNhhwXavUnxP
ZhT+HaKAkdtQqz1kORLzz8mnVDuSGDwwSoNMVXwoHmBoKnBLIiELNG7jrR/JJ3gs
yfTkRx1iNuzJ110+UfKCO/eEEuihNb6zTPBYNUHKwxYA6iJwPKRKUJv0FgGnUG4o
+wMvDeWkGgHEMNh75uWaE+2QXZ2ZktGDhtamVC9ey8nocmJ2Arbx7wqgqTpxuuYK
LSGcjf8m0fBi1I4Mw1pFUGQqwXlr+oSSx0BDQz9SzhB0trzbQtFg/PZbKHTdtJMc
xdG8y6Szi+CLeEuOZ3XMiyuheu/bpGtf9xO4N909MGRHiiqZAHeXfCKLqbQn8I6i
8GvMQn2UvasUvkdP13RQYrwp5Z2YPZ3gk6DnOtkWGgpcNbw5lwu+oU6vrWW1X280
2f78J2NjpvGwCMsyQkCvoEhFn9lutUG/NCAN4SBTHcEFVpcfiWP2nXe/5KUQxM/e
nIBuZtqb8i/7x0zC8E5cLzRpS9WzXef1iMZPng4l2hPo0x58VHI1f50eO2PcAZhc
5kJAQT/Rkoxt2gRUcwmACcKqqx8fy8bv+J2SBxCMj2MUClVNNe1ilJPAvtEsYQpL
91rnI/4IHnWcDB6N6SDf6royahq35o1xQezfMukNrOtt8Cqqvli48dRCTZ2orW3p
lriVOixY1xps3PhejTw80y2Xffdhuc256Dn31imTHwEdCyufcLDJZtmd6Y4j6IvS
7/9m95HGzIn4mqxdhxRjXoOkvp0D7y3tCV7qREUqMIzyJmMo0+9Y1gZ7oboKDoHI
Lcf5vJyei+j0ZsJJUtiRE71wOHsqZZAIrpWV7U1Sgy3nxb0mvkONYs4pHC+OJ4AN
ldnUXoesAMm96XRlf5czmPjLTLZ4QMD7prAaTRWTAW6JrConiveqN8jx2ZnyNKT7
vNyyo0AMnnqkgo17uexn+CBJZnzwpN7hu1kP6ZS2WiFK4w00FSxLCbY0rkmwnsHj
/ewJq/R8lJ6uV6XGhYiczJagQZ+CvYxdlS4VJZvYZMUepZKb5mszaQqqkGA5Z1GS
zqttHC/cwXjWpv0RsSmiePwIyoAYsEMKMRGj7Q6In/sPr5L275LNB20gwBVazY0V
RNRL22QeuN5aSAMbXMUcYXtv8uaaX9Qvb1o0vt75DyfSFLNokeRlsZQsZ8Zp6QxQ
4wN2se/v1n9QKT04VvDTyhoco90BrEf77CilDgzQaXco+1VhcRbFysDzIZkVDAbD
5NZj9pDOpzvIR4CFyZPywaQ6m1uNMGtnTzyQVTsp0+SK4YKhT/5yiIOX+EfmlFft
F7VHlKauyL3eV1mQdCBIeOoht8W23QyNhyIp57GbY+qCFE3dOGLifbClgN5+OL+M
PjN2DrWkkGn8NoitVg2skwtqwRQGAVbaXmmJHQHIlDCFljJtjTMxgNkMbd1YYW7d
V+VXTNxE3a5UKy+++Uo/z8yytLBw3itOV6Z80gc8L8Q6R2kwM1OZEEO2IfH0c4e0
wuk3dxObe9ljME+pSxxyQC/GDIqXLFUKkbBfW966S7+3U58NK9Jur43tp34g/VFW
0pAHnuFIxH7bRu2CM2sHlbdbI3xdvckIDHg5SegbCd6xnDBH/J6ekLlrjzdtzaZ0
ckLTq66yyVidQBOgpa735uQ+QasjbLmm7a0Hw9/2hL/PoadyUHC0EMWZ/rIPuHwh
NHdB+HY1XcsSL4BO62OEXGQZb6/Gq5v00NS1DGtaFS/wMijMFCKL2ckJuTC2y5Nj
+n7YFfhNzTlDlIARtjoc41GT3LYudw2XiF0Ff9Snc3azk/wUnsvoSeoOacFRJvcL
H4PjWwjIy4KKvcwzjgSxEXYFrj9nNHHw68+49iG1awx5MxEwLOfWVZvlNe2VKRi9
tRANzPCLsh7K1CZJE9yFicv6IaKaStWECJEXE4ollIJUQPV9bN3epBkgmC3XPVov
O5E0DHxiMIDW3YnDBCPlh43Q79UYpddZEK7CusRyZ3Re6R8ztGn9xEqm5vaPnETB
0d9pRInynu494cnVSPNUD89VIsCCaYa5QlS8tvo4Uj3paq0vzdwYnap3iUO2Ba4c
l+FXmcYpe2oRXZ2gAbbPW9qa2mHYEsb4hchh0MXvg+AGHI1y+uR2DhHFyMF1wtnm
OnXaCLE2W8r9bUd308zqn7DYs8s7f6GQLT7NYwQS6dsiCsRWXTNQG27d2/kRWpA9
Kz1GZBwk7l0GNsd1DJ0XmO0vOXvwyM04bGPx1PSadSWKrC+Od0+xVKu2vtO/UDKc
1gJcy2DYe5gADCb9U3bqJuHcGluCbbc0M3iTPiC9PrdnIlUuFiVvtHwBqfOXIfNz
2XXr5fP7Q5EegNBmwQ9+5TltQ+59U4vgrCReTKSoFx371oRk3n/UGk/oogSPb+kU
mkKUiCHCTCFzxtDKWGA/91sFnTTVT871Bp3l1WNY4oFiJIMcMVzIWaB4Zm9DhmkC
rVOjrx1wmiaRtrjy0xOwFOf0+OXVWjJ5e+qgnc/KK1VLUcHasMWOHjuzpmdTxWvL
7HLnYKwo+yiCB/xgNXNQgoH67aC5aBTvqrjPoSyiCfdJuQH+CBntK4rFATxtxNzp
dZo9Mek72bgNQrJsJbHbA6qqD74G5UbUCy8edcbRsBVEGtrf7haRhZhwF3C2VPon
FRFjhRs+Svc8N5IEeftmhDwk4UeXEkN3anP3IjPYh9P+B3WqlVTa30hN7jiU+LLa
5zQqWf4Bfh1gv74f80Kl3hNmKWFIrjphEZ2alZO2RzGzPSKnAIvEgf6hZ88ad3aV
84mXHXrSZNf3xqDDCfW32ET4+TKkSMgpsz7RTE2ccSwQBSInorDuSCzAEk/TmFAZ
xp/JAMkhDUvvOQsmnQMc5FLtg7oLzEiv3yMsu4nAl7419XAVR7NUDRQlACER6/Uv
XS6YyPT/FK5TiHwcW3Boe+bIjpVwTp81koa7ClMbpYF5UpJSKnkfDK/u3OyotyqG
lVlyh54crsnHXBEOjMCLp0uCprKiLhISFXQsn7YydAqE6wmpzMpxB2n6h9fnn4BX
hCTY1dzMuJtD9jJdbKe9P0cCh2in4cuFd/m7zEyL//jrbxlBNetrj/j0Rb1aZAfe
HGJIZbXgBxCqmnjjcQMSzhz38N+hF+37GcgpQ1SfUhf03QQbSl15auvkMpjRepey
G9GmcJloK5t17S5PFnp+Btkglzt6hxbRhzj/vFdWabzI9MkehO4VHth6TngJusm5
kavR8zGGvmXHj6XFTghOxsrhY3/Ol3qg7TAzCsMww8M5QG8UhPg1/K8+rhU7HGIL
wK2ssoppJgQAxSx8ly3Ydp+VwGu8lIw5c9YEFN5dpHJGqfRKzmuzWgNqQ+kRsnOe
MrWOmwGec94Iw+Z8lrcwE/EOb50U1LlEljO3ShnRZUUeqdfQa+iRET5lcp9Xfl+4
Gqu8atG66/6oaxCw2yblzdSVOqA3B+jt5h/tCKHDm2M2BmsF0AjdFBit0/uhxdhE
NCWnKVBHzavx/PJEM8J9+9O/OdJsaDFlME//gEr/cbb7bR59g6PllWACLrRhpiGy
qQscxKSZ35aoXJZd+ZMec+QWnU39vmcNahqny21fxozj1in0FvP3rHnNjHPpNCrP
9Dsqgu697JtZyoP3kLG2xW9V32YouQQKSnRwDJxCk0eY7+oSjtvbFxriOsflpkTb
92nNl21sLNPX3eV58Wmvr0GS34FxWLHWNkiGbbMpKIHMOrDrYxxX/9HfXmyMxz8j
tKQbVMz0wTE+0gS4ClTWg8wno2OdAcHdpJ6eKoYMkBBY5lNw2p0Ui++Ybj9l42zZ
TWwRhZW0wyHhClz/iGvNoB3NImK4nnTAFKZm5mTZ/aKJjpYBBxaCTMYsww0oSQyn
/0tHgQlsOsY6xwU7ylygIJqeDXZ+lAz7widRNme/PgTzZ/Jcpkad6rVSS3mHnuvk
/gY0nJuFlZ5lQ9n3tDGsHcu84mHIKxDKISJS4jGw7yB5Cw0RfknL5CcXxDkNUMXD
nbGJgb9gSmqt8YvEIUpOkGf1itHtBLs85NlUHNVBk3RyHcGpaL57BREE74jycS5x
5nGvrVxpp3FX5+Ipr8ImbjGSPizVsGfZQpwiW+nbnI+UAEwcQDkZIVZTeBFNoYVs
ozuoUbvOXLrMgHdqivyqNQsOgGfalwYUi5IjrAx4PNHKftnBXTADNdwtB3Tq/bp6
awHThv+920HZSEUxUJdYj6lVPyM3Gf/BMauYeog8EzZBqZTnoY1gI9Znqd02zjOn
yFPM6AQUJ12I3hNQ+IaT8rnwxjoAtEDd1KLQ2VUVnKi1LyND3m3LC0m1EB+sEQ1E
QahDrMz1LaaMiIxxBo94PTLFJzjzdXVRnsyGVWl8Vh4GMsLHj+A7bPjqICXDCNG3
5egSALOM37wUlrmagjC06MQMLLn+uHk1LV9l0EDwXT3wrjh4X8hzyiy0jkucv8Sd
qu1+o566cSkz/BIYin2XI0DlWOwyNl/p0ctXj6sTB8EhDixIIkYxCh2d7rcQEGW+
FXOZBZH7vVLYerUuVSbvfxiOYpEyxLkx5ASzAt+M3Sav1i39msThsJ2tSJDYcFTG
8V/Zq2+6q2wlTgi+99F68eOpwZvL0VH/IwKj3ax0Igh4yGG8kpx0ADIw57yFBK48
NfLSI2gQGPE0t9CRKbCwvchCUz74cbbpN3/300Y0dNaYrtUB8kwqcx1kH1wTR951
oC6GKzpQBhRiXQP/E+JgMZPZmxwhdHrl5zJReBAmH3Hb+ohLu4fFF8g24F5qM/Yc
17zl1ca01WVTqmRVPHKeqkJ1wUbI71HUzbUgtgBWdSLNyQiZZJ3S+RfFI2qyPt5/
CF9Zcg2OvYhYgT5iltis2c/pXYHKzfcPcFmWikPYpWzmJYsWO3uubL3FzPrFyaSk
OA3nhAMxawdhLf11uz671ovYEaB4+dtovP6tpqHVgZEbukXcmwNvgglMb78xP1lu
qy/cUd+de9jWzUKwSNu499pVM9cJPtH1EehsR1FIIw6ZjZfGEbH5sZrmBP0MOTlT
y4Avhh4WmAPi/poXXCnqf9E7OzeYsib/or4MfubsuGpbcYm437GKodhnuUmowBPx
FjUrX4VEuvbVlvWjkuw6+ypJqE0kDy71cGKWUKfI3w/e92iuS6mInOsCbTrIAmws
0QGqVwfcpvCbg3ssd8j+nwPCmD6MVqjHCrxOBFzBHNfbLgTF02Z0WGYQZMxPNfAM
1Y9txb7ppK18rj3WPSZZkZvSN1D4hDwm/oSol2OOBTD7V4PjjygVuElhh2Ivyf0N
cRHEadVOrSVGMKPOtCcgF4/j5iJ7AfhacILcENfVU909WPnPZjSt5cQAEvof9KsO
rnMZC3woOZAz9uI6++PCJ9XHWp1V1hCYFRCMZg5tLIIiKST4mRDErPZ47B+EyAmt
MX94oWIi8WNdDfweN8yIrtWJBlgsI1OClEHxWiUX6BubQGgoYo+mJMpulVejxmnD
eg0DTTRB4rgiNs7uBN9IpBpsVBZHb1EhPzCLU0Y8bJy+wA0i8rz5/TQxLN6qm57/
nsU9pzWic9wvuC4rU2EdTCqHc0dkheiA4hXKUfAkg/X//P6FrZcQLCJOFAFNSf5V
sDf5AVZ1i6H4pn88RvJ1eK8SBV0nDgL3kTNTHgULvLk2S+wTY+7DGkR6IElV1ImM
zLbkpkIkFXTTtegjxgu07NfomVtykm6jYcsWNcdtWM1XvSOFmmevP+mT4NHrBZlx
2sVG37FtWQ1XMMIK523FNeiD/HRMREQ57GRRpyiEmNxWR6gekQISPkR2Oklt3pot
x9qRGvi4Gx5p5r4GboBW5ajChC9IghslndijL6I25C6wgmjv/Ywj5oNEuCC7BdrM
UZCp8EdPs5PTk/ycEEhOxldblkeeQyR8NOhT/VCfRcFd1suufSIKTT6++oUgUrZ0
FcR3Gwnh+pwMlh2CSbxuyyOMJ8g0I8yhmJN5TRm4scnSfEwgZNRdZKXCOmqvyFMm
6RdO6zhNzXlLud35akaPlmj1W0HN4YLaFl805r9x36VsI2GIMK4dYxEINYVcCWUq
USIZOWNE9Hp4SUrfwBlmGY/eZwqVjBT+Hoowlq9QC7pLwLYwyRogMCNGZ9KARBz1
ssVvY1UnWmCkFuPUy8CsUghkSynEXthnNH2K/s5S+sUDyWSYItDDQrUkQ1HftqGX
Nnsf1qG0CfhvWMoO8VD1F0taP1HhcVLffm2FwxSU784WvILMS7PD/W9Nk4Qh1JiA
s/jnl66QdWt2NzWGwC7cS2fWx7LrE/9RGnzt9ObCrTlDeIQV0zk+By1x8V7bXF/3
4wsD84o3k/b70BnexMo8usNCDuHvOhTDjQN3Gz8DK6mFzVIrlJHHEG+wB/k14vg6
6UR1wPsF5kyx0SvkEl0xdBRUwBwJmew4IB1bSqv5d/YcV/6eeGRGlPC1sAgWaQAF
WSks+7visJDAhy/laIZsmRIsOU50tbTpjPQ7Our+D7SEoh/DOzY4CvBRfVY5dMtG
oXgO4r6K6mSLgywKpJjS0aB4gmQ1GM0E0qQnjkVSY7Fwxd4w3NA22+39Leh9H6c/
zSmA6TvTy3V3IoDyeXZVSknKAj9P+pPR4P8wfUr5t/7WnFa62l4OwFBVjViu+fMF
gsqmbQvbF0vEmY5ehTm2Nhtej0FDYPCQVrbXbEIvlkUXFBVKGmxl9IknTYBP5D0u
UZkH51ueLy4B8WnTO4HHjQ+p2JXuTK1KJHUzRm6QEEMUauLHTbMylMpFqlOn3T3n
dIL9AUo4dHTGhZIc5WSkLFQGCN0D6Q3mwpnDCqBg6J6OD18IbmQ3RBA0RjMgNjrW
WsFRgvyrulMWUiDKzrWUuJq9T193nWjfnb9pvf9INd7i6R52e+89pNtqxqDEzVj6
4yUhBr2/3tRmP0TW5RP94Zb2DxC1wUdUlF/v0li1vIWxVCFkGUb8kXx76/diDJnz
hOJMyAHDrjDBxtb9nAMngzRMzERIMqVqP36TyUE+CWXDvIwE5vVmlWKASYjYpLbu
saza/HdhOwTXEiKpDpawnIuS8JGG+7ShYEyQ4QejdhShtJ53TNlpbby8mwrYn9/q
CQGnjDcQoHCKluUa4wpECeIWprL1BgAVVDjNWqwvr47s4wgO05DvkaFwgMALubAy
m9ffvdNCqHzViG8BMHrwjfTKlo3h8GisBvjyu8y3mtMY420XZxt47STMbH+PJ0lY
PynVY68zC9b99Ql+gPFmUjwvhiWJxu1AgYqXxj8EGOMg3kKlwburH20DhF7pfngT
5FQxz/YuUyPQSg/eh/JwIYXX4CKRKuF3E8kNqrf7eUMEZNJ12CGzw870Cl2WDoIl
xcYOPWfxmtbjC43eKD6n2gHQjuc8QtW4zN87EnmcuxVOUVGZyWJJe5k95nxmxnEr
maclgwubwMMV8+HCblhSfhrmmLLm+b5Rt4hjZU+a0i9+eulQnTKHP+AAMXOHRUMB
TsGR0xIHatgAuWsoAqA2/CxPlUS7lniGpWdX0VvT0xWKAvrQIj3URVi3ytPUIJsw
FTRsWdwnxppZjmJkhT4ntOCN1Q0l2feqyXVm2TotTTg3mluwjA9a7J1wEm29ewzM
caz++hxWDJQl0mfUUsRQtggwu8Pf/f0SN3YuGChfFBsyV0lcvP+/3lrGda0BOz6u
Grv3qZEYJExkHt4PZcBI43FkE7Y0XwqwvNBkdZtAk4ZrRVWgry0elM26WT/uO0kB
yGbSLOyF859xOkWdNoOpLap3rdDk5Q2U2NB6+FjqFaszipADU2XK9CzVC7yzwavI
+UxVNEwpXsU9WX+ItAca2LcnMs37sVnmy12AaKbPd/LxnmXLmjAcT2dUXDtzr27u
iGepxWcgExcXf56mULQpxp0SRFEypHvjp6EFBg4klpRAJZxpbTfv7NgdN2Zcl/7P
sXAZLne+JfaGH6wxsMbIQQuRld4dvJVEvAt3j7U6yM2EA9kb87jjLJGoVLJiLI8+
3IXTD2lK2Kqir9v83UBUMJtb8W4GhSfAW9OJjbbP+V8US9wUyYw0eGaP0DJYu4KO
LqBfaYVidcGGYqixcXvM9/uoXhwGCqOjrTKr/WeFHK+QtZr4nFH189GYxdSd2Oo9
X3KQntj8PqB4j3sDsLdGqIzMLJz9HjjpoMoCibFFJEtkNat4kr18yUWt1ERaEgOJ
Q44n+0YXZeM2nhhBCgUIyMRMOX+xqvoOWjCdnsKypMEWb18SK7Z/0ULId/fZg+F/
9IMQiPhvYm8CJxhxQAiOD8hdoAC6pQSxU9ZrJgzb/iV2YcOMDBEST3Db/FhN9YbC
7Mz0qA/SYzNAdK25shvZgd1+W+7O/3MRuqZcb4UOsmfCkAXK7XIwqFH8AXHz7ch6
9LBLT6PYJzBS/ZGh17mrKfdvX4DDkDC8BMRCxrkOSRTtUw5ECfUyR+7FxHVkKldM
72atlpybp6UV1l16LJ6HvAggPaJkZ1STRR+6tyhH6YGpYQTlZCWxe47hS/EuixWH
GK1GeU4qNAvQVidvA6iq7QjfXi4Kr7ssxWByaEc+S445gZg6T0yGs8vwBxiJebpa
9/eAIv0wfwCasEi2ubjOJatH30itBm4V4I9e+aqSUQIZTkA9dvaSLa3JIVG707LO
lVv+CKiQlOUsTsDIoeH/kapjHgBEKM+GxvHUUEMh07m0rszE8qmDsgAJQqr0CVbr
cfQKnBRHd5HIo2jp5udnG+n4vOhOnlFMRpwKljERa0FxxrxfmaOMM6pwTjbOCZ98
VrluZ/1pzAKbUhnN2RSpQhLZkWT8sYmd98yAErQzsPzljH2zoqvJdR9NaqhcK+D0
QuS2wCdFzfbg73v7rosQZ3kKnUXdnoMo2CGnI2uYhxdjAd+6Zb9InLHHnv98WK8F
go5nS41JUtfAckb89pkRTLywH84UJEFNdZQVD2ztGYpSgfzDgaCQo1OvhTzb11+J
qxDYt/klAGNmyaY8LdrXY8RO3XTnRBOQlpqIft67rVHdZi6Lb+liUFa5Q8ZzJfyx
Jhe3CH1t/cM7rAgD8bOeqz9+zxUpXQfkmkIZNb1SDvKUpNZsl6h8PG9zPv3bc3qK
q48Sw5SCcc6+Df1Vimpr0llDzQD4MX229l7/0OT6pPaw4+0j+UVfqjxLwGNkwzSm
zCs/Gx9NQZdQ0Rl/4eBMSPF2NE8KkVSxx1TctpQ3MXTruCdMNSReLlgMqcIDdRK/
podCgVKLGetbxDKSOTKth2ljn0AEUeXyNWGim4w3FDi3fa6PPFJg1c+S4USkMwij
zEsD9rFn6supEiMiuCItrLv9uKiCROqRg4SiYZIz0FcgOKQ/C0lNK5D8yFioSwy9
emNACtuZQIGLZPQoPe3bRO+a7SyZnCyxLnz5/uneT4yUp35G4u7exSeplAth1Xly
8ysRqi6JUrS994YAocZ7pZeVQWsyDiWz1ucqG6HMgFjdaHrkU9xcAPbqSpiMmE5A
ttuuWWfto+fV6ZYwy27z5ZWR5fqFHdAXRq0Vxvyb05pyw2BokxGq0wGXIHgeY2SN
DDgJdz8843tTe+H8Fod38pkakzTH1cIdEXg+dypn5LXYea6mvNTW+itYGCbBFtgK
3fjMffUovaoZ/AMX3L+ZILRQM1Xg5v9iq26hMwDi9jePPvCgV7gYmjtedMDIoCkX
YP3M0hlgJWFJ7xY+AcaxP+glhSEPtMMyu5JVBNLpielwpDV3Uz10xcUvOg339TUo
Vky5YPc0QRJQBm975zEeHw4cWyfDL0gjj3+EUzF/cRd4pGx9H7G6DrIspZ0PLIao
ZSBSL9Amu16xM/KLSSevJ4Hu23c77qu1TBSzF7Ca+tF/iPR1s+un6Au9SZ4Af4wS
QhbcEd3b8OqlF4jr7PO0b0/EVnT+NGcb7zh65iou6hgAUqHA6glQuCex5i8w0uD2
ItidpBYKsiPdgsfdD2q/e/J3fqpIRAvJtjHX0qQrjFt8u0B67RjillSgWePpYxiv
NsAF5ayTkNSRvqs2bMTeJk2M7Gxw62imKIWOUFf/hg7vvgATzUE7FObYq7Accudy
P5bMW5ETfErvMchezTiZKEhRq7Vu9U4UMpBZ/ZGjaYobGJcTKZK+LLBdxk8x5bQE
8vu0tExQevwBmqnz725KduEF1a7NR05ennFx8hPIGyIbZDCDg2gKi3wSC6YSmKZD
4Wk70hwLDyvFYBkZjwC8JrCNeffUNZK3AqeISwYiW6mhNqULf0uYBCVzFSu+BT2B
8A62zSD40EGg6ITbxAZTPfGjCptJHcZkZMA+qFWC7qStTFQP2tKLnVhL8O57+SQH
nelI0/JeLanhWWT/TmoleuoVKAGWDI4yipWONjqLSM2irDCaJxlozbUo8n+XGF1Z
f39iHNNI2mkyhvN3/jrJObfNu9kpfe6y50ihaM6rD29OdnX9FAB8yuIJLThSCGCi
upHlhiAC7PHIx3CXn5JDVAujiDhYF/VIf1wnj8HJZAG7QpxrE51tUt4z6VTE/4DC
iqK3xZN58pGnqD3aD5ATWkJxRl/FGOmESWgp5ddfVuUKHPieHu16iKRIOYpCVSkk
NxK5fOYAhBLRrXt/M3tYJ4vfwX1O28bl/GWTAraYGvZynYarh+60MsNUle6Sh9O4
AuNAe4xPw2/YdH0Vhn/rfn1tqgh8SQTqSTvLcvoTBWq7YriP3JfFDSvfA8Za/tQp
GDjEvK1/5e+hQ3dznp2HThBOdjeTpNtjwVNViWyVDNz/UBjrdNoaOAsOsnu1XF0z
RFk0AbFTC77fP8UmlVkd507VuahbzsLy1zRpDZw9zrIkyajOOl50JC3DMTlNd0Ep
hUvRBe1A9WAxMx5RsSDgb+Kd0kFC5wBVEh+VegxVs6j4CcG+vT9p7Eu2jekiO1KK
mKJNE7JhNYuIwEmrAy2SlJ/jvk6DX8Yz0qbXYZXXvVcpPGlGOnFF8EqJaeHaaW+q
y8rykni+p94nNRcrjZhecQ7E1l1trI53mXywDTkATK+rnOeF0RWDJdpovtZB0VKc
Ugwygi4j4xKv8hb0brPJHF7yTey11i6MVun0vf1C60q4WWWMQdRO6GeXynJ41RtC
YsrjuXsW8pvfyls0dOhhY9piZS65nDfegorJXnaPEGa2nwCMLzTpv96EPV7ZtFxK
ETNcrrJCSNW4vp2b6DBSogWmOQr7IyOLs3B+EOWH2zdL8CSHWVpLl7pwnLSOpQor
o4nDzk1soE3lnLhBpletR39/DLgw2BrCyYgPM5Gc/u4DU2mdDXXf5eah6ntbXQUP
YxnLPrgo2TBvOZiu/3yYqoxq5q/+FEVj77wFLPE1sdBIh63uhR5BzSBE/TYXv/EL
L9blN3MmGDwddAiW0EUwUyySWQRoMN+FrFOR2eTfE5dtCweV4qUrkwL0uivIOZMm
WgXAq/bj3yVhwLYujJARFPoSga7Q/+Q102nH3MsKZTGGpht4IS1FuUJhkHmu5G+N
8XMDePHXMVs5deSaO5tGfx66KnJRBR+lXLse+l9mR4v2TlQQdYWdbVmIVyy2w1PY
5a9JKUuPGu26Lrg2WIQFpXsblMnhUSoHOe3lypDdzVwSIQMWV95a4ZMxvH8Oo0DA
nFIygbI4l8j+yPYqksdFMNK04XwWHZAbLAIAjCnLswXecqk2aC9DpbS4XUlonz6s
vCBIw/5YCL4fRa/MwWfU5vMLRQN1bAfxEkI8ISswU/FPjq5Q8V0XQ8TskSsuDPow
T8sD+azRSx2twR7/tfqo4Djx/ph956/NPB/SR8dTXYo1rZrsAThi1bjidUcWBmRK
ay2hK+P2iquYWVv/dfqKJqLGO0DRYzpJXSg5DN+/EY6nt38l6/tHrI6udgzH6CrO
f1ZvzfL4FR85B+V0OChd/+6AoajvQnJmAg6aMUsmPd+Hp3ojJt3IqYGOGWaQTU8D
PE0SKgOLORe0iP2kXiyytOuz/go612k/bgJCYboqFx/LSwwFkNYoVNhbA2yPORVp
o+F8rZ43Am4LHpjTkXU3YDpRl8PeQmi7UbqE06b7oZFV4ze/8HKeeBYWx/ARgW3v
VBmYwmcqJm7OcR67DhCKc8Axr28YIVAxjbLfCv93HVQttKnKuXiRvoXW7UZyhDJW
+BRn5oJMjKxLdphRWWXvd9Esrzim1a/XFNocSVKKEWF3JVf0anPHGNzjnFU/OnfY
erGgkOCdoQVRgMFuaqiTsDEjbHEcMjOwcyhSz5S/QYULymZY3pH5UrpVFj6V4Vqx
gHJU4ZNXCIVdHzd2QtKB4fdNvPlXKWWBybATS8fMePJLspbZuakIAEJqdUwmi3TA
A291xi69GS1rSUy4gR+LJ4Fij5svGmwkqoTxC/K7r1ca3a3Sdf6X3DnqvcPBxsDE
vUWG4d5hCfRjGSV20H+uRWZCUdCMPpKG1ni8pl0BZIeWyVbvyrVUQmDLGmmlU9Me
lg978X0v8u3UDQc0OxI1uOeWPsl8N+W1Hfl2V/2vYWXugdVw6mmKew6BThoyk4jI
ncFPaMz4JpYNX9hR1lTn+okl8T1cSNuUuuPNvO21chAZ5EANjiDVodyqREOiZ2pj
+8MVMfnAqX/2/W1pSMNVAPHzqn4CuFvzmox4sZcKyFh8CDIwNe9/Ohled7nGx5jA
SzwoAUmS3ky5pWj0S2s6UE5ZPBj4/Xmfmjgy3Fjw3SEwFkW6SLuiTnYZ7yQLPSYU
p3mU7JlW9IkLU3lnToZ7ey/uq4PSlhV+w9XkvCQgU2SuK5EETJvnnF49oa94r5eD
qg2Sh6h0K7HcB0fZa+TVNedGpHUn6wom7ULEIxWAlmcqz60C0rnjipUE3oOLJhz0
TqjgqynHHBlVVGolavdwglQSjiw42unF77OtZCcSJrvlceYZaNz1cabtmTbV/xRz
Cz+7r9R6UNGTZWYxex+tIh9PSjUmbkyLsT2vAvE5n5Jk9CiP73w7pvz3mf+El7LD
DkbU3Qe9dcpkLkB6BdseO7Fv0+4pF/zjHZh8wxqOV3ApGd+xc2BPjfy8V1z2HHnR
D5Jrg09GVYW1jV8Tl1GuqJQIXgiMl+7Gs+rr1W49zjl31yCr2fygEIBG4S/r0JV8
RP+Qq8Xb6CEq+oeKE+mcK3diEviQMu/Jh9B0YvDxYNzIcfcb/10EumvCVu3kXplw
gdAYYY1kvy0V+oU1eMjcA+xJHWA/cFk+57TeHvWbIxPz45X/DmfYQT7KJR/0qNY9
j1UC/hFX1Oi9vtIB2Nd3Mrr4MaP7bUEbLBTUuHxi3h+zdQ3qJHMfAPIZHYXGTHiz
hlioHtTu9sID02HkrMAeDbe/WSkLWuXyDtWevXQOH8RgPOwoSOk0MfbFt65RKo+K
54teUGwaagV5UacI8mi3Vhbbx0awF94LnF0WtTk2kMbNryRl5igHqdiQtFgQVvg9
SaQUdVyyULcwuFHeICaNrlvaTIG1ib75RUPIB8BnJqPQL0xpxuQLVMx9fG0zeVLM
9SttJpAFUDXl6TD2vnzkyErLhigAitJBGB0nFlxPYgQJAVIytWpmA0Bp6srfMXXN
jaQ0zYnQFBfd2Jqk+g7hxENiWc76soc4iHHYbSUD93julI5dZiV3Zf8Pr9gN60U0
uysBDld9iRu3RHoDldKO+6ow87AlS+RRUmtwnY1Tfaq8a13965Wb4kZ4t8z0jGi5
k2szdOB/hthts0uo7wIeKjUHtx/8Cp2Z00DX850EJVitB5PEpW4NswkmEBfZ9GUT
++z+/F9C9zd0oYeuBOcE3WHyYnK8ZUB/NpQPOGVM0tosZF5cEWpxzWhXh8tYG9Q6
VYHKlMdksDgE5afmrxSO4RPcw0MvXIDI9WS0dc+cgiPJu0plDGmhAmil5BBiAB9z
jEBTWv4WP2irXpVmIJ7e+NTXoMxzkItztB5Vrl5AJEqQ4zyCbeogNlwOfrKH2z5q
QB4PVBJU/oHho+o9mL9HyQ23NpRcjcRfXgGMvgT0P2C6ZgNfVOBJ5B14rf7ut85d
wOpNzWLqBGBaveT5ZKV3mBwkqlM3bbp+ySUQ3H2mVPmG0AB6bj/gEsAh/7raa0OA
o1VKlZHZmj1y+KhwGTDI+0Fr3swe1hqOecbiEwP/txsMJoOsF6Ttio4W6GAQamk3
Ml+s2gI9zDRXMXJB0dzamPuwGyN0//P39BJysPi57NjL6zlOC/q9kVI2ugLhaDtf
imtQ7LmvYTr1uYHJh3HBwzKhQXVwWKZhDl6jKySE31eb5JhSDitf5i59vEGdgdwl
HdWBWT+UzZDQ6nm3ZTfnOeC1fr0efjvM5QSDiRygSGS19+3T1lGqUqZBBtj/54o0
7jJ6A/qsOsBegkfVmmRJOjGC2OC9rDXg9NntflhUcPq3S2kmWx6bHc7PG9wIAug9
8sIw3/t718XSCXSISSO/Pxyi7aMuj1+bChrPxhJSLHPmmvxaCo3eilaY69O+b1OV
2bwo0ardqA8QqjCjYo6z9xFmoiv2r1OnO/V+xMhW1ENHE+hjvJD2aB4lgEhx+7qZ
nKXN1KczHrtLVGwFt2UdqjRCF2LmE+3V3mXXuXED3guBTJDE2WbsPdvZzFg1dDEj
Zerm0X0XNz7q3dNw/hs2fWcLpuwhAu3RH8C0GQJu1TCUvVjt3oZYypl7f89Nhwvu
+HLX169q5Ozz9gOLUwBWGscSsKASTgzJqd8SFUvujOAbfx1akhb6yLSw+LEQwY0y
oIgwtJhZMQOpnVO1PEcLjXtzBE42jOBmHFI+NmAzsdL1bfIu7/Gjc6/7f/sdsl6a
YioJbAGrWZw9o4iBtQ1YjeDeb2NLzeKJRgzwnFdWSGk4kJFQyMh31CcUuBygrY2x
iGhkpHgZNdoc5ydmUqCH/SDNjl4aWG0X7vBFcCwQARFJd/5N8aWuytaWEjCdn/ai
SY2SNrHlmm74kPo9AiMpiM/PPQ+O8onQ/+tgf5p3RLSd1UEGItStdQxw2DUSRwsp
rfwMugvGqpdvsQJUH9or+luAi40///GtS73FlLKr7F14cFQV0cTJ+Lo0BE092z9T
wXfu37tYMMnUzFuZxO5y+KvZU4Ubhw1AD35Z3ZJhG2xReXZmXABmvf9oX6VSBRBV
Kp0kdMFUQefdXKTQplgB+W7Rt83ytTPaY3lvdyCPkzF9UvTBS7AhWedlSxIwPiZt
uliqaELi46lcxhEJeoDPxqEi+vQRrWQj8rlMxBJ0nI3MxXcMAz5r4L+3FxBZMs37
1Go0eAT3u8BwrX/mnwb3JllgPV4v4SVen/YPS2BkAxrVrmtHazx4zyEnIBOBk+xH
1h5vX2qs3c00l9E/TQEHRUHSmOYJX4XtwZW4HaxeuxYKI/KxbB+6OoNTcmLk4o97
lRxWdqVAosLiwm5flHGINKQNcFpbxRlXUHf1JCoi6H/GeY/mYnKDt9xsV5SbIhBb
/901JrPT5t282vUOWVKvu6lrbjPAKwKd/+Yfl2JWy/uC62J/vPylwcvAyN+e765K
YDEbrwNyw0S1YcgoGrplGR8deJpC74i6MDYeG3zCdysZB93wLZJ3U4XA+Y8+DNhj
JYCktvuQ0vklnEHj3N/n6PnpfYnNz4YTasQK9Pk4zV+C5vYKHhHCSsb7/KxRZQg+
HhxVmxApgX0hE5Ucqyo4ju3rR0d9NE1oFjcdhj8sbDPMhv5IYUTgbPZEh5hlpBpY
lxznN/pg5jfQWeMz3wqj4hsKTY8y3UFM9BUfXB9IAaGOLh+V1QcgGz83MhTyG1Oq
cdMdCrSKDFL9uvAfHGmRlXT1AOatRrvU5oi0NF9fislA6u4KmECa4GSROlTYzf2a
Qgqaybwew5DAAh/5IjtkXrImAIxwt1vasY3A9aGH35BsHKtYsIs+4lxxkCp4+bZL
mKL4G/Alk2FTTf5jlW55Jz5alMdd2G0DjFCDLYksYooJK3Haq4Sd9qvwz3nlPat2
rjBmzAqK7Pxef/5JLx133Xhn6+GUi+nYfP3i2xAP6FcYsWC3P4MThPKovoL0hY/0
Ch9ESXBcKIyFjD7aUQBNxcf1Sn2bZKMN5v5Q1j6lnPzk7h8PsMz0CfsoS4iwOYV2
VpQ8jotxWofRL/HFJHD2ADlNg/8c2CBpI/oFUnqFDwD0gapoziU4cGJOe/OEzAvc
RYUSgbtrq6sNQ+gRNwRBW4Rm+FbTQNlfe8yj79UAICOvMFvz9bgjY+QoLgI2S67d
eFodrE/lO8+uOA/AHG7j0K2yX2IOnA4RvUehUpC6NG4of1XcAPy8nVifa5LE1Ens
jxCiaTqfuFnNxIrfl76mMmagfx2U0jRKkfYPg054k6K7Kzw7gQ9u/Ue38rfFIuTY
G8rq2qYepplhrQ7tpCoJLLprgRzFR1PHyf2zBxvYbZjOn/R3Nn5XF+I6RDi5TEP0
I0Nfp96DjYAlHogxmb+pDOckEF/kb+wKs4UjxJtWa1RSLgPIVVgM3KXBqbEavnSD
BQYm1grhLYdE8o1agHMg0RxJYnElEJnd4+eKsT9sDNAcAdfEqohosvEh5SiuXzw2
owXjbiQFh3KhiaUoeCB+HgnJqnsJmmemHfDfZufJIlTvb0a7jgjjZ/kgjwSr+Qmc
arYky68REF2Ip56KhDlBRcASPjPVs2mtFpM2T8b8dpPkUNqqKnxu07Wu7WFAR/K+
M+w2jS6xU/ZwvzCNyPe4aX8XjTFodmTJSI4j/Dv0adAQ+nsFns6tbZgRZITsJNJY
45H2anRbf2z4hWxrR1azukBtbgAwj7r4H82unpFENOCft1bPzEAW5jtIcYT+EJOo
P6X7+I28DH56E6QO0b+FIEkch2dTSUEks/AIjJ24FmCk/2W+LF7eOf1wrysrzYDn
mkntsbKbD01Nx4IGS4SdxFtfcO79UhWGeCl0eNQA47t23TOupkZEE3152BBNrQHC
3fwEvWLDGWP5n+SaDepJHWsFrcfJAnYdDUdVXDhidk1DIj5AskHmy6SK+CJ7NxNQ
2TDKIdmN7gvH6PF5wqCZiKVuq2N+UFUL/vxYYvvjTcuJ7qv09lgRp41HqwCPSMKF
XHgmtdFzkZZIpvEcJi8SidyxnGEsoPJKpu8nycFCYlTCUufl3i4RclvtLgzenK29
Sor6+PJ67ox4/5LdrnXokqiddTX6sCHKz168JA9YxLlW5JM9WXVONqQ+YcTvH/ph
TxX1quOYha6aVUZTPaUORm1m2hJrOg30kzK1hlfqPNZ/WXKI6jy2YTtE4/cNc7m1
4Egkm6nJPtcYYVVQvCICJMYONXsGK59dqukrxVQl0ln7pP29vFyhNNKBxWPLBK/W
8Xa/n+ZoG+55Rri7TW8/JzPOgIh+NI4lk95rCUZQQidLkP2BBInXrSQ++jdopyNA
zUe6V5ZbB22xbMQxeL/dxz/nrqlXpIjGoyY0K9wkwgMYCAP8XzCxQPVyPWrpW7tw
TdhcgHNA8QSmCecsLQVo/Xk3TEgQUniXBGP6+GkM9c3G9JllsVHskKUUB8Ibxp3l
J0+qG9Cqr/zcU0zbPH7gpOpKRbJS24Z46nUlWRg3h4wc81vY7DnDqfasf/RXKvfE
Rn1BJKZptQW8gNwiIhP4M4WS5fPZkNMho3lHYovk8Di5F3SpOnL/BtpAEKSbnrjM
m507FXX9WhBCaTnziRgMphaZm2IW4JV2zbvy2knsEp3u764ePCYN2MLeLBDvS3dw
ZxzCQPx3+rXsFDcE7Um13hB01iFuMIJZMhKmr0bVwMGdZ1j8VHRqcpjUfSLkoZX9
Je3EoTDVYHw/qpQiFGRtCj1dQZ6N41Sf3voNh/kFpUZJJZnETzspd/TeYrlA27Cd
eAUrTC7nCDlHcScXqGEJCLGGM4YNmvkClzi0K1YW6bmDAOpNoqMIhU7cx1xz921R
pmpT+FuGsp5F5kb/FDcjJCSjwpn+7cYKP/e7LzDPPYwHdu8ISjl2ZGgKGAxo93Lq
Cl6ANZUHEEy5r4LipJF53UedG+geD7GvCk01fwdQ0ipHGSv2GVRPo+w+G6V9Xq65
oKofvoFHSYGldlXzS0T1GtVHnFKX8L2bnDor0FrU7TAGK6CmDG9SGPvSHIMuNA9a
XtYW1hND3wWwDtbeiwna0AkxybJPpfZqgBONmH7mlujOr98C/ZZTdXmZblX5eejQ
HZhsEi9jFQeaHkhfZZTfM1cgZlggnvFEVo9YIpHFPXwTW9tqLI2PRWM0FNYXngsl
/OQWFuu5UuNQI83lHZMzJ9cmIuwICTTwPmT1TESkVW/QxhUsKi7LQRUNZJsB7a6p
tbiOc2DrtVxYix812CK6k8rHDxN6KhbrYem0FG/M1YayiwWZIMfuQMy56sLmXEIh
C0x3Isj/SdnI81/aJp9E5hUHxJskv0e6tSEua0kuQPVXpOSwbeoGu/uUKsUl7i3P
8viQcmYZXzzv/B1oDqz002SHlulKCsCncSGRSxfASLr4K5REzWfV9Hz+uwPj803L
OId/jlOcuUM6pQRwfsgHuqMEylVFssSQ87o+n60BtolO1cE4U+PA2niJqiV+8czP
0NbJLiO9EB4xF43UDRCFy4vcKA5OOQjneSEgshK6Aaj+VY4bBxLv4VHuz4qdaHu6
3Jio0y3a9waynoBG2nqXI9qIPbrMSHty7QzqXpsf7lE/khpu8OjoT0NA+7lNT7aP
hLvo7qqop7zqi+aso4DANZEM2SGwHQaPCa1QrYGZHVQNyExOKkeRVgQs3j7U9aYz
Kc0F/FDOXajN03p5LLSlK6GB+GGl5H/V1cpapPWpHfbXNoxlBCRO5jeqby3iYVb3
1jVGphdCjDLkZnxN82FD5KMy7Sj+hgPMs2sAFH7HtM3FJ9+l5J4NjbgF4+5TUOB9
9raPJ2zSSxOum3izYpz5Um7RohDjkhI88hwxe9pS7ZVaXrC2ghTbPrBh6soLWHdZ
HcLkE3O6iuyridHyYWWDJTBkcNleFr7AWha6zLRTcZW3kpq/iy32XP9Dady5TkKU
HiH9lhlqtKxsDxpmEQ9Knvu/81v13TrwdcXws/Xllbywg8TCAqLv3BX2MbhOemuF
YMQoQtIqWGskPrA2ALmOL8LuxFUYdppyOSsSVsc5ZZfJLl68oBtue8baJZ87xeTT
Pew66uctjzS+semDJQei0XRXeWJYE5G73Nvq0X1iWhVLChuFVPTnKT94L6J+kWXm
FtJ183ydMvKnqX/hNd71qiYlmH4h0ab6srPhXRpQaUcCAGZ1gx45jPcwMkIlEXpj
BKrngfKVZCBgAMn+QXBzj7gxjxpOLOtYe4VBk9yftQ4stDdayyyjReDFP8p7uk/K
0jgmtIFGP889+4doxpTNA9tDxWBs70gbiKFw7uESjvsJNsUoS0V2+j08Hht6QhDN
7H2twUqCvoulrC3WSM+GVMU3L+84kLOhjEcuqVV4jmt8a6JwtzERVMYC1qwyYRDO
lG0plHfU1rSj6+CwqlFmAK6ItIKcAVYe60SMuRyDe74Phn9ECZYylIhjHFxtoO2E
4Anl4kK8+GdSxXblh9w0OCxjkswKTi3DUAXlrH69sI6Op6ahe3Q9GlaOjhPH+8A/
HlIL/5hiHlPh1Jg2cZOHerX7mMsBT5pBwcRzYbIg6o++f4D03SiljQsGHRGdqMfW
ULOsG5OIMT9g9wXVk2JK7YRFxb8YMV91oQ188l3cq6418XUmVs9rjwrDm99YlGXW
gNGJbCBEy9VYLIG6EghjQ6VvD9m5KggXZJktDZgJ53rZdvFJf0CF5pseCqmA/y9d
cwEKZlKhjsKVbOY0p4NK+BydKmWEq51bZ7ckPnnFMJ0KlGpgE6XsnAks720Inp+Q
vtVJUJpMQ/j4yrl9Qf4gdWUfpjhZ5aoR6wfoIPhXX9UZFotCBBVOUk5wWVBX5Tq0
4d3hKIdQNVjCfWbETzNJR7IMkz1bs7ezlQNPHW20m2hZ+Y1ZCIofIkhbzU2QKrsg
UjVa8kVFLJacToLQbk2T0yNb6C3g2YO2d1JCvd7kDaTYYn7qaa3PSwWMCPeJhsjW
+7uESXooyhcPffwI147tmr0KwvDnh9i8IhiEBlH6p8qOnVfxYlpMFRTRyXvvPHBq
++fvtzQtT6Acdzq/v0iO+sscWiMNRJZ+efDLn3dC76pU4RsTDy+1UC/pbzlFTqdZ
Zc1ftgITJzu0LxqiedSXgy30tuMKAUNxy63hSgiVR4g/yCab7yvqPpGXz0CoY0U5
uqDIeNN6c6T1UY6Ff0hihoZIJw77WqXzcJwc21+g+FZ4YBRhb5StsrG0lsBvMaow
pZwM3FjVMqKbdCEx7LmtPHjxYo0smDfmyrBpYfMD9ZRTGTBfV5sDNm8pSrcV8Ty1
0XzlrxgrO/LfhGSpRKbuk9lYz8AL//fM7E2/5YtizsCEqA9LfM67ybBhv1sFqljs
iu6cdiOY2ufoDpsGXK1kDC4zbomgMGxIMrkS+NrFd15CFO/1e+SruTrmGRCqh1Fm
xXsKJl12VDXEAlqk97maf81RN21D1m+c5LMxuday15mXmbSkjOIE2285geuKa4Hl
++zmyy2XNngnOOE/lxyQO2ws+OvniizAxVLRm5tlFiGWGtIbbY7lmy9amHjgdCHa
POL+jdl9LMQJWfX2Xncd3MH5vVunyuGvQ2GM5K85U7FHKlLLPK23MwxbDJTvPkUH
pF8003X137CL05wxH1oSfszAiaFOLct3PJqvLpr78WoKUODOfpWCP71vy9VgLnb9
GOiC1m7b3oCle6nEUE/sjymAcpeGnB4mFPnwdMFCcafukPstyUYkrTjc6I+vuBCc
WNLNpDZjM3SCR5VjbIrYC7rdD7qNfnNa+9i8cwT6dBvBsi6kt8do3ls4scUK96wD
eyilTumNs58kMOtvL8ui+gsQE8Tv+54K8BjEgaaTWT0FfRTBBshcn4sJrYW13Zbs
Y7YmImABZh2DIi7/PoXCrLPBk1gFWo3e0S1V7hYmxVfU2Pv5BQm4+bopmTHmGsvH
fAKGzC3B+dxD3SpkboHGBld9j4syKGpgiTyp2woOWXs9CdbqG9L/aclHz1sXAYFR
whXJatX0hlXhxAXPeDalkyWhYQ6T6hXML/tM/ZY2sMXYDL4wJYDsQTVqdxVuYn0e
VDd1C2l84R63J2Luz7QLOvydh/ZCDdjQuAHnfZvIZvMjPS5gFH1x2Rb1SvqJg5Z4
UJCMV55zvaskPhEYS891Y5gXoQ/m+wcPL/BNoVaSB9C+bLqyKxG4JgXIGTrmRwFv
lGloDL3jyVxzNluMI8E0LBS0WqUK5NuH9DhNxwy2hd1qfd3sLdh8T8P9oDO3QqHb
hC8ndckb7xLNArvKhq1NsE6IGaVeuLj0flGrNznI87wMCYOKNezwNEY3zMWq7X60
qBWQng06W8aOeE9mIa/pRUwF+XRju1lOsZDzTndrRiael0rQDe831BnAsnMTNudw
TxzMBmyS1AVXy3A5t090llExj3Xw5hLLviNFdDBajbPID9K7sz9gR/mtBkhUvDXT
QOSAUDmp7UQLkhqpHRcCreaTs16xbmaVL4k0fNkkbbSOCJpSWLi4QJhY9h7xbNPa
lwYOdG2Pod1YxqGKl8UTjwjcwBpjAA/RE+EZPlfSfOy7i7B5tVUM883j62rdwD9b
bvpfA1PaMnj+M/6Ao8lyY5BRMSFciztBrnNF9npthUIz2GnZHoJSYd2yfVXZY+Q9
3fp8axtm+vV+P+ayklEYmNO5FlI5nbN7VctD6aV8R8tGTdMm9/T+047VgAp7z4Sg
+08rUgMnG90LEt1N/2zusCQZJA4TYN/ECUoMIM2x5f+v1xtj3f95NEJtWC6rLgiC
cMtbbZqFo8vxWwUfQ8l+OA3et30TWH0TtP8RWlQaPVRhWWNX1/v5ZtjMzSj1NO+8
76U+RCpxEtU+JLJjcS4r8D33DfQPeL4ubCaBo/I6E7EaKgsxrQVGPSqc9oxiBBkg
rYFFaP/E55k/Tb6sRI3urMHssqbVWCVUYS/AsXxFr/EVAKkaOPigcEYnaCizFgNo
TjXTAxooUy4ddTQAbP7opU8T5bB+g4uWyOjiZAYJZq98fvSqxWa0nHwT+8WhGEtT
nhur7XnX6WzxnxMwWQTRAWxoISPx5EBWYp7w48/tqKzh3t6fQmrR4uwTzZlbdMtW
YCmWnKI9N7XTuVn94QrVej6MWMq7l7Hs7Av+XVlHBNPgBd2yNehyRJQQtGmoKblW
g+PxY4fcGcRU9y8EZwY5JtustgIPalOsRZxTaEwYdRFM4sh9I+sCe6d4spkTOFOv
cFmrJCfd42QFvVgpFKHQtIFk0hz/fhXqWfZPm2curUgOc5fLPa5P/qsrXIfn3ViR
uIHQpZgpeJXe79aEaptsn1UwsfnvihCBfBuX4KIWtwPL1jxwsu9wls/kPEmDYZaF
IeDw+mYWnkbpPqF17SdMKuMC+bdNmTlBATwHM6HuHBjrfjSo69PBltRE7OXS7IxF
ZEqnK4rCJ7dw9n6aLKwFuosdlR3DBuBUQsBPH2pQxZHhURzzczGdduVthzdHkKW4
vJYyPFY3eY1vVOIPjw/oadMSpQeI9e7BNrkhI28X+BYkJ/L5uKwexvfrA29/m/Vb
vXl1SV4u9jD+XmYcPKVwmuOiYhLaG9kG4YHFu9wSsZqvk07T+mOhJ03i9XMw6AUM
MW0vprix+JPWbSduPq5yQmLS8SsD0aE+myR+m0O5yE8iM+06hOzOv4dqqhtM3t9Q
tR2d2V7+bF/RZpyZvmwwTXt0TAHQ60oywUdZ1xgik21yEtS7UpBn9W4TpZ05pnKI
xbDMCxR0pUOTkxmNaWybLUj9VtDKpXNIwl1swG61knY/Tkine4y4t/qTJDlDLm6p
HcY3ZLfNJ+o//8ZWkDhWMydQmwbf8gBJusIZ++V16As0jCZ5WO5Yf8SjkalEIST8
mzVyEIl+fWM6LGvWnF2nm53t+8ARZZyF0v+tPE8OXgB8mmL8W+/7F8Eo4I2tM9Ud
P9vJoq1swCaORrDVS9AsjvehCmCI25sxkqte2gT6sirlbuSfqCK1VQyWRGYsYfNN
LGcyJivzyOZTySMIpVJZlSIgry4MVULMFLdLh3s9ALGstfMmnlk9qJRfq/LXWxuc
VFiNK3OuYtYlfQ6h4dQ0Fp/d27IEEHM+4zigBpjQAwROL7srchkVBpFwqrlp/akN
9z9WGxvMZwTohYIG+455qU4LzD2kCLqTd7pjxY91SlJihIvoI6nxm8bjSV7qArY1
DCDWxHDcpNTXTKltnSEy6aQ/NvOgHpkk7M+A9nUxOuMe6uWK7z3NLiQQNiQJYBCK
2xj1whwPj1T2x/6JwrihBv54S1Mfuudy2/V19v3NZXa2Di1dWmX7oW7iS5Fd5fxh
7yiuegItOXGm0Kz4h1P5XewpR+e5UQOQPmv3MLfsTMoWOUSOHkXR2psWyqhwz4WM
yrGXTniOC08/FjNnFf+i95dWGJIPUIbXHU7lkwLhcXVtlstLs+49eUN87OQtHyjy
6YBFHkZ9TufTWh81MUoZ+Olii6opHn9YAhOFL8DOboKP0pqG76nRcq2sw4BoWoPX
CkOzpBKjO7apUyrUf33bbPmZb6DC3omIIF0Og3JZPEAGmMynElfp1k9LsECCV1f3
uTe2qTfPQL58W5PXzJC8mB69l0JVzqqgh+UPk5ziDcPERHfVVQ3nHTIHoB/7OGH2
et0azJPhPt70Ovpp9jngzAs0Tj5oEeK6xaXHnzdsZCrKPQHqXCmYD9ILiAQBht/B
r1NOYkXt0hr+TK7/cu77IKyPIJq+L2k9/BkIuun76hGyAd/TX5W7XgeLwDRXtotP
YyoP8kXTiBLe6B60/l7cayPnc0lrdAe7QZgOZ3c8R/06c/fA3bp0m6JuvsrCUbgS
jndcRpRVW9H+S2nloqccX1aaOZZok6tIHnff1GYnMcPJRRORqOs2kIh7PkwskDGZ
7F+SmxGHMKobXuZSZ78jnXbTBV2vDJHkNr/+fCvSaTO8Ml3Khyd+cJdWnhaceVPk
CE8bT17zDAH785EDPNbIwGppkD9+bXwt8B4Rc1wjfQJbOYgllvQmkjS39eymsYEi
PSAAzRZf90MunRGxvBtMp1Qyd04oTplngfxSXYgbHGg+cB2DgUE5Ly3yZ2xmxS4C
Gq3o42+I0qPHidDKmsPHk4j6Mw/3ILsARrUrj68FGmpPYrHZT21FTTYKHnNk2p2Y
ubrBQ+5LKdmKAvNhSwJfLCXTsIHW2rglAa1yJN2ZOyttLMu2WHeiHLeXSrjWOEeE
Cb/3zcja4H+ygJGAOgFl7lp5hoUJZJ4zkirhPlLXAQPf35gDkt2bVRNG/gSEosPB
JxKnQMTjpcw/LTsNRrAszaYkepwTXgkMEtfxW5BO2XJG5rJ9Ks//jDciGzIDsWlP
TozDz0KhOJXREzHY8AMD3fcoAP+bBBgnNbe918EKfzOaAATe1jHlZdQvKnrNaaKJ
2tnT9HW33R+fWOZ9dYcS8WhVn940b2aWSyRVO37uXnGsZU90fOk1R0Af95EJQqya
QfFascssF75KfStne9NZDSbD6+TFUmrWDEFdxkGlC3Fh4iNykgYQnH+qPoswCXjz
pW/DdzTHP94CqqfHCY7Rxhqel/pa8c3wVlN6ZGRea8gTanyNQOwvHb0sf7dsV43K
0TUwtoPPXbU6WLbOpZY7wBewaqeomZ4EX6+On96nPO4FUZRNFVpKtYN898Pl0Qio
B6VYaZAWXEAJwD5mKQXs+TSNzMPmK6POMU0Ds9Q8WA1e0Zr9GXpZdFQ3uJ5u6HhQ
SFdSvPgeDNYR45jALR66E6NBQzpQBQApaE7GV4utH21QR+O0SL4V8L/tLDqeFMCs
NR6pA6CRuqG7vjTT0E+GFG52WaUiRwaqSNKcDBqoXampBdmgOhN+tmBbjPvKLTNp
99QRi/wJyOugJ7KgN9B1vNOO3W78LKxZ6t/Dw9vn2Me0uSKixuHriYUWU4ozcjjz
520XpwIiAUNYxsweRbmWq86Uaitsdiuy92TesexRG4ofI4sv6MsKrqsy0gYDuq+J
pKT6SIoO0DOiNAPH2BqzjCgN6RQhElQHW7fE2bVi5yS7sZjvIW3y/dvuyQiz/T09
EiMK934mKIjKpvk6/CcP6RAMsCNCsSfB6U6vn8nu4Uz7m7JmMuNCDcvGwZJoVchE
jK4FyrhsKMPAdCEtQUej36R7UyAIYpwj78+aOB5xFf5FaYJpfzkdqvWqIzyVuRbB
70NmLN/ZfXlsab9UvjlwmtTCW+Zu3AqRqvjikeXczBhOkvU6qtOXioBxDLtdKzPj
yPXVaqSqFTbeRkvdGhvrZGkV9eNRKDgZuP+WgaGm/XW8iP0btK1rENJ9+kufBu3Z
5dEMWlxEpqT+RxxVCCHbsZVgI/W5rl+MqQYBDJsWH6m/lDLiupNCxTWj2nz6FhEy
C3e2CLN2ZyRdMkRtM6FTNv87mhGkibqHiVg4xqBpA6oFhWTkbkKvT6ZrLLUCurqr
jjnqHbvh59lGbd/O4ClUALqjsTdmyh+Dz/PYrb4334YnbLZZMHgP7uu6/3ZAzPCq
aQQ9TovOJT44tUc1d07rJp3MSZFrTrxTNeedRH5WGLtZ6ACrOP7vq0a7bLKAkDw/
W7nyn6ZJC57god+503sSPhNoxOSlAEi56m7dN4MkZ1TecGYR8LCCNatTE/lplkJx
ny3dqYfzmkisKss6hkHqP4gdIZkzwGsAyomTWT7gJ3j7LsESgrZe2iA5LteqWcF8
80JEBa9wdUBwjbdcwW1o+qojvVAibCJbP1bFqv86XxG4zMn1OjoVqmTRSKrZs+X0
mLb1XO+6FzArABGmPDjl879nwYwAqQu6bD8D0qlCEwfsF1BH1GpkeVTDuPFJNFTU
QMLmbxaa4OhcUsEgDiOfXI9/4uqEbCjfbwd7Fo1683tEQ1uh3FygwiJmoH1rbotb
59W4U1kPsk2KdQssB0/pkaRaTfoAnyiwRnfLTvEsAxtNBRUbeM/Fg7roEWYzgBhn
6l/1KEsLOZ5SyHvB6cnKtsS2srOEs4LKIg7rHQDTdqdqbBWvysQ51DR1eYHx1tMc
MOZdHsWHOZWarnOUKxs8BSnVGssLE4+lsIsOuOciGgruCVxmZTLr84D0d6sXOEht
eXuYtZBdmxX9To7snNmmPEiu5ytuxqWhP6qhLF9L0oVlRft/pXd5SMA45NeL8/Fo
4zOPIQyNwiR+FasmKVL0b/6vGewhxEbU4km0FQOvyY13AJv28tYNs+YpROCn2c7K
6c+SJMrwoJc7pJzL/qBIZi15uiNBH+jmMI2OR+0Gn81Rb0FOk7+ZSO0mnWnOBMpO
XJxSTLoxcmIztdLUwCIgrinA00H3BlVsvJ4tzhQAb+UGoOf1polircpkJCJ8DiHZ
qz2drawoaifeJJXM49SPCiD/G16zFYj2L2R6pO9qa/mWtFK/81YxJiH3JR4qDt4r
cceadpeie1+PnV+X8alTPnSOu0pJpKveWDzLZUD98L/a/wBnpLL4SnTHgt2T2rVB
fZpT/DZsiWX3Rv1CudyAgRwfsMUiWtYD5Ngw0afacj+3Vnh86GZfM8R3pctuSUeC
6Sqjj6MXqwCrUs9OKkTFx2C4pNwlH6MjbHEHSeZTEAqWbcF9VRKlJESzIxF3AtXU
mCxfaKPE8Go9OJeflTE2cO3CseuEfthqoZDwCBM6VTBT9LpLnr+WgB5t/VEf9aYv
tMgOhQGB0Vmqm4IYC6tyQS/1ycXcnzrovrsh0s324XOK7v+87ZWQ0woyoDiFt3+t
jeeL4bG6rn3JiUEFzjHpb+4WKd06l6b46SdmqwvTTvkmlXk9ffR3xcjuJ6NBZ+A9
y1vooChqTiFox8l0qe/pYCiSFM79zot8uVHPFfg5zDdVgeDNDjhQ9UO5h64X7xAh
F6LQcrCyDBqJbPNhQfocRYouD9EbUeYYXUa4McW8sXIEUOS51AAD9Q8c7H3K2QbD
4fXl4a3mZmAhVwfdloKRLn82hygXEwQ/TGzIIjQeVlxmkfING93rqHyx/hpXDgZj
Y3tEovwygBljZsLr3JluJuwa74sO2j5i8SDtkkuIHrc5KIKSL+XUsjTIpSny6Ibu
mETgq5hNhQgVr0GrELJQmSgK+VhFFJcc7LrYTzUKQqgtjFcBOP+oCf6V7b1gmm/i
gUsu4bDREwareWXz5sYPOEqD8qEAVH/naSobDX7bBF3nCCV0YBPs/onzuYJtTxSX
YNiues+UVS85V/lpIvWCkKgqbKPi9XACsoVGa9NVXVOLrSZvl7NVFVwuyOM3wNin
B8aU5px82h7DS/5QkhDuw57Gtr75tQwHkMYPyzbvuVW/j0pus92qhgvxqDdwsSiW
NM4wzcybhntvXdwiRtlZbAQVKQq3VVqDQKulof8m0OsxEhH+gsBVKOb6SEqalyNC
r86J8Msa2oPjLetAs1JbVKjNh1qE9nNirvGQN29UMGruXcrDp62dArrDGLkZzQps
XSXOb/KlE5nuMiI9lyhJBdA+RHgAyrHM8lUPixah3IAu8boyV5HC/byibqGBWk7z
rzDuJr05HqJGiYmwHz/lMjKdCLxtFaKnENEfXmwlO8fMuSXqA3Ne4XS+VKb/dTa4
JvEtkdw5XbMTZCoV2IyVkZKRY+9v7llbaX1XRWdNH8jlsy4KGbQyUF0T8DJzWXeV
0ibqP3UobB+jogQLaUcbxXFzGIyhlK0KrGpdGXT0Mg7RqFMzszS/Vxortkx/fNZM
yfJ6mrOUo5ft91+bMvXYeichTCDe73qiTeJleaR6wuWfAyJUhfFXaSnS43rxj2T+
GBE4vYbDwlYlj+tUhU25KYYNBTKYDBpTacfjUliaIwZDumCS0MTssZChIAHk8Z8F
xSx1UNWh8r17H6YnPEFvhSB7CDq2mNx9AVvBDGPUoGwSKzwhDarPLFDSHvUpsWhR
tEZLvSqK1yH4Zn0wx0nldhapQOAinF0oYnM/Xrv/NLDTwJ68g8ZPkNLmdTdEk/9w
B0OcQYr2U84TFwQXKaUpbM5a5/8cdLIQ1D6KjltXUqlvGPDEimjwVj6WR9SBbEUF
Rh0PdDrKyyK9OGSKAL/Q2x+1b4LRO2uaies3zrSG+7t7Q4BqGLcIdJ5zSFOjBjFA
XkqThqpGnucFGolpUejyYhbc1Xj6QYDeOLjDtDjt0inww59setTyLJd8NZ3/cArP
TkODouPPUNuDsjuLmZKto22mQ8ipp35f0yoe03QnhjGQmL4C9m+FsbodaRoBEhHM
qggzdRwXu6X9f0eG6m/AWHuTIncWHhtgj05G+vNhqFjJTTD+hfrXYk2WPqLrqffi
rzAwKKaFQViSQZBkvpPYwaW+pSoa7zN4xCrAQPEFw45Tc1d0KNUc3huyMm2Yiml/
MfPdD5oD8i0eyeyVDioyL2E5hb4IJSFrsxqnOvomR5H1N+qIJfLYpzNf0D4MiF46
XLuyNgYSR3aicPYz79LPtXWyugHxhJhqK0Ma/Gu5Qi+krOrxwo4HXTSOf+FLo7lx
2XdjHG6uxa2RA2YKgfQX56LN1b+Atq4TIDnDxSjtHRidrzjh6Bka6bJhOukAokXT
AzHxJ/73burYuSJy7j/4VUCa5Z4e3nJtfqLUU3vgcgEhJgbTrKHJh0rwnZzWTQST
6IyZz1E49bKs1IW5sjlrm4zHVOYZ44aY/35Sea/eiOa8Shm43gUO08lK3ExKe2dW
oolRVXj2eO88wG+BxjJojGmeF2ERUoWEQaSGd24u//GntwupkUvzFmiejqGtRuFa
pFaRoTB91tg/qF/VuEAaK+Dt31Uh75rzh612G5/wQIgv0fjQmpVxdTjxuPk3uzvB
yNmDN7HIz01mZ1TBPeDMSDqMWWDxY0yP6BJxf25uMbvZvbkqSed5sn0yYYwpkVfY
OzQMP4HZIj8RpWAnVo53zW/loOZZqIe8FLUf2Oxlx35EWhE2sSNsZVERY+rMQxw7
zynLkrDf7Ds2wq6ncfX0GwNq8HgQCLpCWzTMx7muRYBcwhe4NYrvWs6bMBdy8gya
2MAFT7W3Zf6nF/lmYFpk02/VdZD5nfFERCbUALnsWufphvi+TVm4ErkYZseKBbje
++7occw26MapOMdmw1ObogmjaEylUMGXRJt/pKFXE01GJoZam/EGAZP647ino+/7
52O+Ubb5yNVcBXhqT2OBTOc2xlswnC/cm+2qssVop0yBfzDvABOHmv1hcCCXpbym
cilAql1V1rY4pJQ9VUZqqz078fWM2sfh0ECU6qg+YcCMXlRtVJtVlS3bRUcaY+ci
OPMn9jEw+bpQM+/2v/5TxQdz8ULuSF3IYRbMa5MNGvjA2L0QHzwXDMW0wuqq/ISn
PE2eotTPc5+Aatchtv6WhqI9AxhjC+m9dLPUnGl4jRcdnCHVkNJ+uLk5mR5HRkNh
Wz9vW8wRmAGf85vGcTS1bXGNX4x/rWMSwV7LjuA0yZi0CdQeCvWFmwKXHM52p3la
78dH3rg9hmrwL2ulADcpPferobnl+uMIVtzwcQz++5dKg0zw2XB5lreFmxGloPm+
aUDjhNnUmcy1/k9TUGoH/ij46pnMYDkgSqL3/x+i0f8KoH2f0aQ90nAEg34Mz0fs
QWooCdvfXoMimyZ0rTrWerFIkD2oP3wcwsaZuQKjjTp1iTobIHmlCM7G60F265e2
KJ7YzktC7v3bkeqpy1BiVRs7O/+tDHIiViu8kaABz5LM9X/oj0Ehhw595de4b/S0
02ZqK9kqp5FODffQFRaIdc0nq4qoZav3QcPTS1xpdm8s9TbSscZgdyfIG5sOgZG9
hq6cSowdyCp0F4YlWZStnw7MOK6FKkxpIRZ/Uqc+ArbN/39HwHroTj8yniuz+K4z
61yQS1Mt4R54PVPEFPtaSmXP7KQru/tnvLb8fy9aK+TRNYqLpxQS8KhKQ/DSqVoy
9kOvFLGOt9ZEzSsdlR8iXrz3WyaI448uJaPYW7B2s8mJ5RBujAPmKccUKG9YBOx+
iuQwXo5z1dyvruKMqxf5eUZw6yB/Rze+aJ42tKOhNrTmuYSOJoM1XbDUCNaYpwTp
SnCVJxVTZ5thiaa+e+0UQipOydqldDsnZBlWWWS1Bl+cuXHfczGa8ng0XFqfQxrL
hUcyslZbYumbIh0LyNy4W3dlKF/jWRDZrg+NJdWeK5On8LgFOjZiZRh1k0JGHbyi
0CUegyCeT2IeF9oQcxuoXYGxEoWzQn1JoFDHLgpZeOzpXJXtOEuHkD8Yam3jGBuH
CzkkP8/QPswI2FMBog44kr6QqBAy7EE4En9srrAN0Wy9HFZlQKh0UJ0H0OZlr63V
2TIDqzKueqcKbR6bVKIGSOGukI0El1IvRw0Se0UUvrVaf9LVOwqq6sPPapIHTaPN
ah0YGCdRgW2+QAdAsMd6RAQ11HAKTdA9xtOz4vZur4TD7Kn+a2bB5Jb0K+fEtRSo
4C2sMcLU5l5ZrIbPV0E7QQ8IqW01PeYRGPraYHOmY+va1FBRTue2B7hcOTnc5ogt
64lj3yggkSKpcje3PrU6xaeqOTv/9tlgMUgB7zM+RX43cZMSEQOARYdPAPB+eBhL
3X28D4GDuWwpDGE0Rc9Ol2tZJEMg9fuxliKOau6R7eLyUDbgApzLl8iAy/w4rZx+
nBDVc1gL4d9G2n4o445lDdn9fq4KWsQ3l1SXGAr9HLOjlaaYC+LElwYu6FfsCz+i
r7aY5fXGiw1GkSMZ3JQpFyFLUwGge+fjGTALwvEUPjPmQZDvG/E/nCbPT8W+4f1x
qdK4THgpS/vgNcXuk1DepakrC7J2sD+QUPcUnGMfYjE5yAQ7pZyfYJ0qmFSjMGi7
byXYnwkkxUZX7cssDe/6vysU53gqisEEpN9e1LLQgOlncICsMoJ1z7rZ6iMROxiw
pF6ollG01x7jMFk3bolkRIJTM26VEJfpWX6l0vqXHJKLZxzGHTCo3U/dKp6Y6Ye5
ltW+7OK1hrbTrxXvRAgYSIlgta3gXjoQAtsUvzezYPVBL4hFoU43cgC5mDmYj5mr
o/U5+csOuPivJWhhEAdp9/U665SyVmwOOS6rTSjTRFn1YmVOEa3gBpi29zxWnXbN
a+fNojMXRh4vDJi+9+Y1IFyqaKMvnGvj7+ptehmuHTG1RQMpflrbTK0109fBEg9K
9H2FlVpGg0nKoeMz3wDTkRrAeg2P9WH1kq+pC8l+LVhRYzYLlFjn4RAUhxc/+8CZ
U4jK7gcu9HobyHBiLxtwWLYJkNxYdWHFzcR7S4/p7wuRytv4a3VncgSr8bpYlmAb
xGdm9Rbhf0psC32EznyW0Ms43fUhzd6//HzpTxiZ1BLyS+1v4eZfuW2g7qawiWSQ
o5elXklmUjBHrMIzmI/7G9mVQLo/jaP0X3UVBNhEgJuZtls2K+MXo5dqasU3KlrH
EY/2MEVn0NDAnj0XvkhtE8oW23z5WvlvxGcGNdUsbVcC8qNSzrPguU86gHcGd2XM
rOXJ4l73FeansZWdY9SYDFHBmkcxWe3YwEP1mAvY+UtuU0zt1HqwJSg+2K/ZSFOl
slOJWbuDKVfT7pANNehrSyw3Tkb/Ef564ALvtpESnsFMPzf5esNotV1qQ6x08MbP
w7KAHFuVZuk4l0Bj++pe18pjZDLrUs35Vkb1KlPVR3MrWD8quUkSf9KwX+JYykyP
lHrivgwZrEJWK31gq5L4H98YS2j7SzaaFIAPaM9dXUIZQeZUkTZNVt7MecMv9utr
RGps3Xq8dBJ3+GtUsbsRLK7cBFT5KGEtBUnu5onV4L0BC56NxG8AfDfGZjHsf32f
patcI++4x4AHk6vJVIr6U5kthlxIhOrDKvUffleMtBYHxLjPbhlR6/f3TK8C2S6F
ut4iU8vzwYaCYuHSSiLUC2U5ijNU78fOSt4AGLzRvCM1CXfQGuqgqCu03XtDtLBq
oGdIRxLYp6ENKbGzAiy4UeZ/EVk05C13fmVWFRpI0GsBrm80BrIsJjJzKk5UTlKT
MYTa2VnIGZvX52qChuliIkZ1ta2cT45A7cB97meOtiG0glmLU0n8P1xvLxjtUm0H
+RSEEPcXDbgFVeFCRPqg7UbdFz/+hfxn3AlsXpvWxqnb2lWl1P6+T9aCEe7m/3+F
6FOF80YoTN5QJ37NaCvJcOppAZBt65tboIeD+X/Ehdn2ZmBx5DSx7qqjwMVv1M4D
zvr36KS4mJCS/I7DPHxgujHfa2jVWiYwNpWXJALH1Ceq0fVL9ZasKXcLihNkhGuC
SlSHpI/GZX2nLbgkZ0jGPgmHZatYBLxnM7IseGJdUBQr+WjTPu4tXN0LO5LIEc/t
/ZAHa7uV4Y68Ojc9MNIepAGnkUCXanW53IiFdI/6H/SwNio4ZomOzy8j2ccaLHB6
mOTf8A8dY/ItkaYmM2jhU/q5XF9sOIwxWcqlAldZuFan7AXBSnHPw7daOnmuJ/V7
p+URn7q+xs8S3bStGwEewegJrzLJal715JkUoqij6vUSl0dKduG39lLg993Vkifk
2qIEjx7vTRBsfwNtkZHbxX7OpJcNZ8bfjuxvZKMWOw5HW8vZC+wXiFmMGFKGsXZ6
e7T7htrFk1KvYPJ2CqYEDUcLVFQKtZUk29DNN7KO59OxQcBMoNBxqolIXQItSWmb
yTkGeIy9hufXII4d9Ohfqe8lh3yR5/UmKX46tZGPgtoQ3RhnDSiizqYBoS2PMbjf
F3tpgeShnWvAvKgKM6vMGUu/FYwsX1PpZ+cNeSruWzWLuJrg3Ob96CZIKISctNsB
zTMlDh7faBY9+EskJe3tCH0wTH/F0451u1IJrRAaz0kKUmHvBXJRG+qGNeh17cha
yNbd0SgQ+2Xuff1FPMKDbMD05sL/8OyQMLX2fQMDqYMw+ohRRuZYrELDC8ls7or1
x5xy5FijM9wac+pRMhlLUI0+w9qdQNmDnhdrmQTJ7vE63M5+qFS6wonZMKyfv2HJ
7CW4iF6VWwUjx42lU1PomubR7HJq4e9o0HF+rwatxRnhQ4+ncNtG+PqAS7T+yuSp
7i0ixsxdwiw0BBhuCXEywAiQrpfBA6Nyx/RBWMvhZZDSgicPJ6rqx+XbqKc8vEzP
GsqqGu9jXJxevyCv4WnKXGMTo0+iTgLbA0kElVyKZ2ZUgbpVEa3neXq8OK+yD79I
UpXd+YqnK1x9UIO3+RLo/x9JOm7B8cJ1IgOIVxZ3bt9HaMrOkreggZj/92Hvs+3X
1jKpk2y9EwmFjtMZjDO9BMU3DHDLK1ZSRP0si7rFbdQt1uMdnQOR/jHJai4F0FeD
gngt7ttPXuVjbU8bVDKW3BSPY1d56giKQCllbYnzlK2AF6O7686KrE2rQ4iykRyc
mU8wYd3D7FMDmbOjdkU299vJbbkcCbNQZBp0bvqSt+Dia4FiYeQ0DfL6Yll2ERoa
OdzxLldbuy7axZO7CIZAV3ZXdIa/CcXuP/yJfPoFBaZ3cOh7io/1ViTyASE52lwJ
zfn9pjsrKAC2p/acN1e/I2EAJGXzBtk0eVe+YyUiCJzeeM0DtI7H6cKawJKPO6ye
+8jzCkv/hJY7NrUPoszdUtZ8Cv7BCGZQ6f2ciL8jqijGmBqTp9WR/PFBxtatHJlV
jXnp/WkregeR2A8Imj3PCCqpOi2CV9ybm1KAH126vS213X5/Cotyir8Im+u539OL
kWi5rQj0+WUnQB/rDTyld8dj9c2q4cvClSVKj6eZ4Bm6UC3goJvSPG4jmJDW8B5o
ZiB05T7hglf2Lq1s5ysvi7XcLUUBpf9Bl13HHRsYT0qGbQOD4SDS4xjccU4Amg0X
EGsWNbEgrN7eYEqrPpdQc+d2HVNoKdHrE7Ap6Mxf8HqpV6MKCiV+YJ2e5LX18yJt
6C3dXq7EfignNq0uvxiGsFdEoYjXJyiT7wuzXxBF7G+uYt8MiX7uNZNAYJaCcowx
EIM/dLCotwc2lAM9PeX72LoEDTXBIkZ//xygV6wZDsN+Xz/uLOrB6ohPYGfyCsZo
x9mbtu4vIclqk1TiCjoJ1iSOnMT/2Agms3e1IvPOVqvmozrEivsBsNJtOZX2iLoV
c5vjtqNIUgyeCOUrDYNjyTK+up9Y5e/7yk5PQYSSCxuLC8BewB7tsGPXlDOQACdh
Uv0UFHqryNEAExlEwHwcX4CZbl0R8dTWEmIahkPLqLgXU3grCvozE9iUlO9BFLk0
7SJUmHDl0eIP93nlBZUvn+QuJBdhsfJXrI+Uo2Rt6bv7uxv+vS+eGARhj8Nfw+Qj
zoUhfLqypkjr8dkt/bgXFzrI/CimJeC62efOV8WHvk7UNafwzvaa1odi7+CgkyF/
DP1PZEw1Fhia0PexPnSpO0c+vAmWFhB8ZXbHivcpdj+0E/nB5Y67BHRuTt/LKI2s
GLt3yZ9V6QbrtKFjhpI6m8CaX4NI6dyreqRGtjT8uIFMh0UegueMGIjY8q1Ovi6D
cgCXVTXP12TTUYfMnYhesDTraB8R+1r0U9zXIWd//APp2O3EoV/84PiFx4OzeFvO
m9ZuOu/i1xoGNNdX3IkksiF/EDZAOkzzfwY9hi7aouBIb2+PtbHK538TWULVSOvi
APcjpKZzDA6Wbg6JoLaCCnJu6Sb7Zl4LvcpBX3+GGb1YKphnuAIhtD25WY8kTdXo
JdaiXMWYjuCkJcgNWBoBemS0xQjpz5AyoHZ9H7BXiaD9VuGe4k9RgzXxhpF7Pprq
VsoV2x4HzC+E8QEor7t4YIPXyLR0jdtizPFGEOnexgU6fg/rM913UqYin03uybe5
YURbpdgUPnvlzJtcqPJn/b2T7FZDqaYXmU92RYuGePQyKNvrPEziL4v9fuU7U7I4
gwm5e/QniM9UO0nT/lhtLxA0TuPyTuDsR9ZFy0MFbeGgFzmN/uOlTSQsKS+zioll
Y1N8BNvYzyhMAtb77BKRnGdVcfPU2ABwwOTw5wDbU/EbP3ie3XAjOcVGen1zewbZ
MDgj/PGb3xSULhlkmqKXKZO+qXQw9wlD3Fxw543PvQn2j5mxrLBN50SBUPzJxK6T
pnKvYqPBpm0UG9e9mgV+GOwZJpOGudP+rdS8VbJ+hfS6VvZQoKXLEabGH6RkLXmn
w56s75qnGVuVHGiTvrZuK+mR5ynD9XRyIPMX8lz/wk6Ef+2UlFpetXlvQdhMGK45
JWTj2cFiG1juMbfIohNJI9dnFOPrqNVBwHg2yq7QHDJHt2iAruFiLts2a87CTC8/
Bh4nn1O8YI5Xf4OhaTyHhvHe6HbchYN5StJt9Nxo/X1Ne/ggHtvJdIfPGLyYppzL
ZGZ09xm7R/5o3vBg8+t4xDQqfE/dfr/Rn9RIbU4npmRrS6uPOMjteVlwteTgoZza
co7WuO68sbrhz6cQUlesbhfs8FXpbaka6kf2N8jcG8QVGAJbWbVINg8xwCYNNhB4
jB3Jhul+NnVBSSdSjPPb4OAAtTyHrs1AfAZsiyE23nOvzMmMhva5qA01j+c0UEww
clQIn4c5E9YR8QwQVd8oS8yE5A3Uf6mSJQfJasIC6NPrjQkCFgOyzxOSKGsOFPme
L+p7qPv1LmGh9OnQ8uKeB0vUlbKN9GGgM7pAaWcnVb6GtStmJIHhQSJKfRd+dP49
mCNTSDWjSOg88KWqNIQRUn9kE20rwKeK7F/G59o8Vi31JkR0KrjYrqEqfaYXshgC
CAfG8tdZGhpW1wPZydKmr/Qy9Ln8tvCo619Zry86oc/nHxJe2jF3hqJ5nJJf6lJy
yX6o31V0ASaenwDxf2s9nzXTzFBaRBP2GzwoD06mNqRX4G8LeZ1Cc+JPvP2McMgc
9pxsrdcXbvppHYE1G/jnDtdZlknFQ/gujEGu4P0TsVKNxH9goj80Pez3G96eMbnf
Q/ldpBlDuhOwgIB+ricXX1rRmaBjiQhK8/SAsmHSLuuU91sqjr7yEcaIRfqiRp4i
LQBWm0ndq8/hZeN+odrg892ATZH0dwIOrfuNJbKrszsM8BMvSqev/nHsSo+7O3Uo
qAuSiZIB2RMqC10QhXZEwacwzzcjRIfi77tt+ErbIIR0xzfkSqFHjAgNf2m6DCa3
nGvFxaabIsAQHCMiszTm2Imf3LfvMlJSVWz87acvW5T1LbreSpfMlp+eICiyCvHY
oWuQD3uELIQP76/NA1y78EGVWE1SD8awUoi9QwKyaxBIwtIwQUCRMtGSpIhxPnpU
tN5gmkWk+pDxLpMX1nDo+4fE984k2gfhUbUP0laZThwAIFm0c/srOtYRNVvY/SoL
JSPhqUlqyb3s1QjVsh1B0jliAI1Xh8ryLHyKRu/qdDOyr93JGi52SKAgpsEi6xw+
eT5GfEml7bezdGfZCzL8+ljTnk3LubeeUrtwqdVHWohr0/pVWA1PUtHG20/rsGs2
Uv4M5wZ6gmCvsYoJEbuaz4jFvFjRiQX/hxk1b6pJEWARTJ7aDUFhlp3Y50Pn+DsE
WtU6YEj6Lu1TuO4deWDIyynrH77Zd7ZOykVrgYFF18jI4+vVM9g1nsxqWN8clS6U
26fnSRLx/MZxXQo9mCJD73Y8AAU4iuRmyX7nFaDvdNdWg3aUww7hf0YlBESXzt9v
Q1/JnPNoJSfiGlTgE9gAPteid0oBjG7JdgoSMqPF++AemWFWoO8USJaSwK+repin
Wmpr/cDP3m4O/33kwj9D7iCh7LcVAUfBNnvEEEKMZGYxnEoIyvULjn5atcnvsvxg
ez2TFORE/aQpu50VVAlBLwBYF8jDZY260MQIlhGjcxdovKvLnkfwLFDKnWmLHkHa
XwKeIqbbcIZ+GqAUjG3KODAUVqBtAy7cZFi+89inqhQHruvGf04PVdP9xKqnLiwG
FFNeJsbOtC6Jnk/YRLtv+LjfK8yS962248qp03xyZax1pQJwc2C+A/PgQf/DoT+a
WMzr3xC6+QZchXjHRjlo+GK8bvz1Do73wIYmzCAiYEmGAWRDtUYEqGkQqHjSxwrD
IS4xDa1RV4cmApRtrV2bTHvmad6dg6WqvgzmM1Yj7ycVOEWqOeZoK860qmv4dhOA
4gy6jIxoeZgRXGGJqE+09WrO0iz2AbANcQDuvZgOMFD4Q9EtDY5DVJpiXhC3wBIx
hbqxzCbFlrEtsiHFIZd4HR6Ugy3OH1Auhp7NCHYgbhOWOz7PCN4lqlbCM1wYxFa3
xpZJTrbMlwcI+aUiE4mc35wAzWqlFyM8Ba+UdT9zO0cBUyTR42Bvkauc33xtpPxB
ksrtkbY6OX3WJOPjN2th5gP4RDNe/CicSzf9QmL8W/oK9ioo8kIiP/9rr6NsIDqE
Bz/Hqn4k3XrEDp0XGlKjLCShIbS29JnNsBCRH2GsDGiZE7QN+yYAOnmNNyOwMNV9
CLAZGWgqZd8n+BqsBssUYANonmGJGi9HyywFIwHSl1cmc43QR+UXwk4FR319SBNh
XSuvD3cIjWQ8oZ+zaeVPS2+oPIg1+wVl8gLOJrl/pZNWUuweFVXgBfRij0M0FYed
iTvJKhqDqBMFWVMs6DeunS5gLnum9e5G6fM7aFefr8kElxGOnqryv3wAKVo6tV/U
e0W81tRYE98/z6xzpevUzYblKZmopD7EVh9n2LlNcR+A0SttzseXiGYMglehPYfl
Anj6M1Fbs1lGPvP0dHJT9K0yrOldk4svSJfLE547HJ1BFcLgzrXknrF0rMuOLdYu
ukAWjBVWOHEU1N6MUQcsEHlaxcao5anlN2RMJW07DFZ8EjpEnSQ5pPIPVB4aO2qh
glHcSwtBmD7Lgwc5prcSvwOmHp9ecv/NcEDcrgpu6MCGYRtTR52HQIrNcbvAdipe
rs9G7Acv4hP4cXufNSM30iHgg+XyeMgIZUAl+Yv4wq2I62T6q6D0xIdr9JqgG4oR
hoT0D9PZvOCSgCTE03T6riYlcmIFRJjtEezp77l3i5PoS5IbJK+mgtuExeayI0Dw
s7Xe71CkPuhC4kpsndY4b3cRbVmR0ITBt3KUHyqH2h9m2kvGSVdAgwAOtrBleVuO
AiChAz6pj6tGc9Mh9iu9P7lCqQDgN9mhgoFOYLt1cqTf6h9iIoZ+E0b4KWYiPUV5
JrFBj7MRQqUnL1iPdV5cRSFgg+rHUbn9N7MEbkFDHyfQSTyFKp3NoUbyN/XadWz3
QpyTvQHQKotsWh2y+txxaBp8bh5SZiOS2d/ZO4zQUVelvVf3LDDzDkOYyNVSFaUC
Z8udzCidhmD0g47h6Xt4rDyTvQmw5LHFTiltPvQvVrk7rWlEUDD4Wj2NUkI6Dz2u
XQPCM3Vg/vPKowd3OYPMuWbpyyF8fMY5MjdBvFi9vmWKZzt7i1uHjwmEWnIGmKUF
W7uaAL5oWt9wtK/Z6XCoHoq/W3F8c0663wwoFJvN8/Li9lkuHGvbINWsryRvXINY
7s/vsqmsp63tiYPSdMHRXbwCn2CrfPChRyueFd2oRrBzTCv7t40CLQ9bYbxHyQsh
+pi4EyauO+sIjkcRvItHraR3li2H7FfLKphXdMyMqgGmGEh9hGrx998or9vILm//
Q2AhFe1ENnWbKPsKGhAQk3OHDn468Fl66XufWYF6/Q7m1o+gCaUoCsZjnDAV81ix
wQebHIJwIaol90f+9D6PNHN2EicYJoOBbPEVTXzCJuQBeuFomu0ka3U6pveiNFP1
P5Qx0I1hyxMVKOXU/jUXtiBSBDsAQDmy8xIDHC4F6SzllliQL2tUM/8aMfC23cNQ
lCpObLQRqQb14jXzy3OTztEVUT6voLlj676gvlNxv/2SsXN7jV52A9QznkCjgiP+
HI/GYMtQ8YteD5OzdAZruIpAq2BwZJ+cuxZc536KG7WFaScSpkB4sTWDQzkksSHs
pJ3HpGaCb6xJkpI4HikNbHGig/fGUHFLXuNpDAo0frhbVvdHMC+O/nG1Ri9mzBcC
rzd28itdqUs/FX+SkcMn+skwgPdYY5NhrDi0W9rHHbJLxoGLA6OUJS19a2UCzAIq
bnT8XlVikAgT1R1Fi7Z6N6jaGnEY4Mw+L4WBRukviPZ0aKQS3FIHUAGXtmrSugor
VrfZVlaz6E4M+zorAahthtuhsYt6bfWSGZ8XzOGp1NdpTtUiF8rlvuTzFxEnq/GT
UZClnMV8ro8n/esfWYVrBOwp7vETZwV9Ddoc7Emgusn0ImL6tsVrvQqxeaxp9fLa
9ltShpM1BGEL5GYinDTtJrRBnq8B1XRVdgbK71jEQkB2MQbL+kw34QSeK0SYzgsy
xBFFRKxn5PyyNatmNTI+SfNMyKHZ1Ebs6Ggse0VlKmbJT/dQp4qZTsqvSeqzla+o
2KsP0wsv7g4KAAPXlBbljPyIgagodK9ozdX10u4BddnobQeqoMRjzt6POuo3cfBG
T4LNbPpOJ25QYRBz+V859swMNnsmH2ZHh+5QAa53yr+ZbOekoHOjaIt4QEwG7alf
v82i6TTlUnjhsVoTbFuJOmonOlm/H9+i/bgtAmh6OH8Ckgjo9TLXQxXaRi9g4iKq
Jaih9BEKcOvJBWHyVJzJtIvygG90A/ZKjjp9L/xsuv+HcYNJJtMZYEK5WuQmwtWM
KPBcTUkB8VmL6o6B22ANJPuA3pgmIvXEhcQ6UUDGuXzFZZGp4pjGzhpOTFlZfiHx
44HUwawOMRoRr7DF//G55jaWsfQ9UflUZqzAVutECvVDUejDxBU2YywyvmqBZcEQ
Uk0T7mqbNS0W8EqQ2QDyoW4xDZ01I3KChz4rmN66hgljyeuvnJdGGNOZ0d3P8l1p
c0hlzFlV9NWPYNUnCOad67UtyX+OxhESklATKDtN/wOj+AteZkH35BaA5uFpDKdc
Ia9AQSM2RBqkUg9A9yXvKZz2YIFthsotTJFpe8EqKCilPixTKCLduJhBt5BDOwOH
VMUMhH5TQwy0MIw4iPiu5nsZsAiMkyPJcJu7kQC/dsGL02Zld6FwPyoE9Xq6T/I+
yxI0tn8Ce1aHUo+cp2ZuFxYvSvWSbDKWGMVOHM2iDG4J2yKklq7Wnshh026UZkI9
cqU88gYve6qm1sFSGtGM8toxYbPYkIV6sVhx+NnnXkNmVChUKMjOUG80FlFXkXa1
j6pWytxoa0IdRuty6nXYL8Edi2+3eIFULYhblTn2RYQFUpEfJSgxA+go0HXuV0Hw
SPPwq4Sr7wwWpbpjOu0SiXKxLrMmgEJJ7AceYx9K8w3e3YcN924B+bOuaO2vKvNW
Qk4m/MlKwnNLlKrG7WJXp/kzQsADItp8JvwumKfgvLFUn+GD8wHM+FfL17cGlUzJ
m4NN8AA+yPTsnPWW2D23X3xGoo9nlD9lRGzHw8k1xvnL2i9kgH3xPYebaS4U2Ro+
KwTFVo7P2DLJP+lSy4yFYM0dYz3ddW93AUuRa+m6UB9UQR37jDmiZPIyjTEh311u
s5T/h/927HbnXixbM/EcwsbiCiQ8IPCWXvN4fH6aZF1sPL7PMCKstMgfjmOH9NkT
knI0hHHeRo7y8++5bWikpkVvKdugwG9MFDvN0jagWQ8bL/5t8m2dEPSclSec01NX
CxVWfWIKIYG7jLNNP6WDIm2IoG/3qPUgtPYK6e11reFByZFSbasVLRKLWLiW9oQ/
5yp9KfY1vhBl1JFKdNhOs5KtAMRgLEErUMrlThcuaa6aRBqVA5rReM+khfu0Hie5
gtTqIZmF+K6XUePu78Al6jKTJyjrkBWGVDPri58IIs2vPjQqO2+3AsLzxOKQox6r
FFcgp3fNXX+vt9SZTqJT7ruIx2ZodaWaBiOavdnvpiR58M2pAms94ZrX37v91hqa
RdIFBgaDppNVvE6pFUZvpcYnVLzCFCUWhJuXsB7PbOAbIc/1CGpFuZRvAVibC/dh
TMiyCXbvcXCXyHM5HHRqliYUylWs0qsBpB0iYzIC3koONn6Kvg2gbAs3WrDLgezU
HCJp2I7BI6xCBdPRDiKoaYAW/NOCuQNFLGo7+lVYFGaZkYKU/KL/O6OyLRy+lmBW
pMF/E1SZI2J1Q/LFwv0d8ILZV0Nj2wfTlLiMh/M4km1nUa9IFFC6cFknCEUobg6n
ZgcuEap63lVPKTyHjhULyDltUMcrpAN3o3HnXZWGzUnZ8K3Rc6DZRDu8Xr+pDuNF
8jBFXH4Yr4OlBFbWeT+UTqHmPSo9SxSqxqN83daIXFPLa8hyfhRETxAYrK/0iXxb
V0OWRN+MPsHT+bnTp2+ARPxcAWLudYgOwuS/I8Z+gHG0SgEXM309rmxoVGMM5QDJ
6TUj1IQkHVc4EdsYKzx55Vb8xBkXlyOO06u/XsmA/22s+v3HyMbFBInpig5WGn4L
nOANyi2f3N1fmWjeDRV8e6segMYLHwRRRIXIvXVE97uva9xx4aWxc8pYD0SZYCg4
lYTdn9qUGO7urW2B0ZsBE2RCVKrBpts1CRLW7DT/Ghwr6lDZ8pXho0A2MTvdtnsC
ClBVGT/s6cs68vkE3rXoo0rHgMd66kPz52GsUXUXi7/VCSg+C10vxPeV3ioeHf/D
xa22XVoQXxB5Wv/QhqSi5roQFZO9D6Qdow1tMSgAcsMmirxZ++g6gYTwSok7RzeA
i8BT/ZkiYvd/rhknF4t6fS3KfCRwFDO1aeNI3Tlu5adtB3w0woI54SwQAmvEMqQY
r194zj6N4RKvnsrJIpjtXAIPBFK3WkTkj5Xot4y5y//3GvL0Mqi9GUYT2TGYYIWN
L46sutg73XWTxO9D/zTIrCmzVRG1MpMAU/G6KRVtn8lbGsXnpgtoF2Y9tb8n2I5B
W1xLzMP2wUuVNbVTdbxrwEjDTsenCKMS+DCBtedGXLgFAoCBd1oIeq1ItgX8rxXN
p26SY+RAONDaciZUcHk1hnJleJ4VYHaFFqmi5yS67+5sfGcpLZ9eEPiq9bsQbapx
luPRZthRIfpvqcmbAz9F6W3vjoKGc7fbdYh1lmn19EqpDtSBz6C1OnbIdyKXEzyw
WQtr7LMKS/xs18bN2ak8RGhCQr8JowXl2LBvOo2u/VJq69voF9mKvb4UXfVGvuLZ
weyRb7OHliz5YN+TPVrGc5N/h/hEpHJsifRDbTb6UibmNLnyyp9tgxlv2A1gxWDi
hH3FqM6CPrkNZOii4G+cwPToyVbBywuQnfbftJunx1NYgWiqRMD0EZ90SFkxJ9tW
kT3aOIX+gz6VvIIkO6pH9JF7CkS06YRrkCuIP0em6xCxzGMOa8bzpoRqchuy+iMH
EUzjJbQCdu4qV+wqfyUw5gOve9uOq0ki4NL1nE32XhrcpoEbpHWi2cUBspx9Gxbx
T49Mv7mMaISEC/7EWo2A+5m5spoxhMWhMvZ2iA3RL5Kf05FtD3dgwC1bLt98lcxi
pXD3vInYa6R73tvsbqsOT6XigxzTEW+FonhI//9d2dhHozfFe9HOWFSADPCmIR02
SVvpvT51zzpgkA2DmAEoSuVIXEeJYPLOm4TlFfrqgNCsQBMLOLLGZF2KyuD1SPt9
Ax2PkCI5OkVU5xOLYPnOzJlaQyz0EYSBd/KvTXLkguQb8dFNvaOFixy6yRSg7EuI
l9vWpi08RaI920WmWc5R4c7HYO2IJoNiuKjPxTD6kpIx1VVzh46uv68No25FQiue
RdxmwgvImtT1LnjqQnrqMzpvQqVaer2PA9OLfZYVUzAF78tGVA9r6dlTaxmkj1cd
eOEQEzt7qd2K09XnHD2tPDZLG4a+Z8U1Z40qoUSebtxCwZ5ZNTgEGT+0eI/tesCl
zBt0EOLkgQDKNAbhiKKHTLzkhil79S0r2n8Al71i/xq9ANGO+2P0ZPECjqLDPKWV
rKqPVFXIk9inUE7YvEkAWO3L1gAC1EQbict6fN89JDuJD58O7fcb4Mzwmxakmb7E
bEK0mno0NeweV+5dQ+sJGKzj0rkAnlhMGO8qIg8LJbse4if4LKZ6cQGdkPajhVHx
jr1J4gxKa//ExFrs5Bb+4FcdXTMV6L0Gvluez9ocZbff05rIEh6FiBeg8T3D7ObA
MuNNKWQmtn7b0rjkWvL75VgiPc/fvgV/La2KNO4U2zIvVzayaLj/UgvK39iYzwYB
6SfwsIgnnkXrhFPjM19VWUs5KtcKFLmNW84QaO0tExazdSKOaPg/ET8WXjEbTa03
VAxY1BEPSC7YKZpsEqI+H0l7SRG2VdeekhZldXhOKmgNdu686t+lF6GPzjXaSOkE
MyN5myRQH1W2cbpjlBcTfuPU3H1oU4TD083UIV4L2rFDy0iHOgO7aWP5eU+fXkCp
nb14WaUxzvl2yWOfK2RgrYILWdYwIresUQJ9FToPRLYEVjQb7F4cWUNr98DdjRCW
SpWxls+Uc+fE5MkpN7067Omudl2xfrxmbXOsWVCHnX7Gtc1Ik21uOxFlIoqorXbv
u7m2nbJkLGgFC1nsYLZiU6QQbcDSZdwOCAwx7hxI24ZDc/3x6ob7WZpNXUfqS5eh
2+6PQjnElf/+ilqpwutToDKUd3G5S5Hrzr0YKJeFcoAOOl5GQEAswDsF8Cdup9lh
Rdo5ZwT8p3zRqwKGIJLEERl5ZVtVMhNkYi7I55H5gOoeEhNynzW1xRJG3j63K41D
chpK5tf+642MQaMiZAX1FQ7aq5H/WueRMO6orjZzZ8evziC3WJ2113K0LxLWqZCs
45DyatBbQaCmei9ehAVR7ToqvIsns/k0l8f3EYMkh8fmHLNWarsEpHhNyPGuBsdI
Y3k+am+E82k3GFBo6s6a9TAxWzx8EtGLtL/nUiUls/zcsByT3L8eh7j2ew0pApKu
aBBfLo7iwO+whnhEN8zo3fxBLofbqLTONDXrkfqIVyOMngq6vAy0e8A2/eHdKNn/
pJRbY0yNAq6MPAoxf7Nk0bdwRXchao7YYeI2YZND5FGOY7DKqKNOHvg7n2hobUP3
weVgL1merz/RDqA944e9IZ6GFzDpBtINjW17TcP6DMt2ITTjEmi9qJE7/ISTPfRU
X07zOzaMlohYrk6wOriolE32/t8Qf45mmW+8EH0OAYJAOzvOmzptu2LbYEuAXtJe
P6TqEEF2SoxG72T4njoT/WDEC2MT1QZQo/uX9RC8P4TmFK5W6hAXWYYtsfy6vOsr
4xsF+NU8+goBbTUYro8uHnljQmBoKWG0L2/Kp78U+TKUVkbw6ozyRSKVDqB06nqS
jmMB6pZadwKVzPvFgqI2Pyiiz9qwO6YpUpBxdEEZpIGxr8aQSgSaVPhF6jsSXhgA
yqxAPt5cyd6scDAnZpKpfsl/MbYWq7I94Yy9VVluUoqZqf3NN2M7YaZwxPCfSrz+
LfeW8eZGk4RsY74LJSvjWULvgjbP+7CHW/rN4na1jBYhuJk7PJyq+OCiWEMiVszk
nSkWWO2iif3oi99EEFolQKsIkTn1SG7b7t2ncrhtmrtTNAF5HBqUEvly8IcfsQMw
Kwrg61ajLsrme0BsHMIJVz6WILYvMZxHbA4ZdJFR6zy5LsM8ke/0pwQOfWHQ+AJL
fx1rqNLIOWYo9GzaSCwJ824Y0VFPWUPDSU12EegZi09LcZOt2fIgpWQIBPXjNxkC
JpKc3zRujqFT3bl5AU9XJtQMQbVMQOUTgmQMAu4upVc7IFwKy91nfGaot/IyyD8I
sPkhF9nMAEcUCzoJq+LYYCoH2KhWh7zMjgzomr1CZKCCkMO0HUmvsCelNIsebUmV
XBIUMIb8bEsS+ZqdP0Af9bnWcRC6Nndu8LwJ4uhyA4jXfigJc+mVr7/MTMXz4Lql
i9qY+Dw/9UCFFr+wZRw4IEMzDqs5WMHAAOdMTAsEO/njjlQIA3jw4/aFZKkdpstT
OFS2pSTFkMUwlH2F1rKo+dqpDfJ2bnFJPF5xJoJ+M79g6VZdcTPPJisuKoRG++Sm
r0Nhc7Lg2vISI9N1UJ/dFVmV8+QfS8oHkyqU+iaMtEpvaCEvs9dyIpktRSYL4ySl
/zIaO7yKYfMHQjEJZl+buDQtQUTr5+dEQ2kh5NWY4hoSCxpFW5kYOar8JUkSLssv
FaDAWvijRHVjeH4EmqtCPTqeAMl27U6gOXdAMpsDpv7qOVqPiKyKB6YYo/X1dxa8
qRxFbQld0Ae3YO/+8TZq/itZ4TG6b/zbEN0RAg/nj/3pFttxQ3yrag8QOVGo2p1a
tbdiT3gXn8zxeHXAaeSkSQm+ZJR3JEbhpiS3PGkI+tr227Hf43U8xx0xmaPOIpeE
yIhQsxP4VMLoPoWdFyLe3yFMP0G++04L9bzg5zNQCrGB93Jmfxc/oTm9d5rnmf0b
g64rjIs72y27XJCgDH7AZp8jP6LcOfZBb8lr06DoUbwznoAYgrkUSlTAUdRuc+w6
A77BmjByRXIx/9TW/0DhWQlZQrqCaF3sz5grfXO+LuSbpOoVUg1weqoFNkgJZySX
dC2p01AZoHtrL44kxl06EeeBvl5xTeoHAxRgQCebl0vx+/r7r2dTbmZFHiKMVSo+
/vrL4Ht2szG7ke8nCYqI+vyyKfhGTwySa96Ajl6QhmsNzyibXJgG53teZoweSCsK
YDRyWvC0phat62kyMVmggxiBMLz/G0S/9BzpJ1Bmo3PQGWsI15HWACJcoYFwTBsK
Blk0cCRxyW7Mn1rvDtKzoLhc+6O7X1blIoBZBo4Z9MJFvIj5R22w7kTcv+1nWJKd
TEj+Na5iM8ne+G6QNPB9X/+ESUJqNQCSo5g9HmGs9VozOISnrlFabDo4Kxi6abdl
q98gwiSlW2iU5K9nz/wy2wZikrzaKhI3JT2HkzzFzZRyW2tbTdtPHgTRe1n8WKfB
xFHHZolqeDDb9ydmBEe/0VDSaGIRoIMqoe3usjHKlt0vc1tMh+KwDn1/K27WSB2k
vIADywsdZyDckc8A5uWGAvA2Y2nSjPfdm3jdc1RcJczBOJ6FznvSaa1I3XZ5iF+8
yyBZcuY8pv/DTCJkexfF6EMkf5ChNpTA/PmizPCBf6tSTXpE1+7z00uaoJqx2W+U
3jOWGVMGlH7ffV9TArnoDsY2Os4lStit36SrlPysceMYgxTA30JG+OCTNzAIP0KM
8h655POiJgUIF2Y/o0755jZp1u2kQo7//+b9JDB7gBExDMbL/8SxLO8gqO07hq1N
C4PECYKv0J+9tLGsv1M/R73Kdd8GZIz3srCF0vGOATVV4XNnQMJf2/rU5cSEEpcF
UlWDMrPplu4I4tLqWEyFov6r5QtgnkoBNZwA/ivkT+/Gu/CVnM68Slz6O6R1Ftol
Br5AixJ3NKq7+bjXEWp5l74Sh4sK3Z+lObSjk8YFLItUWVc/fOQyD1claaESgbHS
gaHC/I1aWU2joM5Y82vaFDwG/a8DPDfQT6fbg2CHC/5hUIOb+cONn3KhByNQC9mA
hoiZ+d982mOdkuERfx7w5NCo+DXCBoymx5GCCS227tmcqJ3lB0m94SWKnAxLNWcv
KRYv6sTivgi+xPEuOji/MZojPh/Cq3+Zw19WVdjs/T7SqYnxB5sOhYvrtQ0AsXtS
cfGF1a3nlMZFXxmotEu/zQnFswULbpnAHtkYg32m7HOoWyffgec8Z99FeO7BH24J
TJjuqtCApB/tucn7+IfTqk2ohgefibJ+FDrIANPNM7Je7fqMNRrdaVW3U0UZvgMz
79C1dys8wd8NcyUNNuOwEqgRUT3fRTK+xYdmkGtUgDDe6kLRy0A4IP4BAKXBu0xh
pqggq0rY9j18i4tOZA5ZnWQjiyGJg2hec5GrlYFYlhOMcBSkXomEkhRhywVHE5P7
VIF7J/zhA2c/tRrnK+0kOwLQA2Cry7qF4VvXA7AyHvlz2ArTPULhZAe4y3fyJSSH
yWK9gZRO5gLoylW/9+bz2VAIYLvkSKpBHZdsbcjZMwTy5l7WIXImjx5utK0E7rXW
QeqD9ZZ+CjSBcmmUmak6GFW6dOw69EXeSxlE4mJh3xuStYBEY0JwNlcvNxCr5GYq
CVEJ8shOsClE40tA1eHl1RtR0SNFrS2/UiL3jBgqaiAij8B009HeExsTzamJyCdB
DmFyyBR3LuQnF+/CZ6zhfQG4xIFjdR4wugoSqD6Y79CF1Dhtj5u+fuBhvWhs38R4
lZRYxuVIyNtIr5A8qMHp7mBjQh5/PPG8es1wwrueOJQk5nmKN5Kf0eMkdps75wak
MZSK8d+qPbvMrl76cekDQMbn4dx1HLreo8F6/lkAbOcc++s+Zhav8j5XnNOSRV9f
A/iAZV2k4XieAuips7Axcj4J0ORJ23xz4N1Jwc08GuIv0oDOocoMtHreWHneYQsS
jJiXurINZOzSUCRPYrVPoJk5pNrwVPYfS1NPfDKdtk8WXzSoZ/xzGSHNBv+VkUWp
xVky8OS4PIZbTBkfpWIDhC/DGepuXJS6g6dI1Tneqcjd39DteDZ9oCin3nUQSZ1O
QxfZe+n5BoDB0Gv6Mz4iJ16IDNDu+FowtlF3AYrVzAiR82NJZTkAgjIY4+O6RlW4
f0ZjIuSeVCd+jzcZQwFCk2lQw5zMRML/5abxh4/VRTQOhMVxg/egrgHdVKAWOjJw
nnLjm3vn09tMLVK8CwFOXnQoQyCLeACksgNzVVcy9M9yULltHTktVgT3LefMFmtD
/9b9B7p5Jf8vtRKEtP2syWEVh7hpFVx+eYgdPnv2EzG9sD+2H3yEsXqClXB81kG0
5t/iIlp0nIZXmK5zNkttHSiP82nwaw9Decstw937TYT2GU+0RcGXDBat0yi6lYiW
lvwMoDOIJ24J9LWaiDTETf3HKZ7J5VwCzhyk5BL3kkHX5hSMI+GAX6yogAmQ8yHX
5qNOdFb1jp3EATMI5EbCTJPO5uWJ+H6RdbFmgvdVItBDppEvqZaaPAs48S6jA26h
iNe3xWncn/IprhLoZYvTb/FUHqrkQH5EKJzwNeE8NWe8zqlq09IiwfwhkOC3bM4V
1tzzgchvtlLaHYPezof6Pmpy5RgPfSjMUZQF2rMD4kshxadbc9iy6loPtCmZtIPS
J5LuvXL1cz2CGUmDDnFQ1YNCFH/WGGvB9asLgLX7NKNAdCDDUHkWPthMTH1Y8Rog
/9WUtnFa3hfLJoSJ7g8kZeWCv5PsuyOc0bV8ZoFM1PbxYQGV2WZDiIJ4U1xTp7jW
3r0gqwhvbTQxuH+OJbazYs017tgVVaIoecH4eTNEpI/uDxkcoxVXcI0pbRv4Jflz
oBvZ+cv/Vfe4naUXaRPDknKcBky4P5mD2N3/SK61X2hvlRRDfvcpG7xNV8h7iQLh
WDCRLb2oPFDApkx3MRmDURILKxR9eUEoLumnXEIp7BrZJP60mVw1UF/cqHrj7w9X
0Ov782cEMZCobTQEnG2PELGA/x/+ktk65bEClUqhvNnpziHyRTxvJiUGrs3KRViV
T07PtVNZt+FwV7Y+Rx7ZD7raE50/K2SY6pJ/9Hr44yQhwBzQL6uFSRGWhibVdtOJ
CBHo2RKjUMAiyjOA9fAxJ0AovEEQhFEjFUQvrcGd6Mpr1AGsTW2LxvU70Rd0Whp3
t94hka9jAx0NAHEei0tPbXU1zWYdu93L5fx3GzRFY6nIYnnnOpTa1qbuGVWjIkBZ
lvgkhNqzrFzfv1qxKPdG5wljXhBn5jTr8ty+EuyqjYPHVx9N5RZL7fmK7dmNdXOo
w8NX4HO3/uTpUM2f+ID6hi3Vl/ZeQeEc2aEGjvluVKXDHXCQ/0R+Lu3AZtT8akY6
YxHb6vhxgwZbHsaaZqk5yv+qCIJedm7nSYDN1ojmziT9v5Hj562S1//im+p+lezJ
mCkTzKpPqcslPI7qxnACn55RSVVq/ffbgl7r06MW9Y7eJGMCS2QJU+5KvkBAov8p
G0M5D8adcy9wUEoePsi6nUTTYFkHjHaE8oczHMUoHXxy+CxzKfupoGU6N64uPFYi
nH6fNDQ7jscT1lGwdHG/TULqU0gZtTdAJWRAvihOVD+KLYaF7X1OA/j9H8IRILXi
lioXbdFh8ZcYsi45Kwx6yTo2821B7LlpQPW8LY2OUhOwdMXb16z0dr5skNPB3/r2
NLr3dxDoCv123WJz1paVZCnjmJLMsfT7YePukVVZLe55751sSs94odCQf+6vaDHz
pOt1Hsl5QEoXwSOw9TEJUxDg57G1iIX6RAfr5Y0zFY9Wt5lJvTjoBC4Qn3N7AIsC
wPPSnlXiHSEGtcesJ7HW8YoJcJnourMX5zqEUgHR1PTwo2EzcWuMq1QhNSyuOl+M
Gz17Jd5p8BW+RuSxQHfn21hY1tSiOi2hq4nH/rgOO/gpXgZ8AMQSB2CUztjVblUc
oqpC22W68s0o/TFA4PIVUcGTrlWGAvhWYl1f7SaxzdQ1lwfzYNvYDBm2inHluyE/
ziP8Vtcs60tStQovx9VaFqmasHt1B0zVI7NeWKxJ16PAaQoZEmfNI8Jubzd5SCsZ
uQxWG0YRaCjQ+UifsnkI2hBvsdzPj4mcwj6NA683De7MaU3hWA8HLNc0zYhzmRJQ
PT7B62lXHDplQ736jqjb3lDENmU86kUGlHCVfMrkdMGaePx+RR4sDN4YE/B41Mym
SzcP67a1Z7Bj80xTSsdkRdMJYXuNAJCT50iwXdRhrNDyivZnBACv+TjIepVFiCtJ
9Nz2Or62RG7sQIZF7gP6ppWR5pJCNxAdybaTOwEThFd+uxJT60xDQrpvt+q5QfAy
NG1QLbkq4LEGi7772iqZTkEeVX9AmuZDUCEs5fOKnphPVkrAwDtwjIA88ONbvQ6j
c9YOsD1Qdd04vKJis/RtfBlqY2/HEyhqG9A6ADNOUyeJNPkFQVMSRwQDrP0ACsX/
u/pvV5znXMFvHtX2lK9+S6C7K/gWaRhlD+N9UOeUcGGjlvZ3mAxroo5xcD1krMOs
P3g6kgT3iaHURhJ81o4agSop03EOPaKRCAB2Xq5LyucK5O+nzumZTVNuPUg2Y4zv
pNf1NR7GThQeFz6oH/sXg8xPQzyYj9SWp1zEAO9lZGSox920n2JlS/nnatuBLBIC
9EVPuoirOPCG3RlL2mCvdK/+kV07QoaVoML2mCjf0IE/Z2BIxVLJMmuGS7kdE+rk
rUA7gdzpANZsNm/gwbcOA6hL53x235JvFm0E9x19CXu0Kg6vQ2Q4f2yoBa2+XSSM
q9tnK0idpH2C6UjQqKNUMxv5OGNgtkSvqi8w5jhjBM/XWaLR0xDcsXROgNPH0CHk
Eyrmq4zmlbtaJW7MGPfHk3OHCsSqIUANp2JZFOmZvNSJVLjB1RmHr6tSNRR5ksWK
rgI2SHrqUplnisYpVs7z0Quf+lKBTFVHyds/lXzrW3cRDf8yZKrlHGJOU5hMdFQV
JDNEHpIoxfjFmiks1BcwyRvZv6koBWXXHERRmktAju1YjmuHojYelzXCRgYCkRpV
3tkRx5e565II0FCGHyllrudKvVbG+2gZ+mx4GQrXWkC4rKCq/MmHjwOA5p9WlWEK
+R/Jpo+YyaD7Dvy0l5rMNqHGhpGI3rhNznJSOQAByMxpC6Rx1LkVrpaRVi2UQU7J
mIvF0QJz1up9hs6whs9z3v571PIcrhTUJpuhLnSKBVpxZ3sC5QlVnfdlcP8J2LXA
fOb3+OM0/57UW+UABL72HDU8HXDRAYNbUJAIdbscATDYblu0mWZbXFRQo+OwMMKd
3JEW+8cp2aGNjwuBgxyMBT5ZwRagqxYAFyA/u8Jlcy2rBcNtyuIhs4eVpF+1XCGI
65KGES3NvK36wtzJ+dfKxsl8AqaloqIGSZr/f/joNTQUwxFA896fSZp1WDQ6ni3Q
3uL3zouyQzkJYuf3BCWktnVCQsZZ/Wnyr4oYAb+ZKdTWxl1HjDG54sJ5ZFUCaUmN
DqWTHOmRACfgOOJRxbsT64T9CKR1jx0IFBRHe2MAPkb82JXg22vkveG4Wxk2b4Wv
O5C7lomvzR1Po6WVhDUjXd9ZyfzP272vAV7qWlXK129fVD/cKhN/UeFFQtMOYFmh
VoO/bxDgU+i9723BdVcEkiOtYv61MTaQ7Rj4wjFVTDktNNn/xXxN/BH+LPPeFKbm
r7SslJuuBfBXfON1spFvtX/7phHAWrus1iSQxiw8vOZp0vEePxrdaFnzxdgyQqL/
2vCE1eF/h2iWRUPkRei10nKsonoAOvEZbnrsJezQSz/E427oU6+7mAQGBRWhY7F6
i/SGtkJztGz8PIUAThwPYfwshFQ3V4W8sC7xSR+UPbPd0Hd6WjE7Kfbx/qWls+WQ
KzoANeyWmItlNhmWSSw/Y9AKyxf51h8KXsKz75PaxXzt94OSSalH76L0Q7vNw3Q3
vueslOVoPMiyLl94x7x/U59H2lZ7oHhuIHn0Es7VrlcbbuT+CMz8QKc8iIjcrHfV
Gp0hWVzV+sbtXWTTNUJZ+Ow26G0HlkY8GUsri0S4Q3SKQLo82y3A8dPSY2VWbmQ9
X+2fkewdAvghBYNj2oPhYzB1RJd+0waBj1Or/P6ApaB6wTi1Lo4dbHhoiB0Wk0bM
Ew/Y9bejcRREjz87yd8G/DJM+kfYWNf1+u1VbytL54UKaKOnjlRRcbLLUEYbblHY
JRA7rsNQjIZq6xUrkcDmKgcRsfVJpF+sj05y4cYgQZsgzdcSzMra2UINYzZSTGPS
jzjE4HsevvEdiP5bES8l2VEV/ua8hmD9AJMSv9Qz79BQmSZEWQzRkfvbjEQ5S/3z
4oUxZi2POR9vWyDriSt7kgbB4jND3KedIN8kxViWsmmfx+NQqPjLFFZKqwcaEYFV
H+jGDNOv8Z7Un+DajHh7r5/pYtNTHQJIYguoKGyKKIo1tke1HXjO6MmHTSeTvD/a
+b3593OPUR03yFab1zapU7VnQj89nOS49y8n0Yfrkq9lJecTBh0FxsAwYBk5b1xV
Wwt6gq93mG1dYQ0emcF6tOU89LNOqXY/fddXBdiWaNDsuefVnsYkpZnpNYbW1ULa
NFyxtiBiGi4k56Vl753dHkm3e1bixj9JfciE/5aN2fcQ0ijoxguXwKpqk3sjE4hU
QJVE5ngtopsw8lFruMYLxqWhFfIMaVZWKhDjMuh8G9QBmlCnJxngiP1MKthNJuGv
+ASLKLf4JK42dMxQxmx69j+tV0zwp/ziv7F1imco6oADxS4hD8J3FQdSXr05rM3g
R44aoGeO+EGJkC+iNUctjUk0Rdina93O2Rc8uO0jkELrUzSX6My6msrwK552nYkP
rk4oGVrS/1wggRPN4CV4fGYPynyJcnkcF5iQbwHrBi5jZCQmkXUIqG/cxXYFHitu
oUsNQo081IV0vx3nMbc/jPNIqinkJ2Tetji7OodG4LRC6gjMcF/Lm6eEkd1n/0RQ
3s3dTP74B6JPhVVgDNiIR7VlVFuungJDz2iCF8R7eP3Ag0t48T6JM/pv7EbxTcO2
OdLW4hSfXBUcnWg8jHy90b8H0HMKjvLd1TEPFkPdWXIj7PUwcyG1seLxAMMsxqSp
GVkcxM/oV3QwHMtn04nndvUn0oO709bKf5HGjmtoxjSZTm0FM3FSfeF/yqKjIwTG
uPbgC4i3zMzy8aLTFO67qV2f6YWlKf8S+8rY0/BWFsFCgIUTdT00/LUi4WxorqkS
fc5pFJE0JogES9qC0YzU6uaSY9lAmhHdISSWBBAQNfLcva0u47RHQZBVg3OcbEh0
LLcZ74MsJ/D2LEo8WmKvl9HfwgO1DhQCiQ/uRXCuWTLbWTS8rY4Jzsakfypc/WoW
tL9Tbcc02YoZ5wow3C4UANDwYZj00ew/cRG4J4pTfeDLheFTvaPzINCtiwXnNq6z
CkQZgP8ZtdDvKBrSewJtuVKsM9/y5L+UvSYEhwmCg3xlmoRRulO+oq/ULcEeRvpX
EkmgGfbkXP+Yq2USERKL8vj/EkbGgl+ajbldAi8vTj08JYpm1pVfkHq3F0KVwp/X
pLTY3tD4laZeG2jiiUxOGBa1jtEtq+gjjAmLUNthe/JkK/VAzz+thQ5W7gxvWv5R
eBsyhmSwIDdc3fD2d7R5iEQO+w9gNWCJIO8DjQBZdJ4Eb60RRr6pBiYenMK981Ek
K5UOnonj0wFgnpph3BNxcRkUIsLxIEyRpkBPgXG33dSWufU5D1EOKwny8MmrdYo1
WXMdSOVFQ4n9REwzoXtjG9JcWDTnvnL1ImEzHDgWUiBPB3UNyxcWXPPqhesXVIgh
yQQZQWYsX6ZCtR6XB6m9OWePWh0Bvuyg5ZLGdyjbwXd0LA09PXIvgzQJ0HrCITWA
3zm0pEt4OrmlipZdMB4idImwh8FV/KYqQDicWEuA0AGWppNdpQFHyOzqVGL4vAKx
OFpRBbPhGaaa8fxFbnN8F3/v2BZrkQA6fe4m4ip+t+IWGsbfqm8wDEXQuxbRvPft
cZZUIgcJr+E2v6bRjekWLCpuP2Tl+5l1r5Fcg3Hn1F4AMihX+QoxzRuNqdnb5+ns
zAULpxaZbPWIgOg3GZoYwAfPIg2Wxr/ntD60/Vdte8eeo/JqUc1Q/OVptpaYKjIc
y8T8e1yPCgvqo4UMe6aAtIDG9GAdt4tzLq9zibog7Gwu57z16cn8qr3YzuMCStFP
FUIOep/P50PFfzbJjMj0nG/ctRa10OBvWwsBbOkPLDavhHwZvlP15GYZWnh+wjj3
ZokYaTmzPdBzuAQL5qB0Edf177Y4DTpafe4FwZ/DsXXpjX70o90uYZ721phHBt+0
H9GgbX8+lr4HB0Y0fcz1yzQp9btF2bB9gbWag4UHeBr5C5RAPkVf4L+GTchDUB1r
MM+dm6RvtNvjlnbNyrD6D8fC9axCvSmaaiA+/EEY3SVyz43hkA9j4K6kq7NpxFK8
4hwXNBI1V/+psGuV5GoAz3zeYVJa4wto67U8jGPfxhwXM9aFW+RKKyH9V70QVET6
73Xl4ETgK7MUVxcvv2eqeyPNSddbb1sI65CNFxXyT2fwLbzUCuHJuOUKUV2bezhh
jbalZN4Ryg6AsuYStnGBhhzGbewkbWPKCUub7aOm5x7ki/I2NemRJkdBPdF96dhB
g+GDzRCpjS+L5ZzEjAhe49C/DAzoEt9cUE2BU6xfQN5V1hJHHWBfLvq+a2rTDufL
Lmf+8eXpYwoeHQpn9r1EkD9nhs+qDeA26fMZAR+Crgx66pfsCRTVb4sLq82XWNcU
I/XDWOGBvTpIAmY3Uu+boFJOk2ZpCT/uUaEfUWYHdRMVaO9cseHg89igrHVFtqS7
owjdOVT1ZzcGeW0HHy1CAqg8uE2Plcv+G+VzHfaAzMTDK+7N2TzcPDs01uv/yeRR
CaGetWIY0XI75f63duxeQtU/3wX5ii/RiVCSaeE2xCir9MC8dLrhvW+u8onStOIx
WmuG0k4YirD8ZeuKrpJUHw2Qn8yScUmFhwr5b5OB9bzZWz3Fid0sNe2oVkWElPla
J5fEidizVjb/cwgn7YJAZihT2XNjjkC/TvJghjUhRvIY7ZpdaaJa1wU2/nkNqIsb
/0U14BmQP6H3BOj3OIiu0/syinAz/uPGJJHQA2qPydO7UzS1VSR4gfpqBSh5VgDA
AFHJEkYu28O4yrsGrbDpbXHFnf2Suvil2iI6q6nf8dxMi1HeEOXkoZfmbqiwJDj1
Xchr0jLwQjhBaC2qVomKFGwOrtyLwn/yrS7VrmQ7Ae4PLNL1Xxe8hHV6PAYUIi+K
Y/exnUQMuCmByUJ0HalZXSZ39IxZp6dOvPaqu8DRxyGkoJBT04LW0zMacdUK2gEz
g0buC6XSNPCaTs7V67uWl4pFq2v767H5wismwxJvT5f12WHiHFXW0zSprKa0oFYF
TBhQ4LOVlCVpgoCjPIQxSgZs5uRpzLEAwdlxNazN1Lu4JMxIG5RTqGPBr3AV2eq/
j/sZe0/OupCE0wtH/KqYFaeZGe2/gBonpcd6u3rQvk6JK7fCDyACla2MTqZtJwmv
RIw6g7blaUDw490XkpLKLT8xnWl4iLT+UmNM3ReZpQp0xYoLIh4Cs+SSOCFviCup
8VYqN05w7Uez5cIaVrjDHQEVAEeyPTunAMw2ys136o6LhC6PaMTLRVd+QW0aozio
bNGv82TY5NLTgqzZ4ZZu+8q5HClDia19I6xD4JF6vdgMZYtcc9sxBsXHK7h4z1YU
poBYhMmUoJJkQSNp6rGt6YbMrp3vISY/HaSH/9gdu/hgrx9r0NSV6ToKQuaGGcip
OGuwJJr69/bX1OU+a/ym0f7nIdl6R6gk5BLNuMoaTaTGoZpe8pEMjTgW0Jdb5pUG
d4e5AdRa0no/bwAZ7XM4qzVWTB1wnUtBQ3AIIlhSDGSpZCBTnROlAGUzebBYHh+e
jnkP4PnPE532dTrYU6ZDwGQweHbEI+BVG1oZu2ryZz0ihxwgu5fFWSWspwLAhIqk
r1MZhW1oFo3K+m9uDAQtRQ5Kk+jM9pdZ4iKAFlTqKWKk+/ttEjglbJS4drZwZdpN
ERZZdacVcudnmSfo7jxzBT8E7LO3KA4b0ozl+CPTGFdIONOeCm68KYzUuWikee3E
Nu8aa5jHugWrAo7ZC+IYk4UQvKGFFOFyucM7qJGsCOut2lh+mQ/u354hLe9v0gr1
HXt8d1AlRWy1ObnJhHETQGRJL6jpkB7+2kvpWEGhoGIESUkug6kdHuxaAJJkpZ4R
Jh27nfnXExYIX7UawSbS/X9WTUDRY8tjUJH2oxDw1R1H+QIkNqwZH75SVS1kvL+v
NYoJS45/hsX2O9ROYbsY67d8fGLKwb9Zagexgr4YQVoUaFPDN6A0T+3/Y4a2yODO
sOuz2b/qTV2b0TseVlmw3pDZOzlMBsXqYCm4FEABv8JETDlF3XzL9T5RCVipS64q
P4WFYgNwwD+j795cIrJThc8mpaZhJS93cg1purE3q5jFx9AxAbR5fa4rXPMSZKEt
Hj2zWou5Ht//tXjANgOZJODX+URO76H8DX5tpcdtYMuC/bxt0GwAd2WtLSXxy9Lq
z7qiEaFt1Zhk0Mmdikhxaliy+StVb87UHO+9Ufhz9blE6u+4tZ08yKVWTGPhpu/y
WAFrJsh36z3pz9nNaKbjAIQxvTdjHVKpkBfDVfY7vocLRqivJ5KW/Pd+ZkgTxVnc
Gce8paRnTLrMsxxg6l3/QHbDNTZ3Rjo0VhxmM1p5AJIIjdsaoZeZ/8/mOa1TadQ2
OIWm9rDvBndGd6AIsdSlZTHr3XIHBRQQR2Tj192LhqpfVb1Uzz+V9gZ74e1Stm98
u6on80pE3EHcAlINr2L/idH4Buxu/xp4xIkFI+1LvqzbcGLsdZZSLNo6+xYsPRct
CpDVRKLOkD7xC0a56wHgTDT7RD8FiCKmom26FT70Bs9Xa6CZbqfJ674m1OpkfE27
7wQoMaSEhV3VZSuSgXXfqvCijUClNjIBZg1GIxxii3Trz37lFE67qJ8HaIceEt4F
kzuWC3If/0XAwY+7x7tEjJFEx5EfRR5tBcQaWTQhzWRq3RaRtYG+OLvbZfBxbagS
TwuGSQflmBBsK6eOAdv+7OoJKmgj9DHaH1qSWoWD1/GWqlne2jUk7jOZ3+IXXQFt
OaSKScKorDgbhxo/wRFMqpsll7UZKZZEjrn/exFz3cs67thsCKriUEqJnx6PO+LI
KjW15AN8yNs0PgrLn5L1yhnuoXQpVlvLvBwdaBQNNVEu73518rEcWx9Ep3l8TiDs
Nax4hOfI/QSoFfRqdWplELlZc8M5ShMb4OAyYLYffq5kuxKD0C+VHTkH3F8nSbE0
XQXNPhpshXaOs0II9bkqXUIiVUai8J5Hvvm9wYn8VuxV00fJ/tJE2mLLjvAKlLgF
JMMnOqjqCujX5wYQd+o9LEqtE2x7RTGa4pfD6e2UJGTHq0zK2xOGz39ikCmx/J8u
46lE4+kxJv42g3oi3b2/3JKisBkUW4iXB2zb0KjDp6wKg3WN4M1Nj4PeH7ImCwzO
jDogdMIXN2DwhrorOsNv3ZwvTasmLWlg7ppIDV7XdXFxzijMrgmN7tXcg3Ccqwoc
vxwhOpbgvZxS0DVRmn0s+9qn6p/u66hDzC0FcezoVD79jg3iSXnTDbc1kpXvQbaZ
2U411fMUzqCQwERLZ+cLmPXhztpLvKbMYmTFN3upnMo9+1IBscGAcElJGQJb/NCA
4vo/dRIwhR9r5Mkf1EjDGswtGKThs9pAf26nxjRzk2D90AM1fay105Wxo7df7/DG
Xc+8L0yeNFByak8lqLRTyUqYR9O22f9cMJTUSTZ4qePstIYpzeRH2YGyt+4nmPuo
7t1CSnDdQpZFfUmWG55kDcQNfaxTEzDQMKwRJh5X3RjgMOu4ONM/UuAY9KO6Vkkw
5vSIFBb8ZPCt86HYx3L5iKYtAaHP0yHRMFeGLzoVQj0K/Ry7gE6h+YorqwLFP4Ni
siCybAhCgOLiop/Q68+yyrubihCtuHQdeD4VGhTCJ6PkhBOqf/kremjFPZ8o5t0D
dfHNYHor8cpMnCGuBDJYziwOL3j+VAwSQhH528N82a1mldJvkO55k5gts8zAOHwt
TlXHXgrFYlG6LKVWSwWQ2K0Vx5hFLxpuD+ryW/E2GuT03TS2bP21quO+gJA3DkLa
LEeOMY1Yx8O0axkW+Tvzt2F+MF2pjvxWfeyV1eC/e1jT3KNeYkvwEgTWfJFeCE8B
DiUeLnr85dnuLl5PWx7TuxN7crCn4vCNUYXmEfgiBIQx6DrQ0x6vB2B3XhtCUp+2
TZHJAbFo56ssKYfv5AEzx4mDIJsWToYpwzGR5vbvBoZQmiFfY9SrF9bI3gUEc9V2
QRgwWpxZBN71bDYks13Vgqz2GSl8UAnCqJwjgM13V17sEZZd1oCAwCb4jYOYIIMG
FwcaQOfBoPak/r4VuA3uY0yFq2uBTZLa83WZfWQpjdn37tMSYHM42FrnDEekS7w2
RW6cVQgJPhwwmoSYM9q0XtqpepM4ShZxfZdiVIttYPNgJ4Z6oljDE8m6DLBto5dz
2CVSk6ySA6l/XjfBbjmZyPN608BcQtipr2EzX2i+Qrd22sSyENPVEzEbFfVBqoBZ
5GYk9McddJxjJCeEjTCLUeBEtqU6Nfzb49tponE69WjT/NG1936Yp2qGq4ZtQFL7
DuRr2gxQBtj4LNNF6kNNE4wCn6ZR2P7JjlI6Fm/NH52TJIxDTAT96mv1uwmSTzTu
baFmXDdsM7ZKep11M0d4Zvl6pSi5Ya6Y2O9iXB6k/SxqCEVbEPngdPFMvDO5uXXM
J3OYoRIl7Gp4a+L6MNZV6c3b+NZCwJL07P0KsKSg3uE6Fkkg/aB0HcZTSrXvbIIx
De6UOVae646QVrj2vccW/TtFehDMc3papklfGCicmZyUdWu0rDRQ6QV0kfW/jCUM
OxsJasA44ezs1AGi7HJSKX+Ww3G6atCmASdiN4AkvKDM2VJmX70zQIV6loZAt3s4
2yzs3l2oQnjKdpaUL6DuHIEHn227DDAfS3NpU3ABh3Aqw6D5UnOcOXuIoYSlu/7M
7biNy7QKf40dBIIL3ha6JzeII/Yx5Hi0iR3bqZNHvthGF32gakh1uU1B6cm2ERWS
txzxViDyBaZ5cYrWoQJroA5w8LGuFbYkAGQ8a4SYIPoWZTvdoJThOWZBFUseq7Wv
IN9uRH6CA7OE+n+KsvcqjxfA9FYEnv3Lifrd8pIB+xyZae2LYeowjm1QRZsPNfLs
WVnG4f+kLhub8cIQP8gWKoH8eGMkxBZwsJkJbMIK1e1x0pE/9llDtLi2RvWWpWrw
fGi9Pi0Kd72GIoUDwb4SziN+O4VJaJ2BfCdaYWLiF5sE9hEGiz3yYzu37p9sNkon
Qi2WssV/EBOW6ZwDcfx6uvMDiERh0Z0yyaiR2wSTQONqp7bhqzHiXjhApVKKON6k
0q1Yrbnma8IOFekI5M4C6AGQV4rGA0gA07dgDXYUEnAM1RMvOTQrmCpUv7g9OrPR
YRX0n1P7n0hoEFrtgV5ibKzeI0P9pMDuFY6ajx64sqoWsJiqchDPXGVtoqcFz5LL
VZtAeXV5Wr9KniOX5FMV42eQsAYoKkJ8eAPAYhJj2LYR5UnIN7hduZL40mSWtkt0
XEZNi5klvY774cLyFgg/5Tv3SwnbR/fUpUY3BkrosSSnMpVbnjd5193UuowG+yKX
n/Kl2vIUof1p8dea7/ogQAGVigG9hCi+FmH8nfOXqT3DyKYffdLo+zSymvJ5WXnY
cNFgFs07BszolU/Gf2MwdgepHFGZbNu/BJY+UJRcRsTWb9H3Llqh5V5NgEzOT3bU
AIEL9KzpiBv0OFwDuO3uO4hYinbpmpnXZUlREeqjHg9CbxPARNxrgNr8X25RMCtv
DJ4VttkTrx9p+ae4YnMxmmPiJfDoPSSIns+UTph6CxusKzTni2jLynOcIH1NowIR
bpmNl0MJZeNN/wlaxl1y4sJ39oLwgnrOtw277cCdJeGNNfCu3S8X6ubV0DJiW/u2
G++eMmNfIVGvzWXIJA0M4k4fwJeodYUphjIN8WsAklqXvWhglMAKY2fPFnaR7yl7
RFyZL2h8QcXqJ1fa/CC1LeCQbT3VimvkgGY1Dfnp+zoYRsTFMQSOjOejbdh5HN9V
JWmyqzzO34G6uKFGrpt/R3SMS9vMM0nHtdM/mA4CRMD+MfU0zdRGqoIs1nySuoFT
VAkTia2FpacXuecA/QHKPO41B2m8KwcOnhZDg1SZlGy86jY4KoFa3TUccImQwEFR
O3luEXDLQbhxGD76JW+5CJ521bkM8JavNoB+DICMbHdguNihx9OCxuoHRroRMSKM
JOPrB7IR5TxzyC4KmCxUrxaRHHxyNHzSBvDUuUatV2df9b1h4Jr2Lw8JvKxZ112j
eUT0A/UsKLnLI3ycEdD6uXeo4nV2iqAAmcWEVbaEFLRAPwCO3GMtuNCivjf95oKk
QKAohtj58h5ZtBiw6BhOl+3zu1wRKFSUVsFSoSeJDia3qq03V39MwDVeV1Cr6x6s
IpbH7Gb4ToCw6KIFz7N17KyCELEewcoIayVtMGux8oj90eucobRzFah6TDdcoMnx
mSj4mAXqoIrpM21CjuNc1S/TxzV+8d47o6OF12YeJ3yrbZTMfFUYiFa4QE8yDmtl
GxCnxMLq+GHbl0SdhUL5xnuksKYoM0sTa3va4YV/wVRnat4snUFfobzMrkJd5+/4
t0J/C6AUZiKWB5WVOkMC9ts9fLFjOB+4OyhMpicaEcbVxHqJymSjgVquTROB+WLe
ZWTnxs1XxpvtV3GZxS63sw7LL/FXqc7dzzGyuUFQyeJAfxunRZLBL0YBGJcQU3Hl
4CWAJ8gia+yKjWoyMjaYe2vIi+kj+6x0CPZ4dhs4PNsKdbMG4Irs0BQ6cBWrbWwT
LdtuQAALt22PD+ArSmPtzHC6qr70A6Ob3GOLtkK8t4ywLS459JkgxoT2s0+tQLEh
3BNlSgrIFu/ksUw7R9oiuePmJwQYiDGeH75iql3XyJEqQYlN8AGfOWCme380gVsO
3Bwa163tKrqoM+GFZRop0nlWMCS2mdW18RUmJhifYNM8U0PZVC8JXYvFfGmJ6yAi
LvdSBq0yFyxGc4bK89UP7G3ZVONyTX1ERNQ98LQehG50cUdVJq3XmeQSliCQsFOR
dzOf54G+883LTEGFLEzQwFJfhmgB7lsRBKS8o8MuCL9Ko+5LRp1FkPM1j50MtgfT
3yB+xooinxTW1EgcKE9NNFZ/0X51Y6Tcd5DSJPimbX07J3xPij3EcB4NVZeY+DsT
VL5ogOd/d+wFBFLD95u3SMKYrB6RezZ7VV3n2BcmpCSEtKOGLEvSr4NZo7Zp7SAX
uiw3oHGhMjQEWxMTHbyCiyEaUn3OaxjkPcuQJ1HfSjn1Ft8/ua+D3EpIxtxY1Jah
3ghFBrV+E/dU4sU+AkkycoM9aTFwNl6PPymWqC9+JIAM3328QU6BBotC9c3a2qUX
0u0DPvGm11TD6rbSoSCm2kkEGEH5CoKIDLtOEywaZ52WKpyqvSE7eynfOO9zrLT6
gut75Ka4kb7sCYlZJQy2DFfeMsW/ePl6rH4uLdb96pG9HjqwkUfACfBCJFq/ohq1
tZed3rAcza1OZfH8YuQ0coK/Y+KxuGb9c+AG3L7H6yTd+y1RmnsDFvzXQcfnu7AZ
+Fy9zHxv1sVbyzCvi9dfY5dOiPD6BPkHGAcz4D1M20GJOAcq32Re9zaxcZLq+s4D
4OYh1qB4es02hccW+0IzRvK3HDxNqQolnqVVfrGs7Cj0X5pMHdFOEcXhLutXeipr
OiT3LkljodC0BbMZAW5rwQJKXNJ8NoKZwLgVYxcGn2nO+govOQuNDdurHwdc/vQQ
vuam0hDG8rX7CJKH9tGdKH7QO9HMOII5WAjtwH8OOmsWcS14StI87PBYb3rV39zs
Y4JkdLqed6E6uUK7rtp0sewGPtyPFxXFMTTp5AyMz2NqpQqtma82pwR5hAkwuhcj
/c9PRiFVhMlw2+nOpckZqgJ/Yg4v2jhXvU4ZRSimi3hoNo6ST8OLCE9vP9Syq+uW
loShRW4dPDW4CzERfIRKLFoPoluMSLVQocDbNwu/bxj4ytJL91TT/fWhr8n8kXb6
fLtVnNVITIUOXAHfF13eU8i/6D1yLNqn9KeBAxqgtaXJMHgl5GD04F4z2wvrmpPS
ZDT6wmJ0onCWX+0HLkID2Z5jQ9P/QF8oPQ97E+G2xLaCkqgDbinyh3Gn2LVW+0Q4
CznquOUni+81Ig4RYRLiexnGC0XkQUoC4oN9epwg/QEE0EvAquto+Vvks30CayQz
lKTv06sdUPXnS/h3XQIVHuaVf9uTRglO8bNjfMCT9p7gg5vaaZqvxvYI+Rr5r3nT
OlFvuVAEQZd0ajqsD8K2ll/DiUtwflQSdE3+XLRya+kU02LAw9quhPhNW5TpDPP5
XhSclGDiw7XV4VED4qJodBc0dNIH/gWQm7tk/0fH8t3UMwZFx6OyN86wEIsg1nHF
XVDQuEbZkhj2zY1VM2oF2uKQs1fz9HCkl02mUTCgVKWYfNzluBFgJ+z2wdJ7gMvU
TtFRaPZIxqCgcgTsgfZwEaN02TLX+qPfkZWDIly+dA7gsr3l0r+uG7px3dF4aNbX
/RnCDXOIeM2gewEbG5fgGLzVWIJd8eGcRVjE3h364qSswyIqiHLzSAa//b7QU3E3
V41iolRKxaZJVNP4KdIY0OfHc1os1Ud7dAkYv6fJc4p/m+JKTPwJ8PoMlF5gMwnJ
xnHQ/vLHnnc/DBefBOZBXHez/IrJrAKdzOsl9Y0EXMDFhxejBsaj6G9Da3trRWmQ
95cFuqAgLQAJ8FZN8stDTkyfj4XQMKLLifaiA5VY5SziSWgEKOmeTuY0V0c3dCRZ
rrFdpNlWywbtjKYNE69162gictoiJsVpVBTyKFJENsAe6JwlhAWl9fP1z3oIvGTO
XneCFGyyI1dhuihJlU63Y+FdkY33SVMXJ5GG42f+oSX3/T3ywx2fZ9W9MpIv3giv
nxaRi47ECBpoDgu5s7pTA7GUr2g/8i7GRhG/92gkAkHy3OVa3qXM7qAve5Nmd++m
XH4B/BRuze+f/c7njXgVLFLcqGQr2iDe2FedJmQ0YnjNvoIFgasr/7B6lf4AesFY
H15b3lNHSjU83Pc85rocDrl9UjcpMYtsfU6W3w6cx0nM4C6hkfS4LqKVfaF6YDrv
jvEQbPLzeEOStZG1z1QZaD/1+ryeOPuWBPA4hqog+8aqL7URLLRqg8XcV5/B8jY/
EewQAiplHErxWVobC36D4sF5kLfHneOVwGUPw8zMwcFuf5nQG7qrQMAf7/X4podo
oSIUUC9H87jHesv5spVp4iJmP+SYGIAU5dlxhEeb0rJMI1bdkwc2GOcbV1qXRhwI
Ud7QQeacxy2kaBhUV9DLduPslg4VuqjhmbRO5Pp8iFV9wt89kak+CwRfPz4Dn17T
AqdGfGgz4ydieC4HpekekliT4CpSkDLsyX0RZkPI73n0IIKxABsA5bzdtzltYbRR
nySrurOe1672N8DF7s8WQmPaBbk2XSLtRDmaezv2WNbN2tK9oqpUN72GKw3Xbrap
HLz7Dqu+PoK7ZNhiTK8ve99fJIP4vCJ/vEtKmIgzeoBYAt+D1T8RVhBI6Ht5zjhL
ql/Aq+nr1b0HKCdxGkwPWzJTa2I7VW5B49JFnvNpPMNkoOYpX7pVLN4AHt96/wWG
6CJC9cGDYHyr5eAga5Wjt8RuuyxEpWWuysEDpajb5tWqmoYrnggfd7J8SoVshqzJ
G/yJgBS5gQ9VhjdrEh5oxgD/LAnZJeKIu+fg7xI2MlQSyESM3kJIr38lGjpU4dvw
7RjdgabSGo8uJz2wuwE2ce7WwCyFztgHqFMpHpgtOhn5AhKmD18qiGhLOYmMEEgg
VKvnTb8KCD+wFpdiOADamCmnascdGtLbjeiMjY9A+yeQUCg/RehtXmILkh0FGCT2
dNAqTdGosSgsIdhSafA7NwILr2rmJZftGNudmQskyYyt4hnmTOJXjIXcGWoI+6xW
rNrFi8IvlK0sD4cOhXyU2EsimzB1l81iXIvWkBy5TWBpcW2Hn8sipZO5y+hU/CNU
onpiHaZWHe+1DmsCdHbbVaXqaeyoS5aatzyMh3Pe9l4m+5CMajbCSuo/XhdRrwb/
Gcov37glJ6SMPN1k5RPPApxhUYvpJnFUGqU9tC245+QDjno+0pPa5DwQW+IKzCyZ
YoMYWpyUnR/odhBM25LefkYpn1p2GZpoolhzIqoscXxbaxhiZ/YUZlhtcI1JIhP6
Pf8T/WhZUdbXl+Egq7P3ggYs5UTE6OgZ0qTUkBcexYZ3VwLwVX4xkyFjO4SF2WVe
rbzTf/hTYgeVmjpfQsRNW8LeASDNIPU9LFGZpyxt0xkuUEbOwRuIbtnn37l0nLaN
CIgOrTuFBtOzxiEmx0j9yJBrM8B2ZbtsZABY/fZ6N+Zf+Zn/fwvUDr0c+MX4mQQP
uKBxr3wjDB7HNV7u9aCwoyy64gGG5Jh7oLAZHFEX11Rc89sCT+wPy7rDaEQOVUFu
H72mFeKq5JA9E/s0+NOnmBWF3qoJnar1jGXUba1zLm+GcLrWsWJfEh0Vvyf7wpm/
gRfEth2ayPTH9c3bSYDHJwLBWLq0eZwOo8YH0540OF4guZRjou+yIJwAxazupwVq
0jfXJvIjrJZzxzTHKyoMlFkI0JhZ1uC/0AeemZ4f401ZGLfymbcorvs8I8oUJKPf
zCs11AfSi9+esbwQvV32+cNjMPSPR0fqN1IzZ/lyTrNM4Hx5p9vu3AdTEYQlRBhK
ay4z7Y+4j5SwFQZSpnr8pMWlHF45vrJBxctM01X8M4yOYrJ/1YkzfH+wGmBROwRj
WEQqZysDcQtNMvDdxkYK9RmlixXA2GWRNt8b18TnzMbHVXdvIs0PI+yYwhqZ/Mha
Gw463Ix+XzOJ04ScE4LSPKXUcfEchX+qYZKoC7/Fd9Uy/fD7tMV+uoWG62Mb6xDg
gYozwadWxDxR6YfuEJlOj01uMRzysw8Nxo9fmd2YdM+C/L/kKPxAggmMZeHxVC/L
xy9JHvOHu3SM0sZp6kiwuIH59Dr+qzqBqirJfIjlalO6qjievelOWJBPSibTGQca
2c4rz2ULOebAmCY1BadMDm1jGgvmKGSj3G9UrEs2XoLBgt20Qt0oemop+kZHhMBg
eJtG93iIXw5+7l8PRbMh0r+meSf9GbRJBfqrHW1vJP+EBmTlGaV6ubLvVW6E5VU6
hHRs01bMMV+0EIj1vpF9PioJdk6yb1FfY8Xu0xxxuGiNTu8a5cQk3U79D807wHzz
XTeqbSY0vR/lBgsTrDq6gCmcIABVMm7fYcHZ5Whv1JxMKxZITOj5PIGz6R7lT9NH
+axBCdZD2BxiSt/7Mu5Ehec5n9rh/aFFsCO6DY52eLwCF2CXW9/rWWXrnkQEeESP
NygVGsVYR99yvl1UPGwRi2VNXMnyY51VlBShkj6ymtDvEJpcKl0t4LnN8fWuVa6l
r4z0FUWUUFElM51+10uHgyzOhypfmyE/dZtW2lo7IzLt33V5TRyUH8WJgCUUbr4b
ymk46rxXK5rS9DPM/0atUk0KgNBiXz2ke5noHC67aWoL8KK38WUKkzUh9PFrCHPh
MC3Y7k05zbXZTdsMhbvWUDgJPkwQP1oGWhrWUyc6bhAnHqdRwVLWVmn0zLfPCpiG
4IKiU6s4KVrpR/l8gIGnCVG2XewT7LGbyOQVPfHGLAFsrJrzKZ6v0BHj+FnNzb+s
hznrv4iilM9/enzJHBL+wQ//HwbC9D0lTmY3C3l0pJgfUDvVQ842bn6GWQImJBx1
HVmZnumrWSEySwehWFGLOhEnqw4Xo3FSR37ogQ/Dqupw6s6ENUGzLeXi0tAsDQ86
0ZJUNdyW6uuTb0QyfuruY8h6lkvji7Gp2R2oOjBpVKpGQvaGlIpzS4sSu68qsvlb
B/o0uO7Sh0NVsO+GR70MrCjv1JWJHM9fet6gMqT3lQhPxQOquiUUBW9bJW77cRe/
ZJnCYSPc0kW1bNZby3rlknEUoz4CwIgSKFW9qHBBzp+nbCiRfjtuPiHtZuKnWZKv
lvOjKDTLSY9R4XzSMWLc0pG/vJEFDKSEdOqYjpWNLIgBFX0ONZmugKfx6FKlO8Dx
xN3+HMQ+7HtBQp59xftpyq0l44er0rZzpvDImo1g6i2QH6KAESeN3/XWAOveHJJH
ZghhIcAkNVEh10O3jWXoiA00VPqobjijggIarPFvJVZiTYnpRrg/H9e7T3aZwF4F
YkH+gLTM2DvVSyZr8eZh5/ATau6Gif6Flga5nY3F/syKmo6J82mvP15euJiHtMns
gpk1eOgddvLPon+Np295GeXVOLHOTe1YPbnuIPEL+HpZhypoemUOfhiI59bgeID/
kjrYtRkFFFh/6aedz7q6B5MUwpyxkZnSCmmp9ivBMGW0AJwSTOiel/qkB1Mw0cv/
RqaG9x2DQ34QlY3SStBVm4qUSqSSikXrnLSpN9u5z5xcQwGDWL2WkdFyOTC8WGEp
Wrz63m1qSDrid/ypNWKewSKUChofwyJpJ8A6bK7w+4D2a6z4dyZXZ6XUwFdto+KJ
oVVXPrtTMgLCJxhabuyK+WI6JX3DfO5SesrFYmsw4UYe/8jqMO7Ic5rxoCvABIW1
qRyovR7zL0uDrTMN/kSeviRFbeyKDWd4PdddqV0YLRbA7dwX/+4X/2TJuw9E678K
TClYTrxL2GP/rdpqhtEamBl0C2kssB2zdSqJLEt1tITiS27XqgCHRwPkV+5LNq1H
lUQnyS0F5346gwNwEpgY9dG3N2i1XpUsqrZZTjssnHhTJYfA9jVbCOSis4lBOAcg
eDWq13LgjHsdYWajj8ffNQWlcglRWPPFL0z2jpg5UdKjDDafPiVvQbNsFjlJg2eT
uRcO26f3ubxY1FHxR8LjUKfQX/T5IXmlMVHbAOImmzY+OgFhHH54gqygxpt9YpXb
ob9hu78i+WLRxGX8MDHhmi3k8MubZth+LxIqcj186z0zSZbtHH7ucGljhqzR+u+a
4EtQsZ7ay535qgCCv2p5cwtmkjlLp5oIw2KKSdJSK26Axkw8XHMwwQNGV96pz8B8
IakoGmYL0HsL8oul72mP5bXUeWo5fvuM2PfL+Me5JnkUrzR8eRkxhNUZhBmN1LdF
HJj6/W+iHZ42rELh+2gXPBFwdesIQfvKWeDmKe1d/FVkQLAh8bspMNh/WS46ziAi
sICRzjtBnfTpn33xqnq5GBvW7pJALGpkgwEJLHcdcfNgXL0WAUIiS2K92Lr1W1Mc
Kmq3FEEao72apGvwrFaJ7/y6Zd3KEJJiAe9n93/I1/mzg2Ykk7qBVT1vRHqRE14J
WCgZ0TDqCjZOAjpfOxwbGvnSec84uQLGZDKvdqJgChhe5ys3pavLUIZcK3oGY7sv
MJJW94w3OGXegh2gs6337fTwqAIk7+p9tjkHqKnepR1lZErDreYX6bQJdC4kRfm4
adgYAVAsYugErQKgsm9bD15+FhwyugecBVCVNPTGJflUpP4O9CQwhuR4xr2CckRt
J6qJi5jhWflQnDiFMNzMkgQtPlvqjZsPWQzVOHcW9a3qW7yFG/OwNwXly36MtcYU
5yYTHJ6027Fr2tIu8AU3avb/cC3qaZlDXAeBLB1p2dOOK4eoy4xH77DCVIfU5P3l
OD+vX+xHwf1QODrcikV5UrnMMnG3w03IzSPH/hNPNA06NNcCkXgO2xaM4sO0F2pK
bxsc3fKWrSOvlTpy2PzOspyY6YAWvBIfb9Zvz9eNHwk4FaUdLDJRCUQqYO7+wl0O
RhNpAaTgVPeYILF7mFcC/S3Oye5I9Oka4l41k35eFEUg4UgMh9o9D2JpCPfnYEaX
m3jpltgSnqIxlmmPokJv54LlWffuIEcpGXu2kbzEhZsim/U+3X7ffdJrsG9AhaSF
mlYTO96HuUe09Ccdf9pdytpijCEcGr4tjN4CBR09DsUONvbl2Dq6OfeBwVa1ar7/
HxQWIFr5+hKwmjsp5TmJTLWLfpAe0RHYQTnHqQm6Av3YSNRniKbL75ry87DNM9OQ
k7XVjM2hmpA64Qx9rEDRJWIblrUaY2kYeGF+qsLG2eG2X064e5+CCvM5flh/BlZh
byjv5Q9eOJFnjfI2Yr/mdVSIiXCT3ETcDHfGGhS2VCPkRjeVwVQh/P4r9wusMEGh
UAuT1aWrCK/kc9rAQeETn6u1SHoo0uWUWeYB1HSjwnAwmt0uxdiJuMx8BX2OfORW
g8Bnw/DBV8cnfDKymFhAEox0Xmg+gzUnImthSCBlcNmiWqsHxCuxSg4xgIhEJ73T
atBLzMNJOc8wQeMGmJ1uKZb4Dz4ovrrz5XqdezExL/4rG39T/pBrnnzdt3b0gajQ
JBJ/55nw5SPSjN6bkAkv37zgsJz6QCy1zr9kuml8i8AVZy8+BYFF/J7W7CIiwXM/
INJz1/qr9oLaTnArSJnr+2OgRcB7HmzMYZ4rFc5223snk7AZonuHeBWSQ2F/+/LB
vzg7EMjBySyYJa5cK/tNqi231b/iVoazZeNb/84tQGGDfzxtQTBXDqxhSCidLIPX
sdFaR9aRVH/2T1GSyAAe/9s/2Y89yX6vq4pbvSRDaQXO6rhGs9DbHXxerqsAeDmE
h67oDbJIgBwSVmZAKuyk043PxtXbr21lT/wUNUTogDbh60MCxBGeNNNPvC+KsUzU
U4wEh5vnv53Z0a44IaGgJLP8Mw6nowjQX6R3uVg9NsvHzGCswxElEYmFTM+SYoN6
KrLN9gkNFoeqC0KzSyeWGaXvQQjbq4DWl8MZ8Pl0CKAkEiOeC+TxOwPWeOqUAwb3
z5OPTYi5yqD+UDAhqoNJ1pKJE19Bzpy3VEBSVWthHOIkGXgLmzAsZ9c3ZDcjRAbL
iozITjMKK60bCI2db4UUev92qpqtTqP8k/e2MXJ+qsypBqwKtInvoowez6HbhwJk
VUriGsxK/K0IDERRpDaO0Ta1gI11G3Wn5OjyufaX+vJMoNXkyQpf7y/mybexAisQ
jBZri/fvV6wVpZ5EQymtkJUYfVKpCl9vu4hoHXzf60Db5PvFEUBZR21iiKsAX+xs
2uubHcwvUjGePX94Wt9ENTlgDuaTgOBBuo8c9F1G9NNTCmsvJ7HgiOW/kZZxJsBC
DIS0cHhVteN8S7OzLP3DplDeW1OUJgtpjm+HSEVTvBaQyLXd/fRcOF3c1sph9Ym4
TYzj6txtkh1dLloTiVIa+PUrb1dXSfbsUaEUDZTb1NlF1FGZQG0Zj/tDd93aCi4H
McYn5Mj3n/6yIUkCncFlN/yQQali/3gMTduth55gpJnjNTVsIUZAOnpgvcfqtmpB
jYNjfzPyCHdTHtVEReLSh12JLSB3fcKspQFsnfxjw6prToPoMtJ5k1hskqFf8XJ2
c+B17jsJLcxCZPF0DuxZe974yPPIi4vJHWHJBFWYI0+rt06ItkPJpi3XBkA1mpRh
nstHV3m/j3K5kQKeb4q8BsiezEiSfD9E6MW2DQW3XO6nIuotVVHaIDeiP9TuTEuY
slsSJK3HKmjisVyBjsTYVP3s4WYSm6pPl+G0s3FxvLyvzrx3MVQ6XYwELMb2nVE6
/FvThBko3TfkvjaCaFeMYSgpEtM4n/pEUyYks/zaZbkdpbb+YxH8nS+9xVXjD2oR
WSQy0pQOn68nUkLkyZduXptktuXWB0PLFlEfaa/xfK/uOampGYHWMDwR0Xcn7i4k
YwH7yl95mJ2pjoE7j+ODMdXOdqqba82BqwLscUO5oVN8iETiW6hAj6fieWqIS0/G
Cqt8LL+mFEcKfwkEwwzrUF4vFlI0I2hjsFeb42qn/emSv5pz1k1TmgfDIcr6l7yZ
noMwag2f3L+mO/EU8i4dZsu92bQubaJaznouFjSthVMcWrmkaBb095gzf9AHRsRw
dapNRvJGDa5dXc3CVM5Ot7bCbM+NAWuyR16wKKjUMgvxHrMdad8kOtsJyZHTn3QQ
Hl96xbOmiZWTpqnNmFYGpfmbleL1YBSa8odesH/Wkrl0m3LDeEeMtjzXrLV1YZ9m
H8Q7G6f7prokb5jmULvIuk/+6cDQTvGj0b6Rqfs5GFiXvmFjlDWtiW9dGPLovjx+
jWV8aT6R8OOI6U0XLkf386/YN5VHvyP8jKnieB9oTQ7+HKs7g/8VvKn0P7hi/k99
iu9rrssFMDF+e6MM0LxM50QhPYJEgpp15mG6g9cIPeQQ2XmnQQQIAYpvXFOpgxJA
IIhQaoSv5p45kZ+Pw/GSgVQrGRuOTMMk3U+wEwmLltLBMl6qdd1YpGtnhOiLYQQy
gCQ5SYJ1ecDpPg2foedyPE/Pcxfo3ocr4OCbL3RN7lsGJcKQtjoFrsZI7FemyjUG
/t1R/ZG2uOlx0VvtebE14sopmPYaqmkQv8A56zJG9RQAw1BcYIgMGTz9XlN1Yroo
vNEIuRQeEFFeqv+VcHWaRPUcAOj2UAgO+qMC23xi34cn5Kj5wfS5IQ/VeUu+Mu1z
lEOkhAklAj5Evu58my6BFxrsqnQYI8kUmXPX1Th8SzXGfiFMpC+PnxnF+PO//0W/
MWmDxTfaK6C5ljXv5yF2DNHRtpF/7pwDnjIsXMg7fxg7/6vKY0kXMSe4CgZaDp75
mgczNQ6TGzEfruIv8GuwOGofNLCcrGhvCLg5IFPsIbKS4uA6ktTw4xClJBPB/j/7
WqH65Kaozxjqkj+Py4qTDyWTypJ9ipsx4U2tPTjxiKhRhQqAFjCIUaNfu5rv9rqi
TV7rFtNjFBFEVnHSLax3PnC2UxxOaYucg05R6pigfKscxVqyRG4+OsYKpulxgdJV
x/02FrjGxjshFRz1II+6+p7BcCw1M1h+eFikI6RHDyRAlqcDMy1A+l6mmpAbYB3X
g4EHtJegPK4FzuKdsR0k1aO30x1x4YZBE4/vfKtSthKAbA5+97MXTl809t0BqAKk
PHeOkGEusD4dl13LqxCKrzUzvAqlWblEuqfgFyOklG4OMUNJLokXhTQKn3SrIl7v
XMF4jQ6qPVIiH7y1gbSua5Qa2Avrr5Jv7Z/XeEvZlaE6ffOQs6HmzPIiZcPoHeiD
XIF1L+hMYXvPcFpsTI2iSTWUWXEOO7zet8cp4kDLXfuH37daB828v29tq//m0F3I
aHGgH//COvQ5QbXpJdP0Jz3k2xTHhUyxrrnIB1nAzDK0/nFL2lrwc7rm8Bgbh+/i
IZqi7yTkfu5XCNijAJa6cvkjyvf1BF+yOmWLGpHdZPGWjnbZF7Vi3pQGyNz6DcCc
M3MeZki1gEAwnL9jwqiYjiBou0SCHdxM20M70IZ4alUt/9qxD6aRv9hST6VcMpul
iDYVteyciyOln+EAnQ/3HIRNf69858F0uIMeopojPcXfsv9Hw9TEtPyeuBUOceYS
AZ1YxEfW0Y5EqQbABa+3icxUDtpyHx6oCdQvyda7D81jPNZO4WzhhzfzlZDVmNUO
zIG++hqfQ/cemVJZyl0Cjv7gTO0j6zUAZwOStiWQuRt4qPonQSGErqrORpBfp2+D
YWiEy9RhrltQBcnfDDLrjoCX9RaluYO6SjUILciKCuJ5fYF05IuSmsz1Zr7utr+5
xbLWHDfzCItfN31MmEnc+uaSEVomW0fockbeIfcz8BeNtzFiYBSXGOCiRBFyMf6v
x1L2LjTaFsEO+JMsBLkVXzFX3tT5cq+j07asAM7k5+0WxpYLZamDaZ3/4oRmzZvC
nDs+wvS64sZFDV5lQ/f2RtKh7ADf3L7Ut7LVmIBv6WwQZ/IhnOD4QGiBAQGtZF3A
gIZ78bWfGfmLPXgvDHT4lZHOzjS5Uqwa1WpVy9+3uL9+/6hzjClLE2dH7EiGJxMu
E4LmMCWe+iX7UgS2XKkJPNIaoChTQR3OHBlR0PVBDxY730H6+Z9vqGQXxs8g1Kj6
pCfArMomp0us2wDFgV4QkEGnTHCVEmvMKziiotHBWux37JZcXbn2bbaxFx0EOpVL
/CIjJ+ZB8eEy6Zew3e6fmrQjN1EYIBOD0nD0amPyYTL+JjihU/lVfLTiVbQWRBbS
bECYmZFQaRGnTV9EDV+P/EhdlzwOY09n/HS4OAd1N+2xkXiSUp1hSLiXg0CRo/Bk
pJNyqKNAuyx8msVRXGWMhoDb7dXnwLYocay3oEIs80y+gUOAogT4Ihi7OFgGduND
RrjSzBxUZOu7ufhPGpvZdUnO86dX2Tz6VoWRHv5+S9Fxm4jzenxRG6nm6z4EhFQM
k7xYd3rR1srj4wgY7PXWmaN/ggYpPzmyrppJHKjWx8Ewn0odSFHJwl+MX2ZE66nS
6B9p6/BaK/Z4neokehDhAcR8Vpp8CRc+QhgfM1KVpUBmUqLVW0Emj55v+8z8QrvV
myvtIg3YPuiWDUdZfdxJtQ2ttqPVPmyKOmrCs5OBOPqOcsW2J0TjiBtxYn9oVRhZ
Oml3bvpXSHR2yaq+SRJUKICvi9Wm/6paiZbYey6TpNMpi4tIbxbL2RMI1MQO9xhU
gY97wPyL250oLnAlwCNwVBf/DuWgTyTlNDYP8MRBMMFmPXrOFIlZVnd9oA8by6ST
bwmcRJJ4+f4LaTCbYnDB3zPfzkW3wQF4PNIe4KY4NJXnSL6WA6N/FwF60Pa+zmHB
oQO5leI435Nt24Cshlzsf3Ef4XUajL1vt0E59o0DvfIoig9Ncb+U1Egxt0cc7YTD
6jmisnaI+v4SrGjRj+HkRq95EKF6vteS2DNTYH6srWVjzlup/UyxfyAQ+/YW4Gd5
HdKQbJ+2t7STrCcqK7iajA77K6939p1HBl3Aeit11NfiVt4qH1lrwC/Au1LCfrsK
YpyfqszJYpP13jCUckblbgjb1aZT0G7ZBoAwJsmJtswF3lZ5Fu69tT4Tc2xG05wp
olZw+/FaUAle8+tPahw/Kl6zt5SXG30KuRd9Rlt3JlVpcOjV0xora/DPrzGpvV9B
0P+muq4nYeIbp0Bh43Ekj5DdKxsOJusZhrlqwQRt7LQkYDhV0tofOoeVsonJADt/
z+s2FUH+cbUfyfOavhaKNIkV23iGs1Rgwxf5hiVCZvAyqISWscuAymrQo29oFpF0
t2qS6ah+flxdAmii97CF2BML7lC7CBsTLIJJgoE99AluKwQaDzsuG3SoOw35L8Je
mS03k3Ax3IVOCRNkbYWnRQwOHH37CHBmCpjD4SFirmFDdysPpYPlDqYb1mwbzZRr
xhRleI2qXQJeJTMatfA51qfKQyXhCJ0ANoM78qF5yHelfmqAtzMvzZEssGWRra2O
F6P5laLsvPSzBaxFIV4mmyqVagYe8wTA6F3VkuMnKcwlfoIeA/Veo3+OTzjZuQfj
tlrGlmdqM/dW8zxxA3k9W9wKjKYQqhR4wlfD3fHgO3tctNLeBUDtygAI71DUhae+
bi0gQjmmlbHyuNGyYcK1aqIyHOF8tWTTm2qoshH2bh+Z+3y+gTuK8L2H6+fXfU+B
4grq2EZ0Hq+Fwlc3huNgTTtEzSk8Akb5l2FB2CRubMEi0q+qb/YEHZci9claDq1x
H3zV05wPBHA4SdahfQpC4WnAwAqLmOCWt+ZZotVxYDPWFf0bWR+dqMsW2YO/3rI7
liURucz7pnLj0IJ/XDMGTTKpd0/6nxNigzdIXM0I/wWREbtTiFSJDjaH+hiRsfXs
xGLfhq9X3wjzMDQIidzvZGOcvxKsqxSh1RukriAlK2J6OxN6c/HKZiHUn9V+Udta
cnOQ93bhS4v17kQLayWzRkvsqGlnNniO+g+/y4852Vm3oBAyOGsLfi7iDViAzii0
nrZzgxjpwsocTDEtXUhfG5XJex0s1G9vychLxQZcA+JSuaWQTxCN7ODTGTaCyqRx
0CtudzVtGYaVYBrenXfVosiXa4jLO23rENIahQOwDIcTSHoci52j1+4QOXDLmnD9
8l3t6xU4OvD+lKNyp1SHfgzsk6ltbD+EgKnr9UaDYv8sY90CDwDE1ufpOfMebe5E
D3TZ4vd2m0NSL1xoNP9kD4hn3HVR5EaM2LB8onfUonGSrQWsTEh3/VI3PL0KUvXC
Y/o2pyLW1LB3h7m17ZVgIWvo0fNz6ZtWciqh32LpkWVaF0cty14cY77Hj0LruxNd
ZrdLomuNkNy/Lo88sLHy8jUs6tPN/5y09gtOHCbMXroKzwElcLYj3jfrvIuL1WBk
p6oYWdM76gr/nf4Bf2jnIj25Iw2zHyfnQXjH/QL9jYMHkqP4Cg9BdAYyykK7xeAP
sF+eAzZ5JVKOC0Wx8g8d/gs1brUmzp6pMukojaAD6gHLD6/VcNhzNiID3O7G8+KZ
GqFpmtveAneLlC9uEWsuajMerH4beCTeZa00XpUxJPWaevMMOxTPh2gKMJ9Tbd1N
mw4sHIRsCvE8XvnRGaf3sHVoVF0XN87b7K3GaArnYpC4JEUjtpwuzkMDXvjwhQrM
LgOoOLOZxQ/qCNe8CVv34tm43UKK/NZLVXshgZyqFTmFgb0mTZQ9rv2iv9PP4clb
nwi1iLxwoQj/XwNT1+ORuHdhAqQePcxOaF/u2BmVrK6QSTlhfgnVNXjDBUCHAApr
fkOWCqV8pTCEkzubEhH12gLfeEzoW4yLyGWdDE3WwIxZskywFd0xTs8XcieWAZyJ
1hx3yVJ6l2c/r5iapLIhE7Heaisc5pYcHS8OYxY7LUqsRlAHBuEFySOEh5Ey9bBx
F0kn6gdo2UBSiiUrOfmr2XI1fKcFX+iEmsSTR/CNbXdKA/j4A1cXzzftAHkXqFIG
PGnbjKBoU3HIuZe9EaIT2QWpIEkVSCabgRiL1QhqLgjlsAVmS8RkaEh53WeTTNJF
ULiEfp/xep4f7hEBiIrbJuN6Z4d/VnmnSwsXiQwxxdmrdMiq7JB9mhZJkEysP5Nk
WPz98q2dsHJc3ciEmig4ViQS/TXLlleDu6ZFSj9QExirnpCl/J0u2hHeioQVmtP0
URxJM92J7Bx8b5yBTaANkaGJJfDoG3Bx/MBxW46LxK4KS0P7dmWnMX6FJKxv2JpI
cMKL6FBXH1NKGPgPH9UqTopDZ2pEtUfLh/s0em31HgU9UatPl4ozb1dliLM7DpLB
LnpcmgERuF9xQcW6HyOaI41oHZd9zdtYh/Z8TuV1jCoaG6hl+u+1/pHZXUSzbii/
MsszfG6frlfZewTJFmnHF83yYqXgMJK9ga3nGQh9BijdehTLB193YfLl0bx8JrXK
shau05sN6wqP08kCeatG56Oql2eXbcjuDZVaMT4bmS9hGWlQeWE5oCBbK08qOXlo
62fBXKWFS1ldEPhmjpBWyAEHRvFvSi0Udl3/aF3zAwECATEq2OhHppUpIV5WquD6
JbDjjoUx6d49l83g1hMpimFE9mPguiGICkU6MTE8dZkoHW1vYhSw++dNvydUWX+Q
8Uuz7vFrUBGJlsrZSPivR55pqlOxXgOlhnqUnwRUxFQStIyhGI2k0AccGcklTJGt
yE7hFElTXlfE9YDF0RiRMWmL1eMT2QRQlc8jx023Kwh0apYvE6fM7x6ewXx9oqoC
eSrUVngBJYmkNOs0KLCFk8FpF+5aqLWVafJlPfcqR1djpMjCmmh/+h9S3Gr5cugA
9VN1QjAjIh8jjcwCAZqRJrsWKe5VSFnerimoLgvTKCLJjCGAaZ8CC5JGy5OjyM61
s5fcpGy0PPuGgP8mpoV4ZQWGIUpl/nmbVheKhoTZNElT2FxegC7MgxV8XHWu+hoW
7s8brL1fIpRKb78z7sc3CgWDgBe6Ap53JjGDea4xy6ckPetyUiH4CP46esXkA1c2
i+hZ+cVOqMFKnnSU1v8XVcDHxcYCyJc7e8Us9PZh06nStfsfvjSbyZ2iGtW6k1E7
PYLiCQKgBtB+MuEmmI3NU0fQANBMWnip8CzRQ2TGVlZcJvSU/+FF/S8Zf/z9TkHQ
Xg0dITBR3+t+V3XqQo7nzh23f83ZJKSnYJf7BfgjQvQ0T71TGvXU6+UnPv/syTTm
+IcIKvxNMPFjtngUSSSp30Dta9dINzjzXYnPSG82PaDwasjqSy2qad11teejGam6
dW1Qcg+yZccCMF7arRadLhTmRqSpHWXtW2YJGRnNZR91IB8Urrz7rjbG28D4DyAv
0L/gAqbRPXO2YrlVaZ6MCosRtdXUaujtuYaaRhwLMQmVCTQIqjBEMhYfRgSdHHsT
+uG1Ng62zLaVUwqC5zzRdV2TCTeS8gtC36VWu9+o5gNazh6/3aOEyCtxBBJtTwUW
AXXIHFtlYxGjNOBfzgDyzeZ5zCVU5QKFNLOzNAR6umnnzkI1DKfXZepXCTq4gPAd
dNZE955dCfcTO0SD4JOtcrlhuD/HzRxbGSL/Z+VrgCb9zlawATu8me6PtMefPdGC
RR6KtuDIetEiJkwiiQxsyJfM1sUbTveGC72oKC72iTjP4kAdsr3Skc+pTSHfJcAg
EiME9HnvILxXKLivRYoC7UhUU1ciopH668veVeM2K/BE0JH0SM3zoZN/b86jNQcn
h0UzR38mHfYTll3IVuD9SwmTyC5OPY4G0utreRmicoSOktwVBUJnh/q+wDtjUy9b
UqWpfAitlSxHGZGsnFwjfJYx1bXFKDUJxGw41/Azy/ZKPfhpGfsIn0/kdkgS5T5X
+k/o91KsZHK/ypK50ocNbUGCJZnKvef/W4LAhz8dlRuBeoni0l0tUdt+YQ0UZzyz
hLyZJMDUFD59tXsJ/i0166UCnwk0azntFriF3a/gPHecScUwu0oRKwfo7tXzOrLn
79Fp2LVBXf4MriVJEiJJc1qS0xi1Rd26p0fB6T35QaqFuUK2MiVWMRcORrPGyhEw
//aKGizDRNshiRxG3QvIwdsDiqXay/Do/i8tcdfbQZ4fnBJd3n0jZhF6knfnq/v6
aVaoRpVy6AWWG2NyC+JXgMFKKYoRL6LhwfZ1ikJxbGqSPeRgmS/AoTcWR1FDCilw
e0zpSCHzIc1OLQvVkVmDpJSpWMYkLAUlqukUnl5P9sw0iNOA0jLijCerrOUTmfUe
EglXY3bfYmJ8n2wCFgmcu4e+GcdhJetff+mOy7Kssvz3nD9/xk2cTx2mZp7HqfgJ
aUFCNS12U/4w4SRvcFnLmZ8xfb83iv2fln9WAv+S60U+BBhpDQ7ab2f90wKjCA9n
RnaAkOifZ2cGF33oAN8e3nG2PMaMVJREpxAl0EJHbGcPz3+Eiu1zODf8F9gAGqDr
R92wS8QokeDuRc3cqhrTQLy877bHjS4NTnPwijrwCR4Xe33ZxMUO6o53YJUI7DDR
/1YAWLwq7li8Rt5C7PtRgKgmoSSNoCB6fE01V7UMgjc3vCFFLicd5qm8erdsFVvl
a1agKeSLsNAanZUDE9zkE3BowHVF/8tx1w4zOnDdBPzTTFv3PJStmFH+sqgHTGPZ
Jm9OMDxmnExk+i4ltKbA/s87McoRDVY+qtrtlKiyM83MPoYAm/22TVT7cOCXgNei
ADcXWaBM2MizORHu2AsDBZTOVNSbMENaGhvmyzj2vVui1BNx0zCnNIAJKpQrzAYg
7w0V6BpB8JO7s207OLd0M6ViOOTJgLO8ztfo/UwOa2d5FsyR1zbOr2C5lYDfpQCn
dPdlpqlqNXd/UnPpSdh7i5Qj8CqR1/P9W1hfMheeePF4Bul3xK3J0O4VE+gwg2g5
jEqh765naPw4vSfKukjO+3X+ynexFjidPyJXB7IRLeuR5B2Za07JtjG5/n49hLph
c1uuGnxIO1oRo6pgmYIoHz5LLNbu/h2m2JjIcxv8YjF65dEyDTzyEp1cHoAx6LWW
Nde3IkmD8om4yiPnswfMZ2a8a9NR2+utDaXY2anGTvuukUnT/gt3MRzI2nsWLP7+
tiG9DKQBTywu4oj2JI8RzvBZZ6TT3AcDmEizavJSDv1ZHcbp+kpVWJzKbBtpCxV7
w7PMDV+HLWkSWSJlHHudi6NuDldRwfvl5kTZXn3hZ+rJAhHYkg22XOHmA41QV2aw
89jyfiDs8G8MdDTU671dEsD3pa9lMJLW5iBc37PyBK8uEBkXuxy0ZvQcUyBepFgd
IgAylaP+o5ahCRzjs2xfEFvgPxYCHIMPiOx0C8FHKM1UDHAiUSx0HyqztzXcQvLf
/Gy4305ekeS8ifzRctpOkt7l68NquY9uHzoddn29x/VLivehOGV21Y+NsJdl1Prq
bD8+aOtmIZ+aTaYZAnHhcVaZjhiTtXT6BvkPJy1cOCMgczFVUQUjhZu0uPHtIiiP
VI7r5BWueB6g4eZtgsLL0P7zomCpvJUF5+B7hR0sptY4OPY2PyBVqzRiMchMUIOz
rtsYAKGqfeNea0ci2EJLY8moFlrHUh3humvi9NXZILsrg9KQWSCmk7HkoledJ/iX
jYn3eFmFSJToL15sfCPWLFdekFFhLWQEEca6H3jFQLymYhRtyAz3iKFNZvkDVPzE
yGlt0ooeISgaPXbrATwLcDpWmxhFZV6wbt7aY9elMdobqHGPGK93utrfH54Cjlqe
YSn5Uqup1PkmCJgBy1NVaRoT04OOngMZB3RmtKVyi7gfeQ6DWg1Faw/vx8436vns
vfYfEL50i4lfJj/qnWfN4iSUyVMFfFgYx9k8AcRVk5yY2VoFYhMgIPpWuwX8U+Nu
oynHmEcs/kfntR+ks/Pg7d3rHxx1KvIja2DYNSpAPAH+WTOqaqBqqQB6EvKDy0NS
07wQCG7dG4F/v7dmboZv7ECHMCaU07xkC/E4ISsFALxKkJPLTZTdQNCjxxsTNrNq
xU4OO6KeGPTEc9dULUJK+BPQLpxAW3mox0+SviMzZAs1R2AqSgd2Y7GwpL/glB4P
vynLChGLCTb//c/2lhvkxHUk3imfBxk4pcD5F46YqimUf6n/JpPbski3SwZ/xuHc
5Cwx8HSMzB1GIqdFlh1Ho1xfau9iNdKOVvA1IhUEqhLG1bFf0JEQv1P5hLjgORsJ
Om1QaQZQQsssd261/TZuQWg7s+AF1kMvdIUjhk834qASjUG0ExaDIDAVC6efHXWw
6ckXam42kkF585FlVs4lwUCkQeil7tYFBK97ntLttD3Czhy2vfznYqLNI2BlnV/1
KdH3VfTNOjuJNVz7k6jyv3MGNvG4Z0QAa7KJeDdmh5WKenCr/khEs+h5Yfhan3Db
9gjizyhKXughc1S3lyyQxZvkd6P7jn6TPiMPZlk6D0GX7ByZrVzIGC6whq+C+uZq
k5L1kS0gj4jFtujQji/5tmTaOgK6q/Xz6VNWPgufY8xWHozEOYR/firJo97/S8EZ
2jeCOPttKcUM5pH6HegUgkSnqcZj+m+4GMMMMv/cgl52hVAO0rmem7v22KY/B9XC
XwCueWlDHH5HftEykMhqgAbzdY/CNo9kqZrGWj4zxMlXxbnfIr4h0KiAEyQQZlai
7eaMUUfU5NHgyViDTZmYVDGXmYiBqy6Kh45jyAOGVfEiV7mx66DVHcNqmAGGhy5b
4vn9EtKR+pZFBbS1NT4Pi/N6Dhml8OC0WpleDWuigaFA1u2SOG1ZT9/LmKO+QZfT
uELWftDu8zocBzMYr/A6E7rGYfNvjKUE2JRNPqx672mp+x9S3Qp4/12KEwzMxXmu
d+NbyoS7fCYNuJ3pWW2p3/Xa8alGMYkyNA7EC9hyN0SWJw30M/D/IePmivdPklXi
3xdwnul+aIsXZH70XtY5CWpKOZjX/jsJQUNcw8jgGgGLGsJroScbdG1dIRDNmVkL
pDpFn0QG+TAU0coDjW8KP86ZMxX0MnetD49qfgHhBzkQK7gfqOsNQGYXak9esIom
zoyD0LfwhgJFFWguhfsM/TILTZNi7z8RS5rKDrzqRbHeFvv9Xxw1Tx7AbbTcTt6r
wBf/xXYLj5PUv9otq4umc1hu7cL3zBShoHmzepnYXurwT5GzvnS69286+K7W0esd
XOHmSkRr0SDjcH5MX2V5mGNP3Ap4gLYJkREFVS5X7HGmcuM7KILvTm3trTOq2pvI
Z8zdKBGIoFLYTT38e6oNoJUV3v2H6ZXbJmOCTxlFSdkMOfzYYZR1I1FXJ/uHcIqh
QtqgB8fRyg1qBRCV53JjYJGB3gO2yUyQ9gmVv9maj3R4xYMju8kCeiDM6HDJTT7I
ki0F/ShrUL4buwDilnOTZEi3b1yRN3ljl+TK6UT7mEGm61+15LCKix+XtBz68nw9
RqNODr5wIQv64YqYfsRZivaJ8a7db51FijAukdxcFX/0beBAv42TrAyNPcOD8I4H
gnx4xTsfHV41tzaHPOeW/nbUnzzPjdATO4Ct3BaGCeRDQRsVOSJ0TlTkP0vfLSlj
k2TdhTN0d/0FfUSb1j5nvtqPc4mJCzKAWWEZ0y4MpY7tNGn8mKScR7Gk0KFnIsJB
XIzCfrzGWopmdqFJhvj6vPE/zHcudknqL64krI0k2lGESG6X+EQqXDijPz92iRMf
fbC4xzXiCVj8td95Mu949VnmMSW2wsbpACVKVqf7PWY5Jj4zMihEbl7ixk77BXgB
oHytcBIowvSdgLvVBHxxaAFPIaFhFu1dthxtj6FGYrKvfg73gwlkUyod8cogf+sg
unER6d0R59x5aOKuVKsM5KvHJicC6jKyATOL68/wYtPUIXQIc+e5aoWx3Zg5zi1f
UQEpQbbbEZTqeBkmS7RyzOYNPPcbqV7l1yv7Og3W+/S9RlFQpbltk0DCCzsr3hL+
uYmnaFq3iuJN80HRfWiu5EdjpP8mjVF7NV6JikQC1vzxBtzpqhl+RT2LloBLliUV
DT7jxbBitEemSKcnzHynx97fsGQrjIrbamFYd4VR4eqPLJhg477uQYHQGOvP5O3o
BUwhLuJAxFl+Lke5dw3WfG09eKz+mOsLfF+k0CqSh98eTjNqJpwQaVlhDzJCzMLy
pXOZxhfpBZy/2DABUfSc5FpqbaTcN0zVAvHkKrMaIPoDYjfMFpyngu5TaA3MEMfq
67LmfS3TmFGtiL4tKazLwqmLrrIJc55mMimlM9/A1asjXQbgF25KLjbyWtvT3ZAC
iHZ5PTF2TtcIphhUZOdSJTowr2mle1qXmte6WL+1gntIv6Nvi0+ZS7krEqvAhI47
GsY8GiGM/7NztDYK3YQo+Huv8CiuFMrnTEiK4rLClPe0BHYC2zlOt4RTTxa/3NEC
86YA5nrqD1T7Nqjcxu25rZmE77GqwsgQyzRMX5Rtb/0g5yKFKM+ar6QxmbUBzZwy
TYABt2twGMNp+V9NeBMFOu5bOSQH5os8DAv3FBEOntsTv5rsWxa6MsZ0rqI9MU17
9SMPKTVOgaZ5CYsAC0fV5ycn9xjxgR0wpUmEx2UEr8EnzcOn072Ys3aDY7zhkWAt
+4vGA++SYvUSlzPAH11ibkrWp5jHY8q1+P1Tzcn5iG/C3r+NpboEXHlTfkFxHDo+
IL95HdeIuuMsp86Vwr8TRmdz1AQo2OjthncS4Ekozmhd74COE66WxNhSSIWwmr4u
ectN83d2KnVBsKtRDXG1QCBuI2wZBcYoBgVWFIzbyw5HGyb2GII6FPD86sCzuZnQ
CgqqdxtCvkm6zvhhoaMytS9hVruT+xkXVBzYGtMssmAksRKPPzy2Hb5Y5SMZOOCy
tTFbkXtrXdrfSpow3IM+EIRfTXdPOmyMRR9oqNRHVsvGF4LDqHR9xIbxtJy+W5nz
vSiBVKGPvJRAuPJAV/yfmktHYs4wiDAGZO/tcVhlSFBGR/+Q9rYty4Y/XPZzUltU
ujwMKSynY64xnq9NwN3vtSlQA5hVYrm8fjezv/hKltIeCXifJlo2qEIPBB+xttk3
p4Ucs/DExyacQ+lP8C5f/0C66x+aj56+o4LM6YrUKpjjfHKvCilte5Hm0gmBMIFU
IhWosGdf+sdnndJ71/ouVDwSX4XocW2seP1mYZsg5pW0hvVaiMQckV3Jw0iaeXjh
Qtvn+p3/Q+jxf6VOdxScfYloY8CcdZgVlLNc1zavQoohfN3gMtMqCd1/jLZ571SX
tcIYT913ApsSqAaXuePGpvY7yGXeqP8QQGXwVT7ld0uGXeT6p49te+YF7H/BmE58
211lfMHLGvsrvBXeiFy929/Q5uwx6Mp+BpJWb6WqMtO1cGPXtDN1TbxfsA78RhGd
PLqdGx1gxYFAYdjpuVy0cyNBJmAA7/JVmxmAxTLaVPHiqQaPWWllNstF6jt8afSc
W33LuyM8oNEP/CIKD2rxXhStQxeHqwrtnz2erDj9zwdKA2xBKRg76z4xf3bNcFuc
gA3dWQ77n1S/Zd4j95+kDt9xx+C0Fi4T/oG9zVA7/PzRfrxcAWvNOlr6vHBsp5Tl
wGvniYHHY0F7dyb4zs8HKRCIrtqtmvBpQzAYSqs+xAIQcDKRVQV6SJIq48s57Amx
CBqXCMcz1KtLgsaSZ5E5NGc8cjahbCChbUzjYJU8O5yLMagRpn3Uyecaal1n6e1J
X9e4sxSkqonYujiXJ66NkP1064mRuIgzgSF3PPBgY4K35uLk1yVGephvBOKDWM44
QZMxV6peS0qpprQ8Jc3jPMH0JPdF37SoZrooaO7tOqJlb8xvefVnmPLhf0vWiiPY
rj1LNkbhNDIxKDpPeBF7xdElXXIGAjHuJ1JJkyl5fLauoQAAhDfHKBwut5PqtBL0
RZfKTGn1M0OFnroQrYIAZe9oOQzXriD9SZaLdJaPk/FoiJdlMtB41ZQRVq3Xcb8w
yLq8DIfK9qex/HjjVF7LHPPbTkoIm5JSKTauFv/lqzzBR+nTj84QPa8AcY8wwaKG
HnWryMSVq4gBQzY93z+lu+SuEQgGdaHzCh2fsM+eoVqYzJD1bNbY3Ep14qD5vh69
o1/JwdPovIDLWw7O2J+J6pIx/CgYLkWltY/EtPBvNfdNJYrYFdkdFoBwQ2DHEvII
QPhNct/dN173v0ebDuhULIqCR8AUU9L8tWrS4OB6RVUsdAXngJVUrYkC7gumQIcC
9g0Hz8PwRoeK1pWzu7ObIeGk2WnINvtue365dJ2uBClXdvxg0yUgmANT9jxj/a3o
+sLtqo5E3QVZo5YfMsJ/gHl2K/oOUqwOrUg2j9EHOqEmXGcYmzrr4oZnX12PySgg
z9hSmVb7WVxzyoAzIoJYijWDoQLahvntIwwgqe9jIPqucfdas+5poPKoqZHeaTwU
BF4SekB2IIU3k2BmYBLRnX4DzfFZWRjhv+fBsb0tTs+ooh77YPKu10P7WMy6vDfw
iYyLN9N88c5hnUwpNmGDG4vBhPAYgiTISHcMnfZRvQ/iC+dWw3Iz8Gmoy/SpPXBr
EwKgFQVbmPI2YxF1L0b4jKqNtWyjRYtxj9I4H1/ubJiRdfxmFufvH3mnxcV5swGv
x43NTIWeH2eODoltJbI7ZpCCzdbcAykDcgeZGZM8BRMOsjlu10ve2hFMcyoHOceu
vKrF6K2FtyGOkgzni1Z7G4ISH5dXpzK9Q/3s3C1y+FIyRvDL3bj2nJkMHZri7KOZ
yG1btNhtX5xxK39E+Z4dagJwc3AdR5R3nrWZx5T8mXXqPIyr7C+Y/NaOiDu83Cu1
Dky3Covo41/T0Rc4aVKX80TllAWR+glk8weLf3bVim0+Swo4nYwldw79W82rnNBR
cLJYQZiwndt51AQpbxtxZhlOG6r8j/1DHDPr7JANOe2Oc0lqqQaRyEDUkJyjX73N
m+pfTKH8JIguwGoV19EVbWcjVtxkq1SHQcXBWHde/7HzL7AKcWTDlxPRTFlVdhNt
SHzbxevps+f0xB+FHF5ZOl/8hvMNb5O2CkIvRavGmOPrLYkFAik1Sy8u/Nkvgz/N
7NM9WQ3zJfum01uZXV/TGNPXPTkFSQ1hUWcOSR8tm3zETo6tB3LYZ378i/9xpjN/
2zM/CfEhHLV+3I8OUjH8tkUGZX2kQPjdG7JtVU2J2K8rXPQWAKftwh3NDLV6sir2
Rokdj2NHd0PaoqON3JWSwZTMLO9nUxJEZFMmC4BEzvy9PxfWPnX7LbuJJQGjwwW1
1pxT0aaQxpm6uQulOqj9MY1FHND1QH/8SegFoORJdjfyYivPy7fcTthq0Y7U6/Bw
fVW1Pjr2hukZZvzLr2L9xuFHrgZo+eqgdbd0ZOt11Wtfo+C5O/qfA8rTE001kQXP
i1P9KoERfvuWQlU2CuKaipOy0T2Gh3x7NwWFdFUyR5nZTquqJ2JGpLTTKxgDdTSF
7zGh6Ru6ZLAF3FlpBlv47hgfRdfgHgNEWsi4bXNkhUjlUHAkHK1R84rUzlhrm7mv
Sz8OdlOOWDol3+yOGtq/iqxpohcwc6wZi3yltf33/sHxyZK/zx972ngTK2pOkwDc
GADZePD/2BqLOByHwTwW4tsT8v3gET1KKq+r5vtRngBtWuH9uDGlUd7Oagshq3rf
dN5Ksd/2aJHka8spCJzXefQ0ZMFZHLk+ZX4s8QzsxEuPyRf7PuMQvN0odLngMQQc
B0mTEt/Bi/8UTUCUYjHPDw8H0ZvlHJStaCKFP0JbRs8cKOEpDeDzOHWgwtJnRxlc
jlVz1IhFf11Sg8/HFXnpobazXD0XRBBHSzMiNiLqhPUAqpbZldehKIs2mdcaezHP
i2sfIACQqiUUGW0OiUaBnl3BpuL68eFR5u7xurSsO/iQmgc4sVc51fiu7g6GnguN
+VeD1AyHxq3nHFbfUpFOSN4NfnezWdUnkrcRouPqOzJQ9y0SpGQ4GREuov5j7CNe
2FENbE0fRndqn6lE3ZG1p5DuLA55HiFatK6IddUsXyGa2ApOPf03IPgty5yWhzrZ
G2/+RMRrilt7ZMQ9kL8okImglTiEsh0cWup9i8sM2RHRADRMPRGxtfHRfItnfVP9
IeLgiuTLWEqhuYn8+zgOvtSZMDu6PpvcNchUqnkbKAZqOGuYlhT27AF9gniasJqy
GBJkCzDXyvjdzVnH51sVWHhdv4EShcu4m5/KeCvY88m8s5W4NBN4xMeD0C3t5Gzf
CSrYAF8krUEzhYK4Yq7AuCgNOcv39s3HUVxomLnyeHRLTG8ghr51YE3pPlOcPpOh
9CrGN3qNBf6UqTvIrnfcPVLPIhJQnB4Z45iEJuntCnQTPa5JFoosUhLkybMHqBdJ
ZnuK4QZYVhEr0tsz2K5J95ws7W9gO0F5c8l5BBWlUvBVYCAU6J4h1S0BA9z9lQ/C
44fUWlRLrqBhnXIKzsGdx4wk9/Ia6swPCBXJ1VZwY9Zb9tmoICyy5hWcvGMQrpLy
yiarq8OKF1HNS7FsvxVmDclNN6BqO5/0HO92UEDxH3g6DMK87f0buvSAeMgQG/V7
Z46vswLg3z+vO6eC5zny7MHb5ZAfZNkkzIaHgQtJLgdZNLhrqkd15tloWpLXygar
7nVo5FVa70flIW+xWtVPk5upGRWK8BWQYINZ5bFnNZcIFoJrgcUszGejtFsxMLs0
6sE+QHNMqguANUozw2afzi9CG/oYPHNa0Jg8DIZm+CFPT5ed5lDDrRNQo/OaHg+N
wGETQkIrRC39bEAkR2nMRi5y4jBgmDTWsTWhADKTrCuqQxK798YCd4T9eWeAMxVM
SBh3dgm3cv5O4hOSa2XPd4L1juTpsuni9lBFJEP+qBNNbaORmaQDMa7GO3grw75P
kMXDV3erbDU1g50PNkXFH+MpGhZG1OzeXzR4XqvN1g88/MEIMiLgkh+7EJ5YvLQI
84xovlgAENNbnlUFj8ig35Szsk5fBZob/jGNRaPZlKuaYwxEf14dJL/wsHE4zTo8
2IWHOqsCTz5OAdJGVB5sYjjzXixjUXbsJtiHzz4zaL6+qZF4eVYiDG8/NjF+UBDY
S8XL/NQpHM75mYostPSSOTp+4FtDVnKDapfdJAMkpnaMzzm45z6XdGmxiuHI9HD5
Te7m/gkenLHAQSgoUSKEAng5u/ifi2Xje6LLIk6A38YKJ8eWiJi1FxoSwfE86Q9L
pkDTFz75Cj9UJSpeV3uLM8zDup5DvKARjrBGbkq+vlkNghvtOdX39UowDWD7GyPf
QOcjMYUbFG0FfhuyQbVKnk3QMO6dsgQTi+ptHJ+fyBUoDWbniLyDXOMu6gpEmbtU
b7rZVXTTDndDmYOBwXQeBLVBnvB3d/ANeOfpDf3/3y1kutk1RGwMsq3/3meS+Xgc
UCFqIPsVVhdYwMv2HJSyTz7qo8fCLA6yWiKZ6fCam7s6Gb18/HmSqrrqKQLh0uK/
hY7+9zdPgj6pNQ7JNpyfazBtlMLBiTTKj2huHX3NQ8hhtUtTickYCYWOePOLYucK
Zd27VamohTqa2R0FGOR22umtAO3TCHeJvOqWUFTWauJRTTU+xpZf0hX9dNUfImhs
zaw2XtNl6ZhXOQtBHM8ti864GThFRsitQcSsk/nkLNI//j34nQGNpEULflcLqAGO
UMl/t0lL4y/KhXIYcUzrTe0rvR8r3ZqLuL6YZOhzyjDvLr6bmDsNMu6ZVkODu1Uv
9cJnGpud2HB8UvDMIve4N5TZB10us36YCUNOzQhmwZsLFjKi06G/sW6kAGYhkWYr
rPCztGcI+lqum4ExwVFU70jzcmAC9U2bWdpBHyL/WVv8Smex84Ot8ZFtL9mGLiOd
Rak87JyUSN9QRFUCFmEhpKeolvyUKeSAMU330HYtbi2jtQimXcuWaqZIEK2nrUMk
+aElHp8+tVEtHgOY+NrxkYIyhKfI8WwjvBGg6k9rQNMAVOXM6gX2qayBP7dqJd8m
1c3DEoGKQviFFB3XINqdHQakzaLo7r+tKpA2RmAs5SspunGB+oX77HlfOlU/0qs0
VB3VswVVUwXPU4ntXOfKqdAFzCEASky9lTLzl4+fikaAwwr93wpYT6VmvQqKnSxj
bgV+natD/4Z8kM+f0RKPJAI1LQq07iTVYOzcgZviRL7ncK75cFgDX7PQlfVX4+QT
UQEjvc8c8iJpwmhoR9idX6UOCAj9TVogLeANsaimu1qJGoJMkjANffAwn5hMpErV
/90DZbzxYmMLDzNfiyuz82IZvcE4Od9kfUFZtPrrB/9kbvElwfVgXVSi70LJAsvN
ogn+R94/WPtnNbgsePeVy6nV5Q9KPHEc5GJmihVum21kqU0PbacD2pQP7zPlzCvc
6kBWeNAKptclIFCS8uXeYP108ovKXL9Qf6Qah4Qpwa1nw+tKGIx24LlXyQiQgl5f
BcTXuBterE9v2TQyPYQ/P/zZ7r+WnbSSCjvXXs0Kq0izMOJx8YuBU4DmBPRLIONv
/HtAtPyF5zb74JNteaNGoexM+usN4nmCyRxyRX2MonNMZlY8xk12W1pIe9ChcbNT
Azm2PR+o7TgfgJnGZkB8aF0rX9Ws2lZ/PFMZoarzbg4vhGl97Z5Eaqhgy6ayk6UB
slMGRqqJgRsDdKuEIPO8BbIKuNgkaSUzskfsg/JsjN9S4KC0PKBZiFRcwqKfCAtR
9EbL4XGTfn5ctvNS1YGQRF//5hKQOtkw6rTPJnxd5gFeS2h7FRmBzGRs+gwn/pjs
xl37jwpzSHlPFRa+s+nbmtX41QuWKBiSjHLqXz+DVuIeB4xaPiQQExLM2R745ODV
JC81YS35azAOH/UFdAHjGqjyqV9QJ0vfGXfQfCmLKYSfP7FSM3gqI8o6GDHef5ab
Ou8oTyAQmlC5591Rp6Z2ecfl1UpC4ayZOu0ec1Q1exDuKYly26k8UrxZx0YiiJ6D
ouYAyGeIbTqvDnGUnVfSt/V43PFBHikiMQl939g4/RMGXnzM2O4qkuvDD1FtgmER
b7kOck4D1/y/asuQcKjPA3biNxCpob1ATH6rG7B5asudVecFxIL+tmfjjYMs3Pck
VHP3nQe0q2V70C53m+cmVpCkOVqiCTkkA2rFU3VzoXlRwR/xEWsNheApRJ8t94Dz
GL5OMWGT5FJ0C7ZqJsodFmQr1nApXW6evRkl5W+AUZL3dES1M2Nd6daN/mvKZxZW
tRxY6iKJjcldZ3nLAqexzqy+rFyn/BsDmZkPwu6WIIiwkZcLoIx3Q4wLVndSN+zr
+YIW/CtCkrCYG3KF6xBVmUkyKp0NB/unheG04ooNFSA22g+IncWYJIwKxKSFvKQn
y1/FX1+goGnuJXZEkD9Gp+au5LeDbnq/B19VTV4JTFDHZxRG1hU7C/xuxhE7voH7
xfIg+84KNnFVgspTqaG6giWpcPI5UAn0br27SBi24k29u9+GnuvXDouBhTvbGcRF
Dz1/t+DF66UQGWf3Y5ZbG2b7xGcb+I2Tt2S35mic+vGWjZS5XhANl+I9K80f7ggs
hlcweihcHVrM6hL1C1Kwg0purjgaNwM4CHmmkRO6e/rO7E73EbaXohqpSR7ddE7e
1jvDeD93E++a6gjMTch9E0J41X8C3PHvLDXqR+tPw+xjuFIgvLlIebGF1IPhbJIP
Uo7jMHP2vnn/MgxoUgIv+ax3i4k5GFvxopQToDLhqlDvu9SNtyp+q6T+63q+0xBZ
4dttVz+//jmVp1wzFcuibR4YhZniU9YsS3S74Gqr+36ONNS/C9x3OnOPlGvTlssE
EylA4b40zM1W/GoLdhmbsFHrCcxRUuXrjUV7vCyzfpibTdscQ2FI4ElfwJ7N7PpX
ziSFVix3c1Yh637OpioDWtMgztrJZAF5EXPTC/NlODJF1SJmsmXdfdJbjDIxwhQk
JGY+FeqYNvHG4VsqYKkCoer5eOJ7qHFTAZ43MkVCZl32ujW/k4Qq701U1d4ZHIv6
gHRwuo9DHGuhm0S21nNm2+DowK4LY+FuPl8AMK46zzYD88/mXer/pKtMQZSjqx3b
sxNhldoCiimGoU8SgNDc5N52+sH/RBkLAsW8YtVZLjrX+jFF/mJ1MH1rxT03yO3M
cqG04oabmq6X9UhkW1VSS1zHN4RbjX9GeIdNjgsbv/v/9M5w2Id70ZsnF9B4hEsk
ire5Lz+0qz0doNSteZRxEEHYubvrI9gJZTZaE2q4RjMA7twIAG+uvt1OvSA+QXoY
O0Ye4ZhGG0TGhEDV5lpq737h6GecQZu5zRH3hzTqI9ngs1zS6F9UT/rX4RUa/QwV
mZj9qJW/Sft/wpgDc9qsRSsHnl5/eL83nsmYSHW8RstNSRRSpmoHT6Or7vtAg4ST
YTCaFju6TuRkjEN0Y6WaePrANnZAzFFlE0eR+gZL8Jxhnobkb9dVf6k1ydt8k30Q
1xZ/uXmaCnqhtAQUKSTvC0c1M3OYiedTUbf/19r5utuFiyGv2Gb9fFU0h7dSbK2e
wwRbVUPImUitPXPhUvhRBh1Y5bajKzy6/mx3aVBx6u1iVvQ3vgRiacVnmH6QJWOv
UwXpcpPW0OfT1SZlrNoWxu8IcHv0yUrxyA96SQ7xPjPiA7hcH7lUypDb4ANn8iDG
3DPqgV0vELzjeWQtOLRNh2gT8Y743DLO0qeffniRJ/BYhHBXEVUcpLIvi4PR9+Vi
uNJjNKvDKvcWBXjr/q2jSOtrtCR3X3h+a4adq9z6W9cU5nkLTnvMPbCYEmOXuJJq
k50rV2CHSPnYv1TADKboYJ0GG5Tc9WZRDZgCYRs2dAHl8N/WsNGFRXUR3Q09nXRT
5EvN2DT9yu77fFk3kXuQIBt75IjrQEEeiWUugtuUMmncuaokYxE+GZ3Ww7u30n0q
Kc+9JYItS+rI/onSkhijCnFPSTwk3vAQ4gRB3AvSg8AAAjrgsITLgEK/3yTUoOiB
qL87kNynDrp/j0kBVNA+rIo39QMc1oUmP+Z3jU/7e6/rIlLsgqDNnmvSTTJqWj23
GoE4dxwYXPC5Tio1ummrWosnf6j2wlGfV/gwQ1KNvvxq9+GaoQhQ/77GH7eLT3MH
A24Cqmaj0ygc/X7HFT7rBdLV9PLAkPpZLiowPo6DOWOSBL/sAf6PGe1scaG1R0+B
jWXOxlGSSOFYDfXKo7Q4lpV+NlBQPgz9RjQ1WcUIMRCUvc+oRPaiMo6DfghU7/Hj
33Tt+fT27EWWFGHG/UVJ4eU/7BVNJzR3ZRpQa6S6Ijdute3N5NP28HWKoBHw3Yej
mEUN4fFxlsmpOgRN/8jKl2apSb03so6SXE6CqehlAm5yxcFJLc9+b+Kf6P35b5J1
cK7mqKXotcGhrPMuHI8+Ilvxm8WzM1dp4MQZNchm8n/kTqkh+NHcbTLgzsfEacN/
ki5cRu8a6mNf9fWmMyeGIKQMsjf+KHK6X1Ns/rzs0Z+7AGlVOhPMizHIQMWTB9f3
ESvwhYLCIUfcpjaeff5ieDQO1CdyAXnah8L3qpIH5l172+hZ4iWWkQTcQCS3/uy/
jRpi2u32v7vEmmU0eD9rObUim/U4qBqPWRlWyQlXC9jkjS6NI7kvXIECXJFG6E/x
W7+9jDlyrVWj/ig6dITHhersbbnYitL3UvCJJDox6XDtKmb3YgGE3CfpePmuOJqq
HC9zkHtvSCP9ZrFj1a/uT+8nCZOuheztAi+U4Jn4wrevDKythXmOlUTPcFt5H/vK
Ov5f4txxFMMEQxzTvgsNALCwFa6dBtDRivVjtCqUM/USglRlfJFULcRsng3loGHt
2FG2GKV0H+756GSpdUrcgtA/kQeRzVcKjC5pUxAdV/bT1pQT2wW41j3DnCmOa05Y
wMo5J3FGX0Pe3bQ1QhYYhcguZBD0ACaYH1xfsdwdoUzT1zV95qZxwKoX79M2EFgw
5UrgrfOrCpERMumAZPYmU59oef6cTeLVlf/mtxlZh2MlbTRMWF9uZ6hc0JWyriKE
1LMgS9IEVdvlQkx/tiiuAkowgt4zhGskTSiDid2J69rSC6fRwe34Mi1hLGdJq8do
bwU7BDEa/y3GZrmcWQo7Q7CfDCbfw7UAOwPftzMFWzzpAq1hH5EEhsONQJdpSieL
3OsLLKTqqwYo54paGnro/wqeonN61heyiFCHCGEnfrbzoJ73kOb+FFdUpX5HfYky
CPTtDBNV7V4GIkDu+9b4F+GFCA4+bxyHBcIUBZj0AyMC8yDZB7lBX3DOX4AsO9Xm
ayhWFZ8gfFnblpWPipWJ6FpqwgJ8BHw09we31lwdR+RNCcL6Mr9lA57WzLeRsTZd
MGfi1mT52NsAs6cVKODq00euNLaCxAV3Y9X686WLxbSVLaSMQMvI0zrKEwjHFmPe
ByDXvijmmNmqJwep1F5Y7bBnnZodkwjSG4CIyp2EQbUMTH4hZK8ovGZKeKEiwnbD
gkByTFzz2c4CX547xdF3p1oiWpyUccjh0fdvvScH75JL4MTZuOFrfpKiqr/w+IVd
nRLETWek7H9rHEZyVvr8jMuS3qpigp5pWkNJUy8AbNJOHmAarmYbE9dJqf3s93Lo
5/XHcbdMJS40G1nrGv2XqozfvKQd0M+tdSTf2a6WI418C0uy5mg/rtJ/3Tusvr8T
VrPVrLyT85FNq2V1sxkwf/1rQWYlGGxJPEyOU5VJtN+CRWYPAN5wLeEjxzXwUXqN
VxorNM06RCgYMHFYldrNX2wJ4odckwNHUO533qksBvWnhjdSlBZeD12PzZeFQKrm
KtCVpSCEmiOxBZSfjZA4aWhWCRmtHpgGnOzyD2iInlaXl8w2rcsjIPjWhkdZ+SFS
rAUSc8l1TGNZohPfW3UIhOVm5kOVcvzDMSmANlPU/6nK69+CaPnW47Ra2At+qsHl
sSHmqeZEqYrzClN3pWGJKPHCJeS/re7dZ7Y4sG3Wi6mGbWd7omCww7VrUvM1QRs5
LIEFzgGsgrUaqb52DFUEy6Vck2Ayn35IiaW+XodEFUZ+yl7bznIWFQUP6hrbdA9z
dEkwlKapzUYmLSKQm2cNmPLxkJsq5QSPRZyhGYlOk+eT2NH1rUhqQXcVDb0s5ODr
mZJJtH9REl7L165cOH44hot1bTbJ0NWNJ5hLnQeFNwZO5YfZXiGWAb/a3Lf4FXiO
Zur/6s8eu9XVwt+1fFSqF8qt2Ma5pcQe+xEwPqfTQTx19tZ7MNo9bMo73jQedLLk
caG/Jr9/Ssgwusv9EDvZALxOOjfPrRSWgj0Zv0RnwrVVjOb7F/THiNePTPU3AVr2
snhnWnj/PN8zZieXHL1ooTwc7sDUlC32pqhJaNm2llu6ncAihkJeOiyxPGAyLHnm
/RP+/7XnlTzc1mLkAUWvkd2fqHYOfZOLJ3gENqdfzSQkWZP+l7lW+uQLw4Z/+l3C
0yo8vg61El4jAmCgbzxhUWiHPFmqM/00LIVvV/FyHKNOswO1WSKBeG+S2Ox8FX5S
7frazc0wOrjePRY6sVbSOQOuwvszoGmyGRRyiAWHiTeAdueedDTX92UQUxQ2XFjo
xaCDxS5zt/aAR7sDRYG5yt9//pH2gzUCFBMMzVwcRYjk/8OhXJRDFRivkro/qVTL
F589PwHPdQfxf7Cn8v0XlYtVju0/3NhrC7UW+yy7fuHqIW2S3S+TyTm5gxYQrwFk
4DzSccf5eqym29UoAeiwfZEE0Lh1OiD64r7PTj9Tm1YpPXUxy8tPUHsfNnfgTLEI
Zk7Sv+oPoj1BlAefSt8BLC0iL4rFb0XPakChq8Mdsoh3W5Z2gQxKhheu5Mjylexl
YfAatvUnRRTb98rJZyatFgblnQsY4nLmtyLkNDaeWAgpmB87hwLKXgtZszqhdZJZ
edXBGFnEn7vDKUNNn6/CLBE8A7dwfvP76AUf6qIOXXGR5Wm8Ph1AbDSOBRZnPm8w
ykKoLwdfSTSXACgnbZf9jusyNSLA6aZp3Igacb84uDEEOg5sbWcJECYEgpfBVdAc
/hm3TgPuUH9V139yXh00okj8nB+54IPoHRlyYpGB66t61o6UO/+78EGnh6Gj8QoR
ebrmO5+rXoi0IWWTXH/3pGvB54yXEQkBnMTnhin5zNGbY/CtEFMX+voUf5p/Vv8h
r4WLzycPyTVhsz4EisWD10na5ucS0MrJHxqsK1D9bJ3KVd1QupSqKkL19COjG1sc
0quH4MfzDC3KpycfDBk3dDDe14wWofE9zyNN0OVrmHvlpOSWy6MjzaJCpuPJaIpO
zE2JyLFstk0xn7RYoGV0TjeJHnU74vKfuAnBeNKkazBaa+18DNJ/x64BIC6p4jtT
8AkPzShPAYeqnl+XlDW1fcCuuk/ZZR4PsMDzzm2RWlFKz+jf+YjVPwSC+dYD7dzA
+J9vyrX4w5ehCOhB62Z75a/u9Pfl393Ku6xt6NPoFYaYkbH35H9Uo8e1gh/2pJvo
A7MU/z6fNd4ij7/4LUEzjT/E+QdI1N9eu5AaA7c0tSDer6OrzkoMecfiRRfAKp3j
yv64axyPHOzWYPTYUd5lkda3vcj252eETTJoM//S8rwI1vDlgOio7QJsjb8CYd3y
sF49dDuzMSqYi48hcFfddcAImyOkD9RsdMV+klYUEFdI1D4lxoEucAWX26Kzvcil
D/f7WzERTA2g/I7rWPjr92wLK9UBKDoFdsoDz/IKHfazHKex20s3W04baVlg6S8H
oWq22fIFkrhpdPeoYpycnZ9gemA4ht3RCDxEVr8aHrCckQS4aBlLvqKfxbnXH/za
0N6CplFCFsPMJTh0+IJc8o4qTHoKdnn+5kn2G+kj/UWk8lY6u+xx4xGbXlb6Pa9z
X//d3xUP4oJYmoPzojMXXprjA78m5j2gIx95S3XElUcfeC7XU8+qwVYMcXbLpMpM
0B1x/GvInsbeaIWjSsok0/nCHEy85QkZbCibTsbex5nhJZ8K8kB0DVj0ATD5b+ch
lCCQTRy7KkhLa6T6jPv2PdqJIOIgfgGIiiOXpcGoQ/Wd0ZS+Oh68fFSAp+JbahR9
Zr4T9k+/WXjck61eeL6ijvvk70CF4w5MOqNgENTSf5kc3nrhiQRVv73i5Umt9Htz
uxp/V6warLKR0IsD2A+AWBu5TxPIno9OiJ2+wati/OygL675uPM79GabiWklwLPs
46+abhWYbtSRu7ryFpjTz8t1B+02Cibbi94je1pe+L/Z2E6JwUEXq8L+UO0m2weg
kOYYbDqmp04NNtYgrAk050QGGybx6RdlUmJnO4goPIIy3Z0aKGmuX4Kg4qJXAbVX
ZPwc+D9m5y22y+lhWHeLXzY5/0fH3zd+mXpSRsaNcp8BOLljpB0WI2MVptUZrEJ5
VaMInA/l9hbUcIfAPJbKP8XJsc5DOvcYHv6w8e240lcmHSkL0rOFMgLxmeO541ky
xS+wbfv5eUAuOtHLMOZ3FkYPhKdjHGGtuiM3jsiwSyKuZQTzFuU0nYlWhtMoKqUz
lSmSkf1JA2yvU5OQawpapBntufO0w5rAZfsPbQFtjcBwY9uBRhbyMV+gbdhGWE0Y
iERQ3uJxJ3HFBV0P/BILt1gkqBrrgD1BrWiT30BcA0GQwNHbIvdmYuHpM7/a8564
OlktYAV9Sm2eVRbuoEaECPRdSzSHkCVf6215x7eP6JzCPtQ48cwyOzZ8U8bRLGml
agGEf93f7garAm1IazBoM7zn3CjW31XC3OEERcgm9aXBWl3PHS7UMjDJlBUffr4R
ywXUgRwxjxioVyCptWwI/wCSdzlKzIXK19hDw4kEMIrWeKKM7KXrtvelE8heFtp0
L0YEHUYhX790QYn1EdhuTpGx96gvngKFKdYtCxqB9G/Dp5nNRObR2hX+kWv5ggPZ
NScgJehK5EBhacJGv/R/RMTLdND+pVocnw1nNeYmTAKCgxpBxlJqBaPlBfxfFcL1
3YUvmuM4aQ9wGRMVxZRehJ542AGXlv6RO3Wd+cIwvaNBFkE79595xio4Ga02ZM69
puBJFQw/d/tomK5/+rekKevU/H5LlAUyZOWOpwlKYdJEBRkSUhPVb5Td/jwwNaZa
VdLefwbnjKSgnuVR2rA6S12GuUzY+MeMa64531dAZFsroWjNAqljfTVs5mQejESE
mQoFBIerNj7qQD7xwvu8sf+zf/SEJvzek3bj6BJuXk0gfiWPSSXQR08cpk29+f0E
lmBmEg51kxQFpOyL0s484w+8KjL/aKnU3qc5A4N6wzfiFI2R1nKvarscA86BhUCg
dRiO6NcNZE2y4M2KqbTUV7bcZM6OxHGo26mYLnmvo9K8oDdywholJfOj8YkfRYAj
TnXXRsGMFmXGJdWc8D0A1SImYJuqhdYtm0QcNrFKwp5vSBjvOMSlK8T0Tp78442L
SHpaSYYXrck2Nmm5K6E2owXWyvfXy4p1VYbbHqg4PtoRi2E5hVb5njrjue+VpJf/
hOUXkAvv/h/2T75hKz5+IasTjiVQmTRsZfi3X+z4NYzSY7eauq6engANo6KCs/8/
rnq+XPBUmpRHs1eqlsRGXfxXOoitU73dgf8qNHdzP3YQOqs+cyvlaxcFgXob1v+8
gtT58bDYOaWx12oouWcnvuisWQQMpGrE0oblhbVBqDOrrMiND1nIliTvkyh3pJ1e
eDwhCm1JfIugAC1mBdXHr0ADdC2EHW1cmJ5TstCxkara+TO9oUQcU2UsF/rzD5El
KFaFpgzuvfSK8s/J/yvI2lRhrCEhRDRFHPwsjbLxwoisJVf36aiEFV8VhnxS3P9k
KHW94nyniHXwkbnMCoVTtPlINYoqIbb1exAxiNiZlE8w2S5nTq5rLVy34Acy3PZk
XRp5Z3Reosy3JE6V519b1YOv7lb6GeJENkn6vSjdiwvXGr2FUY0v3buf8/FoefmX
p+jXPHZ8j7KXQcweSGsFP0muHM8fOzqMnwcE5nixUMwO/MXTiVud25zAs3GibB3+
/LqF3vp5+KhZRG8g6/JMykfy9G6Ncjrp5Fp6Wvf73kKWcIH/Xl9oTbxta7erwS5+
oTKh+BSHfEEEZCZsKtRODc+hCHdyrZp4JpBq40SngGkGoNd6duf/t1yf5ga/lbvA
ZC1jv/sl9pBC91dI+Gfq5bCeA4f1wOLlxumnOAB8ZqHdEe2/m57l54kjEGM2fmcB
cI/QGlafIwYtShScP8WP1GWNBUNUZYvP7kST0DVbuI/DbVO3+m+TJKtG/hPYaZoI
HHKvjp1HY3N8KQOR2+aNZhVxO4aQn+4Ss2Aakr4ffc33di9EOIpuxWmT7jnGMHi+
BcR/GpTDki6ICya5mebXnsk4/wR7xmrWAJ9UvRdxp6Ul6erd8JeIHi07iqVNvm+Y
krVLni0mcVCEFUyzlOZ13Z3L7c+/hl5I3cHVX+cNTP6IuEbv+k9k44fqVuOXAw6x
UEqmxTNZIUDpU+VWazMR2JD7c9/flUW6SAgueV+5SeHEK4dQrc1bQpusIa559+KO
ezuCEQFN04UJnPcwcScDWpWXgJi8NlwJTRK0zFKUGgcDDDA3oRHyn+IEDWLFs7Gi
Kia6b6va5/QQZCCKdJXkXHzdSe+Tgr7Lipkf65ccK9ssEDDCsjSXuPJCle+i9D8a
m4tPQTPMuIDzLVzU4C1boR9rPhpNe0Hx1gp6b90soO7QeWAN/V3CKNDeZ/wfD9/v
H4R+qMuAvXyss+crjq7fAxjhrZBHYvHakDsTsemHcvGRo8oOp3i7cizP1yRY4HGV
PwOzheO16Tr6ZNqaGUqnI3ewo+S9w8bU9bdb0MHbhYsi141RZUHVgWHOC3hKK3sr
9C+tcme2yD6sQIVmXkooH4+1i6+HAbVqfuXKQ5+dWEWN38pfJWN5VA0o853NhhNH
CYiXv0vBNgzk4ov+qG6DwBrhuiXirXh7su68VCr2CXAldKq+bGH/uD/QH1TWW7R/
res/ccBeGlUM/SiuhopL0M9JmgW5g3oweJ9kgodzmP/mB/ZxcSl4LVGrJT960CZ5
My3j5nWSkxf0CjwOB93QcVIF0WVzTctdcBEsXIU+d+CX1vKQH8YtADGiu1JY3PW6
c8eq/6fOQIfX+WCcmwrdOEJIFFaNAASUbHQBwuCh1OuVy19+TXlJXo0fva/oQsen
Z5/7QPg/mF6YEyFjEr1gIHQKkLNFZ5les88iw31P8Gtt9in2JgZ4uXpp+rgH/MQj
sBJeVZ7ugFx1y9QE5PPZXYtygH9WxdG4BkszOneU98iKMxkEoHPXlpcMBR0nEDfc
J5bvOvxO5v0Uu9dsEal1wBjq8gDax3x2uy4hCGqJwrAFmVgSuRCAlrgr/ALj/ikX
AcuB4lKiQ2cAngsNdzZ8a3XUJJPFkraC1u1OOsUp4WabFhR3sRiOIn+s+JjRIsls
BWZE1luX1jDm8C5Q1xxCcWAsfweA4n3YXP4/vbBJkc070PqHCf52ibE+OeDpkalW
LSsPwqSgzrNU6jxa+3QNN9Cp1EduDbV30Aa9zWHLwMASXVty2e7/wk92cRIZABJp
0RocdJpYrX8EiUTeCyO4PU/lhJ1UI/lbltWE0/mUxYyenqwz9zVgg6Eno8wn+NqA
WSNEfmEPgj1xkCjUsBcBo1y6k5+WKRZxMXe8Cw5Jt1mNOrSjzGhdwBsaf9yYIjJC
Kh6Bg7ZcGJIsMU+XLRQBNi6oo5KxykH5ZU/+yKVPjfMzZpuuxJdQosc1e73aGQ+E
MCoke0n5OXGYR487Bz135XhEoU8cRV8zxoBD5evktjuKODSI+t61Un1XrAWn7sco
7s/EHYniwaHrisjGFmiwCZbC7BZ6iK2Xvhgovu7wyNeQczJrmeIvjCwdUPby2F9j
5IaSP/9asbgsy9LKjhjB7oVOPrlo7vkpRgC85M5MnuJUJ6todLeo2WVwnqtyoO83
Zq5GSOPsXltmLhItfBOKeHSxDyHPCtrfo9ofl7SI18exYY2tWhUpdYuxgV3GZPZY
5AEEAEj0HShsv9FRk5fn4RtedIUzXCM/0NP4554JWaCq6pcp77A8a3yNo3DIqfeu
zttirhg5p1gf9b4ltr/FL3KspsMfleYCX02ZR35V4c+wF9MZR01UYXNr8PszmQJH
+uRvBTX6ho/QJIkvmj5XwEhzsHukNw47hV+vJ+yYN0J0EUNW4tGCV56GzwWFHUDN
NejUbcIFN286mdSaLp9T60rUTLrOIqCs+ZT+uCeQDM3pSGiF3VRVKTpESOsyG6N8
0lJTzeBb65xygZky9N9ASAOTju6JmLAAorNrBJUzzlZL+2K3FN/zLXgbY3NOd2x0
ytWtJwSJk9D55d2tuGVf3jxDh9K7r5hlM6c22jUv1FMg6Gj4H7BYlmjHO2BIstud
JQjKL0MgPAcywCEs2bjjJuO3Mt23tbxEAAcgxMwyXUH1qje2oiBfhB1GdxFYOc85
sXJkg1jbIgvSlH3jndc1h78dokpnbNXt7DYxYbkQSOA+iVJvZhOkeKgBYQ6n4AlC
EkvNuG4su87V19KS3wfn9PAw3diacpZOXCf2jafpFe9l3GcF/k95g4u5ysCleKzF
tM0m84/eDJdLRbU32x91ORMSJYp89Qyy7F1v24fnJneGp0hxQqSFnnpfYp9oUK2Y
2bPkP7dGfd8vABGUkzzJRhCtOv1DLeJpcFM4iS6EUI38Azpp1viHUkDUHgdd3EYW
e2ZJ8lNsU1BcqlUPeH+06MMHqeSgquK34J+qKjPbqiuc6xSXeVfIXW6D/Ovx91ut
Y32uHGS7eFqX7FmYjyXg4+9hEzA+dLklYTP3NRzRfqg3/OsUdNyoglkmDZGGF+ES
ZCf7OJJBuPRL1SoAool0KNkvwUcz5As9vL9zudHflJ03xJAiXRlqQdfudXxK4YXm
mpYErDxhgRg+4o3CW7hkUvNflnLoIggQzYi2ZZWpHbA5MP0f4l9VD8Gpj14k3cvt
n6gHeQFTb07JSGocG7rDzgvRZDLE6eTVPlNfiaKvYA4VDej3ZdNDqXmwxPB8eeh6
5tMrQamCWaJrCTqJPAmFWzhMmDfKiu4wFpV5LdhkZC4TLxRmzmcmQvcKFrm9yzAi
3mnAx6p1GLZ5x9h7Va6shMmTWwevu8vWgmjXncbgZtAr9XTyCGZAop80XH8C8hNl
g0E7MhuTImZts+9+i+6EaQAyUVYY2wrZ1l/QOPNznX2dkbUYYXDDpGnJJaNJQRBn
fC60tzplwvPrNGegqaSq9KR7UlM1PZza3YUFlbATAWuC5Y+BRd/7Q7bLVu15m6c6
XB+RRwTLWOsQjL0AahV26rupJPIh3RNIF76v+I/rOYEHPQpSLb7KGugZ8bO+FLRJ
agSI0oz82rP9kI6WnRpVx3rVd0PP23Px3C6KPcek2aVk0Y3qPtA9mwHgwqRxiNqm
zIOaQRxrgioDzjGGvewPIVf6jD0ULY09E2iAO8bhUWKc1YVgwBRLY7xAIjuBTkSG
RAqD8xHo76je/gDpvStQwg1DujrN1XHvfeYLXAt0MJXMXwhgOOSy+aNKgC78BIzl
t2mMms1sBuLhv3Z+SeJqQf7Y5j6E+ABv6Z2/eIb2ezy39nJLIpzAs5B3pKF0vMUw
wrKLzGv8pwTlB9c0LgXm7eGHUadq02Cfz/qjZl8fZCzafwsdCfoe+j9yIHtLl7nO
UZo+QoUbYs+T30i4vpWwx0QxcaCeMf8iUoVvGVUHIekgGbSeAMj6cv7xl0O8uFc+
LsrYFtq9cZQK0Lo6bEYy50q9GoIhBI8yoy6sH/1ZzoKz2VLwKQWDiKXKY3F99jp0
CvEq9/DJtqbMjEqROx8Sz+YaGFGMTMl6CihZ9GWeka+4cdd9jX8PVI+EGYatT7Xp
bT46Qu6AKyLux8huxgO0/KKFiqlT5dD2fENMpoTFNR2MAIXfD7WwmKOYqyX144RK
Q+2wAObxohZxJb/6kapsSGCWaB9UzJHMl54viOpBFauhIrwwnM2r7mCVtQ4/N8Pe
5T6POFklgnBiDfTyU5FjSkTBsw9v+pRpjqfc2iMM8YqyVrx9PkzvaZd5jpJntoIt
tDEw8BBmQDS5g+i0hNBAZE0X5phIXpslG/UluVda2wXp1hk5vYzHe2SgY7iF1Pbw
EmGqMN9uUIAgq3CPomVhA0msQvBxIy5LuCxOFUgPt0A4LR3VGSAu3iesLjcL8/qh
zmN79Bt7Dr5oL5N8tU3ujtNgz4QDK/pGpQUCmQ16C39tOp6KVKv0CyShM7m0n1lY
iKKYwB0ysBRawI0e5av/z7Q7/05ZXnQcvDQlRQQX55NjUdkecPILQUuwMbxdvl4R
ZbufRjGB6PBB5GOR8spEvqZtkQ8c1quQ79mizXu5i0NZ8vpHF9vRL3OdHVTA9u+P
O/UGqXdqVIgUawV0Yrguww/EiA672Ite2Da2Rhb6WOAFOQS8py2BPkSGJNazc8gK
zKuXRmT+WZGeb+tmYsh8Bioog7OwlvxFSxK9BVjx8lXx+OeKb5ow9FRptvuj//W+
jj+qcu5/1a8Q/4hClWl2SSM4RKaXDiGfWvZ8LF8bsoa8Ew6Uo43tHsOG2t8di6nv
UzgSx/zKEslK+87ttfkD3CL7GpYxAobewiGohpTX1cUTGtt89p6ZESx0QxUtaLih
N4kbMbrEy9I9Lt6LAi3ScHRx11JmcV5rJSVLWKslFHBaD3p9NVVeJg2BYQpWpYDw
RKu3Zc9zJgsVs7nlLz4QhNvzqN0sTAm1W6dTdn8ENxZgnRODiKKUSqvnBgmdwjW1
ENs/Ob3zHDEyOMQ8wz3sFFemwOZUEMjsYVT7DGxYo2SuDMkDtKbp+uZW+J6Rwixe
GAU2b26hLcAlhh3nW8DhhXB/OqDMZPRVe+e2YaSdDQhM68bphv33Uugzc8NqFAFi
pMmkEa5Qu/tuPMwuUWc/30X69eEi8to3Ghz6STrwF8SfoXDimEXwe2ymAJud8qC+
UtxfMlgMxaBaRjiHSyA4dCQR6CxS+wmL0B+l97YiKnzogakOvaXG+A2FLpasgjf2
0ryyxbx/UvefEgzKyzZlGZliYGWPK40noASksXnoByCvfPrHEAA9cbGyZQgyd0UU
EKGQxVKroEoemtSdkp7md4dpalTfO7olGp5o6zrF7+6uCgLnlgRt2wojYGEiy0I7
/7oWnlPdBnn988pi3dSD+ABPPHbMmPqmTl3zBUqQp6yCgVYaREXWkXoj0JWGOx1w
P1/0o6Y+dTaDzxIDUuGEBEL2VdmUaJsxA/yDfghjazSBc+sfMru2CloAYl16QW00
06rAcMieREycCfE/aydHkRhC32bh4aN5JUVeW3uouo8Nnd/uAc+SolJGIVkZvBym
2r0U10YuPamH8yvF0HNYiVhRg5za2ECPctBrFkf6gAFln2TqRmD/6Z9+/hLLlmSp
nOZ11SuNeoiIr+WWA3UwiaqiSui6bVl8UEZqv19zAvGQei+YysFTijhBo5VxrU7p
eL334SOPO/8PNptqMGKYht/H2u9Xda9oWUXP1tYn6ycJPIRFdF8Yk4IrpP4OQDMT
D1r4zG5fCGG3Qahua0QaFZWMvT/LMzcva9KCInNoswkQWGGOsQ0G5xsOLtT0BLWV
p68tIuIfjwB/MUTVv0frqcjccLKKLIg5BVgg+M8ne0BCXSXkZX6Yf/Y6y6N6ybBB
yOoG3oqic0beuX2HhIGJRCPsJcfd60b1Th+xnjUNj1N49RasIgpT1iw2IyV+AtCv
L2dt4O9t/lHhYO+lxYJm+0WGkqGBvllU2JDcXKyzjAiQGML8ssYDQsznSsb+Lzf7
qAmqgoZu7ENQ2EANKqgDIldFJwtgaa8pM99i/K00zYSuHPf0yd6YFOP6BnPV6PgA
F3B1pYrkOWPDZ8VMqjBozGcRyaY3Bq77TZtclc+mn0xQ3ZocTm1THRkb9OURSv25
+jhvv+j/FZUbprBN2iUYV5IeIQGxrcmbH2oLPpC+6dzH/BH2XOMUkYcMH9Zj039t
pWQn1DsnCdBy6BZWiBH8rzA27Nn0lGLhQQc8VkoBEOoCaqBTSpy6VhWhZgfFilk9
WfTRLBXs+EvNlrDOpGg2SzKICocQTRj0bmSvsWpkoJk5UPFlnmskrlzfCFr+tGV5
fdBSZCQXwNqx6IJq6KX5nP+ea6E/4AmVSw/StF+hBvoYrCwQf5fHGTEOsdJEi/Nu
qC7I+17i9rS9D03Fzg2pwB5ZvT8MsuyEUYmfyOZRJBvIoKqx8amR8UabaAqgHLS1
54zemjDR4Q2WvcvGYx94axyScm6Eu2yNoo8GQRVGluAgEyB0t8Eu8begbqYl5tby
l0hs30WvPK67y0Q/MckNx+mAcdRFH8IWUTNbveeWwZ6owKAuHZcLN05qmJgbwE9l
v1SBQJTH/eHYlZltyZ9W5czvIzYUomQCekntQxrjzJUAd3Jmxa+Rk6/DKvXG44jt
WO5lwoZv1E9zjNNuL2VGwmOmyBYQITR7p5nS/loUT6Wg8Df/4MSZDVab+4WDZC9T
BauyJGRiwWnyHO0durqeXgicqSXdPQiOC4JudFI7NbatdFjJtkkMMg/FhTUW9p6R
SWH6BHZKvYw0d0sPYp0SU5zUQCBf6BJLM47k3thAx1g6P/PhK/6qFEZ9Eflk1Xu+
WFsYqafoxwU2gau2ZT4HP6Oxgh5MPTZgycz1DVgas8afrn09VIC3kF3WEwGGwJce
aObgoEzlpOkgJ+GSmCoWTtxbzxh7N9zbkF1Uxpi6G6cTMZvishjttVG2IxGBAf12
L6K9mNwRBs0UWPGDkynW8KLN/dV7+CpxDGVYqua2yS+odHcCICia0QAhTS6T1zYM
VMb4HAZmBb/VIRcOyMtVvIiBZK1uaD6o3dA5Z9dcG8lLmT8TWNTx5zStap3InxxX
9BTRym9wYfpxQmt4udXfgfB4M4j57HcMUFzWG5ZYBALb+lhDjsCkUsMjK4q1VpAc
TfWHq23mCtpDcczM+XZ1Som8HyNmXdgeNUeYoVPQ0lS1l2DIASRCDwo0i0FX3cPo
PTAe6ueL3+fIrDtr5QwbhiOi7OuL8CRVaezZXxfrT2T9+1VfpheLo4xXmS0FqUHc
hUnx71G2CNWeiClXR+Bx3avJnhsVDRzO//SSGKLYweum06npHMlVCJ1Qz0ERo/Vl
5v2p/QErXFG2djoFQEUr5i7PLmusz/KRKRngbo7C9DjjX3C2Z6G4Yb8E0FKUsqCL
FABtwA8go1oZQDpDbqzmzq0ohwh1a08AmSowL07YCUuzywWX9ItFHAOw9Gg3h/a8
Sfn7fytsIQvgYo75SeS8giFYdnWnpu1yrYuJRQu5i6lMKURTCl1pepVLb/xKbyIf
TUf7E18DzXzX1XRMbNZeOtTB4w/2W1KVwLV7WuHn/CzU4JHDeY7HSm+d/10+mgf+
Kz3M2NgW2rCWEFvJqEuD2WdoxQrcVUj+/uLaJ3cPT3AkL4soUaqXQ+WEXtnki2YT
s1nT76IVkr06GlbdwjuBB5WyLygwZfoJpFRPFMMoxi7KXybKm4s6zl4XSUkoMShd
4Lx5cDjHFS+rdLi6gXcTjAZz0LnV5SplTIHsTNsX7oIJlHAjRker1yalBKnQxFE0
s8E1ZV4PvGowEEusZHhBbcPa6/3F7au26LSwAUIV1K1VrCwCpeLBS5jT58TjfMh2
mqOhwOjA4RB26NYTEef+AFvA8ifsv9hV5hD/HIiUY/q9i23NdQ6ypFPw6Ysxmv/V
UdBzVr1Y6CdOi5YlKYZGIriL2JgOsEhb3I0sLLDZAykyNcYTzNJUfk0oMgR2ElCu
/EyE6Kq2pYY0yJ+7QpkkbGy1lXLBmZx2dGRC2yFGbLsOLuzyM2e3CiPTX4tlpH2E
6HfOVXqTvddhhjEYr3ulX2pcxaCbbXmwoqzjNl3ml0c8NIoW1Ibv3nMbOSl5Ta1X
kxnPpsC/lqNL4tvwFQmkR9/t1kF7N5uz3PnVWVge0gUwRCKUsHU7iB27BHaqjqyH
rfZAtwGgDXfcf8hjJYim+AH40KiHhpAEh3cOD+oyYN+vIJlO8SQEZQmxgNO7eDdP
cx4XcPAlbF+ZEVNmVs3tugLRNxPWWUOesKnr+WaRJASt/rHXvi+2KqTjcn3JVAJg
iJUFaYzWGQJhO4lJZKPIWpx822l+SI2OV+Lnpc1MshlMCV1sWjjwM6tgsXFLjY/l
6n034qTECX6E7g21iQLMMvEaK6DKovJd/MzLJ6xIo6D6fKOAWbXD3aV42wOjuWH+
CjzaQHUEQBJP0C6Qt6SuegxL+/IyLchGuwsnvMMueLEvLYeZuu5W9Atd7x4UhL+f
2jnNTk3n+1RMfySCPpEk4n1CA3IhFnHjvvtj573XxOq20St21fKsP8drphem7zxz
mp0HYwH6E4tg4GPamBDSAZVnzBoAo00QhSpV5vGI6ImU+xsmMNUmwQf21VOqs2mB
cZZoBHMZcEvNwVOs3na5YlXAEgK4S1R+whv4oT5/SEkrZal5N6ASSWLlGVn/7Qn4
P3u1hhjTXR0b+J2C8NdeNiZGD2eVBc2XGLWkHRYmnN8f/F2FZPekPnoBuE+QiDNc
PMfQreuQzN4JbTIsobUW8wvK3tXlnR+5uNa0Ze5M+cndtfrrNV1tYtlnxufyjTwE
45e/qvZZBc5YP2hVQTOq+rWep3I3pEd9VhUsZCp1QwSB2DSbWB82MZoMCw1glcl9
0tuF3DnwG+NdTpLht+IsJczvmFOe9DpmKcVDNYjkktIXDnCOHwnxcC7wYOqDdjaP
H5xEwA96PTCLhyh0WRlc5++RNnXRW9osbIpZrsPrLCoW0UU/jHvJAlqK4BzT43Rs
sbuQdR7i6WhbitnXA9ntCJXAFl8jtmCctW6AwTvohmlEpnydX1kvc34tIxU2vxwm
Des460i6/wgJBv0ZgrYE+2ODq/HigqxiTd2hJt4vpHxzxbXB5nCZqpr0W6SCUCNZ
SnCLc5K3TK9+nckKQFwGxOjzAXRRXKqSn76p3HTw6un/lSiThsqkll2zdgXzGH9n
CSZyxcj/p7chzKc4om22GG47KHvv2Ch6orgREDxrdyOOF8rP9cYbMJ0C0YLZErjz
qtvqgc72iISfzQfMZT+lNOr6b6lWlEH/9qaPEKv9UJqQP61cM2IMZR7h42QeMQ+V
BPk+jlkhDqAjh0mFwa2hAHRRTrfIglzHy8C7OZKke44iEoYEUq2QlDa/MkVyGY4L
uvaT4gMvgm80JB6FLbCWwPcSPUWjMuSXF8Y17JIN7TeGE+b+aeNsQyijX4qbEVbh
zGQw7QF0E4LTNQBgmjds74uEQPUDbILWBy+nrVY4RwK1OmcBWpgiiCQU59VONN7c
OcdpUcEr6rqjhRS0J+IPtMkcto8Q/ri6ZlCo8PL+w3KZo27Kc575o2SOpWDkElHf
VexYPTT+J8mZaLC9KTp0TDOFRuDNUE/FLZBvVhNIgRYXPdrEWaRsatUyfQz9A/04
RZE31FOeed6rH/f3DqLdq8H9bH5daW6e4uy2oWEVlET1FNZl2l5zDjfRZPMth8Aj
VHLTQ3O9PSMp1TutoluPFfgj3/TXNoFfQa8u7j5YWM0Mv5w73Zm4pzNDYeLD7u8A
n+RyvmHK+BBH6808Ct3hZgJAHbpyfIkbdg7ZsFThVDP9zXZhX5aXjWjn3igaTHfo
b7eMVk2WpScceiWmBUP//IvVFjcy3kUy46/pipxj9+h/A8wiZpqA5FyFFE00nNig
vTFMlkWu4i1GT6AfqHbSfbojFBoTTLemQyLPZM0uwh2s28btdCJLCidWDlV2yGcI
PhVpIVKTkcIXFThLURxMHDsMhHSvGtHVq6MYFs70HWpayj+DiVLB6/qZNZs0YBi+
ydp3JJAYWLbCK0Vebzhyj/nAoQVsGy7G1aVEjn8jpObgzjeoTzPtfgki1B3jAcX5
0MiTupEhC/Td5vJoNPahNavTqxA18hFTfiE9xztd3Q+WtDt5Kd/1ABAWJN9+arMm
vB7loXo+4c5KlAWZz/EiObYA9D34I+wVIpXLSC9OhzLNgRfYkinMbQpUURjD4oFE
utzrJQW6N1anjkm1Ihi8As817j5TSNSLPFvhG4JdKGrX4eRpwU6hXyPLD5HUFr+4
uiv2UFbMenkecrmI8yYDsnTN1DiMISnhuQdO6Ft6WYpyoKHv7gB06/AkZha6zDGF
ale94eOVpmbJtvoXZZ51wjfrUvqnceg1i93/hQNBu5pTRrseW+0FBruESVTUAQjw
yJKZeXEkngJvyjh0oH3Gv3HMsLKKLhHW/Z/ymbnCNTiPmTnPd3q5QngPG3Jw7JiN
BRuOJkTF0JB5b4G//qYHHhhglqjlW13J+xSSiD66gFmKtEsbRaVTZaymLXqP6BXe
8gzQzYfiI5uHojuLwlQ6n7QZwHN8gcL9lQxNfkTASceq7nThttq6uvyVD/skxnGM
9mJyty1WpyvqhcoJSiaQpeB/aPOoIiMo88o9uCPO2apMldx5fYXJQorNuUizEq5N
KeIhmAl7DtGoSZ6NcETqUwKzk0yLArHz9EB1WJlNRrdYRbFXAL66it3W48LiJP8h
K0VcuIRmJvUp+F6lBEtNvd+S2KN1uXaCYhO57i568zQV2vh4rshavJq5hL0F5ALY
fwmzsZ2x0bvZG+rkdFJ6NP8viqgM5vPCmyJ1Bvzt1ThchvYP4BwTJztjkZOWifCp
dVy2kQX8T+YVkG16x5ZAVbPyjEsAA2GDQWcf2kuIPE3XbpsRbo3xUFTnK6BNocCB
OrLKyVzwgLlGevi+NFd0z3zKjdEFfiE12sUvKChcB3tJkXc8ciHEdErtaErjvwmn
d+MJF+7sbJWOcHFsQciioILhwRrrldxMAgioLaOPmQg21rJvwvFf8P6IniLkuIZe
5xVRQTCMoN+/PNs+ABMzWNbfohk4E+zlLvhdfhT6wXWhhRhvMzEQNsoJpPGk1+cv
LNeWk/DptXlmYoWDZOI6T/twrE4rIwrM6+IwidTsh50LxElsTqh1gYM2mZt3tqZJ
JF/88Tilip6IP0+BrXl9GNyOI9TqYy23igyY37dz5VoymhAoo/TtKbFEe3oOvaSo
SEWN1JLohYdPbOZ/ueUcg6eOq7Tzfw2wcjS1fzD84Mq6F3FDTPbVSPhdS1pd3cdg
1yArFN03dGTWRicDYLc2/CJpeC4lmaEFvfDrWK6zuKDQUvVt9rFoob9GtFZuXUaH
hoaWq7tNrpirQN+BtZwfUsEFMA5eoO74CRFzKvYPkk0l6J62TPLb2BTexCiOqx7M
uthIr8/vZNjQaRY0DOmIIf6ma10/rQmzlk163n9Nb9VFjqotEQ3nbmTh2CTwY3kr
ydL9sLV+qruanao8QDb8Jwl1MFn/q3D3Dw2k51Hiyk0QhcnIMjPmrtibW0255iMG
8vU3M/vPTZaIT6ERMXJuIdRF2OY5LhLEigFPlKlXYyQWaSDO2wHcYDA/hHUfRkG1
BXn+6rRjh/NFuL/HK/HuFB0gtmoMSytLl6r7kny6zSIe4nQ5XxajfL6ZLf7iuFQi
uNQYMXlaVbloeGOFP4mIoMz+UJxcCCbMrCjOTcuoVdy4gMY7hqvAozS0AJH/8l+T
43jKz8xaXQQ8RkLqP2agcfEX5spy20A5n5H3h2ZhN0hbrzPNMdADEu/JUBYpkWrw
bApMrioBqlSbKsTX9cDh8pcumWBixtkcYYNoMpQ5BQftjgcEQu4EdGdrALTPhH61
lXnVLYe0RulLyZQ5GOpwWzqiX1Lvi5Oz/GrJ6CRdl8YclTplEsGvW7FV31VSXVTf
32W6WV7mGeyIxK5KoVvGk8dQNd5n+rv/B131GxTSMhZRB0uc1RRgtLY2pMVfmtE8
4xu4g9RNBBR+xJiH4IBjgeM73CcHtd9z1PtDNmGUFNPv9ALJpaVbgMdkWL0mPCIA
z3NQN3gq2V+8lIBPiyCeGwB7bpqXzfHjkDGSvG29oCCnNKqoOvwhEQdybhUzR8RM
WvByZEJ05v8yNr0m0WY7mpOpv/xtEKDY9OBL105HijmY4cc7dLIpG4MRw0kOL/v6
G9qpQHursdxfgEvMclDUP+njpI/D4sQ0SXjPaOubBH15aBSOzAfn73diglxXLCOz
du6+AmVW4lfsQ9W2ijQVpjvUGP40dYMamZdVeciFWNB+U+hcLTndQKv6AR0cKbas
XbPny3xxGykAj12hhqzSrZ3OLdna0189mj/7IcSdKqxDvRQ04Ye1rZdy17ESkIbR
b+n+AG+wer7rENf+VKsp6H9gjM8IWE/6qcO/LxzCsN8pwqRvU6YShWd6p/oVaeo3
G0BM0j2o3CSbZGzCrEbGFTLZr5G5MyqhzOThazaIsWY/0h1HHPGe3TQRzSVFHaJn
6euCX+fN81MbufMc517SmEgeE2Qu1UgMT75DDMxVr8gS/OtAvvYLIyBOQXMl6mef
kaA6U+BLnATh+KQdU9dJ2FWlt6kZ4OZkTaKUJI9xW8Di7G7DKlgfzjPlZAQadHXx
HmyXEPYGMZIwh64XLzA1plx8UNe7/SPsSVz06HFhIHTuwqvZxcKROuP/QlfXKURf
g6RWebarBV8x7Zuw/Vl/hnBjPHswUSd54HDZjYCsOSR1xdHJq34wWsD1VHLnBKvO
uKSCgzPAg6NY8+Vmf4oDvyWSTcYdyqZBfv/OUsh/NPmaOG1kbMm6EFhLDtd+sMcG
EXXLd6bQc1Ci9VLPFZagql/0/VGFlW41AONkgiBC2pIB/C1PtI/2szFMNPIGsxZW
6UcOf95r/1D90A7qEGlDlpKTOsQP21cZd2p/kzYFvNhGJ4GScdSvw58UggmmPnbD
vOrRzXgZOItGpGpZsL+iLf4WSlo95WQSjdXEovoLqIhTrA88cWT3NkWkQieA8D+w
VjHyTNQJC9CLyKw3f1XPr7X3OfSeBCvotsSWptqZ1kf+WeW/nI30yUXBcUCPRbTJ
vMU/mIZyt2zvqPjb5LIyBsmJp71Av9euiAM0QRZLd/BB7hAlsV05Ba5I4boQphze
v6EifpWBdH1sytx9tDSxPmqTmQ/u2un6G9jY1Lha274xr13KTLZZAvoWKRNiC6vn
WlzxHDiseuHW/1mN/XSuEgWhic8T7m0FQp102bx/pr2wjOrIZlVtyajiFgx5LhP0
Ya6lD6ermBh0cgc8a/1MOwhMaAOk55qK23YvTjfAJ2gc1Sd3WMdu25EVzx5Ue+vi
EpUPFKmAsSSPP2rXNSZMy9MH54/l0whpyEG4Glna3A4DFoWMqrwAWT03rhfqLNTy
ZwRppA5pUQhHlXS95qlh4F2xIYsKM2ERZZnO4WPF8oc6mOAPZ4DptPR1TgTUyHGH
DtcAVHbP3IIJM9W3l7DltjcbCBIRRMUhjihOuDed1aeQHZLmFhSyfVZ/AWCVmnEZ
ZazZU1iLN/Bmbckv/7aRq/jLJfdPJH21IlgtNXanhUd1HfyJvSYhoyx6OAeqrK6Y
+7vCXe/vIY29X+uaoa3RuwVolmzK8g433D42UamGd40hvhSUA3CNBib3lhu/Efsf
nLTXJpnv4Qtv4xi/oMO/TB+y09+/mq95C5MP2boFLyRlblBT2sj7zsWuniMhSBTg
rO6zZGuzaxXo5Z4nyvSblYSyFJhDbeyPEghwIIYCAu+kCY5HMyk1DD8w0iWzFYao
qstuvSqwcRstvPPbnhXPJYm80muKB3lrkwT5bgn4pBxOkzccCdMjAiqLHGrErW+w
Y0Q1iuExr4HajDk7E56XgBvzbw/HdmwP+CDkk+zkHkBD0SPce1qC9F72gvBa8vap
QGcVS8pjOTl+GQoj1rKSu6LTHObsKn1Bx5r1edZZiqPb6ytUvHj1RcuUnWFih7CV
xaSd2+oTIteaRiXO9hV66YB1jYXwjnw5pvgg3xy+XFvqt0bl0CTOIBbOxH1MPrM2
RGbyuVLMhXbEBvj804p2J0GnOKQGv0iRW3Nr/rFaKKw0m+rXZHnsN9J5j5V930o6
7UJ6xxSLq5rjJHyySNflLJ3XJsB4J7OGOrSdEiZVlv9tEOn0CL3NRSa31bqbyQZQ
0dTBcWbmt77BqCzfe4HAQ7JhgmBUoPzLJGGEVYuZBnDwrZsr8wx640QCZFSYq+x9
Pr6H57L8hk3IsZ+nXMldB7Cuf0puM1R0JCAL9/Tj7oE9+mf+UBi+yHBWqX5w5Y/b
jTXe3hdNlrg5cHQh0O3t7iDgbIihiHqeBb5WkFZV3apxhs/BYO7G6R9kfqTrcvxF
h7lZepO5Kcj4G+QyEssycmu8JxnafZa5O/ILQkaFGmSBhJ2E3cv+8PA9FXMAD2Mr
H4GboFOnzpmmhYiPe0N1oMwaH2smfAG/R3XLBGAh5eD+EMiYawcdWU5mCqV9PKJJ
fj/+gmJ+WThPnzpMshC+dvphTwzrnC1TtapWE/+Up8TTV6WQ/b795fE8txKfNM9p
rfIXxkAWbjN7tEfbWxW5LxHLEJE0IhrLvjzYUxFF/eNF0narqu2la1hgTY4N85ec
Cp1dKZAD+Qsdyrxnd6dfSdTiYL0S8K8FdDIeKXGVULFHln3mTVzD8hLrPJM5ILkP
99vqec0jrxSqhqAt0dzc7vI2cT+X0olrLwaMvmqMcw7gn2LDkXvjeoXgzDgCjwSB
VWbnHzdyimBVQm33kBtDRLQ3xlLC4fuViJ5FYo0ZbHELDughtIn2URbyaVlR7dld
P1fQM9860V/SSQlrK3MtZTUugmix+o7mwq/Otd+SGh1gc94BFD+bV5zuTwR4g+6N
foJe1juonNCoACeU4BMbFkv2zKb9RlzRmCMar2nP7sSQpqpMHPdPr8Mbsb61upiB
Xu+NVvXxTtrtSf2QcEqO/n0TPvz0sP8JjIfzDTp/429ca0z6CXEPJ1MDgEK6NwCe
7XnEzlhDBrm2vGwa9iWYYuX8LPEqWr1i1KVJnMAjb8U7y9hnIb54kW7Q6wNF1xOR
zPxnhWwlXEwXaA/ohEhpqkzrAQeHH/HOJDlLGfmWPzISCwr7JSa9cM3+e8JYm6PS
dg4QyS48jOklqo1BcrUo5k5iiCjssTykUnW1cmSOlVgSyhLPA8cdDdwrMPrFjMxB
EUE9rtshaBxZhmEFoqGuFnDTqBQ6afhGkwHxf94ID3pISnzDQiScubkwoexsrRpH
ciSGCDasVuczU/BjwyJdtK7toupZT9y+fz/9SYw6sR+7dLw+xq2uGDz5eCflV3Mr
bJboPgPBeZdWh/zzbOBYYBe7nnsJvjDXOXG8l0zpsInX4Sji4+FHVCzBuPyvnD+k
Aq5Ke2SlptRQGnyoEQIncafAIgYpVCv6Fdp/q5iZvToFlrBiM5dXapnS50TOh/nq
Lxh5pfQBWb+UFIUk7uO43dV4wzt06BEYs1wiiMcFXe9xEDE6owAFQ3KhSkWTjTJi
WDXz/Ae10TO6vF9xRXAud/PajAn0O9XSfUPnBTZGzODJnOOSwQGtXbyhYSQXg0gD
SmkMe6UX2z6dEDfudK2g7A6lanc8vm9jB4/PtC6Qu3PwzZO0QBQB0WUra8qH7k39
0rudg2IBk+jsXhtKA03SHm3zBsxrdfllzkLafuBJ/AV9az+N0MK2sCM3weju6mZk
ZbTBBQDciI1eRveSTJGdQY4VAXycp9BVJa6FLVQeRpOaSomYfmmNmHsw0h3Zpi9g
PNImYRSXoLcJIOF5uvxBpMddgP2QNxISO4pYo2PxXSFFOcjVLlSOeszqwajtRIoi
Zw9ebgeuOFDoX7mHPiQA7XoliJtgV+LwlKJZvHRp6Dw9XfLpkDNlu2S7jfwc5Vfh
xV5GEpfmmu1NLbFd0/92YR3Kh1zZn07Ruc0kGOcpLsDeL0bU92m0T7kLyeGVPQLP
hbgBqJq1nD9hX4lS753A3kUzHhHJ6x08CMKc5LwSLijRNZK5kZ40VuDeU4pd7L5t
IUFSRt50FAdOn1XEFpkq6zGiXtgfj3QftLgf1AYhe9wQOpgJO4FmjIdzgVU8R21c
6jGURrvRbcshfjgW/Y4oFz5/jU2OdvChX+NQEPEoZTbPnwNU8bnU4YnZ6QT06cAK
qeKXTnQ1fYploBBK8NDzLnq6FkjLLoeoB9Fs0gz7Jl7S7kf9cKpoQyMgNsIoKieH
1KaFzfeUcHZz65241yLH12Hg6hnD9UnaBdW97MSI+Di8QvhDZqwkUZlSWEAJbvgr
YRfbV+0DzfxP3NX3XVHNAXq7bQ6RXEVp8/IuJX3TFuxAqXlfjW5vhxKJpD79gxzi
KEdo6tr78t1Jj3ycmdMlCL6tCh0hFt4iuMF+NLVDr9xKWnFjv9gE8pg8MQy6hOAA
2fiNLC5FC7LIx46GmQS/LHqlk/yVKXY3qpUeyU4fYnYIMOwJu0RlxOP+qSD60VNI
IJdwMi4Nv/rYvAr7Pol7HMu4M8C3lJansks8HF7N0USUjRfFIU5Lw45JnaMShFn0
fIKog+TO+Vil4WTbLKck9gMbj2kYIPHOJnR46M1WdOQX9ffLBjRllcvecCmUTSTv
Ys19samCMrMoXJGmTQxwaK9uHn5SdJhiJBcINhpFAsRuAlmt5YM7uJAT8rQm7Vyn
4C7IJXEXtBHZnZ2zuI+P7WG8ok88JEkoCS0mV/SX23ZFTqlKGYZX1CPtrsELyIKm
PYy8Hu8ybO+6tq+2iqgghEuDkRoffHZ1GDAZWpe3gq7oQtrmhpA+wz+gH6Jx7PN3
TT/wL16PL6PsMs7cF67HkhdAO4IXhzAhDSk0E0Nw8IA1BjdKDwFRTYh2VkIj6npZ
ayeqlC/Pg3Gz3sIQOjG26JX/phL8xeeoF5XusSd9b9L1VpffOyFW0RlYR/PY1Tyl
eP2fQLO1snmiPHCF7hnmiTtYmq2qWN4KILrd08x0sLT8cgf4tWUOTPMX5X7dr3Mh
UMtEdcTFC55YjbqX2FUWNo9oYcs+VYfhxyZi9waGNufotpx5A1pi3rNODeR2y+SV
18BvG019fq5JvUIBmnHcHIwpsnbwNnZ9J71N/mK6DB2IZO8xgf7JsbV1lFwBvONV
MMGQm4QAtm4ZDDAzTUvw+1vodFRg4a+o9qV7N0Yjkq3Y8y0IB7gOeJEgpuasTmZt
NqCqOhVLFFSTJH8C3Swy/NkiKMF86xD+NO8/XpWcDiiUa/7KoW6TbF+eQyHdjTAO
Fdn/IlhffS4LlyQX3CMlbHXPVcuYSChjYtJGYLgIFTpcGMg71hBCPnTDMAEIyJ6+
zCvXOlK+N35fK9J3G+mJtvQU1yLIma7uh76kYa0n6GOYpRUWR1l0zBA4sp84LMNL
r2VQ+gKm9PHHE2z1/5Que/p0oHSCxrcN+Rcc/N+uU0dc6lx19BewWCoNzFnx7RkE
MRGB6a/xL6KD6aGwtonHb3sk94VtuGtif5hFN8XqvywQ8QBzpgG/NOFT0E/uCOUr
HgwuUPxn51IjlIQIbxUqIXEhMW+SyHuZ8PyVDa9p2j4TmDFx02jCYFoAfnJDuK3Q
FjyurXfYZwbmohawIzMedmeiu+RCGeWAVLi3e5M2x1bqg3+5nOWPOowccC4LmWN1
L+BCfZHo5lbcCaX+26JSllrtg4y4xeBFQI2SLe7F8NYgtBfjebnZfHCsExFf647j
I64RE8XfWQofFghcYxyLUASePcZrzgwCn6HhFOi77E/MKCFAgAEG03azEWv7kemt
2wB0VogI9ctBk8gViiIEC6BsA48DUqQEiIbaGc6McNPwtIOjnnvPy2rdkaHmlJVi
r6ZCvUVcI5kk1MYTtFWZPAmtUrwtGzuGosTUDoyQrh+kkGSL0s2D4YEYMeXkhhqr
TIkr1ZsJqBr/wPFcuERTE+GR1q01fQU2iZhCXHlO8NYkvEuBf4w6T6lIMFq716Za
KJ+NbeyJAojJ8GN9MVoFhgl2BfJokiEXlYMj5ljg2XxGQaRY4/y8RJahvHu6Oip3
5y3kXNgOgDEhNG7fZAbquNBPXbAPWIU5/drNePCZnkFwnpNjd/osGXcyzZTIpdec
t1XVKtgwr3sOyb5dnosz9xU07yuEfZpvVeuzDPGm0dOS3mXQxydIhiXLvKg2vbRL
+g7CTv//9wxYEDfu5mPIj8N4Y8KOrEfXOnmy1nZoFKyWcz+/JPXizr7f+ozXCa9x
04CeZgkzuMPAzuSr8+1lMsDrLDXtuOgIqUU0kzNFPPZHWvX/kWlHeNfNTykltVbU
ON3PvxF9wUS8cXc3GAS8P8yetmAmqJfx1UGW0JGbiU0vZfT1KVUBqds4iK+AHHii
D3/G8jfTobmNqwzG3Cd4yJ5uGEEcpSpE9Z4Grzv24jOetIok34lQo8ll5LOU6Usg
VZdG1/M5Uknpy8qGKSE2zYz9S5H79kVfmts9BRxBMPwEzoKVJtDxv5pEwyLNSknv
u/CA1ZsecH0fkwqQrTer1RjF6w/5EkJEV3r3oaGGLtzdQqgpGyFNmZPrn/9sx8sP
cS9qJ7dHCiSJM/2CZRgVVusJnm+dczb/+2wBMO3sTex2e3KuSJPIPoINBEwb1y8b
r4rW8oAGVIAAUw7PiUAsWI/Iji6UzNCJ6lpcf3xIrfhe5DTovJsTFt1Ui1vFqvMi
9V8TiTv8ANhZm9wR7hDrhDEp61RS+bTsrWZvk7a7YheVqLrzcofBkzJws93bVeCj
P0o9+FGqnVwr7FdLE4BS+Lt/zsODOz/+xq5O14zJCI4y2GNg8DqqnwZutQy9PFdK
a7Gls/hApNDCyK/COnQQg0USANboJB3jpWYhUzB6erJeIGKzqG6eu97gWx8eusVt
pJ3L/tZhiruAfS7yj8GQ2dsLJBe2M4m8eiZFbiu0WYvH3u2NSxobUv4efShB59Nf
TkqEm9flAvCz8vzDU63TQUpXk2nz6ukA7w1K/9BCugj/6i1CIysxfxTm0PIh1Kop
oKpKpVgoGGaaonL3WoxWiOlp7lryjoOi3v5AfmBxwnOFgGsnQc6qS6Bp2R3OLnBG
70BpsLijKW97i4opQqQNb6mAfeOMo8UJvR/Y6RWteaK9jxNf30vGMNYco4X7R+/k
auOuHkrmMVPES7Zu6DKjimjU6dEEfZmicGKVV0jq/VvQgDgaPe12fxaKIFAKV7m/
LbY31ywmEK5BNPx+8RuyXpQl2iMa3swfeUjkuDcVJgce1ggEvNr/4DWrLOfseDBX
NgxhChxgxTnzbu3wep94tOj08QQW/NmVWfVVET4Mco31ElvvK7J6LVOwJny0RNon
RxRfC7s01aQ1gfVb56MsmebczDkpP2hZc7v/kjivFIHOGDUD+JNiz1fS4J6Y4cKw
rUu6Mob9D8i7TC/GgLtPmGThHWr81OPJEmrYa99lKcJKsiH1mNyhW+aAaJpsWVEt
CYbcVJqowzJ+bMNd4myxxYEoe5xrvrX4/5ywjMRWyyqrwugwHe4K/5+wxeaeCPnG
2VUNR+WtMSXy3/iFiHaJpMBn3N13x2sCgWKGnV0/wMJG5O/O14f1nW9BaIi5N14+
Smt63LV5kxbx7O/sxxlcZQetu8Td/iwFgNlvLFxgmIPNlStPFOrBV47XJJdFjnzu
oDebSQ70+7zDBbAo8DwPARot5ajdyt1ozF9hQfmuEvhNMQy0zZl94mMO+PwnawoR
rGUN84hfr2Ik3Sm1YXT2NXCLsE0/dANycFUvwjyMFztEC8femE31K1gTrGuR2myL
uN7IfkpOJApTFhNvfOVEJDY8LlrK5xKg78vRBYDhX9GVKMhAyAsiFIHFvwvNH39k
DADMvUGlCry1f7zcrWfk1AZvOY+RNUeeiYNZqOPkoBFuIvsCPWviXq+0gZI3W8dJ
UlNNIVZwxnKR1yO3+18RzK5jLL6HeddjMKS8LKn2wqmHtToR+2JabNkIUcHWaZrM
GVynrD1wbsjisiCMXU2iAECy7vOU4y/TiqtQLIDTmxjdGlENJkP8xoav3iiKCP8p
+c/jowawSZbP6N7p2bBshZ4QM7CKbBT6823wM6lfuFUvul8zO1+QTBNknhqK/a1R
wAQSkaFVO3mODJnWZ8G13IJVOmWvk24RArjc2IGac8s2agv9ER4EvdgUHdFr9GW6
sIYpzFQSw/KiAZChu7KLEvBB4G8RdyCWVwtiGeqr7VhzYQ9gzBvXNV7myrUETXRp
4uj3hHJdO+CSRjFvFGACxajBXnfA7MKcsgqEoQ7HPibDZ/8R2ElmxK6rp6YIjcDS
PLPU0Fq6sOT8ia3y3YadLLIZ9IgZiRrjPC4+5FGDE1T/R1Onh0bgzUxucelUKWtM
QNK8XLPnKaVB/oeyhvcF7LSUxKwdMr0PfiA16XLQ98u/wMRghRWH9+WolFn4VNq6
JhX5z1n0lVP1scUETB73YBBM6/SYD32cUTLvnYoXKKDwMNE8XLlyYWoTNjjvrDHI
QCtkU3zTWf9LaKlqn+lL1PthfeMN8uVBSW+fGt+0N+11CY/o90RACssRnQLIMLLN
ew3a1koKBVELaJtxNJDF4LFxMSZ8N5lel8c4PEjfcVX+af5+55P4KKegsJ2Ni28E
TB/ew/rZFWeun/AhprLM20T/UGKJZtuw6DbCnP0F8w7EatfSUTWJIhb7dlPtzu8D
Xcc1yqt1Govab6Wlb7LXIx9d6FJiBhhjRsxXhc4wUXrroXuwjRWUUbmFAvjDW+Bf
uVjuGNn7svfxLXA06BSA+2j0aOuZz6jYhCR0as/OXK/2e805gegWqqYX3Bd9B9D6
RVSwfViE8o6mQjNRMj4f6x5BcrKJ01F06L4sCwROXIUNIbiZ0qQdY7dMbNlc3Dp2
6+vyDEjqEnjPxki233zemCMuCeodH7GrEbi0j/5r2bQXbbfySESn8BvLMtHixafP
PV9g/bF17Rx1vlW2YHONTvL6dtSMv6D0HUxNsq7a9OSYU8OIbbqNReWaC3N+bIWB
WWyAFb0mmd/QAUnyfLVq5LYQwp1J3aSAkCV+Erysm4med5Jb6jXedeJPdVHNEEb+
v/0OSrWM1SdplIFd/u0IN5aI3qUgymn/CAX2D7yaAeHXQnC19BsOMfqJpgdIGA5P
jtxmiXyBMMxcCddUmPnpEwcjDPkTSD8edeULjhCXw8hHcNnBedqejGzM8Qz4tdMf
TZEutQmVMKS+RSe8qGI7EL6OnmH9sfiid1hb2xWqV8dbrYMACr0oy7xWN62RzrCT
jwhHXuvWuXxK6GHjeOxZAq7Igctm0fS/54Xnvv+LJTfi11WfJWOjhepsRCcovi8O
Yys1ar/NnJir4G39FMQx5uj/VmV/GSyhxNZgH6ap59SDGx2Qbmyd/EE7M+XwgXd7
LNJhXjnj+VRHc+FAw+6kTpjSTbEcEpJvUp+XeVaVYHVppf0PtwbXzy7Un6SEm4B+
OxsOW0/y66w710a7Y+wsuhgBzoXkf4BxIEtoa+ghjQY11vJmqfeeQBo3e7F6YBST
J4rO81sg9Kets4MeqiOQDqBTWmrcHj3iVsT2wQDQCGhWVYdac2pxCfI6MY6ouuUJ
ScGgaILxN8AwAqKZNItao9/q/kvrLfnZYaEc8hpBdv3P+VrCNHuUwR5eXOgVu/qs
aEmWsZgkfOS76IDC7keD4YkAVPorDBxEDEAuEvpgTMwfBx9U7Zcl3yhNVj8lcJDi
sir2AWUJvDR/a9NsffGJ/RpGfw4gPLLmkqMY/axUy8ZH8H6xfItohpkSx5y+cINJ
9jNaM15qmN3p8F/YdAMmdaqO/7IilU7tvZi/gCs1Wrcdmepa9sbiFupA4c5x0QW9
fi2U+hqVA3KVxfIcaOtCLu7xL35n7HbwF3pWrtjokWyv4APlnAXOPnzBAgv4kgLc
xYGGy1zIbAtx5ykXAa+1PYOt+LnDYa9ytZj8edmeTR4WmK6Kd2l6mOTfda16WoXa
268uXxT6X7PXoEHOj/c36dBpjOYHkizesiqnSd0wgG8ZVtuJKUTj/ZrvtCnGx6Pr
NGBGwoJexbnwD/nybCMMrIYCshxWwSUHKhYa5JL1XoSs9KztxXQZn3mLaNsiFlNg
gg0GGG4uRewgJDKwsBcV9mx5nVEmJZvcQgm5AGWNbxi07JGl4NpNQNkKF0Mjd85V
t/Kw+fdq6r+ZR8sdG1HZ7wqsv6Qx8uAAjV9Ht92CPR6WExpw+xFsO7qSDUoyk9FL
kzyWReCOTjz8n95G4Dm2WyHkPn3p3Zx6EJ+2MajtI7O8PhqB5RPamvVQykIcLUOx
bRE1m9bj4xKR/KhLkxMp6XErJ4k5yPoxw7RggFGPm+qm5p0sheR55T/0GJoT9SOO
Vi4V12+LcO7/fThYn3UT5aYaVh1cXaGIDSsMuU0xqObRAZuPW5wzq/ZjkNwHzY5Q
fSaKY5WHl0MvI9RhbCRyrfYth5u5EkWP/w+KtJb3g0iCvrALaj5uxBrHGTeB8Njr
a8W7Rvra2uInNS8sUp14TS6EU6EdIBiOhRjNX1NElK9iMT/zpI4+GI9jBliVyb0i
1lrU9UL3Bd2+QxYd2wZRO0O3sKflHKBTLgFfFgvzN+UVre87/j0B7noo2HVl8pf+
Z4brIWua6qDOn/cWQyPQ9Lrb6G8YhQ0IC9TnC9OO8mb8blE/tOSsvV3wh907/FK9
nzxYEA49RoK9JKNdRTQR4SuIRkL4mm09+IYZfTBIT77pCr447AqulVQ3F61ZGJr9
2lgRNBT7YP18/QH8O/9LNCcw0MeJv+GYVlZKm1wL5dsKOaYk3ChUxjdSXWjUU6XV
7nNOys0H787G0uBgIMZ+dNkbW71As4G/DF48FBPRjV8nYUpeJ83gjUwNkv0obD3V
0xrb7pghglXM0CLKtmtEM1huOFWe07Uxy+9sd+whGZIgEnWXVD07VcAF5Jd/Hpj6
iQhLplPIXL76FS5rDYnLr+tdSnIrH+8s/eS0b/FCHCtwExb6SVLfxMHd8DcHmv+c
tDCokKG2ivZO+ZoM6AzbsRaRgalSWrtayDqaSUN3E8VYvgty5odxcugwkqVgp2vT
KzoVZZfXQg52G9ARy8BTY1TzVMq288hDU5BNLNWHSZYYefqo8rblU3PMWU9Yo/zg
NsgBo7mLnP6J9nz+Qc2yDzPXO1ygdYVJi15bEL+cF7TU55Jtne/ZAmZN/MWCunHj
9RYkmxNVH/NLeUbXNYE78//Wt3wevxTJjaupAP8Mazd5k6ABW0BjMWngk91yafu7
gifsaaVVMxPtKwI6091RkL3cCJ/s0dDE0tklNALp9aEthswfoFFyzy3s3lYAkeaN
HjXMR4XKlXaAacMV8tOnqbQxWX1kSimcT3oTRdwU655TTV9HYQHKQT74o8UBcUwW
4jXlPd/LtyNkRXQjJMt4fiF5WBFDJqNBAUQmSUkNhdDdRpxJPV52AtN68mvXFM31
JLbosuGJzpHV60lxLYDgpD6XZDBaEOefM8QxmEFyKNXYVrhstSA87c5hdtPMXjDC
IqGouaF8ld1Vbn9VJzm+cCR7sf8OFF256EyTKAEy2s7VS0n8FmnJSekIgM0M0zz8
dZsETd/UCLrLFTku4+YpxgDWH9xvdVQpXhVZUI5Mb6fzMXLYiQx36VLLzoH5Cr4f
DLgccY9uiMlVSRFy0Z+oGmgbQjnyNQXxKV2wSGQMksVqDCpxFyEps5FAo898qM6X
HiVSj23DiRy/wuaKvR3YpNE3ROutmav+NgX6FTv2bUga+O4MgXMAfbRiA8xFPAKL
K9d3dTe33etgsVAnM1b7YkiUdaQdUQIPQnZE6vhuO9GhRODBSVbCrKNKf6PG2Bnb
7O1DekTeKNInD+9XrMlAvYwGR+puIsT12y6GBWASCr1X6CWaD3jTrEaSGjy3a7HV
r/vReVSST8HU+bAzIJR3qSwrKSNSpt3Leh+Ok8AJznonyyltR6aK1EJumXEEdIfV
y0Gh3BOpKlTNwxPzTb+E5N80JgMT0GSghCmwpPA0O0cBR49rf333mOzXCSoyBHuq
0EqeWWYpWawM4Yq7ro7lVDwJrVKB4WMnZc5ONG+NmBJuDlBC9b5ucMaDKYCZS+a2
a8ShfW/6YZ963q7TRilwgj8cyPqSXom8x+SsZSallgKv5SjC2N5xwfLe48Tk5u7k
ajfltGeA1kmav9RMiyko03zdYxhEC2SVmwROnTayUf+p2LaFKMUGjHsqaDdUdkb1
mXKhTnI/UFTOm0BEP81VCJ2kNQ7dLSqy3sF7NxL90I9s9wYRjMMe1hB+JebRWcXz
S231k1Yh2P4BeqrL/9oVsXrWATIRAhnncdd2JUVyvS0UaH+Xq7wb38/6rXZFvV/f
dzvouZ7vkvNZqiHrF/Zh5SEA3tm6MbOOimF7le2ySpuruuO0AlDR50fgm1QIWl1h
R8Ot0sGzI60nuuzDkD8QxMaMV71X3repwMZXvQQpHQVdvt6HMZMHYVYXW54C4tIm
h3I01uORJ5uqd526dXlXynpCn8KdHdd69jkBcPgGQ3w62sirUovuweLtIdQEbNRC
0Cmb82E+5NaVOnvhfe6MTjkCEmiS6BRywzmJ21bjoiTPmdTCZnaBLqQbweAgb4D9
BL3bBxz80yxGVmo/nIFMAu05va1HIX3cRDVdjSnIeSA2ucRw6qXxFxYkGSI2HbNN
8VsQy5Y0nN03zDv2RZS2Xd8GLgk2cnVHwsz7srAcVbT97VUcEPvgeGIUe67WTqmz
aehyAZubWRtGz6rB7ujhM+exw/9upZV7gJdbdkM9Zln4JXsvwnoSyDQxLTtQJzNB
WAec6OVcIKmQfy/vyuPxsUv/pGleQT/zYvbAYwJ/NTbt94sOzQsNxfTniSPbHcE+
rTjsviZMnMkB3VYScYXM1CsoaBJ1q/jxo0EPU28eZq13zRZ8SHM3M6vmTsY49oXa
TRTMbzulnsYJ5ePfQKbCCxvqIsCQ6fPVgrKMpYPLcM7bQQnZQX4R1FpnZb87Bk5k
HrLZj1f6kuhGtWcJBDMASLKty6nrvgkgpujtdctr9y1l6tC2B59viLj4QaRvDZiZ
HFXVAfY/olDRbgQZCYjeuf8Y6mh13ca0PsLUFVAEeHqnTUzmuANiPMY5/CFdaZHG
d7QG+ooPw3lFa1D2Aw7MLBL13E7WnT0zp0BwGz1dPefIoBVJuItBPznQE7/el8Xb
xc+BgyGxzrOWx3NwacZcbgxq7ovapX1iWyIBDKjBBkOEE5Q4s6Fxj4qXaTqYycNx
6+Wy6ACHPUTzEcy5m2dFPzsAJlvDwj8Q5mFtAh+MlewfZI6vS7MvWkmV3fdxuOKb
293F8LJ/BaBbouypKCAlVp4LgB3anJoawRRBYxudlWbHq/IHQiLjV7DU+AM5LMat
eiDcy7LcEnhzHG3/b7cM9UAkH04xN7sRzZjGFtEVYPNXMS33STZqCcSbu4OwCBq6
1omuxXBFay7F0Ag3GLS6lXuan+tQAeR1Ebr32cu3jTBCxS//X9KX0P8DFcAIRan+
kvEO3EBGEf8stbRZhpJ8EpxTuhSUwZAWC0fV5ED9x4HbcP5zKr3ynZB7NBcGqAVi
g45u+e3sRMLIWA2wE6+BnVyT25ZM6n6D7QDxtW+GuX8bKST458fIQTYk2r4cwEHv
2MFYTOJsFpSBD43HDL96+Rsn0g008tOeytz93QTCuMmX4m/vzK6uWQh9Yuy/7FQX
dg/xtpS47xtMglRoiBv7J/YHA9Uxi5nl1zy4Q7aHPg0UX4svpi6J5hXhWPsCFRsb
nPruX//uLb3k3DJaoRnUB7VAE5+fypWdo0TIa+Mo0UH1JxYL72A8VS84YyKbcLSe
eLR4Zf8BdBZIWp8CtfF7LXRnjY1rq9wTD1KMa3L0cL1DJC5krtau78snBy02imcM
Wg5muKjFt4BwD/HPvhQAaMCTFPyrLNhtw8VoaMtcpqCxaSAtS456/gM3RYMoDbpG
kSbX2E58Vmsygfls1/Ku7XBcRlAMs74R+LJ0dB6cmn4F7SDe5dX2RSNQ/YaaM/TT
R0B5ezExnjofEVfUv7BClG9UqYMNxOKJ7jFKP5C1zJku/Y8D8Iu/AxAkFFAxIs+T
aWcawZxbGWmahp1p3FzJx4llEpfhMkOoZzWJ2zNzs2itgd/3LbBO8uKnMXU3T3/Y
TWx7I3pFORDLlWk2UrChH6+hCgQs+P4LppyGQKh8FSxYbBRo/H9hYlnrVw76sEi0
9caUc1KSM4mDuRRsUICA2Fw9nvQpWfawtKtYlL5KrTIeNcaDV1dZuQKC5nbBwaPR
H0wKa6lWMcJImPXclGcLZq3RArvqdjcR6SwNhvW4En9ll+wS+gien0wfCBsGMt9O
dL7Bu8ygtXaQBXZRamyvMFBGyhYJrOiqdteIUrf6DZ7axU8xuGAA7uGgg3pVyxCz
pnn0SIbwntxaHBfC8kX3QuOwXeNIdaiFbYtD8+9jVP4Y8mMwaoFQX1OOHBfZhUJr
0+K371RbPS1UQm7nUq523CLrOPiUmuOjpiqOZjIzA2YezmM47yJwXBiye+90d+15
gV+G1mMvJqPxWK0uWCdAH5LwSjdngYaWEMl9qqmTjrD2PKlRWNmyf2ilRkoAcUMZ
U1Wkv5RXKcbOgtqNIGKW5vRRwFCvNBjOQ64upWZSMy6+lbx+EJjsboKmjP5BN9Pe
jXFojh7r91NPmu2vPgy0T9FRETmBJSCGlNB6HbKU0SwEeyWq/6x1mZdpD+krW0ew
1MDrg1cnpgqp2YGZNrXiMkg0FDwqmXToG4OnoqsaVBULmMU4+etvWLBfWiwpTTz0
CivkOTafKvmY7PNyq4R/z5FVQLetEV865VqV+4VYxWDiQpJFdtbbGMRuwI5q8oSS
e9ClL65mNnylMBxCheotktczbdKpO88s875fmefGBqbPDvQPh+Kt2nQksrJDjrAt
DDksqIIRueNPUbTfhDKH7+NxpLNtqO59cVTXKnFKWODD2WZAVoYVnkKud5boTX6P
RuThl3uX68B7OVcGT+Cpx0rR8Uqf3F53KyvKy0iE6XT6Pre2+eoDbAWTlJWk7O4A
IxN2F4epKuUiuBPMonbrK0TKKc7eOV+6MLzHAnkHNDAmWsca0Z4t/br1hl/+909q
fipFKgQ7rKHp6ATAKf7WI5ZEoM0qULvJ5U/2zw3X67BklJVtqdyYyeCM/blan3CH
Uo6fEcOyaMOooZZPzZEG0GsDiNtKSZQFWGSYmtLBm4gECXtef+F8cT4tf+jg+6l7
+bCtwzOKqjFiAoAEUDPC7H/eeThnLS/0eUfxUOXkTjXR6utJF8IJCLP6F2mV1qQH
6LkG2Pj+Ju0uPZKX4nuxsGgxqArts+gYp72xpjwy3DZtty3xiWENNs2JJoqWLTJX
cOHsXFSatsT0Hd0lF+wYfowXc9CR2RitsekSsbBcYJdan/dp6r+053sA7YfTGP6h
A4+vSpJqoP6p5cjD79tzH5DxhnaLTeVX3RIBdLtROPlVKbOtPWOTIFSDmrVNWW+z
88h2p3ciXGoZgoXgE4H/kgQeHJjCLGvtxEMIkfgS0uSzOn880YTIQYBlTVBXXWBc
mO4UHB5BCAa38ODzCVidi6n/waYp2mubbFWhoFUqpqMkIjwrDqjg2FYqmz1Bny+i
ij8mZbKVu/GrZktngVBAi5abf7xtk3i3ckC3P5UlvxtJ4Y/DaOoW/y8eR/Z3TA8O
xlufzhb9HQsn20hZbImM7xHQuBd+bK1c2q/84izgRSTKXLC58NJPLQ1SX6/FAVep
1s4pebfygFt7yUkYaNYTdUaz+Sbg2ZiXr7QG9TQ4pEtBo417gI3SMmcMCz3UHcBh
5kDNyD+mSeO9fSU9C64j2nHjbtntjiWQWPCMTNXCqbzMnH4eCW6W7aQRPTD+n2Jf
nxXD0yJG4hAnQBwl08jDP3ycInOKY6GtVdPzvbJWqEcknHcfWMUyQxMQRUMcj2GL
0+9pNc+tJYCjLDXDQzpYU50rJIusHpSRt1G6H/cQu7K1xsaoEIi/U18Vf64W4flN
XS/2j1D5Vo68ZyyimaZLHzQwyF1ElPXg8PcALyxBNfh1bLYqnHlb3twJH7UzPsPT
oyAHM3pCxer4UmNkiYn/qE/jpXGK+xSz18Hb5Y2Mknuw2C93yf+vB9lg/Mn6R+pw
AVuxvcmasxJie3dHF1mrYMFfuA9hCHph8yDGe71naskLGbK9MqrEwE1/WtkiMpeH
v+4fL8iKsSFDTfMyP9vgPby0uGjQWFN76Klc3g2vZolUs4vMlle+dQ5hz6NQ0mmH
0ZZ0RkHu4CsKNeBeG4pJdmrR2Ymhe4OvrQZ9SssSxoKvosmuXzKjPK43HHOoeWh3
x8cWqOFR83QPUyk2kFwxLO8MGSX8ZaMq3EFzDFurQXRiKVpemyZgDFYXDmTsMXqv
uQ8mVriHwr8NtsXU0EL3nSACF0eQCakutBhiVymQbBvMD4HavLEdkcHo1+dpuJ0l
exLMresId5+zT/FszEbp6bWv/MbZrMfxvTto3nfaokhUTsgS8ZdN9NDZC4rbhcD9
zovvWYV0hdsXBcNyg3XT2rch4hnAjaD82f1jAht9DPc/JNCUHc0izq8fN7Ke2Yeh
0JKpWBOYhMXxLXgt2lcT52grl0XwsWzDjRfNF47bB6kP0OeahLSAjCvGgAr/PNqN
/4DNBASIOmyHwBlySkxc7PwNX2UVhweQbfQgxuQ3T/N10wyJUGgPt9rIxJ5G9MNQ
Q1Lmh1tH6HhN65UO/bYHIKeFvjH6Hl52Abcf6HKYum2jSxe/+/zsujshz8YQbg2A
ONvi6yLJXpJfnus5LCcdjaM/2pojldwUh85n2xVlBymuvtUZYajqkFLkLSPZBlMB
/7hG0YfT/1Anb1YrBbICvkG/JkrvVr2c3pOGpEKqJFU6pGQD6LeS/njfExkZZEZf
xGe9/97VmGPZ1UsXR33zRnSJGyuGkO7Zzol0IiwtoJdJVJkT1xIUs8by/37h66YQ
34njQriymYilDYJb+3+zu/iwcoCUvlOS0mdetiLVOqPuc729yEKxbbpUPxt2w74z
JX74QBSp/rKRxhzYVrtefx4pMaBLeCNyrSIIdPP7uxUnk+U3SfoUmE19QsPr0Q9T
GzKN/zm3JHm1H2tQYu3Pj/WqGTIl4HyvdxVk9jiNgYzKS2fJrKMDpF0kDK33Y3R2
7fZbuYu/PknAt690J60/FskGwV8sencFDUehX6bODa+Rx2jkxCyOeKrB5wP2h4Ij
/2SKrZBb6TmkUxleCzSXSF0GfyeHcKf+Nt47um2OL96wks9X22/MXqcueyWzZn/f
xapgXlcW/mGV+1TeAFylyPoDkXozKKuD8AtnEtXgikX+QV6hIX2QyQ0Tsgk94B8a
rjfIwYqqhzZa6Fi8aFy2Cq3V0j3OEzR40FXz8zjYd0FP5Go2qkjnP0SFkTl+Lo2W
WqM/ZFxix1QOm7oEbYS2ukLLq3GdDdedwfePvfrUiV7wiyOVT3Wc7BJrl5rf31N/
o3BTuh90E5jAicrSCcmhWLRHO9716u16CwQK0n/icI39nR4gWyhQ2FB1R8vrv0E7
ZfnvcuLzyJK4pZhDT2FOO1Pt+flRoVbdWnUMAjLxSy6Ek8xkaRMTP/fFdwr5rKVr
gv4jEzqeNL8gW9XheACGxAkWH6nf8fffbdZfSTv/cUmRQUeS6QSz8I/auSrNP4uJ
qsCIYYxAamiy+wmbFrHi4qCoztbnaiI9Bl3x70rsiOKOZFBKGj1UQcoOD9u+zXjS
6Gl33EIZ55EsT50X0wL9qes3jgtSvMwCXzVJ6om8ycHm5sXcRWxeExfe1bCUvkAn
w01DULYPCNPUL7EuxchYeCUZd70bpRyIwLmHTbj8qVQhhO1k3+MpyyX5UFDEhKh6
EaXlLB9bx2mxU6NggKo8gBrE8pfrSwSpTWfB/UO6rL25028d1JmEn8aX+jFR8Gxp
sq4TUiFg29Z1gmvLRoRsEV1TZcrHKNg5DwfEYuwMElLQORTNK7WgshXiTXdgpRZc
I5QhGBLaPt0lXolRDrLN3lD4GnPypCZyYA5uoD68N5jn2ULQZQTZwmst0C/i5RS5
/6LB7qm12g+LZzNS+cjVh/hy17LBj1941sWHIXojiSfNf7ZP4O1E5qnW1MtpYlrq
VyIGSsrnTBytdskldGbs8li/0rdFbO96sQO6UkNcIaiNWm3RHPcWOp5IgcPFGqJW
55n7JHGMvuUaHeflkYJEGZcb83+kq6M/w8N2f8LqtnSxjmho8L4BN/MYw/ltncvx
ZPfWlWZzN5ygfcPslN5+WBCIiePNHF6xq/SShqIrDaBSdKzn7rUC/T6NC1KUrudz
PAPXs3DrE+Fn6Cf55HOI32OPZWgjRowo+TKT1zkw4yDQrciB1Fq9RPgaXHmKhLSk
qQhFxqLCmWQhjocpd9a2LUQ+v3jzbqVuCQPwDiwWGqcd+Dp7se5yCXbXGvS8PDZm
VEqQWr5aeh7XX8fabHn5Vb8bQpL4TZt5+KCUr+3D6Zf8SeQEClPC0rpplLxB6Bv7
K5A8Mbv88LD4eyiIAwxEaZzhfJtYeDKGgt+UQtOoSUPbyY/PPLcxhlzJAMgS36P7
ET5ZdSMzfE2PvUeFsQk/zbWue4uhnQKZ5p/irFAMlN3usNQYoTFaztKrZqGzzgQa
uXoMDHnzbC37s/Lb7kImUKIQCNOxmnuCo2kT4PBb8Tf3Cog9udwp1aiH331Y8Eqw
tP1wtRb7g5Vm0QpltQBrnfRrtFogIGxYa7nu3elGqCancZYOjn/q2kSoKm06aKNx
HJu6mFijE0fWtvY5hQ5HVaCs0HJqM67POCehXTqX3eaFc3nwtwyZheLF7OIYHgay
rSI2PMo9vtjOj/zk9v2xPXneobpIvSHtLo5TisnYfSUpJgf8I+o4sWYELzLX0gva
WzupFrMhZqH5ISH/D/t/EeTNibuRPfzOVj/8bgqpy0vPo5oELy/a3zBmkohUoHPu
r3qjnUjY3lT2BSCA2GIuJG9F0QRIjFJOsu2+K0z1W0OsRJw7prB6G7DE7DfjA5Qd
qsXFsJiDmoBnsfR8LtJ5Zox6pUkv99qxB5h1Lwqjdbb6bSl1itdhfhFo+/fQckrn
WSsnQQhY16K3A7uUCZVqlz5AySXsMw2g3Odyb1vCcki3QnXGPQ5yp7/WT4SepDj+
HUB1XtkJUA2YbMynK+sX7rUoAPB8v3McB2mu12xzaPoBH2SEOaH7AtyDRQJQ/02P
qYBq1rJwRn8DWjTdq4F0dlzGYCwb3GyWL+4H+YM/zA+Q3uoYaiy9pVNDg2zNvXLu
DeUng7hSUIdDH77xZifKHt+tajxpfhNfG0VRmHTSmQfmYQcZL0LwUZmm8J6VSICY
e+vi5TlahksiiTmVTYzilPcxBnmFgX2BZ9ryeCK6Oo7QiM9coLYZRZ8PzpdsCZDt
FB/GegwsK9kD73crdjUPQGjKgYs/Z0WfG192Orjm2B1BAjdHBcHGlFaVImYJmVu+
n3KDZEo/a3v+dkw3UZh6uVmQctgg3TTmCNrc5qOHUYTiD6CSL3vNWgOqZnWD8cOF
UR+7cqf2eRzUfgESQfiQ7Po4u1e3u1Cacm7l6IopwHVdW1MLSGEVa/Yr4APhjxLc
udAq2c1dPiEE+Q03sGX0Dsi1lh0/Jjddy6QoTB8oWD3Ds5z640EdcUX8ld7Q+9MJ
APIzpoT41rfcCQl1/AqweqloS1HkYrAJFP7Fn9PgJx5ovFu8cBJAr1ddj5nd3b21
Is7lH9MYtdGcRzviuUke24O3FtBweOrhlP9w1iKwMl/ULpfCFmgxFdpsmpozZS8l
540U9bCeQl73JdqlOM2hWcNRXzKt5msutcjaENKNAY6ffwU5aIGj8vc9cAXclwZ8
OiioTk00/gNzKQhOAzSQKv+fxKU4eszXBkurEwDTOpGkadi/7tQrZWm4Vlw3FRys
MEbXm2IBawWkyl9CX5AOl09CR6h/THfh1ZzRgIQz3TR7jUw1//hilxQbM/wu6c6o
bLWbp4i4EF0Amrt8o1aXRUkaLEo/siFn0QEycQGgwZmR/dTAs439D1Yf7spk4Tdd
gE60FxSv7rxIL3SGRIrQ4KfaVszasSS84n877X4P6O/6z0lAbvV5ZGt39KtwUntm
2Rvj1uTuBgLLPEyL0xwDDp1VOKp920cMFHgY/OPbE2Qsg24oGqF4mEiYurkHVoSU
6dbD8Du9QXnK+v3Q4AsY1Y5nVaBUa1KayFz2S0kxNTzBAoShemNvcRtGf4COtVTG
fyyjFYtMDRD57lGSt7rwKjWeyP5Wk9MyJYrMBk0C+Gyhcy3lb92niw8AXjsYV4tB
j9ty4Pk6CUL3F81xzA2pHX22iJJV2qAQ6GI170Xc/miH6PkAHJbMgwzCzlgiWEO2
oROPLJumlvzgQgPK/fpaewNMTtYR/YKkMLIYnH1M7PRBJYmDRhVXimn6IccU0cXt
Rut32vHYX9AnljfHgcW+vFwCF5+q2Qxnzdb5oTlowXtcF/xdyvWu75roh1/L+h/B
2fseZVcYOFVKYF60mBYMSZha9k8XSIKlD7qxfHZGj/gukcEZJTD5rLltz7gX1kU8
hCfqysxKOwrwxmrLxMWI5FJp/qxXt67sJgjpCzwYQ/ZwyJO4M1LV5+aKA23HIaPv
FvJmsdaz6bkAU0YHpPH05+27r8enXmqscb2/mXicnyO0uLfGP/LSTSEvxlc8rIx8
lUzapcEDl5i+xfC0Srk+69FxFgByYfO1jLEKCHZzhjD3GTEbUF/pokiKnYi5GAAO
7RNU9HG8duMTTwSwrGYXgjLLJTWRZTRDjhE0EV1b/JTF4h08LbCBjr/a2plbVRTe
l8fVk1A0S+I9BttC3nPW9X8InjZku6GEw3y3rMUYsVcmT1D7RU6UXvqVUGuhmpER
9+4xYbs/VKY0ALR0QLYMzxozQHGTu4vc8yT5+OIAkMbRIyAFaQ5uJ3dtYmsem20A
30BliF8OtSjzp+PON/eFEAutr+8VWa6TxuswHdwQGzF2uleqdZwh4PPQU6ZKmMhh
Vp3MZ5w06iU/l0rwboDw9WFFjSGE0p/9UMlTPOom4Rrfme5sE1g006AqtCZNIjjq
Py/TVQ52D0Ww3xzSKTHwLpii8VGGKFngRU0qqJpGS1EEwvM+QvENoVMMI8nTfF4/
fMbjIOlX8Iv3zfjs5TNVYJzKklrTGERaDA/PLZsBhdjCP6cfnrLqoepyFSkm/En+
EXpT+6m3lib5qmw7QrB9v9/+GzqsRX6MMZt1AxBLappTfICpwJvmamcfVFwT6o+k
zzNpoppe+LuOXPdl+/Xbw/iEw8Coz0GKD5d9syxM4wtb6zKJjU04p/CLAaf1Exfs
WHQ2o0gJJpQBIb2s0mFHiiMhMzTEpiuYTIaTvsByzkIU3oLNevme3kYdaKTxOFIp
d56mlwHm/j04jV+J62nJFt7a2jo5UI2BR1ZpTsYsiB1cZarBMYe19BXr8TYSqJcL
bUfPgXL5s/htTC7q0B4n5oHuxrVnyJuy6dtf9WiXtsE6Gi9cH4Z11R3Sq2NTCjiq
CkSrx6RubaVcXsWryCoq1Rmgn8qtwpChax3uqddJWLra768f85Ci+1/WSW9DZ16e
8A7QOyUIYCd91AiWNPL8KJfEil8pK2klQ8qqAwSbvLSzoOzP3R1XgJrGK/rdrjLl
UJ9hcmLnzAvpS3m6DS5zSLQyTAZrLs3wGuSFxDMvtm7gF9pg1Rk3ufgK0EVZKuKQ
lDyDGblxZXZ4tH5q4+9En7Cn0Vp5n2YMafzwfXCjrU+UaWHCTBeTnloOqWhWU8Ok
8pZKi/LPCc2deC0mBZ7XQcN5+f9EyWWAEq/9ITJe1oKI/r1C6eXayjq7bB364n3W
0WsMbK5/11KxWRmPBvgy6zJhFTdoTnfOyXzbzUbhZ5NTCRfK8VouWjn+zRZLA85u
XhUZQK/UIKUmow69fBok5coMB/oFUESZcp91Nfjerh+0klScJLn/3FvY2Dx9d0Ad
M44jCOo47aUeHuAiRYP4F2I9L84jC1Oypvp5fi7RlVqJ2d0sJ5YpVCscpexNY4HF
ms+tkPuGuSVZN05ni6kAXKbCqrtk8Gt8+xbGHwnHFx07V0fkgrsFACoR0XTrB0FM
bIMQkobZ4V8vmp+JKtg51RV84U+aysM3V/7LHswRQY8DEcrdsnh7yoPSjp+hibEk
w1fQXtAl7aRFJc6cNj5kv3IQigFmxIVMyhRlxc5dNxOfyuoM9bzw9duSmJ+cAEt2
IR1XS60cQmdGsMDCGhHiJ+a9arG9gyYRcj5rG1Rls/esvq87NQ66xDFLlaFccskB
FLKzwyV1VcUJ2Gu5Ma0aQZpz1I8yPXsgIMhTirKVTgOZA8xfY/eWdggkZvC1T6Gp
mlRILfZDx5XvHUdS/FKfi/p8b55vQ8jkGvUpkCFmkTTSe3FeNXkAgZnVzFJW6GE0
Svvfd20HUmwKIXLfrAVC5RtqA1tBja/WAIFO4vXmN61Q3v0vb1HxCUqOAkf4u4To
aUxFG/cn6F6hHfMrDDlVPB7qCYNNNonbPIz86JR+HsGy57Pp6Wff8OQULKh6HewH
6kaafhlDo9BBAvf2vbvkUgNIXSCUQqzourHdv+qiMhlKhr9cvFu3wQHr6WiOpzDD
F6eIl3nC5zMo00OJbZ73iuZR2OSm9D9m94F/T25nQfMK6bJdNvhO336bx3OOdik+
chITUY/uILW5JbC3MWCyCDnhZNLkwfGZ4Yq8fyppMbe1yeNIiTKzCkL0Xv1OGv72
kPFQvAm8YHRGOfLujqP3RVbs9b5YF7HJ6CH53lEzrQCrJRmndvGrPWyZS22EEjFl
PKewuLWpkRwLSv5bQS7eKPQi4ISEj38FK65v63P3u+BVQM1C6bY6QYtKbF2HUFV5
MF2f16dACQqjERYQpetcJxq+WBuGOqZxn8vqqgEVMlk1vhYpLbde1kdcedbDvx+c
PnmkwgM33I+oOl8V6KUw8OzH3IzyH7gF0pStm7ZcV0UWHMhG7mtakgqkFJ0h3nep
/qKYyZA55H+0z4KtUXcGjoXwcEL8ORgqcQ4ENMCh9NXrzO/jUrqCcaSq1m1u+kgi
jfbvc+a7HLP2KoE1JQnzVAxotXSqVs4RVE+gL5sspP/Px/TwpxlMdBtJj7STme7H
3Qk8ZlknxESpDRISCQ344LyRnI+Z0lm/mVNJtODe2KxkUIQvXcokfGZa3GASMF7M
U6V/eu7FG4xpv2V5He9nS0UvFWkeoLxZ6pmK4jP1kBY+7EnXjwffiHo78m1lDiH6
VHdLIkRXjkSHFuJrfrCzBhQ3l/eCZeu0RJQDD5tYsxrvXq7MqVKoAzXUAu4CNHVX
ROHWMMfZczx4yqjNbiIR4j2VyN2VRakX2h7HcflLYZrxfHvvVc71Outkzeql2YyW
zSEOiPnbM6RRAA9EP+7QqioNRZkP6cyN4gaf1qeUzsVW+WkBjxiac3n8u4sPE3Sx
daCQIc41mzXLz7k0+3Xruha9J+0rD9ErMKFbKdizJIH7ujbvpH7oX4++481WsIVk
t+8Bzznyo9qjl/PEpJP0FnUO/LxQTqVF4dQhv72ZUjy413EtW43dlpxCoGmoRZHT
GSx5zw96ZansMeCK0pI9y4SfgQTB0SSPYxmnv8F95SaeVD7cYYCu2CAPgEi69Qwq
SnEXvMtq8ubwzofCKpLyXvGOWPjvzB4DtHmWti+RGRIghddK29mzwsAVU6JyzvCF
z5Yxkl0yKY4qcy8CXMyB+VDN68ozU+Eg0IJ1/33S/T4z6T20K71V3fUnk8c1yaN0
H7hb6Tmt+r7N/JFM2IUFUacstZCUWoWEBAuiYBHQBlxHRubgFY1AS4RRxqoEXz11
HGsSJNfsgGOI0A6zqI4C8uDGbeaC7p8qcg2bPCm+JgxMcgh6Q9mlcJzCpgQgTeKj
1iLZ1vYHJlFRVkKGZ/8Ddqmj6ayJOsFOeeIJacUIIqQfU2EeSyc1Xh00qbzndt+R
gNjeVjYGKIZD5A4g8f4CXkGPgSyfyWbdFHnJcyR84L+N4DMotHvMgunIO8LfE7zn
GL6EpA0gdg/s+Q4xjIo5UxbWb+h7k8tGlm+V1yakFwjtaRf9NH4eO6Qfu06if7hk
G3phSHMw/AL1d5J0j9oFTxDEP+Z8dFl0G6qpV0oRpcSnsf+7pl04jDk6t8ldx6zL
EsjgZ9Yqc5bPd7XyTLQItMziLhBFkUWVKl54zcLhQnHFEG1u9yfc9K7n3H5UEftU
TcOutT79KVvMkOga5O437grT8YLkjo23h489uvhNsuuCM1bSfGtm78i5uFbkdNXm
VAcgHesArr0l/3QffMQ/cD1AWnw677dDf7c98Hr8x3ahXyi/lBNmi9GJ/CI9gsRy
PIewRtOAKqU592Wn9D26rFjl27EunAYRNgsljRmv2iTm08fXsn0CsKHi0k+PE2DG
hIz1bmei1bzgelHx4IlG0ylWeLB79hAYTghUZvbFccXtiXDbwmi3S1Yu1Sq9pftd
6y/v06wbAz5eBZxjBTuAOWhayB79+Ruj3I21DS+8u2R3Upav8pkxs6pTXGArblxJ
Yuq5tAR9/+iMZ3pcF1F2MtH904lWFnhDHqRvz/9s6NS8UoRCqa7yN9qOY/P7n/x0
mR+SPZpZnDE7bn9XXmtsqgAvVdyUsoifqcr11klFVJNqS/YdlNoskWerwZ3swYXS
KMyz0fjpbfoDXRO23wGdH+JUQ7qyh4pHDtuWPurDHlwA8SIV2EqlfQSVJWUz4JdW
VrlVJFZwTbJPN7zBXCQaxX2bXYWHwGcG4UtbIO6lJDs57PFo6hTgo1chvoBip7pQ
ReqONVIipaCuczRMgONeLbBXLULSlnAlf/qsTTtjtoFcV53FmjtBBloA6r64Lqxz
8bL62RMZejDXOzRen3n7u9T990tE4ynKXh3WkOG2vtAMdt95/T4QbkIIt1kjZOYy
mvkY8eY7GDM8RhFzJ+wBV5lH4SVwna3z1BuwKpbcjktiE6GwlHPzsPkJYk57ks0b
jliFjd1yecYJpe9B2TGWsPO80cw4SPen3NGk0OwDXE3r03t9d95zSOspj30n8lGW
2SMBcfTxe2BVfHpod1pIIFpr+NlLOw3eL84xh+ywhQgFqeN3XN2MQs83oVVFags9
svjgyoN2964b6WV+T/9tuw1JsQMeGQR8QgOWMdwHha9g1WyJCrtUEoGt9bcs3nKQ
c69g+kEoFMksUgDXNSLwblKnHy6plxZeIJq+7216c9hktaDoeO7Ky1XuKgO+I9K7
AJJ68q97V0kyetBNSKXh81c7C3crL/ty4soNuKMUAkIf3t27FDOhE/KAZLwvGqFe
UsbiCQWPzxpywDiUM05j1UVjlWM3Z65U0qwPfrcAZVFiVpGBqGZS+Xg13cdqFPVh
x96xCavvk2w9IvffEVTj9XYFfeL/Y2k3XE1siXaU0KqKi5zLAUA3/ElW+P90Z0Hu
/c/ZyPky7zGlSdHNe2a5zM84PfmZ53J5m2MFhhh18CWCsrZGwTORdNq778MzdWj+
t82LEtbJg44QeGIU2IMvsfOVMvk2gGOfWC2s7Hy48pbXxtNNYNZi9SjlQUYN9eqm
G2rSuWNMXFI6JOis/0kWAX62VSdJP/jmnp7Vh4J8B54f9CGPFAzs0rjXsrYmvF4J
aTt75UUqiotmPezBmW1TD+8uR8Gf0M4nVvXdUn2B1WB0suYqN/Qv0wgenEh213/7
34vHPsQ52xj3MvAZxuypWJx2DrQZlRNhHFyFwzzMxVmpT7N0JQtDj8sgUTDas+TD
jjf6RnTUfZ9J05jHtg3xD2mG3XqJ1HmJjcX4rc81gK1Qnes5U7ddFKC6v7slhHsv
sWq89kgVG+wu+ceO8DLwa2RzAUrSuMgzecCO+OwogrTmjUoeEYmuSQPXni69xWLh
KkdglXI0PpUrq/GVhrbI32WiMvlikDC+K3RXaxYor+hCF2ApZvWI3sbKvvnPOLh3
6lhZpK/aug77D+nqpVvBfj0TZBvPcnPiQE6WXAbP5/aNB/fWdZjhK8X7iGj2t2io
8+k8Ylc9Yt2tmNuY4fc4U0aEBjVD3iizxUMejdlo9ZlH9Xr+Y+Q3lkuye78mfDQf
40b/VLwI6GECbvfczfgXhf2ZavOuOxu/CeFHjjw8cRaP/Yd/hw9lgiirHheY5meN
NgolTr18AgEejlRNwppNCdWSHrPdiAg4Gk2x+rjNim7al9RDLC4enruZs6cZScsZ
i8HXwD5CO1zdWHUCGRQSECggI4mueuZD40Av5ilWVMq9qm6YcKHTli4GT0lBX1Ln
S/iSuoDe0cGKCR9phdzhiBwO4wu9Wcx69IncgWIzhQ4qEMY2BiO/2TllNY6Rznv9
W7q4VC92xhQAlHFovMXY749QJi/QOwk6arw81b5COOexf1PbEqq5Z+I0KGj7koA0
ndWW/WobfR5DIXtYA4dN7KYpeYnUK6pBs4mrN2Mwqwla/PzF6Zyk3TMgttqDqmlQ
0ptCkhzbLNE16rNwakbp9PikVXjqIzLxQ0jefNRdNz9AYdlYq4CxY30NH9VbdOl9
bGBMfbTi0zPlcZRiptQFmFBoGLcGUQaQDjge1/peF6RRo4FpfFajYdq+CAcoGChs
AbaVWwYLop94v55Dw2T18aL8pcgH0MrwCiv1sMsXfcJeA7KI9jfp+JwHyQeVz7aP
Mn6vzQaNpJ1ve5J+imtpNgOmwQFChUX6tHNQjJtDC97mMrVj/rppm59mothqsAcn
M7a9fkjZnSWHScRXl8bWoWeUAXgUO+Wgz+DeNK4woRMFb5cV7NesAspHvFPIEZcY
G6v2UpM+4CyyRYyYmdECnVMlMFZ85yyEd7EDa/7tOH2kLn5MXi1fjmhz3vOGI0EU
zLlBpixr+xBRFNMrwKkgFFPJ5z2p9DiG/SLY2PFINHj202Er6IRLITqkYfYjLdAA
quea+R/F6jG6XFrS1oQstqmYLpkgwVlTdygIYvqKEun7Z8l94zJ74j4jOO6fFvLm
3P1nvvdM0/DAw5XEb/ru+63lkHYpgauL8CaGMRbx0wQt63U0P1ic9W2vd3BVgRn2
Bm0bR8wYzBYRGp0APuZNKfcrg2L0yEwsA4jcI1lUNYfuzLcgsfnXSaeFS4I76yj0
1fNVIyM7jFx65zO5dZSVwJPJDFT2Bj1Jl5ThImbOvEKPUxKX0tnYA3gz/WnLySn8
MiF2UlDvVliCytbfk3vjUtNSujho17WfLsuzkj3aAusBhY7UayUsvPZ6D+S+mMa1
x0ESBS3B2v10mubbFxg51HaU1FZ938XgLdCdc/ck5geyktQ27YvgBOwQPFvWjX8n
H6D927Zp5/LlI3xgwFEHU0cwukNT5Pt7wTKkYNU9IFG95fG/oYosg3W8GCCBho2A
UVTLrgaLh5NTviKE2g7ypVsbiIwJh3CIlfFbVcysvSTUBEZ3l+6mTkb3Q3En45c4
cPPIpOFsAsfHZERH9/JyBeSryuyOURJFhbo9eqD+1nqePU6vZBrc47obdbc0jxKZ
uMBOW9S4xLAtvU+hl7hv6hKk33sQMtU+g/oilTcj93sPOGGBkABnRr+IWArK5tpm
/8v+FIKsnrV7V55tb77CGbfw2t8kOm0EPsyKBGrag5xjBF0Twm4t8aW0jU3MCiz4
+0OfCLPI6PZtIJq/97wugB1lezuBrr36p/e0OfKdhkuJuJNg+nvLDA9E0qP+FRsh
ojzNgl+ZRsZIPOsk1B+JXFvPvi5SJZbmP8+6wgrni8iiLWMj9IgjovFdRAdBCB40
zjjXp+Ca42C47ExwlPPJ1J9fdSJwcomkocKMxYJmCzET/7mt8DKVR9+fQEaiFH9c
3b7VygcoOxqcTEGL2WvE4n36JE4P/JfbFdsPJdr6FCOyQGmkGoV2ESbnoEVChdgJ
0M1qYZdLCALSxmag1bpW6IRoqyy2dHded49AQQarE5Ff3Pf4eGhxgm2SI20AgiVI
PH53SqBPxjiPzUlZuLTo2BAniIDutMOitMu5vANLVSQRlpenWlUhx/n0bbLmPnVP
J4zLfbSKx55gGlM9Jvhbspn3OQrS/pYh8ONrSx2Ml1g4HR1bO2iZrQqb4KjFbQR6
1PEccZCU6rOb9DcrCBC6XhEe2BuJHNPcO/gukcvvXeFgq10YmroUbpRd82+tgqI4
TV4yvAe5ylx5edNsyLJx+ZPl1Cs91wsbvQXidpTLhfqBKBzqads+b3kRlg9JVob/
Eg/S/VCXoE15A7wNmdkucEw6aGkBWLOyV4DbrCdDk1FBs0QAXMVLvpnri2mB2FZA
QKVDFHS4J12lONOlq2l+Tu7joYiSanCJghu1t7aoo3pjyLksqTNp8vvIu+CR5sVF
VP/ZbeXuWMI3i5HBEQ3f+giwZxQROWBih5NKNEAUPaQxOC3tYAR0OgprJIdgPoZJ
IoqWG6xI//oIH7fStS2FFCUexRhwi5aW3AFgbQAfauIAjdj7DxTyr+dcJbwBqsxW
0+NWvwEPmR6RHoNjyCXuc9nY3i7TtACkbmnlgwq4QjJ2/UUegk0XgVE35dQBoa4p
eT8v2q8fL6ralutV4jfd8TzMJs+pyDPKCkNm0CZ46Bw/Gd5g6fCEbnDIpAzTkoIX
mVJZDJFLsZbjRIvQl05cTmZWUn0RC1cA+c+OqztbkvPhkjCBY9Q72d2t3H9kEa3X
X3v8t+Fnsdwx3TJA8uSsTScSppkVA7/uo0XrEEG+p/kOvJNzotfJ7lnfUANPWT7o
Zbial7jtOzHoAN1JEkoxj2mvGaCYeH8uhTXiR1kDuvEiW9ThUBhNVq4D4LQDKOxi
22qKOkytXzESzHzrRbWut00XaGzIE7DG/Jyfxg0RH4gzPRgCd4zqbjcYXwY9qaiD
27XKnRLr2/w429jo2uAzurrHn7s4tmsL8rjvXSIBVq/Ixt1DrZlSbDdceT60tWi0
GIwOuSU32IbGcLINt29PzAPou5EmvYoH+J1EyIkC18aiMPOzphST4QHpJ9nkDB0O
kCThN+8XVmqEquio7Ht29SPMoVPsMiN37ThWecApG2+NkhZOYcTiKMSjG+uvdMeV
b/Q/ATuga1F0jzrlxyVYbTxo13J1MlKkWovujfxSgtRzkJXKLvibiA6/TvJOkciW
wXgMLtmdrg+bsZ3xqOAK44vW+qMSc1198gVDCgw/VirIsYEgYi2+OlEO2klTpMsN
nG32luK2VIVbqQXq3VlUVQw6N0NC/DOHarl0PDvq2ZDvFexAPti2uaBY5IKjFkW7
aW9Hq7d1/JDfcE7CQ7r0jSyFOkBIsatGSwB0ErRBLIIKbRd8KsMO5mCTct8M0Lnb
clwOWCKboTToAXgMl/FtxicXU8wwnbJX7mSHlGuLzmbEtjupHc7+4azlckszy5Z/
sC5/yaa89CQBwsR2LHTNcvv6jwrGf6U4ShDe1aFGxAIEL9FD0ZR/8QBv3voqSoUT
yG3mP7+nyGYPC2x+KezlYQVXllIqrhYRzrisP9CCMfVxL9cPVk+5li/0REsDlZdm
W3b0jigkWTkPyjyhgn0Cn/CzFdSsrKbSim4l/NSwYtF3TjgOtpWjdStlyCf30vc/
dZRpF1fCJHaQc/U0RPXtlNEo3PRqzmLzX0XbAinU89mqQ2NPkM8vTcwMOGZTpwSi
EdHL1fGgv474YlbUvbGeitTUU9QDndtl0ucT/7y09kITisozvqmmKRxnu7riUnqg
q0zCSn8jmrxcH4n5pjHSKE0Q61+1ioSXR7ztV91NJ/IFTrceKzTMUljev2UH106E
4CVoL+XGZty6DgcbVEs/zzProDYAi4x96CcS9PUbxJ8yKDhj/PsMXXD/v+NMcsED
ww6D0RX6g353rzvUryTKAfja7KolF2RGPGtbWbmDc5i8WOzQ3xlwhZXKsODf3YfC
/jKs1WGpj1sbE0pW/T0oTcd2PcIZWR0wD+mAMkF75TOGVy/wQjKNahZX526RIjgN
ADNk4P0pFEHBx7+57pTYGpIy/MFAP7gg0YzvuZ8vl2m1eBWBPpw26YN++R3Rtams
wXod0hnyn62R1x1jfuHvxm0cwAXQnOilD3qGdLv/ilxAxQCYMEdjh/EVrDba4LVD
SBT0LlFVtBcsHHB2ROb9JDIH6pMPlkebM5yPJzbSQ9gjX3Is2wfYfQcWm4ZhRAG+
OaEjxazbjaoIhroxAKspUXhcNlwIRmyRLJ6rra11LvLJv3u84ui7Y/98++izmtF5
U5HVZ/BoohARjct833jrb3dJx2cvv9ZmtXFRFqZHIRoVN4VttE/4FPQRaA2oFuxf
gh2adwBtBxKW3KoSjy1X5MrWLNNi3em2RLNBXybvsNwUYWaIixT4wbTrBxdky4DR
53HpBtU+H3lhE0La0MvzswcPMtVcfsuR8E5VD22siqrb5gLqPjdBzsznRjp0UHq0
mlaMRkMUe7r6BVfV3IwyBCeIy1j+JaOQDR6jqymNgxsvFxV6l4LaqJ+o/j8/N1/r
doLGQ3xu07+/f4+0xn+cKmXgLSkIr+UQXo+crHxbcsQu3lNUAKsHUxi9YcBaSbgt
S82au4TYTIjAjYe5QdTHIC83YATlfMRHdJtqjLqS3mrNsddo0uqGKa4YLlToQkaT
B78Ltf8Cw2wAneuojEu8RffxkbtbDO1OxopPpBK7UU/Gd01RXiNxRcxfh91tl40t
Rd1kguf5LLWxQ3aZn55uU+xi/ohBVIEt7TGpE92IediMKFVD7kdpntDqKCEFOIzs
b06saxXls4KsNA3pfUBXFVBMpAfvXXFVn7AzPVyufIwIVBR/bDzxiYja4+ErRdTq
qJHv5P3gPAz88EQc43hO9nsGLrxfxHtAl+N9pWrsmCtr1JnpCGjUV1LjdNxnSdQ1
++xyKL0modOX0c+AHUqJZc4fn1ibyH9P0UYjPuiJdhnZh2QUTyNjjnqBuiy2Pvu2
5bOeWErMeSTNH8QcI/l2OPX4GwHT5E3Xce3sIz08GQXD0Nq5ivinsx+1NDennEhu
6KcmNukRPsik/+LrnUH8Rdm473635K5OqoxsZuWEscaH/kW4C6zaJ4zno1IKeVjI
0TqyfC5mbhrKM2j2JCEm7x/JFi2vwv+7uEhtIcJ9HJ6J/fSu5tl3/WnwQHTO5HVB
oqnTQ4ndbtuOfqo5/u++7/yIJhNSbZ6coekhMheziBdeDJZOVEeVPHu8c8Joz1Rl
QQGeClmX7XwgBmkr/oKUAKvxq/HHRMOlsmLoVF6MAQLiserclhQXul1dO9Z0vk/j
Ey370MYubPewmgublXIBMYdtLWjvuTL1wSuhkVZdjQKOoGt45CVtQcZc/oIoiJew
h/CNZKjuSnKBCdwra6Z7gU7VGZGkuwE97DpSu2M+KCl88KaLUx3zhlnPGaIOnY5n
aW7rSqm59FwDkOZ2cxh/NVKx3gboCs2Jk9Xrr7TLe3ro17hLamBDJB6pUdCzavmY
NYBT/WSQUoGuTVZi7lFSLMdSxIFBMsAbTZUvOmgHMo/dqMcSm4b8YRqRDhI7mFpO
AOfRRYIWFk2Frl/X+mwrfvr44Qmke3OmlzdgLDIGkmLD367q/JN1hOeNvK8N0Xbp
jH3U0zOXezgJfw8z/3VNfR1LRVookhyY6qqgUCN7xHeoq4NT/kujn4X3hyJZt6sP
ykfI8p7PrxyS4MvlBZR6zoJUD5rAhFotuKRQip5drWVM0zIu46kiy7eIJFReXm23
6xnRkFef30gg+CJHWUJNuRanfpvdMaiI2N0aZxn6ANoyzaAE3ZQxdbFb1jR3vhi1
D4R7W1/7uXTFOOYcuiVp+f3hOntLEFCD3FaMQ0yfxOqwLHR/Yy3VoBiQL48m2Nqw
kqnVOLMM7oKnosGxt+UQTFLeRrnJrcOewp2Iq3EezQDDmqRMBepD8OMvOqdeq6Nu
qx7jkQv9nKbHbbUKJD55vI61Onla31N3LtvHAcnZv9PZ5Uv3gUFk5kV+u9VfRR7j
CMlBp7jemS5DoQVZd5JE3JVCK/gEWYJpfpssi65VTKfpatEME4gMSa2VWshZyT0j
u4F+0odvlLthC5N5w4/75QuQvO7PD9uND/nZ7tbCHrkg6Oud/VgyCCuX+tPqO51S
wIXL+zQPFQLjK2VZt+MCMvB8MgMk9y4nkNogqtohAGtf2lukyk1m7+Lipkjcy5/b
sgn+WTVVkSiMOChCzWCNAiEdAGuvDC3+HjC10Ws/5yu3XC9LLCV/Oqluti8DaS4E
ZwrpLe4kaN7UQ3fH0XhI/gYi0c5/Zm/T38upppBScv1BOsHfUmcVNgnxdYJiasQE
1X/xwOkMbk1P3fQZxUirNL0+ka9FQRigQKZYZnTTNY40DX4EmHgUFM9m+UZCbB6Y
ZD+VS9AgXq+B10dSjxT767Hz4HhFQMgz/Zq9vpS6XSNVOYBztOUeQqB12Fs/FUOl
BJcKrJp1wqBoucuJPMk8B7J2Pe0reJ6lhfmLGvFQCdFbrQHYwNKGUP59+mRR2UkN
ahJnv00gPEez2VCyHhU82ST9Kwwb7EIv9XBvyqhYi43jPEcdyrxhLCRwK7bkVLdn
T4P6TNvg480YXqcYES02cNCG7s985r96N1PFFtYZlwNeaq/X0/vXFnpm3YZWmjum
do4E8mrWvFu3Q9DK381X6LPg0RtiI/dUoL0rPFc8z04X778MWqQSwLQdgZFDEvqF
0stWyLsrazHPQBpe49yBCevWShHG1kQrp/zxkN7dQrpYDNykN+QB3/g+7Hl1wCvz
xz8TTonYA8MB/S91QqWD/zKWje17mTCEoaTDuErF5C/IQvmNpZryOuuPUldMmvIm
65RUxM++n6lkQ6kBHzHDKbUbN/0nKWbzhHQ7nMMGFlGc6P02gi0mY2Ytqu0fsNoy
4bBscjuWPw5sYlTUlxe8odkoX6rKEzme5yfmQlmEETesZNi+X8VkWiSCP6WB/fyh
BJ4WBuq6KfcXXyrIt4ab8eWi7Ww/1GmCyHewQjH68m7HgCR25gwvbqz7Wq9JqADq
LQFm5cbUBZo7sAwcXc8EqvHhFGLpRhuEAJbQGoAw6BdBH+bVdaq8MsKpEmKkSokn
73gzGME33qYdQjd1kD/ppr0sOcjbAUOMyXD8tDk3AcHe99j6LSgzKsoQBvKggAqY
Cecs+yEKYwXdu4aPQ3u9koW9Sw+ql9oqSdzfnsihbd04Uj/dkNswZnZxjDYPE3Yf
w5MI8TJdanGBD8f+xUW3tyI/PdIMTEmrS70BAp37xYk0a9bqoQlGhoVQ6KfQh8y1
L4H+OKtPeVOy0wB5QVzJZYyorVLtuccNje559XQJ0vhxju3dbIRUVFkUzd8BIvEP
hqzR3JEOQltp1yo3YEd/AyLp0gsK0H6chPnjRxpIKlcTzXgooBupLGLvbbwF/rFk
aDSNpztCeiNg2k3Q97x2iEtIPwO2v/MmWittYu064jRW98YEu76/iOhyGP9BnHih
UpwqTYfGFZslmRVBi1BJqHoOKq0YgEpCpPWik93hCNU6idzEBKaWqmFXnMSCCWHN
wi1FShwOtUNMDGy2FATlRAPqyH32t/BLwh1v6bNoyZ8nxRyRnHcWy86mp6vC+7vq
3MVUNvzBb6CcJ2+Scg8/n/lO6iZ2KrOTSvYls2kobkO0gcS77csfgm4JZJG16srZ
k1FkxZXWtxiBdu8qLLan/svdRyekMEXIDMAkcg4z93pSKpjWDGiIqEjUIU5heqnJ
uOLVT4ni1Ty6JMf1GZz4hqz46pUb1dskT9tRxx6tszNx6ZskolD8RD7PoZwNsOSj
8n8V6rz5irUPL9sMtGkSDKYVwDMY3tHZZsVocSKSBvREu/sgeJgjHbltuNaF3b06
5A8X1Js06uglBSmFk2O4kplEAjneVBcOJgi/0EMTJhtRVb3tP5MeWjtHQmvsq0k6
dTpMcuofWLFZttdng+uuw1eodylyDIAh7s7/uyQv5p5O+4YDFtE30gkbarbz12ec
dvRquYEClYsPZ34+/mZk6oFFVWNU+vo781ZPQMZ+uXIJD4rZ0ZTxvL9It1dIUk2a
ukZqi+/4dJ4CA3YuCYgtBOkmrkloTURU/QhGt7q1kNwcsMvy21z++4YMgc5qpp2X
cfewq4+nIZQpUrw65l2RWQd+OA6j0Lxbdt/WwIU+a1NZjyvhu7dLuYB3oaOpKQKH
aJhB8sVogz69nMfGU4kQ1yUNLp3INK45+mbw7/PasSlk+PTuw+EXFCzZMdb5/Enf
MG/H/8/PgpfGYhE0HE1e6cRPZMopJPkab6iwDka8tppyIGeCfS2ALxslqY/wCKd5
+YsettnQi5OG1H8wN2Gdnert5u3kfeuT/21NOXeZp/811+T06wEDNOcIP7V+G/+f
DeHWpOI/KCEbhfyXt4+zfoe+UcdWGgnw9DVZQnlp29xBbsO2EswiS46OzfDo/n64
eBW583qCON6CeSF64fmrvzo3/0kNBFEEhQpUgwy0RhyN+28IZaAx6Yx9l4tnoH0o
KE+cRlVHQkfXVCeniI26chFp9XapimIW4moJd3Y/iPCrlCEl1GhEYsBAkb1WZrZS
RUtm3UAGg2VbnZILm+2fdURkDGa8ubSShS393gefZQxc6/VJXwoTyGafxX6Ej3bC
sALwwuXoauKzLGdGtY52m5Pr5mKDl1M6ETz9lxLroqb8LSb9hy2XmJwbXEAvxZ/e
/EJD7l+B0e0JTnkQbtskkjLhvTIo0yx0QVsTVxHvWOdF3WHB6kCgYsmhf8LjoYoj
5eu0qqHNXojO1A+bV3s4DIl4ufUQ2LDyB5VlY9ltK8pRpfBQ7Bx78XA2NAvW8HG+
3iDZnq+3u8BF1boZA3rxNJ6EBovvJ68YCFuNp3AoJegODxCQ+4IPGQ2FRe1jLE6e
HnFWsVCwvFrpVRA/YtBxmdG/WWHmn/xSR4zukws9fIUAsj8DQYkl5SEWlTLoa3sk
4OAwRrGhmev8Cv2iffLm3O5z6M9mXGkIEpNrESeagaz7g6fQ92vQCs61OD3x8vhV
2cAddP3pTLAv421l1v8NSKNUNnk2gFkVOoaW91YXvzVE44rDaDaSw1Qr7Q13NFGK
0Q4KaGOxu5DamzYPDHAmMKBLPMXFZeZsLaYhDYBUx5sFLZ6mWVbhs0Ks5j48UJkx
FvIYvUiOWj3HmKbQBuS5Q4JwnQRPzJ2a/m2cdCsFYwq5F8SWTTJNjh9LCHCiX1gE
h9ll51I8To60QDMvNORfaW/TvGAF4CmpKjit/MSVkzrn5GSIZ6a6nOEbTWQNp7zh
cUnj8SGWnWo+UEjOSDHHPT9KufWWLj1UeuqdMADdlZ8Vo2k6TvM7PUkySZPRBvoS
UWKhDI/43UiSmzVSsK9SWR+fJmL743S3eL/xNfwxXfm4qiSuh77DBNLDcEVXYDfV
ZpeDmzlMDJWUUCOGO64+b1Qpb2I1jJMHahr1gGlKJKW10RSo+Mn+nWaLHChFWqd5
Q2wYgWufyxSP76j+C9nckohoykLrGtEqc6TjD7kPXR/x9UnaMnCXocKL+EHQi4tn
zGsy/+p0GKRP9Kup48NF29trtuIswvwtTHgl59a+UvkiQPFoG10cfWu8y4G8racA
MDp/nf43x6wih4MiPEk+nZG4ZLMfnzOgzpnZEDu5GIFZgyDJhNchUA0WoyA1qgiA
Wl6myyetGEmP6Iaos6cRCO1xdSEQrBaFi9ynhuWly5nTMjOOXSoDF2tRkej15mKO
48RhajBiYeiPvHcVi/dRA2DEm5Lg1UfkpngzzRUSPrnmIYLR6r6DZKiSNH0D5MOj
bWr9Z5grI/MkZnbC8RDTxfSLSWg2SNfw1zYRtmFDwxalUmUXGhJbELg9rvA5/6/q
VBEyyoK7C08aTu1E+EqONq3Isvi9fSIS70ih3Do/UkJPwpCLA8ZBpc8z1SHXr3p5
avfX2vDFFSriDTYwVbS+yeJ58AVRbJUQrTbKnrBfaelOte5Zx6ptGs7T5aAx3+fj
W+wWQ5eDCjqSJqWe5MX/UIFW6LFFmiCgtPx++I0rt1khSVVg8v/r6bcyFAEq9txW
K+w09Am4b3B0iUW6A+B8kzogGMg+mEi4I0VUx6HabYSsPtGslUIhooheHe+SSo/C
ZysaxbaUDpRUAnyp21IrNmXQPcueEXrRmfdYQ2GHywOX2xTY8MV9/ErpKy8xVa8w
kh2UUMvRPIJuDTM3DEY6GSvsCuGkuaQDrpfHqOUY+EBAMVv45PAZkrHaqAL0JMNM
uNI2WMm2jBNBU1y4EBeEgmxKOOUnKFek2KBJBakLpFLDh/bd+DaAsN2g7wlQKxqU
E35SrwWdoMC9SnRgQo8U9fJdZQtdEpADMaVde0ZOqBvPqJ+PFY4ygUG+HS/tsRiA
BDh7hVgV3Xs8LlAO8hPx6i9mm1hl/mxq/25TrOuChsPMd450aoeh4cA+Gwg4V3fG
QQFi3h4rZ/xjJ1Pk6TsjblR3i6QJpiM7GYg3AGy2xeduNnkfZ5QOrNPNtunm3oc1
iUD9adJH4K89+cNw8xcv3TwZks7JRKe+zNogf0sKIi9zETINgXwfIucGcQAimxlT
pd0bmL3ukEHnBYaMa+IGGveut6SW4wdP/ZbO37/xrG5jMsCK9BIIxT+pPdmtVCtU
u/Ft4ks+DfRFOTN67IeLN10uxxSxW8bmOwxSDl+apXzQy4if1dUw6NnbTYO6slQb
rMR7ullbBLGAyFbHaJyNXkgb40K0+ZBdUHrHf0uetLhvS4xbK6Fr4CHM5cTWzz+2
8xDklZONYxJ4BDN3J8uPXyCzAK/0yE/LmXN/h3x4JDnQrb5QjXylkxqxa8beXGJq
02xOP8633JAHACjpeaLTcHaTygpSK+ekvFH/FqClyqKFYkVZNRoHMTej47Xbb75H
T9qBaLSmT5o6QWj4DpK6/C9L+DeEuZFlEw52lO6mtIUny0M64bXgOlks4D6GLTKC
VRfAbauP5Gw3erJRaX5S0t9ftQeRvaYN9+NoHT9zkHE264XuaT32bD2oxwheG5zc
TDjhwQ6I77ywBOU6IAtIrKESHSEPBf+mt32jGmiXpXs7BY74fF7H6GpR8uTp5iQ6
YCqzN4judf2aVVO6rphL4MfhN8d4Vr3CMQKLpDbvGMYon3iIItcKJe8DkbWQB0Sz
L0S/HRezs36J1Pi3stros583gCau+kmpTcaYCvo22DmQ28/gifIbn/1WbjWiNrq0
hrS1mVABlLw4Xlud2zy2Fgbn6qEp8GfPMzhtEtD41oXeZwkoUJloLcZv4nXE2Jza
dhUTgRrqr3fDb+sv+bRX98v+rGfyrtkuWsY1/5fMzxcbGhW99kGtoSXcnNbE3f8l
duFnZVsIWgQRlwX29GjaG1TaEGFZilOJ/WhZRAwyPU/Zj4XPwXcNyB4d0b2pGXhb
uqhH7yNNysWaphoda7vT2DNwEmbDuJTnrNAjMpBLkfbqDndbBlugINKq/BJ90epL
ySuwA5GK7j20rdjee4MmETyzrmaVzwHORdUHS0lgDRbe944FoZk4dWV7h+Zf8+/d
t44b+6SW4AQB18wI/hoVpL5XXIdymlyLv9IVvYGVl5QlFFPbQhmc5HacGgul3j7t
/HltVsMxgjb4ukExiPG0rzasZDkZ+vdKPbCP1GP+9Hh487pUXrs3d68Fm8wG/uyk
2JnCArnDDQ7a3HpiPmq85NtaiCX+7K8JB402/Y0r49GArM+WsBh/sRPL9HpHaafU
3jh567nY0k/0N/DIClaoixT1oLl0FRo+LPKbS/app4HTBjuwhXxHHw1AV18pcZGu
K0JxscSxSlfsdvM3UZqRl4T416rljtCaRHXcUt5N2cILIxAZXkSFVCdJPShFGZpN
+QH3crQmRIPout6eQ+I0IorU8kDiiEHpbFsNAaK9wOkbytIWuVTdiEgltFzukO9L
Yu4JxtcuapXCwWt2sT2BMJXde8oFhJSJHTlpLtC8NvbI4pYbMX6v1FUhmV++1T4U
Y4P+LNi4MClDf/Nrre/hZGmAfhWzu3DrRar8YfNQ346nRpcFgNeTZEs1oXiLQYE1
dBKPU0fJRdRSOvuiID25rJtqJ67cMStKjSsVCLaSVrTV0TiWqn2kPZOjlgb4zn+O
pIO8I/1hAfb+xttEI+hkfjmcODn2ZwDv3FHY6G9HctU4PjmLv/0Wixl5Zr2sfeYG
p4yx84GjoDNWmOLZ8TWFMzPuxLQJdn1LfxQSY6X3kzGqqhTO8Ps3EzS4s604UIL5
FM4U55Yi8oGLwOuVIOHQTUbwRPa0e1YW6XYPaMdCVwCLZt4hZDsilACTEI0UN9P+
pVopwiEeKoBrcpskXnQLV7d7hEAg6qth3Ad/F5yvuKL7ZbGZMStyhTI4nyyq6u9y
DFk4bW76gMp7nG16P2WnxXH1pAiz3N/sbrEdy75+Nbc2b/ClSOU3dJmV3w6c/OzW
eTU96G88QQam9XJW4IlqupvK+xVfrSD1xxdn1tdDz94l/2yrX47N5qeDZ4BBRSIs
tX0rzKXNgszsTTKM99n1HslRCdT+rJNRRevj0uZV35kCm18DwAT0BrGvkq2zS+tW
WS7vkfmoF6qKkZ0V8U8Z+NxmsyI9YElLYGv0/wswelsshi0dJgteCey1r5qvj+7C
uR/nzPrQ8R90nuuM2PV8fas7m1MthXfNELsXujB5cVG/BRXKZpgAAoxuMSzTdNpF
HJXXgj8Ug05Hiakg6TWO7fMHlYlFDfW/8QR25QbSpzZssIctRJ2XVcVg5HrYhrGW
2cpxPCs/lUof9i07uD6yDwdW9WsYHNkow8JfZH3hgpmkp7Kp+Ufdu2XpjzgaH+3o
ZZbe/o3+7E2bgxckcGPXA0yto5+osrVZ7h51ymp/SJ/W2lHr1d6y/r4+YjCMTi/J
ZF34v0N18VZPO/e07/8bRjQTIp7zuCRp/VzKQw0DE4pKLIUlfB4Sx70aG/ALUOIB
vQT5j0GVBQUbDdTgYggM17kVKC3eIIEnVZRVRM0VRtWVbJ11MLEhXq7PHJlfOZR+
dfPeR0k7Rcyttb6WeGHQQRMWOZUl+oih/lKyMLDF0UL+oEcslf6m1b3fLatfHJDs
lUlw4ND5Yz5IaodckyBSehfC5Rp8rCyynxICWDlQlbUeJp+DmR2TmNFF9IcoFkhP
vDff/kiBsu3EsgrP8FkakR70fzzreY5vY0PFYJRdPVdgWPMn2WfQ2Qq9tYB+0AcZ
X9ILuggya4BsNnVzx17sOCCqpFaF6q4CSp3kt+JmVZ+Xy8UUTMRreR2p+mzkD2N7
tRIZf3yq2/VuwNyAQzX8JiRjm1NAPL7uJ4BzEokJEpcDuzaDZmUTPGZFadVw1AzK
u8x0tU6xhTXfdnr8tSKONha+xYyjLBmJa6Fr+9CZdS4VqxoCIZZOTZbpMA1+7vcf
FOlWnwP2z/w/QzBm8+UImO47qyZoZUphZ9alkE0awfqxnJ1yAn9YXAM089LCtIp1
NkBHrA2pUUpW3cPP0ipgILyFvNz6TCJw6RH2CZLTLKuI4vWIg1lv+g00NI70fDWy
22dGMgMS1v0JRqmwHpSQm3R3S43cA9K+Y1hETQ0eknFwdaysHwgSpKuPhfuw6cCw
M7cQVPcWbtNLmi03QvH1N6jDR68w6saxWLZ8O8MC0gXydTMVr2mvBbJ6+oYjmtNS
mhontyZOarHAmLgDFWyBhAYkJJsglPkOwn6fmG+u05XP2FSQCtPDRwjhtclc7etI
PhcIVyxV+xKyFlB5Vk15yCJ2Ap8EmUXFZ2hRaoVLB7CCc9DSrnPlzAgEDQyexVp4
awTE1xUJbz4h8qWJgPWXxzccKOmM45KYNqhFW/s+xWWPMH17puY+MUF/HVKIXIKh
RR/SKqq5blayKPGTYG2x8L2nIq5hSNTdRIDvogxdq+/bFajmubCE3gFORk85HUwI
pUqEqf0Ss4AasvonUMfboIvQZRn4QuV1N/nJnHKan7UyPok0++i53/Mt3ZXCrOFB
9EvQbLTIknxNJ5TygIXxO4PNjMNCuDmEjQkERjyN1SjLgGao0tngx1UiorZds/l7
1mtZGuZfFDV8d1WEDY4tnlXOqw+xdKWki0umWsVibcTf6iAobheB2A01VtM2OlAU
IUUrQ+JJnnvCoptV99lwgsZEHP0NJ7+6IbZRnsSEFYSuvcrZkd0MaRRnJXYNPttd
WTyf3hqhlSWavfjMiL8CR+f6EQ9+6OMizaET5oU4Ku7ypgg1OnWPVHWNllSc9SRs
yo4oErnMeiaslJEaO3MQhIIVqcAv8mh2sVPG/zOgxJbsIChSFmJuf+rtp0PBjAx9
VbPq7tdXKefgYJVHU/bxexj6z0i8ELa7zNEAKuhp0IXb5NYAe5PLvik8aJlZJfso
lbJVUZhlgBDSeepz96ayv6qJMX6Uo41zlfc4hmamt9rcu/sBzu22ZsBd7CONR7Ap
Jb6xf5+ZuSdcvfpyNfbonbusYiTFs4mSTksYz/D4McipByfy+tGQ9xTuw/cWMkFe
5OMrCg2GqzbG8/lH/kmnS1ClMowaJdsHwFMRgcaOeapksYZ+w59fs0jYLXEMxGMX
BZ0yqnPnJztICIk6xJgTgOBYlvcgP18V6k4cF412rhGfOZkaIG/Bs8/m1lkS7HMV
lVVN2fDP3XviSt5s8HJ/FGmjIYlaSxvL5CgeUkgURRQ+AGgh7MtUc3ErWwqe1I3l
al2oiulEOWleAf9PMxN/MS+jbnl/hfQ+cW+wtmMeHDdvkN9iwdFRh6jrS2StM+NB
F1xKqw64KssSuWgB2nvC0WImEVVUi5WsDqMlMxRJ64o7NFHy6nQaxPQKxw0ZiWGk
K3KhdOXjIEbbWS2hztVB278Go5JNXm0ov3IYgfbzjzi3y7MF04q2gvUBNN047ig/
IEsyF40g43MV3fFwQcPRCFZNbfJNi5EofGlBpcXEYahwwgT8F/m2TYgVYALqeRWT
6ArAUm3dFH28pTXuxjmNJk56HPFeS6SITlg/GKxb2KAlvWZyTXEGOpBt0pQxvWyt
jpv3hfo0VbxdXNH99ebi0K65lIjq3PHn1hxAvpSlejcH6htT5FejUU54mkRYk96d
uSAPwnJHWTfu6ppS/6zxUg33rurL6j7KA81Qid9Wyt6bWhLAAcYR1gMzhqC0xWv1
hFl8h4VTI8AtyeK62d+5HYCQgZHsupARrLe9MYS9mb58QhXhFhCKWyhJEI3Z6+AZ
2LUkB1ln+GmOZ+JsanFj5ndUjjlGddhT5QDdnVDrK7XolqTf3uVU/M8Y5m8kIgdy
lFQtEt/Hii26yREuobXsZl3/AkrQYcoChXt4gLnlq5m0l+0CInk7umUhYWNpnkHy
Olv8FxQVqG6XYAMhjBXH1MJMSY0qnBdiR2t6zGww7jpN7teqalpRL3lS/0/3aO2m
UlwdnAG7ixQWEZbuyk+vc05gDaUKxfJ61BTXDH8nW8Ezhii/ULI7iNxgLWtEar8S
FZgqTG2EuEI0BTWj6NSHcRNvSZNkKeymVA0O3Mvv6xYIiCqNG+b7rEeYxEb/rwvY
uC8xdoYaJxtSNEOKc/zhyOyxYVPb6KjvJ+cGOqoHZZhl/aHMWqDGJ2EJ1kdR6wZL
GIeimS5J0orP/b8cwt6/4LSGB71Ov0rG5QCXmQcSsvvjSak2wUQeqGs40ojONSYg
taLDs74z3E20qtIItjWAuyoRmvabiPQLz5QPd/Q17lDYuNqoVOHqm04t+MZRJstO
shh9cg29HpEeCFkDBJpZtkC7QhcL2UD++eFRIviqjnV+0pz0BtQTMgQ+Vm91lcEE
dM8mLqkeOS0lgibyIhfyWyS/udvCAPGgi6SiBuxC7iJai9oRedQHQW6xGHp3/hTD
PYW/VarQMtgujHa22W6nA+FxHH6VzJKRn5DowZtX9AnZTpHCaz28bcbqssJk5luh
Xllhk9D9bm49LP3ES8C9dkSIoX0SOBTN+Ceq9pXY1wgByWD9nB9XBkLBT9dPajIZ
9cUoKjJW40AfQAuWNkwxtE3EGRjaxrPUmQXod80LUpr+uXRibDUTzWlikwQypxPK
LoeXCRtTAksbrG8Uuq/40XBODmyRHc+oSWYkJOFkw5iJKiWU43ACnDuF1qfPnLkq
N15OoZZHYTyWTzAowwCwGMS9oTVNaQR86QYkacs7skjHu/f0wIOAzpAqG2cz/95a
XkH15XGYKerMXnC/v86Fxl8w8jP769MRgeDrLa2AmxmXehK4xRLJ3pkwRWGw3YvW
QQ+vrSUc2gYwc9zOkba543Jb95WwkyPAT2/kAvoRtRYooSbnCM4sNemQDJXto9WV
UD6fv4OfnwH25QCC5FjSOd1HL7DIf91rqjWqgy+pO3ix1HLXoE9gnylfV+P9lNel
bLCGDhiykf3Pv5l6tUoRHC6QHcZMG7cvsV/R6G8q7REVzlVurQKwypPVyV+jL/6j
RzcwfPoQh3P5q6zWjABesS0IA04khAfVy4DT/9pzrt/js0JvACAn5rqu7sCrlejm
9d6iiKl92HN78slwFvMoSXX8vlpEA00bUk1UvO6MJGXv5w2LU7LdkxDToLWe+S0S
U8yex3Qz1yJpp79f/Rp1c3k9KALXybwHbPqNVJx5FRcAr+gp/EOVVSBUTNDdnoei
cLIs2oZiNZAEEDV85w9NP19W6FDn+fKclK+CyGQ0JuFyDr8FnCXi+DFOWFxAxgc0
Lfv8KxKSgVdvEM1/ry3rzVXzvHyu0qRIZjiP67vEEO1ZtI27aYujmasdJVue7TAp
WmTFZPXh2ANb42QkEK5g4OBlDF6NuJlzmE/myFPadpEaKkdgsHD4BsPWuJIXlIs3
5nkpMLf3I5nL2tjht0WtLhX9wFmzUHospCN9f8xHFxBDNn0ptGDVNDAq3ul8nG6x
ybOMbnP0OCit7xQ0Dv34eWeCL8tQHnTOIu4gYjy8BOFJNZKk7O4IibEJTaYWXRoQ
cvkLMdiNQ0rbtnvmXKAcNpTJ+KbSHyj9q7JOtA3jUz/mNkpgH9RJ5kA0YIMFP9SK
0YUJhXIzbf4TyjLestt18Np5NidToTKCyr3nH8qdD3x1FbcAuttEADNLRs2UVR33
D0F52o4FBYi2M8dqCiaA73NfQEVRv4bHt7OrdoYaXDoY691r80DE7tkNBTm4xT2r
uiBo/xTOA8U8oGGoMRN6ueXwMCMY3+WezGSnZZ/Vi2MGQMbKYNF1IBkBdoD5m4Le
/3V44DEw93Ru1krZwckZybCJl00+leDwcQJyU1QBpvj0q9nwi6jQ0Auodr7WCb3K
JesBimp43Hb2OWOdSCNtD5gAA5FuQBYTXe3lo3PUAhkB4Qj/jBBE9WUUscOjz/0w
+7yOvCyMm6xllVUKYovOsmsem01scLf8Ot7RJqwvX95j/SJOERsl/TVumWkqZrbn
bvAjyRlE5IwNp4+gpmv4rwTlMSqbzvSGM18pz1JXWqr1CK2rDi/izZ4TiWpyy8Bj
joUU+S04NsiK/QKAW2x4ZPapemTP2kB8BzkDgKRQ+WXYA7I72dQwwwWBrilMp+xW
qiR76Gf1YcfTmGra9v6buvx1z0jTo4iwZnqiP4Cnw3DpggRan0xpQIgUVVpZ0HeO
1jWNGTzD/XNjxt5bM32MLAFPUvd8CswSmgvdRJaANga0iKxwjyhQYG3fFq/cvHrB
BRldOZEBeiChTLjFcZv+jB99iNp4cDPMbR7PebgRVyx+GwLKnYQ6/WLlEVUt+gZk
qOPXO0GcyyhM5lUJi91TWbHH+wvV5k8CTIqI77zWmNIr9ba78nGlQWwKbXy6ggQQ
IudaPqL2NXNkNH/2FOj3vV32zRAh9MAZKZb0luXK4rTKMBS2odx2574MajyVEIxm
+KV3NbDYjvwkfjGipLPzRtTA0qxyIBUFDeXw7mmpV8zrRmtZPZCsKC+1xxE7ZoEQ
OuDgduA4op21otj0QSIutxT00/PlWX0x8tKA5nvwrvKyefoHOq/YOPcx9Wi+7O22
w2gsOnruKW7an9N8ueItxMoE8prDWb9adgLJ7Iy4fFXtMR3LtXbctwDfGDGdCn6b
YRE+VgV1T5jdyhcpPWDPVCOZRn6bKxPRf7n4zKH94f4Ow7XD7kWYgLRP7MstJRQh
c/1TLJTZFmXY5FZeXUT24l7SfrSlZr1vCty0S9S2zKTDzTn4Xz1K5zON+6YulGJM
bPFmhtJOnks88qTCyIrGbViZnXx3khKfh1SqkOfdaT2bPYlu3u0ASGyf6jCFr+3Y
h/h7HdTNkHWGJEqJEdZq8pTrPI+d+gijykJhIcaoAPaYpB7qMTKn6EjUYgg/N1dW
nilPZGr+2WO5n5HjiXHGE3wsizPUfQj8G8BE8fOZs6/GwR6v+o8EAIUN5Gznganz
ZtXHn6yCoCj540Z0YWiBONgSx/oJmJlYlHQHrNnCYy9NCg8YDX47qiFqB4n+qxOs
tn7ldWQI0aY/+F/eeUDlBVTyrgKIubp+hnopSLpQKEsAXfHYofVBs1szNZwHsefC
nUIFeDyUyxE0+zPTzpFzNO6Bt2Q+vIyiIrfmqWjOZuLbxOOCmU4d5ctQFAqqTtLC
VmhNoiZperzRdNfoknWsxncOkmDgQJwn8VwyoN6iTsiymDwFMz9ScMDnwDdEkgNJ
B5QZlFrNl0gZoh+Gg5OyJpR8XbhltkdKuibb5XWuqzqaOaSO0hippNvHFy6qT2EE
vo/yvLjH0mj5Jb+EWRdV19BDPxfvLP8US4NUp5LPiJFz4lwdNv3z3xaR+91YObiv
K2qWxb8zU+id3TpNRjwd2bkh+Wb2go1dLiUsdazbGXQPYHR/ZD6QQS/hHKN0iZHI
rHgbIu4P4bmKMo2kdXTJYlEaeuHdwR1IxGqsgAMB/1CB2zFSIFY7yO/lwmRVUlT0
TCDCdrE72WrCqm5nc2UfY/uh+LvIjA7vM08Ci7/mXWBMwpVD8YD0CZegwQj1kOzh
Qxi2MaL9IgNI00hEgzUzI7bfcdttmOaZCQPnyURJmzgsKpwm/HR2oLFU/zUu0mBK
/M2W+1mN+rqi73pAKFdO5trQf0GMz5K6IFBIuaXx7FDxly5nqGFCadUbelIl0MVZ
rWVqRId2e2YOisVAcRk6Dd533dC05L4B24oPxVvT+Nf7oAJGjPqLYIF/K6lfM6fp
yyOgvv8vMmr7Sm0hxTsi69yMIYaUIwKj9r7aGUZYuVH7gvzHmuE2CmAwM3VGsocx
bR4LfD5CSjDZDq4n4pzcPl+lUoAO2PW5GYH9UfOjIkfjCtQsz8TPnQKn+58ba/Xb
oliJa2eNmhBP7xiZG6ZxXVe4xaJd6M6z5uY3LvykB1TTGHkYUOLHIFWrV0pdFID8
FLA2MTLYZNB7BfbL+gcODHRRF3Let98QqGdKy/hkkMZeZMhPG5BjNd1lch15IaMl
zHTJz76AItuAno6HePpcOJdkfF4T2jF8aU//YQI3hULHohnFbKJysKVulk6vsQH1
rHtLQX8d2gkA4BNCg718kf9RYIu8rnlssy1z8BGqEHAeLSQ+OMDWrGrny//TGJET
02UJQjcBCafC16ThkRO7WJ9K1Q5tIJPKc0Yf/qLIavlfIPLqpGBjulumBTJVvgcv
xnJvegO8rsf9am/lmQFjRNq1svNr697jWkGVfsLM4u1r7uEmiuDyrnDXyeo/wsVl
wC1DEpD2f1HSv7PNTUaOIdjTXD+f7SNQa2f9Go881U/pFQ9f8fRoJsAKPr7TqD1W
FvABadOdWH5X7ZlUnL1xnKWgRrMHSHB2bgkwH8VNAOfkYU30V0IjGhLoJsF/PITh
ydjWj/0iTI5NLySZXw71s6KmDXCpjGW/9e4s19XNZ13uyLUvkvFt/LXJO0dSo4Uq
+04gpnMlA/tk4fOhvG1dRFssWVIzAMmX8CPYA8YrVAyTAY6zfSLDXO85xYhvDQ46
+S2igmrB84cz1UjZCCos1OxX80LiNmCHoLZcusFUt3XEUdWfUDyL12N6J/n8Eq3c
QPp5ozFwaroznwkdGWHw8d9AlF0yilDvquJnmlnvIsy6G6hFiUjJspE8XsEJWhEb
PRHkUB3dUMtDDUQu0prBC0IF1T4YSqpK0E+lQZBGFsxVANDAmjQXU/KE1t/BHdwL
PmlSX6lYQ108SQEIOHbBTgdbHdQntV9YoFq2NJWZUvHKm5DGv4k+ZkBa1TscYjm2
N5GJ8Xc1ypsei1JlXIJItZ0vvdKTsMxImZ4tlCiGoMitXCluwj0eKTmDL0wmj2RM
v+hAcIZ90NgB/5wUSnbRD6m/96v1TMeBz4Qyg+lhDgclbwfnn+y6o32YATywGXgD
OXfqY5zcjt1VGDsSh+q5FP/STLcQDQ76wY5ksLRfgfEpfHOHT2R9SMI5DoG0NAfs
xQlU2NB0TtVknNJ3A3fMBILn1HETxiwt61x1vsgRVsfJAksWi1lDgvyMB5Dz8djU
pmpGUl+18CS3F2kAUGvaZaGQdz7EeTjumCry49mVO6bkxWdhZaQc0bkhVg8IDxOv
g5QOh8Cp5eULdw8SlwfT7PDsLQy3ZsYBA8KKoUV8AlBOeAEyjFsbfymr4IezaGAM
k7SMiE01gGC9gkgZD53SJNSa7x00bJee77/QnebueHcR42OFpURCp/pZ+F3/UKAN
FXkiqpOqyqhn7HdGD1QO+aneuI+2SB9IXSf+xIsGKZnBnL5/EPm4DuxPMIEacP45
9+jWENB82wgX40agFUp+RN8HhMgra+YWdcOGfux2bxt8UMdXmkSFeQWE/MYE0w9i
xFR/TbvjKtNSRYlYetD+cQjhsdxpP8bdCz9Fclg3LDXwk0hnV/8Nk1p0mhQPkOIh
6yKs9RKdPY6IwoLzjjiBYi+9G85WSrBtBZxJYI/OFgCk7QlkMhxpEU2Sbx01zxDZ
3rwC7rHGfU33ONFFTjM/dJUbR9d/M9abRg+C9CehjK/rfAAfNpGF6sEMQ9mP8ZwL
kdMvhMQhL71szVbPFYppQh5OoIsk33nU5U0g8zs1T8WFfFEKFmEk0XGaFmLii4Xp
QNmJPMB1JG1ogm/LWAl6rzg9xeQbLH9YUVeh9ykWuCzEPfMbbV7a9AmC/L8yx84B
xZt0pgR99YAfMgctSfSvbsdvslqHGkoqDUvQxt0npLhSFANccv2oam6QYMOT59n+
b5tl0ow9uKstmiO6K+Js3pAWOgsnlR7kG/Q/cz3lS443066OSjo5euyxguxBMBZj
URb5KnwAVEUaNE8E6cYOWmugd7vRqpk9Izp2enRTUvB9BrzkP2P/JUqQxKn7rrib
aPlWNmks9n4+uDKeyimOTXy/cyJ8gaJmwACRR6kbQcZ5iJtiLeD2l7phS1lb2xf2
qsFR+zxzo1X4+88dtSQoUMzHDSMdzRrC2c/tn9+VfbltqviydpoVZNi7ibovtCMw
BinxVEshIu8CQw3YcaHiWtY48zA4zuMnCGyPN/JAUIeE27L7YZaXYCCV5HNEVETs
ERbamjK2ifClRfHsiuOsW0vhYVm7tOkBJKMY9WbCsAHc8v4DsRx+/JLfQEFSgfT2
zBMzyrjlpp4ajMSiUjQFsgwrTxRj5KaF9YduPAPafdtU6md3PIOLqq7+mnRD/4lo
+CFdGWWaJhCzMXYGXsZx/yZ6enlEQV7b9pPKgH2PWul14AyGRFvNE5M9t6iYj5ME
0dW5pUreX6OFqN0ioNjuOA76Dexmot4MgZhMpMq4QnYmydJt6FAwA3Dxt3oz1qKc
pcPsYfv6KLI13gOaFbETaBxTLXfOyL4w/RAAxb6OA9baKnfVHvsTPBJNYHOBthg6
TKbV1ubwlO4FnL0LhoJNdz4fDLQzACsKvmj/2HFMygJWmugqaT556ie0j/ce/rXG
2e25ECa/ijXKKAqFGKKkAl9SuRJw54n0VXbFgjoFuoiTvveoYjqHOAVb8HvMODW4
tQMa5YxqIIzgazgd0oaCyAdTQrConLG5CRXtwYivAzwFvrZfhmzHPSqv0HMr4ado
XA2756TKMtBRLEHC9zG2ApwstfklekUKroGm3BlHDKxkr45v9iGFsQaTkbemCsAG
Y0Iv8xA+ue24fSG0/DQVxpvvbsP+2J6WVwN3oLyUnk/sROWmkTmomBXTiAB5n/dI
soGEEU9KNssmzaSk6j8M1WZJBQ2nFfXbJ6QJkKISJwXgT+K8gozExo+eqyHPl4ZK
Vnm3cI7uOptTb3ryBZA0RjItR3h/ROx2O+ysX9nZF8zZgwvanKdNEcI07tCT3TZS
To2xWj5LkctjyMoBXPgBSh8mWWQjdQqUmqHp8J0FUngjvzMht9iSzv6kn3r8QmRl
av1vsh8rWLUiFvJjrLQc0Q9ZxpvNBMOpiUMGZb1oKfysxPvX7IYAR9D6soIWZenM
6lSrt9s+lSe3NaSYY99I9BZwEC5YWvABxiBCJAhxVoAHEbz7LVYe7sAZaaUPU0UJ
qa+l+oRJUDy5yRitD9IoniNHSQjH2+i951jtLm39CnPLYpABeEbyIyEtQsrQxfI6
AqxoXdidjMjsqJi41XzTqwX0P+DRolSiElu53j4MgMIrQPhKVo+HzBADv4bvmlzg
xljXHLXbHBhqlBZJq1PB+GZi75WfUbUSXhjXfc+x3htIeStM1Vh/03rguWnnygE4
ok7LYkimQG6N9I7kYfIeQg36wQq357Z5YOjAn8UfFvFK7bE4d96moj1vIsBu1GG0
V9xQKozVasXxSNEzjJc71h4l8EnyjRSgXPbrI+R3CAhX/Ow3HTAMajnbbj+yGk9O
E+gcthtkNU90t6x5VbSSsOIOPdBoBGC/RBrWRj+payr/B+AQM3FvAsWCA4cQ2hni
V+PF74K7MoLMvajTiCXEj5YlwGzsRmM0LDtlycksKoxyXhUzqbg2mjmOc1UwVLRa
OFp7laJnQZoYkSkQ4EHMxDdP/lBfPtsjJitUWf4fTQuG5GPO7T4U4iZdbd0B1FJv
izCu9o4pS6bgg3WZmQ7uUaiv1PKm9bZL9SEMtu0F3gIaF28H05fw61iZBMaSbMIX
KgSJmrpxLm6iQziLM2wGdfC920rl2xhkHF77KR36i3/q9f6E5A396TG3wINjciDE
GVTDcpD1vkDK0QziaskKL2cgkeENq/sEBZOYG3E4ahN4LiIHnrAtFxLdTJyY3Vm5
OesKNha7plCGAfWB8CvysbXCHwJF4evAfosrL7i3cptQCqMj3W1jpX43ENAuh+u6
MIBnsXJY2an2RrNm1f4J3vGBma1AKLqw1D1hGeri5HaDA6lUVPTgDrynUkp1pq4h
+4T/6k/vvigSHZ8LQumSlWOFPkcULRLEKKs1s+P1+mXTQi62gjH/acpnqd/fDQgx
X8SJjvL/j53QU61cGv7r5G0kQ1KVaokEdr+Wb6q2kt4XfrXRBWsPCeMolQ3ptdUb
Wtu50BbpxD6KP8Hlp972ra7PVJnOkc3Lhceb5XsYqWapG+7ohJ3Frc0DXar3uVQq
gSERebz+ubBCCwbsssvcXnhYy5HBtOVRqqngm0fYtQS2OVchrDEEIDZcsuWle+nR
NOt1uYRAc0ZZ+kZOCkDimjZZb2oBEc5TYpV9sokQi2mRnIO5aCO68m+R0UzTt8xu
psPZ6gh+ubPyhnC9ydX7RGJWXlJ/cKAi4ST11aYcDP4Ekfa75U6j8yCDOQeURbTo
cCPIa8ccC8LNeYPUNGMkSYZtY56oSD/sMiRTSiRrk4lcrMnEvIO0cLDGLAMpDedG
C/DJ3Dsr0FCcCH8zRzt43W3aCDKu91buKeNsD9LoPgyJwfzfif2fM/8OfOfeKZyH
B7axMcUVyhUy2F6OKpAyVx4B5/MVrgufUYqPkXCs9rjWcsZN77IU1kMPcVNkeRzx
kspn9215XHk3IV5afIgC4MFW4zVLuUJ8YvaHy9j3E/RV+3z3X91xyG48a5SHI2G4
QgitiSfORb9oSwQNhGKQ646ufjeJAeuVV5mQAY9phFi0GgRx+WLqBbXfyg5wB2V4
+hx4Yg/9W50mnFjadASIlBE1XgA7Zbx9wPo/N/NYKg2iLT+oIp3l93thT40iWKM3
DSaQJlSEei27oQ4prZKA+D6KKwfn1XMXYvvOlBfoaSgs2oB59jtdEPBBSUFoz6Ff
XtUizlO2WMIJF/PSvRubhzwWimv07O2406HDk2JhI/xAD2duGi3248hI55VJ5cLz
4nJuodLg8FV/v1P8NR+dgRuePQJyxvAp/V/eZpU0KdMmv3LW+Bg0C8yaPZ4+jQLI
tXS8nh4iiNnWXPB+37gsD3UPZAo/yJ2oEKO2ZaYikl9u80/uE2uPaZr0+4Cl/KdS
VJKV1T9ZNBc2m2UsR+5TD8ViuooCtOU+Y/05+uOky8VZ5sZrIL3XSywNad+ZNj1x
3Rv4fReYroDpCvqr2rCKMq6xL/s+4fXz42cdPrP8vUegSuqDPRBUV6twqJ/eSA57
IisXKgVcXUpUlkdU+64FWCODLeEBLkhujeCkTdBRtAgwmqq/D+UOV+eX2zKP7KMz
M/xAhGveB1NERhvYr3lbW67yMTGlZcJlga1Op8euZCIZrRIUNpXGWV+877tCAPt6
99I6mcAltlxGIyPIESaKDcWv2kizd9i0Q1NBDbvv0MDoD+u91PQFRz3gZYajwHK/
Hwk3/uPgfHw/aw5jsciQBMa3c+aT3Xep1GAzZeJTKGFZ8a7kZLoKIBoZDQdMg8T1
nrssHytnI9QuKbjcTEN6Dr/DkqGjOw43s5MtH+EK6ItcCfQ6p9D6ZjdiRvpSqRPN
AN6Vv2O1QfjMZDTxVncrilPRsCrupDsFPlTcJ8pp9j7VAsrTDBAIQKGNEy/8p1XY
BTl58cuf+zUsD5BGD1h4IVM7EX8aGiTOJtVPC6dHtsKurJ1HimOqxah4AMmsZbmX
eMWBaCBaf/ZJW4z64N2gqL52Qe1mHWv9ZH4hqw0xvVYFXTQVTuWTGI2808zwdamx
b3KYpMlAY2hIUro27vEs5k1Dx+YB5Gb3fGWEDnTcdV0gm+sC/fLaatLpMh70LxL+
sUJuZeBjozA1E4ihugyI/JApTYEOmJP/nGLq3cAIb7N3caltCI8qkAeLdX8yb0pB
2r9aLHCxz4tQOKvd13B9qDM/hW8ceFJqcWGaFd2jAmNwbrQy4ac8+LwpggulLL6v
eOP/hWkc00Vswq/0HRDsllDQTtichKlKsiaYK62VSpOMV3j5cgZ2pmsinpdABjoL
rwNeJNdnCJqLmAA2FBOLaV/Sp2B9uUIhF5CSrFemXipOxV+ryynyze153IFqsRYn
U9GrSgir29O9Ka/Hh/B+CvvK/xeUtT+N5cfjhzJ/buoop+JZua3t7Rz3f4xsYfk1
7cF33sMtI7WZRCyV7/EQu/RfAUq59BVaJs7SVNtG4TRvDz1XvwFniWVKB/VFVu7a
oaEB5ntlG6R/3/aVgcCBZ82jW+CuF8pnLV3TYu/zxrLugzIhJodXyFWvwkLtT97L
iZQ51AMIIlG3Jp9q7a7hAngBHKM/Z8ConnC4eNUL8AmhxJ9fI0tdnKqV1xTcIrBP
F1IJK9D99mEeT6zTDoKtYnoCRHPy81+Tm5qAPBdFchu8JFXymNF5NLHFJlrtd3pe
wMAAFFgSKDF3SP7v+pwzjICmopijIVbnOlM2GDM/Y+4hu1O7h+MIPIJ2ql9avalp
ky04BGC8cCsDGfchH0m1Ehdr1WvAt/YaCRxClKZwDkvt8w+PwLBnINjeGBixLuQS
BC3jaKc/+R7y6VFzJZg6f8IARs7bwC5jnS7mUTLmAm5N2IinXTuF7T5gZZuNyMAr
tDuVwnHw9u5hfrL1wvGNULE3KkzX1hQ3FfofvS71SEBOKEf5Zlcll4517mx3WBMi
VkHHvM6MAlQ4eKfWRNGBA8octZfXpWQcK6BhMN7Upd3gn/UgfISc3GTWYEeifNB2
opHdPS5A7WcP5v8Yvrj56cQI/+NC/VlRLz4i/ZrksPHQ8Y9sldRPIZyOrRfU2H7q
eHpc+ecP2VyLIRJB+c2yPLZ6vvPPDgHpf2zHYfAL9P4PeobZ0c6hV+WOR4cKaG2s
+SQq2UWgCpsq9qNExjSWp4kaMtAxzcvv6vrhu0EL/I1vNyVgdnjHlEOdrqRybXvF
SdKXn8L1Mz+emavY/GUz+X8UzThUV88MNCDR17XCcmTfbAIgXJJQGEy7afkpFY6g
nN982VJmtTcTbv6EyJQ0N/VESmuPsw4c0NwI/3MF3yRSXdTaE9Rjf/w7F8mGR7D9
CPTUYkgPinan62al1O5U0WoGRYu1OLd4fxGcu2ThAQ6pjuWP16udclHWgWZ3Y8qO
/mp43aNOGAj7jjXJaZJHBwWFmFEXLSZpAPgDCkAlDAp53LSKu6dOJkdda9yR/eai
9A+rPUNeRNSUba1I5RhMoviDJq32DOs5BK1Ehk3dlp4MnwHTyozy1E/Tadneah25
0Ii22k6B9QV4LYW7jJ8U94c+miM8vUU/3BaYw1qU6t7U0HcH3lNu7neK2GBEH5q4
X34oYdsc/f0awtrAijOrR7AxtxVm7SRqV/KX0BNYYeeHLf8eTxWipg9ZPIXrdkEq
PmZi4G08Rhwj+tVk8UexSGPAz8UmM3ZOanZm7qWbfLmUAyAi+Zq+Ppj8nfcSUraC
zRdakhQnngUb3f2uAdo1M7TZjbhQkpajWFXgs7k2grQKzpuRIng6m7atDlPqkq2O
Spq8gV8L7zKkDF0iJSb+uM4bv6w+y7N/5EMmOMFYF/1No2Np6QOJ+RTuuIwl0kVR
VtZilVhA6VyxygFHna/5qrjtnGy8apji8x8Ej70M50WYd4S1CWnJCQGqDtwM4qcQ
N0T84meTnq1yD/YtpD5s7g1fiPWhpKzs93QKgLZQ6MDT+OzQZ3UgUDeUDBJyP/yw
jB0BH4gopjyY+Mc2Ec+XFGZR3SSloV6X11moA3Xbaoc1PH6qLxE4CCDWeBXXJKqE
8/hq/TiCinHZM0+35KKC6SDp8vcGHYfKU2q5HMxaxqtYbkco1ZXyvwChulgZg+ao
m3oksaXP8zutzs6uHcY2HJzBGIPYtqoSwv6n1Ck9NQLVsfzuzqwcu73rEpu8XL/L
+xlUA67TtYRw4C2eYelsN9QAMrU8Q55kMgvh0h73BrSZFXIjuam4TvDRDfyFm+/0
5vFUmDojLho6Qg9vcm9GootIDA1DX0pH/Oa3Ux7+x6LfoOESvzs7hFUVOP5uuI3k
OiRiRXPnjfdgy39FUUeQMOTCduxBqU2aIExWlYfqNlUuWF1csW5MiVnBl0HZKJw1
OZPJNZ7542L75Apk6P411Zq1H89stxQ1L27PIq4Gf5WdiTKZqmKTCI8vsK21YlI6
x2SUAAv6i0VfrnSx9zT0zK/ZwslyovjFrVjyiN1doAMrs2SPZLVzgs/b7nFTcoJq
81ddTWy/8ds/+yPr1tuql116xsWIvJXdm+hUiWEXiVQI88MAWNK229cZsGwhSPCn
3pfRVVosT51Vr87ecBDXExPGRqjo+2uqIX+ZCoGP6EkED7qPq2bMF++msOYjDXBl
drUPOwKnGyoz3eeHkS738ytQuJMUn87FBJRvD8/hvM8+zMto0yqpTWs1ZX6lAFRw
QuohQPaDRzLjxSXL+RpRutgwehiKtF/JNNfnk2gx0F9UhU/7K4t5G+1rH+Iy0YZj
otX3S/QlDGTTXN0M1+fJqaOH6p+kqwDI+XrDSeBWMMY2PLuH/yOhF22rfN4BgcFq
joyUIvNQG128rGQjgVltF7q/l/I17qiWfAwKIB95NcD/lIiqrE4UPe7j4KBZoMSf
xSGPXRkLWezos9+o6i5BIuB0CJnVIrjWf9cRxl3TcX5nrMVJl9HJHFdUfzl9gv41
7cOmvkceGbdzVZ9uOYl1KsAwy004wek2rRt6lCH3JFSt7uxegLaMj9E1VtFqo1AE
ONiiK4Je6HwuByWwttRTI1m9ryiTnV6LNFyMTpSfmReRXp5L1bE9c9i7v/JVMEc9
PV1UxaX1uSYUIe9dJxXcwgNdE9PGEe0ejjeLU3eenyko51yhugluTZEBMiu4kaOw
Dii/nTVqRuT7HV8qj+6zIbfl86wOZvrT0mm7/YT77kwBKJiA3jHCm48EerrYpVnO
VUi/tjE2ufi1YCld8Jllj5Sze9MMigSCTEKxQ7UBJW4ZLYyCQddVmcGHhYfaCSln
VbFbYdzpL+qgVsl8ejkirT0JdXF6CrZudJRr7BlV4/jxcbJKra8165OfmFhHvaz8
QBm9sYqz9jnEktPcZbRHuEFS9wOE2jAup860jtTtmfPp66yKrVtd/ghg2XJllBtG
kBj2mbdyZZuidYfVSndmY66ebhGkwnT9YIsaar9h/6izrPPGn+kzClG4cgfkhC76
Z4Vl5/zL0W/hVVY4S1mhdGUVbRcuGHhgg9kdFcgGAOvqg6XiB4V+6A1xBHTWzL8R
SM9wx0n4HDKzb3JMQjafliUuIQivdR6nl6HmGkSSs6ZENXOO1RQ0l0qyPyzDWUfP
ad0kppScBXEBcLbRmTyU7jxDdn9lXtVWJ6ef4k8To202sYcdudJv4YxoHy6wX34m
Xau/OaYl8hPDKnW4kM5jfPfSpXlTMOvQdvfu5CnqDlXyGzLBOSY55L62XZgTboUq
6saeREDuaNuCs7w4mqkc13lFOTdyEZSB+QPfy+rNBIlJCN2RF73pC3GLGRB8QPd+
yysTNF3JjccdZTjmIs0BFjluBxR5TId+FYQaeXzYKoF4dlZunWYTAZWkg12fl/hK
r+eVjmkLEU7sH6rYDXtOgETd3ZcLjFgqgk5H0/6KoE7hxs1x7k3/qOAoyZ0YsWtB
iSsCrHUMYQ+9+csrlLuAmPDp/Nk9OYRuTTJqByVuu/XVJEXDt1PNcDoVdqW68yW4
64I1FqOaqz0/SmHn/HbN/KQ+VgpFkH6Du3CAhiSb3c6oCoQxsbc+y3ciFT0wMxkd
Mq66d40AyPaFwVuh1WpN33dLL2jFYidEbSNDDeXmAPT/YNjicQZ0JDZmjfKDhhGo
sntwGWBihku5/CyudhrjBefOaW3C0lTD3cbzA7PIJTytbFhYapEloMtJN3QsmC/O
c8uFI4pnv2m94nlQgd7DU7WQbXUZhWT0Yl34eLwgNKfyoXFQrFQxGbtImc01TGWd
2EAcserR8209bf51BHzDhoyrvMpAU3pZS0FdgHVoQDiK5rFn2KD375sn0iTA6uY8
bCIGuFXb3Q4+555BPT8DuVuxEbPAuZKQ/+WDBMGYd6ecCBgFF78hdXHUjiuqfaLR
1gAQ/tTV1xHT2Sgljx851zwHHUupQfuk9nay9sdUGp6DpcXT4uehYFgiW5/C95cO
NP24OeQt73Y7O+BpmMJUSUmoCEgo6gPE+i5Av75S6bCPgLxUENbXM00wngUueLWo
u794kJztH185ul4EPQC7buTBbkQ28jH3kDQ51Du0eF4uNISBOyRmfada8mieKiie
5mNnct0q5xb279oDfqYpiFPRjvdlBH/0ybwr43oC8vkafjy/EnKIm4UbKOXN5wX3
VZbFgZl6CxZGKuoQYS9hRewtQtbVCdyZ5NL69JBRlONPMPAHl6KFuCFxF0TZCxJs
q8EGAIESqi4wXYQxnigiflndSjUSHKKAG+eIlpfrY8uHSjHgd7vTmW4FzQ9LS84x
47L05D5jgkhoWjQk6GJ3Zn79apscwOHRseFllyRxBaZWBxCwlGHhMEkXiDql6RQs
rRFtYF0ARIn4lIxbtX81gqhzmKAHwTRJt30cbSvy2C20XwawBTfwymlAV2bI1rAh
4MxShJXDwMqUuUA635uNaKzf2/V9ssJt5g2PsGbLEcLUp50pq27ZoKG3kCD7KugF
7iNTNAwOiv4czwMpYDRRQzvRbwbM5UvlJm0eUCc+5Y2kpicFSXUkmk7DT+9KVr91
acpdms9CSHAf6qR4rQy+BDRlOXVAxveRwu186j/qSRHi3eDzQoXElYOcVYG7+dtV
1yN+BsS/k7M6GT3Fl5ZijC4MxUl8c7xOG8PRYe8hYu56frnlxK615g/mWeKf5VDc
eAVn5zj22Ui3pexjVnSRwNfeLIxhgIK8rp/GaHHpa24sC2rrsejOSXMguRoBJ5Tj
B7LczpzdC2lDQlw5bmFdbobzJvZTigLrsOqfKt5fOwXEk5XyJ2AS/aTTPS+mS2k/
N6zKTw2QHYQc9OuOoBo79G5U/q5prFpcNVu6wCQ/408+j5VAq7q/3ecXxoKLLC/b
VJUvzDhZkyq07T9DzInZm1tOiNQJBnia0Wh64dBI7C2JWKBZ7s3+UBndLrYAgGY1
Oy4GiGSAMLKZBhXI8V19lFPvhkxvjKmrgDqqyurHw451MMha2RdG1no5Ql4WWp2I
k6nTStKqgkGM1O3cQYqCM7B9PKj26K4CRkmckSYW7VWxMZhL9yDTqLTpKu1H5OHo
JiEpYQtpXc8jNbnhDlroN5F6ADtgMZMZPRPpzT6XHUsxSaBJ8CIGAlVoYJS/OBAS
VgUqF/zMd8TOLcb/o4IAk0Ckmw+8I1y5CV2UlfvPzO6XouypfhlLRR+MoBdfvC4/
/HMW7MiB3PU/W+CseqIb6ALSHOW7JVfmKtK8kXN7xsSpgEsMgRrlZSbWZiKRhY1K
VR895D+2SRjexNfvfI8pJeCF8EyN59WDFargh9nImYNU1c1Uzunk6/iv6U5igj0/
z2ohMXo8el9X9TyIBhTu71j/vMUQKjn9NR75E9Tw7YSCO/8naJ610Zn6CCtMsT0E
WV75dKOyVFmqTDqCyGm6oZYHMxiGL6kSDl5Pptwk5sM91lF89QhRPuPI2gJ/qcjS
nw1V4yCDCA7dKkmIsCSRyDAX4/2nTe5c9lHd9tVmZ1ej9V6jn2L181CGx8vfetEf
VcaQJvKQiLndHOvc8r+nEyniv+u1rQ7CAasCajCEyX2J3BE0INu7xDd5qSCHc1Lc
vs+23I04Sk4Hw8fM9lUpIQASmxVTasPedGSwUP7FdjplYTd3ayJfNYzDMRpH9dSU
9atL/hJyDzIiTvWtFjPBZ4AynPi9UV+5zOUAuauocpK9QRdoWS4fjZx0G13xCoDy
JmHdMFI5klyYAYE90o7v5VUw7VJaAeLAE2uSpRVNgk0YgBETZ7NRNmRiKIlPNnGt
vqhSaE/1gPFgwtVz6pbOM4Z1UB5BtntwidElUlsy9oFuFxlg8veGs5NXFva+J+Fu
7VV3dZ54TH63XdjGXIdlJjZofS+BFNcera/q9l9qiweR0fS2tboBv5jvfC3H/SJq
O9sdbVuv1t9tg6iqiYXEAcNiZCb4ofKPuAEZIvvK/tb97UbC9hjsdqH2C+eAhE22
XDu3n9v/RZqOxAlD62iQtWU+GKTjWMTNQ4MJU2uVI6dIbUtzdNFDruhQAKDAWp/I
6cORtT9OavxG56vTLxhEJKI3yXtMQbOgwZDu0wN7M1HgqFQMTua+/kOkEyw1CaF0
KD6+be9AA8Ra56X62XUIMCiBAR8HL73jbBiyWzrOv5OGc59Se9is6OE84Nc39b/f
6JN9Sq3Ii2C+nL096NITIqhYy4BBYwxFSzrrSlJ62d4o9ykTm90SJAhSTLy7feNF
o5XwSxQ1vefick4hOzEbadkbzuIUK4VvtjzJVfaw6AG8Xitv8Whs7R+8W9cUbaPo
InSuQlu3lL+yix+hp5HNcpWRTl2wnw3M+v/PYXvtwHe9yj6pxFtQ/8k0Of66ut3G
YIfpT208WcFN3RS3jukRBqgEVUtSvg11dWVkBOkgroGtW4XZjfXov3GkJt/pJKGR
BITrkt68Cmzl6ATQ/VM1BCFL/jpun5vZCEYHEDmkVm7/wgumMsow9dZkdp3vwb33
CeqbU5IsLRwP+J+TfdNk0x25V1GycFgguoT1WZVGq05eIG68SJfptBxTJkXs4R7s
9JTNrWcVfsDW3KpjXwSXElyOy07mR/MegYwzyT5DxQPnajAsRixVloj8ZV6BZYcs
VKcYKYxH3lThtf3A11kHy3OnCA2hbBdQc+dUkuIlqYnTVZeviSyfvInwYpw8ob6F
CjQzVYm34YnRovOG3wqAmLQ3HkVa7qmHm6jQy/nSwYWXsdgoT/VZpjhVO0rSHoGn
y1pvIfN+4wer0USLWw+s1lOeF3GTkU805gRaCQoOwoRHN0g5yMEbcxBKey7F7KM5
uJNH1X4cHTNT4aQU3hOCI4b1Ne/0cXFgYmajoWdERXDBcKhM0Dt4+EI/ntYI5Bkv
ZXaLvK4R0/VLNcKxOavRnyM6m04dpcAd7duppESxS+K+ryYU5vZ88Om+u3S94OVP
yNN0q2hDWxnGk6tIQwgwfrgmqYfBFR1AakRC5N1FLddGPo33hVprAzwqGw68uBNA
W8okEjRv2njJsYoHSEdktII0RASxnorNjZuHSnbPZJPBNwEvU90TgNTMgxtcWA3Y
ddVN1fS+fjcgQss5OnsSZI4HTOJSykpFVhEjnT0g8LMt6P/zKdf5bQHen0XqZyZZ
LexHw8YJ5sYYbJQqFu1JZJKLIpMD+at62+KpLk+qCWYNCSdR/c+DVWBj5l1QlWk7
pf2vUYeXTiizNC5H65PiQI+OBjsVfDR0Z6dj6eHTae+266PL2elKHKGzdwo23rQO
FbjPyl7FNRmcTCcEEoevc2JGseHG/rk9sMprEv+357uvnjrNcvYez+yUrgtQ3V14
Mk00Pa0bZEtvqiub5sgHxFXgw6LkG38KPaR0jklBR4Bx48mHW5aVv4GCoHnSQO1c
ypXUD50swcoCVSENjjjDrIjKUgCi2knuI7mwFffYoDJEMwz8f4BP1rZWUCjPvADN
m+oqBz/rFWWsXgmNU3SkVBqlB06fGzKx6EiHRrkaXpy8jMSdGVNy9eMltsUPKOH4
3s/on+aDygQJIthOLVK6lldHINSKEYziuhyWSU3ACmPr9kChxiqR7svvElcUtmD3
twSbunvRiZOtEkxqy3b4j5WVtTPkimcMzCPa9fBVNp2WDD+cgVTo9SgBSUnl73QI
CeTZ5a2u62ws81WAOq88YRQ1NITBsrteEfurClFyQdcmsaRZIHertkc/YjhG3S7Y
9JlHtYFJ7q8k3GwOo9jimfXJZn+D5BVoBK4Q30qHIhC5AAmOeTzIpKdnxyOTocgW
atdJtxUr8YUc9ZvDFxI9N6WWfNvNxqph2mR4J33qMPSJWpBiWwl/fdK4u0xllOXO
oVDgPHNwubggdMpHVUcuFkq/Sv10fH8vJ/u0lHPdMvB7GVggkuQ3PLosHOpcobJW
RRN5VTNfA8ejfVWK4OFW7JL/QyIdSMFIVw10M3HhRx2NRcEkAIEWxM2M1N6bdckO
hGqDYPKtRcIsKUWUTr3O+DLNUehUrzm3JiZLrO0LNL+eZVrBt/79WvOsdnmLc92L
x28FepWCB6DvHPrwpBFDCNAGBgmAD9y/aT3LTT4PQs4XLOjfAhrUPB7Z/VcM3a5K
VE6wW0Akz8xFAYh2pEcBeJvJxcal/WrKBa8ZFcmCm9G2j5ROS/KkKAkxRWazxdtl
pH+V2lJ6n+sdRqwj3PvCz6m5OJl4B6yeMfSBFtiRt830eyOTRQe3Y3EcO0kTYCqR
TG4MeHy/R6aiczYY4f/8iEXM+81HSl/AmHeH5PjW+dXZwKLnr3DBfuLNqtclEYSq
MqydFJlNjWkzIiqsoj6FRKUSQD4edyuOTpxkHHuN4+d20TIyLWnPajFeGRX6p2qj
3H0M2EzQksE42wFu2VMTjWAg2dpbl+0Fo++GNJHyG4YIkqycGXNCFozyeLhdcVyF
1joABYpFW8dI6BcQBY3R/FPSEd4mOUGsiejfIDXRXUkxmPcQ1KUYjQLnlTwFrKdN
Bl9PWtq1t9jkMjrzL4endZEqovoaoxD9lLyRD7ZZR5aGnR+rJLZqXegDmimKUROM
fttS4rO7jKaojU6NHmR5WOrw3ucVzCX4xuXPmaYfdSlkpooAyPe3bAK5jWykqnIv
bf+9IIcTqGlG6hzGUvoknh+YSmSLhGDTQW1hcD6R1bJV6jzmgyrrMyWSJlSP+zrQ
E/sNbKjuDDfX3pQfxe25UTyoHWrKPTKwEIfngVPCyKGBWloUbs4bZc2WsNX7x0Qq
h3Hz0GhcsPfH4uC0zVjnhS+w0C3tu1v3kUNGlVodPRgBFiqPM6KC762kVkmOIl8P
eQSEri3IIPT4VsnR+rniv4iix696w12YxnHUvmqLSpUuIkVcNcRQXvipwYx3vsoM
6ravIyaMEOdoJpeWixnTqIuR511evKsLZW2LLypNS3d+aPY6pCrZmymkXnF0qNLz
ah82jX+gUZS8zYJDIN+WdovLBijIlDBFJAvBSYR1P3U7wCh7yaAadIO/k8GvfYvS
T5aLZ5K9xgG42fJw1+vHsEA+saQO2osA0iLnQInkXeBblfFM79jCbjbwCDp/FYp9
uXpBgz7hbJLIBQO/DUFKaRTrWAXeWlRp2QJng2kdk8hlHPjCRqqSRfMbq9AjxMe7
wO9xTELTchZiB+zifdDTTEFgDj+KpOJ3zBwpyZZ4aZqvOf6le2zKhfciP5p3vXuU
ryjd5YpZglqan+Vk9rzB6iYkOOtp9DfnZ2Oov8DGrY24OX1BDZr29Z58Ojvjer3F
688KzPN4AbZ3YvHQucS4rtwl+3wDtBhKBtQq40ywXAJB0G8fxsTl46DBpEYNo4V/
Wnw0zVIZxKa1lK0yBLOmtUPyTFNneoki//0JUAIscxN/wjVOn7oXoHI/nSEscz9K
Y7IwtiPCgm5vxZv5AS5sFh1Q+iona78+wkp1pL+44N6riXhl5H3AROJmrQsNKLpl
jsBLsu0qwYtaLSL3Qx/ov6saUYA79Jn5/NS1psYT3QKoQzUl4+V/ErRwGfEJIseO
cXux6w54hfmWt61bC+iDT2+uqDPbiwuJhlPEDQdza/6pHLYNH+pxz7XercyGtcey
+OAzAMjl1kBqdE5mdZNM2gZZTL85LqJEI5kNWubYnlcDKPyjo29VLM5AkXxbfUOM
Ue8aUVie7hqL/06ESZcU0Vi1E0rQv0TAJwACsxUcNT13yqNCPbwMtQNWKHYl2uns
QeVqjvTwtO7/+sj4C00dTtukq1ZEHhZr+RaXIAu8vbNrnb03P5HsV75rLwYw5/q0
rf9feiDtel3oF9GFfBhl93Cx6hQiFdV8m2i/0l5PBM3KC0M7hpvhyp0Ney/u64rY
XBjs7JAtAxyb2Tx7h/aQKQ4D5xY2412wioCuiylJxc0QgsV/z/EHmbB43nv1ZjXD
MO/8vYmwQPGN7raf3RSvG++s4vZN+Lwi30tF3rEYMZiGJnb4Wd2x6eAZfolyZoI0
Fw0NlBFgivYg+XM0xQ8O+eVMtZ+QzrYGMs/Ffr73QLXbQjcKcOvJ26WROYquV8Fx
XGhsicqnJfxClf7cQeKA7GEaDcYyYSEWMYpNpW1k1QrUUSdRvPcth+4ity5lnPeO
zymYvyxKcUpQSLLnqoE84g+5MOrz6Tm8P40BWQp7UrtZ2aPLiih2MRI3mWQ8sGdA
lOJRlHxqbqQsiBqurx6p2S2t9Ps0goHbHOaXwzX+jO/V9xhHHQ6iBzVPYAf8WMLS
vcy7GgsoY4iUfdTqNRu6AuPhUb32a7NCBshwtjMTmdv3BK3Cu+Havc4ak0Y1TgAk
oRxKl7vBrxSJfdT/nxlM6IxUtvwlyhSE4UdblH9Y4f7aHLRVH3FWdiyaUKZBNdNN
j8sbv6B623dVcDYn9QeS8aqUG42Goa0ZwzXsulbHQdIUGCgL0PjZYtRZPxhhQd/g
gUJvfVr7tHF05aOnRN1kj6J4bMfGNMN234v3W4te+NUo/YE/KPNy6kque1J6F7tV
7KcZ4HW6ZFbxKEk3ktUHj0re6TOgxfDZfBcpK6G5D1g6GC/w7CIvkvmF889Yh3ld
cyv+YitK+5ltCkDzWlYVMi3af46fG+PwvNpsWvgTKX9T0xFRt5SmwPCCMK95X0y7
w1IBufuIv1el6hylF75FG+k5xKLWJabqotA7FOjFSS9hDReuF7DNEaY/4EVnebPX
BK35RACcFCV+r00bHNndDYMWnkCpLKyN5FpbIjtpNK4JPjoxaa6dz0TNAxf8T6iw
1rXulg3WqBCAarw/YK0+HoR9yWU+8pbzxH3QN+lUmMKe5TQxfVi6fjp2/5Uikzmh
ARI3bYgaNAV4BzT5q9hTW+bEDVra84A8puM3mkXWB2L3hLh8xNVLqooVoCLIWcle
Dk6zwlq0xY19kjWhN48nYmeQbl5uiILHqENEcdu9IYXx2tnJf7si1yApHUyqvRg7
oyld9+CMCIf9eHXmFasJFMX/In7cg93J1v4M44c2rAGyZ4Y7jMQpDtADbH1G/DWk
Zpf7S6kvnT5h3TCSeBEK7a6RtvN/lAo7U5Us4+M1/vpMiXghIsl6LpZqvVU/aoQO
9YDJsbpcRWr0NtoXziz9TtjPe1wqAL/Se17me3X9/T6fG2Wq+YYit06buZcqdZUO
a/p7l+/yQZsX+ZTTnP05giggR8ALU714B6y+qxotJI0cjmvVYEMGfVd9SG18pkg+
csw1sJjbAfrOcLha580hJFThz2IQJRaaB8hJWkP59hQGfyL6N2WmWxHhdvQpbKLm
26z1ZObU6hbKntVmoOlxlp3JDdHBV/exSRNDZ4zm1rf6XeHMg14jLRJpi04uIrtE
fVC2qNeeE1DF2GnjQF+j69imzFbtRAt4SaLoRcnPzuzwuWiQAHYKvEx7f8blWpVI
3eUNzFhFgUsveLQMN+pJQead0wbeMtsSVENeYiMatFAPNDNX5B2UoieSrTaxqyhx
wZok8gODJ5B1Qd49eJu15FhPXyiZUiw99U4L4oN7nbWKuFh/WsykigR0iM4wirmJ
PwPcr5AiEnyaPCosywQGBHB+ly3tVV4xvO1R1YXJQMVHgbXKoecfQrzNqWLynv+m
WsqfftK09NNo/expyQPTbJquAXVYVer947eulz74Mpz/EQW57PnrQbpyWiJgpulu
2RwMlewjjnC5K09KhNhQ28n2OGaV2kaiZ3POxWz44J5oY3gSRo8HGWfXsqLOLOSk
7CcQuHWe05MgwVqWTPowidDim1+DlCEY7DpLKHQZqnwxRg40zjMZML+Gmoba337y
QeOXyf9R9Q2LlwF//EiwDbtMQUiu5hZFgyPuXdmWhNjP+LLWmkAl8vsycHYwDTmI
EFFyuIud82psFyrqI3o/1zrME9LbtFlH2vmAGpMlBepZ+Lk3jRIUFL6uf4jUCY6r
dufbh6wqypuuwLp/KCPF7k2YxxYWYASQrc6ZRDdutKmK1URbkbzR2SPb0QYa7BvI
rergZA3gCgN4d1fmj7aRfqH3gkZlmUCAEjJpdUAbSZARX0qW8mHsfsZR5KFTmVfw
aba8Bck4Df4E12Q9lnd2h/hG1C+3Yjoz0Xp3hgTOe0hNaHqZOBzUDpVaIpJjcQ5Z
Oz4vyLiVsFl9abr/1ufEHRCWSdiSpFlu4hgWPuuyrCnv5V+zMIC5hB+zywvuEV/p
2eO35ShjCkOuUS0Nu0fwb8gaXdK7+vBPIb235QtHyTd3G4nmSt+RpxmiPJmb7Ft3
jEinHANf+jpJdpEGrfFjO+CNXKkIMfaTrSuumaAhbxJSOxWog6MyOMUoXAFky3nw
gf6vSFD4fimyQnEe8SX6B+3PNojcFxSQCWb0/FhHM0Kw26PlnjEI7sy7rsldgunW
mipGJkOntIzD7G+0V1LDXMk4sXnRPvPN+31ZhxpAu1EHQ/jZofObJGgu7FR238IK
+RvtqR6EGCAZMci9ipmu2YWu1j9UI7HO34p1Njoepm5GVDGMgQXLQlEo8IALr0P/
xArlMDkL7mSNnqahMmw49/5tEuigJmceC3job920HjhsigeIiW3ioC4P9/zm4322
+rk1TK9POQAj/7FNzX2sySH6deIc9AjLLiBRlrUNzSciFOBWnIMs0JpQRKHHLGwI
HZ5VzDuE0ROLC0RNuBs4bfC9EhJkesHAY6eR1/zomOGynMJ6nnEcDy87YR6/0mdY
fC3BatQaKuLr5xBx6C4ZykJjLYx0SbQVI+71wrq3CpXKFdc/i8Zj0oToYj4jVshs
AhdTRrMF/MWpr2aBk2riXkm3CDw8XgERmP9KTHa7SLUeAnqBrnAiWVjYkuC26NLD
rKkoa50XPuh0fEgh0tpS6ey+DATUSvbUjTTinj5xoVAj2jiiW9tgOlr/Rf3aCpv5
RqjV5XbM8cVo5Uj1JZmiH0Nuafk6M/Q6fNNSA0Eh1CejdcWzuTUwEcYk5EzvoZtx
3WLQShp/yewWST6kjxDXxJDsQs0n560+TZNOF7zC16SdwnzNSx9nDjMSzr3yGIom
07l+Q9Csjr1rKfxWNhnGgzxP7+M+xKC5ivh4iFsVOAMZ2vbGP80OOK62jCMonxMc
TWVnHRlevNdBaokkJh4UUN39yhRV3IWiDsxJ8ubE7mUgd4oAF8UX6SWcPyjl7wAc
rT1Qf9JBvMlEhD6E7AbNV770rEzAH7NFTE0ZURaSY3+GDHrRnZEx2mzXxvDGMiOV
YXdGMpRKTsfEcF+ZgwapR06qPRVoQQ+rK7zTjeqNZv5Q7bvvcDH7PlfEq8VsopoF
Bm9duYDfe8eFemdgOUEPaNj3f1Sycdz+VzZVmS22vSwwVz1zlo9IbPcPaaGsV4Eg
apLuWViz/ROdwd3l89gfqI8YB0MJmpidodWJGBvYvEWA1oG/rI7TNdWy/wcoio+O
I/G0k0F3O3ew55uhff2QegK0BdhganojHXCjz6YE7FPyoSWiptUWXYIp3KaE0rjG
9gbXc/W1KBlVgw6a/AK62XixA3s9h2OWNjCprM1lbHSnQ82lnEsoODJJsT0LWuS7
UeqVdZJB2M+Usa8uNy1i120Wpux1J2nHFhJJqj0gXGIYqsDuK7BvV8uxykd1V3u7
EusLSiXdDclS8iKT++0OqnhbptIJ1XjA6wjfjBOWu92YCUKJiSq6sMpcCpQ4Gzxb
YVo1RTI8twzTe1xh7eCbG682A+e/Q5zR1spnYdvgmWmMHuk3M2O4xqdW3gMPH83m
JEGWN2CuANPAa0TaD0bKvZzhxYTLkcHlq7PcZs5UCnpGa80hWt3BrlkghugDHtkY
9fsDxXSGfUwjaHUtBjNTtcv12nHIrXmfZ7bpTcZrDuejoRonBkq1tqY1knP317mj
MWh1rFSKD4YX2KE6Tt3qdNCO8OQTEYUABsDKSDUkrVwP28zZ+DdhPNdkRDGmTpOc
U1B+NwJ8ufwHxY+dum2KGvU5ko+tvQIo6s9k2XU3kZ+EBF/VkK0pO+zJy/0RDGUp
XVrG627Rsln8PugyZrwcZtFSqyW6XZvlmNILfQblaCLZhGJqRBkmDAA6eq0fknU9
gl5GFWH6ok1PLTw06A1xnj8B2ZEB7Ttt59fW7wSVOV7yEHq1pGjdukbTEb1d+9bo
vIrKsYKtI7+HGi7ZDz3cBwgUsj6GdyNse/x+y4boyca4+kve5GHKRu2AO21DIIKR
6II6ieBFHoTJikWQei6fyyVovtAogFBOUOVw+4LuNpMhFeOQlQk+IDnCNu1i2KnW
U/CvszkIlehXzPw7VC3vR6D3KQL+6jZ5qcW+IjJs2uyaL1pVpHiPGR+wvL0KkZ9C
4Va9q7tuyv7Dy8ptKsldFOQNg5rJeoYZyaDZrCrdTTdnIddwJ7ZXCO6j4wkKwPoT
v4+EOtIjM+3vrDVB5PiBDIk6KyzPhntc8d+dFX6VKM4zG7ydGiV+88BOKxUiSf1T
mw95iWKzJEhZqtnuSKN/n1kyfN5rRgxzpiSqW1+QCPkPTEBfFthV0iLNTazX+dIH
HBz92IBa7W8fS40TmHsqHW2fSQ6PBO8HgXvlPgICGHLEx0O/b5DUSY5IlBcE6WXF
nsqTfM4RSjVYrDXKcMPsT3baO/H1UYw0If0GiCYOaid08qwoSL8jBPyYV1D+0wT+
UoVsJfkIM1yA+iSRq6o5/G+KGNd3qy+4tkow9/t2PnJWz9voZct0keeKYNYuqAv/
B3TFc9nNju7YLoNvB5xnqfMZZ9SPlGt5N6njyJsOGx/1RUFETO/jDWi6jDm7LC7o
qchBDkNlVoOHzA/3l6hU09khtHNphxpoG6YVyyVrNykzFlkYaFkruUwZAf9WslYX
IKKzHzOR9DUPtWZ2/rxfjXXA2EiqiS6hanfuED103q2e2Zi2WCIQSBLPool+hrrB
mTOGwGPuGfxp9eN6FYfJ6nRUGqWGldwRK82AXeL9+zLlcknr3l46temR68z/oYOC
nTE6219+Te7c4lTihxHACO4finn1TudEhtqk3YAEpe9DltkmR7xaP7ImWKmW611G
KjAJ4wl3UXOle8dSWTCXMVST3d/t8HfNdPmTHRAw1jIlf/dog5+2y/4ZUdrv7cux
N4PByZHheDHsxSXEvvtupQxX0+Q/7/u94P0o0BdBYRRWFv7FVqsw+40UcNrdc+r+
NpqN1r0U44X1rCUmwPUTp24psXle9nvXMgjkYNww3WepHQJQd2CgJ2xBxn6coxyX
2hmLt9L2kRberenwF9CfXZlLNvggS/Xc8Vj4HPWpA0+AUcR3FjJNsFrWxT5DrEPy
Hy1N6hJ3Vc8dN7mrHRoMWujjAjCIllwiMMC1jYPG0bLcSHmeig4kVg+imfx+SyU8
1G7BQOM7P6jpO7iWJ3Rj2KOHexDTi6USBnpvSJMJoG5Lyts4nfmvqpxm2mOkyov2
tWUyYY9yEFnl5WgZfimWYyDg5wghnF5e3Gp4i7Vm/N233mLeCPeYmKCabw4HQkd0
sK4qG/3EGsUYk3mQAE8ebOPvxbo0T1HRbLV1FNZnTnd3GeOwBK919RuTFxLDNzs5
0RNiXHBVYLFrDJowIVNlnxIVYG5P1VkHYQnyJqJCSuhva0h1h54JnzfTLk6/fxFo
3SuBY7/Fyfc5MfM4e2ucAKD/p2x4dHwJBQU+Qkp27BQ1ZKkSfNdHiYQ7DUTp7q61
/YuuupjyYNttDY8fmqybP56AUolqLubwU6CDimJrypZ5hHzFWe2Rc+kgT/6qKMWg
yuqFDOed78zqsvAW6Xb5Bkz2RhiVGr+AilrgT4rNd7Fz/1tCW9i+yF+NcSyWLv++
vVh/GLIiIWmlisJbx0bMOxacm0RKLG7sWqGIypC9sbLXiPMLM/Z4q8E0jGKnMndd
PhraNQaS6rPg8a/eEHntKa9MXfNf11dqbl2zmVUJqpQqzO2cvQvCptnGM6lWxI8P
ZqUng4m0eArEjv4DZVC8+K4VJT/cGICRLjy3VSL9Z4oqVnGUCJeFeVbiyjd7BYDa
5vLK4zsRJvIGqm5aU8SkIcZTuTWNJeWT16SGn8TKDTtLtygPMQpT5ccYt+VFgMXI
k8fTj7jkX0DYeXUBjECtJYPTZh0pEoYgYsmiZRGkmiqYSjR7tRnAEatJq+ikw5hF
pHWXnGWFhPKbe46Dfsz5It1Gj9HZxRIzgKOnPQI7RazRbkrl3G2OmtPrcf41IQ4k
8h74qVeIpcQtZh1IdX040I0PycHBNCUUJ48RNpcO+pgPDiGSqCHmz8sTsoM20iqf
HXux12w/OmdUEF9sVIVJhve4LLcjXPnrxbpjtLatsBgkusoaM9DHq9l5sKjc5zYH
m5IsuUyxEeihB+WsTzB9dvjKsrfVKPEiilLp2unlidjy7kNdiuKuAe0qNXnZfKoH
+Vqfref3ln0Uq9u3DiJHd9Zpy/tId6JFydbe0npj9bH8kGZhqxTLLks/jgRYUVZo
Arxzf8YFlm9GxzPXk2aKP8aBCy7j4zqxshUHe/S1E+cR3eGZfWkqNJiMks1SOoWi
kMBxoA0T3PZiFmav5LmiHCwIP30AIzN/hDJ0n6AS7HvBfY30m9w9qRWO6oxfFnED
db0UXq8dAz5FQ8RcRQduQ7lg0rNxqwAOHeXMwAwbRgOfKGbn7vMw7eTCOmMgesRq
Jq20GTHutSVkiKufznqEFfNUhcHlZpEykIbU6RrNYKqdfo03FCurAKulzjkQQ0cP
65aLY6eysSMvqsYBuxZYktsA/N73OuETnXPZNDN/F8NVHiRZzeR2ziN9w0oxnjAC
60DPIgFpNmhHF2H/NnCctKK7zcwp6WoQu1Eb1tf/DlYW38cyTtRfCNzqk7BaONMa
x54xjEboawWhc5npa+G0l1ytTKzoEoOBA16jofqKRrtcVYLNc263DtYDEgBzPnVN
z5CjvUCUKoDnYXwRAVtpNiwpjKpGvTa6lPwriINYN5dFAFzX/I3bFZq4rtPtInJx
CGTzvToN0TSwuxfNUYWIJrcx7rkDa1dBhVSttEpevtLtU/CT9Pryu1NfKk1EWSdR
5O6Aa4+ytcxsx+scrYuLZhBDA8/xB58U5HktzmtshAjj2hV3jSdYZzejQeRWS6p3
dTnEqkK0XGNbIUdntSXWg2U0ghuZp/bCjM1nV4733oStDn6OctmCK89hXACetomF
Cab42Jso7KNjQXsyceJFtzMnpQSyTbsKsnWv179fToCfPG/ijsgPx1UB7Mlky38n
h1RiD6TY4+xCGlughKUkKMT7EEWzJd8DjAh9Xe/JzbJUlpZ8wXT5jOiV1O3EwnXl
+gvI67/wP/Q9nQPnhqJxlxZBJCK2EXzHWnpTVMe01Myt4FRwydA4nHKkM0qqp8Tv
CYGK9jd55k6Hns/XyTKYckM8Ja5JdE76vw1VUTkvE98/h/PgjgO2t/8JNWi8MLn7
R7AYjMFD3avFa1XFB2UQ9ohtxVC9TzRW5oU1M4oTNClHYXltTfCUjEQusgzUjKDI
fxpJ58oTaV+thb/Hh2Q6sDObLW51lz/GZ8rcnpOM5OxkjfhP/AysDbfHiNZpyurF
MDxu8J6ghfbfgWrKK1sEbXg5A8JpCPZ1IY+r6xmRC6X1IQdQrRRhF16e6Xx1+aXS
+zBG0pfP4VWFfJIPWIJjxlbHyRhRcPwe57iQRhZaDZD5z/1sy/6dQXhoJAhcPL67
KG4vGR1eFK+rm/CT/hJkcDcSNfsv+Q/p4ivrq0qz4NTnemw673Ec8jZVs+8UlRsg
HjNpkQqPJjnEUQ8mdVXss/y6BOfnOPqpMN6qx/UeOKR+v2uZD9kdpjXf+quOJLBD
nNJGaAHJjOQg9kUL3LQFmFgcT+MwXrGXvf5Aljsj3nIxB5KWIYHCETvtWjQV7wRb
GKsaWrtFysPMZ+SisTJETzEgt+RwC2419Ngy2AtUh4dDvaA+n0nb74yCIc/joZPK
hS0ISCF53PSl1CmMZSEHSILOaqLhEfglDuaw1mYxuBAMbd0RmSruqG43GBpofYSG
YQPU+2BZfJlZYD+XIFkqQuIiQ7zNjJE7vnlbQTbGACcMOV8IrNg6siQsTPlikFKP
EybUMOnnvDnA8psO3RYgdT1PosJIQSAuA7mAkaWKRJQXfwOElWBQPF1nO1kVqwGZ
q8AEnSPHF6bO6wGXdzYJp1/hWjyRpFnBiZEef1oA+JhGIknj0b6WHx5ybQMEXNhd
JAyLUs+4cuyH+/+VthbQswjVj3zXVH0IChk6/6T4gkMF+MHv7hjgu7WWf0vcw6F2
ecZaatQcIr39zqs9++aTchQuZmOdCa51+Ok9AlG1FD9zqVPA149GPGZAk072Tt6P
Ok9n2vvOHVbKaZRv37kGUq/PuxHkB3hXXThWhMspyERoOHFhXu/XNlIpQrSyu/Kn
5ZCmgaFWYtYSYjNQ+hjWCCWCLOshbZoCu3Mn5iT/06Oj/LaTi8d3BF1EriYMvB+T
CCfyjUTgdsTS8rDFMKSNiS8o67C3H5s6ykusy273lOeG3wy1sSiGdZ3FKyCS4Jup
EBikJO/Tp4/NX92HEUCgfWrh17zqd3l8aBXZX7xIuG9cClGavtHXh3duK25hPP8L
qgAWHgEnrUSMR0Z2qSCWV40D+7c0a4RxTTY71DLYcVpp+EoOuFvrYomh1SHI3pjM
QX+IHnuKcAO/TWOUO+9igbm6KqPYRe0Be1qU2DfOxTLZ+w0pNBndlHIggerHFhIe
mwhynqi3NhLU9XbdCfmy4J97Q66j+/8AALEWBXkJDNpS+zYvEWWCB8Nu3ZAxOMh6
ilnscQ0y05NcKNDlBNnhK6jyiUHkIAR16K9+pHsG90ZDi1HBGpCYF0H9q9d003/3
ESCVRpDcnEstZVzPXLRoSiUxxDFkpjzFjQNwBildGpz8SHezElIUkuqXor/yaRQX
IplfhOALZkNtDvyTmANJd7wtIrvqfnNZrVe+S/zVcZ8vL626iPgzXrYWnN8JuIHT
OzzmP1h5Dmw+sugormgDYXepPRVhQ7/dOdiXBaXflS5pzOmm0BBOx7xveMJplGE0
/rv47b4OHZy+scXvYT6eTBbiZP8arEtRCHTcdwJ7c/GlM8q6UtQ4SJciyXg871uD
bPmGhcqlWwe8m9LEkRXcGNIAay5MyF16hcnZbxEugmhb9P5dIraSRjV7ZeTe8Ar6
ZTUY98nmiMCV0zzJnP8owv79KHVUZhV3I1bTm6ZVe/6mxykBRdYV8qKmDFMu7YG2
1uLWa0QDsybPgBLYMQEc+btpzrdn9xvgBmx32Ja3EVcz12zsXfuVA98D5StREm16
P+fWyPO7CUlOWuNJsbiB8aavChDscE7l1WGNeRDCeF6Mqx8NpZiK7xLleH1FIQxd
5AfmkI9WeJlFXKlziM8EzGFwPNfBtEGqK/8ZY98DTamCPvJzZeRGLqMD6dzI8Vis
whEfuFyCkrdQhcKtghohHWp727otk+VUw3aopa1gpBNUEX7mV+OxIfpr4xjTDYBD
67tUZRe7JtGGkIcWnATak0lGJVDDakuhRPdvgNnDxZesQlqVLlkvcbleD10cNDF1
mUMIkoy0TXPVXM7RFpsb94ejYKhD3+sdJN1bTAN7iMz11QR036+KKY5490VWgr2g
3xgsD7wDGQzV08h41ClKbdXU39gAAnBfOPQe32pQ6KCDk/3e5IUTapvTHvdoetZe
G6V9ipRmOdWzWH/4AXtczZmMzXju1qCxhHSYBEo+RH24rCL8nECkLwnmBGyH0tUn
WvviGEqlk609ry/WyuFnq2qJgAnnRB6qM4sXOptfcxgB/TnsLChZTllVBQSzaHCM
EjsIKiIHXHyPXXNpsXivT9onqNZlU6Da1bq7CLrPqvz0HOJ86xMEXGpSWVJSfKcY
oL86qSd85I7i/4GwzqgMGBaAqfoq3d/57kjw9qUktzQLt5aH+9V3q5yRdiOqFfpV
dpOAcXIIy05q3o+7A5W+edhZigjbWaOwOMjfTqlMx2DpFZHvCpOavG+RuhbWdDDM
7Jm/nEO2BqbZMmGxNQCYqFtUpTLurPoe+/5A0GdrZZQN3Lzbo8UDW1hXOYiHvzIi
2KdmJ/SOTpilvl7EFVqtvBNqxhpwE9fwAakSqB4dchHuIdehu0ZxjedlmH4qDKXo
eVdWxp+MA+F60sK9X+ARcsy3+CufjbcPhb+0QPk5VCPvTqKNb5ILzor8IxPSJFx2
1nnBmkhXhYV+bhOjqIYaJ/yhxI3IHUphycqRiwCKVVK2aPtdVFQH2DgDCqNGWnV/
/1bxiSICMh+fUFO72bcEm2szgVYuYRVCPizKnTEbzw9xdj9U6YzQD6mceYwtQ21n
8GMLIHr82J5lCv1XLges40Igai+Yq0VeWDLHFQgllkUKTtE1Z0HD437pND7xi9qz
SSxc3BZGGPWdXhdH/yngtVjTpBJ2PvEOi4SPXUW4uFSa9bO6xfYl5MjHIkHHsEaL
fq2qxmu+8N39SCi8FhaVVak+JhNmHeXa6GqEhpkFvLEjT3jPOWbjQPENmxBKTKlh
/SSJ16+pu02sn4rQI0VVzsLvD1osRWMQvp4ELVv7fygZNXIduvXCyK5sxmVPtQT0
UKoNhbmdN9zKbH+DIcmzIvkrL5HQSej1xJnb3lLhPHB4/Pn1SNKiJjl+UCcv79wx
BB9JY3xzWT17ovTD4tgTlL22PPQX6nvZT9vRr0gDJHGICu2sj/2tGm6JYK1GfsiL
bA+7jATGofZET91d2Ff6dcFWqbPDfBn8jTlMILbpzTnT2d0cApSYICv+Mo6w0EcP
O74D0JfisaMnDUW+3h/QZNq3VfwhvK8mZ/LeLbmQZG+r/F5sZdJcxlAvIRXn9DcA
lL0spfCQYJAVcAX13sl6dcecbqQ50L+swckgCfaW64+elThCDwMzulNSzUb6aUgg
XtXTjVhh3gAO4BA8ovRVXJRNRvnqdF7JLxqDhrWN15/OsFiW4EmwTHcsTb8KFFXC
AHiSvtxfvrLBzXPYtFMZR6+bkUgDcPLfTEzp0wD22UjBMe8UDySRJLMSU0j1qQLt
X1a8e1NdB9iZSwWmayAkoCV+/JjeH9AyIZv40Q6jqLtz8eT7IO6uFy0GrcDbJuLf
X7AI9vtUKKyj8JPfC1W8XtAhBxQzUBBPrilCBSeOJC0e4Vwdd7//F7pCSbxwswBJ
IHqtJjZBC5l2ZKk361DdRji5/7IvQMHtARY6a96H/wdnt/13qkI8VeSZzCvs0r5k
1X7pDNK1kHF5D4l28tlsFZvBr7qpeyph4buZCuDLiipiV+qfbHLcF8L2apETe09X
898uzB9CAW8GeYSezflPB1oaWIpATp7VyqrWbyoXz+u6fQdhHvVyqQ3lNW1ztsSX
9jZ7EZbhRMuL8kYHEfnEsCYHvYOOzERkeLJNbuIJX1/RpfORQFbnxB32aylsiaKk
NF9Fs/PgZ0geyWVcvaF9cNIM8PZAG9W4j4184P2Ap7bqVW3meQUxNIAHWI+iynC5
5KtbTlmecLiDMZTmikS3pd7aK0iPuRwqRxNmiJ5MM+ovOGywtpss5V0m5MHw5FA7
5rE08JVmjh38zUWM3nRiJJU1X462OlYK35+OMJ5L1EgqtB+CiznD/4W5fKU3Rth6
VoTrttxTjC50r7uvAECJsdI1dVoJ9xbDWfEOHZvY6mmelu0EgFjvipyg5OwqKnjS
oVfYS1s2i+7PJjW+ADHHwKsOHjmUR2Nu4Dy2jfsLYg3FEDRTM0P6TBV5A44Vak3t
W2x2YC3sYRb1eHarsVQrVctF6x6Kro/2u5odUcTV6MOIhBBSwNVHD+ftuw2HGw8/
/3/F53ixIgI0cXG1EfaH4A9v7nLd3VuNVhSEGK5ih0iQ/FW8wUSoMnFNCVPxdnNb
h2Xzxbl7f1J4seq9ZiqmeRqmqS7JB3DN3aNCWNvEPZ/jyhaS2wEHMxdhlpWWLqP6
3lSfRleNmBcDQlH8D3VfDjTgthIdDYJvrIq6SijT3/werIHPDZ5rjpvqlLM4uBUa
tmYmbHcz0NVVh9tDmiVtRMNKG5M77nnMRmrIAPNCeK5uRoCyyKVWsczKv8v0wmeo
i4PZQ9CyYF6SubVd99t+PuJGAHnstgNL6ZEUB+cTkTVqFFOm0JqKCEE56TGiMJwO
8TOcgpptqe3dY6jXQK1MdqwNHxVd/iRsmCajAoDNztJEGWyER0PkOYORHqMOXg+C
LAogGRGGcl+k5twSl2H5pDJOpAEWWBTn1vGt4ssjaAo+HfJg3QqglQkCYTrwk0Za
llBNtGfrFkDK+OL99OVRXRNknmrpaWZ/jJHt2oGZl4IP9j/vBWecX70LYy1AkYXW
dJdWbNTmGH/DM/QZFpUvq5cZoge0i1RDaoqyb6UuoD7Ekz2/ASXbGhup/p+t7x9Y
5ZkfGRwcsoVQEZWQD+kZcgV8qoc3hYqB4ogxr4IU/lH3NVvLwU3oFHsFc5BqE9CN
hmExNrbydADU61bmQiUzCrOFnMXcILOgXGivAxFUFPkrg0ZBE+hk/KEYBvjifbEZ
HtQpH6DN9ilOMGDugDtv9zqoR/jOIT/c+5yNB6SQ6fGx0O2r29mH0L/RdjoFu7Qo
tLVl+8Y3TxMzEi/a2klwi7e7pTgZ9RhyvfwnAlqgkSMiVq/p3t8ZZulj05YlTh3j
gu5re2Pdx8un3rtYpdcw2rvxf9oaj/CjtXfzTlZK2Etm7U0zJfRnkWEZG4BAG7Jw
JC8gS1Vo8wn8Q1k7/GWvL6hcd6Our5utgpvAKBINc6vnqFGirqBW7/+RRywoovaK
GRe/k7z5lMLf4D5DAD9Xz1SlE22FKbuW9qkZXXf8+RI/ceHqblCYrbIKOU84PTgW
HkapBAu2VQob6C2xOYtnjSKe1eYL/rWk2XYp7SABy/dC3IRH/H83IiYsbCY5FiCr
152xXtQV1m51Gu4W+KW1xwVQ6f11uF+r+N0HhPfkCg7TCzzZ1COu/negVqEsu9F+
i5iUKjZHXUANnZ9jcpwvPB6lksswz8GrXk+yqWrD1AIgJJuXR9hgK+yb7qfX84Hs
WQaWnYJfBebdtkqEQuBoQYMO7DdfgJDgeX7JEqrEzwPB6UujmUhINqgNjPKEo2W1
4lTmXgazkmO21pvCT/MwemvSXBRNNeY55QJbCfzX67XjYdjpYYw5cMIQyBR4T4H1
kkscUEhnWKXG8SxIYGkRKHdgyx0I36wo+wWlNQ1Xv5e5pYuOxY0SoIgz1wvrq1Dj
3CvhoDYn/3ddA/uyxnVMQneuAjgKu0wSeAYQpniJISYRrpGL+OkgA8Y5ZPGTGnSR
2SmGF3LNilCgmFW7jwVZ40OTjWRmTETdJJovMHCu1cTFJZaw6ALXxCz0QpslA4H5
NY+W1HFF4ZyggZ4cUGMYTTrucMTRB1effaaoXQSkIQMm6j6RHyZ6buGrTg3A1l8P
ayluY794hu5KX/n46hHKYGxedHDUw5uMPiIMZaKuE005t4T+NsQofEABd9Ki9B9y
Lj5HQWzTyxwjImFGQzqYpN5tbisZSeflY5nYlyzCxYBFZsSTtOfqr7HCw/UpItMi
nKVyBpz4DwGumJv3Ny9A5BDqapXOISIGTvqk8g/hOFH+1L3W3RLGf4lIiHT8Sfgb
A+Fd74bg2DnhtyjLaimat5V672l7ia8QcMyBJ5iAVqHWu2AFgQBp9rkUA5QzKTkU
nY92NsReck3+GW3/+1rE6wRI22MnbZsPXGCdgNArtlTD185oQu5oWuCpdFt4uybF
LtZnbbKAW4MfeF1r6M9S3gSAHgmTlBgiURKPgqnkCiHaisI071KBJvgHHynEIWak
qNiRUemi0fMXekoPAah1KeEgOqtajhRLDvML2z2sHVouBTC3ku/zw9M2vOPyo/pX
eDJdqKpcZHXVpHHqR6YiHmcYXmbgfMpblqZL63wndBj9GKpjTjj/fs3PppEb98W/
Osw7qgQ4WsZpIe73k4WtyY9TqXsanvI7jsxCk886DTDmmYghd+nB9rPb0BkqrFbE
oGw5MyglID7jOmEGb4MOs/1GrBhB1cXiEchYHkWWeGFrzkgn0eJ4NGSZT47lSVtY
UhrUk503+W3Kk1CusTg3vjseagZa9ItFbYzjthAUxcUooNQ7Z6b8s+601t+7yHIK
yMUdbiPBao2o0K8VfkbgjgPK91+Vwr1J7xyM5Z1qxq94s9Wis8yCeYI5YFw5nDAz
msh4IT6sitcT/gbCR70CVxebmqntuFUGIj96Ux+69UlpYkmzAK2necdpgjW7PQv/
MdLyKJgcvhAbw1F+VKGtQTCzT5puBsXIygcmIFYg+r51BCHvsgKXxwqXQvaKeWtv
9rvw886UDRGipKo+uDo9XRIRVQJqaqYz/mZn+QjU+7wgSIHwKLy8+oUDsiyQAvGU
mjpj7x1tFJz2EeGLPnMeDGiuUCQcax+FUPYxenlsEkvH8KAbRR2YsHkgglB0HFUG
GbBL1JmEKQqPt4S1YlpPXf6jItIeWrUCbNvtPY9AQWcTu7vr6qA95Ytb1LCiZcsP
bpyDgQwLT+UeAqeOYsRifQdHKUEFbDHbKNAdhWTnRok/LFWCrVBVvC9h2/8M9Jt/
pQo8G0GnLoRxuDXi1JDXpuwOl+wXmHk+TegDtKW01K5s4QCb7OuS6q5UoFzlarss
RHhwUoEqETMIEE5iwGZGJVxJ21gtYEZEtVkUgiZEkiYvWTOV2ERA/EAU27KN4qnA
GuwSCARjyqx6anYV8qqPCeQ8lXhAxMhUEhxacQ6bpD135/r4eHOApCRSVMcJMhDH
WkhOYhEPGba3Bt88q7mq4evfPAVtVs7wzJ0iPAG9GAYL8jTGOLBLrp0PD34Ua46h
d2qA2WeRLJPUgUrFivtauUzqsHAWBCgUngk/FrgQFqDgnZpS7fq0frNVwnr5W/LL
6prq1ftL74DxVgIsQmQ8wF44ZaFq2kzo5P0QM9Xwxl0NOsfAOgNRVAE2Q0rXiZO/
XW1Nsza/TxD+m1SfRCNX6so+BrmL8nb5hS2Px7Ua3h2Zb2OhiRd03ivJcO8qneOy
+jRHgNuqr+1J+B8Sl1vi630wGgGxfRMrybay9pP64pBkqYU/3cxHx0QyeqkhShjN
XHAAIL5Fb1/q0q7uFWaNhLqLHdUJeXY5L0AQnclPibyOUIdmIlMqp8divAcOOODn
gglGK5wWFJKcRBszDq23TU19JdIrndDoxXKrLseZVOmHkRCgVzCHdDSEj7UEty71
lUEpit8i5Aw5fC8jA/Dv5nHr/NjJ3JgatyijvpVPfzb65jUE6bN2tvnEKYP/CXuK
jnNF466Kt+wKAYheLANg5KrvD+vb5LGztF4+EBEcUosEQUOHvLSlQ/fZXpJT8wx9
1IjzpC/8DsF2Fri5bPIIfUhqSpU9dt55sgZGmkxrmVZJgK6oi+JbIdzvbqqyuVWx
XcIbyaJ874vCWxN4VPSG8MeFk6pyhibhR+5gEwYqOrWxiZUlOwRV7p0C5C9/NID5
2mH+j+qSEWUdsd9leUbNH3YQXDKZaXdsHhxHsKfcvBX6TAGeeRf6nodfy6oCTA7v
ok53n7X+llQeZiffYsREucpJC7A2gyvuWM/B7b7KhT1KAvUdbf6zP8PCq5939gHf
uhvBnN009gRRUG1Pu7Yq+jgWRnHjLS/spiEZ6SscrIK10dfZ3KIraazeGYFcmANx
5MGATW8NX40RORJm4ZyyifxxztaDNTzTS0zhTkhyRhg9Ryed7OeyptLKchvofPvH
UEGt/seeyhZpBRb1rO1n65yobNLjJxKaZM1KVOQre3sdz5W9V2oO8G8vHQ5KylXe
dmH3FFALzoP3EWse+hBcb2T3YIUXldooDi2KPlynlSghfOm6oUnjDctOUxG07FRx
pvP9COrdRo3GKcwMpojRaz8Tt8e5Nakz9i+manroDJo6mBAXuyaqyUpQt6NE+ZeU
97y3jX5wLt72zMBQ+gzQAnPA4lw9Pcwv0vTEFIu/deojHoPaulcuWu/+QGDwNNn+
imivqDiTK4x22Q+OV+GdCvvF6wdR8pYeotP1TrLIWI9eeljd/wqqHkBVlj7i1bAo
+BZpEC1xcW8qUZgJfBNr0y7y1iDiDczrYkkp3r+YCw6/pDaKJuX1rAy/8gobolmk
ifJC7G1CXZdoKVFvj2y1UMIArk5yjnRbX0Ua1yjtb3ConrbvRj2TApuVA/71qJ3H
dq0R/aL+MppN2ojMNrC8LnOH7LLolyWNNrN54dvfE8SiJb84YeMUof7K2kN1y0nK
g1Qq54Ex6coC++GBJ2ZHeUX6mumo6F7iY3S0u0xcbydc4TEIu41aRqG0cpoRiqYu
5Lp/ffttc8XlgAH8TkOEpbwqKxKQnCBFaV9Rw6RtmAFD87Y3TikvQa9/a8JEixk0
D04M3QerI+xeHxplCpFMudRJ3r9QHhSAiGuhmdf0tyaa32uwYc29qyo6ARpK876l
mswPCoD59rj++caZt2J1UdGF9BlL6PFsH9cYsvnjq1H8gx2378EMyEPpNjwmrNue
C4zYtI9ryPjCaY62w5gPIelQKjwrza1If/W0qOfzk/rqz2bVWPxjzV9NTD8UV56y
2X1R+G9ZAjlK5WItOQj5GBjyQP5+wfFR6bj2FRR65aB89jyDUXbPaViPw8SbnZpJ
QKXz8XyzSRf8Yx4QnRqwBYefFPfBm3KAfDDm+QlZF52gJg6Yr3SyvjvX53nJwzCe
56QnZuOcmtMCwPwyEb56C9e2S5FJO8OdYylbIDZtLIg1YL5UOi/s9UuvUMgK5imA
0qtE0oJT10vWmWm+2tWf4tI7r5wPnN78IUkDPD6639D/dy3wjN4YG2/WQIQDJQX5
isg8Vo7jARQBh2DVi/Apy9tO+3g4/yG/007CoRj4p8vj4erCsnRh6up6nDgCcTEv
OlvJHUQwsUqj8qiIv5vWrdgmTQbuLO4gRSLWJIXLRk3z3rOZCCHwbdzQlJtFKrvI
Tvu4z2xIraUdJGRJhZszgZgDR/6gps30iSWt6TAwSjKauaWfzzH6RcEwxXI4z7J2
wktEXP10DvEqesNCW1oLUcwtw9kfzeDPiucNXpp9HtrdWvbVLqJvDO7EnsF3depQ
Tg5DN9Qdy51q6SoBWTYufM5f+EFsZQhmqBelzp0Zq9gdJFDUrMVEm5hieL7CEAW3
yhxDrJIJoQBs7L67LWcvhLn9OAW3cy6MWtnAwZEBiH/ABB+KpLaz5ILTLd5rCM+h
W1Hjfd9VEQzn7onezNYZALHdkHMSO2vY1ruuN2BaEsDHURblXmYiXY9xFqdC2hSk
DvyVgD4fpLIl5UO0VXTnlBY7OXwPxCovJUtoFA06C1K8O1qxIDATEccr5mxEFnKA
tNNZYhdTYucgkXVRX6XQxgg2OHnGo13QlcG19aUScT3xaEuxUo6J6aln1VFcsCm9
DhqDB+vCZcHSpyExXS17MUHzjcy45/6hbx2k6u2cVkfokjNeDfKA8GPt2Tt10aRe
a7e0xEtIoiP+y8UvWKgu7zGNXS7Bp8Nl1sT3UdjtxgifHD9DY9/zqfgJiK9672dG
PqTapmFbl9ns9X98Y4+ctLYd+dRW2VoH6dbPORbSsxMtC51NzM7WpKtg7EWGR2Pj
ysfoYSJPhw4qVIc9DblNazfArQxodQHiDKqUtQ75QnyoA7hoESFQysmULi2IHjLV
epmvi1IZVoHviJfSfoKOXbHD1QOEIJ9nD3hkLBXt0UigIcgA/r+/evo/KxMHdw90
pJ0EBaVfNLityh1R1kPYm0lTVE1E7d48VMPngRzbBJf6Hpg5tTklzN8oGgCtdj8a
uNJFc6ornZEq/ElrBuX+zKDilyQX5VDV/Kv7NAzqW0YjhwPMUefY9KbpMfL/SiHn
bC1b3BQb6rzn8UQS3jzXhograhhCkordRLgkBPhxrnngpUJheZgKh6I2k3ue+XXX
WxwoSn4NGT+qHMXxcoFaG1QDGNYMsE0ejTS7YInbJTyFKwCXZkAuhLKa6W0saMvW
VLueb+ZN0Stai8N+SPTV3+DtP89oOXA0rBm63SuEgtEuOym4dvh/AQKNihll+w1Y
RkPHwtAJsNV37BPm6fAP+pUYz7Z8ElnZdtxAODJNXS0j7gB00UafM4q221AYnL7s
OmjkeG/hPmHhXiYJ+EbR/lS2YSSakloWKg2nOR9vR3d4cdo3QQ3pVPbp+aO6SCCh
Guoe00ZGVHYpUPDWUng4xEUtZXnr10N24BHPCsp7a5jTGQKxflohml00svuMQHab
o6zdtaiKX8Qh8tqU+c4RmM+V8F7mYm/QbL4buOp9O8Emqk+CTscmLDKSSQC0U9q3
x/37gJ620C+u9NycEKLhh1shI2xsf7I1UFdJkSdPKk2GlyZSc6iLG0ku0E/y9fn0
mZULNeoQNVPbOeDjYFx84cspnNf0dWxP5w9B6r04bnC7O+ja0vj+efWFfO8eSYDS
w0ReN364pbUx+c70QYNmWdBAvrqFnpgjIO5fv34TipBDY6K9Ipuq4hAkT9p6L7SJ
Nh/Hmqmwr7kSA0KRhnjjotvKG4YA/N2hjUzJ7xdx8b9Q7z6X0QmomsxtCO6ErSuc
q+ixTrhijuj3Sld6IxdM0jqWQNDzzGg4SVKPQ5D4c+OAF8y62Bnhk95ksI39cSNp
hzKnkqlCgYbcrL7jI40+QXX77dvoGXWwlqqQEkBVhbzYEqlfp/21gb0trvqiO9vw
vKPfyydxRvbNqzZaa6/Wn5SkL3YbFRUnosLYbjUxoACpnyO9Gz6LbsNJPkAtSG6v
zJ+GANSAYbmKKu28YZWEuLIyJFXYmvD6zpsnor1Xw9f+eEu0BbDAok62AKRK2PG3
ko1QOwo3uIz3FfwY7CNl63KXkaJ21o82t38XBm/pVijiAEyJ7c/mDLuTmmestiPe
/vS+HZGgSruCLaRFKhT75IAPU1SvXkyVz5wkqK+77oruV4J5576AbKYK+R3KUbNk
Aqru4XKOJw71xjVUXhcIrMS1vo6MjLsbnAiNr2BGR4QUypx0UOrEpyoKNWcRUGka
fM+TOUJlGPZo/H9f60zRh89MRgsIpjFW15gK1C0KSzP+uKSDWlNdrZrMXEuUVXW2
5anmRiABWyavHp0ZvfALeV7kfXafpCaR6hW8XTIiUD6sCGateUir3iEEy+QKXBgy
FC8DfooEtYuTPt+ZEn1n/FCXxzg4fVzUm52lekGXkauS7Ftkp9S0y8p26HbtibZ1
p9C/c0STzB3mtfVbEyK1M0fRnPuo9/EkhUF4SWCCnRvkr+QbZYcuxnBUxU5zNkWm
uQKcZ+PVpuw+2m+exMfNof/Ib4Ze0DQGL126xhworw+jjN4XSX2jmeGJVwu6XbGL
E2a4vo9BOOmbvulbW+QbYOCbFKyzRRbLx42D0fGgclKQmA1R3RyAEWIiWwxkcwmY
NHMJEdtnlx4lBQRodZWDQdNIjWQxAzZbbt3YO3BLw7XvoYX8dORrvyY9kRCyfkjq
wNtgP0MYtN8v1LeFPCSHZ9gYaMBfhwtGChosa91BLb890VF/UFnvH95HrGsnc094
dZAU6OuE0AWuC6kqX5nwfSpGyzsYXmASAc3Ex9+eewpeiIWG82jDuVnVl8FBnEL7
FWv7beRuvjt1VA+OJPD1dGa8EJw9Yee6cCJFEUPRMLVmxIvR6UE+TYYTR6BNrBkl
4qMd1Quy2MVRbZtPxQs9bQ9ZokjAwMSAGONMPmj+gz708D5wvzyqiFefm7rFegD1
B1FWoJ1ymWCV4JYuEOy09kb1iiIFFzJ5JK/qzDjQSzGDqpdZ2ZxbWC0loDk2j6/V
AqM5Peuu7I1MXbYk6PyPkl/WoL9nkfcx2txpPApB2sVFA5tWprvl94gPKL1YXL3V
wGnZX0vIHOqaM6t+HvK0pLt7Z4NkKzHaozlMrsGDqhKgq3H0ylTJdTc1tzgoTZbA
Qk7GG060KA3ZqxZqqanVUwJV9BJHqCL37BRCMfZarRs9JIkwbVK2nAMQyYQX5KSV
JpV9OwJukouio03+5xDl+iyBKSRS8RC432LevelnpnVO36XxDm6vkLSFmGZSgjfx
BC0CVkrDQfSL9/XUs1r1DVQEZlEPqHoUUdZc8ylxPiyO1aXf3iC80cKMGxKf2pjY
YmUUy1n5JKijozWl5Tr1+ibOrmJ9cNRtMKUKYiAFfROByRMzesEPzHtYEXX7fWmd
b0YIqadoPM9+wqbXUBCTc2n6l/zgOUBh0XO+ENFFvJe3FP44iWitXEkpsxSnvJ09
kBcI9iAYSRbqD4nf27DOOevTyQ1XRMt20clsktfQL2CgG7z6/1EEBG3RC0MSiNqI
ia70oH6M+3NTmE5aaJgQKQYCJz8ky2Md3Vhx3Qzwz/AZ+HyrLsYqDjSKEW9WVcmt
Yeuw96fZURfo3CO5/NcF0qFCnzamtM3eqT2C4cl4JCa/3C+GHA5nDeo1VyBGoINl
URO+eCcvPe8eg+28qVgQQ8v47Sz1Ng0lPqsbkWe3VoKxOrNAjAU2M8rihoQk/xD3
jM+CmMYf/mCnU+4O2R+q5SHhURnGk/ZLTR2LqZNJ8PHrNkHY0UL3spNL9khSv1oO
7k8hH+4HssJiD4Hs6ePsd9ZluwXJasEaGEK9mLxZ5kmBus6lG7FWKWtI43CxFPQ7
W5ug5iZ9oOJdpHki5939H6Lkh+IDgBMCLzSnSPzivBAeEmZR2we1dFmM4OfK3AFI
4YENc5Ns0pAERywQX1wmgBTJjGraLwMyurQWS1bbqPdJNlNUTOG7b6fzvKkaW/Pf
VXn1ykv3B2bkDkdoOWzbFg6yBmPpeEmGMoO98SPT7TSOwXW6b+mKFH9i/G8RW+xh
rkQ/oO650xucAxFq20SRHT0cH40R4UZsvbdZzjwqwwXosXHkyDs4ZAHvZjwunebk
L6K+n/eCVvikL/GB8NzW8/hnaGoiv1M/hqrFTYRyDe4FoYI9P1sM6ZNYaJAGWO2R
pBumsZFS6Cvg7q95MNsJjyXd20gniXQAl5RB6tPWf0OaN0ckI9bJYy61qS7VJtGr
xyjB+vswCD4Y9Y2degN+fjaT1NGah8Z3HyQ0RgtBPNCiVLoXRlnh4pSendZ0dC5a
ipVeRIvg6usUGZ6SXRN/w0OV9jq8BZAgF18U0vr9SAVbyvFJEfOblM+wtp9852mu
fLu6mnnyfCPm+E0R7F1kgS6K4OFT9tca4aoQNtN6BN8Rv0deTC+Md/gUUdXnTTw2
uEhhpBek0MqhVs4BYSjG8PHWFs/WgbI4WDAIV8P47Akp4aNY23OeWk+jTZP594st
qAOxEEy8VpMAmnBzvD/GqWC6axvIMfbiNkL/ANOre4O5KZD7LRf3p7pp9+X9Vs5l
Eg9VT7TXG3VX1myWTwfCUyXoefUoHbyRReo1PAfWS/jI4zkCXXDfKFyq9k1iHUB0
br01Os+AoTNNWYTh4oQhxhZWxDw1TVUhyHzsjk/zVQeI4eCaVAH0Y2x0p45RFYFw
ZuQ5qclx2iePNzDsHWO/KeUJV9f0hE3jaJIhmFIRdO4cZDhqpdvTuKkzgI0AfLQz
K3Lhu4A+6nCGtBCsZkTBJcp4mvzg/KMqH0/OhG0GluYMaZRcKp4IlTrZYUg5MOzl
ImJPIEBBbN8lmPdGl5kkAhO3MZY7N1lI7jzmKzYEu40huAn0QT1ojm+0Z5A7xfEP
Q4umy5hHaqrUk1KJwgCkUDTR1zkNtCRDOyQK2Hw7lfWQq7F4TYZrwFh7CfTeh++4
q8EGuG4qGP2eSa/GLWL4okrAD365lU74J9I3FA64FHD4ZZ1qJoP7WJpR8YGN6rW5
oPiytm+/pLCxz0UiOc0juLeTrStw8LsAw4UgI2q7PcujEIv81XCGYgMJNt3AQFxA
itnjt2OfMeXNj+Lux4Lwwb3rMfC/+XkDLw3Xg9N9kNJ1nqI9VK7ZOcnyRrDeri0Y
j52XIEr6IiATbYr37zJMkUhxtT6EcneS2rEPhcbwP7+NvTW7qFqf7W9xNznc6l/o
R1s8uQHqclpi1RPQaq2du4ju/WKtv0YIfZ6xGMY/d2Uuo00c0ltMAxtRHw5FWIg6
n71cvdfQ+UpF3a54PMoxwiPbkXL9mYiyFVyJVa/fsXPOuITkeAo1e4B6VO2BU8Uc
xzN+eZVTrbxzN/2/5ZoPTdjIuvRWSFTp/2YOaVWBrAEI2zt4bkBUP2YKfB0QTMB9
N0Py5B7AwjLiTnjGeuMdN4BXE3wQMImTdgCauujMUV73um6G8xn6twmfxsWTiyzM
oGPYiooao4hC4eRsd+rCPf35H0s0RCl10uw3NeAMoowql3gVNtQXgRwnTKWcuzIF
xhcRPenUMz+cawgveHtQFxQcOiNpUwINI9+PK6dofNsBjaLVtQdj3qFH0Fvim361
Y1l14JqvMwbrACxHoioTftsTVIHYBVqjkI3czbTWfVOQYHJmBv1YuztEcSx+6JOB
kimyGUdXS5jbyHGeVENzIh8YRaW21DFuuC+oXO7Pmip0qj9AE0epsYOuCNnX+Bxt
lAZw6DyZpT8puVAY4L5gmNQ84U11JpEq//mlk+NXAYYXQp87If/qeLHvY7CiyWOY
BbyLRIOi8yAMDp4HlznXruE1EyyFhI0TmZi74CQqK9y/UNUnuWdOGaS9UFNKwclE
coeLIwxPlTmQdnLTIH4zCgZODUedtbi7dIj2D9k8D8LIt2Azh/X4WXt8twAf4NyK
Ls2itcKaqn+l5mJ8RsCjlUvWh14zgwRFXs2I8wyKsDnefrEkGHamIfqHbSnmf7ra
kXUYXSOmIBHGIIp3jSP2PjOQbCC3/irDdF0QjAzkXdiTJ56KKjGQmEx816DC5S7U
BXGFluAT6pm85Zb0zk4VtYMi/4FqUsOhHG6SWh1qYF/0z5fGVz6oOMTB2Plpvgl8
I4FjIcRuN7MAJ3v8ZVH75B5P7VaLIqfVTXIy5yXpf+4szY6KQd6UPlY8O3sYhCEY
799w3ozIY+6/4B6s3wGvmVy8rfyQVjdZfKFpYU6Wb2kQ/ejWew71zBy/VRufxSu1
99UvvAU3cb1LY/O3axzaqWbBZe+HKWlVqymbACZ4heIv5+1FM58D5uyFPqIthDUY
QprVuLNIJYKZ6+wgm9JvarHcF5w00j9anHtZ1sPkDQAlQouNIfoLvTcyu3lWMWUi
HEKCbLd2bMyGC3YtkOOUVb0ZiKjT19WmlDXi6DHwX52VfdluG89PaWUR/+h1H2EV
JEkKHcAywhCN5mu55DAJ/s03LoCz+uUg4/AHs0AR8vD+bqkNVn4JIDeZtgLO7R4L
215piJdLkj+WggXQkMDOnWccUJwfjhMmKeWUBjSQeFuPoQoHrwrck5K8+t9XPQjS
vNieQ4fJQ7/UXlgyRFHzKGbXVpquGzAvMiBVqKAzYX8GlN+0L8WU/lPOo/VAjhQ8
QEWfZTEvXrDdxVboyc8dWGIgAuDvUL2YMJqta8ci8nvmpwvLsF01uVqZ3cStnsaX
OxJ5EbJN2FbWTJjW2z/S0WDLOzAV1YI+rxqrYlAAowEgc6ahW/zgDkdF/WMT55qA
+dJh9WPxfurtu1+600rYw2EFlid1Ky+2TWkBBktDUFpSTZ9pTm+MUd9E6AL6IIHh
FBh4mYq6iIdIS8u6yN1VF1kFHqN8neFHwSzbQb9wn2pJVQwr5DVLzLUDEb7egA5H
guzuIbO/uQCYn+zwPhEytrxSLPRIjsH8nbQuIb240rlmohujXUDq+BafChJBNuuB
H63lP5d2JkQg0Q7W8MvNMsDhpZixcBw+cf1F5Qf4UZKtJp4dcCHuty2jifpWqeET
FQfiaYqSgL2lyFaOqmaQKW4XMMxJbPInVUyMyGY9xf/glMKN7U0Pt7pSLKCkrq0Z
zN+7f3Tq0gTGJOb5G2hDcPvmGivQl2OK4ZI6CTToyuYHNu6mSQtWJBiXXujFOeVG
JgmdGNT12PukLdugGIfHZts+s966mApgWtjJ9UJ4cgySyNkeiMVUP2SD4ZqBy6xJ
y0mcZyqMV0AxIvyYBPjkVZCwTrWRvtoZgkHXQ/2stkhWGwQ6/mx0LOPvQ0Wb3rCw
g8V1/H938pYXkxPjZ2uBX2aiQgJbULDRkwUNZ/NFPQeuzvzNzxis5sUOxE9dbPEd
gp5cGqhiwE27iLI+o0bVMcrwR/KRBcEJASA36cIbH0mOAn3e4z3Z274wTDlJV+S7
Co1q9thLG7KTeQInYAByJ/1lZisAMIVgWMFcLfb/DYvvRbbrokVvXzdAAh8f0UqD
jm72vJYhoPAN3+k/qXySFHkM/KBSON2bhupVKTwCjbaOvCEnJyTQXXhj8kSRqNoh
lGqroD9Mviaii12hHbY0lvyEDtYT9I7Tw/AQOsdSW2IGwf0cSxAroU3Xwvwp2mgk
aS+sHNM/dqX4SujRYr3yXldm/Bmhv18pXSD14BRrwNzSAgIKtntLMnqcGZy+xB/D
OiyzWKdqjnT3vRvaZGzYHmAzd/lDb0lJzLcqt/7WUfDdFXakf+OkIjMZpV9JhJN7
uoG+BJBxp8ezBIu+kUqlRSqK4fUXfAZnAw1VH9Fp8KByBzxKG2uM9NUaTnmKAkOd
mtVCfPGXsB5yG7mG09NsxiakJah5KA+0r7jtWsH62KtcZDHmaTqw/cDLT+/E2+Nk
WXvtFy3u17x6/061iAyCx0RNRulfsrwx5lpj/6jCNNs9KsqwY2wTZP7H6mi0VvsJ
qP6IUSTf1jEDH2JDldbjVeyCx2s1Hj1SKQRsiWx1VWQix+lAvzR3bEZ7h3V9vvQo
O1QJ8i91gZ9Kf0Ec2bg5pHuZ9c6FtboaBZ9pZuW0Zz/CraxS8R0VtxBUGsNrLHAk
OuYOFVKfQIY45fpAcWyjU7Ug/rrxfmAIqgszCSyL6AsNgLnBT4FokFWpfOghWkp8
Imz92sdEi9F2Sf3FCAxzucPgFyT5lXrNp/JlvWA2D21DyOgxh9FjJKDDpaXbgbAB
W7UhjwQVpikjp304jacB3mXk8NotXm6D2gghbf3Do3FoDX7CiytysDE7Ph0Unlfy
ElQMw+0/+M0rg+CY41Av6OOJgeJFGlW9jBZWS7D62fZgfBvCMnEc7K3RHOkUrhvF
HVstDKWCIqBWNEx77n8NeA+DWpm1khyGmo4LdfNW61uZ/9tDdlvh9ZG7tF+hkS7N
Y6am2ddIL/J0EZBGUrGFAWJov5PAL5l2DQ4V5tSR5aRoiqq3rA1PgYNEgyQuXZkK
4fJl6jKCX8gDSmu41IBF1kkFPCsYD46Fry7WCZ7Z9gWeudRqjBAnliZzsDFUyeSP
knUCBDaUIz29wtjVPmtARF+EvgdH8TsgqSS54GC2IwuHO5/7DtJdqnCI8NgnVRSW
4d94qqhILKeoL/F8O8RZOk+h7VYt/GkHTBu5d8zdAViRRbXmoNgHnguz/elbJjWD
dLCbRKSmPE3w4KO0gUz8GhA5Rtogu/n5vsjLzvKuoJ5lci8cm7cNtkR6EXURWA7j
MM8hgoccq0nSLbLqZIPeCVzQdkWB9UYuRVOpqrUGJ5Y7VyGTkHDCogqt/btWbcVX
VeW6degT9rSxYWCoIoHTkjz6XcTGfRushlWcgA4eUIfV1oiD7F5uKvPpQD600Igs
CywarIXlDkoAqIJXy+R5dwY2hrBnSg+hlUAzyv02++fyf+Ootg+Ozv7hJ7Wb6k7l
u4X+IR+JjhMXZXi5Yw2tb8WryVS8NAzwNv+fvlHqm+mO2tSH+i+GPirbCBCNF2Wx
PqMVdvbVuYEBDuwQ2q57qMy39vHExYdkgPG4cwCmmrqWl+kJ+hHMC35OB1hKsLm2
rOq9nOkoOdPIOa9sHwvnU4HbrM20mwF0nEz06ppb20GfcJNK1OoXM/0Ckfwj5oLp
seAJnQe2zADLJRQZs4XE33xhGu7NqFhO42v43iriMExvoQNq1SLwRv5U/80zs4TF
dMfcfQlZqzH3Sw8G5zGS0d0PgsB597AmYaEt66vKVk9TXSidOLGF2u4pGHszbka+
VnebSwWxdk6w7IB3uAk1QzGMhdWagtP5zB+Vd3LmFsbIzvJ2i5Yuw7oGP/3UMXeK
WmORXYc6q3selkW3Ctabw5/3IuhNCSBl4HhIlNZoiu39mgGYD8dsEbh1STEDaspN
NUFO6sAKkryQvPZnAMjpZ2gM2Vd9k+EbJ7vitDVkOowoJ1NOIo7yTEsVQRvgBRCU
nxJRXVMJDrV238XMGjCPSjv/KRkwKoAWVO6Q2CcAlzre1TS9hlDPwPPeNXwKxF9K
y92BpvuzRKIFByBK9XkEb7kISCwBStQBhmU9rsdzlLjSYoU5dlqVk35xnUJtuV3f
mVDw6oIJ4C8gMeUbIZzIvm1YYDoLO5hqNlTI57bmXURg6QFoeLAXTIij+a6JoP3n
lTmku+Nyiv+mVkUmqMHtSXzAlJXj7hNx89RhFHTa4ZFJ2g7GRD2TRGlMu3gvoH+0
a5bc1mYfsNLL39Hg3oNYd4NL98bNMAmmGkcPX0JgUSFHLE4wVeOrb3G6gRV96jRM
2flfJoC0Ao9PzQ9NfX2Ia0Z5ctIDon1DweBdvLTtO2+29yFDqFuNfxtKfg7ANWJ6
plGePAqhBYMDhIbpjlFOJ2m33NrY58LDw77idnjPryTvAG+QT1w/exfDm7mzLrae
0nyA2BuPUDxew3xLmz8DGqva+a8f2cGzZZKQ3WdwJO2qU4HZ/paFM7LmB1IpKk/w
C/jyG1rPZ4PLAl5hLHxtkj68L0r3eW2/gGsKm9CR1Ai763P4CD1BZd4X+dUst0Hk
tHHiN4ugcUio/PcsCT1KUy2178gz6rYKqI2iH4CKt2C/dlrO6qXM70sRdsaxk/KR
ESe5/5FeV3P7a9/F28uBKo9EVGpGkNkeq/MZChmN/W3KnooVhCYUKdHASKlXBteG
ufrnNv8oMtNNBqFqye2O/DfdAvwJIrNcke3uq3nTrBHhLnXBkrmUXiu8pxmodoOz
o6awr5A68+vqssA7iIFeyC9sAkkO8xNkfpgyb/iqGD9XJPvSXLzsmHn45+ZKyH7q
cttTbarFC7/b6HX2lm2FNP1sIKLaUI+rrgzzMPYNWcdFUfNN1Dqhw5qiW1Q9pu+v
T607BAhxaYSTRzfcMoFv9p6Y9apRCofuxV51+UpOC9XtlJyg4CsdlIwgjV6SPtEs
zNNBbqTA/Y69rgdsQC6ZmZmfuYiua8uxfeM86wibHG1sP0Z6skL+46exFKgLNT1R
rQluxsJXzrEYdyqXVplWwu08VejP727OlTkPpA238hjFl1JlvEoAjmFkPrKXmO6u
UTB8bIky6nMqBMStoEq+8l6hb/SGXF2YZ/meFikEspfVPfj+4ldCaCCTqtQgbdr2
3FVIIq4KYUxGgRINNjbpIVfWWHHdnSsg32J75mLpIpLJ4Rcvi+0nQtJ6TSf+R+gM
mhzYPU9HFDqKGBE+ObuawlHLPzNQCMsdHFDRRvMP9UCJFCepdIwWONZ0BhPHbsB3
ZumL7U6L7vKb1umctCSyz48FWtBZgcKwONPJnbpA/f3WtIVQLAc7ViWfevAKbWQC
AX6csUCSggfwPSZlbRdZPK0X+cqQfI7iWaMEAkeNwWorkIv8j+uqGCsodkuCVRjp
ua02tpwbG9vIWDAM7v2DdqEv8Y8RMtbL16xHyiEPp+EhxvJkZXjDp5WN6QMWecTH
tODQrAiuESA0KT1tvJCq84o0vjXyh/zjxWslS8CCHAkzJeSg8RDuVufHyKwjtH5t
HTL5l5z+s9th7LISfP2kVvzWoxyrJJ+ux6Kwu88gq9zqLrnAQE8apWbl3Bf95ayr
3bmM5okXk7xRU7NHiXDTzqRiSfqal8zP0hcIgNeY+7acWuEG8J8muDe20a1lCf9o
SB3BLUQhwNN0PwIdoA5tkGOfTGaJCidDotOXXDWUa219+jGJTDXtFFUiwCD1TDKc
pWLbikyIgTQxRsu2vrMef/f7puIRWq4z5XOYJUDq9gw4C86lnp0o8QEuFYq8w5Sb
Opi8a9CqZHIqlj6jhGOkH3E0FYLHKhOlKnKXVjNB04z3uLnsR4+ZiM3RWsYbw2cn
HeTU51DFKi0xc4Pag+rQJtkuzgHNVCmfPEw3L2Hfq39y0Qhyr/tsRpKG22hUR/V8
7B3XpZm+NaCipx7as7MQCVStWgWK+jRFS9O+mFHMyRkCKFrgAKN0dBfwn5L24TRw
VAEgDwl4DHz/c/1gFEHmHadgyFkFk5xYKRuXEeNx8USOOCeUTD1yEgZkSO6G6ftl
C+qVR2HfArzyYtna5341EZPnkaN/DSq8bKRFdnEFGXgrdmSrdZ46Hg7LuNW9aKiI
AEbe6i23oIkGSfCY1kmAFOWcxvLN3ltYJIti5YbI8skpq8JYgAVF5VVLEnErPTen
LfiNd9P96h2ZAniPaNnP8NOk2LZocoSGQ7giPiwvWI1sy/5LlF/iFotfGWTqDNmj
quBenCox43A1IJOTqjdHhe3gzNaoXByrELauK2gSszIO+1zhX1mkzy3q5an0Bv3v
7H3EHW3vQ07ySJjPV3yleRWMFs5XpBOGgQjLZ2BRXjOL3FaQgpIUgwwZoosBKY0E
Lo6VoRbsQVQkH0PRLCKfbu2QKl3T/G9mnM1qQthO+XwTdHpVTccmFy3oSqqbGdNp
4xrwhTIXMck3RN4FHzgbjwADTFkgsLPrRYpVr0YIl/5ialo4ckMwTFK/MZ4BevTw
u9f4NZPJjOXD9RI/1rRgDou83QgDyaEWUqatzcLwZTKm2rAO980BS9WSUqLrFYeU
HYWKCXrE6juIgL9fKNYIktMuwKLZCJSo9lDMxmyE58godwxaAOXIgv+y0SkIJAhQ
4h1JG6umPvN9C0kZS4eSb2kuU04L22llLGi0KSeaTv9rNW1MmCnRAVtxasRQoYP0
rmElfTkg9lPYt9r+BLCNJiJwf4DmX7shtm1uEiNnJqqx/U4bZ8GplQsts0PTB/K9
uzamvIvI/7j7EzlPyWzBubpr5K4Bcs+fefZLU3txpteN4eEeFCTSGGeeWFseVZEJ
qH4EuVlwz/U/fLL5z0ddxsEC7z9z9yZ3AmnDTWhh80YGnUBGHxuTRnxmt0/QnCnV
zvLb3UPidxBcyBTXRdf66TgmL62K85hI4/bSsJ3uw/D6TCBUOl62jYhIvK1diWzC
o71NwLLdMLFM/UWC/fZ+TZtXaWz29UNkM5Kx7IzqGBf8pGvV+WVKvqhAcd+HqTIt
DiboHrqgRf6ARHeH5EeDEmil/payw7VNZNAxezgmfDJZMCaub7ILtOOTpbFoF8xT
m8gkt63obRE6dru/qpY5KpEG/En78o6zV7vtBSQSfRv6aJwhHlyJn9UjCJrviZFj
EPAH0G2SA4N0+wG8+bpLP1Xotlm8aofmacFOiP3MOsKpchfmw43pvZFSPgP3qxd9
vQThKTEAe5P77ZLFUmUlZkaw4OyVZCCNmgmm7V2yca/ANSvF8KXClGafKDB2r4JD
NlbAlSev9GIawIykF/HQQBNSb8SQ0JmItSewWiT7qvdsXLOL/xR/EEYpBx+mPcIy
dQB2wzupXczVtgl2YSKzPhklqF7+Bhv31cgPwPXG8qpwnLtTBmG8EsipBihU0EXw
cb+91B56CJTgUTzfYm7nezY7X/mbuNQRtlZUveAaYr/13S8jvp29aAmi2logByTJ
iRXisONULlnJouxUSWBlBGINuekgxRhzRJB2AhLAwV3BawozSWpbMSXIPNnsB+PZ
a2dzvvfAFG6SuEe8p1Zwku7Xd7IfTozhWCceHkhBxvx/6tCdk1IZxHj1S+V5/yzK
WzZuLdV3BNGFTkLRQZUNBdVlbLg1ytksImEWh+D05ZCKTlWOHVhphdyZ1u2xscmN
2Hw6/fPPWNorwXGIfMSvPTgpdIaQdj41PkbodVYPjZvcn+9gKUZp6YXb/2/h9Xpu
zyrryxi8b0fh9XXxRaFY/NBJ2FWvRxQY/Xs8XjuQnGjUxeRd57gdIEDKB1s5B6QH
geEsn3LZj9uyoJG5Ps54NvQqU/8avsnXFx0PJioEgWVY0gXwyotIn5f4sbcVnvtX
o77Dj/OzKq50WNUIIkw8kR1EAvpqzQt0t9G7a5kfSA97sZUkvn0X7X5XcyTOxRKB
Pbglm8r5oORojPZMMSBLY4wuymbVbqS1HvM5TleP93UZiTzElVxPfUOKrUoxWC2S
JRjuBiQpxpU6TooJlkoWU8u+iLE4OJ6Hvfzm0T+UmdR3hJSLEhxAKnqWiA5yDbxD
AbA4wz6zZWk+TJRAt0Ca84bQ8nrtBbISIFALDaUmASEO5CHX3149T3YgNRiD5p2t
A74OuiK+szEHxvBtr5PQpgYxOxUTiFceT3MuRWnR0VC8hk423q5msUd8k8DwM4Q2
DyY6IjYBczkFaDFMhWsUB2oWU7UJlx2rbs5hFORTX+8wYRBG26j/BOgXe1evYDyJ
CfoaOxawSctCALRn3qvq98wCcH9lfgs+kmPmxOTiikHpN2ulJwpyl6KIjcDhPUhW
qnozvHUKqhcDY4z1STjtRbddwabQ3d0c8JaOKcjiXLUGZFmmwVdqQQW7k5SuMv2k
SrIoZ76EtYM2Y4f8IOHtTZcWNMaK5ZQ59dKIzOrppmF+GbBbr5psyi7eJZL2sWoA
8G3lEuaQ+I2/02nmfZ8ffs+5isFeZBV0ADoyIGJACtBVztiJ0ghmV7ErwHooIr2M
eVtRrmaSUd7hRg9Tn5x48p9Cc4tvoXZKrVAaNZqq5+/FdQAusNqmalMIKNPx3ctO
CLdG24nLy4QA/CGBj8OvZ0N02XcvbNzpuuTSYAAff8X5OrZpV+UL0w4E2HkWIptn
MUoaFt6a1HTiQDF5NAfYkRuoqjH8ua5GBsARh7Bmw9mWkUYfc0GSa2lg9boXr99j
vsP06FBtWIkGCsW08DWVWZcufkaRUi8CMgRwd8yspAotL0MCWK+kYUaL/ASwDTtC
xXp2MPZwRdB3F/Vi+aeZYaqyxHSHSny01AIXuq3yTW2U5ax9ab12bNb6cv2Hqa0a
ccerHJOvQha/OWDhY0jtj6PukrdQ6Sv4oxdnlMmr6tsZLZapBJc4m499dlrok/Pd
/ynBpywz+vwFV4Q2aSz95+2ZZPP4qR1KpM1Ad5ltIKBlNSWgDuMDTCLOxf4/3bpi
pzpWChceSBnfAfCjornkH10NDYLq6t2gXoazO8nU8VtB248lI9U9nRXS25gi/g6B
mKOXtFfC/ogght5rhJuIcOBr36zliiP658YQQWhEJCPjWmTj2bkHUG6m6/TTPf97
h6LevvLLYk8oO04kO5NubV2q0nn119xeUQhP4gXSTeZj6sL+a2oBm7iBEJBM9J1d
7YJaX5mP1al3aJxmqt7pjb5pOR9AeiJea9tGWxmy8MkvvUajparAIeFDhVychnEY
50T2N2wUX26gEnT8ygKxVuJ8vuxIv+jqYyODVhi+ezf5BqeRK+vk67yipBEyVfMO
andQOknC0hTnUvcXwr7ZqcLRiv8oLLolB8//KsgdeHcdId3PkLkOqKOn/bdy3ZwK
Ga2yDuagVH0aOIe0+R/ZYzknt9Uf9AziJY9G01qZg1MZmOlP7arrOrglYC0vYJLC
cL7dUHwxBaQyQt4w/9/c6tIZCja5R15JE9oa8fmXZVWENmty54kI05CephSzf3wC
KgcvAo9OHEVGPXIQbsP4/KsGu+/alpsY2yMum+kJTxZs5LTN4AdzRFOX2Utkbi8F
MZoKPjmmyb1Ie5UUzxp7UoSxIRX5ddS3vYU50Yb1EclsZnWWDy9LwsQ8lQyv9Nxg
ZgsEPVRuJqC1rPATRFr4BiaUwGh5FW+YT4qo9oJ5p+PU5KF34mVDYKHhPfGrAIJQ
4WJpsOwRnhX6NT9kWlzWRmKs5Cm0U7jAcbPqrT9uRX9ALpYnefjApwG9aJjLZU0K
KkmPtZjpoHyvuJzay6p5jTBJq/tL4CrGtfYtrlWi+2FG24c3OEkoqnbK7l9WfsS7
9EJ4Lka5IF6xT2MXBpSwGbsAfm8TcdyRXcqU1Gedhwj67r/uZVvpM0pC/hvGnFml
xpi2XXZ/QPqrr5ItRNDIsxxw3iyTxbn6Ku0QyjtaisSV7xK0VmWNnD+OSpiTADJW
+o1Tm8EJ7iNKrjBwOvlkjPXKtMeZ0yFfQVPirspU5ncnhsEegblXLQurt05tjn1A
D9b9l/beWY31UgnrJ+hQBhec0nSBk107eiN4PVlQ/4EAGy5I/HQT+ncywfuVyhpx
4zKTIqoyG68OM5CpVetdJAO+7f+9QjPXKrFMmslUZRFyQk/UVjZAOMcyQy+/CF6P
vI1lAqv+uF81RHIySEZ+rU0PLwX75EsJMwRa1djM9B0KTpA6HrffLOhpzabDvQED
pHNYIRAdmw/foY3NuJ7AA3Hrd9oCH5Hhd1uxqsaC8sgNhGLnt1P/rA01PvWoAbTa
7+QscG35UADHDeUc+cmwoKEfIkMZMNNsicX8/MllLuEw/NscQHFpqaQ1hWJpDpT4
El/V5X5zJoroS5OW9LK4/qQzzsX1YzYHSVYxkylitCshY1ReWmmvxhO/HQRYkSo2
M5R64HG54zSjEg5EFWoN5DJY2vv7u3GzkuKr0T0xBOoCaG3WhOJQJfdNY7ZNFTff
/C87GRJKMfHNAwbi/f8e32QqV6FgG9zBGsukPX4/LRQG75zF8W6hv9LWvT5oyCuT
FjjTO3/3u8e6ilOVAjj/OjCi05D6vGB3yZGcEY33XNINrVrDk9mC5h7wUgCuEefG
cUro8z+btKS9sba5YKGC9Z1qThzsZqn+y8+6cKQknUiA+JSctovScuj/CDRtoY9g
RTrni76Hm4A6RjC0GmS9HkjA3S/kWjI57+tFFFRv6oDyoXrE0DWJWRLj39uxe6g+
2bsPlUXTuWNUc4MQMISQyE1XUGSLKMTdgD2pYWUMg9fRBtu3fNNyuCHBbap8AJut
kZQL0QDMx/D6CTqq4LZBARnzizeCcOAqfMHu1oN9WRRdupj2kxH/rsk4D+z6Z67/
OXF2iWK8YcOBOA3DdGBzDNwUDVx2BZRd7V8V4WwXnLURzDrX10nqIPvIDLl4zeGv
4aGflbdaeJcnu1iSbLXIaY1RjAplqZy282/ICds0TxfxySl7dOg2zz8BLP/g2od5
ii35BNJweYr17R0GZAQplbmL4HIsU440HgyiYwfRuoeODJX8a5e7s8hodW8R1fUZ
AOofnglANmlGThStX7Cic9/73N++x+zho/BCA3y9WZhEJZER6Plm8+/LUnFurL0j
XLG7Y2EqjNO4RO6QBjOLqU6QASRGMey7pEDJt+pLSO7Xw/xMQDIe5+0ZKkNsD3g/
2JsqAyZeH3QXCLRROFGnlS3jBcbNr0F7BuozP36fUrgYU3y93Bns7BSd7OseEPKA
tih2IJk6gUvqniegQkr9FCOsJb1skjZwo0MTw6Yyda6YG0a4QWD0L9KHIG3yAg1z
+5DUX0NPPnondB3XcAVqms7mp/mCOrLrih/joOwQNpgYpfsKYBYQQZZ1i2VuNZ5R
XVRNGU+ennj9IQTtV8rBWSBjHInasWv8f2M/6b1+iIEqL0Fr6SMJzg9DmViVg51x
E8zegs62ezPgOPut5dTBeVDYvh9QBPzaml2nZF4/q81uiEakIz+eiwc4HQs/1H1C
pVL8DgbEn0+vMypfOXogSVpdDuQWASQFF0rZNznyRm6xsHeAlefpLaZf25Q06A8L
qn+teI6klk3RIdM0ITOqrgvAps+XcTpeCCi7i9EcT/Q7hOTb1MJDfnWK8HAGTjyn
uZvc/QRyBDzgjqNl4DFltQzz3enR8JFa6PheEjA95rO3Cti7OQr3oSG1ur4THKi9
StMe7ige7zhA8IPFg3g/FdFqXVCqRENHW3l34hZeW8CvTVFX16NhUcyHypC4wNd0
vGGtqZr49Xts0aqQNrfEWW3v1Qd28Dad/oRrMbSBoMR4vti8DvAIe3vQjSsnxpGk
YWUyfsd3eSMlifUty++7A9Agxt72DaZNqITUZ7/80Xod7Gft0GiaUaNbSSuY7jUv
4tUlcDCyQBzVaOGZxxEkUhR6DGKz287YvGbrkgeMUscYViVmm130Wu34bHaclSEa
SbzprRzbcG0mmSzcc946Ci2m3AQqICBojexJ38dB2ebpG6yLCnhDQz1at7rNJQ6y
g2L2jSbHhqJUCmvGv09HvBvTbjVMJ7TZ+3chfs3Ms4rORK7wsy8+8ePkTjKszsnG
mRP9u0EuJhPNxc/TCTNKWPlYfhfQiPUhGBy4714WtzYleio1576m2Ndh/trRMFFk
d19PWrn4xkown75xkamYeTCmD4DNkKkkST3zdwrhX1DYkD+r/EmH5Fxpbr3g3glD
RUIpbbHpXvAYw+8Vg/OZXvKyKDp69ysdJ+Mb/vDi76ROA5VEBECTB42DmyO+Emfu
zQURs/i5y1Q3o4GYcIcDEluy4lZkXevTSIliO0haWCxpa8kkvP7sZuOmBOi4sbWf
uruT9d+0HuRVZTfWOMcx4UUS9SbQTmxeTGuKSuhwDrw5WM24vQcZ1TeVVazw8eNu
uTM1pPMez4lWqVbzqWDqo5512t4CSekBpguA5v65fWNYoI5L8Drwv746DY6uyunz
hMRMGNOFGPMr53Cn+ficRP++G/flifh5FMWNcLMkl80aUJ5fFSjmL37ch2PackTG
F0XphYRF9FYfITV1v9kKVsoYy4XsUmb1f4PDvoQH8EYsJ84Mo8WxvREHr+CYd6PO
M2qNftzcrwTpGV4N9pqLOJVGsFSwQs/hwf9TUxz5pjqKlMtX+NO5LrFLE7jLVBwm
NaSYCzM2qtkl6//1xXy84Z8sIYaP9yPRFQPrK1u8bgt2q30lwP49R0v0psVuQpBE
6C8hK9QaqugMTL1+IJ/kuXL2LWXoNzeIzTEdZYordx7R1TdX3LvdHhvEyYta3HP/
l85ACpeWCKTZXJk8ax8T1WjIIBKClaznV8JVJfjeI4o/1oRykKezbN62rkX6fWIX
9NhlwpGKdzsh1MR4+DcglR+HtF+aVv1n58kPSZkV8jv7mGWr7+KA4pPKbknN8rDN
5oVAxukhJVTtJSr8fqPbBS5fgarBO+vtMTL6s1eTH4vmXRYJQT+zEfbHj/rLWS4E
Eqr3uWH78oCgwzOqEu5tPBMuxb1y1WeCKn2h9WH8PExHt0EBOvwmnBW8IH/yVXR/
h8Bl7V6qxEKIMwZLlYur/KBJsvzdZevOYKeY/A33JXcU8n4uey1Lf/wcxVLDrqD3
NYSWZOA8FmPrx2SkBrrmZtWqwP+TPxpYU6ZamZPloh+oN2EokTG5jSr0Ys6TZueR
NfX2cLB5FcxrJmbeCSpWRpzAvQHVkZu3LhZ7Zo49uYb/xvFgDLGdhx2xOfTkPQXi
9hh7wyxg4Qt2LCJN7qsSMwFQwiyBGdTPLfCL/H37tOSXHEC1Y+dT4+3/v51xS0W3
oDRk9ZwpBmAs2IAJDWMAnC6QPAmL+JPLVjO5bJr3ZSROcJVAdDXahTuprEDWjaHu
ajMjPZXUS+R+6UqAs4R8YZt1JYgCOCrE7ewX0xeHUbkhxSNEht7TocgvrUC0QYRh
txcAZFDE1EyS04iwlF2kyMvN7GRYoJIlATCMKFy9dJMQJI0KixIfDqiTW524HWdv
iq+i9W6faxKHsQwmovtgdxDBX0mOneCFqaEdkU/0Vo/ThYa2EW69bSG6m5Cqfg1p
pebM3pXXTKVG+7alsHSUBbAv2sD8CFw7YImbVA0NCqvBl+Re5wtqhR0wVZXZ7wpp
UYsYhpOb5AMYO0hLOQRtyJ9KPKU57YcahCO35jWbH+/uRPcA7iCnZwFxv0o4WW/D
xx64wnN9LbpiZkWfuo+C+sBZgOzjUUZzNWrIqj5VGVXjf8f74a6SskKOXg7s0yUC
d+f2vlakrdt/2AAy+vZ7rJr5qMZ18hzHkXf3DHGX577qLdu9pBIycq8pJ3HIHMap
c4//ml7NaLJp1LmOB/2TiJ/2A9Ghqy/FTGZttWomNgtPGeEHjr3QfqTC9Sb4YKNi
c5GeqpHLB8TJPM5pCRtBoGobK/NVsORqgsjN7exWXTqDNugZCuJSPo4orE/yZtfK
cUVjD0GP3cDI/XtQ3IzXOhgyvczQFo2iHf/aKaZboklXNYz/6HKI69mUnrwEZE/U
gwtdipPfG0SSNX50haod0Ob+9a/X0TdZVtiRCrDqFuc+2laoVSiYrrUKxAzAJ7SE
5oFGroyCgtjGzERfULbNF5+QeIqrkAn4og4stzf5sPZVVAAiZ6opsyow0Ybf4aCc
yI5ysjCw91ROJsagkDBdVdhzIS8QlaKWywq4W81jXvB088y15M3A3GsuzMuGq3jd
4jvusrHfRAG+pvH1supNimSUOJnBjU8tIDsxXxZou2G09sU+MdkEXgquJJflEAVY
IaaIGCcuQwO4bzs5y+dHMwDGV4dqN75THGKSIoHJoD0pIPZRzaWD+oPeSIWHoOHc
tGT6CPYynhFZbhTbgl1ZohVokz3r2kSRo5KTXBpUOiypmqdnJhX1KnIbFRYUdT3B
neJjy/ZFLHRlxbJZNxvBzLAIaYRXYXvHI0R5C0Fc52wvXbXyihkOTbYK2AJXtZvT
ziyaK8wRHCNfWhbYedwMYjXaXBEh1gT1Odk7IYx4QhrcePys+i6d37IT0D8tMTAp
crGqiWOLWR8gMyKbuF5+12xNLDqMGIvO8zbdjZyynA5PQGI3O6altwsLxaf+3mET
J0aZ44TxmkumUxkhI+U5pZfPHF4sT4dAVM1EkHYV9T2OfiEpJDplEPcbXEhrHnXR
Ft3QobvbZYX7PUmWaUC4GlYChPac2VYq2zPdO4IaHIhodBsFL3OZuthvhn0zW/L0
i2EXFHi27rbNeaLn4UEOvVXhvG3Gnt4RlyvhWzEZCXqSIfkDAQKeWxvl7zdLrv6z
+qXumqiK345dpZ2vXxk3yJDBho5Ew+22JoJ0+fQiMo2R8WnOBoFvEXvMlT8N3yPG
Zbws9Izckn1GHTNyIaIqiFV28oEB5PpIxjaFAJ9kWmmFq4+vSInLAG3JxOnLUqYu
ALiIfpGxA/0nSybDphtjcyMMgBpe6LsmUTqvpdhEjq/3bI83KdI3zi63iZRkNA5o
PFhHJIneDF6qFqn3NWIJOzywT61Fd0bpqrDP6boG641xv21V2X8x6xL40t9uhFVb
Xl36VEyyITyAH6jLvoa0T5aDNS1tG2NGChf+mEdI4pk+nI05IzKgaj51NWEutnqM
8FSxu844Qcy9rygIs6kl8M7eVmihJQ5nr7py/mY6svDbfETNj9R/JJ4tUtwN6b/z
W4/9cbkEFnNRXPPF+cbP8XNQKKf6uNzMVRzE1m2KK+V8X7druF83c6UAXjjuSjU7
OPqzmYCSvHCjJpNuF7DvYRtaJ0apvSPwEj85cbklPiCNXydTH/6i/hBUpCr/O20p
yLx82fI8CVPKjYezgheZpBzDN3EVhymduj0PQEvuqdfu/0vx1wD+d6+YYMCBWnuv
jNNn1lL31Zef7vIIpONLdEV8okJ7zly9WxHB79UgFb35OGf+Vgy/R2+vAsy5lBf7
MKubWOI+aKkEyMsJGfoFU4WlxdLvm5ggG9ltp65XAtLuKzyVI+ddM8da0oPo/J8G
ztCD2rgFX+1tSy2rAj6XwESu8OySaaq2UO/3aZcyYb/u1+qFonviM7h10oYnlYRh
7OD0S2xZTlrBpKeG3OCs+xqw+UJ3e8cDnSCpc8mBHjbGSpXf4J8jJDjdwMyo1L3u
BodtuvtzZgyCDubZ/VEpqUVRVtqLy/17BShXSnLGNWX62qT0kYPXbpZGhtWXijEc
52VK9AzyOjvq3PmNAZShPENN88S7oetbfnLw1oygFapYyitQeimkS21YsUqHrab2
b5zBLksiHp/hebZpb9dxBBOZPDyH8VlA+9nzLUrDzSO/if3brUjkfEtlQLX44VdX
y9oCQbJQ/Qof8nRzAgZT4InXSXDLt79DFc3u2OKGgAo4Qg9wPy8ClMQz6w1vTqc9
vZvZBSuQ9iOTFu2bguFYcoYtg4p5RTooBv2Fe9hWtn/qScSIDVFrECinZwCmwLwh
GvmpixAo8BwD8lg8Dr7v4mUsZmbo7bgNTcleUXJsbdBr2Wu+cIbH4iAQpKiuRtFL
VcNXkliEUPVLVJr+oN1h8+tv/r/6tIi3hXh8GIKqOjsJ4tARcaNidRiQ6svsR6aI
p9GBc1vXaPQO7ursNnu5v3IT1UIqfdv2xAu9dz2vY+5oJcabVZP3NbDvlTAa3EQw
sZcV/sl/mzUX4L3wNZn50i663dXe4Yh/hTBcGfXAs5/CAOes5V3qnq8ypMH7ki5z
d4N1CJaSZEvp3crp3rqFJQGSG8Ku0brvvHnddvWPdOjBE4gn3D+SxhFZGaHbHQBY
P8aw3CDd8FGlgrtEoMMhlyqV1qeIkee3KKzweoPVRW7PXix9mtxxNjT7IxMxcthT
R8b0Q+U0+/I4DB3jfmvt7f4g9px1dSIplTLALda6C9ndutPgtuuiGyHsNTppzhHC
8rLvZg/129uBB97s9xtxXHfyBBJDPLofd2HhIhCS9EvMERX5BJb3I73CGuBYWJ/Y
a84WnDPINOkkglz765gkefZituJSEm6VicckINr+hsckpMVzhwfnifwYCWNTRRbo
asJkZNyC5lIXA4UBnsqrras2Rl9m5olTlatlDAQTQ+j+TVBwa92zA5NYqMEtAnDA
iTNlq/G5phvN7GJhVUI13BoGf3dxFuf4NsDM7BOmffF6GY4Xl/JdA/L5gmnuNg5e
WBEpC0fG4SvuUroaarRbiZ0Im2NHj2/BeevAtPDpNOGjeFWxYJhN2fPqSt2QrNKu
ONUqd+qo5rmm4MMuAGAIZrKU7j5ERwnrcOfAN6k9Gzn3RpqdYee52Pt+qLUEb0px
mFWg4guWBWrtS8lxtM/8sHF1WBcQZFE/GekM+OM2KnTSX4rdZ/VNbFBuuh6O+tRE
cw5ln4QtW7SJp60gz29NXfsgfoe+yN1E1B7qM+ZftAtzQttjVxPt2TCVZP/hC0Tq
98s7hs+HwOtgmBX5KU/ADH4lUuakj9fqiwf8j35SEYUu0Qy4Vp9KvTdZVmUJWqUm
hHiPmfpMeBKa26GTC8jUYS+vMGdw6AttgeFpVwrNZ+rHCB/9BYY+FyDLJSHcUxzZ
kYgW7RlaRoy37ZrgnMYTDapbk9+p5ehFjf9oQ9oc7htylhbEyEcD7acMXZ5CIZXE
15AopMvWnEpnQg9YZ2/pR+9XDn/yoTKulGyQzl8LZNOC6eFzzm2F+FZNv0pg2u0j
wbmqUmAouDVZDudtFvz0fQqaRABHgfkeMxzm9NiUDVq88t/HkNTLt1TBUyYyQd74
yZv7pmP2BOv6iUD0851+dnlxFr4MjPMDlNT6FWMv1AIVGoCOlvAaax0vIOyFz4Zz
JeyzlUCl7NIAZSIhZ9yDoocK5+AOFWbPwGW0aMjaVxIV7C1DYbGUlHl8NE5F8JFP
FtIo6JYdjwbXbVFWnkJqPKLo5Mdl5n4zUuT6xJLpJsjiYmLHmVQETtmgEFHLaO6o
5zPe4AEc5qHsIlkRpZ9vZlzYwX6D5a9Dnp2X4ezr4futYz7wdUdAkoDJMU4783DP
4h98OaBY/22nptAXRnJbAj+GkCN0fEb/Nd2RisTvFRwF4bVPjXlk4y6tXqluuKIN
hEQoa9FAYebH3pP7IKM6JYbmm+zkzCuIobUF9h3BMbESaTCl3pt7dSRqOyOblJ18
QFD6k3oLztV2vSXoBiuGZR6gI5IG6TvmqWhMr0BQXv2UM/u70Q81IkJb7Rb+t5/z
tA2JFXCU9MLeEF6MPYNg2jm8kpqO0cu+LGYcQ3OGd6Hrx5b57Tiqvp1DUahj12QZ
3qtv/FyC+/cWUKvuzuEiBoQcHicyJXj1PZFjYVYqEUpQ8O+wztu6BVeSztAbB9qh
TbdRP0KtsqzK/W0+fKv1rfOs+8YYxQgiLCFXUp6jUbs7BuQGbFOrdsLN94V7x/KS
vCq1cf/qoId8CxQ/FaYcU/ULnmyRSG6eHjFwAxXe+hWJUA/rx9uRMm8IXF1myYMd
ZYFgabg0LKxc6rax2FtyBJnTExeJNvnhd/0Z+p/j7hclGHLhgqLuwGulRTqpP7wm
Z3OAcqVha6ZjA6GpHA+FUJrP/bYYd8f4i2iIo+iD/U0TqphnhOfVsFcrh8cUKJtL
dU6mX+5f6tQZ0TitVNo4WvsnZBHLKZE+nqbG1PuYeW8igxL5DzXkg2ToAoqIOmo4
ZAHjpN/dS0sQa2XuW+o5fv1yAaG7+wp1bzqtjR8Np/Ce3nrO/Jo/0TZJMbR5+qnZ
wcjLDde2rL9zBHtFjLbZuyohyUigWtWS2DYOUAhj3CjtEtHzhK79CS8mn3bj05mn
nGpHK5or/oD0b7NXjVpmN7Yu/EV8XUWA+bvzCn5VIcDfrHVTVrtTGO2AIjqf7AcH
J8xUfD8sCnT9fE1HYwpJmNcrljKHs0HVlfSRD7zZg4owIzjFghNJO/gmfp/b0ssN
H5p8d/UW5icyuXQbSgT80XX2kEGkfybb+Lel4fDY2dhDLOBVEgnUEtGELUM1It24
dPVX3xqCvNLQ6tuaMKEGe3MJZemiIk4nTsguW+rHTyHkzHeHDnsiL/4G7eLDnVWE
ACvjQ+StNlWZrLz6EBLXh+CmcGuXLHtzFISsZ/8UV7Y00QPsqTMGf61yWJ99Lu7E
1T/xNhfA6CouKP8KAw5ypJ2hD+6cwsNMkSj2cTJ2/eSgTDvJL2xkqhlt9OO/GWji
/fApfY8lUFEIi+y1G9OxTyDIZrZ5Uw91FvjykEMDADHgkdi5891KkBPDqCbnhLoM
MDhdA08k4uM/LUAKKeSQq5BFdO2DhoJP6L/jwZFJ4Iflc3HJLxsHQwVG88TxsEFM
FZpryX3692kHJP3t2GLyMTB8g9gs7okrXCtY95gVv9AaUCxAzcgj4lx0UcK69KnF
MBuCViXKOQO+NOrq8KLl1mtzGe2nPW8U/8Y+R+eaFMIDr6cdFQRJJiN02IClA+Y/
4LdrzVPsFsmQdd4dJSoJc9TyfpSmElFHP1HWh55lZ1aHeVsydJcRZLnOWMeeCXXF
zllDe6th5of3Smb5I9v0mOR/yO0Lhh8rQZD83u1cIgoT2LuPlo5ybX5KoIZjOdyY
Nol3mixkX5QPyq/V0Bgbv23kwelmgU7onVV62h0LFQhNMgtvqqqvbuWi6dhlfNnC
lZMNM1qLSad5TF0/BXeaWZhb0bgJyUZPFWjZN52J7MHZoi6mgHMhMS/j3HfgYZWG
qb5CrhGS5D3wwvIY3KuO5ryVNQuzUxoVHPjRkxmToQmGb4XjbIHSi1C4xM0F9pil
aDQBoFk5HJZ8QvtUSt4Urb/3I1yI+Z3OsVB3gq9wTAk5M2an8d+QpDH+vU93rfp+
iaPfWiZCiwYxTGdVTlLadagLCzYk7AaKMnue8FKc53HDeNE/3UozfDfTgNCqvGcI
1M4cV7TIDygDs+iL8bZwd+nRB4ZEKYRkop1ASMpxu6qHUoYmfSQNKMwwJ3N32asb
rk6KE01WLPHSXwZWsd0Ffv8DmEKP1+4C+8k4ZlcVchWxvUIF3tAjfrKybzApz7M/
Xy2jOb3wwpvs53lRWgiBwlcabVug9elf9i+DmLDIgvnEDvSgO7ILGCTLSL1tNliT
znu4vtxN9J8bgJmka9Kj5LoDUCoBqZrsXppnutlMFH7nTJJ3A2EFMbuzoedIYSz9
zv/0REoMwvc5cO0dLN6oDeCKxi4dzK9EKOqE0HbZ6PpwTLzCwkW1m2c9zxaoT7Pv
YIpl+BLuNSYGQAPBQ4525p7zDJZw9fRcA9GI0+BBw6BQJbxlqMgp8EMW8ileULfj
7s6RnHP/6w/d/CBRrcygRuOjtJYWXamax5GavV6oex18IwCsLdNifIjvmrd85gkg
h6n6ZrArDKPzaVHLkE8yrGQEW4Umy55mbhXvTjMr3NKoWVGgFKFeN9XnZI4Q3qnj
zVdaNjBoKovm02yF4lmcsTNKH3O1RFC939cKipGG1P8HX7vJYl5z9mpLzzh897gJ
TNF0aAnjCANHrb4ZVhYBvRhVfKn7gCdpoLrCbQdsc4oTeOaiKbI/rKGMt//qZiZ6
hdTdHK6ZMyb9zA2bxdjcKg7ogx/oakKOCV06kvxtlKlFx5qIm4ko759jDHu7+PrK
6QuasLovhSU6HWdTNn2YT4Se5RV4rMmd5s2gHimL0PmuGWYQmWxA/KwO9xkuRs8P
i/Z/XcpLifeqa0c8nf3eWTmaYd6PDLIm6VKaTD/wV2xCMu4G00deja3qz2bcFJYv
pikMSSwo8UJAd3Udd2W7ffQ0qWt5yAAVE2KdiVMYej3L/HCDY7gYRgnQTQ2zJglN
lPFtTRHULpyovPh+DgZJjAzV62hSENBzrGbjNiNoCotsa4W7on00vNEtuj2MyWnR
GIJfS5rDps3GHNrqrZX4xKtbfr9GaNWKL8/R4O5cc2p2xGNvOokuPcawkrH/lRuk
9n1GfzgdZvKWeHMd1tuWDxWVjJYow4Cbiyf6tgrG2QkPyYm20Bk/D2KsBfMpLk/1
VuyrjS3Tye871bKiT0IL1SGtsoP3fEBX6gKberMWjJQVU6cMzFPs+MrNC6gRLkVF
JFBtC//EXcd/7CgIUXpZ1h6BrqhbtGOUB0pUwZWy6gdyFQCevsmrPNPdTpFgk0gz
xgi6mQlguZ6PwzRSlay/1E+HRzJgk6gP6VhDLk5ISZdz5Py0BP2LJURsmdMcoNGX
U1mLnpXU8OSD6sQp5irXXAjHFq3zILQDZ5pcYh5pIGn4Dh7fT9KZp1kKrPwxNdSQ
crL1bE1hP0fGDJg9ju5HrHax/SiykELfm0ZVjESSxvZfRzx9zTQ9LBkzPOQhzUig
PodHyGxnFa3vIDZOHPfZcZptiA8DDXsrRmxaIeP319Vzst9bMZekt5Rca8gFh+uW
TKYd4NuKNYJ86w6Kro1myB7qFhVAT/+8F8va6JT0Dn5s20XKVSz3Nu/57NyCJEr6
iVwF2OioY5U5GdUcQhSTChI2y/KIs9bUyEumyDZ9zuqADu3iCvy+W3wqYfweVPld
xQJdHEQP/sEvukKHIDoecqLbKB2rdCnc4GUfwMlUdGAlDqmp/GSVw/Nzxrtr+Nf5
fGv7Io7mlM6Lz2u2FN9jratMaABHQC1tCiBvJ0a2PSi6BlzgC4SMlI51c2vvIUfP
O5oXqnZtrQpYkHVoCgmSqxq+KBqxRJtpYyMcMy09w+dYZVfh+YB5QalzKoTUqQlJ
uiL+x3sDy5kjpxyselISj4kmue/CE0TJGzzsAcXLFBHAV2stihHZ6C0ULl1fCqLS
9NpmXOPsZfkxYZiX26L4x2+hrnVSVJd8UyBsQUWoHO3D3yOiprYw930UpZdZLH1O
OFMuFSqjlGRxualOcgMouhzs+OvElKpgTZWs2mehWsmbxos5344viv1daIvkLOrY
qquHuQBc4K3dSvaP0R4Nf5tD5o3n4EWbS8zRUZpI1z1kMtp7coSVDZR/2ymiGnjv
F+51OW8OoItmwa0n73sy3HmTOGJ32DWGJfINX0E3W25ymyHRFMd3fLCP4OC8JzOY
U2QE5i9e2Kn8HIwlj2big7hudCWCmH8Kv3m1Na6dGjii/OIcn0RMfG1mmUjBANPp
cF5rs8lRYQT4UtnOxFh+Ms32YfJl8bZtbHVdb8fe+01unDNl7A5mIbutubxLkfnk
raLsU2sMAMhuYoE01Ruu3QDrHuaIzNh2T/tfZ9RkK9RasS0NNjai+aU0UIcK6xTB
EuwSnWjkuFTwU+76nNEE0fz7KUexqpOnMDzk1Vqw2DaHx8iUweoJxEy31nJKkvCs
oCBME0GQbbnYh4pIvAtU6wbqsAKvL6Gdwa9c1+/I3phCkdmnFzxDlPUarnQESlwM
npdDWts54yN1nAKPkw0UAmCQYm3XDmr+hS9/UYLKMEBvepz9/2y6LsZKrMaY5nDD
9P51XvdzFRZG6fZnUus6Q6pmzF/GluZkRuJX7r+womoudzNbKShjFzUG109dSO+F
C6uwLjJOg+f+NoBmDn6dF/lJaVfNSBAKGMbbeduoPojlYjBksVQ27Za5OoI4pbWR
MSbNpt38xAywT2PMCFbkUXIar6zi983d/VDisTH4VXwoee0rOoPpIy1FI5T6AUmg
qkLwNmsMEiii1hbXQciMXnemMsxXB0iSx4lFoc9LAm8MUDUEiYzX5VzHVaxlfITq
0YhL9SmMEqg09ArEyWk6QHLvw3xAVHgxcib+vT2bz30ZrmDvFJjSxzwjjYkMMZE+
RlIPH/jz/CR78bm2Qd6QqfWwx8bdFH+4iUIzli/mD6eLddE587tsjqMuHbUO746c
8Huewo0jPUcXVHjaHgMjZh9G0OTPXXPBQmacL0lyTK+ys+f4SkxNiP/KeDrFJX5k
Odv3XYcBLg5gG9NHPpbamQQPGcdl+HcEM/sCtlElC3IA0z8/6B2id7GPGvAveSQY
GwmTD10yOy6LuFRk6oWJAgha/aY1/CeD/lIkSxL2vslAD1V2mglWdXU3YfpL9QIC
3DkbrQuwn0iGAXcA9hnSvpnaoxqqXJR/cR4i5T4Ie85WlfZfDSO6bfxxGcX3TnZv
i3YbvjBXsfeFBve4C2w3KRcrnfcHbuYIhw/voithaOFJI4G/n7PBGaEV5JPjluea
5Ll82Kjuzx3rFCEpHYV4wLRadK9EK0zLyNifyOLmF8A5+pr3u07N2i8QgrsHfOQg
A6BOsRiggA/l+8iN/zHOqTBq/X/8aKk0OgvPQWBVW2Rcby/y7RVaSVx1DVbFLNUC
UbWqoHv279MAmn+ix10n6qfZe0pSWDCkKil8NQQwBmvHcoU063yhFHENWnjIB/7b
N0vYsMxuEIoaES3ZAQb6amdO5WhBDMp8qpjYcZ82CvT3SnyOpUdEA58OpZq6XmPD
LAKpnDbZOp7wwvJ9h6MpA0xUNpKJZkDazZ2kb2o050gzgWRF5j4bLO6SZWedeuo/
89ChAkJ2r0vYzPEVdhvEeBriKcOvdFOzYKEua0DudQZToznr2GQT4kqCOu8VJYpb
5gL+2OjkpTg9XeK29grdJfjNmHKAD8PAcWDOCquLmeomEEDCUHOn3vk987Gqd12A
ZdQFBqWAkHN1bkJboI5oP4GiTFQtLbH+Pk8ECoElFUMpFOOgbaRJ2tXfeSug+0Xg
ga7QEd1dZLpGiKdxQbG4935vEMCf65plrfRUKoXLPdvBj2SGBkQOqKAJW5IVfnNQ
ChMjXMsG7nAJj/fg/cmrz7kSuqedNzKoAf92gDik9icvcxdC+edJOpwS2nR48xvv
LsRF4HbztBkPFU8EhYjubSPfq9kd9qe+8Ca6EGmX8hsvtrsd6BsGA/MLPbMyYuzn
O2WDXtivsL9xSY+H7YqNIWTZQPiF14GnONFIMRWr7CrbQlqD0QSnAIZa98o5ekB6
ILPl0j0D9oMWasjfryYQEIF1GO/kmW49FChVT6PGCX4YRr0TOfI/CgiiYRRsZC0R
v2ytY+CsH+tzYmZMLAbQ+KISmIGf0SRoyFg14k4pc8hnc/iRlpieIbE3MNLlN7iD
22aDNBJbwc99Dt3lRMUlHhB7UZ1UoLBLC+PRasstoMOJPEixfLv9/O04IBAQu65P
fdw0pZC5GScdCVE0MrSpUxxRBe19gCCQrzPi+uE/l1aPVWnlZ4buNgN8oD/iLiy2
NjKv92HWmjcqW2EA1ZOVjemWy/Z+f5Bp69ioJ+RsclxR0wE4pe8mFTfUbPS/EQLp
MtLQ3DLkqlFPMIogFQMBx1BkvzuhDKtyn8qjj5iXJZm0TqagJEnPgYLjpKNfIwKs
N7pfAdPcL/XGMkl75U6NTiFUeunm/R3d6HC0kKEw6H0Gp1Zultfkk+oRZOyWlSAK
x5VPQmpxnLorl6hcPnywbFCBxFfCaX7fWa9XTvpfAvIcQBWKk8mGA8LRE+VVmBnF
96V8Bf2Jl0OTE/3xfnTh0JRTkunwhHCAQhg9vtPwygkrQGlUj0Jm8NjCS1xaEGam
Ad+kii1zeaVIlMKTTDxCnf7C8z/NTW8JP0xI9InKkz2mHeeZEkZEcG0s2HITbcqQ
In6FnRuTzOMft1rHwrK9Mt+cqr8KDh/8qqcHjLwrA50fXNDHSXHW2RUJjm2izdr5
lviXf+OK9veCsCzFxRU7GiW01yz34B0eB32asnyvZP1AXGJWdXupUgiiFLS6Um2k
QGW0OjfkhHyFvENVa12YXj350M1Cg2URH2PiBQ5yLsLWDUtB4Nv/YE4AZ5ZtGCEO
IkPTTrQ+1Rro4XUsJXBm16VmCTgxpYwdFtOfbyB68zl3UrPk0PSpGJ7t1ANrXUqf
6GgAkYRbHcZYe5F1MS66wIg9qu8BHkmsQjM+MFMgcAS+UUhXw5cQVJZmJ4Tm2TSN
CPL1LQZzJJrSoYOp5TGs0cpc0uxag3VGbyJKhPwqi37fjSrfT+bsFOUpS+mE57We
ZEhW6W6CdUXydBI1t6F0lp9av4Orpn5g5bPw1YPxoogPyqG5bq6uDMKG023PngPg
y4B2pCFGVDxf+r+4HVOKI7xIx+rHVLNytnn9V3cRMzqRdk1MZhAL6UfcIsQPlJBK
dRJP9ro0BMLNlWKNb2uw1qAkTYVKWau6fa8+ynivRvlpzfH9Q5RZNUQxETNeXLDI
tPSD0rQebBt/hrFm0ZA6fNRVJl4d8gbpNscVPaiDR9eFGnljFg/ZK1SwVxl1Umty
QlRKSMSjAV4pQUFufGUNR0maG8EbkH7Q7kmOhbSrwixgG9W4kRdkpsVYydBFI1Ne
zTc5E5RkAq4SuMn48gA9lE8gY8DIqIzBhWkrW79TtTvxCGHz8enBJKZN2nkl3Zn7
l0FUsoAwyhs+gnEb7DZLx7O6gGpjHILOhlBAkz7ireOUrow1MtDBiOSPaJ0rd0Za
QW69IxTF3RpWp6A2H5ALgJq7JhJz0jZFDAjTuV9DUfVcjpvku8GAdj0KUH07Nqz5
bhn17l5da1cjNJ7ScGHJQnYZixTmRbI6NZRry5pesHN0Mw+E1CoVBd3QBrFrpcA3
9h9VjDc3nfErStQoXi5PBHmRPX0m254kuKy2wfRWWM+cMz8Uvnuf0RyK9XYoBS7x
2vxa+OrTC5/L7j3TyYmac86ENrm4h3EV0l0scd/KGm98Ba9uxA9JAuS3kpj3El6p
peWfRE3YMrETY0aMAzVQ6WHbxvjlQBrJvYDTLQkt3FPcNe/2FDHARMtMoRaj3asm
yX3qwY+EeUGK7sladPH4G3mzZQblxzU+8kcNvk2tSkqfHIj+e9PMnXmOGAT42O5g
1rxL+5nbR9/hVNDLQYrEbIAh0R+T4QFWrSz+VTaBg/TmwHrUS905BBMxavs8070L
iihHa/C0ODiHnASeoR6mLGxZS3OtOtUyG3x/q5WmYFbxyoVgBQTPN5bhHy95cZ7n
VUnt1m32rN/zcHRbyh8kBqiz+hHlk/bx7fr/BEVTYVv49UoWFTE+V2mxdl2ROg2h
WnqdQhHbVGKSUxCOHzD6Y22zCeKew42Io0vnr+0GfD8LibqZbrx54slFEnZAgLa3
Hqe6N/awG8Zox48672Aeq8ygYY1LAMRhXyxgIUcuxx/eUpEE+FqvYzMuzCdKmmV8
5lgpyAdRN7f2/5hCS0XJSYcefb5rMEbrKmFFFx6TfFXgXDCpqccP0yrTVBydV24g
3sTytaSbPGVfdfhvrqBMnBee1YEPg5ATRDiLRutcklW08IBa9BPc9JCMw+Ve2rGu
c79GWftwch7DE3RjzI7aACo2ltzcx8Ek1fA3+bixWyzW6s7VVpAdfNEkJAcFrKNO
eY7ERrTEFkzYtGHOMRAmiB+T7sFDrgnLO+wg/3R5OX+I+4Hd7kzvzLCNsgQJ8Cx8
9oc0/egcjnir2Y00X31oybozMXjbzvhvlaqnIoPOd81zzP49fB4gOHeVt2cYTi6e
YAlIQ2w21UKvztatSjQyexQZE+44Ah2Q8WEXxfILU+M7LnRd+OHEJiitWFCVxXwp
+3WXOJNkg2bgPs5c/fI9DBhgtq9HzQc0UJmeU6CYNDYCIDyt6QgIMj6dAPDRnVCk
q8gjRn+cbsre+0gsKV9F9Vksnxa235kw/BmgYu2czcp0FMFxuDECbcohgw8rUqaD
OpFGE4DS351t1iieAIWDv4h+0byO4a6eectTLH+6K7xOlJCzSD2IzkprLUKKstfm
+rEn7rUduZxvxsKyZkqNxs8Bc4Uxb3KyRMitv2gkEIFBTyHkJA0xDvvTwkmri2BM
bxZhqGAzBcDlJvqQ6PmYKaT5okf1VIfrBDsg/R1cRgc7zdA1DjZIEhRCJ/sGKjjE
COu+5HepGP1TdeDdxAsISqhqkg6U2nIwrLLZZL294KhHgYlAZuk3j4wCANUe2nVe
/fjj9CqdylvKFVEHCpQkNsHT/c+kdPHCsjl73C4vNqEGdZRQbpj7N2SxzldItOCW
MB1JLWyECEQKD3Q/R4bjBQSdhEOAR+f9L6IfX2T0xMzUq1E8PNlmEE5QVH3KKqcE
R66Bk5uU5J515NDq7j35138F010pDSzMrX1t37bVLgZXK5H44c3kCd+q7VyzR/AQ
R+ji8z4B3cS2y5+LnPKDvvdVbmMswuFtJ+unwKDOvIRDkJ9a2LKZY0A6CrvqJOla
AlaH3Z+I6DGnghb0Is3hVUVUF+3Xut0ajbYvq+wWTboz6eCsNhHCL0xmUU9puZdt
OHNPipPzNchpu2UU9pTkVGKgTWRHshKuyei6IIjJQiI/jbXDisun0yDRR7W4/dvs
XgBr952AYVST4aiZQ9xcv52nlTYAMIOwfQ5PD3JCBY6+141X8efnl6nAYGigiaEG
v7H57+KUIx40eHwO/u9T5nq7sJfeeNBkhO3EYxJitxqC3Tnsi13DevS3sRsvHFlv
yiVBjvgBr03zC1n/RirVqU3gySEmBsvj+yFDXAW8z60p2ZcBqtYGlVrvbcbfd+Sd
57/FD2XAEM8HN5M+1yU6VYtY+1tQBrTC5ch1SDD/bIFbUnij2bfR5VRHKg2JI18c
uHYnzZHVRy6FAgSHRY4NjBlHQDviTXaVBaXWLFLRSkKZmu/WBlNnCbolKDIiEONs
14kNblkF7DrD0y9e9Whx/1kkX6MjEC8LkpUtNJhomln+o9VAZVdKpffVurHbfApi
wUZlt3lqXss6mR2lXEafRJ5usST6JilLic2e5zxe4wOXs4a+Xb71r6fq2b2ZYqrL
vpmliRPQSoHEFY/m//6oQUXHh6/PTkwKAdQz4D//QFJzrj9eMjmzXEX3CB13wM12
Cf3cebbiegGCpFNRG9caXPrRWA/WND5hXtF0p6lpF9AK0CfY1yoQQBsTA0A/D4m6
YxByJu8Ul1YBl4nNkx11RGjlllwc5TN6d9HJytN9Rl0ize6QKLzQaYp0Ds2AwSJt
UU19xb5p5CQ1CQuO6SyGk5X1HSCsF1ahxlyEogZYbu6KCkCcgyGe3RI+TMKJP1AC
KPItwsIsSjUcFlPQ4Tk1G5+VebW0NbY8n34xJbHpXq1TS/c8SUtJmm8n8Ih247aj
2PYcPzmTwph9H9C9S5xmyjIR/lLoZABfxLrLeQ1vEBOp1b5xduGJ6bOHLryTq+8S
YRNzmbyBwqH5m9jJpDUF8SbH9qcfwu76d3dgu+Gnk756JarwVnOM6flcUCKoMdGX
AwExnRQvyQnf8R+Ules1DbcCun85ZYYYthXcFlhoWg0BPFhyN0f25ps6/bJNUMcL
rna/gQeLkOEROzRk1scm7Wm88sWFFRgdXwDJLjY4NH7ya16oDbRbo1C/T1wpap4K
nSBc4d1NWwSw/3mvlJ3RA4G9e6OLI5jVYm2FSWm+iSl/Jd37T9DsfFaG+Z+0cKoa
n9NezrZTE9XhMd/OGqZVl0B4IYmwQ3ET6NqCHxGlt5grSmmqAPunPtYGiofdweYD
Ns3jwv4D/R6yf+oyuFPX/nr5sC+2P2JDnsEdOLAd3+LOdIRMqbWmbgiJUdwtSK8t
ve3VeWoGwCm8q+qtdyTuPNqXRzxNkru3Ke3i4kFqcSZ4RlBUHA2nYUQmA171d/y4
tn4S+M3xFBkPZI6U5yl9+RKwMs6qA8JVK082ddvdv1PpGuZtZ4s11OYrY0gNG1wT
w3CYAXKggiJvojIBI3NLgQ0Pl1L9uln19KaE89Ga1BzLCoI1ljiZzPEg+4+Dh59W
C7G/fnpZrLpJ/n4gJIIjg1vAGl7rQRhGMhpflbQoi3s1eJakgxzUBQyCoUCQ+Y4r
scVRG4y8DwKXEk9XFiaKXL+8mRl6BbBSN5qommtCrYIFhakyMNt/xuEc0z6FkdGW
cOL3OYdMKNw9p0JfS/6qUfh3wwOCP39N9F8TeOOgOGtJrIgZ1kIKn5D6Uj7uo0yy
aPDNs991JkE8CcOwHR/AaBTSWIJa3/BgIzMpAlm71XKizztS6amnfni6nZnlhsnA
sweUpPlde4t/unmA06KAxjxh7eZchBt1zMsjOwFE6qKhKgmvij/2Hd08FLYNQ9x9
70HB5iiznknWNT2Pm+sBCmoBx7yNF7+SUTVfo5Aej0oGjPe+X0TL4mqaAIB2HOcF
YLu+6kxrkm75hXRvpvCKCC6tHZgdaAyBrfSYvwHzanD7Jlqxm0N3HUJPcxTBcmn3
xyKcqUn9eXod+wLiVMPyjNZJvp/neqAccGkRBc2KUfFcvDWjnq58s0FFUCMrgY4D
55T0vt4ZGrjJQx5b8CnreQSzMp8N29WWf7AsuOnGzJ9BkhIqzNMpqeK1tBqX4FJM
7UOiVkWdFOp+WmNhygByZD9tV4HDFoP4T26DtiPTTJdSdsgeVHfPrki3u2nbj5e4
TL++LIIR55ajlJoo01KtnoGcVm1s9MElBZjE8rtQkUwuF6FXMj4dHQaxRoBrQlIL
6EbLanhKgPlrJhyWqVCEAvttNlxm+qyLVd2g0Y+svOLgWhCCVM8B1GyL6aane7gE
iHg1MqoJDs+EtuSc9Bk+AdxoYoiH/6UHGlAjyA9eKHuIQeOpUzyGmbO2rRhoAlZk
8saZDdtOEmiONSkk+LVp7kQnFVSgEUL95c6X/+dRUOlhEzGsqYteq2ym7u7w6ffN
Umxn0afFCMBQt/xYdBK3VVl8PyACmU80dAEvPVH10GBB/TpVbat2nAeGHprbuxIt
XAsozCKyHoJ+9D3cTiwTa+5l4+658hBjCHGRjgtjeDGJ9ZumVba/W0388H2rVxL1
lCXqcTjCiyWoDEMwyOaPmgYVP0wLBi+iQrxjJxnTQ8n9DMuEjC8QWN8m+H8aOOEY
71U8gFPktdwbspE7u16ozlB3OfhJIfUnJT4uEMUkZnyh0AirsEnMbBT1TS84tuqh
UQd1QJAF9TTHiyma/gJSwS9e3/BsuNyOtdmq7dy3N2Mtaaf/9YHQUmr0MF7IPh2F
rpEwDaKd88Lff0VLgb42ygVEzlJ2F3D55M7swuTU5nvgEW62WnMjfM8l3434GA4e
wKtVW0O+684aBhBjiOQO7FIOTDkoGZ2ls6rHNsNKq56RmyL9NQTEaNuK7uYPVXT5
LB2g9r28LsomawOOIAF5JUw9vm98rEgiVCAuyY52Wh/NAw5PzDpQBwKN8L0+M3Hz
zSdR+hGrDLK/CWpT+NQJcxL5VvWstHo85WrEZUIbEn8q5SQZnB/HDlE8yihjkm5I
pHwW9bkI1gT7CC6Qaf8JWsHpp3pLllerP0GU+psRFe2PcbwSPKebZGCEqo4wOS4X
gxLa6UgwUpKWX7cQrwymsOvj5vh1T0r42VCjdEwcMWcLnPYmM0OY4hZAsXuO7mcD
fcIVlGyX/fkl6c8e7a9bu/J226km5T+A0mAS8q2yZtKp3bXV6Zn6TQgZJcjuJJ6/
+3ksnIvtDP6VeXDT47Ncva2pjPhgsMUwgSc422xulfirvninhXQo/2dPYKUBxal2
JEU9NTwo14yJ8jP1iLFtxazoW1PeXXIo4z1+zCc5ZJPQaM+tS/FRR10FXjvtdJJW
/9cwsZJBMtJRDjxOWiYgQmcJZORIWqc9puW+ElO4GKDjG+BHlN1ctEhuQq5mvonD
8zkstrWaeg+t4N6krBSdRnntIkKndOiC72bVr8vRCDYAEPzpCubLd4++e1jdmxgM
ptzizQ2Z3l5JzW2ScHl+BcDQCFtMkcyzNUcHbEwUPmBNU3vcnpL0ytBJhVAd0o11
85vcd716nGASkQ8vzve9PLZL4jK4DX9LxWWcviLHXWYPwi63rbp6VrHA+PLAxiYv
wC7uHlBrpnnmmI0NWKYR9XLs1zicU2CE2BUXDIPhI1ayp0nDo6Otp14SnLt6ZZkM
QyjeWIzAKtU1i8X08B+yGA62gGvEyu0iM4fugsPZtSHJRnLjO3ZS2CNMTS7gBnMo
hkry0Bq2FL9pjuObl/3ZbgjkuaT2DCscTnukECnkw/mCfwkvfgMmwjkaYDgkVZvk
1n6VxPYGlFZKMscUqmi67Ow7KOrGPMgEr7fLQ99pE0+wJkyOG+d9VIcINmE9IzTn
6rkajsUB6zfjZfAhMaWjXyn6RZ3mU9cpd09bqqZm32njkA4kCVsfKgtIw8UrTet8
A5P7Lhwq1llRuyAIZObxIzmj6r+1jwQPjgQ5jrqAKgiZ9ZLtyEAjnIyZ8VmNxQLe
MCcsV8vFXujl8aEShTtoPxYZE2S+Nrru+VQa98rGOspcGKDzWp1LATuXU2sqK9DA
/ka40/ekvajajxvBJsxYkk1vMpS7fgQDg1xVSAKm/09Yhd+y5ze4kWXCCz3PQH5O
YI4B7g/y95GDOp21iyD+OgkoaN05QDwnra9vilwufvXDdxuyc9xi4K0UTBRED/vJ
L8Uoezz+jxieaRLSPHXRhz6CFEkbuMLYJpNCK1DlbXmmBGN2oxX6IgcW4NdFp9by
ACJa7N+W7kZ5A4aE9DTsz3V2UdkHVuOLurgeCB3pf8L+Zmz+p9i2bULxTCX9DMsN
djsWhy3APtCV9BIRrhQKsuf796TmdmAo02xghTGhusxWGBCAdGgLGC9I/i1EbS2c
EwouFfXbENFe3w6Z0TucC3dwx9ep83g4TrAXryhI67T7mM+WFExX+j9C9Qo6ahCC
Ag0fXEeNnTtR2wHZC8nh2oHdSw+ylX4FS1CMNcXW8bY27eZJEkEqlQHLlNTYl65Q
Of0s1szgAUZV2OT+Sz6/VTSNdoOPsUUKN/vXwfwYBai1iTjRBF3Wgra52CuNhZlz
1wlJnhH9RCqp7MnaC2vNxgLrW3hmo5OxKjchVshHayKo3/Ybe6DlSW/Px1lWWpDH
DhZHA9QHsyklOzNchQwyezt9W9bsAUzCVk01nbHx89PjgkmwALVsmEx1mXUrobQ3
9lqMfrmMBk8emDx1m7Ga1T531g+AHBK9m8EE7SYGilkAYgmqr+k1xD5nHUOxDqkc
5vSXPZcSBRW7hoIHONthCY/EG3xx+ZjISQLJlpXsnX0DS6WLJUrZs7ztNuFTDKJe
dmJiVh6BbMklo57QziFqoPaRzt0iOqq7THigYeAO6CNhDWqhELq/Pta7le5w2EKE
g8XsPBt/iFaUidkAqLngIKbU9vxByeS7/FEmrp73iewHTfeE0W2hR4MPgedOgXD/
HarbGBtMiwnjOupaASCz1PdHNvsZUmr0Tj7vAF2256Xh7MZr62XXTDTgz5wdg5Sg
3ifw0j8Cl82Jv1py0q6Ax5JMiVik7AR4lzqJ5LAsmedbjoaufMHCQD3P8cY2kV6U
TaGcwKXAjBKrYn/5PUkh6BHOq4bcGBXHo8v3xaRVXDoOs9R2r1QNEGTVTCnhii4W
BlmJqLVpjdC1mWzGprDWbXGj05JBYMDHejfxrMTmVx2fTvP9vFpLeyA3NLoucvfU
J4o5ikiG2ZySIncsV/ds8Y3VsWafwt12uCUJ8/fqtfyFRVXmHBSjD0a7qXfYCPkz
DkqfUyMCVArVJ2a8wC3mGAJ1ExwEmdghQEqpsQyE8VOimrjTIVL5oOmlPFcsqL+H
JUpjUtssi51b7I8mlrV4fR+aubK2M/UwmVaOCtKzi9YPI7Ha49Skro0RbgBGJFf+
EtR/78+tGWr0znhLDJaTtxhqwoydq0IsMkT1iwOT8tGIlKk56OSwvdo1/e2I66yf
I9Ymw4Cw65nGrSY2PxQeGxV4RypgcVelzzEn+35GJgLnne1Se8zzxuR1GC3dRdo+
5kwJUfgKYIEZcqyCcJFSJa8pdZC3qeA5vuKR2zy6ov7CXfqF0kNylEIQ7D3eo8+S
H/LiKALmCwKfKHBrcmw+NeQv5KdRU4Gzxr2QBBTw0g5zXjscGFCu+oeRVLdDfQEB
rXFAtYb8krTtXDVUi+H4zTj6JO1b2Uc6JjtjHpfovfD6ryKlK2XLlBgbrc1xPHcr
bdChSrKZ6d45SLDm/Upl+VSTEbz1gQ++qiyrGnCGFnLF0NbkRN4Umejevid3qQGC
A+NiCAOHmWrO+whzgBgj9pC3bpKbUsE5wSc+9J4FaPwLUYBPpnWaSKaXWHrkb3yk
asFXakBaBC+aJmCha8MJyNW8NzmaOME8TPEMdSf5gdiYETLIeiF/m8sWJgtJuZm0
wxnYOblgCRInQVvnbjFjsuU0f9MGIf9wOGjZZg0ZWP+XBhwlUzs2m2+Im1bcJLfe
MTVK2IDNYeAdItaqfVKfIpTcSpGmpwh8F800/BlW5YzRfC3Wlrd6iRYuJy837ySU
L+XmKgF//xddZuEQAYWochMCb10H+g/3noY1oja7yyEFG2+9gTK8LjVibPqrGEz/
G82Kacu1wZcPxBx9e4feSuSKDJ3vev1sKhWOwnxhocsl2WPpZsUB+X3VrjNeMwHt
seUJoVIFbffoSO7AfQPmnNjPeeL6aPDfQdP+1AO7IQsORGPcrayRh7XHRa1GQLsM
EQ+JPlIOtpjbV9oeoHDrF5cPjtrP2RmTsjUBBSgxHOKzCaUUlgR2epm4rVsc973C
B9SvX+CzOFVUJdXGyi7KBuh1tnnvzbT75ASCag2snvKXyEut37xHQp0scePXVXjR
JX6HQciSz93W+7jGY8k01fYjKCbzY4hfR4SlP0Et4O3pUxIPI0l9q+PZ0Y4/0IuK
18hfLBnAivwWPQdIqQpNCfDY8GQGfnsdwyfhjQaVClft+TzjKSOPoH0Ed7LGAz9w
xtRHGJCpOVHkq0GKeis9nAthxr/YI6OFku3ryYBcGUUodr+Uef1xbOBY7zFPskky
AwUUqFnF9b3S0FMmwAbtSgEu1/zu+HBYV73TjNspNQNux9Yr3n40Mzi8P4n5pLhJ
ondcn+uJD19hXb/xuLO4zxH8+xwHBbVqihMGEaOHHUSP8BzhBumQ96IjJQ1YE2lC
U7NdYMXVfRVtyCWJbzwvyFALyDGXKXNHHAlqYRY5ZTXsBCYeL5DnMWK0sc6qvgk3
8bLVGq6zQ17iImyBmjOyZGUaL0Cj+O+dMk110Ym40+VBRFte53PzyqWsEQyC/N+D
3SnTg0Tgthhy78UzYZdSArbaiiVw8Vwe+2cOt8QUTnfcTw5zD+TqPqzFpSmyOjs9
LNl03n7T+/uuojubrL2pC7jb8dJO5/nyQk5baW+mUPxXhh9DOVctYhKvLc/suQJX
DucMX9DgjxjjirFlold3B8mVQb5bq5BgXfy6MoE/zj+GeqKpqJggM6csoyNoIlyx
CPEC9fyPsd9ayE/uXqo36NL9v+bSvXUnGG+LQfeJoh4te+QTniKDczASUb80FtFs
mhur6yxkSOdmmumBF2ayM/5TjtzBmR7py7LFS7GGc2i+xZGgGsjp00LtrBji+J4E
Qk3/qwdLHSg6nJSt9twUvLYR+SFsgLYWqWEPLP7QrOQwSIP7ZxTYBcmogRsnky1Z
Vi7tkKLpsf3aOYz4zWFzoW6E/uTJ1pPaikj07Nd01DTjky9Hlhv3f5mzbtZUu7h6
SCBGpTOpKOCyADj+28cPXQYizzxt/QZlqexno45PwYJDkv8q0nBqfFFx02Fn+ZZW
ebLwSEOASWYtkyKqEX6jus2cTrRy5vUPlRyUJRiUA2gC95Q+Lo+fo0akxIxuxfLs
jaMd6NHemC20aHrNTs6cCGJ5A9FKgUIcedFwMjY4iWiB0vhQT+gOLuYrZC4p9bv8
rY+kqwnLoMW9ioslEL0CjBMGAr1WK6keM05N0ft+Ji2KeIP46YsDXiGsPbhqFzs1
kkMpyDBICW4qeadbF9V84TK6kvJUhygdVJwov45WtVmTUZafMQx7jnT+FXDoaw9v
aPkRSn+QsECUOj7vqHhlkdrdaFA4S6rVCcLkLN0z0rDimXCcl3fTXMSP/Gh4luG5
EuU6sKUJ6jukKgTrhcXNXvTw4nAY/6T2RnkqpwXqUJmiryxMX1bBQfBGasBwS/dK
9bFkb5lPWeOpDkxJKPRiRcE4HGNFFOaoeZoJX0KtNyHYm2wsVThENFCE+dL5CWaH
fzrZv+UcNML2HCBVCr5RkNtKHaS4gYbW3oShSZMOlIpH/HIcyTDcm4XliwD5BGda
FWdoPn0qIqmXZ1gNWRXzfGMwYdevAqgeG7Kri5MQPH+4FAEEWSXhRbvW9ERDbZ1u
iJikdBhA+0SzkBLrWyct644o/d9gxl4zcl+XRwaO31zfEflo+fSRTA63X2wGaJYv
xHghOZn+l2o1lPCKUf7qRTEOZvr6VBGo4xecECFE7CSHbyTffVEoM1OgD6Z6daKN
HimxZPKP+fuzFkYjVfw10k6xFoXxXuEons6jsNaARhDug6yK7+Zw7QlW44Ejtraa
mNuhyRq54QXhqijZMy9kEvYnVzIieYje9yDvvswS+wUxQIEqiwVuHrKOlAWlQ3hr
Q0mHjRDtqkJjrvjDpExE4eGKN3k/E9vQAuBOEGXL5j6R//yGWhon+cruGF3vRZsS
naAujyZWbaM5K3ne0JCBWQi/kVsQcL0/9zch70JRFAI4cZpICJAcbYbHOgm8RRO3
R9L5Vef6p1bhitbexgdKixI7w4hVvHoK4MLarVaDrAsK4nHUMyjtYa8iaymBc2NQ
WtDiFeTLBfh+ISNX7Y6CgxmJOLEZ0of9f8RMCkiRotQ0M1EWqDOcA/Hg6bw94L6j
LLem7Yy4rxGrPgimJGk9gWSvwqaDtXEu5dvUH57Wjsv+zIEdnqiIjDxLBJ9YLA99
Pi3JZjA/hgWBgdDHWIAaHqIbuStnkpHpHzmWMZYRrGkQvLVze42Y06J38k/ki4Sq
wEWNuINRro9FGhJXAZmolhh7Q3anDFqR9kB+HsbhYKiRBZ8o0VFJh1I7xof3n7hq
1zafbtCFK2LzFz+cgtJOJdfB8X7xcIsK8txumD8/5tUrMN0Iu5EQG+3FvAIEJHNy
RPkcul3xNceKl+SzDTInlW8btFGzIMeJOjNk/IsNbMuQEtr93Gk9KW5wMSlIGhUX
7qhuaiq8AJrToGL4q+dimWqQWVONcwdtDkcO8ehQz4bfbYkYFnmPPLGDS0BBr62o
1FT6j1gq+BMVPVwQ4cMYr7i+lSXdGkzgc+xGUGg6PG2Tc8NtrS46lw8FjVlEjdNF
oJ9U7Fg8k98A9MVwUwgIcTtsKqTVpEEZkDKVS+On+re3wNej2NzmrjEsKS43aOGV
lEiq0gVgzphp7qFkU8ZmBE8fZNXE8z0NCIn+nzWX1L/YlAWRpvmFjPvtDtPDNe/m
Wq7LRA85WAvvoX+U6v+0roBfcUb3vfJmuGqCuFD9g6Xp2qUy0ddk92p1pHn9SM6J
cPYoPF8fI+IOVEPqYWvLiwgoj7M0r8vEG/dDh4QdV3waoRmR0ksLCgs66/C6KrVQ
pPEStlgwblfII8xC4QXvVnRyhMqdvIEg5vnzdgYgAeBpzXpuxaZPxjp7QgLvGyX3
j8Azo7eJFvZRWyJh9crHvX0WnrW0n/2/nLkUTDRTDqp4HbAQJ/11pz7YOGPcoksY
APhw8kiJShGuuGRZq0E6wIKVHqDic1ZsNhskCB5KR8qRQs98HapyObEAEdejWM1f
hhA9Y2qqMGuwmrVrtKgczgMeWcT90UONz+6rNnuR0vYu7WIbumNDO1fqVZu/SH9G
gqv6dV22s9M9DkozzGIS1lms9nSSoBvvn7uLSkSxopjRqFBgVFvlg9pu1mbannv0
37ECe2lByQVrhMQr5C/OUKbCQjcoCX34PaIfOGrt1uupXHsEZRKJDKgNfJEWOZO/
qzF5Cl/FXQQKwjfZKzxsL+Z8A6XwwZxlwSJnqvEEva3nQ86rt7nlasAyted0vpgp
A8FeNz55IrrK4Fj/j26kRfGLTg1pgPtbnQU9gIA728c8WzMp4ZF+wk3y6n01XFMx
3uiG66iBcFnQ0SF85N5RBmcCpIWUgAv+2pr/z347v5Z1Uf761arpG0aeKU4yv0pE
Chzeum5mqNEUS8DiPIHJ55AtZR5T3b84EgJ4W5m2MD+/iwv81tQFGgkWaEP3Y/8O
3f+IRR65EG7oVmMSP9d10W41BYkCf3FpYlPgdiLc+RJxaPeU9q8YG4Rv+/FMqieA
UMoAXgnNg344Si6YYB0Y4DBP/oxoWilGXgnhsL7GYpOi7XzGPpBo4GbrWwSjlu79
jKAVndOKAC07r265nh5OlEjk/bWIHXlSbwZq4MDoLQd2F7VCWQA4y8LqAlR57oKn
o1BPbGJm5umRNupsxD+AALVWmXgfTXqFr2rbhvUfNyAquIYRcOAfugrt+w8RkZVb
1ESks4Ly8xirsxvvyK9oiEsV4n01yVtHneT6v9XroJENlrch2oXeHZFBUNnYDFI/
x39uPZ6f/ZD5MZPqnhcfnUMpL4WEZHHTdWfOWrHwEUM2BfNhtE6Xvb34QNyFVXAu
pT00ooiR9esRWHfrpCtHZcvc6hGj5KKyYmob4Ihc0UvskfW3jlGhZNP2MQ0GyLxe
9sjvxXvUbAuA5hg44l74l3u1c/xGT07/AAqL3xRfy5EyjyWEfkjZK23Pp99GZ4Bb
8u0TNWFnoy3yv37g7n5Ep3ytJmxkJYQkOEtGpTRGxwHs9SLfNOibkG6qyJZYo42B
MgqgOv8koc0ejidlUIgcJ9J2uAUHjTeTeuu0IKb8BBJvydE3HorW6u5PN+7LlrFV
rRERgj1fHR80fN2z/4k3Jw/MoqC+RO+a4CoP4nvpLoT/LaYUf5h08ukDm+Sr05rn
l+v7q/6hYFVcsFUEY0+qwFpWUQox/395XqXUPueNemhEtPgi4E8TlHuR+0GKY+I4
kdLD0+aECLv0BLy7wJ5W08LHXZgnRQts8w/mDX4Cmznaw7Zv8GMQqaML8Uks9z/b
2gxrRfkAZs5NZVEReCVjp/sitZb15OKNkHOk9ZrpWcFU5SdZW8MYcGR/zZV1u+6F
zlJDYpn+MpRGH+XHMHkPo0htxHxBa+Z/cWfExThKYqVf2Z8zGXIyTyTr1DFhY5te
eDMTUTS4+uAacPhAAuY9OpktIguagg6DheVDVhjSE7adJK3GJ/1YrVSxR4A9OBcS
5HN3WQipLJWM6vaoKpwxiyEh3B6Hvn+DZvV/V27iunAdpcEuRuG3b5VDmeVdecq2
x1LqoT5swgT+TqFMexqGsOQz6P3/MLbUdnaMpgle1uNKTwxB3R/LBoj3CZf+Ia6d
/C2JDnBe89vo/RNf8k1nv5PBrVcy3sUjtbG0PMt8IgNyQ9iQOA9A6wbwPcCEeNlf
B4q7GWmGi5jYuiPRGYA/3MBaEe0Cekfh9H7JUm/OM6LBitgvtMIsmprWKpaLAp3i
2vN9sQgNLfNIi8htfn2jjCGF8d8B2jZe1cevkhBtx5+WeAcYKnCbykBdMsrLfUWd
q3iVWtqguthuH5SMT+fEp04TQ97rFe5IoYbbtZ7K4JOUYX/9U43PM9WjLd+l2KoV
jPXm9ntQ3r1YQy1oIn0OtFisfohlsCzza2FzSf6fMW6UAjtOC618PsqQPgh/3/UZ
WD3wTX1cZ2luYR/S654+Ssk6PusFARaKWX+PXVs6yQW6E4BuLDi9ntZ6eLHBwiOS
Rt00sCDINpkHElaONkj/MLM0F1GUlbKxKCU/5ed+KcdQL/hXe3raZ4fkI91cXZZt
XVrKHByCv2V0yKCzhBUc6idOSA0G+QSTX8TE32DgaPca2rXHe7h1LRurgzbmBTaN
B6D5XezeigNRyXs1vKn8kxxEsr/uzeKC+Ug2K7YJxit0TBH0MGQibnan47DmVwty
0g+SKtydqsktgRcgao3wzTRQXW9XBQZcsKu5YwZ4x/Xr8AF7BAUw1BooVXRZs93U
YZBUcroRKhjqZoWi5WbfB3dYjh+2Ng6kFhvtNkQWhAvI7Q3Og9p5Mm0yls5pJpXd
H91nDZy3I/63D6Wr/GTLFsO+rqwCZ60TvFAZfintkdvyG4O9Hjg2CMqiF5T4tEab
vp+ZpWk7rV4h+WDUVkITsvFStt+Q13404xv6qOdnjoKRrhgIqLCXs6mw8Ep6es1N
cafhZPktqeLXe4m1G3tNBj4pPWV/V+UjU65gzL2umYfBRtmFFCbON7+JwPfq6HUT
04Im10K5xqVjIlrwuTLI15N1/2u0iyau5i6a5ooXlJerlEiyVIkKfL3ZQ2iFio+a
FMbjUXVk4xWR/oCRY8iNTzDrFpza00m3echE6ssUTeQeCGwTYrILsUO1zZwcuHH2
3gd9C0L4DMUQcUdxB5Rp3UQv5IBw3uEn3ZSBImEHwczyBZWgYegMCqMwtRdHq+xU
0LiNvexRnPZB0jyuuk27lWIWk67Q0ndAQmVM8gHG7oOFOAGQD7BUhLUluo0BEQKd
ckNnlT2QmSyiMfZwPaRzIS9cx3N2s6p+/fdRIojrbswXBtF1gzeSHcjZ87kxCwVy
K0o/S2G7TvcIPCy2V+MHJEkWntwOykul575SlVDQpnYPD3Js8LPY+GTnvgF75bW6
i4CdR9savvmkzuz6Cf8bisHYCAedsJN3eNiqrFGiekypiVJJo0EzOlu14rlKQMOf
MZOTOr/mJJvVsN4lSoqOCOo5qfGi7oN9XZHlyjKhQkEznBXO6H9Vo9W4LQGDbNMt
kBnELrTD249qhXKF7uNhbWZgXOcCUqwvuimyfQe+wcKw0Pa1qx3TwrCNNMYMSKMd
o5IfT1dWYmc+1G6ocdX7d1PvviYSaaB3VUBp9TmS3p52nhSvAIZlzzo2w11+sJsz
9IdhLKayl4bDzZqURYcYzx+T8eEIwYMWfmJCZt/5yLVN3CDigBJ5lIJlDMHweE8Y
qtjRiZozpAq+ghURGNnaXR8yXFhT5agVt4/SC3JggJRs1kxUKwBKEpHMevnURVXt
zUCRyUr2wUcgHws7P0uh6tJpTMVJZYLzHTqKaGVd6kVbsLF2EECSJE9tqvzEjwxH
aIlDZhfmJKc7gcZpa+LXJM4NClgeEkmdi0qm1pVSv9yW/TCudisdybADfUOFZ0Iy
vjy9JgjajAjdV1C5mnKwzLP+Kar/32M3l8jkJOQzTOg1urs2pLcZsjg1sHO911Fm
IEgrMo3+ZfOXcOhAxuS0LbbSyQxQNbWcDhXFe1Z+0bH3hr1n3+e6wA7n+r1cVWiV
87A6ofBEFn/kDmRNyr6WvVk3rrslcXc1eIzqTMPB1WNKPADnRRe3JVydMjqwRoWG
D/9NpR3DamnDHHZu5sfX9Vex9wIFPwwnpfcIswtae8sOylsSNjHncL1rivOk8aAh
YvfxbgEACQVAcFSM+cDOqD/4Co9YDwamJhAyZTGZxrzyCTSs/9v4FAhRpWbTJxzo
c6QlitND2ToeCwmAB8ag9b2h+iZYxXBukM6p/v5R0ZIfOtQw00MIT552V1QWCIvG
+bYEeqtmqtQXDgNJjGTvMC2zKNEW40RFF3BraHlK8ZWKI6zk21rhneSg1VmtJUhL
06ko6BhtwlVSovf/kXW4ehkYtWJdgisNW0Yby5Jc+A9oxe2AaI9VXhxVZgSGEmgA
UnFfVLwC1VdIrccqfipk3MQgu/xcCOxiYKTIqyfp6D8+Ps8A9ZXxzlGh49zf/nUz
oVklzUBVPNjNGlm4zrwnag3wSQg6Qvy5of7XySomJZoi2AREi9Pe3ficfUUmfjc0
m6LCMCjF5ghw0jbF0cdpOYORJZk2UORayLsM2VWiQrhasvvj8Wc/r0a61xqCx69g
3ALMjjvKOuyFizfq1Vh4TJlq/Orpn+DZMIg9hcvh2ywRN/fHY66c+vil7PNsL48z
aO6/O9N5ZVURENv9wg4k3zdpOGHRfAuKJNUZF1CY8zgIz5QPcC/XMm8VmaD1ZkMo
yiggbdNDajJKcf6np2BnClvjSKIMlpPtJrE+zilRQ9mx346rfSc5mPmbE3XcSRAQ
LS3AuT9nqU0Vzb5s0deFvKYQKhAwJyemiX9sOkiIiJg1eUkpTFCufIPpAu3eAZKE
dxyWO9sFh2ESLrHWCGU7tGC6y9cL9YRvKq3dz42GDA89zDFtxafQ2DpQoWq6EqfQ
Bx1IvzEQgvZ1/h/3Zg4FYwoRZnFMfhb27GLNAntpwYo7hA8IyuRBZvbj7NQp2G+6
IVmq9N0uCIFVeDTHNmVp76M26xcawBtD9KHPr8DlLzPAULNoqGQ/SAtF+CAtaJJd
iWvtQ/j00WrDkOBDpITFgNFBd/UkMpDQxTuxY/3mP01jzPEV+cfWoUoyuGhfDECe
zm3J55hrHg0JdVMoiRyL9FSkaV6nQFPVYS1rBxLf23U8x1HCnzgHYv9CFq3JiF/O
4SZuBvck6MDfOAof1g4B92XmM9bZrCMdcKU5Bt0p/8qkaBHO8golC45CPHOnZLuL
9fpM9Ipdu0vZox9wOjozVFw22GzLO33KUV8fOIB0O6br5XXyGexyXgEp2qChLJDM
ycQh0qkeIIa6jT8qo2I/1EMYhJWPHePP53iTtGW7mDNbub2deMWuxCqr7OKU1W61
SUS+qkOHD8pxT5Bc7eW1VdCpmC0emJSAk3IFtB1PWIlNz8qu2rnjsBW70kR2A10S
P5tC6xTeot/uYah+yYRCMl0ji3l26Pwc0nGpjwB3XD/WJ5ckiZ9TpwQD7R4vGPAa
1pLQ6a/OydnoFfTl9N7jXBXUf/VuzhmonBitNZsry6JrgYthqCj5i+gBTqIBRpn1
sIPZJKlXRDXxlfXb3jVrqkJCzE9CiHodl6TQi3wsy0WihGhsVrbwZEvD8pY34vPG
gtRKIpVjsIEzwXSQ8T9MKK+kS8hFanbZm1vQlPaCyJJn7r5rE2fPhJ4m7xzSWzcg
I6I3LmworAbTwkHFe2AnmCAZhZ+CcmMNHCzP5/X19tgRjQxM1vnYDBviTChAAAtF
JYqVeRzr1OmDhgRnXxVKF+dtPNqAi3C8K77B+KKMVeje5S6iKT/Nw4wZlnVzb3X4
yHwRqc5aBvmXRQNJBrBspu8gP0+Gj8c94Ea1PTNJHfuf5XnXMfpIDY46d5URXdOe
VLWgKcrQAJCD23E2bs10BjMd0ArU3/LQ7WDrf09kuHBy/bPDLLcElNv9OJgttCfh
Di16HvgQkf+z8UmEdg1SNfCIqUTOuMuGqsb3nWf6U8GQ+oGPSNSRbi7q3DveTbCU
t2WLBqrlMtQXUIh3wUfUberbhbCiRfiouC1G37Qe7YLXqc9ZsRPOI0avBoExW3t/
lRKrrbthGeBfFsXiTV3XR3TFnZ4q5aWcSbhFGbbYBMkMYdj1gWFNDtLA9qyXNVb8
3hy1VGlAC8BH1wCBc3LuVyCjgXCSdO2fcDL8ZFOctYiGZ+VKMbBacd6vZC5pswa/
Ooq7dsxjIe3PvtXyIF9+tM4WZe22gDh+XLT9RafDBxKbHmOHTwyVcqdtJFQqmSi+
0ruE+Zv4lhfJJ+qtJcna4GL9oPOBQ/pQhLQpCButWthqFjv3K3qxs2LFiK8KwCt0
lfaQiQDgo0w736kXJDO3mYbcYpf1BysmCHoVp0FmGgYv5eEqh6o5m7tm+ouZ8MRs
XpxKnL9xMRXgLuvSTd0l0FMU7Kq7cyjEUtjXguxYgzVUIRTK4u880TJa2y/JW5FY
pjr7Dd4yg5uz3H0zDjMnQ4fzu9lSULmJ9Jwwdtl6xPSsixm0VO3zehTAhFOG7BAs
mTE9nroG+HSG/fG8RkYPxVoiE30Rs+KoObOghLx/zZejR9GzO2soqx9WN5j+mUcd
33wtD4VsoznoN26jSAG1jD1u8+ZASXCns7BSy0tMWgs5i0xPjBuVY/Gx1vuslFi6
E2+W1IdUKkv/mGT556jTepX/x1E3+ZaUO5XE6gqaZ5lN6AESKxhC2uGkNklDZRSp
BxFTLM8Y7hSAfsd93yhWx4HJBCI72K3hpQ7oupvrs0n79kyqmE9nPCx/qXGtl0RC
Bx5lrukfcz39+kjHSq9vMlEsptNGlbHaOTa9Za4Pqy8WBa7aEd5CBlPY4UcofHyP
+eSxWID1YOPb6NuJdFzOwBTew0RVD8tr5YdlkOJGlPT16aKc5ND6+6O67Hb99S0V
aNEUpbAjUy74lb+qto2lglRdddd41BZ356AGpxYFJ0uKgHEK5Gov4RPUtHWyfSuR
RgnY0m4NaLSSHX33ZYouKd5eJw6o6151kvlzZKfBXXN8azkXmHriPCAiVeQ07BcN
DNGKi2rIGwzSMY3FwKG/SxYyeVYw/Q+eIijKBbSvNp2VxmI4mjeAdn3svrSoDlMF
aB9bYIi4pBZdPgkeKrgD6f+7WCbz7VewQnbVo9XVzPt7s0hL6MRnmke0DkBlpkKw
nI9lZkwOHd6XScZoJuYIzu8xbesmtHwnbg6zqA/LHmpgZSnl4M+TDVxAQDiLgGiT
BzjYziRse9fZsKKfsJMyuzUzZojYm7uvOC5jV6RzyWdgCKxx1yLazKv38gQfntVM
KQ7xz/QuaNSYYNEGi1IIJ8qbhKAdOG9DbLRW8doLcTPKEKMCNHPDQHFgsQ9MS/E+
MLwpdRp9QVCuCks9KOrltghDbM+1BWIcgHYXW8XTngg+1/ff4glRwzj1idrZDwqB
Sl7vU1wbK8GchyjnOruqSrwLNDubx3HBvztsKLMwOIZPPnq82zzU2+iznUlcTEHX
Qqgx0kHkrq1IHjvQjvEC+V/AnQlfHpK3z9WeTuep6BCn195rnJuyh42ueT0x+oE8
UjTJuGnpO6X5musanbYMmK5wMNN+TuIWGZubxg1goxqF/obnGkQHS8pwclK9PtkD
vtyAiJvEIxC1bVOQlnK1R4ZtRlTWPYou6TR7rV2b4hMNYDSXH3NDbyA6oJMyf47W
xGdxt2Qr27Gv828Ft0jLu83x4COCzL8lCRguHNSHSuJECnS2bG7uBPiV5wmWz7Q8
/1jpYPkYMfwBVuo2zybGIhKW4gS9FdYIl9T+Sr/kDuEZaLf5nklB/oo2CRSq0gjO
e9aM06484FSny/avByUi3vOoVXOCUwN+LpJpcUSmMVebDwQ7D4X/qUufeKiLglaq
llXLBALQESghOo+t2FyOWgZgDuYe2w7JN08m8hUcxJZ2DUwrCFaxe4Cs1ntFoVSu
qffQwv9UaBO6XUHcHPDwuaHgfqkZkmNjnijzr2iBG0q8KFHAqqRQ6c428QPPDuQ5
F3mqvOluwEgIdim6ccW7y+UYJALmjtrMbByF9VWL+113fUhevw8/iY4DQT62Wbqc
sYzlnOx9tpOoL728t/qfIcGUUFD3lkSqtyPpVTP8SUaepzkDKIID0pMp1RYaIWE5
im7ZuT1a6al6swDCpJlecvUap41qLH0P26c2APlmxXGnZLiZsWNM6g5gdp9Gbn5B
v0vkAzTlRoKmiiG0Xde7+zmklassahXxwnoE9fAU1ZoM5Hgm/Rj6oyv8Ph+T/u1d
5tnvfZTfxZtVvihNZwFMPmA5Qup1k5qxX7DzaB3Fhyz5HZX9cBGG8BRACDcUAotY
LO67LfRuOYWHXEbHP66bLF8GebGLL5sjjXh0xbDeQ/0XTXvftUB1vXEUa3kjwEXu
3gaxSglu0MCZQWzntC9YK28ddmpnszH7iuE1/nVnhARfpqbTYmpnZd/+ZHrL62Gb
ebAZ/pRAJaQTmsP2j/QfcD6M5aNNkjGTuWv7F006Y/ebbiDDM989ES5/XU3Nc3DG
WUmTdgQu8mVCjAuljliLkS93vgs/KQP0MJk2lsz5qUFUE0AIvUa/CK/VQzkNqjdQ
YLB5Ha1IOiHbGwVIl3L+epZEEO24J9jIhGLlm5VCIBAM7+VrMZDyXe2JDy4S3NvE
AVPbOgeNgxo7QDc7ZhsMroVXCpx/iKoYV81ii505lfbarvtQYB5DEQIkq3MUU5bg
FLBG2Elw5t/PrTPM/7QgyA1zOOEeP5GYPsEOCJqzdICUacaoBuAKkFNoo919oc2M
8+5viiHNGkbLXF4+x5RE5NxPOKghsZV38t+40QFwxiQvUmquK4jya6+mp2UH1JQi
3tEV7LDlQ0lUeDQ5ExV3Q1gzk896vqQPOTKVp8Tjs8HQYRa+C+NqUCtr6TXl8Ycw
XBxu4JfpZQm9TdSJDVaMCiYVNI1DG34l73qs8dX0Opl5+GkSYxbOzrVcGLcA/vx/
Q2UwsUP5rVOvIsfgUi7z4PUEU5RHD1AaRBxtV8qKdgJb1WXNASryudbFlSXPgRlA
hr8vY3Igw9w5lcZZ+c9iGOLAXJiuWEtv8sQe8T5N36yAQ0GzjwgKwXzVrm4sH+Hb
P+eTeoW/TrzeLUkTtDlVYT2TVLJT0rZaWQo3E3uvFnqc+PW9h1c2gSVVTUhHV/+i
qv77/PApTVUpQQjw5wFI5uQhW08m3nEzfiuAJPlGVmrw6oJbt2L1ZtbST7/gcJ7U
L5Vj6iNwNT1lhPj/CjFjxYsGpGhAGEY6OKgLZA7ag27y4YLBccoiR2CbE/MZXXHp
pg6JqeGnyUuwP9RzaAffHnEIE81qts5P65Fgb9luwEVjYsg+tNcthAn1jQnASey1
onZjP9NwdXdt8k57a9fTQsdLSRcTa86+cLp/UlrorGny7c2wirAJdm5yUS3jTEdd
VVPukZgHFkxE7nn3+m+tg04tnEwrBbmohMBKHjLxvEVAtGEsiEJl0EvBZ6YvYTNs
Murz5qVU3vypq+fbScphSYrbLfNn1c3IMd2a7QX7FloorrZsl5+6thtVjbnAqt2X
/pAtJnUoSputEDt/hnfJMnGCl0uQ9oXBIuxDVOJkGHgLQwMJ9i7cWU5jdanT9oAM
uSd160J/Q98s3wT4WdXOifURRYbw0NxyJurJgyxOScw1h+vnCTb7qGvEPmYR27yR
PX43nO3A/VTkrhp5iImm5N6YF6WskmD3JIDwSnEEuYBkBLqXXbK4kcubmUnYHtN0
66xmfgko9xQtFWkf7jFyva9HEYpWcqvJb/bH1mtV2aNCE6kxu/k8d4mH0kw28Zyp
EQd7QnjhMv8qmAntSsC51DHSb+FfSQzsb6DZGnY3bumRY6yQsKVcDu/JvdG81ZY4
vUSAas83wuUYpfEUVlo2LrdhqyapLvEOiXi2cX62okyVRWST9VxrUIeMXp/UY72B
D+mKnCZ4XATGegnXaez1fnG+ZgORs6hClRGlPPpqSVFfea69gMDZjQa7d2fEmtzf
cr2oWx+At7YNbNxVQCAVIC+N93oJJ+uP1FD8zfS0H1iODGI2We28LOAD/9RPZaLr
LKuzszo2Lt1/g4ONbj2oHbCQNetXPLrKplkRi05vtDMQN5l0+qd9JyDY8H8yWera
cFhIcVD7bOSzITw003dSf9RekEEq5VKdkr9UXoYuzEzJ0PoFimAiOEtbqvraiw9H
OpUqA+zDkjLV6zda7frZkoboAwACMzAgwZ9pCgo+cPnbjaF2MZfT5IlGh7SOJ16S
0F6Q8iPWqFguzWbLE/iMvC9UludObQKY722rf3DU63xmemaUH5MRHzmXPgEDcrmA
qS4sXgOU/zZGtEOJXntqSJOGAzakWZCi269bDFroqzLEPWDSW6T2TegzoqkoVQZa
kNt97ics/U9mQaicuXJBzZfy3zwTvRYVBqUHf9sKnRjWc6a4TG7HkU/Ad4V75/+O
a5saXPXVs3yoS+3tzSdho6Uuaz5HPintXf5MzqVpNQ+GIdd1GWzlqwHKb3aXZOWe
xVNxRTHEXbOIFIFx9DkJfB2QyklWmLy5TPu8KI6dIOw49xrFE9xIcZozJ86Zxdu4
niYeHEodlsHgzdMlwoSvpozfGEK8ddFQxgxZQ1PFOkGRVNRDdWpydAP+zDcGFXR9
wcdAhYQd30sUcuhNDPBSXXMDHswM7EjUce9OpaPe4AqsTtErZVngiujSbJtk07Uu
1XYZf+El4FbNUMHMEnbPkH2ScC+GC0mVtGIXQMSPipLzgDYJmo41YIJRNgHu6kJq
5PUEAen6lr1yJhY5zNKCFU4U1I8+u51ViWqmlSIwM9Y5qoPaJD+vmegsw0pxikNK
ymAhTzi1QqaQn2SRWuPm5x18EUDQH9gVaFNN2yNWwICi4gb/KP176ZTgwD0NUF5N
rsXBo7s0MsKRu7xz3pkM0J/FiyaEY6cOqZXPnlt6y9HDq8292N/WPbT5jKq6ej3D
CJz1q5Q4/59CZfm2htlqQR+1A5CRg4CMz/oRslJV9pIwpGMSTuasVQk4SXa6aRad
mwUfbNVykZNnUhIbIKsVCiMsinxc4niR32ora++fs1T9nbdAWpGsGzE4yFzcHaqV
lvZFvpVX1kHzIO8YeUXv9PCqs34pYP8pe2UobeH8fvFxFLL3OgOyx7RG8WTwnpvC
TSTt7ouplKsIJhTJFNakZfP7U0L4GtxjVF8SDmmeCa663GBWIe4lXGUzEKRipCbk
WKprprxzNU5U1frfxUT0G4GN9BAeQuAYM21VX389gUkLBcr/sfzKKK9VBjvNvEzB
tY+Ky8kvnfy5gYRVoSvttscgLBJcwucImpi5yDvhSXy5eWBowAgZ4M0LwOgWSFL/
xKoJ0mpHYNmAU70PsYbYRqzLo0KEHKEDeJgdtCfLxvTwj7yoBewJHqedmHzOYQEW
ZEp26gw23uFsCVWkdT7XV0mzvjD0j+hVgGlFO377WVlTZbQCYATBX/E0Bz1+j5Il
O6a6oJy8ZbVYsmcxhA5Qr1DWG70qfqMFG02Te0CeOVYBfhgh1arn+Q7bENi5gGRj
afRga5zOzv2nIf3w3TusxH5neStZBBU2SI2rtwRDMt6q6ZEcFkN1eCC6hcKYkFpY
MBY2BLvJaCjImF0i3XVtXKgkqcWdJPybXyoR2Rq3SRR+0Vkwcq/ax20UlZ4/NRGx
Ndl4w7EnksgX4FluHCXW6XLICZmybJGrQSNvPk9LZHm1qLL8yKFCbkKtAq+j4leW
iH0bHJNQzuWQCfyjItjnyP/R+Ja13GSH9MjPzBurGUGViRWZ5kcb4XN5VdNeVtLk
OQWl3o9+dxqmAjcLx26ZQ4YcFzVtuYZ0Fk2szHzias7EyZbiiFfGDlkJRpRR5c9u
WD3FQNZPe5V9u+5av4JO8cs+AXQj8dqhW/AaZ6IODM2Mbdzhoz9CncAPFM1Q0m+w
g8guQarvHA9aLp0vHM6jJYb5eke/BaFKAgBpJQGETvSqLG2YinjKZFmDMeGokgmU
bjZo+7CUoGUrvzstTGAnDJk7P8bznBalWzfX5TA2AS3TtymBxHXJt5g8shLnxI2x
TIvsqH1G2d7rsvQdRoAKAWMq1y40g1DOtv4sqqC0wayIm7jVBP9qBdz1gKf2OWfk
rHoIDscCac/CuDUGhzjBiMX2QhkCeUI3Db+axNOxIC1bE8hO/tSuNPf8qODsAjwi
hD4Uq6XZeNFLmot+M9n+6NePuXZ5R68wsdcrO5ZCVdTjtAW/e5e229HnEC18SFdC
Vksyz45qqzehBVq0uLdcTvyliKEhLNSy0zTbCp76xWJHWA3qfBaHgWmiv3sTPeDE
rPe9Ci0ZlB/0zEkCba0UP62R73lr9obcQyongGYhB+IYWV34BQjnrnvL1oCFlu68
cqddtutthkRNVrusdgG7gPkJ1naVsW6NBSPTcEZf3FsO3Sun4w+zmQcDgjl5SC6i
2BRt35ePEfYy0KzR4fkSZh71tx9cwaukRNGb+T2DXcwoDQP9Wo09FMWDFEnc3Rrj
KFJtYsU9s8qdeS5BkbHJIpP0MlU4vVosRTefY+tSn/tEzsb7FDeaEBWSgxXmqC7K
i3GgJFXwkjQhKDa0Nul7SEZ5YZlJSHZjbwCXCJ1O4q5N/oFM5FFbNj26iVpThPp1
W2Zemd1pS1MNtkqn8OAAsshu1Olc8e/P/CMw4TrJItu0z0izhaLHeW7U64hQOF0P
3J+3wTlvjHOxCCKdxC93qOx1JCng8huvQj7I7sw8iT+rWO5o0kN6NMfroJiJAoKL
qPDTt2IDtmAKvezpuFxjrCwYBo+pN+FF1nLl8q4ynoCw261pqN6VLkRCkgPjMQvj
KQSQiVXG+8EIZQCjHynGS8k2vzKC+uG+k7jJbXhqnoMU2ppndccDWIL17x3OE8td
IVQOa9dQ5heNk/YF/o6hx6L7NwzAnoxojz8uvQtHFQ5WY42TEru59C7pS+vUXX1C
+H8mpkq/vGGINrB6Xvexq83mk95fcY4Gw3GHkCdD6B7k+gs6sZdufQtKe/poAidV
4ibfxq5SSJ7exxAL5UwnYrZOmSjZOJZRIGui336sngp/pfY9GJvem/fiH2ytKn3E
055EK/nJXg3LVzM52AkajCJq2++sNYbkIP4Eaf02rNsAJW7lpc5+NbNGtmAXB3J3
LMU1Kt+KXAMKN626jFD3hnddEM0pVVzAggPVBWhv2ei9oNyXtb6o4CJCOfp5lpFL
6azQ2dE/wcglKkPyQHkWVzzX+/5FatfmiX3Ot7BldZD0BlsWGpcL9kn6wP5jAagg
3tMltuLYzNJizhMn7elRqyVppzEKv0vAqlBCu15p7YSAvHanC/OTJz6NXMfj5ikg
MLsDd2f2gCLk5/52I6EAmSeANGa/OMEDwW9UjQ03udy7rJ8yMh00LQlY2C0gMl8j
pcd4XMoiz8aEkFhjq49SENey+Fu/qM/Tqh23O7WGWOFdfBZJ+OybJNpFMDeP9CG0
B/VPwM6l8/nWAu8gZAOSMYMtvgorn6+cGazT15dQJYBfKT2LHbxO5Tu0x8yVrJee
HOLC0r6YLcplOcnKgZ7W0CjqP6gvp+I9E6AB7L31+EP/Bcd/xSNBQyzt70CO20fX
WRxWrVzwaRe+kVZtu8GH5ZCCRUzLSA09xw9UAx9ZiO6ngyacjwEwciiQcZSmdnpr
zO1t/hqO7bPrCULCmZ9oIICTocjdaRejbkYldVKvthxYxn4lvuUU2rHXGvh8CZGk
r0lEi23IwFC8vzwqqnJKwg9J3cr9NDt6w0gvPiWhtkJU1iEzG+yzrnlQ2k6jNGpY
WNEdKPRoXipT2yo47IEWSKmPbCvXERR+DNpZrnobVPYKKyb4NO/AcVj9kFouClMu
EAJCiIkrx5rb8XLqWtJ2k4dvcH56ZO8KwvFvtUyMxPv0dzuD54Va/qi/R/257Vv/
Qa8S0f+uSB3BORKeDHtkfdnMHUgrlmFM9fGeY3LbuOTVB8SP95aih+hMGzvKYuyN
syG1bkBBfExSjkaCFeheGskmdh7zAZFilLmYi2gEy769HgdNgoLARq7CUbWK2sDq
tKuOpMRwHYJHOa/+ag0/kN5qv4YsTNzYt1ChaBjuQCTqd9WIpUNasu7dhoRYoN7r
QHNBuvQ8bE8MDpRbOeDiJsd4nsN3QCRmEXsm3AHNpm1Tbh2xce6bSFi9oG2FwfQb
xv0Y+OIFUkwxGlQcNnre72PCxbnDwUksAQvDTypQoEnfCUpmobkyp022shGePHOV
HZKK9T1NZe4mGRRWED7Neo5ymBQi35Cplgu39NNVKi15twX5PC8UDU8Bb4/vI3VQ
sXEgvC32h9tX7Ods4+YRB+Pk5bMosV0pnZbNH8ldyMBc8gUe73Q3lHM/m+v3Uco1
0c72hujs/mGFYadyHNGDNwI59bp/Ol62sk96dazGNnm7mxXiJ5DgHLDy6NjgP+F2
SyhAC2U3FdhXEF1MzzwOYJisZNX+I0gYXgwDDnr/Z5aX/9TtTBMArlRaleve3xYD
PiKkY9GznaGXz80P8OKC8g1BkeyA9XdASIXyrfU3QuToNBvpKAr7spGE+QSShq6f
lqRBVIGaMofy+yvD3nEjeK5eHLJ8gBmvH56JTnDHSBEGTzf5QXnG+/zPORF1cGjX
J5pyA4fx98JZgd+mDAtj85K5jbRx53wY/szcCtyEs9SMnMVzUCnqB/1Z+E57I8tA
e1li36mzshSeE3z0l6MuR/wx/dR68tE+X5ErWLuw3tTZPiShDAigkZMG/PT/Dfjd
ArDvPxnLGc5msxnQZElo2mEyfn2W+e4DCEpwH2x+QqbJZxIlHVfezZd5czRxiX3J
2HUcmEaCEvAcaqeKmDgM9RJOuSjNSyFTN83xPl8betuhMn08JUWSTKWGptDY2l1L
nZFIqBuXLe5H058q0643bGOFhnWLaw11wdbubklYHeuI5XNJ+R0g6Gxp7MP3yGTy
owL+y5zQRlt7l8alJx4Wu0DqewvB6sOzkPxFq23SKlkoZS7I60/zO6D6j1QAaiCE
11pAxpbbvEdRI4fjrEJUCsqQpIbDBm97bla312dN/jHu1ktUa3M65BwAM1VB16I5
T2XeiPQemxoErXOjvOL3HU8rERveoX2HmnKyeiti40CPlTXrEvVBuk9PllCdjf1J
jrHcoBc+N3KuHfORHdgBldiZvq9W7uzZq2vEesJzpBKbfDaK+RcTpK9WweAqIgLH
dTER10UF3PlsgikwwftkBmRg4iUYcRSKHC3JEBn5vKivZgd3I/7Js7G8/WtNdIyn
k+ALZDiLDUjGi6x21BPQZEAT4Fc8dOVk6YSHxXSh2JJ5IROzlG74T6NBdTZpq2ts
x3wmonHMP6vVOEAaGb8IJ90pMT0hiSj2Fji9mXrKrwWwBUuJ0a7AzemrdBvXBlR7
zN6/rBBRA9uA3f9E7luaLbFSOmG7GbM4YTNyfxBjoMXX/4ZaPXpUSMMWYfPa2zvm
NyW9TPdnu67jI4cBC4Dx/gpcdpqrp0LoQgRBkigJXYN0w0s8qnCo8IV8hCieBH4P
HWmtk1JUZNSKn4sYLsQuqqUawvJRDQ0cQj84bKgmSdMyuE2/f1J1t0/jVNZ3ZnMY
kzAMu7f0d7liTO6xKy6J549pUMFnl9Kb1rwkaoDeLdt9b7r/+gfbhQpO2Gs6ShJk
7fM/rUClMwKSKgaRUyoMyIyHxUodaBn46FkgIn/Enh1jJd5Pm8UoVEr2xZesI7Vu
5oTV+1wFaYifaR5YeEcS+WlB9nkyAkL98eLw7v+Eenf4SBZ5UAivfz11ZgwuBCnp
Tgn5VcdpzuFIL5/9FLaW/6GZzIY9uU+yL57Eo8fEsQfv6kXy5qboowUiGB7+c1TC
laM5bl8STZlLJAqqNtd2WLFAC4ORJuj299ulvGD1Lqqa+XqIUbhUY6duGvaHFDpj
TwrOuD/O8ksetpPQNrXq95yIcCd/oo/MmmiQ+odw/T/LF12jT2TuwwG3dKlJ3XYv
xp7NV8+ueZawAl/ncftjMKPxM5MDdj5wczd8Iop57jg7+CwLCWGObHrGBG48UcxM
SNaMUF4EUfN1Or8gLWtoo2OLZYj/00+vVSePbMA/Hp/ZpPqEjTb0QKDKQhW2o+kZ
uweCPdMfk4TXwc6qUp/xY8/+kEoWwbI5FVir9CikqEu3eho1HwJKaLuKQTvdtPlF
oj4N7qSxp7J7owK4+MRwkNWp7DXurxJURjGum/7w7vEIY7xxk0Lep0jCq//pf48A
yq2jzzioFjEfSHsuSjYOVkNJxI3/YKzId3KbCkU7U/4vALKD69woo3yS/RNAMcrg
oOx6YMSOOG54iHjgETj4gJ4ipsEGgGNEiEN1HztVOXtwPK2wzd8CCCawN8rstnVb
iMgClrfUlQT38IOupFKUkj4tPInhSnB3YGqf+HNhUFqo9PCrAHddf5/rq4uFwwUp
7HrAt7RlcMYDg37ZKncIWOEA3ad7A8Z1u0S/FlURFCNF1uOVjcxsingblRndUyEv
e614e/vldpaPPE3F9N/1//Wcn/4SKi2kbKPfo1qUFV6zVP0loGHcOX/tWvp4gTTM
E8/fFkbSiQcpOoQPajRf8Gyi/L96CA3o8kws6eN95jKpCNIkeKcC6f4KADHCgUuL
s9g9xsA696Otp4fKKidcv4TTEVLV1J4G2LEz+F67xqZQy81sToJZWSZwhMKfLTVr
AKPgaRMYZBAwkD0227oQQqj0v+SL+IDJNJfueHSL5gT5OSsHxhVP1gZ9GOwgSLmT
JHsYWSPfSdtO0gn+VUe6vYiMsh7uXotbeiNOVlYJqzH8gH7HzXZtM54/XjcjK6Wj
C4TWa7sOOtrfJP5zN8lVIR+J518ncEfLcseZ/O1TtgKez3AjJlk8ZT+9rIUtlR7x
QLq6aPYugkxlcEA43p/U8XIknKRFKovcwBBbCgn5EQ6b3eZOLfJpnCf9zZEmrBMx
9GgoJp317oB+0MWBmSPaUO7w2QqCHI/Ahgw8aDAyCj9JH+mM86ysNO2SRCNkmM50
sk4jy1VunM6KLsk32mM05k7g8vEWV5ZhIecY3JIfGugW9PY9r2SafwcntdLOYFi2
YWIXoMWB3UhqhXf/riP7nFSDsunHymopnX6ps53Kn1CBmfEDw3Ok0LBDcpDLXsY/
BvNarP23TvcfyjY/d37MOGTPI4lMPdKHD15hDtNZ+cKi573Lvr1vRVI+jGrgIjum
L/vL6n4XH4AWDiJQ8tNXwgC9Kkm+fwPaXPORxgAcF6w1CAPEOGWsB79MKKmzUJoF
Qbu/SBH+496CbKCsnpP2gdTDy0hhvrmuB3OwUz+wCIjtpkbMYKBawb33XgbXo1+1
6M+zNo0oqDYNst4Opi5THAlqghyoobFeJUS2H/RNUmauo6GCStlUrCHoAkglE03B
ksMYpoQCzPX7vPcgAMxZe7MWyXpryLqpm1K4yrcdEJD1iOw7qy1zvU+lroYo1wi0
HPS5KnHi5p3E0c2fw5gwnwfGC01xQd3uC2J5Vx8i8Hy/m+5n49LWgpuFDVjD5FGb
dAYLIg+5xe6fZihUZz9r93TPdJzlVkAYKTrufwgXHTT7RwnXPBVJzYlo++E2dAkc
/7cAsSKjyBVMN8iGCgQfUSyUHs1bammjBDxByAW93BBITsbV7rxLiAr5KIAWlQ+A
3D9k1HMJ6AL9HGn+E/j/anHqfezYHMGx+kLnFiu+QUdv+uKh4bVcJ7VL0ZT7Azmd
Uig5xvtI/GP7zwomC4LwFfAHwMVXqk7KxCNjdzXdmD1xtaALGSULR4/kKH+Rtslt
xOuiTQoCEieOV2td3QPIdHZPd0zbi3ccP/E19F1UCVBS8U3+mg6xNXil2sAfAK5e
DfJ0IenYCtlaI0d4mJD6YrK/Z2NnUTPdyzU1aWPQ2nLUDb6i7P5vG4ig5kMYT7Km
v3lseSawJPdy+v5oU9zzbHLenRqMyBvz6hzAJijYRMxpTuu4t1Oj72Vng4BTAY4e
S+GSSabd4gluBwVklgs1XedG5m+AjNPBhrk6BsrIzwp/eWFIPKyF1sn0Y+Uclomu
EZ6PpH48q9uEdoGhgDs1Rt/PTLUjOOtzQ3i5U/yADx+UNfu0L+va+/VSovpxeePw
wLmyfKFswABWsz9ml90CwZfb4Ejs3dzmq2li6BuA5wojVyVNY80YjAJV3C/5d+La
egIoXlgLbAIt+fH+cVxHn1+mL0Cxm8DHC58wgKrMto682nm0Oc9ySMVOQemKAnv0
pH5wJ21ZkQO5yLHpAguWMy9mIVfzmO/PhIp+SuCycSJ7JqbC626xCAFohBJ6WWuH
2NzS+nW7iGKlYl0agE9SSsGoI/WQNX1dEmuXHhpfjpBQIlvdSFxcS3ptycCJv43V
vqf2PeExUOhEdd52sGVXjqgOmR3z09esTnJx9P85cry1i60bHbv3cr0D1RLxP94l
qsOMU0Xlo8QSOT4ZRkbbzbEzJ/b0e3wvzSSgabyp/O9Iyefowoc8hfsfxAX5FTvi
A1p9opMHJUr7DdOidJc9VLBBE7UiAP/S155JtK46VP7I+V/+uD8pjAJYk40Z+WAc
Bpwmt2fKIst+ejcblmO0foiAD0pfjaUS8NdQTzZUlYcUNKtxfAwz+zMkjic1+zl/
UkmQF01AYcv8QioLhiMEQ4iddn3SG4FsI52a/AXm37tO/cZn91AGl26mkhoB1Knk
mV6fZ2/qRn5Mlhdt8EZdcERMoI6/HPKwYfgEeVf1JQbBYbhcMwKBCz4MkTNbpMKS
L64fXQ3hNqrSaeoh2EdxCnDVAIISTh2PlIWzs2sP0M77w6pecZnQ903qjAjoLDQp
0g1CTAPcETQnf2vDRMwd8+vYBGHEbGxWAWXMcjDlZPVATVUHTmiuF4qbvli/LDDv
y4v8Q712vAfjq+GEYP2dn5umUMZy2QwQSDcxkD1Q8UZRPlalS2I9r+QR0voAA78H
/3Uvv60cSsVlEhfWrLbkLIjpl5fyzFa08yaeRVC4PTHu30u8UGz1mm5nBbrons8S
UPJ4nx+rLqY9erksTGNcPbVxvkQBXFCX/pxFnV3hks7Di2uwY/VmRmIuAA3imJMA
qQmIGSXFJ6+f0uTv0YWjVe/LI1oVUKQFVMk+3e5a4/OQQ2dxFXqY7IqSzzmfIqb9
v4H522T1Y9CJqV7Cf7+B9o0mBCqghJyGQU420a6x04NN8gi1eo6EqrKfBgPrdCw+
hdKY2f4m3Anrsee5Rd50spGy3RLCyGJwPinB11p65sRXfE0qqY8ZEL/2yWNs5okU
kZKwQa40YNCw08IkKHdRZoU2YV5CjZls2ET7J7houia71Aw66dlh6/+yWX4ZJ3P+
8EzByKp+qK4PXgcA6hE1ISYjJYsfjVpkEeoS4uMsIUVmEyO9x40eOxkWpmeJsG0+
0JdeAKLnt3+VvMOsMNiL1aSDGrwULQwEyZRHDAzKDchEiFe+17OC80ZXkm09+o+3
RAfOFdTW4k60RaGS9wK7aPQdEnpcAg5rZE6a1sdE9zQ/MIHGXlNBnEtbNI+6X0sx
RkhCv3ivzo9SXUwhqxv542dL9lGZ3MJV3RjH23QjiGIoafvaygbLTB64/XSzLvNB
hlD1ZeH0bmmpW9NHqMlsCfCec8d43OQLjrRcNPC/NHxgaoE7bN1qaXhHEmbqVyaK
76bIa6OVCcPb2Git5pg1U7+rfqinOFStE9kcgTN/wtmK/XqChAHb8NfSfoztsxvW
k9mOcyEJE0PVE+ZAwogA7GGV2Fc2oVWT4EMIRq02CNztODqZd7NaCoqqEjFAAOgt
g/0OvnJjP4z5qtQ0xDHg9nFvvjcXNvHj65ZTM6DE5I8/VyFQTjpgS5IY3g4wWmNZ
0QY1bYKy7XW1biJ8SddGHTUUC27q3C+3ns2qRkoNDcHZMN+oX2zRIHDArqWHPXPF
wn06ueNa9Tl98ix2Wn4accYyeLn56YCecYHUf+dpztd9qKtlTq/pvMW2BVbkgjCV
Jk0xE9uRcYiUhzMyBN23PXQGqjvpG00VI4XQBBIkxzxFuTCaNsDCIQDtZ/U48EiK
oXG896lsIX5suD4EBFOKObRPTsNpm0mwf5GzDLQAIH4+0DfhiPvulPW59MYDZgJF
LdcTGN1B5ET998uWzvLV+D/KKDHu8H0HsM3F4miqMEd8KNTjR2yOti/k8aV7utOm
rv1cGAYsJ98jeEJXpRH+r9mV1M4Wsz4Fpe5I2Gaf4fwkEKTUnm1yRpkygy8AfYJH
7Uj5U26yiBQlXlG6MCr7cLTTsdf588HVR9wOq7OBaOrO9CIkarKXeVjJTBtAs3s6
rzkNpium4JOArcpqgpAV8dzyqbQTT/sx5b/MAxd/Gl4XZKm87yj3X018cbDFmRKz
p16icNNpl03OetzYEDJUHM3onyrrPdFZXwlalpaI775MlUvpuiSZGsX6aEDg5SFm
0E6j9oaOuWyPVo1+Eobs51MV3XEMrE2gDrDWzTs+W/w5XErpI1+HAjbSDhawTGTL
ZbiWatUc2RmUUHEpfF/cRJ+jayfDrHVAudv5ycgY35U8hbdNIgF1HIFIgS26Zx/V
y/gFMRD/vr3J5jk5MSjjuwJOSuAUX8ZOEsGQVthBnh1bfAlNvaKypCk8DlLfoWGw
uaCbmYVzfNBvOLRwBtWxqpKDj+rZS3JcW7ut7rQfu0KbXzfmJY+cQDweVHOYEz5y
XtuBuQ7SJOdcQd/xLKTj10lb0rDVNx5vcsFLK9prh2rVsdFhnyd5dyQiHC4dbvUC
L5uOvSwoefyG0LgEl9LiLwo/50LGtsTKHXrrbKOzzJx5X7qeSrxVVduiUoXH+VZr
Qv9QRQVDVd2AKXL5PZohvcGxJ4Q508X9DseaAYBlRL4Rn3ZKHHMPI9GYL2yelMVt
7pjUcqaeARI9bxGZ4eEuXOnWfuFGpKHvqmko0qjJWJKmUyGMUFP8gg2oK2bztGmN
IojkE9670UIyTInGgpW7kkadfoJYePg+MKhTX2Q2XseY3k+6SiSkh5fzETwQU18L
9V12Rj+ihhnprKxHfmkcFzOCZPg6rvwr+cHYFuoGRBPh/R54lWsFbXq8SchCzBEx
luS8/Y+J/DUkFE8nPSIh67XJg3T56E8WMQrMyU2bjOf30K0DRecspuRH/yqmfW/D
xRxexc/TeunarJOotKMhef3Cjw2AyB7WAsHsoTQN8IOmWfwcuBYK14y4B+Pbfqr+
LvhXwx5+39RIpiEuQaiwEPRrcuQcJqqWdvzJWe5D8bAoL/k/TWFvgIIMjJMx5RWP
Mqt6ydmidTtTtQc24sR0RDsFH3v523sR9y8Zrmac4qk01Kg6bMHDQCZWwmuzTurf
a+LPlEmss3llcAcShYhV87ZU9/pV2U2ns4u/0KFUTJZ4fAPWZWuy4kAD5FT4muoh
hXhVnsRA1pyrkZ67rvVxi+SIXgY3bBsDkgYrGmuvuHrck6WMjgzSdCqSqEqxu/RT
hGathIHHxa2iuR4kJhHFCMvW8ueNBe69uieZ+Fuag3RauwaC/YFM9klDsi8BGRMr
birO69VsG3U/53Lh4XFT+Kyku12GNher+Fl2XP2npY176B7FaeqKBabsXxI8sl+D
wzoyGH5W5K58xIYBYBxJzsuq2d8FXnpkK3RYv98rfQQHvJtolEq4l6Q3MkrZlUit
e+kR/mSeZnVjQHFAaPNWk/HVU/KwC3IlPyXII74QYrfjuD3WNrkkGsxnp/Hem7uo
vGn+zW5NHyokKKe+hOu6ODKonDWcybDJ+bNEeQSJ6AycUoeFwlHSqNQq1+HBtcIh
jWVRTdcQiGi6mYYxnOf4fZUQ6owkH04RY0V2EI2XByOU/neXx2cINpmsDNRi0jpX
7X/1FB2lSy1emS8ltIjRVH+YIgqdZnmc44quPdy2ZL/68w/DrtOkE0CkGI0yNQrp
68NY4/pu7mdOAtOD3rvrFRtcFKHiSYDGyB8ZqesZSlAon3J3R34M+a0QHkpwfNFT
Gf83Ie82cKJyW1Axkt0lrOUArrjd2dTtIFqHrDQU6Enyg2s3oJklUXsGxDyXawMu
PBMfdU+x3o8p2rdPuHHjGNtF9GKny8+U7QPtJ1f0sj38eUeW/aGbTkhJWCXN1kT3
DosbZ+A3ZmOZW3GVDG4Tv0my9/8Uej+tcMOcferbQAQ5Om3dYTm5AxipO9aaTWYQ
MXo+Di2ssADjPI6oohPB+3ZyOPVeKuzPP8SRq+GeWz28TqaA3DJ2mBlCgVC0QcFb
ctq95Qfj7WxTLPE48Nfd7qO2TckaFdPqEtkZYuagssg9W5V/CCuBjlu6DyVgErzZ
Q95eeha5Z8u93lOr9r31qDdsINIZYA0w14FdPCL9KYzmkb/1PcUlieNOi2aIsGc5
N7/tDj++wKYwMeywkoJzG7GoOOe//4Uj3nw9yd6vS9qfy+z8dPGDubN7qi/y1Gn4
SkkrGf81cs0fabkz1WwN2FCwDAGRyawPnE5tCYBWHETQUI6ljpN91xoHN3s9jr7x
HoroeITyqqvOJ/22DM2Oow8PF4EtPPXur1LpUUZjAjBnKU2RLBzR7bq7ODOmU9gv
Y3rxV0InzuyiJqaFHkXfeH/O0v+Qcndw1RJQkZnygE8QVFGWj2o9/lpavHIqPMSF
kBB1ooLa2yA/Sh9N1Adlrqjolh26He6F+usOx8uMdKHhcGd4l3yYiJMCkD2fbUHh
J/zxak+y9ilBHV6Jn/y+MqdlemsmQWEp0QaeeR09HxVkFw9W1gb5xKju3nUIYLAu
blRBqfG0DYfb9fRqOIle+w9AqePeZVVK7eIb4FundCOAGOvHM4BQ7V7YPqHAkAfe
g6RYVKfZ909mL7JICeOEGW8Oos03lvyDnBY3UhXMe+r+cGyvhOjiei4/clfeAs0r
8ABbhWPgKi83RJyy1g88DZBQO8IPpa8eq+f5HXadMS5MibnAp/AV4Tkq2mVUvAxw
DmW4v7McdyjKDTN+nnY1F83Uv2iMfI/aXNF7JaeXJ5hekZU9bjY7PaXUPZVsYQtp
j29JI8MkaI6rwLZB+cK9CwpDONSDbaWiFMxNzHylvxyfzhnj09gRJRgOoZHA6jMk
BxSzTDyVrdEf04yImUcQ8RognGFWVFU85YPlznqYPUb8SzfKAudxAu5c7uq2Hqg7
zro4xN9k60RFntaFBEcTNwZaSDqXKmC9M+utK93e90x7T9EueGb+aSDy/sEzWkTM
aln6uc0fANPOvRhIfvQTLdNBf0b1XYh/DK5EQsiYXN+/kGuYyPFA+KKInYgRAiII
wgCKod+Lp7MjgEnGi9KsSSSQlHEOqD1+owPhCpU3M0Skd+YLgf4bANHMHQRbKZZb
DsiPPqZR6Sd+b6wuIhACK+R/d8HV/Viez0+4zAIIJgrW1J4Uubj6qcE0+StHIFoz
zYl0b3wDGrH7mQHveQV//UTThIX7+50EpHjb39b5HjQeMTn1aabDOuPbfazDQRA/
LfhHSrMjaRTDeUNn+HRAEq86bTzvBYEruWIg5G2CnsiUW9dylqYChshYXSH0XI3l
MfNTyS8iiBxWjki6kHIK62rdmHnUdjPabqJLUT9+FJ2tNaxZnnquBt8rvrZ5lC47
TBo0N0AaDju0ragAn4x7iMHmHaPIlzzRfCoPqiQ6VNEUatLEEHeitQexusmjWyPl
sLfC2jmJVFAsIOclIwsIIWTTSnQKtTWGetGxsmzjgCMqJ7f3yTnJNJqkuhjVPpeg
yPXlL2kigTOFDuNKwzVL0P/K4K7VKaK9SrHrmhB5354o0VwPzOt/jqThJEiS1hTQ
v9Sey0MJlHMBzdbgEELW3ScR4aD/ID98EiAqw/se1s2xcbJkO6jYmYvqdj2Bk1If
StRh9oPb8R2o14gZLoVtSmIDt5EKm53qBjQMPLkaNg5d9R7Nezzs2J5NvsAJ/FPd
jl0KBCLhpMJl0FgX1zOHGcqBKmqrDXgeiTNsUYPMyvxtpSrylzRwBlAhodIxV4yE
QIGwbir9lLxiwNx4UoMG8DQ/WdIs3+aI9uqStvzfhhQ6IQiZXHnWzQLZtZ1mJizI
kf2cSQHzc2zJ8HdtYZSNbvHDbZepe1/rgmik4EVeFYiJVb41kyxUHx39ppyVkg6K
Jqfqa2VMNpqMNGjIIhuL0x/6F1RPPezXEstrG63v3XG/jgPvhnp8CrxDx5nFD9tT
NcjAAuB7QeWZK3iw61IPHgEGEhIGda3t48EpIctxRBCDkxparDyd6sA50c4nSYn9
0fAB3UkxtfAHjOJ43y6SY2rFVFyRPDsrE0sGAyCS3l878jyT0ElFS7QaeDkCVp+C
BwSsou9f0JBCRG24ANFcZZqtJGIYmoQUpwuQ7hpmXXAA/NrcQXLyGSwtWUvTHnNr
devlghbwhSmRUpe30cZT8ZEvu46h4Z5aNpxzxjGIOhg+/TevZEiZwcHBMdSn3422
ZQpsspOu/xCYdQ5gqCCO0Q/J07ZOCQGsg7Ox++xMHm1fcZnlrr98FORO1BXbvncw
MJAmqziX9LKLoluZzW8ENu29hA2RDCPdFc+pPnHr/0SKWxNrKc6cxvXP2HaqGMiS
ZAxAr5WBqNP7ej7SBHAy0l+hRRLWmubKVKvPh/Wal+bNhYgEYcoXiSYLyYgQzIDv
7F75cDU7OtVJmezACx7N+Iqbcw9g/JaenI+WxX0KZuSlyQYYNBJFyL1s/mPFGi8r
cVF9D/XfM9ZwScKsNMXKxg+qVfAT4CecyDHYq3VYi9UXRt8GNgeHM/F67JPM8VIT
7c6X+r/5e6jbcn008/cnGAQHjkKy8OjuRYx8ElWwyHOpO0TQPJpfKeOHKRWGZEy8
OHr1RTynJXlMJ8nUWsPCrqlW4a7DUGHQ60u14gKbTxbV5egAK9BGBsgwvpdagHs8
lIiAqJblvyUqDhyV0rF3uU3Dh55gCEJJUaBGFpCACmG598QGjSyOB4I3KXZLcQI1
rTfZVQZ0pCTQpzbgIwtWdCTQ/VEq5JuNi65JahlZQOWl9/98P4yblWeRv2+2DRMR
ae0iB5EOikermqB15qmWXoL0kUzo/BIBcnwu+krP7I2P9qCfd7DgbQfiQz5Or/Rr
4jKcJoqT12tsLGdUuDuxEJmCbhigxK0xzFoAQDJ0MT1v4nLvIrAFEUhANl4w6l3J
Cu9nyQdbxDkC/SjCG/iKxlmntfzouWRlHj7D/RpuCqH4H2TjO+qAFMBzjQNAHgzd
qdHQhYOmS/xHbAT6RmZzXKHSOLfASz2o9CS37aEyl7zSAtSKjx7AgHMMmIQS7Xg5
WRitQ/exogYR7oQcgMjXgUbU8JA95Fiu2H3FOr69O0qcq3pufC4zZRwQUyZpP1QC
vOBPzPMu3atvaUtw4Np6bViLx09ooAXpX8UycY8m8JDjBawRHzd9iEcrXxy6XkN1
TMI0lZ3wFCSlqJhKaN8LKLmFZKBMVfp53InM2PVU5V3zHf8FLHlom3jkYD8+SEGn
vfXWq/G852bYAIf1mSFy3ZQljS0kkjTPKeUm1sXRMcUMlP52zzBStQ0UK72Vn3KH
1H+1YBliutfVdOFMPjWyHvP6FypZ4yVot3iQIO/J4d+apm8goYW+WYls06Xyu6Wm
/Ms4V1wfz4QKAwPASHstFKq+YF7A5f9U599YX73ifKXfGWNf/DksZTDzGIjSyGH4
JcwTOszXVyjmUOnsAL7SzjoSlhSNesUzjhMSerLOjLP0Y0osN2yqrT2h5Uyk2cpT
ej3OBEptGshJGgPiypomcwzVpARb3jpLEuL1iwpXnqSooifDca1dwSFMM+qTmIE/
GO+ZzrvBevxyDpLJOCuDq2GZ8Lm1HG35zgrcYsecGmB0Holc8Ug2mOMUW+giJemg
DeOVxKxAyJDYuDztGMzG1dWfl4D0hJ4LpqoTK/h838aqZGVXSwvp6FZ/53pyU7NO
88LA2do82f9emczpSkSBgXOVHq8cXR+zQ90W7L5An5RxCyZzjvMuaAvq54TJXhLH
0+x1Cj2gKYq1NgLTBRP63c9si1oWFu8wggMzPiqxMTeXsI+KExG1HTR3IKXY/B8Y
VyHj6Fa2yZToaJGsih386viYHtYWSENCQFwqmQX7YHj4/5g6qX5GKny+eaoKgE8V
yFIXQSbE+VtS12F/7p8YG7oEwcTH5CHfwmNrDSTLaZwJIuZDbJrbw089OexE2EHF
ufI+1vgHT3pPtZ47hRZTLU1V3RdFSZNYk/1xCIDiV9mWu9o94qiEt/plnX6YQaK9
vDyWsdeZHkXu2wm/mSe8CCQ9wPS/2M9Rq1wccLfHaGbeZ0jFrT19sLSY6fQ9WYSo
0BHLfQMDZ99O1RbUsuMT1KzeUA7bOX0YbttN5p3yY0jQKV2lrZ8yNs6BkmeVPLlQ
7PC4vOFygBQO/ququMzFpEgtDJ4Nsi8ucpiXvVf1mfOGwmb1B7oogmnChBPzwUx5
8fzqvDG1SqRYTxg0/A7h7DWXriblATZpCBQDC1UTWaYbshLfbTZ9WDD6+a5GSIwA
nql2VTr9IPJ7QjUauxWMO5oE2Db/Yf8obPBvDp0VVlVFEoQ8pdxviEbwJ2jgcfA5
ToIA0ZaTIIvExSsPX/aMZBqZTaFqv2GKhbfJ0hEBqGAk/V6KNTU+zERbqj37UpTI
54HlaiO//jqXw4g8UVdBFdWtCzCe33vlXAWL2wctuFkIuJ7EFkQY//pjknXof8Rk
he5cSRnisYjXlf5JwddUCVwysxn5v+JQsxqc+96r5EmVZvxptZoifTtVGMkWN0yn
grFupXS9PN5mQ6x/8hpzD8xRLIaGUrCu8zEPWK/zEy0XcySak053h2b9DFh2rJei
nmYWHBJldIJOBTuoRbsABofKBiRz3reAVv3lB2pdYWv3tcKZlL0d2aR3Isle+RLT
avSa+4XIwBRbzxEKyeGaWA+JiJK211b/Rz3+1OLLpfW1gaM/io+7Ltt0M3GYLRIf
yCMtYzvlRyCTWOkQ0x8KIYGN6m77ogkLj8lW67vHILXw9SzvxQedd93CKGe5jShf
tZKTeUzIEmRrgtwLy5HA0DDIq3KV3MPBOgSdq+gA3z6Lik4Jv1jZd7UirOet/UNH
CBKI9O86Og3pkTNGbt7hNOBZzLMbGvggXenzYcFA3yU5ih+WKMo81/t27dX0kRqi
3mH4TXZOixb6yYGxQgRFEDAuODNJmXzO1p2buHtIYb+lPmczPq4seRkv/RopbJOU
/u9wUBVW1Zx7ljaDQRQgoGvblbVwv8PMWEztZPAI8SHNqPBbyLBHbxqHl74j+uCa
yQ39F0uYPntstHfbxZM30fUgspNb1UTpQfiP6lFjgEQcmWpr32a9PUkWGIxnCZO8
o58cEZzksQMmjt6rr8zdWpiy0titmx7uM+N2IMUjhEZ5BiHCf9B2QswhX3mX2G77
PiO6Pd77RaWYQsrMFNPmCfOx9baPnJtdfCBciLuENXdB0NsLIwl1TrAFXocOqsfF
Vnbsf28ylhmnOS8HqIEYCB+V/FnziHbfVtx0tvRTGno/zHOYGO4gmCVTuhUpEQ5k
98KPCYlXB4IOkK0ctip+kSxa0BTGpKriRWjMzNwyanMOJ4F4RnHJA06V6h0uRJS3
ttO71aztbeIMpoaDiN3eWImzLy3mcioLCz1w5GDk3ZxNQtv18bZtY4G14v3n6+mS
Z1f4eHrYJUGIyoQetQLlazIhsO0rRHNHKuSKaZV5k9amkMWXQ7c1qEj67wnsJwBZ
j5pWE7vkrCQLWJacjW5rIgG02dw5NGTKtC/bHEMarUVm8FTlfuBM4D3rj69GXNNU
7N8qBw193Z1jgNKbZVdMA2FmTXoj79dqEMNFuywV0HttxFQtsmmqjt+LK/c7cQ8h
gGgMAZk5n19zY3O1ViAlMlPNvJAZLEURUHxrkdQehC5bGkDLY6knYp9CR+BLvr3Y
fPJRZYHFxjXVaxXDRMo/XgoToZzW2JhiVfaXcIG0d5mWBHNASH7VRurHqWrwZzS+
/5ZkPM3kGzLJ0bcaQqJIItepDIFi37W06DKgqrCMYMiauTxnGpuCezawwAyRwusm
KWyWBEN+ZhZ1p5TJ+F+F5k9fYCmp8PTkBqbmp/Z+dtne0DzJTsXnfnsMD261M5rO
q8AfgB7+XwoS+rfKvRk5c6mm5P5hvoBa0CKNbbn2i82kMXBYY9EEijgXqasu3aFO
Rdhy0NE3XusU8JtgR/fJitnyXjIj9T1jotq/gq+VklMBacZHXRv0W4vJ3+05rP41
ix1H+2H9cJMRvuzRVag+dLLJddohGO/5WIB+Jf8cmEIfF6snDttdxlBBNyJrd1IQ
AZ3czQKP4PCVyMFvvysS69Fs8deffU+d+oMOWYmR04T6onRjaYRmSVvyJTtDYEc8
e5jo676wjwNTtNRZyhgGn/0VKiABwkP719iJiL8sDiuBhBVsGReYeZwrONdxqdqP
OavJyTx5pMwodeJTps04my6mMgMvY/u0elq2dYNidqe0Ow930rE9RmkxYwVcwPEQ
Z7LSOC6AXV51qCBBa04Sye26JPna+LwQ0Sil6isYR7BvWwDj3gRtpjNx8acQs4J9
ms96dRlRPUaOsZBQPBg1Z9IC5KqXEL9OeKq91syZLg9fcBiorDTj3Qsnr/vVt38z
C/TkkvU5RQ8GW71Hw7F/q+RzxEWAI3VX5lGKAsAo3vFU+ok3FRhzxJUIofQgNBRb
FPYWgZG9PV5A5y88XcKmYao5PErEimvsZMmcT+f4xQV2GbKoI5OIJgt01akF7gfN
5nXig1MRLa9c8ucqqW5INMIidxZ9GVmp2zdzWaLTPkUCS1zLFtSCqjujQBacqV24
sK8HqCwx9IHbidmsV86J5sZw4lyeyca2jJ9dQSS590juUbZBZmli5D8Mze43KBTs
Jj9QfpmCgk7k1TIGknGk15xW+6oV/PHpBqIOWRCbcfopKB5SWMRUOqlzWPe4GPbh
nEVebB9d2xf0fD7u2kVbSv6vLr0I1oacEdU5bmlCUA3xvvkKhi1Gag1nu3nK0onX
SbWLoM8BbJ01lqYyQMwSJq1O7nlSkCUoVvqLSOxHdiv5Dhr1eTaX44RjAD+gxhBX
0b8OVaIjpV6vWN1ahxjG/sB3EF7e6P2REGkgJkX2GSsF8nizmNq2xth3NVENku+Y
WcTrjI716ywICwYfxsO+9D6H7BgWxe1YUdRQPokuFBMfsuyPxaFxnuIKLf2g5bSp
OK+FPoGDnp7OHsgav32ciwpV5iYcWXV5+9I9lzD5QClR83HvMQfStmxebErfPD6M
PYvD9hzB/rE/iLcuHAyAxoJCMEDFeQHjkQj/TTu+PdMt/T9+NUEx8Qn572KjxdBD
XYbWGvvf+zjXxs8h8TO18V5Q71ILPzse5eABpxnHuw187Tz93/7DUfdY4f3Zq0Ig
Z/7P8QbqTf3e88SEbOVRy5VnDo/9bheCoFLeZg5LRzlsOynUhYsfbgUNopubRia/
5bPwLWkDlFa2zv2XW04wQnSUPbwu7BytkcULSCJ8xvhXXudBJCiwmSmpeMggadZ3
93KYkdurJFpQLVi/4qdncPtXw3DInRB11PMcXjneWpdTHTlrXHKYjjmZL7MdZ46P
FsXA4yLGinqeUrO8hL953L6Z0gKMiH2zShesUvDPWDVvqa8Z/ZsxVTqcR1q/aIc4
/ZdiU9XVKipPYG2cW0ra+QOsNfv+zr/JPWc6NHN+7Yt8zTVg/0FOM8GgxjjAi5nx
nQEH6aYzSvBIri05gQKHUjOsTJm6TTn8FK8mxRT5Q6TiYIIi9CizCyqZ4Vjpv0ce
AZ2L1DElaWNiFr3mP68TYjEnTn8ByIud248aFNyeFNGw3iqL0yXQ+TAyyAamopNS
E2QRyf23HdePBoPYY7dRKOvOAD6Pxavmobat0WsxfoTkwW9yxdNq/O/CJa/ywftD
eqc1I6pOEFzOtr5p95Z9P3DikJzEqAyI+GQrAps6N70BNgJGQ0+GdWQZvlmkbV24
4FhEKx8RxfZ4EtbHti19RSV27veA0L56IHt7P69cr+y6egdI8sMjiFis10gH0Mok
z8gLsq7MghMsReZzu2bIp9373ZuWJw+FeIFapGYH2ci59e2SpeN8hd6VtcYGJ0wy
N62zN2MszRA/bflc7HCFmYdb5bRdQJPOC26rGbJ89bNGkrjJhXJH6BKGdSzw79sP
XAtOljbrK2RX6zsXD6WwcRSfOdRj7EmwJrCic16q3AnUGK3fD3U20AaIVGKYdjXv
xaxYnrbOCgqU4pkJP16/SNW8IRMFkBttnxGovm44AXnMm0rNiEopsDyrSx8n8R+i
acZn9S46xw9GW43LjHZScMRI1vFoFHOAfEu5oZlTkeBO5U6q5pD5Ywix9ekbx6bQ
rAoGcdYl2+hxU1dsIRogm/BhtBS/nQmPk3Eoko+WxKqPCIC+KUuder/BwpSgOWDP
ZAgJMECEoUlvcdSZDfIVMA2jYIyIHvmFEn+icH0KUhYhYTTYrb626m9COLifY/io
6jkI2jWezR/ulxDwnjnywvp8OI1eAsENL1ZhA39r2C683WldXh+4lQJHoYvr6aEc
m/s+YU8I2YJzuupYx96TGnEGTT8MdmQg9glOsU+W7bBPXlQHUj3eSRtasqydIIBy
8bG3OYpr7WUXGBqqYjEKYDYKdS5UxDarRuz/C47CY4glQFvP8K+TAvJudIeGf1cZ
p7Nd7ZBVx2zxp8i00dJGtD1DmtE9vziVi2+rwEa1LAs9Rw6oPcosyVlq2AW08QGF
mo8Ze7Q7eABQ0rpMaAWG8/CJqHxtZrN4xg+lFDwy/e3ctIM8q+0flUH9IvPzDtyn
1C1Mrx2AnC1QcSp1BgnIU05wQQA6HqmYvgjEysE+0brbKrp+Rxx917GKnIQjv+DF
E/EqGoSdlHr0Pa21f2Q+4WF78tGzuuevHnt7dfhXjLdbllsIs7JfLavGez6QwYpt
RBlB4xkZ+bDRlOyzqt7eOno/EmQG1ENenI7XuS5e6wP3/gXGK9h/n7z579VR+p+M
gSujlrwAMKQuuLG0TzYipIE4vYN2D6XwKw6UAIRLsb5HIX+WM93k8wiXi21qZ2Sl
yw3m9RuSmJtNPNiqWsBNNGAhRVjbfyVfD8JOMbAgt/Iy6C+95jV6B3EceWe97g8g
ZdwAjqDk6ll5mHPjvuMvmDhEdWDx73tC62GWAAENHdGEZwFjU79V50UnwbiNTH3D
utAsUfMOX7Ht4hjAzT9V5Ib3n0lCCidXQG8MiJfG60m8Z8aLQDkxjEwBa8YzonKM
rWRuhp83FqvzRBCQUwaZzOaI36q9luDiAijT8ROM5SMZdotEhtIItSYwxYOovP93
mpL9KZFBGlxQDe6A9+fKi7Ohk/8XP+almpVwHsZYDgZnuaxdpdKgIBAOQn6LnLS6
bE2XXyPnHCkvS8NP04ojH2vQJz/x1MOHmGESQzDrXNO+NpHM0ChE7S6Gjt32lsAf
Kh2ULXMUDdEJ/XyIvrJf8cMHiFAPEO4T/RVNaWeS+9DBMRJZAD6xliSmv57aldI7
vpETHbcin4kde/7KxnuhbipsfcrafvWU7N0kZkB+LE/AuEorbisZRnJ7GE9ah4xk
rpPBa3oe05UTNb0Dgw6G5f19CW2QU62kZQ2UI1A4YtFLQGUgcup3sDH8aVDHWs+7
N+fNixZGlwgPujsrY5NCwXadbkMpt9ZNkuRppZk3EW72HZ/yfSgtdYpgU1pQsbHk
edNMQiFgEQfvf134tzFAEh1WVDhNCKbyDDfAWNfRKEfc7J4VKX90dzjho4ddUPDS
5udLHyamUEgJ/vE3HvvWL+GtbZofDFgRJAYc2IhJ5cXt7QKVMadn6ICtnEjUt+Cj
cbWosBHRedZAyQOFONhv9Aea4KtmFT+3iYDMgaQj6lJEpTa9nlVpbUjVRoL0gtLw
QNr0Ug4dBWvh26NP7yzcPGzeiwIH7218r/xJmWRXFErnsjTpQdmxLGSQgFsEj/6/
WIloCkQBwZfXXSg/khZcC1fysMgR2qbdKHcqp/qqrXxZc7hpWmTFBFs0Ai4a+YT0
63LmdD5LPhnQPbvCrqGZYrYzKIO0hCIAfPXNcqhK9nBr9soZkb8Hs7AlvPVW5J6P
ATKA42oUc9eCve33NCJhsBuPrsTrghMa2kqRooOfCcQTfQdutOZfp4sK4nBQ4PJ6
MCkPlyfmVAB6OIJuvLFtvkG3qfCzKCKPsbE7LRXoluP02gw+XrCEo8TPVNY77WR7
4WGb/xHmfi4PAMo/WESDB/ttoyyxtGCLDfe/A6dPVMSzd9QmivSgThMtrnu11/Jl
PSSdt2h7ejVnDF0J7bZ/IvsUoLYI9xUI9ZAF0b0aGeBcwUfEGNP2gLXyoFVH0yhC
nODj6eka7MScX9FVsaDUEauOQ5xfHFYAIF3xG7/L43rdE3WHDuCXcmHPCCMm+Gh3
W8dDniEIrkD/mnHanG1BgTCg1fPJzZt8E8xYbywJ8fsIFI4200vwLfYGYl8vNLhd
gGBogG4d1Da91jbMG+vMkyKWZ2w45oiDe3LuCVF2mg0QHQDoA0iyRXUxARZcKPbX
8UJ+L6WZjeV41yfIWFRXDfk2K5dejr0WjWjJL/cGBuBKUPGk+O9/aeIqTSIFdNL1
2LI33xgFsaUpeWR7P4cCcZUY4n1MJANbzsWP1DjX5oN2qB9M5RTQGYrUFB0bz72/
B724YUzuPqxQb9VSKP5+mW8SNO7nAx3MGhbW8/tFU2rQ1pdZ6WUIWuDmUtj/7BLT
VCmn9b/YYJT6N2Z8/xTWgmZ9HrOk8yqaZ4Aix9mr1Mghwe6TT3nzLFNRTHPsFLzm
JmMSWhWw1iMKKy6PpJ/Phws/EJu4yqOSh5PhywdWxabSjsXHlFFe10tb1QuRhDIb
BJTqmis9ltMeNfUlrVXb+AyS0bBhoeqGKa0P4mIqQkPdWwk/njV3lrEwdoqUa1C9
/HHXPBSfdNTjb4Hxw/7xJUlb7UxINm0NLV1J4Pj2kjJEimUfo/T+YO/PO57QY8a5
d5AzMFStWPLjeA52fkQ+UPT13KuGqj56SU344u6vknV9GLyyLOYAibL4hlxoEUZz
f2u8rBCTO2FNH+fVNscEnygrBQV67pNtRNGqF3cWT1Q0x8xmCmUDmisG13oDaGJ+
f+7fOxzEpcz1JAs7/+GSpLz4pon4KJOD7xDSMxeATOO4gxk7nulH51EBej9xkSwD
P9fjNbnX0W41aDYpdDcgYFsM+tCiKTQkM28trzAP5k/faRYeWLqqI8s7kzG4g4SU
Zy8oR8OYvCYbSfEtVqVxCfsBzDZHZ03KlqYDuqYAquJP8k7ol9FyeZVxYj4JdFCB
O4nS8gcEHcOk9IFDM940f8Bd6IGLJq2maRTYRq1NBm5blfokiM+aq3Eki/kjSqJI
ZD12zkr8lXsFl81TfyaVrdwPJAYJKKmAmNf6NRW4FAw+WWBMGBFZYgEgLUUoJvih
vIF7wNbAAsrUmWp8UQV9l6/+w83+SlpLri4PsgwEyCkgAUBVR41P0Pc/gChhZuFl
mAncZ2jh7DM2wYIdSvDfvuzAMin16jHtosVLWjrIeJlKHgoSHdd3xGmsqklW6DsI
mfwh+I2K1H+DX6u0lSglbcWis7gGvlisaXwOWIvEZaNClWPo4z7Dts3RGQqpCUm8
JVgJr4UB7XkQ0RhgfBcUJOx3KF2vd06IVGk/hLOdBLmgpLfK/ewDYkorCdKvwDat
EuRVQc7Qn0z0CFq2fAqNyE6/xBF3BzQ4sXU+lcXiHh4PD6xTTWShjPkpubBYBynE
VXngrGWYdWlYxQBSy4UB+dhPXBjOWmznxYmWm1tXj+aPAuoX+Uvc4Aj8FRVTwWMV
TFosrnYL/ex3bCW88FjUVD95wNBAMj3XWML1b3KqLwuTc05+kX6AMJBGzac/yExS
Cs110Fu0XhCxN58CAirIqeUY4hTCariRdp0ptauhH+ItUWrUNzwygRqvQffh0Ltt
0YFA4DiQPFTS7xfRlKtfHXpeyw3rEPppwQX+GSwXrbI6YgC2QseiSU0UXTCYxTE5
vsa38H+4ICCxjDyPfAVa3qoJFcHzKAVTsfRibV4Hx6qZC8ZVAano/FvqvnYgNlDX
xE6R0PbNbjEeGn81kStqCijHwYVs5BsBgTwijgn66y4e4fiUx7g7qsjZpZhmL9aG
4BiX5jpG9x9xezEtWjpzi6/4Z5TW/fZM/gfmtvsc4y2vVqR5FH1nj8hqz5DtNiNW
Bhaz8lNNm6LLhcj9X38iKKL+s37BcgftimRZ2ZXRJcMczTymr9NIVhCkDJ5Jvmv8
nDD0oCb+QJaYEqXqla0+didTAql8KgroNhMlhlOGYD0MhvhPfKHDMRn+RSE8RzeE
m9usKBVTVSJkk96X3jXwObw8CC45fOsbV1eKzYNfjvO5glU+SokRH0l9MBv4tVaP
XpPWI5x/mvCuLxiWNSUanxCvyzu62QRsRPJQ0isEXVnvYVu0B4ZyU2LFPH59qb/U
f6ZmmXLcmWpOCAf89Y+HWQ83l+6qMkSN5jylDhH207mKySnivRyFvX4i2N6XIadf
IRxUGyu+fVCemdkapCpR+biJXAxJ6dsZQYbYAGraVngpA/GYg6fB4K2fv/KBv7JX
OuoLHgRxxP+UemMEryjS3YB0sDB/HvXwBMQF31fwn0Jb4IrDti1SV0XDP+EQG19K
3fVv5O4EsSWsG0UrNstN1aBXjl1URHjB+ive7ZIaBzeQe5ZKVSYPgTP8BXwFm+M7
sr9FlZSZDXkayQg/XUCYNsOTradKRthFFZSVoAXYzO+JsgHHOi6lINkGk9X5XlhV
QH3SApu1O1Q1X+WoGCB8hMlyfEtlqnSHrnE9DrizoLX8uRltF61vepdUMhexKeeE
wifWvsY08bt1bBlP7B8xOx6Iuc1OuJcQnHXlbmNyOdX7tSWxnU/mynOxY34WBasr
kxBCIkacAOvwmtpxzTfnjOYCpIXKg6eEalvEcNBbsCf2evL9LKk9m/uPxbbrHMdp
mBgB0mvwoKuLGMnIukAnaRLxqlPjRKXHlZPt3Z7VOgzKOfrwR74B+RyuKlNxwo5U
dbTYVo4BYNI+B6KpnkecL/zPbhg8GcgoCVk5FrJJM9XnNeYNIWGNvrcbe+oLpaOK
Jt6LVa7NbQUMpOVKSQx1wcwDAme1X1F1risls5s2tCozkf2GQY9jh3fVVOGIkgWb
uoix2GWvK1pOd++dOacj8Qd6mPNFNGj/F5Lkpy+igRwum11IF8JKgU8xXa0DycsJ
7dubYaMfHphilMsyENK9KGCIXmUhBD9lpSoQokGdTL73vx/0RwJv2F4jfrhRtl/B
E4qk1VHk4nNsENgGRXrFI5qcazTO7RTpUaX/B/9xOTqIHNU0EfywzDqMuAuAnR0R
asjGk9F4CAZ2Rqa5WMm90+7DyZok4yPtZd0Cc9c/BT5yQwYpdTI1eWesOIZCJmUf
XwthW75OKK9dN/M2rkXrCWrhaM6WVl7YjP8g2TvYoYOjLlT+tfzo8tG2nl80s/vj
vASevYIRhQ/6VNKqYY0I2UL9YH5WWZSrAkorBw2olb8I/L+6IdPeP4TnjaQq5Dis
1i733DcONNZhpWORJ7NKB0LxDBvKirkWmqKHQDMg21GxJYtIQz2mNnab4H+0U8j3
9pnYEt8n8/leWtvB6C8F2M+VONowEJeUN/PIrctg/Tts8x4+kMGIUiIJXycaY9PJ
3RIgOwssZXjED9jd5nxXm26hV+q9oLt0u6gllKuc/zXc6sZSY+3dle6DoKs8MIyZ
FCNYCG2xeuHYRLB9XjaP/2pLUKR54Gb1z1ODzbCR/RWJZh1A74MFKXSRF4DejqBA
zhdEFW0BMNuCmrEkSMvMGLU6PCgkLLJP7G9uRH7vuRt54b6hWMxJE744WI1U+/K6
yci6pxgXLzMKcHCZVmtt7cl5pI0WR3UBOSMVN7zt2GT2HMYaEYkSujWzniY9wmq4
I6CiHGTCXBNonizeFFuAN9oqbMLSJ5wv1hxRNx/xddekZ2F/hq0AAR6NX5mJWZQ4
DdGxpHpqDt5lsK3v3mkV/6Ti9gAOqz/M9nJLZqzhr5wItP5zctNe2JR0BQGhYplw
JcO7CUBPFoLvH1m7zg5v/Y46GcW3vDLDrUcKSefoHbnr2QzkYTX6N4v1zRdrVqVG
YOLigGOVRSVJgAvPva4FZeTQwSOIkEt/ISZkHBJA1Yezht/7Lad8mtyJ/DNe44K4
4U0YmfHeprMIVao8Yxb7dt2i4mSFh25opVIfBoyaleEB/sRZG+pqmxsvGR58WEDZ
8vqk6rR0P+5ePu9NLqL4fKn4D+hTtXKLC6mwo2TiysxU0NtZTFPV5ZIqyYwxvii0
4ujrZ5XgCsY2RKlZ5jEvaHeRvedewne/nPrzcNZHPvAcl4e0ekKTqgXKWzwzSVSI
MYOsytdJrjaXtXUHqT12SR4iwBPa12/xAUld1fa7y7om9HOUCoKi5Wawcjgdma1q
/ZMniMKaVU+MdC/zQlsMrINZOT8gVjetZmlMmB0ZktHJ055WY69z7aa6grWW1ocv
K6GHvSkkQaiqttbtq2VCcKOxC0N2mAUg3q1pscyQHU7Lbd6d3L48xRnT5RViF6mJ
6YWqQPNF91yI5TdSromwGIcB3v/JDIVLO+FtJEEWC78tmhPPI9OC8IJMuX2OVaOs
h3prG9LVZqc2lE42lIjZ0pnc7KdopQzfg1qNovA1zXB+61NnBJKIloGggMXibME5
HFGSJjQe5WTr+DYLTQ8IkotPpt3+Bs5g0G0tIUNgctCLG2iqKwqpaJhicWmUUDY1
PT06e3Zkr4HZJbTXhQNl0bJKe/gtdxQKLeFhcWLGU0eb26w0v7+Fd5kacXH5DHxL
dFXjq/eCWt5yZlj/nZxQkLLjndkkS1Wx0CKKkUecVtYDanYf/FajX9focXsPvh2/
F+exHsS8n9LpWQRWDwJg17w6xL35vQIyTv+N5D/XOTUxSEAf/Sk3SAOTmdSyVOmf
YggY7wK3mIw8CzPU3MJP/IUCEkVZd+w7le6L+JNuLSDPr2HU5ljr08U0wg85//Pg
YddxoC59isVnjYZ6IfqtIOZBliJMLJmlR7lMwb6IkWcKI0//e4aqWct5dY2g8C0d
+5YjssU+Y+tYQ0JloNQnhDzliBoGeYgAQULib0BWJ5BlNPxh0Pono8LQIZ83kw2+
ckMxi0Ky5/vCA2+llzTTo23oHp5rTfz3J42kjzeMlqCpH/KeM3/IiNw8zCFFJHu8
fsK66fcMCh+Upqc7Se8Asq4N0+WBRIYNNS0IrsqKVot6o9SWepPCQtN2iWbHyGx+
Yrz8npmPCp1b6KY+ErCVduqCWVG9D4Z5cFv9MfYsZWyNVtRNUkU0821knhyKUoUi
eXVxmAfto4G355J5qGCSf1lUOKSwCHY9T9WQhQ7elysbpGICK8wqWFFW5VxUi8Uw
V1YlxTy7d9hPqUfzxvQp2Fpo5SlAjCuY58x/ZtjSf1itDLmo/dPog3dhIZAZeR5J
ZOp8gHtKpyzapMBKgibzWiul6Ffl1WTL098aR9GCMjDxUyCdCjqFNmfuO/YUkGK8
PuDEmSZhFgo13QJT4uZX4B5VnGzyAWjVYKRQtwD/RKUMOweVd1/Y93efWebkh15O
NIsIcTzRM6NK6WAoHDpDczGMPmzL9rZa4DxB5J+diVmByLhvU2Rf4vAMN2JlU/DP
aLLJYXoMJKfNh2rz4RlnSLZfSrpeS61X2q9MwbDklbuGUFB1uwiHgm3sX5b7vNF1
kx8MrWK1dh7GUaD5xIBtQNquel6pzs82ReLMZbGBa1J5Uam2if+a4yPyb0P1qmH9
sGD+Er2+7/oZd33EoKAfeA+9dEVbSLJry23fdd+an5fgU790vRypPCeo0Lu5BLL+
fLEBSjubP/syOGf55TPp/2tPCp17SUKDliK91WtkEWGm+2y235GStJBe7mis+qsx
+249bc33ffaBHEf77vaokyP6Z0Ksjqc0ePMllQo8B+nbDxE+ETRaNsrCwz/cjH3F
vAL76G3+3EEDGCIih3oIa65VX90yNjB818pr08aMsfFWqbHJJXx8jiaZTWhB4GGc
jaOBuFYmlAQKj5Y7MQfKFkbYW1UNweyLVtoMatcK3P4lGpokn6nffNca6BtPLQVZ
r4AFZaCV2sDPbxl69oAWb4p5ZOuWDOufY+rDCPktE7v9UI1+IWe88l1QhCbyDyS+
cOc45zkGdE4ZKs8teUCAgSMJ0jym6URKD+1CuKArdg3Nl1zV0cujqPBEHJjO7nU9
lkVgHpjc59Dbf4IIQ3ofa74RXDKb7RD/5gsZYUcGNss5wMEvktS7i6EPVeYlEpma
naDv0ezVj4tHB2kAezsEsU8/shGza7SkH+9Yne8UdWYmsnwnzJejiRjQQejaA47k
ifN+P0+jpI+6r1cvEAGEkew4d0EH118GcXfDgifIrKe6iLtZJUMePQfvzV4S6MwW
2+AWEkeOB+dYIF/26dEcW5Wd6rPvLIk346cCIchlZl96C3yCXgiNy7hiIqtoBVh1
fx8bHys7uH8P4CMUrvjMEihicbA/WeiWBhM14+/0a2y/49Y9+sv3mXobJ3nSWDyF
E8R3ugaR8ECSBDNxEozpBvMpUN+uqzwDYt1hKaMfRn05HKISt53GNzp+DC0Y4cUh
iqXG7w06LslimykvLGEo6RL6gcpGTyevBYEw09fJIqqYtfrORbHSszjFaE+CtCiZ
9C4Jf7W00UfhZm0jSFHMXu3TN5Y6TvnDZb7rEgSJJ2mVvbXQ5PArOQI+LuKszv4f
Env9GNmWCGYxer8Aoa62gvK8nwqA3VDr7auKL9eFcyfHtE2sra7QmZgbayDV2u5D
bKn9KPBZM2Iovaq6Tz/9ButzvCXNWVJLdhAQxQvNZTKeiQ+D5Jwgd4p+ssGXMJ00
dWYDE82ibxt+97NA86S89lErGGAKPD1oQ3Y9q9B0CKq9y6p54UVXLkrAXDoYr8e6
TJL+1t1nUL13fxN2Y84PLklXNsjqjFB2ca5Ao0DOLKeicMokqV7HP91wD/pt2oY/
v+oQWi60BzQHXfBvHqMuj7O6NTmLv7AVGBhCrLZfMU7527//ckqvlP3oB/bGQ0E5
BbWn6Funyd1aYykVFybIGKJ6HTKaQks7rJTv6Pkjdpd44qQ/1mXBTp//tBvpUNNW
2I542Tz0tNXjmS/VedgGEmHk3Neb3lFuZELhn91XKgzpVnnMF13MKO6viB79r2w/
/9oMvNUt42PlUcwjcWgH8kszPivixVw9j0s++pJ0sZhe//fvjHzjzo8hLZCDznrp
atFVSMBKrGE+eOCHk2/SjIJImIF3PIz4kLg4uwGFK+gdLKSNlk6f9i5A37TpGQJD
eVM5BdMjboG0VdH5b78LG7GsoP+hLyaTnfoNSXaZM6NZXN3kJ8FCXeraUAd78DuN
umGN1U90BBrVsfhZJw0T2gPhRmmHtgNfXaZ8+oEmD5huQntFmwGdxhquryn4RTUm
3JCRX07vIOu39x/hV9pfTdXyICN0moFvAHHBNTSWOQDCbyDnfKQyO99YLccUqCpf
ko/Os1qoG2tKIeKChsfcTSn8VQJ+fRnNleRjCX9XZml/5tqK+MKAhcUq9IdiFw6s
6gL/tXvTYYiHK/b6kItXmpBudV8wb/33NnCao4ThtQkS7r7cO4TE5XrdXcBkGHF/
jBEbogkvrz1EYpV7u+a6OkR9U9pSd00jjamTuIWz91zicvItHDbh8SMq9qr4ec2n
3LRUc+2lwnknuVgfZJUMGzVgDVyrcxBdqe4zdBFqGiGfY8lB2ql54vTQBj3jUZGi
mHZeVd9xn8155w3FrKo9wouXA9rC8M3vDgJ30dt6yiHPQuOo9vTs6gWWQ1tYQP4c
V9/CeQXFGsJKapVogBtay2xGqbU35e55fN9/KgZKZdloMq97cPfn3UMFAYjp01De
4nyfavWQBaso1gjTvKp3r1VoM7LBRyE7J6U3FgluJknJ0DP4JODBxnTNUaHCKVQx
gE7VcdsIazlI+gaXHIcr2hPALzkLA1ss/yA7MqtJMzSVPW0kXaNm1xY7HdUJHZ5r
V2vlZ2UDfZ3dWBUzbp125grFwIVWJp7/z7iz7q+2I09Ds5fCEEZjj+RS+xKMJZ8m
UPsTBul6qYfNaGmri9e6X2jPcELtAFLbDLaE5FA86eilBcn0oP3/C8QuhsLLji+e
u5BN9ZQVdo68qoPztrEiE430xnyCcDlBwWofQvOIU+uQatjrU28XgYBbSoEaberP
E5PlH80nYMGe1+O/+91mivGfMBigMJJLp3s2R41LiL6MJ1iNqKZfyVxX3ciKGDai
e4ZTSD8kEEuQh+W1WYvKtw29gFOMU6G0gQ2EM/zd1b6G7GUaP0ogMPnC2sZe5UHv
1EMP5zftYg29ztcHafd0o2ljLBqd4hmTOY+wpc8i6nIlspxBE7FGCH0Bb/c8rAWx
l/eo15wjURLE/+bVMaa0UQmiTJ3gc2/qPnZri6sqsG8GRMlTE7IzJuquf6E0CF+M
UE15e7587oIHZOqfAQ8uK1fRj+kZzaVXmYqw4vYVAifMTjEwurUidNPPAg+jl+n7
6qOg5aWCowL//DO6KAJnStY59T7gqMYRii+LkZwpDb2h/8hlclrtsOk8sjTBQ7EU
CxqjKB7H1XRgGpS2mVHGNKT05SF82wdzyxjeOBVoNxFDhfIsEmJF/6WfI4nVBXbZ
HRR7AA5NDP/LuYuBlYnicXXsvkjiuLta5FkFwda0PNt4KC+u5eukOFQssKTX+4vh
8K1q7koyPzYbN2dJkAglhn2s8CPS9QEw3mNVVHYbgmD+35kvpfX6RlFZyALu+1dp
ZRX4lNASMFrGnq9kO5v11F8ETV39W5KX2xhuBiaTjhnN8CYrXtFzSCIm/09Anw/8
3uY+kdbktQZImHimY9gLO/yS0mK3ESkdwff7ZJ9le9LgRGPLuafO/RCdXcTYXtoN
3zAVzRadnX9YiMC2NXsQwnttB4tQtasEW8ZM8+VsALqmis20lWFzaHIvZgTzm/oO
UKpSqfA6O6tDTibCGehXe9Jhj3R80CCgO5A8/cqO5BidHdp4lurQMH88Dh/GQ9pn
YtKrQqGLCkGLVQHNLVonruhrJH1i/2W4lq2NIAoheoriZf+s5kPfX6lbbMrKGDz3
en/d0Wb5KfkudydLGQUSMg5/MI+MmY7UwD5HsFrpq3dp0iPHUoW1C02EFJTQxEIW
Dh4GxPv/uL18AbzuFN8159PIJxl3P2h8UVBJ0sx52Cup67f/H6Vfvh+3hULRwJqw
JQPDNcPrUFSpCa5kvq8hFfez87z82KG9JO3r9KxLW4AR3q6aQGTcRWNNfl6eAsiZ
EqR087T5SrWzYKYzGZ7Z3Cwwtz9Ddp7WvnzQOWhOxBgIUK4ATHW+J5DJcQPchvg2
0UpwL4l3fmIbe/Q62EDpjHtDCoTJc0nrFwcENNAseWU8MZ1tW2OYyhDYb8huxvAM
qP7dJKdyZoKh61ajz1zbprjueFyKXXu7j/QEIBKMi5kr/hmNIMreMrojUFpOJe4O
TZEC7CG0pIT2jpe4244SlQco9wb4F/kvoNnWHhRBL7zwL/fLdSjywbN1/RYh1Wto
HkzIcQQ6160PZtywmiKdrlD5CIKM7UqJiNMu+XBF/WIQ/ErbUT3XF7JoKZlSiKpn
s+u9AXTxwi4KZYSsb/bipOGr8Lgy365AK/gmMvdx+A6Ekvhk/JmfMXOZ0N3GPqV1
02fvwRZX2gtMokG1FjMsQ5C+ADyMav4KrPpSXd5wbj9WyTYZC1l7Y0MfpZvMd8I+
74iHNiaRSLH3o1nWBRm0Jp3vO2WQ/ItFhAe+gCg/DYgffKqOJDEfEqf5OUjGgtqH
iTf9sY+0d7BuwHgMgXSlnxw+lowrsmnLl2EamOaMXc6yRu6KzeK87WPj6qnp6O35
rOiU1d1zsidLd43vFRAYwwR/fHxE3IN5SzzV1gfrKYjW7R0IHOE1z+8v3oo4RYEa
nhng3+aiiSeMhs5ukFz8/h7rx3iQhf8bG60SanVvYfq6O4wDJIhrfirNcLEii+3b
Ft2T+12TeqwW/eH05EPGDD74opAVrWbKpLTBwETmErWOg48SG7C9d4QghneaT/v1
VSEr/8nwv54FlikK1EBJ519Ku9GwTDdIzObfoy+Xg0shBmc+a8lqDrrg2X9pYSXE
7xSxjBJYkuTfnH3o/eNwrzo4jQeivszQG4sj3SsQWnJTVZD94DCLuYr0YTI4n8wX
sS/zrpIVPCc+CLS36AAy79zbpqiAtjHv+x9RPeel+8Mj+6jGCGajz/tToFGBY5Qj
JKodw+QcQz+4QlLoxpa6HQcrq7uoj5MpETLtSRrwWK2M9QJfa4VkbhULyYvHvD+q
uGtrdS10qXak4gXzMcRNc9Q7bXYqnhkpGyt28L8fNFmHSpj2RLtYY7JTLZoHq9DD
QRAC4NnA05xkK2V3p8KImIsYleUi10uinYzDuWaRwVT5QLAUYpZ+G9Z8dwdbItU2
clMH/mLX/BjrRwNtYTwIV43eFnIWMIg13C6P/nt95MEwmlSFN3bAMKgskOWi2Ivz
OMrOi8BGhCYjcBtBk6tsA3hQDVqooKiclvU1glPI1WLb/fvss0RsFSU27ItbNQFM
9TC6+Kelog+lzRLhagACuqXFwRbl6oewmwo6HSFxurnmh7erNM51cJLKN53+bWEf
zN7lweCZE54eMnCS92yg4z8yitOdLFWopab623S7R4xqHP9WOs4aQi+fB7h3VE2i
Rz8NYoNGnH9NyalWpbKaXokFISOTAj1FOBWHTovEZps+CDjTcpRmicYkfhl7/fvi
qnPOT4RttkmqH3JxXghFkWgslEQHtk2y0x4mXseEvwyqypXvev8GcyedORFTpt4q
KINPSlMU1mSC8XOjUnhBY9QZL6WGJUyoHC+YTV89O8SUUT2u7zELjWzuvV2GtCE0
s3+0KQJCFj9NV1GqJrW9Oe4Wj6y8APoKlAnbN3TB8BIATplwVd/ILLCCYzssjsr4
DbXOFLnN5XBrnVFhLvB7ARGxLhEn8WNLP8f1j3RTG47ghUni+wec5Sr2eE8bhT6F
YjU791vsyaLz0JoulR30rqWUpKQiW9yFl+bajlMkYVAPLqmXbVVkOcklUaPftAPG
tqLrucQhGIQsmCNO3QbmSNhnv0ny4Sa4OpLxI6g/qXTACVuSY8Q4X2cGYqluBbYa
AU8XV6GGifv6vt9wdt47zYaHKwE8lPwFxARSplVd6mrS1Hs28YvOidJifr6bZycy
oiEva970jFCzeGZds75d+zLKGCRF5TmTvhmTfitfmNl7v1nllCVCNO9yWgAIb/cB
Xe9sqZP4Nqr3Id1YCtGlPlGvbaj6bIpgPsc+qKdIooujR95GfEAWLmjAvyRD+0Ri
yBz6kVE9uVNVkuTeCal1ghu1t3E8dXFix3AEdUVF8deBdeOKcvr0ujh7wJ+5ZV4b
D6oukiTn/nnir4C78bKDVG8+cGQXayCtFijk7ok4t+dOefEvyp6wjcu7rOTmIv7E
7LzbwrMKFH+5obGjrubQ6HoSZ51/JmmcIDpQ5LlSg/dJc+vEVJYdJU6spAkwJto+
RJJ5lqDC7SKYatg0QWTmupfTxHEkqPUBOnNtfujKOrBkJfHhETa14Ktjbf0tH8mf
NZA53BhtXtg2piX9gthzohW900LR8x7ORhj+PEyYZZGaBuMfD28g1DACj3SYZ2le
8fTp7buulQ/NqDt4zQfj7EvP0UdrBZ3aLduK7GXYwokHq97Q0WCIvOKKd6z4ra88
vgV8m8HGmfvXyb/dU3+T/iIgrtT3ZLnpHq/+Hc5a5qjvf418IRxlF2E8rr+1T2WG
MxKVbjwD11VmPKRSrHSDOkt2foED2bFAK91vDp65NtoR5bslfMc67dPiVcQKSkbV
GSpLtXwF/VQFLE9ugPRjYEGdl9Pe3nk8gcB1Gm2sdbb/678z3Aun5nHxGgvlXA5i
BRUE5kzR0xr3dtp/zv6X3aZN9y94TCzFjG15rWueBqN7X6abpw9fJa9X0K1P2ym8
o8ZxjMFblZpzcaa90fVbwMH59W6V7GuVhPZ7kbddYq0sStm1uOLqZjIHpq1do+px
vLCtrkHAi4H8ixHaxgUfTFc4j9XMDI81LKjOOUNzvnlE2LAyrp2hcHc19hfF8KiC
usCCSKl5SiQ0NZAiN1ZZXEmB0VhBPH11BufaIPVTrpdsMUzvN2mo+XyfuPRq00e6
goC46e5QC6HQtv8E5es6AZ3I7tQ+kKZH50oPpzB70ey2r6wdPlU7My58sf6WrEp9
jt9wzw7c1EkLVP0KYfiph3+DeqO6AOrKdCCjVgFsny4MUv+64XLGSvqv4eM4Mkqh
ES7T1vVqc79U8wEymGemooIPhjQXZPflEw8mS3oQIU165t75VjZsHg8KAZRPQ/8p
Ye9NxaZ2RPANaj7Aox5tD7hhO4l0YTcf35uRkcNFOwKpS4np59jSckbVLV3Bt3EZ
NT91PpRMGE99n8hymOkhQwMpZveoxZclgznX1cmtlmC/jkumAP5I5Oozms2XSnIY
5FmqGcpOdK2bYVPy0gk1+YQHsQ7fGidPode4C8Mg1RcfKsso+8iHLwNscgj/k0/R
gL93L1HE8puJeMPt13gI0QlIpBbsEoBbj8NDDg6zZHBQnhnLjNefboz7uqO/GYdu
X361rwXjYymRMkGkLeqcbPVbXmFToPd8E3TF+VIjpHlmLFuHADJz/kEqdkQYkkZb
dpDRUczT45ZiTPb/R8vCYv9/dzUW0ErwHiGnM6MmZxowPnC81/+axgZdHVlUHfk3
xTDcL0VqUXOE5ot1faJ5KmcuDRk9D/faRW7zxByux/+ZH/ga6f0gK01U4zPXmO0k
TwGV7wSeBZ4XUnGIccxKCmUIRhX3eqec61sH8Vj9mwW8JxSfBsJwTXdtCFcK12JX
YNs9PI0o1i1kKhZiEoEzi8xspkmJPNWJAN+n240ib548oqZBP18C7u2uYj67niD+
DmTTKmx5OmZ66G3Cun3BmvTmSApQKvy1snE5WB+zBBhUIkYPCGK8X3HX2c/1741N
VQ6FvkPs+wlrhMbxs8lI3ynZhYc821dkM6Z8CTsrk+ZBx6Vx1cjmOTIJnWEEOGRK
+iMsi7i1TxS2WKtWFxkCmavGvKgTkBtcOUxmuikTfvT6i/xqk4VpZRqNvElm3OQm
YF2+1nnlamO1LfHzr2VQIwbJTuoFTD+0or4Vk9kIUFDEyO8qexX2rGaKlMiHENnp
Xlj82679AgR0kEiKPTAdyhg3zYvcqPEY8VHEYhlX5kj/N6tMNoqEWysEnownYy/3
hn0woxlGqIpP6L6TeIqpLaHskbaCvKyYRBIlIblSNh7a36XUdL5B6tR9zS3KnYK5
WSv1MZCrTS04XffeSN5SwMt+fym72pMIZyF12ExSC+njc7cbPNtrDumaAHOa2Cfn
kHwVWC2t1aIOQRv/1NmDIyoVBXORTQi2wu/b7Xxa3cDeSp1qjStqEpsvA47OSXcF
U/OTbgqiW+JC77GYmc0KipthBjdGwiPdb6n5lBRFqhV7Q8ilE2tTG0CPvJ6AYUSn
AwWpYclGZO69mRGC82BAxpetGhR0rHpFJVuWFdH6WHJ4TSESg3BGmtVk5WY6/2qE
Z6Nd/4AWxYv2LF4hUObbWNZvhXhI7x+Pt5Ng/Et2ramWEubWf2AB1t4d9YpptkEh
jp7u4S9sm7MzHIJEuGyamnLt5Sf+qMo1KqZjUD4bS/vghs5nNJTJfy3pwmykv25/
b0HEECcmhu6ADeX8Po03FUy1eavNcn+OWjSaPCYq6dEffB32P1XTlyzU7TxfSBUq
Z6AhQtu0cCclUs4RGr+UrJofp65RM0MpY1fyIn3ieU/hFQX339zDWH7lzDTs7s0q
hxoYgBEfvI7Muuoy9AZc5NCMis0gvCO18dlr5C65rEzpu71lKWVEHH2y4BcZ4Yy2
fwzDs/vxEgkTX93rchDZzOQuBTKNc/pJTRl4jeQRGAMtXODiLAES8AP7xzX9Fqdo
kKrLx+xx29q90en8Wpav7/abyGtIAixqjMGjDEojTAd3nFLM+dfzXlSQBf0Cy8jB
lZ31IZ6UUaE/XUndmgMse4Fxg5L+3VH8iva17QbUy0IO6h/xvYIiVPh5YJm+wqD/
WPH8mOKRLsvoMZ2IdPftQN3HixYNuZ1L1YPRvtNTIQ63e0f5J2aXh4PqpnWoGylK
Q/PRtTRW1bIu8unSU8ndh1Qouigbfm8/IMZTvJMLUdACSE8/WOUAAt7WOcnypxgn
OZe0ueWpx2g0imsUT94iz8I9Ppo9DFrRIwfsf14JxedcjvtpfR4+YmzNROk/PPyQ
9x8qBRfLfiPo1xZeWdPc4Q7zk1mVlUv89+u5FNhCKRBVd1ttFhnaeQq5f2cKieIO
f3Y2V29lECezJudCgmQx7Kpef11hGcS5XvuvG6wWirsEUJDlXLai8A1gVXK9fpV1
NKdIf37YeZMsJD/Vk4ECWpPf+PVWe/kwGzjSz/+0lWhpKt51hQ2V8Ku15AYYmJ+a
iDC/ELUZY3gZPIpXpjzKv91k9KVT/Hjyn89r0LC6bKBkTJkU3dZk1c0aqNlvrZr4
pOKtjAFf5/76MaGQKwF5HkxoLBNSdr+lsF9QfcUhCzVLvfAKAzASYi/HQpxZ5Ocl
brE528aKnb3KzJgI1QNASUYtTGTIY10G5V8ilDE4DbT1LqUYVdnCs5i8y7bhEBNv
xRnnYL1ar/Rraj7cWC9DMNzg6BB7Oy68VMxGHT5kd/CrMGgNWSO5+xDOXC7K8NHn
Wh/g7hGW7gU79Z8EvldFtCfjYS9tQVeaKEtv6Jw+cCmBCn7OUXkeokN4fWtNQtjP
A+v2g7ngn4zwMOaqKtI1ARiwaSoIXiX3QAa986TsSJ78CYcy+qOjGViEpKZ+h5Nf
guoLB20/jVXd1GfvOdVNDKtxIlszLFAG82aD0g/K9Tnz0a67CegxKmXReLLtcFpf
1IYWDYL899NJdSrJ4VBL5npY34kXcUs+ylRjZV/puVpHWQPD1ZN43QSepUj2AEMZ
ca3WLI3A8ZucuyCoCQQHfJGLPQxxzCKl/kYcP+3rgsnvWPYhen+daGkykXJSxhSW
QXrTS0Ufo3bdB2cyTFWLzE0fzXpI6goCrkO0k46/voqQyd+xrxsU0yOfgwjh4oDv
q0FX804qZzoV4KKCEWN04C9R4jMZ605j5ntO2XJ+Slm21IdjaQuP26KB26nCqTTP
WYdEZamCoRsXslH8ILGUs+wvWilApm4x+i5+spSrzHVeM9EwBiHt4haDkpAsvNbJ
z1yy7C5bVJMa3QmeJHbPsRk+kgrKtNoplkBC3XNAf3Q1xkmS1/eKZuZsBYawKCS3
tGoSC0vBz2rEpjOeY/bv5A5ref7Ui6X55wBcaDIqhq+TK1OCPB4rNNPTTtizw2/h
9duUHNWLjTwlqr2rxXXvjn/IC9l7xqa8bCFkFa6OYKea0vv34EjVNyebcFedkeeA
ntiCT47X1ZSFinKP25DGBK46qCLAD4SoCLOWICqjUDjeHdVYYp6UBddxi92OdPmk
YnGdBVKq+qNxIldU++8KQLjZPhEGlvBKVlvmqDbEzww0vR1VflRZf+a5/oQcnlb1
g33+5SckLOeO+7KS3H2E4TvgWzq8Yvc650HNkmRqdpJPVYpcYFvXX2fHkJ8O/mqb
cRJHKfu0K7En6+bJZW+fETsrs15dulEUv21HjyhXzzkiu2H3XeStyTDfTa9Q+3FL
P43uXU9iU2ZVwyKyp08psmRCxaPSB+DH+KK5f7+fhCq8VTL2WBgdSU/l5WTbQ6o9
iIZWsF9ArGCDSLQJ6KPetUjBBbMhcpyMy2qyyzCOoYaFtvl08QF2pZ/SQkVzfVhx
yYS2Fu9S5vtzzIdIxuzMIo32D+h7/UbGLSW0c0M/iIFGFf4yFKMHIFfQeg3kASmU
S/GuTYvH2xckOWf4c22AEwghA4TnNhuHsK5WkBxUoJX0hHFKHlEZn/lSr8ztGigG
e6MmwUf4wZScYUiBlGcJ4vPrwi0/A8rBhXHBTE0g98rsKuEsdxjNStZiaPMrDixa
MYRPFE890TgK8jpVzPK1LTK4RC9ifha9pxoQNEcn4+SQYz1pd/AdvfJCawMUZp8Q
91nzgTGDgqj+nJpzTEknNf+UZ89ylhr1uZPVOy5khwfPJT5GytHWtN7cBaLkk0Fv
q374kpA/6LFcw/K8GWww7PtHTQw3bm1MbuB5x70eUoaGxY//r7m05qi+Zwjj1mrk
xBYENbUusdBBszFvPmqpaY+51OLNvTcrN5fVdC9fMEOuvOX/IQFbN3Jso5X12Gty
RHcVmB7ORkhPmXIjYyiVff4PxTtlF5dy7ecxQhTsSAvC9nK3eUqN3wbyFE9I1UTx
EGilckwpnyqmATAAAV2HWVlzSqV2IzDnU88OfjphJrRXI4b8SkF0Wq7DLfSkjzYj
W54S1xORI+YbEmzGlAto6WYidbAWIZRPrJYErkoo52brSpcYg3OuPzrmOAX8Pu1U
L+pkEKSp8F2tT+70EQYLAUyLaznE2vrtoW0SQA7p0JyhQYjzDSLTDx3zqO9DnZYH
tnocLKesZfM2zW2itCZAbRbYpF0OETdCHYooXoRUPRAgRrUchqeV4Cluen6pCswS
exxDewJxD2QOUePc++KITmZ0N2IWZwbdvgqGndnLzrt2S6MauIAhUyJdHnblBwZE
qyfmDHOGF4beUCLFU5hYx/nWXFMgiXvaQqqqQTH8Kgg/499eZwaPTAB/ZGK/Syxb
jV8tzBf9FunGJ73x0kXiq+z1Jf083YcorQ4L0CfVv9H0KAzfOuoQIpoitaUpMIk2
CsOrc3cUhSd91bpqvgKKQeI3hDauFCQplPyp/QGJqpvhC1bYM//ag0xsk5j7EGUw
+4IHiSHhiPR1XteczSrjOkipR6L5WvSf0Y+jV3x+S8wKfZyC3G7BvcslZl0ao0VN
/5MTEGrGPntmn5ZZoaJmL9+apw130Z8VWYgTyq2FdPJApcPenPmTvMuTURk5IXjs
ylTQCKsD84M0qI847XhKN+aI4u/jAq9plB7Zw3q63L4fKBIiTZ2NU7KjYhJZl8xo
WBZ4rrCftwU3mjarYpjDZTQ4GeAmh/rGad04+te5sWIHnttXvvgRd+WwYksbPRm6
+J7LnmDqwJnuWBcUsq/KPTeIwaiphqil132jPYlb3WveMo5MMa24tOGUzyaPxaYO
bnmNH3YspgvNQQnh9elaOosDXHpX6rWPeJ11Df2spKG+vhnLUcVB5wWlGnNjCiRy
ixYOzdxcI4qwb4JtFpqshsfRI1QxldPbPqunK51tlPxTt4X8puZIP5kKfevxwu8H
MTGMtxJRtXBiejRp0O8g/tOiZN6KJSaBwgleqj1rt4fUfKOOur591+Qqjzsn7HHb
0dxYOQ02E8oOM4B3UexwEb2m/u/d1Fq2VaegOJiSdibMCVM0u5sfSTDdsaWGqF/I
lw6JI4vIk8WfduBL0lJxdE4wUE5THBcJly+jGvav1883BvpBmAfCiqZjJx5GuOhp
cKqz0TaCMBgCWtYiRfczMqvfkaeM8SUUJFI46e+6bL2+5kS8I6OZsF6QLadk6ABH
Mi/fCNcKYIlm4VVrVCn+LaWYGhWjAbmQYFSkpOKvhHF++eccj2cmFZwlvYDaoh5E
CNO3dHjxZYQhubxwNVXO/hpIX1ZGKkJlVrWGQNzrKu9e0R/FZVc6R13mXCM66di5
aFPd95PPcF0CFjsC/pZEOv/yI2PsXm6uf/qfZAWLp6+nwVRLz6cRKeemRAuRh2K3
si3q2Yp5fl7AMi5sTI765OkFvQTJjCKdYp9s8mKkXLZf07kRoUCffChAYGzhO6Id
WkfIbQvO5maRU6e789OPZx7mVCCwII7WIgNlKvG4F/Rv5dY6kfT/lOIPbP1M0rLi
urojv92i/6eX8cHYbPa6QFn0Ghxv5AHvMU/uJJA1M5QDrl1m888u/w4J/jsrf8Pd
LhV+l9WN0sXrnMKEJfJnhbhkBLtmxfIMTTT8obj9dmaPD8Xob2LPicq5ksB+dfbH
Bo5LN/ELaTMfv7pOq6LkGAYpWrAbS/yZPUs3WoX7iAO1MEWcb3urH3Dbndb2YR9p
WoklYIicGjV7Mzq0UG0nqzqgz/IhUe1TFjiOqvFExWU5uoSi3n72X/5CLmtlnqtQ
3h5VjV3cqMYxQq6Zj9qtYbeZzPoejy/kmEfygp43nr4GRqC3/Sv6lEmEoHdl6/HO
qkdLt7NrYEcE02HnYed9RT6jGHAWrGbmmEEacu2wj4Pxnt6DuIbzgc5+2Sd6h4tF
s/E3150GhiF7ZXeBQrrUnCOVwAKlaBWD0vlUl6OrczvP2NkXPCf26Pz/IlzesmX6
Hx419ZKdK0H0p7vD5Zcxm9UW+0r/BC+hz5OuGzGU9+5KmBSQyx798FfYKTr92ifr
dABk3tkIDAbreo3cNZBKMwKmPnjWXC8l3XdOKpu+VQJygwbHPpulOW76FlHqivQC
hZ06p7cdf1rfJGTF+PLMwIUXcF9VGCBLBhgfU51Ttz12XzJasrnEm5S+lTf7KPup
dDGn5HQt12PYA48fvsdTRdEAaWqLDPUfpsr7uKLMnA29VKUYSU5E78uPyDGFqfAK
XeIBjy5SwMf7LikD5nWeIqr/eUD8AonvxrEjpr3nf2nEHlTqJqXoJr9dt4kzlSI+
6xyPanLe+iCC0zuQKlAbAaN8DKeznJNUbOIKAoI5I5Y6NrbxFUgm5KxCvDT9+Uki
tJH4lSbXPLJqeEfx8W0R0AfAJL4qv/AKwu9QlxguvxbGiYtEE1f3UlxTEIQjdDET
MighgDGiA5/2nRoWhSzk8/zkRm8c+p8tCtxyNT2S2tATGmlqB3G0Bui2UPx+ayBy
W891qV7OFIC7FxL0KUvdtTLCTHhmBB8oOS5ErDfYZNBA1plHbVCkiVbRwHsXb1xS
6/6c0TNjFHa2FRdIAB9vdO2VZN9aHL1HzEZo4RZY8EhlGFOo6+nwGX1IiLut943o
oMf6QqEhkk23iZ8BllvtFKTKFlh4dDCNu5tKHrdcS/ulz+2YqKcLY4Y8F+SxI4GZ
lsbkFRVPABY3fnzwd453pKHpaJe7T6PAJ9gWd77e0IgtJWFFQbDez+sf9mrZT96k
zYLXqi6nJ3uNaAfj7J5hdCh13UCHmrkeV8NjPbS63zoEigsgM03XNIcxV3hrDD+a
1eLsF2deOzfD4MndOlKtBGFq+FLGz9UWXLXrglNL52rx1BBsXeis9BPoXtYfCJFE
WExL8HMrcK5WOz5PdvhYien7HEJ/nwaHDQE99HnoW+hpkmBaAoR+iutJ2//obsJ+
Z1u4VM8QndqnQIOIOLMKt/9H/LZfVjbpRvn0uwQ3fX3ahc44SkMdGyhYakxpx9pM
TQLjokJwJRc0W7p6CRhWshHV0UgDPUZa0ltVeByl2+BNbPOi8lObWWuvp7VwxYB/
cUi3Sqpmh4bDLG3/5g/OpIgpcF3Ytu+dZuZFPWlwTri2PDWA1zLUZc6Toseoy1pV
0rRo+KztDuFhOvYz6hTUx3FKpn3UXFSPNFjQlBbf3REQkfQ/uIitbr9iaymAPDPz
lqCX0zsvqZwSBo8XrZuNsPUYVxZrLMLBglvi1kyFcXl9W3ZEM9naKLg3nkeAPetd
m8mml+lcw9D2NUuY/dwK32BlyRMmNPcvPjk5hauZXdZRifmlsvCKcx8WWUnXOlp/
o2zptL5yU97di+57ZWXKNMtBkZFFmC3uc1XX2NSZI3TURqfJ9AhXhhcL2F6Meayf
4mT7Izv1WHzSfIy4M9QWknTifUq0s4DhLrJ1CwM4jcQOQAIR41C55/2k1vq19RZq
s82xPttvVCq341RrVnM9cIVJG2tbG0bBKWwSKFym390LJNaR864aHzn0ZKt7Hfj3
nAKIbNZeudUBBcYmjvPqv0JrUyRkl4cxp7DEbd+f7IZqkYqtmnH27JxydX2lEMAI
8uR+2kuVkC1WBjse6Chsn4LoWkeKUit0/X8Wc7yqhBdllzjRNJ9fxlA5ob9AUyLQ
3AS2TWYXiit4uKyjsCfQwWKOqYoI5O0Qr4Fa/rkX4g/1PZ3O0sPLEBsPV2/9sv40
yPY68pogTCD5AQ+iIJwjnRpm0FPdrNJZ7hvW3dmXSN+rQ5cKW+3ldaH8BtI8hmXN
oOp+OphyajOuCjJ8dcmsU8RDWIR24aDUEVjSP4KAlUoWFokldIWzP3trQU0qRROe
Vdu+PVRRHGvV6wA0iLffdaSMIBFVUn0WK/CV59bEUusunjRLHjmfjAHoHQfUc2Ze
q9md9u0hamkyb6HCqbmTiFBJXHEVL0ZyAThx2TQyAt6oZg94bIShj9ZqXAWrc6ON
S73ylfmu842qd3vtp8nrGEnA8XMCrnB/A1sfpbeVcd4hu3iijEWEOyNzZ8JrTYFy
WUHT0zW0aKGpo39+fKQGH2Uspknmbg/fPJ8UY/2Jm5VltYBZ637aDQ9ySUnRGuV7
kQ62bpyoG9P4p1MXe0yQeaAX+6K2eQmUo0uWx0tIY0+/W3Tb+3xLUrAc+O0KuHzR
oVLT1mxgl/HLk0ccXCJV4BZliWKDw4phbfN6s5kehbLwVhiQDtMzeCRkslNbd546
x/ZXnJ35Dze9YP5aZpiGcT3L776XqiXfiVUQigbA5V05+JJLeF8sLuPQn0Q3Sicf
lBkPydvjY97Le2Q9FrTwKq4gjFoClEDfiJh2eVcLJM/s4/DokTTWTy7BvqiIiiQO
TV7b6a1yucfojDB1K8iTaUYnPL7VMRKTUrAG3YFCVoep0VFquRDWBGbZh7LHX9SO
Xxtph3rSqi4JD0y6epmCpT2h08V13VXnoO+31Nm9GhpJdb3J8lxG6VwYACARb15A
SrPSTytJoYNVmNdGm8DXEgCYMS1jkUTB5Jc+eD8NptZHV961ZQUql+DTpG3iM1Sy
WpuLYfltClvd/YA/YD51oJN/J0i8g6SW6gJ1uySZv593dDPN5vj18+Z5YOsl0zZO
t4gsy2uSR+kwFIYvxDd4wpB0rQTlzNh8HYuSOmXwj2Q+siWGKwR6NQs+4jqorlsC
k6kzoRcQ/QS4VO5hXa6pUsZWGhl+vh1UmfTqlaIdQTrwDbuZ4nbh/Dj0LxUWgbyH
FAlmN/kdLT0U8AJNs9CcSyvzvPf2ztVTQqqxJW1B7trjofbifYWipmLAyO1xan44
9EwEHvqDgoSekWuITg06rVIK5fH2IFPmAkxxrnL6bi2IQrBZjpHdu3ROcXTEHR32
O7OoEmHdoC5eEcChgBJBLzTnUW1wqw6qg1LIP7yj+h/JzbtGS1JtSi+lLaIoQsJY
sm9SejXtS41vz/EMkAbbXLXY8ST6iCznTFtmvJmVBecv74dbilBjxL4hx3U+STHL
hCRV0NxVcUdlYZv6vfCE1CH7hGmjvRd9c0IarRfim1E7KLSymGXs33N+U/QrHfLU
wURbp6aIsTAxvn6zuPIatKPvRJiww1Dhdk4gI7N64wePTJ+/38jsrRGHf61pBiFB
IlQ9A+pAR6a0S5OzcXYyWaqfy0/Yr/7Z3CbVNvjVWIncagSK434viLxREmQJ8H8c
6i4QAIPx9wvX4CKtnVaGKZneWut43EQzcwz50K5QwzZ2iZSicy5GWWY7E7WH/MnO
g8AviMc9YX+dWQLpDR9LFO1UfYSYJAWpsVl4l/cp6w7JW/ogs6JQWNgwDPSDLjYl
KqMbrEaaQXYZrBC4CcakOq0bPGRcB8ULVEsxwHZDwzHxLPcawbqCL44pVranatg9
xuxjheo+RObJ5J9cdkfJAeCTCUaTYsdDNnirVOReq9tQzgo/d0Vsb1aavL2UR8wf
VLlgIhQo0QInWVHb9W6W9dVMFNLNTRmd4M7VPYzinl6ojx+O8yuiQx6leZPdHdnx
FGczjR33SpBrWIO4Ogc2VszeWfbKYdKyoGwyqPpef4jZPH6fY9YR42+YlqOhek6X
Svd9W4MsSIu4oK9e/tFrpGHVfWBndW3nKa22WtAKvJ8kLEHyq+hKiuk8wHkfj5qR
m/PzJLMn49FX/9pPd0pcSqkFSm6EZKelndx89VhZIgYTeSbpRy2200/yTXloyezz
KRO35wzXs711UGZITTRR9DWZHkJurYZhJpxkN9RZ6Wk1wj3csWnazuXAYxfcI4zS
7xhT1R+IBtzV7TCmRDcN3tsP3lL9O7OJf0qc7izTXcdqUjVdT3I0N5NyVCzTI9jD
92wjEvVeYOzR23G4McX2YA/GY3D9xortRdJbxR969xYqP1Q0U1rp6jyVcVN70xLy
fzZ4+DOgUogql9C6BYbzolU2x18Ps/0AdnRuWJXILWzHvTdtZ47MAVH8wPHzxnWx
T/anIa5hzPo6fIJFrtvXiC/FJs9y0kcENJMAzwZg6kmib8OirU2tJT8pI6vFu5AX
JnwAgKhSvgb74ff7z6hYKTBUXjXajgF1EknZFHGVG5GFD9nJj1H1Uj3BbfPrP565
A6Wh7kY8metLhCHl1R1v6sbTAuiDSkHYN7b6EH5dBwlJfHb8zZ3HFyFQ2qAL+Psz
JcmqJ6sxbZFO+d0O33BgFuAnf9zaiavEceNxgZ3i+4Nuq9hOzEoQOwiaCl9iWuwN
UbHwoNgtUenitfWroFIvsre8HK606sqrwANbBO25iT+qrsZB+31s7r1m6GkAgh6k
bjbZWRXdf/CSpZ/irIdUGGs2ORUg/g8+Oafo60XuBnjn+qnK+2BblVmg+F+6mt3J
6bTyuAIQMGNq1bhYVNwLmbz/HHHtyGaLEuDwFMQw+wbLytwzChoBC5ZbsIgiC1zm
3YJxuQK3/kncM6GsdyxdBDFCcq0FC9TC0wh+DRj8BtJqO1gOBEBSGt04U8WxlsWr
gBVayd/t74aoQ8VJQ9tW+FAymaePqm5djMe/2AlVz9lau4EGgbd/KpcujxFu1Uda
XNO+JP4A98XpCN0uzKP3uC/F8xZSBAleKYATSYnJ3SQHAgyMBHZOwswxbqqR8nvg
rIeevZUbUzt5RMbm2Sy6xwU9bbzyk6CC4TqF7qjxsnImTn54ruBdtrEtB92xXUJk
sbzD95v5Xrc1UtVvLMhgP9+7O/IqpbKdjMIebR+c3DgFNO64V5jyAK7jP85NjBvv
ao0CgP31B25T9BOKgED+ADMv6XPU3SynHmJ80hPd4KI6xurLSEcg2XE7kmXAr6F8
4MyZMZnGshf+79ZiuxzELs/eWNGd1ThJRe9EbTlvQhTcivqirQRu/Ppj58Yxo4Bj
FUxbyXzQh9Mfn36dMuAfjr6a3eiBIK5+HTedIaKOPiwWpLRQTwB6ii8+F9WGmC+E
wu8brdo5NLlSozo3PW3rK4JUBq2XE/T3vEf6LWJRFf8pq9c7ekMzHdIwu4QU3MG/
SLV22eXKbqHDDl3jEjM0OMH6fI5cfWQlPmwkQI07nV8TBF6bvVtH8lRWe8z6W/y5
gs51rTb9F6Ic1niQ9UbCNP+X6E/ZwHoUJZo36S2fgYL+v0cXTMo8tlBP66WvtdSF
f9GZJ5GBl/uAyya2c73Fh2ENWBPO1e889n7XJt/KCdNiZMdOEivbBifu/VNLA2AM
NFlNm4/JYjSYYwBgYJyJl3BuQnziuhBAd4wo4ErwiqtCO55JxR+rars6/8S450QA
nXs1IPs4IP8RPVy/bJVcqz1H8XqVF7U3JhAHFLIvYFDCUOAAzOc5YhDZmIL42pIu
erdWis0qdHvnxkwKaHlOvVmlu6QV+lqoFrr7TIq/W0pJzbX80y2I6sUSE8XHPWp/
sxPNg7rB7D/fNh1Hz6xrqrfR64AJF3BiqPM2NfCxggsece42d7UtnaOgCIlvHUjm
7J8msRbbZgBersXdEVltWGQmrueSjjmwyEVb7md+09GRpKJnBFzzaiZYdg8TQcjM
4l2lldAcfiA+ddOV8Xs+1oCtHOdrDmRUgFAuWpUsL5sBLGa13FoLWafYBJUKWu6i
QcSrm/8Dg1dAcOcHFY8mRWuhKRiXgEA6WDixBiUprcsDfGNiXM0MJI8h7122GMyR
hTosQzQ8ovirXeYPMOLUsYQS6kbnlYr7Ysm6Te9glrTVE1F67Jw9hzjHsDvHdDIT
fTpj5VYJocRhLxU5IdiXeGG3k62lRNAJwKhHfO/WY92zBWlbEeRH8Iz2d5KvZ81y
36M+CaMXdASRb8OjYn9LBSZBG1PLz5robzosQnkGCWJ2zPl1h2JMwlPQ9SvfImS6
wJ8Gv699GnF3jsBWICN+TYyZHFS/RBenF6gL8wbEZehHXQY7Lu8mgYmVi+cyKSFH
RBQU+w4unhEnMk8rbPuuDnZ6vc1VSGau4Nvn4rCpZdIjF08SqPZIf3SojuQPnXvJ
sVWqJt+bSP90qD7tQZzW7PXx6HL+4eJoA8XX0IgG8ypzWSBOUxRnQ1AwNeHveg3F
gJO+oCcS+L/vfMh//XvQG2URaf4EhXOlf/wS6hZPiHDwwTNp0WVP5PRBbORBVV5L
6NrUJNEn6sZjlyFzaQCFNphxdHk7U0Iup+dInwvQbPeW+Udg6cWYVPQGwtLB/nfs
t/x6vTuae4sqyxkvnLxY62M6fY58L9JVPP/zeZpjN6TSf4p3Qk6wL30JaSP4/8Rv
xdk07Mi96GHTcq7/6IzQT+Bz8jZYxKtXo9wdqipR3xuowW6+xlZZQEK1KpBHY9K3
d7/7oH/gOgZcal6kNJOw3Xi4GuHtSMPIww3qEmQ6DXptL/YgY3gegJGWfRgSljVI
4Q05my2es/06F+Vq8TnSXlgcLMGhKMs6OoY8tpcjZXTJGTDKEjwp6iM9tB1XUYGw
H8FhWZKRDsuDM0xN4Dtf/KcfFltljmvRkhlaPvsRRIaj3MTeYkzepUz10l4zq9cg
7ObjIz/eG4yOE8t4MkG0hSYrlICEGH7LWjrNlWcNHFAon/W7+P8UiIyAGM6CuxPd
s1ejjdtc2efQRFyhFAP34BkQYfAfItUEpyp5KPxoWBN6nOxw0Pw1tWH5Yzxg595g
6C4L4+x3w4pKboYdqop7f9MIPpCwjcKJ+Z6tjhYt3zU+tUhOUsgw0cDYJnPsbkLJ
CelBkJN8oHXGepXiy98EW90N2szYu/ObOqYWl91hBNuFU3Dn3CnZ2jcDfVjNBKBM
V2LVsTTW+wt1Cd0MKOlE8Kxi1Xr8PHX0zp8kf481sGW8QCA9L24VR3UXi3I3iSaE
0N/nJky5K388f8Prm5YMVHeB6gJMuqZopiLh9UymfwHOLD/Y3hPaZVccXaC68ffn
o+RJ4V+0sTpKTmZ7FLw/udG2JB6U52lxmBRcpKV91rKM5T/ZwlsMukvnj81ErtNR
OWiVbduXhiS5NwjHiPc1sOLxOLoqXa7zwpXFY/MV9b3ne+6UULW3oh4kFB0uXNQU
OKrfUXrbkIdxWAaIRiFJ4MorikBYST9tqSahXKCxylOehf3ArPADYrjnY67CuILS
YO1ETxHbKKa0xtJhGiNGI4ZTXaL+/gNu78dQ9a/KErUkwyB4jRsbvg/zmFGaVm2s
jjF9nsNrs/xw9JW5D6vQvns1IQgjpLqtLrndSCYvAmexxBoTbVPyjLy+iD0C5YKd
oDQqlwnjf9aSXE//CFWrfDSdnRRoBeXNbuGdduJJVifUQDCz39fvEVLulFlBJUwl
VXTeuXujlY2Kqw8BgMNqeqXR/WweokofYZV2rieJ0pcnK8zmYtM4EZWThe89IUuc
UfR3Hgt5BeD55BmaPHTTa9X6LopT5kAf4d3oqg8yuXWvidi1uiOBcOmdGUYpWoQz
BP8S6RkIefZ7YP/H1fSLaLSNemT4GwBSIwlAimbUnUZbqS6F5RvWlR5m3iqtnp+V
HCNSqWHo5dKIxgHm/Zak5eAaMqFYYt7Gh9Qu7iDCK5oEBrA0+X8lxD9frLbis7kw
Wsm5oZmptHOOFq8y28HAOIunUy0QM0ypuiWK5HUFseq8xy7rbrSDCdYTy5Ua8yXx
i7roXxJ6qhcKw+e1RgVQv8aFCm2JUCrl9TA6HZHlxh8sMh/EzMRXIvwOZbYdu/tl
UIzUR008psu5RxAbvlkLMK//QVie/O8bY3RFpELuxlKTzREjKp0WboR9xavKKZpr
MBUEA5wNg5AelDekZYU2xVITkRldA1588LabgUDI1b6cZDe9gxEBKW3QWnfDP98z
50jysbyrq6nBCxkgkGQoSCVixF5Zusb9yfKoqcGeNrUBdDe2Y2ICCzXUOwDR2x5F
4se0vVtlO1h4OpeYTWFH5I4+X1fd7S+qYbP2CQOMotYsgbsY4k5+wwlKWVYrsPFy
zIOmpBYt8IrlpmhzWetVDXaseZAQjUdxVlK9HyZK3AVryiBUFq6i5iEIchdE09Jg
CdLzJOQjm04qKiY+UVIkevLat+YLwlK5BghiyakeXjp8nHvScs4JdVCK+X0pg15i
iyed+lM4gvo21GSLSrsZXSNzktrbPwOk3CEzoQVSAjvVujgUOyFO8F7Ko+SngZiA
aYnTeUd9cK1eg5hMBskbEeq3i2tbFhqnYns5Dbx8+tB7NBuXvE7mEseRiJAo9MPt
O9YksUGUynxTLRuwtihE5LTDryOpMOZJAYJN0KzRr61al/e9U/GGV5DfY6Rvi3EM
7uUSjdT097Ihmt6kl4iZUqHHO+YMbq3FFz0uJVLGDkNP9lz37TLmMjJkpv0/NzxC
qvE2FRyg+W1W1nLbzj075PgEKbVDGFdnjjn484gGrX+jJGJG/PNBp3h+tpNGr+n2
gik03uTu5AI80qyG5CAtUTB2V4r1DnG+ykFdLwX9RJ36nrCHdF5YAk0yu92zu8Gy
JV5+SW8kjpCRI4WJvDAEkSOhSPMIW9+VgNX9T8IGUMviiZ2+R+VwjguIXp6tHMhg
mIYylVTCqLm8t9zLW+ZQq41M55ADkQQTP5FRp5vBPnj93CexsKQNGSk2En3Nnd60
y/qLzL/CrRq0KZCW2OaTwMFYw2V5r1Gp9aZgDbXj3vTmRrzwDP1pKVpFyQERtqc/
eP9K58gt5Tnjl3EPVlz8zc7d+L9jU9/g5ZRyvQ8z/FjquQl/1MKO8gPL6NTNWVf2
FbyX8nsWj4yn3Zu3y86N9kg6C/byCwQpcO/Roqr5u20utESpAYRipM1sIoxXcoqH
JkEv9eXStD8/95k+DPgaAfTckXzldr+BNvLY25XHtWVb+3T3OFPqlCdTcoK7UZcR
Aoq1pX6TqDCBbFDngnzyvIbOb8PgpANqG2/WCDpHKKGdDrSs/F89TIaAx8qm0n5B
2wxHoJABdDCSqewzKlWx2DoeNFXeayRfOU3xAeTSGVNYwVqpAXWSTslrqM+dhnxE
EOMQ/uE+iaqnSzqAmByyBdrHUp53eo7SHKQnGIRNO9TczqULN0THDsDXHczPY0I2
7K6kwgm+/9G9wz4tMwmGntgMzbsRHenIMlM4CkerKyirkBbRtK/k7M5GwD6yBUwj
8lTe/OffAwGtx/jdLNaolGUsxYbZl209M5Bi72mt5558aoa8T4s68pnseLoMms4T
dj5XLC3uFlq8Kag6vob0HuPq57hJmK63ujnUz0y0k8RN2lRuUNfCSGGuyE4uCIFC
9tIRjXYRnSA1IhlJPQHAY4T1WehCo3GdJb5lnpJAnH8gWw1FqQ2dnxNPmQ+TECfC
9ZsJGVjV5Gxb1ONsIrmZ0C6MSe1BOrfqYN4wPW21Rp4KZQulmX7OdBvFriIEZtl2
+IVqJk5xW2UkWYsIRyhKrJlyUKnMmrgJMAFv1GVkyTN+TvYzNE/rG8HrmOUL+cEZ
JYEzlJbrKH4jCXw1NI5zmZ6mHcHpX0Mlz+0rxloNwtToFmXlz0TQurLSsmD9v8ld
BtqBJXQ7ILUl4CRhuIbItmyjonzvhqDDo6jsEf+rUPJmwnK1trQ6ZF4BOThLhdHJ
ZWx6IyoOCvLek1OqMtpO15LdfIyxBuWU6NDR+5hFoav35CyynaYYk/GceKCPdXGO
74JlZFisSgJAsHI0bK9guc8p1vPYwXcm2/uiKbJ97oDB5nJDvrV0DDpA+rE2JooJ
TOlPTW7wvM8C+xKmROEH/Duc+tvsCWui+7T7sdiQrpAORA2m7ABtb0TyIIlntesr
UjBkqSFcklSKTG3wQAFLhIv+gYdVndpNePkXT85FVPdb08/e24hM4fiqkzqHC95j
KznWI8DMZ44U9X7CO1FHnMyZ3LtZKcZ6I5Met9FNlpOgkAFLab+ou+nKfDJSq85K
oEJUhYI0pcVCd76e3njeubOstDiHZkRAlQBX2GTk+pWbI7goDXVuloUY7Z7tbC+O
0S8C/b7YmZeiRiL5WdfMpTTMFsN5d/U/xvVAv8viJdKQO/wgblDMn9Z3uIde1pjK
/B7vng/WZm9FZLvL/xjLNdtYpYhqYfYkbVY4y9v4r1YEG9+gj3N2+zBJQOgQths6
WruaIKcjjiPzj92bNXzvuzMbyR/7juWHsYkaF4kwwpveiw2zrAHz3kLRCdvXTE+t
qT1sXz+f5jL1a8YJ51E0QloCBT9MCOuH9muQrhDErYcfezjzqFzplaEGCzsqCPBF
ll9XmBMvl/PFSf9sb24kAHn6UCQN91PTjdGstClx2SDyo+0M2HtmHZVS9U+Naz5J
9SnYDH4OouIu/U9X+m85Gq8HXvuy/gNc7cOcfcWS+dElyLJOlYOpyikk5N6xc24n
cL6kgVfeKNj+hT0rx2XXuaDn/NDaT2Muat8v2yUJUqScI/qZ/kAvLC+UP7oR7Wbp
GciMjiQboDkRaDB8WflkT/WOYg9IFBnvcSEOxYFAILAwDqQwjcrlktv9sj+KHB1z
V+8sbv1uoA8M75GWY8Dekhd4QaV3wFtcsiAeOucF76H19I+EusyMSSPOTV2+uCie
lFDV79ejMCzHGT8nMHzYkFSHkptvn2gsXEMt4QNRivZtQIn6RAMb0uWmZCbIBPsI
trAWb8nZEk3bF+dObpYI9DhjuId+NYC53NntMmaAAmGeVlL34rm0KZ2BQYwlpynr
yGFi07NbYIx0fQ2e095xq2wXsccIJ4CUBz/tY1fw90CyIuWXr7FGNqbMb73ZoAXT
Fin7fZe7WDVkeBXInlcS8zu73+foNCV5e3qv4m9PilAyvk/+8Zmn/RwWL8FMnalE
jv5eoYz5ZwrdpToWbAkq4UPRcEoBMSffhqv6/zCilwbZIkZPf0yXmwn4iFrtO+TV
sSfpeiclvYej28XBntDm3F2gfQ/TW81mqzmJrR2iHyVrx4IrGdKgFPnv0D3yXo9h
CG6ZPk09cUiSZGWrHBcsfcyYjoGPr2bqdreRYY8U8p5IRgNx8rD+bqVvIF0zmYZA
RctUw5y909/i4Obbo9fi33ReX6KkvFOTdGX0jPPLBiZr3EI5d5NMk8pNRvqk3zrR
4J6IuowCgpbJ+G0iAp0yKzj1xmO+cIDhBpD17mTM6oxAmVRBCKVIhgQ0yoxSe7Zk
gaG6sF208bDXa/nPJ8RFJfLKv4EsdXadiH1VTfanX+MfJTaZb0O39HzH18StX4n2
ghRRH9Y9jFKfAA4lQV+LIBakBdm/KH6Y8DDQKlwAELVOksX0q1hDPgUzwyxtdm5G
yC08hl6yvXp/o0fABITzm5sHaImfZLYPPTAYXJxziHfXRXmS8SqCm3xFVEOgHnbS
qcpjbCpBxLkTfGKMghg/YjGuE2qSPMyr+JByf2DWp4TATX8PK2fdSIpvXhm4+WLd
mxMQVmSacIYYaIeK7D+Ir1p9y/sniMUXrwLZGxB1WPorqpQXs5OTz2GsjrQYXC8u
A7D+kRl5CCggVbs0hsf78dTcQDgz27xBF5XGz3Me4X4F7f9w/HVZ1NZTCCFuAr5U
minb+QI7fwu8qyZCaGayAQOeqec+fOtpcdIoJ3ECVQT2R582519RbZWFPdqS6+MY
IrKuqWrGjUoIKGjPmvtEnyYKrQktgWNLtjXH9izeDLCc81+82EPoyzjTELFYKB9Y
BKoycbbhHeS0D0IQyPoc6I52GMHe1r7TEMm78uwIvjT8qxND0w6P1ubaEiFLt4RN
mDz3tN41FzMvexgiI2DNcUfwUYyJFeGao4y9AIW5lk91P1uh4XiX57iynmu9FDHg
XDaOTYr6lLKxXrklURyVmJzlg7anSwiVfFzofwpqLcRXdQ1mJMMKUA0nSzFyyeO+
s/E83UVuRa9M3RqXsmjdaEy4ShhSrZf+71qnT//Q2Hb7Vxwjk3mtNgKRLv4UGxCk
dUYjtoq+2ar6F8hKKPHpSGICsUZVfreT6fAgLvyfDw0tAxPwoWs7fg9rkftsNecD
5zEQa1H/W12EnDiuiC9auVX720rSilqdb7ZiYBdHVhQU2fVBVD5Kbi4UL7BuKUlP
t31EBkun0GwJ95ZzEJxvEkUbMnh5cAZjAG8AZzd3NkVPeNMWA7lQp8WCoa2HqgkZ
uc1ForseRTb7FFgyw1u+4GHHwTi3/iqzHQM8kBFD++cJXkiii1O47MFxFJGdPFRO
ufjuLl1iAthRGTffpk1KMuHTde5HwyoM3dGT5AVhHOtRPMtJpUeJ3y1WzdAkQFBp
e3l+ho7VOpFh50exDpgjrsO85/cP4bSggTyzzfEbRyco2OvPX1xGpwfStdSJaYoQ
80Zhl6QTtdvh9xzTypIfP1K1zWrmhETcJ9h9VwY3vkdK9aabWgWx8kQwtZQZZbBu
N9Jiej/p7vR6eOjpGyTHu14akVItaqLht7Xkmxl9ZebstVEVi4fY2YIv388w42Vf
fwie+N+THHeCvQSHR7O0w4fTwwPazGQTsWssmFqjN+k5ZJJ4fr3LUOdPW1Fj6/Up
k77khQsx0RVj9sYI+L+nLBymJOwwzhPyGe+02Qho3wa9REfDfPsWHfLmkw97gkjK
jQlHeeNnk9qKyDTBBxu2ipggKoF8K8o50R+NCEJ+tD79vNyUeVMQ4dugvIn0qRdb
6+klDHzlmIJxC2pydHq+ORojMl9unqwryZzvdZ2Ln4/aQFkW8OdD0rpsoTS3cNvA
jZiOXWKsX9c8wUnBejtRb3PZlKhQaiEeci+xPc7Amsf9WDxsXgeX4K5N0PBhB9xx
7gPDDx3JHsO7PKEkG1lR/OwXZqbYvTRYH7gDbQxa1WIfUYg1o2vo1HzHgdNH9F7c
dThRlQ9dYvV/4FptsoKqCEWAwPbNYsKMRGXGJUSVjFeQ1yI9e0vs1AoJT4NQNw3G
Bhn+YtFWJmDM9R7JdHBpV+vQRDUkIZZpAomxCqUpEclfxg8xzwZ/dfaCTLcovh8d
gV8VqZXwya6cFhxziA/xT0MBafXwpZTTj+cMJ5ad1Kn0ShN+cF9+T3rmnmhlOiIc
q84yi4S8AIqEsY1qW/mGaQHidwCIhTni1KLmQD2aIPKaiIh0h5W3Xbz8G9ajEria
WHbAyFd4rPUjzXcr/8km2B+eq8af9sVmT3wPIYjDb8lHYY63FTGqGIFlxxxFxKgq
RzuuJJzonxcKa9ueWeO0OPT5DvutekQU1Zlx1udvV+dclVNfwLR6bjL9tBzFR82N
vm4uJJ8z4/YGtaL5icJ3i9NoA5nmD/aHObqEvm7b8XE8GLwD9I4z5s2rakzfUIHC
k43KjdTo35/R+Fny00PhJkFyhfaFhDaPQjI05cmQpyehUTJBu9Pzz/nLsrf11zTN
UQh25zSRaExSU4o5tsDYPvaa0ERovuQ7DjVP1AxiZMxg1uVc32u0cfBtQ2jGShb0
3WCKvOss6yXX1tepr16WTHBs5pfxoZaHR9VqadUOBsrfKynX3sBrbDt0SXTSMwHG
S1cARZrxfSpJ+JUsuDnaxgx64O5ohjMc0e0vCU5jlmJTCV3DMKbvS8nw70Z5X1sd
h77Y7pY6I6jckeqbQOyvMjR8rGhS55ZhaWIV/Z5cK6ZwMnKDGFP+T6YQ7y1FoZlY
sMrPnG47IXhUwtUawkuZJwNS2BXYK2Y2SjTxltKG9qU6bvoUYkYwxP22HFaMEG08
q2MVh5HhgyNuQS/YjtnCIIrZIzRy5rNXjZUlbbZFv2btDop8Zxu5xpksBKiRTvSs
57lScZsQ8eJe56Pm3mnqRWlJjnTKV/GGGXUt0dgG3EWlTmlJ0pgsnnhJJGKhPoQB
BVGNkr+thAgxYivzdjEuaID63wDSdwF07kJsTmB1nFyviJbqbkm94CPOMlykIWRc
BQNFF9hEPWdIlv/hiUtJY1ylsvQgUubpBfMXbvnantyUX8ZNuMKnC8XbYnHiVZZg
MhfkCaVOpUH5kH9ixvEksTApAwG6VZNz4GmmetPlhYkTOOiRG+E/X0rvvzPBcYNl
3ghWMchI6GoTJhERymugUFEljKyJsEJ6uZwPgTq425Qcw2w7WBjRC3S89Z0XbAs9
sVO87f//1rrJgygPEHM4sZ+QlmnCos2cFx9IOpRNXPmNZjU2tEltflmjl1UdNjdZ
VuVjW+kiZWj0CxibxUXToTGZJFGyS5eo76r5BblhOgkA0bNlwy9OxOx7zxTomjxF
HV+HJU7lne+VdRSWv8FguSXRxYUrLzsqbRFQkSzu5jxoJCoE4a5QqLFu4QjxAp7n
aZpNczRSNexzlMA1baekjX21JsLSOJy2Kvk1JW2CvaEd3gjfB8Z0QioPQYFENLGk
CtvHfeMs6pr2nUuRAiCkbPaHpU6Ymy5Na4xHawzDKzKWB41h1/OHKXZN8nX6MogD
efNYbxlVyTrQfFrwO+PYz6hUAoHn8NZrgy63uQE48TyuRxIGp3QQc/DtJ7LPAFca
UAbbUxFlNJv/o0+KqxWx0WkJ9fyl0miS2k+E1rQn5TLO3Q9LThpBUcc1MTuZdIVN
9IYNSDrm5g8REzGXutjYbfHKyDuFzCDP5PclGoBa8EWZPEQYiwM3Kbe5HwYws/tS
aZpgpnThDqAHJ89iDqrPQyM3C835svx3pYGf4adBksIctRdkcOHzRXYACDHSee+Z
FWKa1EEwl5XlA6qLuUqTjFP2ZibkHjPReoF0iEn/IyVGNxu9s62JtRpLSxGwNqJP
ze8oQ3xHuwYw19Yc01J/qfT+cUw5ZGD1nw2ekZz3Lxo4B3PqQV4mj4xh1/3xlhm6
tni1Ok1g0shu82qWaZsKLVYwPrEtnjQkv6yJcWZehy4EeANiw3PnF/1pj4GnuziC
3poOfjz1VXCSt9KAJaPyp10gEe0P6WsjqjxK/OWmgFGA8wk1NNzG3ERKorJylo9h
dEJ6y6FtKADAJnt+GS47UqFbEoeYaCGgG/9lvS2KMWTRNTtQs+uhTJBXxpLgxKE6
GRNJkZ3/+MBNghAvrVUDBerAmVhtwLy/tHHEMrbAB2zAS51SELwm6LaY+C0zCvzX
qyNBqfWp+ltwZnR5a6KypZO0GCvlhcMiS+4qOmVj3+gN8bxMJv6wxm/B3DMdtcTS
fS2zgM+QNL6/gMUUfo5DwK8kIjTjCUYejb0navuiwQ1lZLOMA3ceaHuHjbRWymz1
j3bh737vhEF62mRVhl3wutJV6YL5MrWng8T48Pet35TRZ1fnLor3ofaVc3hT6iV4
0fl0SH4TkaT60oGAUhm/a/vnAHdUJk9Fs2f74lbzW0QBKxf0kibETWo3vosfJ8t4
6WJz+LxwonoJnN3S+TU/EADF0Vq7Hr535zRAyH+EM7NJ+q+9Vlu5q0IGpfwLgM2c
Q2C9Wp/2H8/l2gRPhXonf3Ue4ygPwYIZ82Z6xRTj0tGCtIlLOREA86VpiOgCIGK5
YN9IIFe03fJ/9v5e9w9z6QYm2LtA5qWL73/PewYul8rv5aPTOyF2lfH5Bc6wdRFr
fBu/pzurwSMdaOOhqm3CA+Ny4YlvbRdOeHb45Oy2V48JR3DHw5RGN3kwfXzs46KY
iv56k0Yf+UjK249nnJ5DNew33jxlUX8rGHymRnnzvGLKhurBqf33XTgyQUuMcc/s
WhnuGVqPogVvj2be31BxEYKTzPgmHrFYElkyFjh+vxos4ZFhYqRzqS2ZOxtLu5HW
Lox+8El+GVIXIJju/7D2q+AZkcfO3Fm8nejU/VZkYoIxjsQyO2wqu3RXBpVHlDmK
C08tpXhYkRyP05SFZHlQ2y9NJ7VQ5Z7Z/RDiQKxR+Mav5u3r8eKqtbeUjEYjK3u2
j2cS5gXEWrTXjp95XlJQPyJh3P0dBQylDxnCGNDuSNERcANRDX6aMKBjyls6W3t6
yZrKnw9ouXoIRG7oiEEpONAn/X5C0vbmM84R094lGC1pdAL3F7PJpuWW8TfASgYU
CpHMq8ewRbx9yuthhgj0Gozlpr/j6Tnv1jMh7vJEHJvCK61GRiulRsGia3l21xBm
mJyfd7cu4TmDnpjg0bL0jCkMCdG7zvsQ6uDq/m9rvIGBnIg1cDcr75ABIx26OUUI
PZrH6rO0XoCEQKyS+wiWmy0n0vF/4dw92ZrhQ25e+L4hOTQeSQa8bBz/zPsdj41Y
lQfSoFZuimJMXkXsBV7kkl0DXtzq6R0f24M49NsAa2Hdzi5iLPAwsgtN/Euew8H2
WMINDOXXAsq4+nRK0zpGYgZ4EFCdAj+5uG5q/K8II3omxOFpyI1oXvL2WDzVgSFF
bniPYahuy4qFaTkQESky4BZRksNcHYA69JF2nP51gvBJ27XzIjYNfgwq5EuGenMh
yONfMOtw74N0VphgKoKb3BwzVOYgi7v71XBqOxEmy71guNrvUfhPCbg95Tm9xYaz
YTaqLUd3aBA1YYUu828xxrTNy7LjQbg1anUkTFzZVyqdxs2XVq2MmrTfgI++RTgy
h4KEt+kj+uvou1/wI6Ppn/i6fi+A6EcccLO0bZI2ruJNnPyihab1x8eRo5uzrfii
2zju01HTUukRxisDJh+b8dBmn6kTt4ztjK+toaWAjNrHW6VnPS4ffa4dimx9e41J
4jBq0x4GAKu9HLTqXh55xcAFBtb/zXU2h7mDbfYldwAqVLnA8nkvGvw6U8nUXZGH
nn40eGqfp3Azr8myc1SSZtwzpGTod2UzM+AAXUn/fc4z3DHlqkD+Fd7gBQyaxYpH
kD8hzR8Wo6h1101U8vPmyPdOolMUWs3iVgqXB81NWcYRph5uPo5zat00KnPuHQRw
SkTYnA1/fmzqzbzLuoyxFv0ytGP7TmgSFzs5W6NrM4E6L/d4LE5CsH39ObqP8BdS
F2i/MUw/KbkNNTGqNKCjQV4p9hZKrlcHFBJSpFjFQu/ILhiLoTeJH4IejKaHXkFI
JB4dQwXV4+iadneX1roXlT15ZCwFTCZp8zpQPVjbURmcKOA6pxCqFgQxvP3zpyNP
MEAaGqNCy6G5R5axcggGC5Iaj+TKdo86ec7znw4E84b4WprxDxm2sscCTKzPZWvB
wKip2a/ln4ud/FxMOGywKkZp2PwlW/07PQjbdpHfUDWZjRzjBczUQ6k44HAWqatr
NbsZjFFCvF0gTE8fyJ5sIQ8H02GsAgaVzHi89Uclx/HfRy72RiuIFjXYWOrGcYFj
xAb7NsxdiOHXW4WFNKzrCeCPsKp2/EZ6MwTrpv7sNB7Fd2qzNozkJ8Jyu74ovdKk
EegVs/ESAv6BAQYMnJwcqiPI8F/JfAFDfYlj2Z5jIjxsvlFJFhAjIelbGj81xzjD
9MBkVVWfRDlSCUBBCUIZxRZACSO2p+Qz1nuRKlabeQ6Ru+jgs2Q7EWuxaFgl4xnm
tiWNVS7wRD7ZvgGEKANSt7ebaNO9x0KAQyx5I7lWy6EPxg3mBURCOIGMmtMuVFDu
ukINmjysINiki37ge6KMnxWo+CIGd0Kx0TUDLfN+BZ8UqpV0a49TiGMZLM7wjPkw
zmi87bAAwvwBnXqSKlaQc4aA8QYcwjr+i27rLcR5wYbGrilte1qznSWV/XF4Ro+m
Vp7tL7BitGvzvaAtAqNGKcbn6s2hOlZSlG3W8WHtBqUATTBhf0GD9pl4BWxoylqr
rX84/wIf6Ck0+4g7GBUFXSMiGrTAQi8IUhNzl8dFLr1FhOyaOuaVmM5b++jhRp5A
YkrwGSVwD3h3kK3Fx73p7Io00J3DUGOyhB1RTQgguvnEIhoWZphFNmsdUTt2CVGY
ok7tYbNWDcEodRbH8x6CYJPLS87V0iHA98wsO1Ek7dQg6qOSp67pufpxruZKkqmk
Kzy9xjpihZO4dLT97HNGcKBB96JOPiHWscBUSkLH8788Uf9WD4/WbZm3cDr+EVri
AwWA6MeMZmM88NgWYf5QApPMOdHg3eqp8LF78gQKNARvtkZqX1VDuQR2oRXAKv4g
ExIygO/txjsW4k9H/JZz/cxdKLckLR2C/Lz1gPk3NMRXlKXwzbMWmwdLvovZcX8C
6TscQIM/iN85uSN2u1UwKHtAKB/a8fk6b8ZFqDxrFuksUzHlIi6DqTm9Sh8RrQIW
ybVK9n458ht4FTKOqnohM3zsx24YxwDLeuIKFwUeFrSUQHTsdJrtVp4YnzwsdSLz
x37TRurK3n/ypD/NdU/T3yY6dSVrAvmmGjF0fAK6S7A26Z4Iw3akDxYGddfnWOY/
IBZtyw+5WiNj1cF0Ex0UUSybZXBwbRCZXi+bWx4RLmydq7sz6nIv1ELv0q7UW4y2
WX3qW4aZ1EPHv06lgjT1HedFxziETUOdt/SKs8Z4FvuPVUQ59foa52Ki0oxAl7O5
EHI3azJwuvmeg5DAEn3zlw3etjksTCifmWkUMjnmSPvB7aSxRTwRFKzPbVQ3XBxp
X2w5Rgl1EWIGl/MRAi4ADfaZjELmdSkGzG60oAUSG0/mXHY2aiEvC5PLi9FhLyv7
Zx9bd6mLorxtX5yfBt1QlgA35wT2Eq/cppPxOHrRZf4EBhxgMMtCgWLUBgaRgayD
uW3s94gRquOo2s6cRDu/ePGQfo8lTt8K7OyYW70m4S8Th+tM9DA05W/UdqTSY0EB
as7tiq0coyZWxesA0Bp0LHtslEOundVlUJbjJYtmfFTBVKXQ/Ya+XeJMy1ovUHo6
qLr/UlnrJ/BgkcXcRE0r0PUzTspANm1ZYXE3bGvO2d0INAZw/sK/BnXHnUvEzUVL
+jaRAmEyTLSa85nmkMuxnyY20rOggF5FDqd1fv8ZQeWt87PZgubAi87FXLUHRY+y
XywmNCI8/33fZKqon/WQykBOFuWReslRHe4e8an5CagR9ZKmx3BT8FZvMyhfg3vE
yK5T4EEBlc/+/tVCZER8hOlpSOK63JibO6lJib9XzG/0OpaY3WBq2+QkNbFazwLI
7NeRQYSBRIzGix13DWloTPpgCdrJtar3BcNlHukCrcguRfqDaJ2LXYjh9K0rW7Ig
TGgKpfWciBQmAce4Xj6Qpw3pKpScERDcMXejWqyXptdQZOhfEc6BbkRXFCyfzJtC
jl8R17Ttr787xHK2vqJ243VwhMbyNHXEjb6vFdGbUrjfScEJrojGwrAqN+VJ2RNE
VSc9T4VZECBpYmPMUQmj88aD0HxzYLV1oRGwn+jfgdmULudw7pumIH1SV//LkWRP
LiU9qi4UQUw8s6xK+GaX2iOWt+wL8tpT9hJlKxT/mI8UJEASogiOe0OdomuaoRCi
TgvtM1fwfExErYKwx6K6fTHBLxJQhG+fnsNxWf2lJqsJMefY90yhU7s2kDLEQnWc
xq4UqZgmSIiLJnODXaXOxf9tNMjbNKdBLqYYJM4oOAGi3qWTIXEDaHuOBYhwpNQj
EpRJNxs6158jAcefplXiLBZDoMDGCAhXht030KwVrc/wjFrVjoAi/U/CfACdNg3Z
LosTSJq730M3YGm58LMh2cWd96q+wLTFoZfOhV0OFmS7nSsKNM+5h1eDIN1BcP2y
YSjZAYkgGMdskl7f5MuFZZTIjxT+r8xDti+ieYuFIXhdmamGo5CSEakfWXsN1f4j
OLCvQ7jhNrFRjGE1klgRJ2G0YT16wDcL3qR9uJMesxs/Bp3f6vZqiKKSeiPSrK9A
gi1Bje09XyUxwJc5DjKTLFCi+x3EWBZK3v5ETkb3Kp0W/v7RNy+RSa5aPTd8RaF5
exDNiCWoE0kYGhk4dqN5t/rNRzb9xWIFdIxXo2XsEI42w+c31xe95nNTRZ71K0rn
JZjvv9Bq67/3dHfkuGLWsR/+gq2p6XTNFu2m3NwglgMv84rkW/cSd+lZS7viT3YR
1V4uk/4R299nEYZXHTMWK64iJA79yjhDBjuYiNvo6TIoWoIoQUhwgsiAAk8DsWvI
lVIiia6MPweL1OBNXZqRA2N7Wc2Ot8Kyehg9dEFM6Hx9W3GSvBil84ZNkbQBfqCl
HQA+V8DOpC1oUJMzLJDNFihaJZqaOqM2JCDyhQ4wj2PMxqGyHezDoz+Zxm/Zsocm
zdCRpEYVrIhavp2M8yCgtsr005ssH/npmaowsWoFk1h0ysbXCNBVQ+1UHNsUck1z
w5zjirg8hDuI3DYd8c52LY6Xpo3WL0Y8OS3ZpH+wikLHriG/Q7ASfrS21POAgQBE
HMRNVuwjcoXSIH/hAUeWI/uqp+zCCQQ+Ycbyhrt3FAhQj6sdxbWQkR9iYx4PdaBO
kwp/oqTNCJISzl58dLVG8nczTiwCXfavsD+QrZFmTcZ6wEg0tLSZBq5/CJNe4uW/
RyQRutD/v9oNiP77fFEb+tHF6dxwnipneKhyCutABKVlXS5Fn0WsSF6UKSvjbX3U
5AXKc3ofPkoorg6OZ5IxAR9pKqkaMBSQnvFYg7dEGH/rcxhPOzw0wcZ0dSH5niGX
cFh69x63RLrv86mmXw2p3f080d5jrWZwYC4ez8QYS1cAmFQWbccLj+QokR5GTA55
Subz0slq+oSu+U0wpAvx4TimdctBgtcVKFWRAx1ec6kg8sy+MoaPoocKP/mgX3hu
CoaWZr9ScpnP2Z18X8c5tCLVHfYRz54hWUPp/xIbUWLjEr7LTom9iuGE9tllzXPt
AV2uxG78pF03qe6N+JdIfXcN8kRrOc9HwbvqLcxM3g6on3Hq7mHCBjTFuPBUaNG7
yxyQcOAF1NyKaEChXMuLMz5V6wnl4LzFOtJQaeu+b0P11NaoYgabIMAmwY7kang2
ESH6Wbfyiyi/wplwBbrUdVl3AZBVe/1Wu9oflhBEbLQsIC902xRCFpHTQmEcDVXi
29HFmcQX0EIEdwttMOVkkdrSHx28Zg3nuEW2/6gokN8eR/LSI1/pMreG2b/dfVfx
Mb0FxseRJQlkyigFpB7KPk5mKB+Kv7Q5Y95dpqvk7DKk5Of5soheftlRFs22Dcc3
yrCz/9sqx9pa0pfGIi87F0S/NrHKvnfQ/YcRLMbc4aVXDe/osvPPO2gBvR6NDZZA
j3Fq0plZGQyKpKiziRBfZSpl6QOJzCVux9+PbeGqZ88OjhkrfZfEBOF+QypxrEsh
/1SjXw1nFMhSFMhKPXdBErwO47pwriV0EI7WMk/BK3s17Q8nL5GtS8xZwFoYcZxv
L/+gJx5d892R54D2Vaz1kLonHt6FEip/ayjwg4doFWE7DfpQ2mkhcnxobXC1OIXL
V/1u1a8AWvNjCdjJx7gfH2lo269zGZHb9+MXTwQd37GP1vybh/ighZmgGDF9tE3P
DLpTeVdPzCJ8UyfwlelKSvWc2uLp465P+PTZ5pO4+PV286H9OXWb32oZry7zvYzg
vMDB/97VddiWGfxBCGcE4WlIUhEO03+qW6ZqyrBOx1pjD3ytK9byVehvbYColzM8
2U7RIrYpWMdC5lvOX5lyO8gXEI5Porjb66qISO5o7ZwkTzL2NURFiAXKkVMTKDqB
ZzN7d76XNByZzVTaNXdYNBRrcaPWEhF2DUqImsS9v8tnS5ypbPbbrH+fWCNVi6R4
U45rhfMpMk0uu88kQgJWoQn8HhKX12R7AGbHVQXP5Lzk+bkk0M+D5s1FGbHghbUq
G5DW0KQQvfC7MsxxkCjX5VV06zNuQ+tGr3lKTq48QVoDtc/o1jy+pctgEYGYd5fq
m8cV5seuUE9j4/+Y52TwHZdbAE8OqglU9qhUItkqE1p4y7ZWqubbg9VIPYBhAvDs
4H1zsL5S91Q2hqCppXDMQl7ocSuPv+Xr8D6hJqVecy3+ZriJUmLd+rpyAjEPoBGR
T3Y8lMUOkrZfums72GzPNftzmvEDtBikt+K7+QnjuHZaXwTOCzidNi4dFRskZo1G
WCAhkbTM7oZtKzbhBCcagRNzkMNqrP3x0lnXMVMZAXHPtJxkY0P62JtzNeM/PM9t
LEA3jQxDmlBIl9yggyyxDJEsuSVh6HwmpBiopPVxmnsG+2Cn3pC9HGXJP12Or9I0
33kmunrwNmG69Sz2ilY40yhVm8L1bFYS7qNt2QuYGapC4eeGvR+qHSp+b4b29DpP
FvN4EPi1sIKVMnsE2+pXu8tt87SVjLUX5MCFFszd52ZknnxbaMfDkgtLRRJYXBk2
s0fwkzjn6NovjDj5lQLzFzy+0S3w1XtgYViJpoOPAXX+qeaumfd6KIJHZvdWlT0Y
4pPFwK0HfbkHphQDNHfi/zkH7G0GbwzvMGtaRveM1PEwR9pVwZ7nKRslm124b9UJ
ioYxTmH6bSEZtN/YWj2c/sUXbeViq58mjVGPBfERVARS1QBslrwKHKVMMvawz1Xd
7Uj+gSqZxMbxVl7FKGKpVH3OFmkIqQDvXLOIZ2BASo4rVuuo7oEl6xSbnsk2BuEc
2PrFCmrErBOYA0wWqLU5ZwdTblPZsBMXzaRzmCceyT5nbnBGodHlJqvuUiaH5z6c
5diNdAjs3yEnc5disgUsUvsitgZj10JH3ltKX8yMNDtteN5JP17jKEnE1unsLd3q
YB5d0PZSZIIZGoD5O7f/m2tHguehxrfgg32Ebzy6cqhuD/6nKGxlvQyQnl6J1KGJ
JTcZSe5P+Y+wJcn8y5FiYXApvkixeyA0xKZZ3Sb95NXrSdiMG1LCkoBS+nF5mkmk
tiQueUFNgXdNV6UfOxcyVG6HgxWBWJjbhv5LkKltbhuGFCswIPj8qprF+RbhC5HB
u28j0geO3zdAFbpLGjqIgLw+8rRHlQadQNvnNOFiylcc4OD+lO+gGVJhuPoDqi/r
FsAPKaqHLcAfu72OMTbcv8bi0xSYeszOO7pvLZEJv+nFd1zm8HWOPC1GVtXAnXgc
uYW3zPrYw1xlAyGQ80HQGB7ZkBzNghggcF9sdVhAaaduLzA5D/8q1WuFYzwiW3SE
kAlyxGdm3mZEuGAIe5ln9wGEdBk+VTEqUFueTNKPqrvI/J8TN+CZER54TV3+5TfR
q7ytdL5OU6VlBYIdBPGlqhnHNsbWHoojOhKRBVyt/UO7/I1v+trVCo23S19zKQ/5
UX5mz2ray+1ETrngObo/l6f03vvI6W6mWjfJLyErHdNvlcjuM+Pfjh+7PmQF53gC
UhCWgtvY9O093Xa71teLJaSiVNWS3JMCFwfa0r4CzIEDl84b3wAgUhz5A9942B/b
CBhtZw2T4AzNzG9SLe79xZO/ooUbIDvVzjbXG2M6p4+kfcCap7KJ60cCHpGP0ulH
VSJwygkURkVzxAZT2cbXVhBchXKOUw3XD3PBx3ifBtyArhYmUA0OLeemxV9LFtc3
HeJgp5Yu9VE3J5eqeMpOpky/H0Pc5by965TJhlymoZgKs79Z44BIi9iMV+BxrHIm
e8BoxiGK4n5vWQHK2l85pN0R8OlXVkxYHBTkAjQcRnsQCp0AAXTR0cuuKJwY29Y0
rWCXT0c33TtOSZLe0jlD1UdXYe0v/Ne9cvgW7IC+qcv86pk6rv98zeu0nOlhF7Q8
ARHm5b1rAruWwiVxbnJa+4T5T93O8uAtSmzVQ9JJm/1ks5S1hvm8iNYZ4CaZTfay
deFnlTsZDbtkI+G3mpnqt+FrjRSWUk+NiKlhqEtgLmKvUQsgchX+tgzC1JHzRMU2
iC0gF2WrbPTPJFeA3xrbVS2RGM7COd5yzVAnad/XKx1CMyfSXyECnvjTOsNho6g9
bHGcKwlkO/J9x+HfOYHfgkl0Bezw+7+nLeWVdCb/DaQ//cYfJSbRZ9jEDfHWabbV
wE2ehVJgcFCjylT2vJCBKBkpujOQKfYl/XaDecXpGB+C2QTP5czG5vSlNxde1pGP
l04rXwqYyD4/8VqMOYTGej4rriNtHDoG6aexfaNo+zI5ZbifUl1HT2k+b93GcHDL
TV/fpcxnHDN485cPzm2K2+nvd3Kpbsn+fjNLwpXiKnRvAPPz5RLTgM2Qjq4/HNZ+
RnNbnvxxQ3piXYVN3sbpVqLrybLEBYAlxkI5GfJsC/yOwUtoY0aKwbl8YxbT6FiM
5eqSMGkNwldtakhdiqAsNjcoyPVvtjfEV9RalIkE//Jqr7DZkDgG3Dwo50gzmIXz
h4PzVhesjeTlqXbCcTJ6aUQFkwugyiTiRr98cHTU5ri7QWCR7DZ9KYDJB4Jf8bUs
sy08GoF/NdzOvyZBPA7EGzQelrggLbDT8xGl2C7KqSnPlrBfe0s1M+I2GEOB/l4N
p4rp9var12TyEN2oKJdFtKHpxVOGa7130rA1h2qC6zbNw8Q2A4tCm1Nf37jo4EVS
CXfF9BJFEsaRlEYEakdKlrqUl+jgJN7ODPPp1eG9GzyRTjeaLiuqpXZCRv92FwUP
xqmCaTdcQM7tw/fKMASsf0wVhu+68W47OwLv7IuzMBxRXkFv9cNL+3HQ03PJXuwe
wSwcfW8AprVMJ6CAYZcBi596VKrUPNQRf+g1EovOp40zcEAhkEUHNI/jmucCu5sY
GA3akl6inQPxFInJLtsFH1pp5Kh95VFqwsp/DJNdvZfYQxNI61fxm7cj13OC7RH6
5SCqRCu0Ci1Af0nnNqjQ4zBuFpYBLUV/HmbUDW7DRZYQdkiOTK8ZDGG445stvuhd
UDORF8ZNg4l5HdYE2MH8rVhCnKXA/99oBlzzUItQ96GobRktHkNWdgKMzxhw+qnn
aBEiqBUk7HqGquTr+iqA7sivKXhigCt00Leb8ndRl2z8EmBEuvmQLfLrhtnpPKIg
5IkCWUu9KmpztuV+joQMT/t/FKd14avDPymZjN4W0OIYGAsV7mqm2Nr5lgusCmw6
4Zs+WZ6/TRARSW9PdvJbwuuesbJ0bH2lLm5HWwF5QR6y+blDaK3IZdWEkb30XImu
CPzKi5HqrQ/egroZqu8SiUdO8WGvbBohpUmU6GeQ1pZrd7HxW29nmJNesk3k1TqW
ZoYDOEz0s56DGUEzhd9HWykn2WWj/143Jlg5QiNnjxcetHX1Wzas9zFtxCZ6ZaWc
seOvqSJIJROV0dQ+GS9SclYcNchqmDXS1GCUAYR9gfEspMvgglq8V4Y20gzI6Fxb
92Jx/KRbYdqzdf3TehDKK2AzvVXAlzfCTXdG9zZJlUXR8223iA/PYMnD0+U1Uh8e
12LH7VLbcGK4sxzSRc9SYfXHs7/maYhEET18xfMvz+/7tBkGqblYIhlW2/IyHWw5
i9bQtPd1M7Y78jOMNpKC/Pj/ZuY5cMg9Rh+sVvsZzA14d5c+COwHleOj64yyjAu+
2p+e+Zp2mUPTXS/xgSuCZLXDpFlmfYoPuc9QSImJmqZm/s+yWZCs6sGcNQ3xhFf7
Ohkwva5zMaAulgg/WTJ9E44dqoydO7FNS7pw4Cb++X3Z2PBxvv9T5JXA2FgUJDJk
8LIvVpdWPpRGdRxDW21Z7Qf9rnnurM/TV9bxk910MZnGvlOddiXXQUDYLpSXIHZE
hX0O8a8IkRV/d7t1dgWNXOKvZoPyzXyUb+Noh3wwC69SkxmNk2QcRfBbqcr49SBi
nplHoh3o3ThQ3PkRhP2qHmdN6FES/cmxWSFxzKRPJ3HjO4+czh97hrmaDTsRdV/h
4TXlHj1uwes8v+zqZvu0t0t+km/VRi83ajm2i2e0/OBPX//Eh7bQxZM5Bn6nulaA
Be46ouc2jtA1JqK5fyMGI3q2+4/oCnqODKKRJuUXgpxYNKJMUXZbBG1yDGtk2/lt
Op6L0k1Ynn/BPZukWmSCBe8AkjOxT3GZhATPx+BpeM2XfOGrbwjxfxqIFnhvOCke
RXxLyNlUr4V3esdiv18Q1Dz+Ubrp6n6kZHuLsADGG/NXDmZ8WHn77eo1L0ASSL38
dIOdXFYEbpLqTqZJApJiGz0bitdozYXufBVMX/g4S/mv5MyWeMrG3iyDQe6fykTo
/GdI5hUtIwKY17vhU85eewMenkiCFEUIkFA39spANaPrYwNJxcTyIlp8Jrzn3mtc
2umkOJzFA9/ty18ahNi2iaLJNzPNotBWIkMEwGEz74AES4GPm4a9LKZyUo/lcGPL
LXtCjj5NHE0kKde2iulWWAk33gzog4A380jNLSytj8tWd87r7rFlEsy6P4L7W4+t
gs8BJVi13bd3CvAMa1L7O5HpRe+E23TE6d1Qxi78J638vtWBv+96lHfFI8/RiQ5m
q8aYvj0Wq2JlNmk7kO/meTYVglu5T7Jm4gRwynB4UV7Vt0x0fNcD6rtidVYApldt
RpQRHZ2tQDb2hnNDzzm9Bqq38IJ7omWoHFzk/jNXCVAbfDNyPcGpy//doSw5kQmv
SwuMoDt0B0/0qSHeeS0TpNV5MQ1wkQl+GH5pkBXhyWDeXP37Fb7xkwKtN9J0svDF
/1FF4Fr0Z7XLzCWmOGvZ9EhhvO6LpIxCReUJGIS5jnb+qwRbk9SlWgtKqwh1WHrf
0WcxF2b9UdkHYhJ9cBWDNbxQbFTunaJtC9Pjpl7xLMyUn3d2zumQ22k8Cf+uifh2
6Pi7sHApVh3SE5R4+ilUnRoHjVu+Xdfi21hXmXNo+B3SEkSPkZSTkGy/OXzB1+iF
59t2JhMOi9fk0Ys3/H7USTcVQDWIbJ/n2X7p/Er2oMrLuy2dBebXHE9zFh4SUO83
oIiR36HcOW9ErqRVWvR/+xvUsMsPO8jJnwfAUvDqN+tTAKVvT04atoHp2LO8XY3+
tbNRPDAj2mjHg2kX+ldtBLGueOx9u6EmzS7XVAXJiNOScBPJGrpvhCny/6Rl63JI
/LZTPIb8aRXqxdnnjvpKf6cJKV9FJr+9nSiJSAs21iaMdnAW9AAaDq110RomJw6M
aFmbkkicGQQWDAN1He2f45Ye3mENhdoG0ZGYZP6JQKa8nOzdqXb0fP6V+/7buWk8
u5WFdXGfuTxf8ag0BmwJffJgXYa/zYZjj8jYJl30afFMH4riVZF3W3dByC22qDEJ
Zvx+sl5IMc0He2cRcoVseXhSIQfbMQK0Yw9/UVk8A1mgu7gdlS240koMeeitFv2J
CkjNYXgEecjwErS+gK4StF5mfR8Sd8SUeGoFhjmq4JK5gfgDikkItwRBLUhxE8Jn
j5/SIeBI8WeHGr/uW4o1sK2YeWmuzrNEg5I4WY02gptwYki0m86GWKCdjVUTkWjp
jJwt20/A7xhaeWcx0ftHqQtkxfWwgsI5f1ZaQJkMNMDVtLfKDD1iAmBOKEyULO2C
IKlbdxUEaf8+q3NFWj6qvurOlyOnF9vxpnIA+fInokVHtMbxiX2wS14AtuHiW4IX
W4lLmZtKDgwSSj+R3w6/N5Acjy3cravG9u1cfFnLhbpAL3DB4ytAYxgqvCjP3lO7
0amk/UqrFCG0Jx10N7GTC7Gyzq0ILQ07ixQOM8eRg/GG8M6gn/bOe0jNq1OZFHFF
O6qGxrQyN98GeROytm89PwPchPCadUyl5U2ZoPg5OtyOW78fODKffXTY98lWcHMV
Aq5uajP6jRZBCYj7k5NcP8Z8T4mqufyBh/TLxDrFcylDgIwxa8nSaTtpO9Sf6b0m
o7lFp3FNCtZtQ5LGxVaRzkv9ZHp0NIolsLnyFENFrj7hp0ola8CzIwN2IAhgoHCa
VGkS/wEQninN0v2z+H/iQopSy/KUgq6OTmV7fPINyYWs7qVxPrQW2B4NE7rQe6UP
PspIbY2SpeF4IOWHT2VwyHY3e22NpWxNIhmKu+ci7jgOgShaL6k+jl6Mt7jlOO/G
5Jj+7jzRZezq8bvod6YFYCuVfrIpCq4++G3HayCcvfhCLWc59bdV8Y+sj9M7lDxM
2CnF38Tt5Bwmwcfp/Sd9YDNQhMgfpBHENZIFqDZ/f0X4J3xiKC3vid5RG8+SgeUD
qasrWZnTsBG+2cPnrp2yvVrAGfbOtYyNMXOqbWdh01aGtT3/6jlBliWp/qHxm7MF
bEKoQ4ygFd2iBk1mJgnstJ1jj/PacM1lNlcL7nYa/fC3cJ0OZtw6yXQSvNHv0ayV
eLiJIdSK+iAlQd7XWgk+5+ByK775J9Lx7RghR/zPqsVCxi66A5j/EshUkbBIpoBV
SB6gfqJ0BCMGVTgoLmuBSVxZZ3bvxbOzLQGv4Pmh8rFp5geau/Wne9XajvMGUSWT
qIBPsULmwHyuF2vrN+NwXRiPrPthIOrirThkF/IlvKr6/mCLHpuynKHNdKWs6Jqu
n6yUqBySo8kG1qRd5K5d2dpo+0xa5e/6Sfm2jrfQCK8issuJztLbanN/HAtcDlnC
xHyGMDzDRSnPpTn1zv3845/uGSpqWwitdwGA+FE91UZNTEVZZ5OW7pzsiAVuWq95
1JRs+Vk64hkrLackcAzkZZ5H9vp/jVD6whUfGoCmL4PRTbzcbPP2ZupliQ0dgCGk
l53pGQ8f+PlsORHoDWACU95dh/cWL1JQH8HjdBa64FPBZlFK0W0U7FrbUQoC84X4
kwdWXbvKVzfiPdSvRneypwjQDcFKN+dp+zIext/ciVyIzvDLDtmlTXDonVxVc60e
mbwtzKShlby87iWM17P9Fj+uq+Mo0MoM8SiHFO3UVNjwSDH1Pko0Tm3IHXG083Hx
MryIbQ0IlTWuMyssJoo5Syp+/+YYJKkL5CWlItRNzk/53/YlcB4yFUH/+W7aHWqQ
ioCgzIlSLBsOg2yNki8ctLzdlH31qPjKfaApwMCUlinUOwchlSFiaQwzcXzn/Qw7
5KGGWOGXupMXlIB9E+N+JQVrPy755TpvO+9bj8vf9kxAMFY8D98OLbwUN4zSE6uT
GSjrR2hBiK2sqhfm8gEB0dYeUoE/bxJk3n3P/cDJBYhQtzMcO/zoBWUCTdCMh9DZ
0MM1w2l4xDYX88mBYfiGgXpioATrtROJy/zT14cjM8Crd2ArQ76l8KBW1iKwByOx
OIWaehulGc67Baxh0oYFRbHam9XcXawh1TUZMPw9gCffZfs5eEwLicGwdMODC+Sn
G6OsinkzpnjlqiJqsGD4w0e4vzjMCQriAjKmnT7/oxjzwJGE4n3SARoAOM8ve2qA
F+GDJwM95XMdoxiflYoIjAlmsG01RzlU9aOJgsCLcfb1RI8zcfIUbT9BZFyBXCle
flimyplGGw1piny5B+yTw778a1BLFCUR+yHqyJPzMx8iWAPGVIGhOHg4AhZFWwGa
6H/dsLN20obOdCX6DmBbp18VbFqxL8Mglabn9gMElQSuopqROgScP3pbPEDoh2bs
9oRezI2k/2KLR7yHpZ0q1iTgXsGYeJpldj9g2Zb2L4OhdClbwCBQgtWSMb1loim4
tacKfPEwhd8MEWPEDuWwMy4KSTnkj9YR9w9f6yf8LZXIrqTMmVqbRNdinCC2uTLY
yrqejWQM54Sjyf7WoLV1TM1mrje6ptqvfYbrP0bP0nYgJTSxO6PWf5ZdgfMmxKW3
CFXyzKkjWN1XwOy2RS0q1bfIqFcnnZs2sWn/nAV2AD3WFO7NIFtZ+lKZmXvQD6lv
FB3eaQev2QNZnntt8XWmjBYWJfHJYya0lvmxG+cA9FpiVLRAWKRs8SFjA6JKrc0x
A1NRskCvKhIfDB1Pcc6Et6uVk71b+eFbh/SQEv9TgIpfa3U/r60PZnSfaTgBEV0o
vyH6Twx9r2QKUMVxy1Jqn7eMOphPHV6bGcK95XYGnzwuR4bN5hR2rdRxehNPDlGa
sjLJbjCE9cr2e9gmDgadIh6TZrUvQMJzEtMybgnMWdPwQ0GMzRoptQos92eTVevd
UqU6cNdspI7/XUnPEpHMQwHb7bqkDSo4yUEzzSqNlDG75kKtBlZiB3vMk/zvZtFP
fyAWxOegWrqB2zWhTGN3e+iLQ7Thh02UbdvubO/DXM0TnH+cvtffcNG4a1grRg/F
mnAJySqcIZMkNNPDHZwhBDbFhIqrBFKt3F7KMIDkGEQJhiPz7BwXjYCDOwOyGol4
V1yM4zHJZ2IpWNgw+aTWI8wg8XaPPKuh3isJLv5xO2gNbn70f0rPxer6c0LCxnA3
iB5OMU9ssNi9Uabn4MuuTVd3LiRbLoPLZkpCCr5S82RXZXTj84wI3iVYUo6jN4iq
hmwEY7c8otewk3ODpMBoLYKW+8tdxXb8ojv7VKyRk57kM5Db7m6Bc8kX5dCaPK95
NB5tfZk5Rsc2nhYUGgEH/u0uYF0HJWXJrzjptezQPoBvPGwxR4reY05sdTaBWpPO
WGYUCQAzdITCsJ5E0EyxgRJoeysfh69Cnbohc1+3wbRTEx4wlmEXYSrTOno9Encv
EiAojXJ2xxuzcMt5yxreHpNaIITodQo8k57TKFLEj/Turjg0UFxW/RW6nIPy0RYh
OwUFzyNhU1KfDISCGUXJdJcAySpMXKBKHg/D49WdoDja/3qKHB3PhhvE88xFiehw
Dk4BSgqMfNFFK1h/hOUkUSCGh5oYk2qlL77BOsHq+X84ACX+CXheoK3BDxeHBKBD
SUlv+cQT9CsPYsVhG+YkVperUBo67c87EBrYjz+oR39ljzwOw5Ngy9kruM1vrByD
0400PeDNPS95iMAoA7ON86AJ/ihSrifaYFQP6rN2Gm3QT7tuX1Mg+zh70Cc5PJ01
DL6zaaIcppow8ygSpVFi0EvXLi5IhIbrwLQPgcZo5VwgGGvWcQ2zvSUQ8ZRnSP3R
KTKDpHLCd31SoRFB4OC6/VNXZRV+Pjmh7GHU6ULfmJ1Qr70ymr5SkpQWH6DEWEr+
rM4YRTQRfMLmcsy8PuFLqoxpiV1kuRqfdngla8Q5rZnBwcgto6NUKdv7ah3D+nFe
1V5hpm4JYGM4V6oJkB02c5EZB50ZM2ybsxYQBLSeBmfSjYtsJS82Haw8xLF5OM99
K+wXZ+yMi/5cHADpaOEqKWzUUM5zqyA+PR/Hg0Wu+GBKVsPwyVGLf1UgupgE8S3D
6c/6yRbeLR9TifKPxvFuCMJGEgKsvbNcf+lGshdYsvvWvXkMlAeMlI8XtRWSGVD4
vMgoOuQquLIZjRRgCn/Zxc2ve9yWYWpujKYtMz7kj+Wuib66BdrMveNzghE9GqxQ
kPchavhTSkl8Sq9yzQX8VvwQ+A0u7s8xn+1c6xZ1GKY+6dBt38uRA4py3pUX/KZr
UUuygvF1b4Hj5FyZzyqB7mBc21aZtq4gtjC0hjhvM5CI49dLGXslesZeNOPKuAbI
h3LB9BasSB6cMDVvQfGY8aWTYZw3exc4mg/OhdFn3ilemD0EI/2cUUwpw4f7tfra
rbw5ASoBpWR+Fof1X2svZSmAtHFbihI+CfbZQKZcNluMepFV6rMe4LRr1cwI3I6C
kdQ7P/NuCBDsJdxOFkrDukOhXDJwWY1GKA4jDRwE1nODArWQxogqxvCz8nNwakHz
A6cpN8+rARdon4GoRmD/z2x14g0fxaPKQu7ugB2BwUwHGkrY6JUlUR2+OmqxXY7S
e+zWike6yj087NbHz5anGiVKWz/JjT72rVrZifbxy9fDW3RXOCAcKrPrzWrI3IcE
PSsdokgN4WSHQ8ixDJxmoPJhDR3rruBKooyik0Sv96+jo00Ek99TJts6gRWyG6y1
rLPsChxtxg9X11F3yW0xke/mwKcTkteN7V4z2o1MhJ41ThQDyQvIByTBu5S5zh2q
Lnphojb4qQRVG23WeNSuv+f6HcaE+lWPIbj2rcD10cGSK7fzZoBfHM0fwWGNPe3J
xsfFwvVjCCvYmreuseySrz4uMJEQQwSVT6AkKJjxfMjtvpGhGNPK9SMIIeodFXo6
VMtPaqeLvDOxHqwbnp2GXfnTZU29il5IP7kgRpdSRrkZ7k+NDKAA4qbHSgnNJhHP
nuFMlIbUmb5opr/4n77bf7cEleT39wc4XE/oo811NKOIFefuP2U3J3PHeOPHflAR
JFNk57CGFLdJ0MNygie0JVcM22WtVlbI+6sAWby9o8MukK+tGL/yi3jr0e4arEUF
JFG9Jx9ubnn2LpzqabdWMF2z5zprg72vbLguodqcnzkQB20pZUqHYrkEFEYsor1Z
iH7Ud1vd04YTlbhhnKovY9lKiQmbsbdaMt2xhqklg1IsvHYdJmUCQvqYH7k88TUA
pAVEswJFosncyWHRqtCgrGI1dQfwzJ8C8HaOC5yL5DsOeWZLEzFChhe4AqrjMU8I
VqVKGZq8cmDPfMyvlJ4au0ea5h9hTi3bmwoy1aD433Zz49bdPwI+/EsxYLMVdaDs
AmrjUvsVDSV9I10sb7VofLzKXN3gm6uhpcmyk3f19fEtzcRWJwTD3BSugimcgl93
EJZ0geNsxMFtxBDbjBlGxtckK/WDKahU+4Dz094/9Ot+DZTX2WDNMzJJ4hSQZgvG
P6n/85Y7C2vYMsIOJkPGRAr5/sE/+/RMjb+8gcCuUAXwv+2QFBUt1oUTCYmcCbVM
fGEkf2SXDys+fGP6DJLpJfihqpC+iA2UG1mAuwL19aRLVC4iYoynBoOVQyZPVjjk
Nmsp9+hqDlHFKXALODJlbcC/ly9BxCkIxmmgvPW7oIZnoznm8zieqmm/yl+4wro0
PpNzsfQbo4Gsj3simvi1+9ey8ZOknEbdLJ1i8avyz3jNyyIiyzsQI9f67oxke/W6
VX0mukPy5g/1kd2ZfsHJosspwQ4o/cqxyJ/XUaRaXGIxrY7Hk3jrhPIa96xs3Z83
ED80E4ZB9uK7WO2+ZUFn5PJ3THR+VwWU0kJLAQcOPM3tOtIl7o6hz13fI5NJ9QqJ
f0VU6yb26cP4aYW4n3PeQFixklexO1ojRIEJlWoCPd5JWrj4gWjimTk6H6PZvHD4
24zLUBCskwpawMoLwHKpi4Y1WV6S3yj7kgk8dnv3EJOG4vAwGzmNbWm6lBmdYQ0i
ZXIYktm/gfLV+QIwKvEMk6ydREAjavs1b4cLBvBiDgM+j/4aTWKybjpWXMUORlZr
ekdXfoMA2o92nJByI0EeGGiOxwlHcNA2xKPkLbuw2aSEZvYTllktB+2bDiIVUcy9
ofiafFwIirjfq77Pv5CuT7D4CqHXAXjuawQ2dwUJG8waSa+QGPx8Mp5p42UNxyYB
RBg4Qk2Glq5rrwZLHDPwj3g544JVKsRplWGo5Pgz5LLur7Y3yvaL+owv8gloGJMF
XYYif7GpcpU3ru+6PNuTOfnXJ8mYDm3psBz83t1H4x9V/OXs6s0o1G8riqTYhsA3
k8nTORIj19mRscCccQhM7kCVnEjrGAtDS6y9XPunW13eKDmjLW4Jss0gj9PdT8GI
R7UFIR7tuHQ2rzFtGvmUIOQXohLScDntf+NPis6hxpi7lccf1vSpOimC+IW4a+Kd
tlf9ZwIvTwMzzZexD/9cn7NjxXHAfeDBdINrsdnWOj6fT1Wj5t1yQk7jeBifIQIP
I82f0S0GFYcGbSHjbK3PGKUpoA6Yvft2rilAsbyTqcD9rTe3g63m9IOYaAGUQztu
waYyxRd6z3EZ3BGVgYgu+RAF6r/r/v5acpmVb5MLwYIBVsSsdb4Q8qOfJy2jzH37
hT2+pF2F8rOzBvKVBXUWChMllyfUNKyWmv+7DPNzy1q86+WExzDdgkSfMxy3/PzN
oZIUyQ426EKjH2xomMVI/qpZ4gm4k6WgvX+O0k7el+I3Xjx9FyXnJCyq9p5pulDx
xKaG5L/C1HiOXVZkXLVTRdWHCVEIM8208GvWIPdOQr4ibYlni8dJiQxtg0Xw2GQg
w8wL//r7VVbyz2QZKCjFgjfHlEQdy5vH43pQFcXCYGwty6bhdaO9gmTWPOqamuTy
8GPxZn20lBQDjNzRzNXK5gdo4NtGibdX2qB8kSjP1aPbTGAyMc04ux4PYzKQvKhq
1HeWnCVdruqC616md39qjyVLFq+JC09Tg1fZhVYWEwDhlnKgah7Mat42n7ACyiXi
DNO3MSuyX+GMDxxTj9U4GYrJw64FhKUGHmJplV05RzYdi0o6B39FV8mm8NinGXrq
D2B+IFokk5UQK4I4hItC5zflO6K8BM67BSPVLV0oyvIqFVH8PzZT1cv+StokQIH/
4ABarA2mJ0d0eFmrSZtpxo2blTfoJB5YX3yUg3olo/zR8eTxwBOZURfcXTljWiay
ZlxvPdNNgFLlTNpZ5zTAwBjRXk2GgCaumwBBPp+t2xhaGPO1HzjXZKM52NeewP34
+SKKnBqVDYYio0716qTA0HEIcfrdRRsQIt/yV7bEtMYRXWbABMtVWt7zxRKDCl5N
uC7aAx9C07+MJYOG/PExuY1PTkudjsf9MfkwpkLRkpT7kTWmIMSelihKHfnzJbWQ
fanejpp87aTKLuQIf9QaWTUTWU8nN9triG0RsXow0LIIK6gAFa7YxtmANFhm/nRL
Ug9myx7Up7fMeJByL3keDdDMFBZvVAxNEnrLLoRR8sPoJ2Phs5hvEBqu+AoBFMab
pSPUECrhIJ8EsShg/MiOSJY7wZtANyAvKF6MpQ82qBEGVtOuW+LM+xcFwYebwBsh
Uph5F7Kdzmi6zyp4pwtY33sUAKDPNsnhW1mUI/D/o/3mEUOoBw/Xeyf2/MxSfz0l
xbTdNbQMG2CjTnWdudH2Y/gulFDiWnqgsXjYwzEBIi0axjirJXdUqyCaibswRWcP
fLquhglpOlVZSKdQ6wd3KDOYGyZB1TGlV9BRgRSc44gYvSxfJKppckljizh4SKWN
dYo0NKb3oCQcqiorVT3kIJZdXqMSkgrZS1Ru4Anx8S3tzJOXRGfaqQqcfdAoYrai
+zAIqRntFCBr61K7qOabvJ8fgtoBuNemxSYeLUVGF7WI0hl7h9P1uqezcsDD/Ocf
zCMg+g4eFFe8/OgVmkjaTV8XNdJU33O4FbtkMpQ+7zmMx30aYPFjN2waoOol2uyQ
3/l2xWLYA3arj+mjFJVotic09nkCbkfl5r9mSWGk+mjDtIPggjH8WqPy2593zilT
XB2omhXMlslHANL3fHomeNbq1F3tQWkhNbXAQO/s0XRjVlH9UaSXIhzXf8++tvRW
HwVkarLuGSxHQS7drAOU5oK49YORqW7fQ72sUpRkwOlCCJrMQYQpXxRXczqjvhOb
MdtQkPPrAqKAhZxrbKMxmrRSQXNUh1Zbr574IKTTf1gYQHVEJfn5vn9Xzeey6unM
o3igaVXf614B3m7M8/zTWSnVNeniqOzMpxLJfui4xsGzW6/JYb1QRIvkZIief4tx
ocCoYfuSaTviR59d8/tixqrq5v86KuP6Lqsw+qzt82kQ9G3FzCaVaBn82K4N0QXF
WeflsM3N+PGb/JxrxNKy4yZS8H62BkJMF+aD0Omf4M5JEIH+lbVUWb2uhbsl/XnA
aIRuB7k6pjIPLVqaVceyM92rroa1sNslYyCBCNlbEcwT3LoY0DBMb1urEjPxxT73
KfY8+0Oc1xrVvsZcTJa8sKtXbLq0rxeRDKH27ERlPnZISMbDofuyHYfIiZXmdI9k
X7Eq8ilMHtZNvgQAtv5jnwitzzckiFMcEcXowFcfY+1YHkMxwVGANJN5ShKmgfKF
D/lL1SEK5mPZ3gHRIW9B0BWTtbrPjLhVm5UxlgyywXpfBmPlI9UudcRPrNofk7GY
d707aTuIWYI86+Kn6neAMSIozsQOaZhTBCWT/qQSOt8yetrU9D3FL+GG+Q6jsL6h
yq0ZJfGc4ULk/ixuLuLG/8fEKvInD1V6IauSyV1zbckXPXLjNzlkmoMaCBg8LruL
0lQOQjaKaVWC45MgzLxtK18ZzllzC8DPBXpOIjUGXR8vrrRQfYEEawpCclNOL0Oe
UTY3hZI/n5w9R/8zvv0aDHjiDiSBk0fyOL5ff0UgcMVMzsqC+rZVKHn9l3mfmDVE
/efuj/0V18EbyuCbC36zzjpnErqb3tmm0FKD7D+nidQ0zCmPlHeWCYivDBQyFjvI
S6eWs6cVEi1dT5cwuxqyw3lGmIVdKQAxPDjxMo+r0/xp3yhGYEI6pf9ntkyXofio
hlgDxWit+s1N21iCB+gt00hAmJgYxlQQC8W1wXyoPR3ghOmH3ZsEDTeWm8oj7+bh
ahCS0KtZNw+pGp+4n+ZaGsTPfiIqs7fJFEYlvKgPeFGMX3SYY7bTuqB5n5wIMkF1
MMzZAyzug9EC54zJtoa2xgKU41STxkQpWVQESAAqNRV1RYaCrxJXUJO1cVfINTEI
zn4TSW4vb5qqYMEVKbRzopGmp87IzKpLgBUh1YYfnM4CkrAT5m4P0v+T4QoMRjgG
D7fxeZozt7Quhe/fKonoMiTUripGaMgAs7dwpwVwAdQ4o5RqxnINByzvrMjYXc6u
jtI5pwQbQGYuI253sNtxW0QjKVz3MbnY3zLDoqRHRg38W+1CgwyAHvkBptjw+jcA
CWpLTZCEIcHGS/UkBKDARalx9H0EXGLIpd8cSt2xlXqog6SYOB77ZrDNnHKmiQFv
cBaYioSrmYwdzOZELxzX9wTZiV4uqHlPIhnpveCBHYbsDYhyVVsHWJmzP3CRkH6r
EMb53DQzyW8j0Qc6AQ5dE0p+cFUapDpYUgeJnCNZf/KUnm1xVH40nv90pm4bvpjl
E4R+PfnY+qVZzHMZOiixNFukBymJHiBlSD/5//p4+rikPTOXfxa/vlT6WSV2Oz8d
q5MoI4FWj0KQlC2r52uMoi9bvI0rEB3kWgIcjxjTD7Ja/Q9b7d4sEt70NCa9V0yC
J1f0kxKfrIZertSg4OjOJG7FiqxGpB3nkPR9GUOrPPDHVGbmRh7TSIISrvzcLXyL
OzTfzsibSaGqvxPiVlZqVgkAWeSdZpBXI8Hg9oqiEWzzQycAyys4VQ/++4YyCyLK
/JFgiamFri6PJ/IYERV9IfEXPx21FGyZQiWTXAWP7ZRPWKuZ7ew3ZGkCIf45I8w0
AY23btBGH6GP58BDSxhBy9vtUIhxNXp7tSKB+eZM1NcW8Afn2nE5t3FdF8NbDJ/v
adAXAD59M5taTVZ7BDZqnrlT5dXHpq2kgcNzGftwMrQv6LQ/ua52SckLZRzjLroP
ac7MsuPuMThnT7qgFc9ZhebPvld4CcRCm6U5WYDsoNP/n/CriycMvTK2l/4lEOHI
dix602Il25PYRTtcAfX7s1NoXJlMqqLLa5XqDJlbaZmnf/6om4gJSSEhWRF4W1cL
CmIFpry3kgAtSfdKYSruQa5cPSAS4vzIx0BG5/y5t2ebRIRx9jlfOV9guvViL7Rc
RMzxxGIpIblUIYYujF6bESKhpz3Ipl9+F4E/lvoRHuAKuQyH90y9FUqeHbe95MgW
c0uJB50eLy7q9U8/88IpJoaKebdcptwh5X1HeFh5cNCWBub98ilsBJX9lT3vEmYE
oEoJITSLMyr+P5RvRMA8dRMVEXC3PdvOjLVx/vSFZ1xtmPk+WfJMJfL8ryQuKlHs
gBW144+cPUN8Z0lhgMohtn4+BHkiTVLDvpbEKD5Kibbhe73Q7e/mokfHaj71hBxB
bHzWFor9H+lBHZ72O3/Etn2KhIL9wIlO39/6/JlmWNvjVj3BPK5OHJvsVBDYaQLR
QVZBb4izEDx4263+AGQiwb1n3vS+v6cBAchsUdlFvrd0YldgmmwpQyI99+gM5aQ/
SWlhZLdM0lFDt8aZjsydQgcwCpg9K2cFqU4u0yn/0afLcLydCei1jF8BwhrwZzWP
LqsdhDLADxxYHoQjnDpNMaLFJh0DN1re0HdwIKnx/XAeKcdoo9a9jrQj3XC7sUGt
qPXiGoKiGGxJqyr1WruTW8NFOf7+OmFwgY0B9GU5uwQqr4u+29FwXAmLbEYfT58P
danY0b0P4zU7xDTyU3LYAMmORD/LrhBDGLYE+jgqC1KQhrOorAD3nZZ5fJdeFjPa
As8lK1WwRAjUNkuxIlY70P2JmBbvlf1lw8MyGH3+KMHrd/vrFRkmHIAJlB39hPmU
Q4T1CTY2uOiPTGMuAgSdWmoq/2KfnZ2UvfRwK2uEPLIbrnvhzzDL9871blI+LnRo
4ehk0k0GhPLuSKuUmaZWB30mBEwnk9rgjSIb+14G9YP9T5maD6q1GQFUz6NfVjFY
oZAhX6lGrNvem8U3IlqSEtsh4VaRl7Ce7AnmDdXbupOsvyW0xyhM7+VTG4DtGEkS
S7Dl1K/6r/YZaQfBuvB5w+Ct6QUuEzqE/fSQRJCsTkPqfpLEJGbuhLcmaHfgoFjE
J0ezFWEltD8kreLJgBVDze+lZ9QzGCTSfQT0UK3jrxpqohqiifBbd28QiPzAiWwk
/fMCA/2/pNrZHVTlB7VTmkm/lJHFo12eQQKRQ0UGPAqnAjAGMMVFmC64tPdlZaEd
ddMM6P1cDECGit3afLavmzAc59PzqYb5eAIr5eICIN+lBAGr/vIpmeSMvQ1Q1Imc
P9EDPtxaSxP7Qtlwl3ndYp39vC2Tg+dxNIjddYazuS16x5KBpmwKRpOeerNlcgO9
hYMs4PA88ZrCKwdMMDrsB1Ftpz53jhIZUPDh9gjCCvP3qSuW2FxGaHiwPz709EM/
YDNa2mVASHMJ/XJUDfDcUNv4zWB3e3+y/4jPR68kL3t2W1008PvOCglUGxyOpKtc
0LBcTnSGf2ffLwkKpgtQIL4+M602x9WWd0XWLIauam6NnjKmgIswsZF4uV3EAU8Y
U00bAWWyuRwpM50DZI6/9B5vr3OfC+hEJdjNNAaMMe70Kr9AiYF8hgO45yhgGmJ/
2zh66Nu++NIRAxr91vejAkTVzk2f5d3wjLNdIF99d3sJXtqjaF62WU9mzvv3QtY+
BDHufDl5hxFGOyAG2m18BAni6wiwoaYAYrSiS4p/8AmmUMYYriJ8Mk9IRHbDs+rY
oQm7yEvwDczllGtWkEc1f54L6FX4tQSXM37ScZIVIxTq0RYpKaVZcO378ol/c2HJ
V9ymYc24SSOfNOyijhqiHrn4PkfHtIQsaBM/TqxFoQSYKpY5b+9aoQCvxgVYNxBW
0A6YLcXyBm9eec6Y2asKj3Gc58aCzfk9xdY6N2ncHnSuWHfJy2LUC/huopkD5prv
Zw5TXwMSzZst6iqrJpDyW1f6B67NiASCCEhOnqkkC8vhHPmSEoXLLaq1Fs6nPXZy
VMkSLQPkIcgryLSu5DzL0PGDi5EhZb2IGIj1rj29mJBcvUZJLLfdPVCD7Ebwvauq
9UbB+np+yJKskH1/Ae7QwQhbE1+2Y5Dl1UBrUOW2cTKnkn4GbpVP8FIeYUOEVyeM
3X9XLszQYBzhqJ4MLhUTvfVMHwn3PMBAgLYObD1avfNCZ9OfUbMHkHmgOUAzleqs
1sBKfSmgNQuphGVcNMI7aLaFbH+N5eL7BtVN/fg5QT1ybNwn4xruzLxjojDONzmP
JJu1hB2XEFkAnrIuhtLaZdpkUeUV7pfrHeRycLuB7XpVTIj5nrh8IZNT/p00A9ui
4TUa4nb8DXDsoRXB7f1zf5sBbvrdCWPbtr3Lj9wgcCaFVNrLw/vkeJ1bvnv056iy
si4rKhiCXvzBMf5bRALH5eAgCsY8pUBHo8hoNnCtdMxxvOTQVZocHIzUvHyfrNFR
5EvZpR3/vi3D/JshyA7B2I+JUqtyq4Crr464aIZKInu9JYQr2TTKVUfAh0F3y3gr
jrFDWauU+2dKQetCx0pvtzRyQZu9bCNPsvvqYVOKT9Z1qZrZzT2tqaYYo0x9Rsuo
58Fs6tQaitPfvKNcFOqpK42f5FwN6xxrZVG+G1UfQxDzjHXMMfsS54HlP8bRvlHD
iNzI2zGETC224SzgqMzMIcR5ffOJZ9JZu6SfYTKbZZ/cjFjuiUxXi8rVdOtF3Y5B
CZwLO9tGXmYYQkRkKWn3FAd2r6kuv/DEpHD24zgaemcl+ZAcj2f8RmFKNopP9A9M
eQwy/znSjozdwgxELRbpuEtv5qFxasjZJl0SL7830aspewGmYOXnw0YdgqJUY4RP
uPoTlbxMOm32ChBOGiBAblI3d30IQM9/5+Q7XsEL1Ansn/A2NYwIhxPccqFxGqih
syJkLdo65xsJ45j8UxB0QbaeQYzutwqKQ0b61heTR6kgJiOjA6IR0G2yKTgDAmHR
VUYk6YIrFJE+oZyb+gKGNYp/W9YugLJ+d5mQiy0fnWIlZ5WMQdZdA1v8ee2tWV5t
4HVSacSy3L98Uxi10v+FlPMWWxQOj4CTrUFp4VWtW9zavxiFkKkdag8+CKgY8TL4
/YVkj+K9Qyd5uMXSSsOLEvqJqEUqvwr1cdvr0FFgNxFzQ209tp/5L952dWSgiWXS
iokR6eac0FfN4vDKbWd2t1XW8BMjWBWfFSl10M8U5zykIlQZfHKVArEWcku4XiBq
wXvyQN/yuXIf8mtd/ANL56RFy/HGzHOdS2oDZgdjsr2JGiy1cI5o3ap4BBD+OAkG
UcxD9qEoIuJjygz6zWo0056e0Le6gt5JznIAlwyh3v/qurzUmQKb1hnLMBGjZCI0
DUySIVo48Zx6ukkamf07UQD/oF4aXusH4/gB2ev8bmAF3XzU5Nrk7/kdwNr0gSii
aNfuCVDHdlWNfD7axxH7t3df/RJtyqGeghaNqm/kF2w9XH4Q0iCTNXJJKkvxi/zT
rKcWkCOL7ocOeKwK2cvsMrB6x4U/D0/jYVjCDEUjPHOi6AmPintWi9+o6NSP0wXR
srYE+NPazzDs4WaTEGECfc3rTVi6WDHgpyis+iFKApwYwFr5wNDEd4URFcKtchNL
rwvJBPv+d5+NeAdxImMZWblCMYvyC3ffRNB3BrYIM4kefDwlV458QFEwInAemaI4
nn/8TZEEgUhg7TwURKik/BUidePzfKk4l/H9mskH4bXlAlh9THFG4z0IdY3beWI6
ar6JaXOJgS053b6p6/6EOTLdSjENk6tFfC6kx+MGul2/L66CiVhw5fWB/1g6Zpit
MfpxCWob9Ihhbi9gs3CNmPGyP9WTRbPzpNO0JI0f3yuxh1HeRzfQYqGxWsVCCxDt
H7jLFxbWxUUlFUPEg2lfGnX6iqDAYuJ7z73Cc7OoQdnTXc7PhdJxMtHTHp2X+NXF
wtAa/KwLUA7hVHyjXrCPrYRzJ02MOncvXdTV3x0c1H8BZeC0pB7x6kCRTUVdnf7l
jY/QVqW5aCYtvWLNW4sd2zUpswLTRHcyXHz/kFQnqLg5BqsA2E5m3TgdgFgo/w2C
wprpB4MR+97OEYlZaMH2nSC7ajDle2Sx7KGgY3Y7nqZkuhGiujFImVVhMX4ajeij
XPDiiCJqyH8Z36YsosZolSLNGrZBCdfckaGliAwpYwS2uPdnmrteUrVrT/r2iA/V
4O7ZKbD7FvKjwCjnyS74QuM6r+3RuEJ8MQLuVzKxZN78LrR7JMrFes/VI3WG1F5l
L5MUGFj+NYOMBPOuUGQXP9HsL+d28r2903LX3qmJyz/RGz3gRMkMRMnR5tRAONej
qGCIdEcsA3gYQHAkO59R3Ymkslnbp8Xzczum2jKtDz+EYvluJmTGUt1TqGb7OSho
13XQfKPHmdnn+QuyunoU9D7mOncOF6+FNWBpxIXYR/aFOReY7kqbTAj1eAQUj08K
TqBlAgXKzHE1+qX/CcwZM6qSROUyueDK5IJQBAbd6hOkVhUgIkXB6mlEfNILZLQQ
+ai5XaT1MMyNYvFJDsmNiH1QLf7hMnK1gP7q2qDAy3WtHk/BzoT+P/ZX3SQUa9Cm
odwoZbLeSZHf15g455G/dXNALh8CIGG4G4S5yj81/2eHxI/GFsZ+Q/v4ifizv0J5
CzH60WndbKY2Ml9tMS2whIrK3ohzFfN6jxNG4e7528vu3nWwDxqGSnGs+r4E9R9l
zsL6qyqW6nJcvkov+V3tjc9IYTU9hJUMUmwbrhrpPTxJLIex2K6CfxPcbFEqTgxD
Yu3/LJwkWMsU3J2mtjQtVBGEwfJoUH8SdRgXb8T1cqayOY8Kl+kxA4xgjb80CF3F
7Dkk6HW0oq21d8DVwJapL1fpYCD+TfgYg+1vLIritaKJRmzxz/EXPqz3t6I+lU0h
YxZNzWRDaY0CCKm/2aMgSzEiweuOGiPH9+UwP+AIXSa7a1cV9Vrel5hlJnhxx0za
PWS4kM+MuC+vwRSkBV1X+mM4K1kJ7ACJp2KoRPRwc3ocTEVkkBRxYPzcKR5oglFY
7qmSvCeXazoTfaJlK/Or4EiufDP+TeAj8QmVc5T1c0ti6sAaJRabDJTM6neP/ZMT
EmtLNUm5yNcAOrwMT6ffLvy3BwODAERpEZJlYs+v/CvaV/Hb6LF2o9LgxseLsFNf
4VuqPY84eFKE6vxc9egbDDWVbIQb8XhBZLdP4pQOqvkqG9YicQxCPvpltDT8S0+z
vnNunCPAmIEZ02OzEXyFe72o/gCKoQ0e4cfufdhZJL8xXW4m4Ph9LzspzWiYlGN5
5oCCj4IvVx3RujTuSvpBpcygU50bx6uG4atyPNuAWxf2VIT70A4Da2LA5dexsjhM
oK3ugzmsYnS7wk5Iwz1RHNgZJ/87z8GC4FN01YOdMXrD3fSJv7sv9yw3SURi2E2o
CnMROO+LaZkrHa+dgj4FjEUYydp+m4lkw9yqiu+W8MMgt6MYGSgArsLPR45A+goP
JcQA2wSn/m5xE3d6y96873JM8nDcDBWTmrHTth9wbuJQ1RCRjk6Mc9+ZmirtnrAH
An1AwawDd6FHpFny8prgCPtXcZfL6aEno9/f3yd0ViWYQBMliTE9PR6satDrPb9q
NL5Q0L2qVVZ+X5qcbQI4j8/mZWcLYbnYOEwLXdzNE2H6EMXEPSX4i2lbNmtBa0Gi
0Wxk2NEGFV9QVkJ/wlalLUDeVVH5lZ+KvEkQtJ83cDNI9IuEee2ICenkQAFeybc3
NHz1vy7INwEhvvULHEs8tk5M1Ay8kv37wjihCa7FinM4DWLWdzumf6QxeVll4Ppx
/Ypj/bTWDzJyDbYzes4l/pJMgHAKm2kz3C2wUGmBSyVGVTN1eIC6aNioXXkjdyVN
Q0qo2dOAe8gU63B5aeWAcUhtWpk2nvhGKqGb/ANQ2UJc88/sPAmUYwW2dtishJky
vvELt6GC2jkZf6nPnLweizzZGnZi0Xe+Xi3bENbyCU4zRM1MrNN2EGaVhmsJaYR6
vaok05XS3z+QJW/7ih8s3UTh3t7g9Tq0ccCo7OtUhBbZRMMvUAJNQJqKFO7KDkNl
B/q+D71Ar2TeZ9mKm6ZGPJkeSRk95Z07zYsHHExfwPYD/cHF6zhbheVsmAk2doqO
KXLQ1or0R6Yv80CVTfkdGIHUZB33AkFo85T7itK7+DKyT1iEgG2Ri3ngf0EoFJoL
EZ4P3KB4etRJ5wvb748vOoRyrhwesy7DkzWMf+8l6LzGbDcGatruDZR9BEOt46od
LxqSrefX0x15zRMvwT6HSUar8E7c4mjcOy6Q1TlnncRHwaA8VdxxY80nMF3gMKWl
TaGXaS72IyGYeKIENb4lG1QUk0mLfKlajPhUh6Mhja3YZmV3mFLsCx/7TKBos6gX
0gEyW1YkxYemh0eAmfP7h7anRHOIOH8Tsg6iICiaZ21n+QzyLX+WFGgLsNulkEeE
w/PlCTeSmk4clwo72asMBf66oNsff7gVMVVvYEB7NdBBZ63ZpeitiWHSzJTA93kW
vVD5gUQy/lUlTPAZWgeIvvk6b+jtZ90bNj1adIRvcBT8zBib2XxfHuA0yYGb1013
DLwx6meBIVlGIXFS+AKvm+gwg97v1vb9qG7Gtsf27i3f4ienjzGEob8p/va9hpT0
5U/qlKeMemFvevCmrSSbL9/D3UOmpDeU974VLRzqJL5i8np3Cklu7spM/MsIE9xb
MNJUZcPUq2xbYATM5yVJNdt/bvSCZ/rbnUPF2wUAvLjH+D54QHztoSABo99ZdDZT
Mx+nbKaAHx9SLd6BkBTzD0cZ5RQxSFjqzfvelYAVmmj6h/2yufLENWCxZ5I7UAP+
aLqqxgZWHNt1/Ivqx3/oZB4svlak8ndc1XAckvk7EF4r4ex69N9k6SwkU6IPIXmU
4gEjxXzDLgu9gdXUvv4kcuKQMMAUfmAk4SSHABqbQZQdi1lDij4PXaH/L5Sbjq8g
bEf3FtsIF9/02tZNHAK+WN0theZlA9nN4B3LXLSzRQg2JOrFbxbS3kyHnvEJDDpp
7WOecPhi+7zwmZiZuySJ+VHMO6y5E90dl7v2ug6fI5fyBXQfu5kFZNA6lUXxX8gN
mwmiAU2elu7U+GPWAjovfDcGiMe/5Q6YzIyIXaUShWN7bn6dt0QxCaIezYFJKjG/
Oscq4ZW9MR4bTL3bzvBYUIxR6ydtUjQI2ILQgQ52vbY+BdM6MYJkXgq/lAzYimdh
kzZjPBZeRXL6issUoAW3+bOZSC6K23oAshoKkjomQwf1/gubRBJ2AQ+t0STa1v1n
W5kiKnbTD78sZhkCf9wq7wBQB+dJIDOXFQWAIF2xR7Ch8Ho8XK5eNoiwFBLIWcbR
Bqe26+rtSq6EV6RgCHc8m14rR614emAJDzO0hQadYz6GTCKrVUSiy18646U5r0+G
sk1l3UXGUHSqeP7o5N8QE8QtqiCV/BICPJBqZb2mnAizsKF6P5txE0Grc0CrV11z
cQDSzahMPQ+SbszDY8etInL61rrQkHNAvCmVrvNcI0q66haocbrq+8wbZLSD6w4H
62Z0KvncNmrobEAYUZ9+1LaMMbRv2Gg+rYgkkrf8IqPL4mAkZzXhItDCUzeQiY00
li0F51eEXF4Anqhuy6HpwPcNVmZaa9fL02DJYIsGe58kttp8dfhtzdMUgBpRxiC0
jcfEOaMdROIKAdF8NpQKACCSEf/Apb5BILgDfFosLiIt2Hfr2C+xY2EkBHXArtuB
wm2naPXqX9lp3m7lbT5CpI6nxXih3qaQ2UhgTgLdJqS56mKO/jTx4/eRIqVtV5lY
YLHkv28mfMHOv3tb2BMptFWOJTjr65yxNi6OacGmTGTnBdmBqS4705TIJ8bU8LDK
cVzHdT2iBarubU307MJOxH1j14UylPamVHWpmzCKP6JF8uPMmImbJJXXOfhTolQC
fyoABolknHAKLn/o7aGEVdAT8CcSBgjxKlXhVnhdUCNdSDw//MgS4NsRGjTcipFj
E1FyIR+wWjPlD/MavoA9DuF53J4XJjFxUXME3F67/kb4yfXQeru0N1Le9MmQJIIX
CHY7OHjEGmfiDi9fwBSTpOph16XAjrtqSYseMwlRVXEJuGuCV7HALDCNgC+OczvW
vzfZ8O8yf50pdOzPCmCMtETdx2RUElxYloegEvFkmLADYl2ZdGtoeJVu4bPfhBdY
ZAAqjIfxZ91dMsrqkrNSFWCkWsGvUJ7u91Eexui2b12nj7epJQdWPDJ3DP4Fvrc9
TnSv7ODrtgDC/SyofKa0PeYcqlQ+jp7FwXpYzdZR7/aJzp8IxjG6SugaqnKEwGGk
aCi7w/OPGakLM6BibUa6HBcLHpS+vX+YY3aZ8hNky5cO9V/n2Zq33/obfD21Boyz
vgbuK7YNE10wjyHGirpoD2MrFNA8G3zajy4jKyV9VKDRBf3RcY+kRMKpk4xDaxKO
D7M6j88SyMOhHaG+pOEl/f7Cb0+m3LEi2tOED5v5Zze8sIvllr9FD6zQ1AvcN3Gn
GSk1Late9zKHI62vqTsC/FnVUQ6v23GJmQd6JooNyqsGs3jNtqRye+z4Q8gEwIt0
gBtoV48pZcBspcCVaPv+kKS8gbX/hLcqnlJiCdt6PG1omvJWfV9nM4nxyxWb5kAr
Ru3sl+U00FZFSNrI848KZy9FbSorV8GXzEj4F4V4bcmiVHyI0IfqZahu5V22TnKr
6+mRjGzYl2dqAJOrdyVjkzsZGqL8bF22UCnQWV70SHhSJAnqp+bHlX4/36OrvRaq
pPRcRju7PzwDN5SPxxACk0enEzsLFaTbqjdwIu847LamoN1gISUss46n7q1fwPws
tXguEJyce6+WETgkaLDEIZo/ASxSwjPyVGA7hr9EfaIyzPOIhAj/7yoxvlrT+vjk
8198MF976TX9TzYLTxHitIvl65AkvBI12HpcryevoaLpM1mUgx4cmE01cQeAm52/
c0G0FGz+NcS0Mvvc+c2rkrzydMhzADVJF9xVPoNmJwlRcmhBT1WNprhAZQUufP6R
/NJOz0lIg9SM0KYKx5Oa0aMypLFTNAZiPEQcKU4sbIAA5Vn4bXjq9Z/8NJH14WXg
wh0RHnhxAb6CiS0Rxc+WZZzuzazkvMEiH9/ufz0QqdFWlXEcYY6HSuUzAofAn+Vh
ki6N3FKa8q8vIrii9LUVI5iTBBzUnCMCh2iQG1l6+eA4zK+y0ulSEEPWV3xoXMr6
IZxKHn+fNoUk4oNcwimT1qw2JyijVKdzV304QLHKFq5gOguNN2C89wF4g5Y6NmjR
QAB0+r00HUgPP8UITUvCVdQg0gWtxO+l7UFnbrp9F1p1m/0CpZEZ9NWlEah0vjI5
L/p4JVMyH/C1m/E5f7a37KTYzgoYxWCSSbfRLQYk6vPGC9LBmIdWs9QtAa/H4QW5
Jt9xtZvOQuTINOK0/1rkFIYfnagFBYgl96gj1sdr+SokFCX4DlT4WJToc5DEdxvH
H2VHKYE6h/CWY3nI28jcURI45rg+X8FGGhoEGONfMOkKKYAEMfFiEQMpxGczzsi4
5033TQZZ5YjXlE8l3LU2WEYRVmVj0IEY1x4VnfjtcCAgpccbaTE3Lzu+iX2qzTwJ
Hq9q0/Hr2KPCGtIbqK2RTg4KXU/u8hx4L4XL88ptNpd/I3X0dUOQgZtj+Fxvsw4L
rr5Ur7xaUPVLUHWSBubfQNGhIKUjKXOI+1ov7EOht5qm8gRmdUw3Vj0VyJuGIXFs
2dVuJFl8mwIverYgzwzTmMSESca7C44d7c5bH8uL66b7tuKCSdqUmJlYJ46dim8Q
cADYoM630HCQJZ99p5c6g8kbhIK/AX5C3VjnyupZdmXdsBOBN0Tg5Bo+BTVHplF5
lOF/5WUy6yyjBJkucWlmiIqwPjjFxruCfqQ8zTRR9nKCPNtBmtRXmRk0Vad8Notv
c28xWeOIhLrfw6gYWYlh4Ph95GK8BnWjkqWmfOZo0Rlk9fKRZzPuIuiBvILS+Mxc
eRSQdpDWGZFGV1hrtwJTuKtrhrtlrGF0MYN0ByTRFimqMdiehfCdMlCd3rDThFmx
LyayMoXKzgmvVIkF4stFotbZnZ41Z9ihmJWXb733JhNGwD3McNvQ025zzC6P4663
MMV3sj6NHeuJ9Nkh55qTeiFrATFbXONlBYeLqxkcczZW/OUW+ilpX4K7dm7hdbym
AsHcV5WIPGIg+8vTT24G+V1Lk5zPZKToffVzVfrBL0pNR0lwJMiOFOp3ftwN8Phk
HsgiUrNLLntlHQIP6Qm9Pzb6yYT3CNLVQJ5n5XiDiZKCiMY6VnVmP+vcbRetByOw
hcXYBkM5LiHnWWGT4qtyOBaYO6BJC02t7VQK0Q7QIn/xEOU4qtZf8wLZPh4/Yoif
XmuRUXSEKCTlOkUhCwr8Y7CKsRoHUJO/BGwSahk4vS+MjjS3reRaosrfVsfP0taX
GbXFr08AA6+BgVeYwvb/k03FV2jVr0POAHqGile70tXjiqgEsEUIbk2kP548poyU
3y0JXuiHls3LPBs1t0GBY3O30Kz9TDrXKmTaVeawXw2vz5nAZkdty78JEEZYcTJG
F8UdSx8tEKkwpj01jQ+kUwZmfhg54u5+xyze4eaxQ5OBBOoaBjHr6r3WbRUtRwqM
oX7JAN88dO+31mlThZczTFO5QgRlP+lgND5zqtxWD60eOPsVFhQPmCvHmoeaoehM
GJZ0ZWVaMUHNYxJTJpPSKfLPt947zGu9yDh0SDkOYKzleinNAz6eI8InSJLA+LVz
wb7MOcqeIlFmau/xAXhKzGkbZkCjou8l1hxWZwnZP3FWF9lli/numI0kYMIr0DhY
O0ZMTZP7SD8OQlZK7Hg19pWC/IVi0WiUMM7OpECSHptYf0RRZiwOULHFy0SKABEy
FaN0xr3A9dC/HLxPtqulqQFrFDlYX8EG1xmqLHv7KcHbAWO0+NJBiFhL8we8NU4u
oXeeknc1c9jCWiimznDX3ryF7+sU3djC+aBgE+ltR8CxREzH7n9lwz+KdUhyMPmi
5Ie3eQlrwXyxFmLS/0IXxQyIZq4GZMfbjRj1GUSEj8rj+iCw6TAgY/+qZfXatcsW
XHA/NTmaSNNHkEFUz28npLXU0IeY2Ar1UK3YqZk0qutnWBZLmbz28qAQ1Vrm3pnI
JmhvSNAtsbsGyGPJ+hMus11N68jtIBeJldOewSU9w4YD7qgQYYccahR6E+hF114R
L2dTHvPWetlCngrNkUAap6OmUHoaeLBiPKT4zJ3rFCbXzWgM/FUUtJzFa8kfeeT6
ytfhkW0B5FOBhkFsY7U5sr/3tjlcMuAYKQem6wGmO73wZKnbVyZyAuSUTx1K1Z6s
PDh37dCzCK2bbQV6HWAbpQ+Nn/R8XysJg5QySV3xiTVbK1w1pY0YJDwssh7tbOOM
taVAGG7+4noMhng2+L2IHvl5bFTnyf0P8Dx7Ig1WcY0rZ4O6RYMIfQhj5ad/aJAH
nrqqMbdIrNEP2LsNE48ibchq5JYhlmrPNxalayddXuhKEsl1+PYsssGp0dKfI77g
pdIh0rngjfqJ+ULjYlgVopvfw/++m4BXVrMpEgjS+0+oja1frroziIug7+KLt+Vb
jZaX6PYgOq0zASwygVDBSRR3yp4zj7tjZ7dkMEfudRWsVZu9gkSDPd68dXEbqAkV
fk9z4kZOT95XSYB8GTCFp6i8HnsPLkObTxVzDcxGW25yzXpoQBVUi/ZCt3kIQGjM
ReECaOv8qsDKYgkZTkx4ritD63My6yKsHiGTQz7JhvN/Lmk6L6tkgaMWTKblrB3K
+gyyJiu0gTEI+nFyOUaFxNmV7R/aZFdHblmVy1aNPeeuVAISJzglJ7hW0l1y9zrg
reEHXv+VtjL8rz+nGX+bb+d4DNt48WGg+vZ6zDtzHlNBWZOeXV1WEreohSgHK72N
z6BlcERObGG/Hn956KvVMKBQr5fJtURLPtKq5z42fAjGAxSeeuPGNFbtLWmc75VM
+VSb2O2pNdLHRUK+f/1I0u0p3u6h8Rb0aYvV7C8SGXV0J687Pl7vz63cOYCzdWtp
peN2TUW51EpAKO1BemRnoyPtG0vQZyIjt8keZLAoTtMC7uwkphsGo0/TCV4Pmlff
4OlnHUj6rksGjRQR1bNOVxw3gluNXcCeIKos/nqYImqiE5dDGGp6gS55lZD1o0EJ
WjPyRsFUYmY6AGom7t3L3A/iIDbBs8V5DgCNlYhIusToLbL5QJRQvatDhXAm/+/V
YrTAYhAfMAe8r4RKW7XPQ9B/1TQTrJoUfkngCZLGQacdNpRd5Rph8jb4dG9BwhRr
hCgfsS3NplC9bOCXbdvUBlMcBqLZxnek3rKNKnl+QrN5r0wb9beGXT9TxUCL+QB+
/vesrJAH325L9AjyCqVi5+UYQSIK2ylk1Acb+P7R7v9V2AaQja/8jbDT45BnrC16
l6/1zvIZmWNQPM456NgjHLGq8B81OzL1v+lRhszWgwhZRMHhRW2Hx1YR6Wf8vwyT
Dj/2WGcOf3n81f39SWecN51iF5eQh0FjtAqRkyvN35SZY2XtimVfUNGTwHUX+x3p
7KEauptpuSD7c9XyhISZJWIRvDvHAMRDbknltwGIGHlRp8rbWbuodNtzSlEuz1CC
1Pw/03yeze5kTabXGnDc2/ofH0CVUyImE+eaCjES2n0FRMqiFfer5fSubQ3/TuDb
W1iVDtyvUn7REFSVNaEBrJ5+nvIu4Ifdkcu1+eJSsZV9Zzs47IV6sHNMHs3j4rB4
330KWTfadKTa2NrW5RZpulX2pLldpNKARjQRwDBdFBkH1fumMArR01GZOp18Pz1H
M1+3owxO9+8aNk91mzEzuAVr3GAMVR+0Qs9/1rmqVB/L+wpTv7K0xxTy5EFqbdwJ
H9fG3wftYbBHz8EPPoBp+4r0xc0YWLgE5iC2PjwcjMT4gtj3RdADihrnXAqSRlPa
SjgDxRm04mGxmaB//lnMIUiLkfB2zi4ZD51EFh1cDwgz+YJ6sGcLHO+OljK20GpB
IzX4uKquPBCD6etyEdDnmiRGUjWb0A/QZe4z2Q4GS2LGCBgunYBOu9UCUFLfYakT
OO1+EQgbMQ/jHKtMZ7oHXuT4Lt4/EVcQHTeUgDgaZ7oLTZM00YxRPNr0p/4za2AJ
UTBOBO8wIBO3oTAoxTR/P5JGQEMExdy5HfK6j2BoX8uApb9aAwvH/3YER1gxTze8
r/eIQuKcIgKmYamngMFxLo87YHXetO3t6ipWq3iSlo85aqh29dVbnA0NC26Hvy8/
w1MByIc9Rao3ac0WaUtvpQTPAjjVYk3GA34wNK3YAivwK6Ty/4bjikEJBRLW5s8P
F4r8WzaZIf7YX3axtjARwSrMOAPfWRz3Qlmh+VhRR/Affas9aJqt+G2SZzPQ+L1Y
j2XIRZUyX1d1pJ25yEmS+Z2kyr9xy+ljAl+6OtZ6sdAByGwBr61L951MGNPK5I3P
+jS5y9mk6pOLbvJqwMdzcm7CWw+Zzz8Tx4VD0vfK1P/VkjLOJM8mbHhQ94nBaz7m
50EUrYOS+WvA3zGWt2MUTq+H/+g0tPkrgl7OoNbcGFRDpOJDCBmADNKmxTis7qH2
aJ241AJt5LiVBTPbwxG9xOJNrYGtVrOSbkubmz1IadklUBquUPg5qR+5TWOMbHPw
IhZNjXvO/fNt6Y5KMVfHnpyXYa2JsgnDVQhEG7rK1w9ETuOHBVmN+15OzXtnIlE6
VGi+cHupVyO7QHmpbIJyPo4F7Djp6N/xS1vy769UKuPSC3pJ3CYEF0A4dhKF341I
TTCR+VSZmLgv0mbkejFfdfLaRN3nHA5exWGPZiqy7V3z8GTwyJTtZRM5CV0jqLA8
4J3h9MhYDizzeBANTWp1a2c36IvBQpfYWGIBGprQW72kwrnae8bO4oNpnBM0ywSp
8HEe+QXu33ORpImVVoc26otorfBO6kSsXXNuA5VWb3WiGgZjx3IUvfUHXx8SqyKQ
3VfeK3TR+JD2jzVmlr9YqBHb18bxsLVuha59zyC1fCyGfM7nhVIxA3vQo3DvXDKm
p1eotk6H+RmhrlrOFrhUWVATuxqOKqrg9ttudmoBXoNDJjWVILLUYOBNQySt0Je1
ZD3OYFtjMrjClsb/iiFMi5QsErk3ijmL7TIZgTT590YvlEjKGS1HbUzqkKeoScND
jftjj8aR6PO5KeQ23yylLyR3osunYX8amOUD7J+LewRjJ5TvIOa5mtzZ5S6xzhsR
RP3Ck++yvLE2fBQnGgZDd/IOsoI7sHk6ecr+RfT9w9XfvlX8m9y+OjctzslX4V2n
EUZRKuk6j/yOVaFguWz9jLHQF31EfTeGjaxktGxahIXm2cPINuNMajKKZLhmMzYB
zYyVdir/M9cN+QR82K6y4Y0JVwtqlf/lFTnKmhpfZlx5yhMwH6FZ+IrccKsUgu8T
UIaZMW0eRX6PyZDeptjcUugy1PPrxqMxnXtBWsNWi8WXR4+Nk+EFmokoGtk3KHfJ
osujbOU/6wlZ49mbBAUXDY4RSw9q+YFva3PgNlCrXevbgwPJULpQ1DjQNO3/nHPo
1ROOxy2+5MSCHDhCHgxhI8m+RRmIoDanExFGmaTgyGwAqnYTJpo4N7i2TYrhPgKz
Bfo51YsbjsQzDQQ+Z6K0Mh5Zf+jmhcjACa5aFv7QkEcNGoo750/zZH3f4LRmqcV1
2hj5WYj1mCXssZF/tE06Jx5PtzDTM44DPTkzKmiZS2crQrUYBYX5SIn/avtxtON1
My6cZPARRnxFgr5ic68C7+4IwWG00NOdDYvsOcNePKSFs1IsYRDuHK0ITOwjTTHZ
U2BnMhTASi61G3bJhvf5WWNYcAnhH4gY9q/uLVsaY0US2WCnjyt6HJlJWnREkgtP
Ir8DqSlxxmoNHOx+YQMkf4vKRF6O7qVVq/YwOwUG+tnSdC8ZIDO6jZbn7sHdv8A7
zP48/+XyiPtdw4dPt6NatyWP6YHrA1BughcYixRc1omezw2XSEFptgjTwCigaJnQ
RHk2Ct23sIhN2AOXWDLxukXieK4ir4uyXrsMtDhslCfAOLdJ4vu+Um/vxoLXO0sY
Lr8Lf7L1uQzGNL7wVr7gOr/AP+hX/nTFhAwoRfPGoXjpCNtU/ERRAfC1flJayKcR
XATdDZqq18O1GyFv646tXEQfrHtqwW+3OqbnfuE6YvgrK/PI65vki6fnwm0v6iOK
D41K/quOl8SggukuI3TmeqBwt8l9DKAZ0KzlKrgyFMyvEOaO4mclj981hqEQl7JX
mNSd24+8/WyNoZh9ymILO4etVjW5BpZvUsIVwD5TNWaDp3hlUN2+RJuaS9COf0ft
6Sx/ufuw/ydRlpzra9Xq1lubSuCLW9SQSthHizEVKnZu31OY/74cdUu3YRuV1L9S
RcFj9bq+/+2stiQQKkSwwjZ4WFGQbZvCE/pxi0MgBxOZiCLEomLvAhYt2D3Bg+Hs
yfAKeoQ/O17oyE3Ob5kPHuSuG4fNyYkXZFUjStg8N4+k9a3W3e5cPe7N3lf8OcC9
3tGZk+C89zQXn4aCXbwE2DuV5xWuWZ1xx7AJLRelsFu3dQgovsE8btpb+G6SOB0n
hRffEztGzLYpL/nXI6i2xCmYQeaLEOYguTH3j+utYL8iZBe0oHVC7zOI3R3zK0hE
oJ83n2lZ4p36x//bLRRJVG3noB8EqeOpPBNowED6HXcDnAVKjHafTXvFrylmfPn1
eA04oX9iVoW/wuA+mSIGq9vxvo2V7WZQmuuqdF+l7Q82q5qagRcsJvHeGjOgWycM
MvUc03qUBUwm71Nr7Ur9W7I743Q/qs25nYQ2cegJ28ALeOAWzLZUCvXTcjqeQ8+N
eJiJZxw2hw4ZQxLeu31aZmDASmvDCbju3eGEaFehKxlG+4GIm99nd+47RI+UBIkd
nL3EC7WB0vZu+jPhOmnmvbH0FapxwIf6oP6jPNsqU3wB5HlZ0JHJih3u1XrRkygJ
1EDDFfDATXjJR8u3ZfySYTS9dtUM/qJ42UGKt1silvjcoA1B1/kY0CsFBrbnuciJ
GyvmfecfzaZbuTCRqb8Vp92tyxdDqXtPlrissVFw7U2Ysvmhy4qq+63EJR+dlyV+
gXg2DXZCzVDEKtrs/ZjWsC4HNDvXz0YNc2cIa39XJbjnZ/cEfi8tkhKOmITUaDUH
+97HPG4ZTwt+YHAQX/HIDEenxl2v1xZF6is6IJmXBFaOUXQyhfh2pB+yf+wvDFOK
KqqLaQ1g9oMQ9xjQwr3JbzPPGZboX12QRBg+SkQ0F0sxpEuENEv58+YtG20GzV/X
4VusaAHD60CUPd2N8TlhGM7xplYJSbo1e9bJnlkvnKsJIvyzg6mrbT4n05pipjYM
EJ443wLTy1ZlWRJiWMkTN1xEDkEyysLpHfF272Mc8a9lDLpHtpKoiTivWwM9ZEoe
pfF9rJs7brSeCfN47zUfLfroRkAoEUbOAkD9xhvJZFWPW2xPcJW4k5gPgJAoJKKo
cprDjQZBrjqotbmWi9RFy4irMI7oxh1IwIS+6saCrhnGjstk2P26JfwdyL+EJxPS
uUX4oOFgSO2orirjUYql3VoEGtZAHRMGE4XMNaL+sx9TerBzaI/1XYGjzFUihsij
lIHasG+wp5BytOkR6U54JMEjyHjHP5Lc8BD7nMnMAPVqOOYATuPbDDqrWoKN/Q+U
IhosZI/RyjnXl1nf265zNG7LEob3hk4L8Q5JIxYlEeSUb3muL8BYO9kHXCPYlV8V
2FOTWQX5h/szm3uSVHh0zBSzaoUVO56MZmlL0Jspc/GAgo2RZVavyIE91JbpdHU9
NngKGa9ADpujdaj4VrZgmUJL9wbP1CLzEgarasKhpoSfrrceM41Hyd8WDtU/HE5L
fshbNbpDgzRc1y8CTMhRothzxZENv4tu1Qe4zILDdBRqtnp+75rsVYu7eS9/IBoo
ixa0QtsA1AWZPJagLXB30FwwLpaGvUhZV4fWAnKTwZXJjUu7ADxuy4iB2WpIvb/6
8S0mKnVgtLeejGJZRuJio3kN9yXgndIqlc65xiXoisIVhJ615gen8DB61e8rpRjC
h/ZHnUcShWo2pdui5etsPcbI2tLw9HGg/sEXVCU1DA4H3470G2Kw3DQZD7fBUi9i
239KwNqMD6gEJgh//S2Kj8Mc0H3a7YKx+mjFtERfnWx4DwhexRnaTe3QS7cbtbPt
/zRzk40nabpB7hu+DxlCGe1NRuR9YItHqpweTTRj4DQdh0gCSJhoOBowMlDTmXvd
bBJBaY4wiw8lpQLFLZSmEM2TViLzWMb8zeWLGWFIx2FwD0eGCVZrcFvIPF2217sC
S3YmNOUnAzlLMLsEYRsDG4Y/2Th2GxnisLPcYTx6zYKSCEaRmsbou2QAcV6n0+dL
Sxlpm+uxr6oLLKl5xxRytPafw2erLWa0aF+IVA8OqWPwdSaS1PpiyS8N9cXfSxKD
JK85McVlgxrZJh4AZha5tJocsAMn3huKrfXPD0Oqghey9xq28dMnBnKDvHIkjJ0c
tra7zbsd3003DfievHePf51uy/2QnUThezyHYWFzqdFD3pHITMjswtMfbKqa5b8T
HF2eWwcVt8530pQ35DdzNnBUquTyhSq5/pLnuEN85i2g9oXc+hRGT5e2P77oPv/3
C9wItuYXfFPML48yakH/9Z/+C6MukToZ20T6nCTXgqSFihykiWkKPrDpRWORJXFW
FTr6w5htSWslmikcp7aZqToyMxXSjSCqlumWjCrRmmIsb3VQyc55iBaEy8fuSGTs
W3ii6yLYY6rM61pzESB8/SkeIxWbtpXwD71aZbsVEM1/NySQGxULuDOxCyg8Thb7
TQPrqdD7FdL6o5IxJmnq/iQo1Ghr9ol3+5DQzeihvZxnygm4ol5+Obc+IzYOQ0u9
b/A4aquY3ZFJLGVZEr3vvmRwYukfcgi00bjEDGkyVh84wnPPwx3AkaW7zPywHyzV
BP13oT3N5ZeD8iBmkuPmPzDEbSVTjUxNM6b60hkKoq5CFE5qCw3F3zuOQyu9kC5A
T9zz+LLEUEuWodY0fC58t0gKqTz34txzFRX1AIsEHqZQS4gBRBj92cRS1ZD8XZIC
psBx0UfWA+Gpz5UDDwyax4KjXisPfgSG1K8ROkiYbgpEtgBvUsI3sSi2BhXj+XOE
aT6a6UodPqdbyyd42FVHlvzb0dG5hyEPd7kKHtZJHmJ10HGPFW1/2BtK+uDXTTUz
0L3cH6vDtRKJCwanO5qb5RNWtFebxzUOaHQ6//cK4rAyKqiLHC7Dr+oq23I7YnY/
x1gXxMhE4LsRYB7aMniQNQRSSBRgsRUzwokW4DkgVFptbAPhNMC+PStG4PZ0fnN7
NCt20+fyFGbWCH6WZhWY4HhvTxO7MFZN3UURrTkHAG2Gu3tVuz51ZDp5C0f/pTgK
DgM9VMTz3t7sE4kFy5JqeIX+s9lokeI/9kgJi4mMXsj88g4KvoUso7CQb/Yk1IxS
I//nlSvdvgWU0mt42ls/G3FC1Wt+O88anwWYKINOlXXb57vp7TtdxKrH3VJRqpis
RCxd0C4m9mSSVK6BlDuX/86HhYMU8KMyQcnIRQUYWQtFd7WvDk10mZFrs2F6oWnK
3fiNe+uLPXuBwxef71+F5I5JugGNhpnESShZWUQK5wMBa1XBKEJ9c8ARmX1A+n6d
ahO9nvDOnfypARzl/6UWpZxAbVG3bQ7/zg+l0FiuYppHGU9pjcLvLLmc9psyybpd
+fZi/5mZzFLURLde0a4xj7q0PBb0B/zOctkN+/Db/v4b/gufEdEQJvF/exBbdIgR
w0jLzlxB/pht9IXOhZs3JnJ5RCLjLQFGpzTJTw6aCCXdcLNX10vDw/o29jGwfrrz
Cvl4h0hfa34xnMtVe9Ke/smXMiCB7FnWIBHDiNWA17f4PB03lsrMumLhN9+dSpB3
CCpF4ipAUgU9Mn+zy0JZiCkMhV9XkVtiGFFuPNYdXKEMsnU+n0T5JSqYtRB+zprZ
iiM43bvWvaxUDPJzlxvNm8epMji1DHKJzgxy/mJREI+aVgFQewLwekxDBzbTVsrX
p/undd8G/yudElbYIHsV+wPniehhhCP4LREYOkaLWAd7j0ZB+PgbE/eFtElbxuxk
5UlnXJDEnp6zkxCiKnujdWIwU26y4ZchqQx+5CYuK0GJE0/oq6Xn6UTmmzLeHZG5
FySszpEaR8L67a6W0DCo6C7H9E5eGAkzV3HafwGdOsF7HuCAzGWK86Z/2onK/k44
JdagZadSkGDUt2DDTLqIQcHUlOxL6KSxi3GxMsg87YwyIqkCe87hbNb1NOCci2K/
OoCeSaQzzHpbITyadhCrw/aqmcgGqYvWdFBHiSyABg/vdiOKP1nZ/P+soUQVyct/
C9D27CMa6OozU6qoqy2vRs+JFz/tOgIYhLlCFYQDfJi2s4Nz3IGyVPJc+vOf1OXP
K9Qg0AIG2LZVJv8h90vJszFxFzFB3ORa1U9/89UP/Owi/Ius3a0ZUyliJVChLq12
3U+OFoT8WuwJgPjV8F7dIUjNYmTo/7OtdL11HqgsPkaVvl0ongmKkJTLu2PWrcv3
ENix6rVbji6X6FyURcSF9QZkgcWvuBW2eRmBEjf0XN7DR3CwrLna1VR9RqLRXpUP
5Ex16ni63/QN7AE//korcwNncbFk00gskpaBgpFcQNyzapfFvkwbPWKZAl7T8n1u
CRYEg35OHOlJiVv5bEf5J4cjk5xAoy5U6Ue7n5wDPYbbLbVa3LzDTE0E55ITJBwg
u+SiZod0Uy96dxZ1Kwqbyo6hIgD1favuRd9rHUel1QBkIujH9KOeqA/8yIF4R+hd
Pqtb8O1H6LX4Vw8gRcHnBx00DHgE2JBNxZwJ59SOhFow8QmBVlugGzGTCP+2WZ+d
A0WXADtElYLlqOkQG7cWV+C4Ui+KKqcDJL9oy6NhEitjfVEKoVVPHoNDkeUrs/LW
Fo1/1Z5p/Tk6NsxNBjngCqtv3Doa4xy/x9AFHadQqP3SDqkAgje82MfDN6rrn6Cg
xAZUe56B2RBwtUpCrHKoRsJrX1ClbP/+F/QGCwdZn7YgIau4CbH37X4wBUpvyry8
TxJyxfUGW9inDO4GBWC5XQ7XMIiSCt0igAvRDS88+vF11YYlGCkD3Shr7ZFSrRBH
9Hz4faOBqSRDcoUHoKAwnB/yHE+H6TH06k5yHK8RCkSGZZUBK0D2OzJkfB3s3BSL
BDaoM3TyXOq22Kp+TzgwNY9bLkgTDSS7b44dTBiq567yCw3rMUvWUE49dQ4FPWKU
QCBf0rGJGQQ/UAecsIPLJ7hQODhS8MW1AOzfvROFANNzvz/6vOONqR0PPuW3BMPJ
ozg0rWxgWCnLE+H8bnH4k1PHx4D3t+Xz4RMNlOgEV6VYMGf6J3SU5fwFm+uUBCeG
VlKVKTKpr8jFZCAEjkW2G1w4BXAxUm0z27HGJ6vbxgGpInuLHgJTBieJjeBaA8d3
lohu9OE7gjNJGXPZ6a6QrhYD+BW/gTyNL7jhmqu+Hm/Qk4rwVWgDCrVafNWTxnX5
WpUpB2y3b3hj/U2cU4a4ze781G+n+QQfYf7wfcsticdl102YSILdwaCybtlXL5rO
IJI6cCp8rsoV96Fr7xK+/baRPujwuvoujwnvGZ9c2cy7yS3AWpyt5m/lqwl+aByu
9b98RGZ6UNlhSsTciAN9vtS298P1DlH1O6HVb7uGT1qHpufyG0nk8DcpjrNuRSOS
MhFuc4pBCpxATghIPlV/bzFUM6ME4EouP7D7b/yL3QcEbxv7WXeJ8JNzMDDshngH
rJp1pbJN38JYnu+OJQzutn5rQGugVBuh3CvrTrf+BzAMj97EbXdtGpndILNtd+XI
e2SODjXw2AW9VwHb/EjNJHhrBCuz1c2PxzEHF2a4PYLy3QyZcIQH+XgPjQLa96dY
xXYx+cWTrZkjRe24UVCSuewJfuxCH4qCDdxHy8bQNt3N5oA2OCYlBGuJ8zgVkRBS
gnbGeyMZIK2cJ4CzdJSZgNqxO7Ed8CNAOh0VGKY8wJlWrxM02LCfSKTBkAVdHVG+
sbtMKbz5lDQj+hW5XJFt4OTyyqgc3gyTedi7CUtumg2cPka+2PyR3STxGx4I8+w6
7tCJeHAAPOF7P2ersUgbqF6Sju41fBgI+uFzj3tcf6y3P3LGy9i34XFHQ1xAVgqj
b118jXsiQ6Fib9PWUB2qeR/9i7b3uFbBUV/a0/BkdLy2Y8li+kZNGseW7OpEV932
KBPGCA2n66z4UEj2HaJdWFYQgTh4g3ZX5fLSLeLDblL1LB2w6X+HecA3JH3nr/Ei
JZIzFplJszIB/QdOwWeE05TuwkNuInutpB9wJQBfviMJT34faUD12ZV40UOS5RCE
Rbn/X5Emtn0MgkcWg+KR46QHM+55wM8yOwZWuNfs9XM2eZhfwZ2PnWwpTdsb17W8
GWN2mmjSXq7+JJDNwCytymNcA+QcvIXqxpN8qguinQnUTvCEkRVQjI1LOjua6qtn
z8x+1H2MhFDnZFfP3K6HrteULXhYN9xD/IB0L3jVvWLWQe8z1EcQSxXgOsd5pdQE
45moKCNeZ90ZDZ+8RXSjqkTJrL2q1A0o0cegZRBzrxkm3lL9OCmeZaMUocBFOYUA
8Jd5w3+nwB6rDjvaejyqBCK+6tsRj2mcEDpV4yVHs9CdRSW+DS0LqOnO4ceM6aUe
2/CdMDonXWRt1KVjm08qgB695DtEQIuARLKmmMBU4r9C8gd8LdAm8g2vw6eJwbvf
3tu/fY4JJzwD1EN8a/8WZqNkjJ6ycBVvGpoHnuRqfRT0SFUAC7mQyCxvEsfAW2Da
SgTLAgz36Im5n7kgnncCz/xWt507CVkeMqitwaJGLLg1cQOfh2oSinHIX/1qCPjY
UO2JPFnufHU6FPIblT7C4uj6H7vs0cwuLJYc/DqkQ7M9iC9MWa4dg8xUfUwoDUng
jtVAtAFPfDKrgkkq+6yl+ut4IarxrxvyWsYJ9TXDi9SqSPPPQxqbfWimZvzqVuT7
H0djnfL4rS7A2NyMQXklTkQqRV10DKiaGA5wRzyzXSbJEWYiwu1PWWPb/f4t2xFF
qhqF9oV4q7sHva2wzjwapWN2uS9Ayoa6J5ol88tJJPRcPaWtC1PVvAdKHYbh8ahB
yyS10CssUbfuM4XRgz/4wFJUSIF4fujo1MPf2Vw//7Rj7qmRvNymXcIB5e5UgeU/
2x78MetUU1XeHJWuKfOzzMzkq/mkaYBowifYDmEBJiqdzsYyAAfKWMjuwnazHYoM
9oZn1hBZjlXs/YB8t4HM6hNf8qjQXjqP9/zUmr1zP4TOej0dWJNkeiHZVL0Nw/q6
6773GVmaNTccMf0T6+9Bk9QKxbGeoM5ZSEXAnKqIDRWKmHe2sHlhAXfq4hjgC0VO
cFzD4tRNIi4xxOG0Q1/XPdq8roafoS+o8NgOEj46Y/6HbyJcBVDCjJPmM5MRn63r
0wmi5+T5OP53IefSsEYj26+Z/FtlRi6he9m/5564+5i1IAmchLwE1qFfg5o4VODY
FikTqdXjM/CMktvnaj3fPhpM/FWSa7uYVOL0+klx2y7041kiKyyf3kJNcjN2WyXh
LJQN2BZ6hFJN71aUv32L3TvLAzQ0OYm2E1gMqpSfXpVUov/2t7AsfAtLwB1CL4fe
NrAaEjCQKQ5ht3jm2I5B8ACjkh0q4g5aURrRFKR+SGGwoQNGIFBAlxipeSN/uwem
2rkHbluL4Gi1DT4/7mJ0ZxYvg/yKsUtf8kwEgWzy0rR/crQVeNyOgih+TKUbyIy0
V6GnbuEoEAZhL1Jcqymx2OWclwy8ROaElPS4x8AvRqaEB5XIkDz35XKEMlqeGMMb
Tc/BJpV9ArpMSs8xceU95zVske1CDtKJuAIa37FKm0BsGaMO+KHCeFRl3wnAh25U
LiK2ImNdSQ51jGccRfQNoGK7M0WeB0Y2k2NUIgyzXgPxYDI2A98SQnjwbfbLRP7f
EgfJkbal9wkb4Wu5GPd17nMRi9aW3TjO+g8PbU+V117+hKM8fJBiLv9ZEKsBppeh
45YBL5mLeIdFwRovJIW16Ja4F5LN2xOloS1WziEfXU69CCFD78mTuc4uGUhjE7Nj
d82O3nTbeWBaKWkTMVjo9Gjn+GoMeupJP4ZVe+JjuZfhrtma+DEHvJJAbGsep03e
TQxLUrHkUsf/KTd9v21VFlFpObKdcXuyG9dgj/xk4hMiaZQVximlRzbQsFoJAh/I
OyIeU245I9kCr67Xba3z0Adq/QPs0ZGJ7c79csLRDeWFeE2ga1vB1PM5IQFCFwg+
yXBjpQblt/RcLPCwOFkqoEXHQ3VTIlP35KDUOWPW7VzJso9bsfuuACqJRXMP34DI
sma93It5yJY6AB1ptiLyBMSFSyUaerPUCaPE/TmCsTDuI1m9RNhGRoqK8pdkljjL
G6G3AUjfAFSPZhTa6YThosCag0Co9PP118qmFaND1eAKytw925wmmah9F0Wggf2E
VkUdG89lkbAd5wF48As7G3ivTnsvqdV3Aw0mmYHHK8aZxGZUBkguPSpGiTFOXYr0
FGSOL2dxxmCng/T5dG/1q5WDg7MG1eMBbYxP5VMQszCDv5CxDHuV6bw9QohLX62J
BztEaD3AMATTDXqRMz8dHHl3DQlsgsHgHfx2PXbF3LfNYXNnKOUi8O/HYxcH+JGm
73wfeGueUliRn7WuDoOAnJBtQpgGtKwgnmj5foFcCGlvdIj8PmWciSh2miOj0V9e
tzniTI3/yfXllu0qy7kRemalB0v879VHmKDdhKrD2/eXY7M2LtlJ7sWQ2AewyN1M
0Fi+adgiZg1GF8yYqO3d90y8Ru4eDwaoDehTACVKdEbqmQyi8fqX/K+3jtiyTJSG
GSi98EbhY/03aLQJZk6uuAsXc9VnW0IVuTD5PYQ0jqsmpbWYlLBKJ0Y3L/NGVg05
/Uqu2/eTaAVVugveZoOgSBcF8SDT+DLWbubHVnX8uMSUjHeXMC5+qFhJ3koaAZUz
tCdwpXNEDx1YlKxeVEE+/QTOMUxoxK5tDdDV9QxxNSAdX9tXpD+Cr+kedwXSkJwf
Cl9mFBPxDOoHmSVvWGS0y+EtaVuUm84OhFbymuWJ+bQRlAnhWZ+sagjxA51PgWDZ
NHFFBoeoc8lufPpwbebKyyK+diznj2lgC1oGYN3SDooqeDPvdTLV0FpQ71PuCIpj
uB2r2extedicw3d7LnI66Dq3Zw3cuhHdp38GtEaQ3BmKxlUAExiBzhivrdajH4x4
rSHjhQnaPPXmrxfWyamQiGfTtIf1af5zZbriDr3sey6oDDJMYXhcKLKWEGmDjDxu
ZkNQltSoVki9q9XWw0x7pwSuO0bQsIwFJl91kOkB8Qlz8/BAK2i9JH547mF5enO4
kEjjvN1qQZVEfY7lTsNf/Tm4Led5ggD6EtxfEGk9z8FXdFpmDf8mdmQo8kS6trQU
30CdFHwCtFb1HGiYSI5bRhQMY2uZ8HMi76TYraV9sJs2jSKJCA+AlYqBH+6QqpQl
WRVFO+1vNQDQE8EMqs5eaQCfXf5zGo4WnJdiPndMS4cG0MmTrBznQJedoW654sr0
ISwifiYg/oCFyTsaczl5cN3AZnJf3E+SihyB2fl++PfS3p9po3C2WhuWhZtfU+/D
x6/YT7MG8c+/05K6FbjsZ9jo29ueWVUWV9gjLqzyFsu/8PlYgRMrJl/K6Rx1Yrn7
Fv5NF5RaenzucS+4DNEmfZj5aT04PxvD/VorArkgJz9mkTzmlObWyJ1Lk1LkLNnp
GH0I8TjW/+g894OpJnS8IgAJMbguVYt/biNte90aziGSzi3+8eLeWteVOm1/1QbN
O8ktSG0F7D5/3W5BuDCTilXHDrRjPrNvyrZntowrnB9Aa2iEitC59aZazq2kSTcf
eUZMXQ44CZcsF8pFMMHtcJeZvSL5HMMedpvIv8eVob3pwZ7/ifcuXBoZZONShv5H
JAzoemUlMFqUV2r8+NmNGyx+yVIZ8TvMhZ3fQn6DW9+8KmGUjeFGj0XCOJnvi9ke
qSGN7X/kT22tp18ilfROotLmMivWqVtocEhNWygqo8FjTOLyPQjaXeiS0mwtpkhW
ZJJ3TKQXZE9b6G25s2nIIgjfYe7YKjtCEJ+YEOX2yaDuHAVMoJe93Kaqq+5T+7LD
Q0F4LbnUz9Tz9/GknFAZo6IrAcokI3b9EQJGdAgb4KgpXJjGNXw8f3/ElwGhxYaV
mdTL/FvCdxC/h6EWCBltFCktPnkYGeFbnzco8ljioohlzKxG4PvRzT0DCJwgNhFy
ufmcRoI7MWYZIVxSppIMgmwWsx2kcrDNCfrYZUzvk2LqUljZV1rT4We/be61ue4b
2wHTisJdyEB0iNN4jI+pgwC89ihA8+bIj0BQiR/svvu5IStveJ4k0Ehj2Tw+E7WB
8nSjZq7h/9rM+Ekdu+n5HG5yCvz1kUiEBZuC1dyRKv4NFLoEuyZM5Cf2vkrQ9B9x
LtuwB8OT79XwZe/pD2ozNrE5mNg6JHwyK2CdXIUeG4zzm81BGq71szJ/IfGERx3a
nL873BqycSLHv4MkZlxcNn+So6/yOxzztyQGZLi8HENQicAz1xdI0K74RGyZxu8a
J+AGof/5vk0QRej8Hg4/LaWSZs2lTVmIkoGBh5Q0fYrkjsEhg6oxssjW82xXB25X
Zdb6+y1aRm160l4KBh8aOAr5ET67NQtBMYTg7z7F6cpBxkSbk8EpTw5GrC99OYXa
ulF9bUNsyAtHmz4Ksg+yroawvqGRebun7HMyuOWh3vzJ5tVFiTK6wQW2ODMqVqn5
EHB1EbzsYWI1UndbPQxteyXfKOP2/7pBEtwZXcnq7+N7C8qopYKTqj43sQTlq2qe
W8rTwL0RwMTc5Ujh3qTBEXqrsFbn4zBtnFiMaxOUll+IPkMpNE+CKX2PHpVApfaH
pxvPga84dc3UVnPipszEbSd2snpuX1VQEZ7/TYbhh0Qfh8p5S+EnHry4I9frD/U+
0NX8G4i+GFEjfXa2Oy4N2rKR0j4OR7Cn4lwtGeqIiRoDr2/H5gETSgkYUR/UnTay
7pJgT0L26wxQmj2XGu3nmeusfa4BQq4pxF6FOLDKN4RTqem5t1awSgMliJ3GoxDU
T5Wk7jU7g0uGnIzxbimjbtpOCMLO6aZgGp0wv1hpGJxDQ6IKTkqAysWVETianvrG
iM72ckMrRF7xIwd6w98KEZnD6142GpEEZtpxd1Qw/Qj5Z/+LTU913yicycEdHXf3
ZZ2ojR5jXwomiLXVf91Md2aB4+V6TkiWk5j8Rj+iJQl6bQ93MrY/kkczAcV0DYhZ
ix8TvnSSerMyF/l5JRf0LEwQVIXC7woY17tMpKHjcoY8WiyYW+c3/5LT9mfCWMTX
bPXuHljxULst9tmv2ookbyQXhtImUxRCPAwr/9h9bvTx/s87zcMd9HOht34GNTGk
F55UmMuo80KFHTABNX3RG205ZNn/M5znGvpdDc5WQ/E/RwpdhTYnSaKMbyVTSSHl
kXh+CWGs6RQI9jOXRCc7XrTl/rYWN89Xh9He7iZeg3YzCiWH6wwnbQz090KBUPxu
jgMlJJO/HFLoom1e/cKWXwrtDteNcXU6U0cn/asfThJW5FbGBrLDheAgsXOx0MFO
E4wq3lVe3L3m9G2GJ/SAZ1yU44d6eJbaZY/d+Eo7jkAM457UE3hr9KBpn1bElI4v
kZ1E+RCjD4HzfWHMr8dhm4RAYpa9dhLup/NhepWt3lR3aoo0oDftMSu1PrgvYlgh
y1LE7MTfdnGlL3NGevt4zPJkTAj1DaaRCDh6btD/v95wcUCBzL4GMJJ9+1Wkiwfg
ZpZkk1ltkEWVhTWlfSgsGRah7Q+GjDkC9QU8br21SoRdef1aO6TD456iJEIRfRG+
699gVsCy34aNDbtVte45mac1OmWZx6fIu2qprLDKcDG0Xjna9RuuFJg1/QD5f8YN
fJc8Umo54d30ND5/hVSZsVAsRMguZSqCHhUogWp6oGeqYvjmsIenSBP5LbB8aE/4
qj9Lj7EX3MJtrJyMZ78z8mnh4l2vufMQtUt76u/G5vzdcWDBm12tuk1WpGrE9TfX
WsK/pfhWtkOExPpzyj9wGI2Trp7Ln73yo7V1IXlUOuK1vcuEDjkCrGVJTtO7ItWz
wggZ6yn8ZH0erojtN/HKcTxshiMeKhNKwc311NjSGi/ophJLIz5Z/MidWPfRLqd4
rPf7WPN+QZwBp4a9uaoVwG0VfnI4CVwDN9AuF03gVX0uKi2NE2DtTk+I3fltsXf/
4xpXIIqXDPieUOqD7tqI91TFD9oJLfg+Tg2VHg1deEZkjt5QJG8iSyfYrvOgM0aY
BIanxDb320f2fz5WOAOe2yyN1f1oXMb350jH/In+eCwTEz839srlFJDuB8gg+mYx
vi2M9ERYZ4reoTWPAv/QUiTZs8X7mo5F0ctsbWY6TXRiPFZ89z7ogqA/SVbv1HuL
pp1xOekHA8Saj4zWeU75R6uvFQjgNHRTtbY4JzTvYMegedBZ9TIdL01oAWcFHWhB
xDOZW2Sw6MVmqNudyzxCGkAHx3KqcpXGiWRAz2XbFm8S4GGSw9E+TIgdNSnft6to
E+ghaywVPcHhbdBmIi0wDYjfpIJR/5mpbOKUz1WTzu7sRXxwuFoud12RgiSSMICP
pIidVCkfLNctROATI8s9J5ocW5Pza5B6i3A0Epqtl/T/kUjfHX1L6AJs9PdYEG3c
XxnAGUBitP9S2YfcUfogsFiKFUwpPs/zXjkl+ZjndKMPUi7waA4wypBNw/hXgBt1
h3840foXuraU2Ih/IUUfTdySlOxpmMJUngvpAbZ2ryBHy94v0ox1HVdnMc/9Mcim
iDR7QLzdXNB3bBVkvsdNrFlm8uoeg8s4WiNvItB2SzRZtJOcIItcC71X/ipuY0BZ
e6UogSE+1e9lH7S/rUZQm/0/qPTQYzaw8lUY33MkYzyEIt2mQYc1ELoFPkWeJzPR
XtYzT0E7+CYDBcopZBjFOCuKcrb81XxeJc+SdnFFTGsx+OavNupRdmdi3YUK/426
dWBjO35g9s8KA2DCkBYhIrcFAJ5D/yNJ1s7WJOfpe1D6lGlsJKlPDVuUwajlBQEo
R+0HfTsJKGchNheOL7yepd5JArLETjgD6CuDIHmgH3TKcgX55fFdEpFazfuHPb3d
Zqb5NFP734n0ron+BpyuNktBsCf+u3SNltknlQc4liMu+z6n4VjG/zbrM8M4OAOt
WtGlTJNqWwwXN9VfCrcId4GYJTdvCCoyvZykFPJ/F0OKzixKX1NGf33euY62ZXni
e+qgpitk1SWtUPJTZA8TpFqjkzzA3TIZOPOOnw9LzWoRLAgPVZhx6JdwODUxrRE/
bHsJmY1xLsoMl9jMOCzx7jO+1BIIgUJrj26UWEisWoGST6YtnVp7wamHEAsbuOrA
UhE/DoYgO1Xz0oaiU4Jf1hi2dCLpKQIz+uc8UzFaoGLS7MAylLYPvdmxOk4ryvXA
pq2QnX4q8jea17d+Uq+vcJGfTn4QceVaMEBPoyUF4HYZYc/KSnPBvFGZewB8C176
s5WabU+dTdUs+Z77SqzvhJ6MCC46b9+BXbBiAb/U2GExhQsAs1k6PY94JXu4WDpC
+1OZSBaR9j1jPWLxdkxjWs+NG4RSFbDsfIayK2dsoHVLEo868sN0ZJRIXkF2HBQw
L3OuZTe80iI/rlLBhB6RNjPyF1URXQaKU26kDPevXcJuPUzHKgQ/T7v9Tpt8RkjE
WlOqeRGUOeFc08ao9c6adhL+4WvyBSMaXlbLPMFbm+r9Ev1As0lWKMg8oK+AhqTC
KeVyumhO3ecqyILQP9Ub9S5I/uuinvy/52zYYDrtM9YtbLknEwZ4y5uP2Wl6Rm/J
AyZfEWdq8DlnwomP7NS7TPWCcaEVkudGODBmCkusmAdFeXUTYJjT5AvILHad2gIW
iRgHK/URH0v+1r0CfjeC/9J26GuzUm+Z+sOwCYjcgCcQcVqj6/kRk1HP+pHGX9D2
llwp/kPNWFXmElVTGU9YXfeBB6SpNCVNJr+3J02hX3bUNNbX1j+OeQK4Va7UBluU
T79E654bGka8cTtLHa/WUAgpg/ROl0lfUw5oMal/NASR2fZMcsCL+IBjvaFRPxSH
Ydx2HtbrhgN/9WRF3wvbpn0rCnfKPF9E/aLicDDIJ8nArwbMNsevYplPZmVHxhcn
7IYmhnGRfr0ONGFOWGtqDpDWIG32yM7GNA3nSS1UwJ5FZNMdQoXwFYdrJOqjLBAx
Le/n/cmIvXuJvHN6BOCctEe1hrvyCyIb4dBGWDm1WmM8y9lFvZrwWpfBr9oec0QT
PMfydju80zp+zhrIw2SrXGoKTYlxE+aG7Pjc9BhgdcgxV0abAQLdJ/ZuYSoh6T2O
CMW/V2AaY07+MTfCmcyTXbxPUkaa+F9VJl8xTeQvskNEMK7+5axMIeqyKlT4PSdy
EzSedGX/1W1/ywHT7WAFkD+KyVZbNiwWuy3h8BlLeM0ai8YhhQ0OXBNNwBmrZIZk
JdVJeqAa6iyxBYUQ/KOxMQQa1DInpEgvLHWTGVylBlC7Mu2s7HDcPu3cPrV/km25
5yGU/IwgeUvwf3y3fEQ76BrF9tr23mska5oT6PhcD4OCgDkh51Y0LeoXlp0uowim
EikXK2V+5pIuabpgJtPRCtzL4T9TSmVrKsrGvu9oHfeQq0E41UW7HbcpEhGWft5f
RBoZLgVbV9JGcNTZzgOxd6aD9ujaa/1rvBhIQCumTJOH3SxFYw35E/KGEnicYk26
ttoQCQbH/QTaprmVXQ9wGdHfDKdpzyIzNcy+pK0Vb+OTE+kgXmrwUXRMlQ3uunVA
PKZu0S+jjfhtkyRMiZVbGR13BX/nIVtHDUixtBZknr4ScaNX+aMvm2+g1H2txokO
fU2hwOUVFeluGllln1C8yHJDb4UI+TDeISbtIfX3yF3qGg1QRL5vQq+5g/S89u0D
6SK30Slir3F6qiCHUved3faB5e/6SYMSbq4d+RZaXFfe2Ll3cLeX63q98U2XFX8D
G9htXQoHvifUWRoIUSgp2u3IGSnwMDlYEDBykdf2gEv/fV8u7zhBWkKyM4csza+A
MHNx93HybeCVGsiU5nAD9zG7qXj87eegizYoco1fRJ5hwRLhKNWCPt15NeTWZSDh
ghZxU8lhUW8wB/pfImvYG8hJHWIEWJnqFGvf1iSwAqO4aVQzcmYNRHWlN2WQ3Y/V
V3Y6B0s0wlMXCXVzcn+wCwlvgJZHvIXpvxzTf/QDrj1i6Cw4dapWXpXlh1sKNcMn
cvRkyrj9S74KmOhceApUfoHH8rPhf0XBbSPyvfjaAsUSfca1f63a0QCXdgKGiKTc
0E+I0FzjUcUggXlRZO4e6f9Z93CwvHIEFc3bNBEnsV8TQoJ1Rn6n8R/ugkosJznV
IDZSBp4461368fg+C/Ju6jjMuzg4JtgkKcoiEyHfPMuNRA7QbJ5JqaAjsQMmvcx9
x4Mca1OU0KSdPJRw+AbRhdJC7+UHeOVbkhhL8EOlWWk9B6IkGLtpXLxbRqPRRnA7
NABSNlizCzgkZCsAFt7aHFr638G5ALbRYSX9PF6XCuorD1Y/xeQ7wsOX4hTprW8C
YPrJfvg9KA7Jp4+kDt3aXSh9Wu7zb7bYqJdQ4ovFTzUj+RS2dVmr2VP0tNrsf9as
wpGtPFLsUiesSATDIrEFn/xxkHrwnhZCHCm1oo4Qf5LtsaYsHZWBq7UnFTohBAmf
K49sQotel/EOYRoN0q4AiYMx0o/tsxE44+SQrcA0xZVcm35IxFTt5gbxEthIQNIF
fg2KCEjEA/befmxi6T1H7offpa8Mqje4c2PWa8CutxWOpt4a7drPDdTa/BpnAYMS
UTaBOVq7FSbnKp20uYT0Na6xorgbRvMnYJdVNtrN7U7DfKVshQXkw0GYqw2g0vsx
1kY9Sx9+cYjVsKcM4ycMgtXfSxyjd5XyTk/h3FVlUejZyHF2yxM0zyxlzhc9fqyZ
e52esI/eaiHCAFJLvkkBPsXLl/UhhLn81hyvKbyVzuU5tvX4YhDvbt+yvJ7pcOBl
CAUMi44AQ1LAjW50hV8Nz3Hlu5gofm6eFbBcV8s3Xe2bUTG0vfFwwsUEUZ6k+8QC
wu6MgEhbuG0ObkrKHdZo+NF1kxYfQ+KybQ2Nv+rCqlIw7VqlzgYmEH13htEjxYPP
9OZwDH9kP8Qh/USO2lEDhSz5bV43lsQFsUcujAckGZdg4GasFdlHyOwvIemaSb7R
05u7+vE78yhwaHg+wvp9YPBgdYfYIbiUAkXFBa8pEHboSIi3NlMPp3XMwVzSYbP0
/IgUQsWbvhosWavOceRXfzN1y93SSD9tKA5/MX6TUrXcHRvT9ISfaalBjoh0/oLJ
MSU1RdAIMWC4Gc8QXQFa2d6J7p1vG6LPJpbEVaZ9ja2aoBsnrhMPs6vGm7NicIP2
2/yNExXoHNl/cn9l6DGq0vjh5MVhnsRrbWdPmR1XtwJ6ol/A+PsTRaWWAwzLwgeh
lEcg+U00lFPMc/dgFllaiU/MeyA3ouWupnlJP7Tu5AxnvGHWd07ym17pkmM1emV3
b3agXiEtumXWvVwP0m8lXVdnfBh2gI5h9QzDRCNexYZZTB8sbcvt+oG+T8x26JLJ
CwfxMHhmCX3i5NVuVO2AByDnITcHWUDENm1oJf8kqhyWpF90X1+BXA9pqLs0Cyib
S9xfpZ9oaLtPKqzP1b19S+4F8PTdAscpNRAKNWry1TAp1WjM/KvMTDr/Ej0om3AF
VE4L15XEmVgRKazm+SDHsPu3+dsqOF+xNA/4EU4zsmlcvP2C6Bz+C8GVcapDCVbL
V7Vqh91kFhqM0xCaKon/wKxRYvV3RfluPeUYeAOk646uOesjiAYRK7ehNHo//7yr
5F8pfGRtSVd/OXSWA7pMYKqVU/zKigfMn3C/bOyRtrNscIF/nJ5UpvWERIU1NF6l
SXs14PsBPAVnEGhO+39m6O+W0lnyKO2gkPHw1OEhUS5P3rikWQ/jXdF6kuf8reC5
EHsHwOhCKMIxgxbuqx3Dk3QwWEmgYpXgfwrjryogF/zJUfgoKXmna805TsfnWsSt
lRi0lLxYEPYUDRiPLb7SsaNG69e7Nl8m9MuKe2DMfWd78cjxsFLb936CM+TU1pQE
vGYEp37FnURUHsgNv9kfwPTEBZ3ad0H5qsQd+z3rMvhDvWmNgCzlyOZdz/xnINCK
KIIHNvpm3y/7ksgRWPzAx6SJiTSOLLe1IByeUTojtJ7bEr8AgbTbhPBj6Z/ANugT
a1tAklu9M/qS9jL/ZOanSAy9wStJPIWbv4P3Tyz0dkIN9iau3VNezeMBBtq8iJYN
RQZaIR4utR+52h2ZR5l2WTffHI6Cgp52t/ry0WagM2jZEHguoCHsm0YjNwbVyA5X
EUvU8OFpySbw/hq9ljcJimFHtgm2W/cDpWr0kr8da+0zpLEJIOuH0rZUm/NgU7/r
OGmMOiJY9bessK13oB36/gfPbxaJeFuvcrghlR8ZvvOEu0m/+LWz7cL7JGJaCb7h
VkkZBxAifehmjWdCM3OzbpfcJgE4T3HIXEaw9+bY0RHYBO7cRxX0sJZMTwb96W3T
ciqZ+1YumlcOYuTHwZEv55iH25BZlGknnmVhwsw/y5gFFzgE6XFXIZbydL7H+nmI
Yph/PnN1Wr3rOLajAGp1CtWOvVbS/0WEd9rBurJBurWSwSgMLcvwUsWOgogs0MZK
N0t9QHpD7Jjo/s54zAO64I/JA2Dmk6p48MVS0AjnEk4SCbQ/G/r9jg9R6Fp1+psK
I4jTQ/mEBKRwGyT1eEPJ0rS8VCDgO/buekGxqlKQLBgcrzhJDs+PXam9s5RDAEU0
akcYwCAWyaLEvqHzWeBtcz3UjAQ+9ZklvZLfKSWElrcQ17clrFZZUP4eYYaUa21T
L7oNGUAVia0rOALfhN9MJfRmgz2mWhJcbM69emoYSkaGnK747goCGNbSvutyaVqr
u7DQK/x3rXLQK5GnMroi8bQEuQSAR0Y3KouFdCDDfyPvVTCpHDxZvgtq883PKZwI
gCVBERh+jHv9P8Z71VDUd/v0Fv1g4pIz+xPE8SCITDrSLgkMnjd/xY07UiQUEa9i
6ZfCClKbxVF1iVOPvYL4vUp5eUOgdtuz2Ywvo8S+goJz40nLExl/F2voYwmFchLu
E+qNTdX/2aEdYoETxK1s4KE3/pBRQcDD64w43QetUkogFegTSKeOQNWdI2V3KAwz
6HTgqv7Wr8bPRvaoYBys8r24qCXs+Y5Cl9pJOYKGY+AuMsF7q+UxrMimRNT7FCE2
woxGIhgwWbTD55he1z1AJpDIGLpZ/a4WlB9Mz23bFw6U3D7KpKNVoL7cr2VIJZJi
Bqp2ULnIVTi+zK3dnir5yeVpz1P7KaYYGGuHbJ2SrERyHOVLN3sdh27XkjkVajc8
ontUgIHqFPO2YSeJFbUnFTt9HCaRD/K3Z+QVUBAeA2HBaq/gi0TJC8S+Uq/60Org
Hw95oClnZRI6xk3Kwp7TT9WylgR3aB53n73nsyrWtekfDg723oiSQNrwkvz88/6T
be38NnuiytpuhkPELr9OuPNZVGDoZCFb66SwgUs+q6X10EXk+N0u/l2lZ4Y4bsIP
OzotZP2gZecGJU7tYTRR80sQa1xzesA9F1dNllC/hha3crjnvA/EE/eaKgMqj2he
e4n8ujLDiXBEmSFI1yBK111BTnjdpZeBgW5c4xFv1ZYiDuNcTLaY4rw64aemyCYd
r4fqOYWWL6GPApQynUm8bKExvI3BVGpK8ruYMoTn9Owy8DVG6U35meMzG2QCpMyI
uhHIxepUfQPWyA0eWM4PJ4K3bqm3GIZ02GNT24ZzH64xEHotbiT8hQi8o3gXAqMr
Jy4Fs0g5JHpA+BEkFvcDLIBCz3pTqO0reEIZrx8/ehUGRGhWcSLtCD2y24ndql0y
pzJDwSta5cpDe7EcKljbashoHwBlttkaYMA/lWIkmxqozn61oNowqPjmZUjFV43m
uxoHOgQJrsosa1NYcGB1eR6LuALyb/ERVg591rVgkZq5nBjxSA7APrz47onPnj4G
sDDjQiyE3s1GQ6v+OOV2Bfak03AbLJvl952VsmbnPA/yiDGD4LKieU/bmPB9TTeo
BGnihrNvfjX2uSIbC8ivWCOlOkXOO1+wLC7ZaUz25EbR1H2fi+cuesQjQmBpCGUE
k+cyqwlgDcF9hD9o5EHIdR6uE1mj+XhHozV2WzhnLsUNUa9xoNThJphtSqTgt9Lo
+ToKQ3p+B/MJlnPq2vNImoC8vTZEgc4nhaLWUEKQHrFgUcpfEjlSIMrjJPSHd1XD
+XziEZ5OIDTqe8PB+e5wPi+y+Ohyqd5t9Lv+46aGDL1CAJvM62gedYmTe8jPxjSM
dzpPYaqUEE2z+Mm16V96+/PsdAgNwn5XwiVSekgwrOC7h6VpqUUgMIc0wXoxR/+7
x1m0e0EYmtfmv0qP93IUG4elUc/84EIiF2Que2DDiytRxUfUCpGY/bkpr7MCHn/S
u8CJUAtAp+UH6+k+oqRp5kLeJWDX3ab76zp71LDbY5Z/qhZ4Dlf09Fnxi/FwAYQN
XTuHQ3cdGAkdayipinZ4bXIBaDsP+4cEmKeH5ppSctWAUV1ODcZLgguEWGPzcKGk
1zuZdS5lGKhu5SIP2vk+xkotLo9c4FC7CT+IeUalzBuJRZwaumnXXbXel//o/x/4
DGt9QbzPZN8IO1mUh8TNQ+in3qR0wuOm2PZ0g071R/AzSOM72s2dJbJHbDsnlyr5
ZQXUpPmGJ6Wp7am8JNh2lgobvnkik3ru36AV4CdWHP+HzSZIFhu5yNnlAJg+tPC4
ek0l+NBMtsutXVbdcfKsaBRsj0RtdhDF2U0cTOmZRSWLacYaSu2bJ7DiP2lT677p
jwlHqDGwByMe51S7QP2T3gjYko0fStMC8dGEf5YqRjKi3ao8b5hZgDgp3ji2ycFm
K8KHLb0qeV5w00bRk772/x8/wDOFWVxz6LebGsl/9ZqkJ05Ez3kTlvH6DzYDWvKJ
y565ZYYNVP1uhhHMuac/keBhqMyD72LfTHcOOJNx1/tK54CMjPYUOoGQPZSLhxIQ
/Z1ockd3FAclMIUMxnNvLtmePQWIUecfYlqx7pKVqpJVQ++EWBVd70qOabidN7Q7
Xhfbm+rvnp3L71XbpHq9UbvMJcBqARiKq/I9EM/KV/9rHzvfgRVeud3zeAh1PvfZ
lqtr4wAxP/PcLGgbbDQineVYI1vT+/CdOvOEWuRV3UbXDretXHrECKHWFXMOrttn
u7nr+jkt9TDm7gLWgElsaYugbVM8wXPGlC6eguuV9gbuyZaesvW4X0BTKe739luQ
824E284zrQvK75rCfzM3A3tYvKkqRUHNlInMYiQ5eH1IylcYYPw5UoPfcTR7pR3D
tGXf8/GpqaPG1cQlKKoHdhCJGHMTpvPXVN1Qp8UjjD3ws+UdsL6uUL1h0dEmWnJS
yC98NFXCPv6TvBThVClzJk3wyPVDREQNvWSQY0un+UpE4XSJNFd7CzkLvzTUOD3k
Zs7favNmW0sUCNoMpiebAVvNrqQmDmJyoRmnYr4uDxjScU+bt75hi1su2gO/oaM9
cKDX/VFPYAzQ1yy5OJxH0EO2MlWquH87GTWjThncY5WDfvtXYmKsMZDHD4FoeM13
QfEUcIxl6q7zrSSHCxngBenWwGZRg2RZ2cY/YcV3RtnWGuGerCzT3f56IyGp5siI
37/2Wg0+LUOIO7U344vryt2q/557P8qCocLhQATkAEb8PWEL2oAgqMPKXRYW53kQ
5jwpRBC8a/3aB4Nv6i1f7qzPB+R4geEMEoRqAgHSLhQPL/CMjiKSKjozjzLGVMRP
V/u7gEtsPtiQq39PxJ9SUV8kDdO1S3dsnPE0I4BJ0OGUGrZYI6i4UINcOTMiuyTM
EGeHnW6aB7JHaaWuJ5P7r697HslEAKDyb/BCqui227VucuJngKy8A9dYrEQ3dJMI
SSn5Ga9arpEbJQsWFmLZiOfX9TbxBL3uO5hYZ+fcTN5N8Og7ND/RiksWtpCNq8p2
vvSzUsMCBHZzcG4wsh5yru+/aBR33uZFSuM4/DRT1qfq6RLa3lJ+kCx3B8D96nUZ
iJp30wRs6WH07Of6tYnnC+Sk+o6GjtSCqq8hrHKuu4yZ4t0aaZDbk/K6787myvva
wiRw/RIMQvF7TG3kYEMZN9X2KPmURz4DlL4GKY4lqIwZEGWDAOZwCy7giJViIoB9
v0Ah/xlvO53zYwYfAlrY0AJF/vl+OGwj11iFAE7WY/I/b1gFTrkx8VvuV+d56atV
3DquSJBrpoGrMlUwTS4CS3nHPZRQdHERmRCj+tuTnh75eXBl837wcfQcV4uPIkMw
X7UoOT/fhc6G1Yu2mKRqmBtZ1QuUDhYeKyiwRHX3EG5zkm2WH0/O6CLTrt4ea7ge
xti7WGdB6jgCiY9d/mRdKpjZO4Oqju0PVxsr4rbv3muBHJ2KGejyljNa+ME+UgvI
j1aFmBo94IjPB2kgoS0jD035EFG7D1PNq9W9o2nncwwt9i3GSZwdXp+72YBHERUp
EFzJfh5wWDzygE6FRsd22GhIAfKP/3/twULTEZHEcIh5D6y9dRrYPXlkgIiVIIXI
jrlhAHkrE8BHomQCWUblSJAzSdQ80Qo4CbxVTyjz5SE7FherF1squH9xcFYmpItL
W24Jp+oz6JkG2sUt3uzuaGiSWCxRNXUEOr5zv+ThJS9H5kB+qVr29ZUg0m49muJq
+L61wK5hSKrECVv3Ea8v+SUxr4Rohqmtc9/0CTq2tayG1ktIZR5RHtGFUsEjhMGA
oIjsuknDWx9MBZ74U2m7XjWDYeciHKu7DI4LsMIlupNqAL6AP9R81EJnRLCNSW4b
aoFfar83FJeE4ByCN7wW/efJcVEhPuhfVt8jIF0OgjZi3VZsQGQR8ovEEO6HLwA7
NPNaEgoqOlJSXwLtGATREei7jSVhSKlXCl4ZSxeVy9j6LEXzaGCs1YUSOn1hXXpp
Ii2oQlGtGgiKV5fKKqgBxIUw7IUAZI3ggPK3cpZQ+ympCAAlUfdSJgu7NIeL7pVn
hZI/Un9rUa75rRj4k0+kCFSNpBNJ3ADdJ8C3Y+wYy61bIugWAp4XrRFc/idhggfL
QFDQLBqIAFVnjBHlfQVw3ol+OW7tJWFQxspK0i0Ru69adW9HuLKEm8WHdza7Bsz7
J9VHqaLLH9Or3AA1GkwQimrg8GHYGbUYBGXfxavAXnCXrcYhcM1J+947qtEKtD+a
JFK5lHIy7iYyy4vjPNnPozpYthd2XlWFQcGf5GPtxTzEGCQeiy+YYdiw8epZogeX
w26JeRolgyZdptIuA7fTGi1F0KNKuJnOsj3n68PrtcmpOdwjq5z6b48ZakmhuSNg
4bb1A95bpnPbBndwILW4+p6jjDoj3YI7x+myabPwCNrYBhT+rMUjFUopsH0SLknR
E+QUc8i2ignCpXYpKq5rnNYm/QGuo4HqM+uOpDOvdCteb175qxcGbz/+FPUrsvmy
D58kGLblljcKBkIqAvDu96+9OVEA9NDdPNPmmt1p060hH38osTgdvaBiXJfys+Tj
KYkSQ7MW97rXwZsV8yGFkkkExpFGC0SnicCaKmyV+TjrqYaB+7m8/9e8sOL1Frf+
AjjZIybDNGUooPOFtFgpdXovsTd3La9IQjxMwa8HaIlp0EV/nLnbyxXHS1DulOIj
iPhtqqtiXjMJl/uADtOhnsPboJDYcQCupkTYJWeUpvlxOX/9gBmvaO39hBlWfp11
GoKdPRLYJewheV0k3LPtTtcxG59I8frs6Zc4054uqziVwLD7FJgj41kAf95on9ZR
TV8TA+Au9XffvEyrDyFpL3ouAtbHT5pmjeG93Ch8+RkRnrs5yo9+/VqWHBs2b8HW
ZzqGCtxC24GP4aWm00dJ4+d1c4PGTVjb4YhQ60Z3+gmrX0aT9A42VHBBB3VcdGDF
Xk7aoPATj6IY2CAq3YUIYQBhz/b7Z0jIxDBvSoTgpv5fPtPzhwL2qnh01mPA4m4O
I7lqiWVRPbwuBFoSr6yFdY7cQejNXO/CtS3G9iJpA3FJ5ih4FTviBkrnf3K933IN
nLVvmbHnrnO3OcGNxfTIhn+djAfWjkXpRHo0FE5qTLfciv/W/QnnywXSOmFJGwcS
PvFTcJO27F7ydYhUTZcU5/Jyk+1H+i6O1MLFul7lEVVN3BvnUWNJqL6OQXroVG0D
UJHzrxRPk/UNTMH2ZQZyunqC+wdMGjHnfaPtM8Map624K0t5pjRYAPZh1zJ04EYZ
itMa2Gz6Wx72KwZQewpCqoZdLV+kFW3Q2S/qlnJJA6Lu84oz7WmoNf9Rkn30CA1x
bnipCbBfxHesfFEgOaHiY2uMmcdhKmiJXYHBkIbHzDjbZifJmrjWNgM6XtaP+Cof
MBqsJUhq83hS1wWGYKf7ytJQth2sTNgNjimxznI0xJR8dTCrGc+KuP1ftsJQpbod
tlXsq6tuOR1z5gvIniGcRsesHlLxtY3I6yo4A/cZg1fqnKv8pHryfu2oksWsNxvw
0eeZpEMWAD+aMoSlR6UxdWHaNCsmW38rAq/Bw12wimvmR53gDqV4TsPrNyk3MuM7
7YkgFnXFZnhP8Lo1kkp6IKQ+wlZoxQkym2mDho8Eo6z/jwIGwb69EocZ93RcSk06
sCuyQCTdbWdGA2wUEZeW3c0rlJztb7RDx8vaCw4+HpelBkPxZESOgznvR08G1Ga4
lqU5U1cgjxbQhXpfwtwi5Q22fpZnYos64GRuBykazGtCum9WVC2HwLTVotMEfnc+
rhDRvQfMHin/KWSB8gfbjaMz+Vel7Npz3U19sM29GTUZ87NGb+Xu3reASGgSDl0O
eoWnDfcN3auYBgN6HEtS5ofrwPrIp4DriOVaFxLwNEj3UkS++YlJhzi5NtRgKqEH
XUlunnDuoGnxJ1aoRsQhwrSd5SMAgoWdxN8DlReRejVCCr4FYgPofJIt8dRuP48L
R20y9OZRFWujF+/tMHxvUOTTGOHVeLkxhyDc+ylJn0/7dYuGXQbXjBvKhWdC44Qq
H5AIuYR03dnQaIde8GmG3sYhk3iSqpURzgNfr8jy/Xrpk6dBHPU1cMPS0xhNUK8L
OEG83SRSw52sjcSozGMotYjtGQEqpp7LNRJQBkZ9SFtX3dDaQvhhKpqPwIxIBCXt
2bmJPY43xSSE+AeKaYpgMgoX5qLgMlWjcIK8m25ZGctXyiJoqReIoj0Yi3/VVhOS
dV0mL/rdWLWmIWj5osmSEiW3cp2BN8HoaepY9btpVB8AWy/w48tQksWHWSVsFGg2
IjxQTj9sdXVAM9pJ2g2ggSvh1AH/Zs0JP62EenL95GE46syC6CwP5XAY7PDNgyT/
Yzy3Odhv+IDC/SR1pot8ReVdHE6VDFW9/vbG3pkj5bhTZcp2YJ3+foEGwo0p+jSz
IEsKKWgfP3nn9EuICXMsogdKytsAMb4JQ+rhjRD610GbeadAp5wzYLogF6nL6MB9
AzDL6I8/UEcd6Nj0QNAWqnqwdE9KrILLQcVMqSvKyf1qXCD80fl27Vy9V0yToebn
aCppqyw7bSxFpLnUcBbEpoa1hLNSuQYnsWkimpEzCSgr+tPOfNNUHPiDpp53msdR
4E5Cg7BQKFKUqVV5JA+cNiJeH3fwsksBULo9cIF4IxqJQS9plY/UB+lYxx2VNk0Q
lmiZv+F9+RA7mzO/nweKOXbhjS7YppkOJV6TcqvYdxktD1jm7QiyIo2zHTRjEE48
FUPuKC8mdJmiTjBbisjEd84zzYWCrHa0MLPJGogFlTqtn9aXbWATtzgSDkmOp/NN
TcYSiZqHQhXgh4QaXygWKiNW9MQwNVbPuxryJcD6OxqROB8Otri22aEKLBN6Lzxg
S1s8YCo8Lrco33jIFthega2PuqNFTkzWOFgK5yQX+f3zqSrL0qvGVqbIAR+ENBOf
29qjp1e8zKoBWlq9y81E3pQNQxF4WXqIVnMwML1u+gZdFiP/VkdBM7PiaIXzcmKE
KMr1nMaqtfEq8Qy3hAPUS0Te4S23lbqR/qNyoliMQ4vl02ciVBp309kX3rpIPyX2
GKWzL5jGF877Kp1r9UGJclAkzdD4wIvFAFIQ7ffI51Y4dB1lRPKM2wsIcDtbJF2S
WCfdDW2Z8E2OT1gGqrzFtSfMSPyBgZDtpvlszK6mZkphcoqJcz5Ldx6QznOE2hGH
IpxfZN23VMXDFm0WIOXy1SbkT69lbMuVqiY9VKORaFtI4ywU/JjQ58TAhpU8FWEx
CET/q8rwGRdf00V19oAEeqpX4OLotc02aSP9IhGUxvVWl2ezI9geF/WvUIl7awZT
Qcc7l1cInLKW7UIVNEJFWxXApApQv1oxmlt4ux91CAzFiwHsTRup3HW9TbDqoH1h
nPK33R28/n7p5MCFVDC1WPftDQYDcRSIMad0Kr6HDkXGq4YLaO5Z6IeJnxj+MBzL
f3lNpVUABU6q5hP+kBvJCjVMm476TPFG+i8IOzeot58Pf9VO8KRWcVjRkPVBkipm
qh64osa43Na1MUCo9ExRZcqnx5i+rw95EerqNr7719S9gStYGsLqf5w/GQveG1o6
71AWG2sisGsLmf+0lPlyjv80Lvyb3oesK14TL9V9tdV1dEDcsa0JvFlLggi+jfxv
GLWLcVcTKWi695TMPSS6IuXcaz8jdrrbbxhMlHk5kHYpCDSNQZwnU7bHKX1BEkIO
5HegMzIPCA4MBz/SyiqQA155yN/Bycq6pLc1P0Qcy8DJk5i+J7zMFRt8traYrOFg
n2nJ2uu83FwG2e9mvYS6baLqMdY+QKJdn6AuFFZ7WF/OGALrLrSDPJZHY+scWDt9
3MYUlWta+HOtXFGBW+7vxWvyp08NS8qkKsemME6G9jnqBX8x9opMD//o1GGnSMQc
g6s1JT3hybWQ5SkUk8LX3S7/LFQWCb6pu2gIChmJBpuv0RFDTc2YMSkOl/OWG/Hx
TaR01LERQZQh7jLoVFK+YTOf/XVWyaIKM23vhJSNMxpw9buUa31HCRlkmJvKdVs+
bmFofe1fXiPrG4GXdTePU4U8OY+DvWQUHZTRKbHD32lygv2XaE95QQhvQq9hck+g
Zf6xXSCLB628MaUSxDm6+PwRg05fBHUqmp0Pf0qtbtXskaSd5zsTQFJckZkstG2L
n116/dWs7eQgJwU/2Vq5/846xIJE4h80pgVsmLiJR/0Rk6MPZrTPC2cYGZI8jFb3
lo+CaDD5AkBC5r3fuE7ECcSKtfAsJ4U56aY6eAp6gM/VhPXSac1/J8uI/ql4dZEL
AfO+dtiYzJAAl1rBc2xmoBYI162W1mKKfhwjijFmhho6eprClJXp7KbyECnMNIwx
3rDR37COpQ5t3B76HoT7JnXYiMFzqWHKkCzMAkkVwHZTXBwU8QioXjHxh0XPhmPA
GgulQqHNhFj2FPhrFFyC+T8kCfLqV0/n8m7naiwyO6or9w1GDSagaT52B9Fs+xnO
cTNJaYUN6cLIbsomFhWqQvDcMcZtVuP5gurwSJ2ncxVnBsbUa9r2xDyOPljE0Ui7
8LkGp9WdKHrjDQbBBr9oXK93o5iGOSH6s3h4gk6l5JQwfiVeAWQR4PKEkgf0cN98
3+3JtuyjxUrqsRkHG5sAdqDgRelB1sdqK6VWr12g3MKZuVEOLUKDWcebVAa4mRjL
XUNgahlGxjLUql7F3xyutGFFz5MXtIxVQTNAhpfrnJ6glaLQQe96s/W88srykl/s
+MGzoPHB24BTDP//nUDFamPjK52RUlw/MA2fWH7f2s1Ryf4VdCdPG6BS+8Gc39Up
ijQ7KGyerYK121fgAMRKovp7R5kETnMq3cPeiogeTqfvY2Nll7zLvBK2+x7AH+vb
uhD5dBtLYpmq5rWRhXQcYVlcNv05yPYo5qUaeHADCCzV14fYcAPCR/mZ2On/UXzL
SWgVuJ80+duK7RpYHYrMk6sNkkt2lRejjrgtgpHEKEmrTLpvWU0dchIYvc/7tfCM
vDrBMN25qGhlAW/sr2iXmQiQnyYB5YLmd0qbgNMA5K0QzHYlRJwbDEBRisuMSx1c
yFI+Tz0yJ9uys6DSP8nHMy81EFsDUXO2qXBRS4pp6wSujKm9mkHNC9+d/Eo4X1Kt
TZgmP30rzOWPpGgaolbpBmcGX0v2SRsCxtoR+TeapATSsbNZRK//0RVX4uoozny9
NSDP0rZH4FTvNrAE2aOnAlJPd5oobYhahQG8nWB5Ski0Cpp8sz627QlbIl5g891m
Lafi3ewOX5tP+yFU9nxc0JDCfnm71ecQ4MulwTBPALsd0jqdCmI6ye0S4bLPdogD
soLQSkPTXvDT57yVUwsBgxSebv0lD5q8aSWNAe1s7M0OsxZwK5dF3B53G/hfHku0
roBKmwPEvfsQapJ7Go+XmXM1b0l7NUnKa0UhscrHrCpF3FJnZ3qHaIRWSsYwM5lb
3SrQHdTzeOz7qWza8LdBV+DIS/ZhJcGiQxEccG1Z1AoiWHIsP6miJ8rQhSckCOTE
MwnqBlrd7Und9Oht7yPItutzbuCTPl+FSRkhgOT6HwfruHkHaaDBm3B6ApkjPt4D
xkjW9G3oKlDLbrw69IQML9CtMItHVxtqSvOVAOUtNk/URY00PD0MtALHEgWIQ/gk
ZgmdGr+QdG5DT/gtat2MH3l+rlY96Jqu1OIKuQ1zOcZkmvuiuEC5V6fvkw8eOoIU
aNLQ/v8O2n0dcXgld6qxn/6cL+Hc02R3jGyJgHjdxafInhVScth0VtNVl5hQjZCH
4qxta6fd8qDO4yYqlGs/xKZn/qcjIJC5aV0SjG9PkAKXtmOSlU3oVuYuoGOAo10V
o2EuDd+1V3UjhAaInAhdQfORFSBc+wVG5cJ1OBWzFcBp8zQ3h049+LKUyVA3qmWo
sYxRIAPrl00hj4/C3wclFTCkRyi3gF0RygOtMDjKSF1U0MWmFY9iBHUNnTqXQ5x8
9vm91rtfnPWpsNaSYaL650B3F0hcT+nb+Jx2imWV3EatGSRfh+ttBAejPYDiVXJy
RhyUGi/1ExNMFYWBmcKEHfuGfDGjwKGY5CfLXK3pfqH1J0LAZlT46hyu4TdL3uIC
tUzSbhodO9CAUUpEIPr1ExlJIumRH1KOAZ4LNeXYHBh9rvELl6YojCQmqgS2Kwxs
7U4J1ZT9FWCCvWQ8cgtmnPxTtiABEkGnirDVOU7gbEseGWafg6AJyqF01djVA52e
892GH79EwntvTxiipmYsBPcyDl7yP5ewr0iflYNwWfOnOmLuFZl7MCK7OoRYagIz
8ZSfY1Z/2wLRBkwRjf7ZCSdZ2PXH8Mhi/aOTawRjnmBAaExUHpJ+ij+PjdR8DBcO
cSjnXiBN7hIbp72JCFpm7Ydl2Q1a1T/nuu0zxjCWwFx/Lxv/1T1HXNQBwxKsOuI2
9u5yD7bK2qjOC87jkHAu3lWlFlM+9TdtAuJeUKiXC482lONG/ogDdehqmn5CIUiU
cvLk24AC88cc3bOtNRPG9hK4jg5GXhV7jnSOL5Uj+d0dGDkwAmXJD3Mdehgmh+6H
60gaH5KiYe8Q0NQHV6aEKb8/zeAx25I1US3c1JJYP2vE7q0JWrBvcel10VLfc3Tp
pcMJeS+U2QlkJnk9KeFZXLPWQcV0vYuZmBghCJGwPlf6knjG1Bqd1qHeG7mcTC+B
YjZPjJs5vA11ol9b8aS/BAR+LaiAeXLiYfUXVsUrV043c1jKEEr8YO4E6AGK0k/h
LWVsF5DeJp+tRE6BdgF6qo9cbUgWE4TqooBCWj4qzyHOEEI3X/6pOKaIzYQu4bIY
QM0V71A2hcEpusR5iY5sHLHwyc1SZDvfNROrCmdKkVHnnUd4mvkRR7R0z4c0D6iX
QnccDFRbSGD0g9oGngbSBAeRBi72ew4wHi4pjsq9JTq2CBHsekHYopsjRynKaro3
KC91jNDV5T2z9uRQ/3m1KTh07MVUOx7M+v286E7NSI/gI1nQrV0LNznSn/A+s/Kc
2ehdQw0KBbCKxRJ0VbaaZPYFRjpLtiPJ63X1l+JApQVRriTvtAX0vAKSvVqtk8gw
5aNMyjf4oaw57QC+1An9Gw7QunmSX6UXfKj/Pu+tsTgyJ29LYiKicaqEiLFnBvWL
Y88JJ3yneF06KBZRnSZFG8GiM/cmsqR5E94CNZxtBuXbJDyrRXqETPkFdPLpivSk
DqfJ+w4vFas2cLHQiJQOAy8aXaDPb9ZmY2AaZ5gcHJPnVAXh52LCmIX19TDC+kFF
FYqxe2sEsv4XaZKuAxaPFMV60hia60VM1NUKN/ivNbz4Riey6gMEr89gdR3IqerI
uvMwh4RLifVdTGGKBGBz2gD8HTGLf9vl4iy0gWJ3yxfsMPfS5nWOmOdRX748tGKZ
6N5/qSoddDheVXqwP+oA/H6czQq/wp3prO3d/uMHt6MG6RKRb2O2xqSuRQwqyuUj
DQ6Whdc1PEY3YzmVy2rF4Y3rjYR82wC3+0qcEqaVzHzgBlJizYZQUvGUFrU4iZHz
Wci3gmIs8ce5lp3yVK8sMXHzvQl9nBH57IYVnbxLFTKpyjdqGL4R4cysDIu2UIFB
oJ9yn0P4b9tdoZ/9gADSmnAhjhNzdjyKEUlyZfW5ZgeeYnKQA1Tj/LByVFHL5KMA
2w7pnQF2g4go9Dw2k/PgfgRJ8g18PJJz6BK0eNFW3l1CsGDug60Nm4V+KS+ToF4m
iKCrxTYxHthLnwL93tpVkzXGwb18jjHwI9BKCcxMX/awPw79LBhvrnqE5PPMibwi
kLwn7atuyg+cbYhKXUJXrCsCBjRPdDcH+e53HzSRhlZJhNIYM2w2QFBlKX6c183P
WT2oIoZNhlBD6I9hVfhnWdMgxpLn+Q2qlx3Qqsx9xTanYQ2E+LNLamBixRdrdGqh
n55boeWAs3d/K77FMs0+Ts5PXkw0mX+2fcUp9xpXHngKmgOuQ2caHoqxFdaLcvMv
87cHUVW4B5lECbzJ2RjMlaAgQFN81enNXkfmgEyxFvzV83FutqKzdrMuXOJmmACg
3YovP/JYeRBT5xdvLenNAPpC3uPPwn2Xt7Mv+ywbk0Hm6QLvpoDcR9mB1srjBqtv
fg0XQeNUK6iE6briebz2GNZZ0x1NKqu8DAr194ZIXAU+gUSy5RWq4p/mft4vJEYs
gS5Kh+nQBha1mcYZ45R9gNxvQJqUc5l593P3FcLvRae6Hp28fwPSP3GucPqbk8JO
ir/mVsO0+uJM+SqHzVTPrjrMcqbY8KBM/7T2UPwXren/fx9XS2BX/sM8p9oPYmoB
Ct3VM0ywViA79rJk9Uafg4gjNGwHMBU9NVDHq2SuaKFV6YqvmrJtS6FJJOpKQUax
qIacYRNJQNGaLOark0rxqxkg+0aMrQ3KQUYZo3uIU745ANWIQ0IR6eFaJnRvT32Y
/zB7yFoD04PxJfEBNGyd83v31T6BGZSloCfPdFJa5LDiK5bGiWNK268iz2aDZUpK
kJVPdCbAvzBcXlIzvBQ/PGKtqGFCntk2XnMZrvdtjU3d5cFL+xCTADtXW3Z7E0ll
Om9moLalymKXO5nyd6YPJ8Dbnz9epYDE9jDhg8Y32zlH8X/bwCPGTi0ukyPtN1lX
GSnEae74nUyOF0Bx5Io5VCpMErGEfu2r79GG6xmWQKzPFN1MrUdF0KRjCdmudBN0
cpdAM9wlUSHHMMhapVqVxPtmUvVnaT/JwzoANvmm5OZXhKTVufiGFtX88kJkyJtP
1l7i3tfNGwxaNE15qLPmY4cjuJVB7du1DzlJDzU9hhPH+4n+qgaoYr3GZlUl8MUF
kHWa51ko8+CxzQmq9JYMlYi3IDhYSqRCJq4afRmW7j54r0zXd6Ss8arP1PYxNCsh
99kwAEgRAxnzFTXdiwMnoVOflk2e42kqbVXvfHjHcWjzAWDwKV3UUJLN0XQWEVJr
Vkui1xz18eKN19WtLRCZWBniyPdXeRD4nbXL0uWf56y0XoEhZwl2kTH6njH8hw86
9qjMVu14oDIfImxawJ5DmT5TVgcO1nzlt4YTgpHlEv6kxkYoUf1QBqOf9X3yG/02
/TwpLVb7IJfZB4XUY3RMUQhy8UBAvxpzotm/ld16tuPxhhBeVSGPDLXWBde8gbVN
pESwh4Sw8U8VXZ/nMYDSdl05kQpF/CFF0MhP6HBd0u33me5yazYsGIlGOWFnsgYE
B9QxnXTEki35b1yB35eGygL5NqJh/3S5sL5KMpz5THZYJLU2ENL58CNURDgdArBs
5lqVz7/Ukvaw+76JqEI1L+EoqK5HHN3MhKDN+Mc4qxJHWRLtOl+ba06q7FfPm6T/
b4BhWEiP0fgj6SdZqPpwaXSw2T8RQ2fJQ/33b3ICVyqLDcwsmOEp2lQ7YSIhTFR1
AH9tcIQG9KNGdSlMw5qTfRd7q5hGBrXOERc15znVSw6qsOhw9mOEqX7n4z7u7TAO
gdro3BDNlUc6JnYfgC0U7JyDZOr0dEmIPlEYDYem8Qysu4S3gH3NYq0poHA5JUM6
uvXkYdcNcBvV27kQfTwj0OB833kLy69Hgxly15Frgzfp8gjRwmdVmP7ZViHU3OgW
GeC4hKOZRo2cbLf+lkT5lgXuwRvtsfVxwTJQIJMyFGc9zjyO7javTk8zopWMvJA0
utxHL2nu07dEe4xk36DBYKexyYQdUE9mOG9ceNPzCXYmelBbbHiGuDTDgRktDNBi
VXgeHUPoyEdGnsjbYBXwSeaYti3YSC4+riPTJFdbp3LOj8dIHOBBIqpMEdIU17Zt
jYtq6c1pYJ+Ft4fR3+5Sp2cgUOsr+ucK0eNat6il08ayQY6U5NMDLyxn7PcGCUt8
a4R6aTBDQmnkMKBCWZTKP1VYUZU8Okw8sI0946EfbQlSJjRgv8KuNIXjHUw9uLws
gRipRNV6PiiO5D3QZ9/piN+Beq4sq9+rD/FL/bGROKmvZM9yf1sikiSUz8dZetyI
wQrwGBUbR5IrBT9ccJID2/GNR1f5+fOqQ76VInqKUw9zKORkDhiKkSIumvb2qQGB
RiJ8YZB3jC91brnusmbQSPDfO6Gc2KBre+/OgEzM6AuLnXj8DVOP7XIb/z0+r5c2
kFJ3kpNo3mQZUIo6gm5REbEUnCdOK9gk/smIoMJ+ZAms0XoXprpndsPL1RDKG3/i
oxyauDu2j4d4RVJ6xAu4Z/IYPU4UQLxQDeLCueKiZw9udT9vr4yPB8inX+jLAJ23
orJndWR1MZh+U3VwYfHftHO8kqfj3zFidcAYohBipdwJlPx2vg+YrsVCj2urEw8H
WmyhRWLNcJkYWR48a7R0CoL3dJH/A4E714OIjFZ1R7PyePDTyqzB3n3HKcLVZ8PW
o/J5kVwPC2Ff83+XV3C9NHj9CywqvWVZ0M2gNH4ljzmcJKXxjpSTWidjnqARBFkb
Qep4JJ6cTo0KcytqiZDPtg==
`pragma protect end_protected
