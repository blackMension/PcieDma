`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KlIxHa7PhALSMJIP2sOClTWFjJLKtXTzh/P4uvi6S0oRJI0ucV4hyB2BJpa//ISA
VJSdltAD2J8DvrWX60JfnUEuLpJgiG+CcOZtkYLKX0J1DqwKZ5Dn6S+4xGDmdgz/
BGsZ1Pp0h3aEAHmIiviKjIxPl9StgZrPPtDufFhTneA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4096)
/oxONcUilDrIzTHgxBdBX39PFoAnJzfNmUWWLtcZatGWpcBU8WAkN338cDBOWnFe
PQsKoXrW8iUdL8ywlphX7WjxtdpT6cilscUZUP2+/VR/QQNOTdxTazus8G+YryXa
nIq7l1J1PytZGaLFRAEeUi9rMoaAOWlxFiC16RlxGpGO/vHvLz47esDhjI9oHqzw
Fuvx9U1JaHQ6cIi8jhXgthlVyB6IxTwCsYHJigJUoEJktBHlSbLaHIshQzIIJjRt
visggnyzImCP5i/kpyBXTIUZXQeg7NhcoSB4TGqmdWQDoNFF65hYmkqepwXMiUrQ
OHX23LnNX3D+mVu3uF9/lCKBpt/J0JGjuHaM/WKkjxoz+NPsxCRCMGEGbL5mqjad
uy0byefx5o3ULm9BuEup8hRYfjRGpLEn++2tnExcaoRgMjZwdJc4/TOUhWxhX4bs
qpoG6cjum7or0uzWR5b3jMdVBgXf8k/Ct0mFhoidCHn8em2y38aUDd6iwTYyh1/U
raCMA2/BJeqAv/FMpUMh/8MxPrTN0Suhd/8tqu6G9TPAcxU14ul28x2reU89/l49
h5QDW/iuLP90jkVlP4oIqxcFtuC9N4gU0Zglzfb5E8zbnrLQfzgXYeLPVEmZaTGt
c5XCksBjdh+iUNcBYW2dvlNTk5SD7PcVdIOFQRDAjeb2cNsKc1DNxj8dLKXqpin+
cQAOx2r8ZOn2anrpjb+CmWd86s1j2sXTzJWqrHzKLq9efR7zSiq1O+zvVgQRewCL
Zq/ZjnJY157r4HhM9aj/0eXv5RTIFQR2i3em5kBZu2+Y1Mhitl6QsLSJRAj4kBk9
3mw854bfHW6FMKUmUCHgI4m2df2wZas5HLxqhZf5vOcbRTYrg/JqQevtp1Gg5nJZ
gVE8HeXx1WWs9OWup9Y27F3Ahsh2U9hys8y1cErBGV3dEyaMRJeY8ItJ38Dpq1UF
Z08aa0JYY58hjYSiQGX7LfbuSCAsKqhkHt+wsFvRx0RkLD5HqD8y6+qRUXf5yvbz
8G1Ux9MbEaLi5JFrAvAJp5yE1i8GZ8yhGcKrswXk77MZriX4NFn+uYUpCsYSNrcP
sCe6f2KaHr41EBE0PeWiujqquVdJwFhoUmlCd2KlrUOGRtmNM69frlKFzPZ0CHo1
d+o4bxhIxwwO3CgboXeb7wV3du59H+D8Sjvdft7PVCEKtwXUtj2w6bBNKJF53N7G
72728a0WSMjT+ZtHMIWEmP2PShjB3QTCiU344IoUyR9/42KgycaAZUg9UthN4Cqr
p4nAADYyDYN1wo5nBjvCetiYhwoKmbNZMh4U1aJ+HZCdteQWQirNI2qyO4IJrfAS
VT92ZbKwkL3B6ybGkTNcW5tG1qAs2cQHmY4XLYk9kybWZDmTDJcgnSRDQJzRnwdH
r7p47uzfMSdMp/pp4zGNTZxuAT9JXKhO8RLU1MSnVtMbBnWcIQUnLH5j25QPoM7Y
gQWOmRiw4pgZDbN4DMtyhBR2f38yPfZuhtEvFY44Daf/bVif1K8rd1W1hxIc7U3R
GTkjZkrl0bgaDqaIeQsz22s0d8QZpz90mK2iMnc+F+8Uueqy0XQ/VtkVMMz+kn5a
22v8X1mU0VCXfUlZ/ORqprUtMTWo/HBzAbEJ+Y0xN/3XzDY8IDYX7E0QeI3O5y4u
L9JvaBw1RVW5ot7aOg+ayI/1Ds/BcYxHDRxbl4lwSKWVIXb93QY+wW1Jv0qD+WM0
0bkf9JHM1k517xwcS/56F18JRbR1sQBnMNEsCYaE2DrOq+z3i6W0Dww9IMnEpsP1
acW8AOxQlSTSPBEkpCiMXlYQiIoXXK+BuBlCSf0x60m/97HRwXIvZNlJoDuNZKMc
MHNlyDNtMtED4pAJGXqhQgbzVpFRmypB80HBraqGaefuDLXG3ctgZthR1w0gOY2k
ztoZBIJpm+eFHHnpU6XGPs6n9OBTqkoHNQZp4bw9UtzyT1xy+dT06mrU+wuL6r3y
cPtjtjm8QNjgSD0ndwSJX5oH9AlErQym/UYncVrO9DNPsbEkZzA3qP8p53vTpDAx
XlNwaaTy68wIbrXuESumO/y7gM3zBAqZgIA4c9dCIS6ycG4dNqYk/gqREn071Y68
sJYkj23yxH+YvKhZrtngTGSgdYe8QNIqwMJjqhSKLtmkliJGAe1BCPx6eufx8TI9
OKiz+x6bI3FNzwgdj6tQxpQXL5WxmNM0KaHA19AB7I66Iw8Mtf3LeIVhjhTK5FvS
uZw7dWCjWzmZb9RG3HxHQeQ+/og8G2BhOM45InoAO+0nC2ZA1IW1MYj1UdqsNbdt
3OlimfEjm9D4dxVszCYxkz8ffxZZ0QKdaSHKAWXAdbtdgWiRGPqkF6PiaVxHDxJo
uCaK9NF6LHjtQCOuuylWzyinf051bGSqrtIh66louXcZdUn9YdLGk/quFxbU/iio
cCNZuTexrjIsJ8lj2oHWkKcda9i45grsuOYUtmfbHpfa+rF8pXV7VZ95VJIN4paK
shAmNSbZG9Jcc/n0pnaYRHiibDuhHoFz7TdLoHOcrUmFwjir5IxM8xCaHK1Kww62
GnaVWZML0K+5gUVp3EdQVe2dWi4AvxIdi0crepFA79t54+XOshjycnQjSq+hkxMy
c7fjRyKZMCSULD/T4Dhaw0XQTCbkP2fvfZGG0LtCaw6+QCnJAbdzJnXGeIDU5Jdr
4hi7Qp4zZi1Fkb19S881CSPmmw/rlQfxos0htMOmf8entiR0gCmFAVfq9VBWZwg4
qVkJhaH0RCZGwlluaYE7FpMcIirbAZViOixO0BKvL8/m6J+sj5N+9zuLIhOJtWQq
5hmcCnupVMdUMcgjLCwwvYnk43nutq+5YE1DcZ9n2cFAFvPrkhwWhTr7LWcx4sv5
TFrqbadYRpw87aDFYYhTMdJpuTxtQlpUbCxrB91zqUXh1cVWa9d4gfJH9pF9Z7pi
9OZhdtGWf9Om1XkdVRVTr7gBEjrkpxITWo5C9+AD1MFarJ2RydPhsDrYu6YXKADL
bWGwcza58UjNWoX9dZrcWqDH1eOT162htRVdkqPpJAkeJrR5m/lDyS4Rbas7ljCa
7VxiQkPkFHhXDKjxrQaA+KcsECgAi4lIhI2hbC1wOhHr5r7acKJNKlUplPfaMprS
3MFLW7XXFOb5ZBi3zTQIF3H92gX4ZbyAM/0GTJgxImWxRGjRfr+2mWRjTQpoqLds
Z38SOQgLwh6z7QQWF2B5LgPqBw/FNbsTrkLpgCznas7GFuRpzkO1kTF7HU86CZI8
Pf7HICnCH6kZzq3EhAlAQ0BxPJCpLF0sfTZrpnTLM4JQjIgy6ZAQDDNOsZn/OKup
/chWHCxdKNwrNwFkiA6glEUf+XMnge06xV1jD76Ob+NuWcG4Lyz+7HTfg8lWeOkk
dEY9pEiVrRxmiTrIH4ftc0MI054qWInNu69rMKgXIXOWuz0DMa2gfIlFUjCES6PL
/msy9hCyjSUoKoCobvRFIBigIjq3YhuPCXZgjuKL+/wuTNtjvSxBFgF5hYUb501K
Mo2Fabpaeo8je7uTokgBTXMOkS+FcEV6gIGjKfxPjb5aDUAA+YHan5A0kL+eCRTi
LCrEbjEMTMFhKieMOdUZhQ4nPUYX2IEGQZ/1K0eaXO0ufOFbZVFAK6o/s3cSwnfs
66wH35sI4MyfqgdZgR4OjX6u04wlVCYe2JjEDjx5eau/JmeJqs4XYeZIBE3DdEeU
LtAip6iwkXPwpWRRjDlKqfpRDLP4cSUgFGiqAIYeJKuzxr92f+sKZxxWuX78Pr7t
IP+yaYG3iyyKOBTmPKNk88WuTPEEGXCUT52jLBiNQKgXSG/Hij5dFz+Wwhw3eqGz
bBkwygFAvD97rzUXpxgr/lSfHM6zRROglTeZYG+eDLq2Sh/qQL0ZADdm2MkwJZTd
oc52nfXMpOuzF9I0oERkhXjbmLorDwqhOTAe3r1Yn67gxJqaLPMChQp93o1312Af
NHTuk0XiQTVeqOhdRKFOn5K91I/ZDUKZnE72aIsSn8nctyqTpBrfRd/+ng7K2xBZ
4ymMpKW2ZWFmzL83oqke9CKCAwx7yqL/gl687bZMVfEgiqZ+eizAqR/Gq0q2BAg4
vzoQPVyHzC1ORV8a0Gd0FUmvrg+i/+I3mehsWg1hbF6XHMbSai5lFJTuIN/0/dqX
hK91jxo3/06LipkU2+JIpc+Qbxe6gwLDIOdLIZ9k2CtOFYWofNVVHkqSUGyDS5x6
d7CejVrZzlGIrtJ7HXBWlonqTmfuLHAl2YEtuIHRY6Oo0w6KBLfbr3k/hh2co3kL
QhjVYe3OcwtWeq2y3v0QMAU9E4MfMYfcetSoAMvanovjLoXZtPApJwrLhbrPvCkK
cndZp4qR2mdUxVUPjkJ8KxTv/hVis3ux5yZEq6qIdJnZQaItnD6hQKjVrRujGbjn
a+pwsskASKaVCK3Z5kBBIA/3qoqpd60ZRX3cqA8JOGfCwq+NM14m/Hv4Vih2jCF9
K5e2blWorLsCUHYQGQkxR7gO88bt3/Di7LoEXuZLHfNi4Cs4ScTmte43O5MxtulU
mxFuJXvpXT4C1rJFxmduWi2JoLNChzmrWGHpCr/QOqLJU/E5GXiENuGLVtpsm5jG
5abYpxKd0qhW+MjqDHOpdrqnmCxv5hkdgeSCgXEh2XEyK9bfdeLCXsQEFo7yqygQ
CactebxJpJQQWFwlepdF+LWyXGVVvuFEB0VYzo9rfvAaEWxbJu4Sazwpmu5mrgwU
qJtpF4iYuTBZn8fcPRP3ad+l0LhwR5psNB+fSGT4g4JgC8mKXOpXme88IJu2o2sa
XiU1CwS2+AT/fQU10hryD1lNUlgwik+GQueRDg1vQeY7ayISbXDqP8H+X8HIxKri
anurGp/c0oJ5uciJX1IBnhMcfHIM6beCD4F7YB/PRJFHvl5jc/Db2Ahh+6plPaXd
7yAyM6TltUP4tjAQ9hnIH6nkeBuj9TKFxPUmUBIH7l9/qEYRz0FFsI9Dspop60+/
GHxVcp1rFc5QUuhe64ta3RYTR7kki5n6wMSAYtkfqPeMPBAHYWOmtST1vwTS3Ekx
8tPl7plWNQNiUvo7tipAH4ZGkpS+QBw5ycCfCxWrA2JdLsHLe5g7FaTOkPzQ3ATT
pgWvF/VhDm1J9R8fBRCl7VOfdvbOmWGaRnCqP2cVV9duDvkridVuQRB6XTbjZryv
CPIRGCCMh17zUrAbrZGF34iUgxm6lROZoy+ZWhCUQe+Uciigq8mD4e+IX241di3X
CrLfRbcWb7sQG5y3avSLSRHrtLhSBJaAO3bwbNpcJOrjHbw9XhkiKyQIUTOPhJoM
mtrILf3ny3IM2FHk5Ek8kQoyEgpBaZl9mm8nzQCrZiMNcLL+rZN/iCTfnCydVH0s
yYlO9m+MtzYZ9aoSUb01LkBBMbxRgafZi7sGDNBCJHp0BK7ZM62TWu+vWeSvhQtF
kzfYhy7bxH7g67k8FFtGVA==
`pragma protect end_protected
