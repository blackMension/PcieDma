// Phy_tb.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module Phy_tb (
	);

	wire  [31:0] phy_inst_reconfig_avmm_readdata;                                      // Phy_inst:reconfig_readdata -> Phy_inst_reconfig_avmm_bfm:sig_readdata
	wire   [0:0] phy_inst_reconfig_avmm_waitrequest;                                   // Phy_inst:reconfig_waitrequest -> Phy_inst_reconfig_avmm_bfm:sig_waitrequest
	wire   [9:0] phy_inst_reconfig_avmm_bfm_conduit_address;                           // Phy_inst_reconfig_avmm_bfm:sig_address -> Phy_inst:reconfig_address
	wire   [0:0] phy_inst_reconfig_avmm_bfm_conduit_read;                              // Phy_inst_reconfig_avmm_bfm:sig_read -> Phy_inst:reconfig_read
	wire   [0:0] phy_inst_reconfig_avmm_bfm_conduit_write;                             // Phy_inst_reconfig_avmm_bfm:sig_write -> Phy_inst:reconfig_write
	wire  [31:0] phy_inst_reconfig_avmm_bfm_conduit_writedata;                         // Phy_inst_reconfig_avmm_bfm:sig_writedata -> Phy_inst:reconfig_writedata
	wire   [0:0] phy_inst_reconfig_clk_bfm_conduit_clk;                                // Phy_inst_reconfig_clk_bfm:sig_clk -> Phy_inst:reconfig_clk
	wire   [0:0] phy_inst_reconfig_reset_bfm_conduit_reset;                            // Phy_inst_reconfig_reset_bfm:sig_reset -> Phy_inst:reconfig_reset
	wire   [0:0] phy_inst_rx_analogreset_bfm_conduit_rx_analogreset;                   // Phy_inst_rx_analogreset_bfm:sig_rx_analogreset -> Phy_inst:rx_analogreset
	wire   [0:0] phy_inst_rx_cal_busy_rx_cal_busy;                                     // Phy_inst:rx_cal_busy -> Phy_inst_rx_cal_busy_bfm:sig_rx_cal_busy
	wire   [0:0] phy_inst_rx_cdr_refclk0_bfm_conduit_clk;                              // Phy_inst_rx_cdr_refclk0_bfm:sig_clk -> Phy_inst:rx_cdr_refclk0
	wire   [0:0] phy_inst_rx_clkout_clk;                                               // Phy_inst:rx_clkout -> Phy_inst_rx_clkout_bfm:sig_clk
	wire   [7:0] phy_inst_rx_control_rx_control;                                       // Phy_inst:rx_control -> Phy_inst_rx_control_bfm:sig_rx_control
	wire   [0:0] phy_inst_rx_coreclkin_bfm_conduit_clk;                                // Phy_inst_rx_coreclkin_bfm:sig_clk -> Phy_inst:rx_coreclkin
	wire   [0:0] phy_inst_rx_digitalreset_bfm_conduit_rx_digitalreset;                 // Phy_inst_rx_digitalreset_bfm:sig_rx_digitalreset -> Phy_inst:rx_digitalreset
	wire   [0:0] phy_inst_rx_enh_blk_lock_rx_enh_blk_lock;                             // Phy_inst:rx_enh_blk_lock -> Phy_inst_rx_enh_blk_lock_bfm:sig_rx_enh_blk_lock
	wire   [0:0] phy_inst_rx_enh_data_valid_rx_enh_data_valid;                         // Phy_inst:rx_enh_data_valid -> Phy_inst_rx_enh_data_valid_bfm:sig_rx_enh_data_valid
	wire   [0:0] phy_inst_rx_enh_fifo_del_rx_enh_fifo_del;                             // Phy_inst:rx_enh_fifo_del -> Phy_inst_rx_enh_fifo_del_bfm:sig_rx_enh_fifo_del
	wire   [0:0] phy_inst_rx_enh_fifo_empty_rx_enh_fifo_empty;                         // Phy_inst:rx_enh_fifo_empty -> Phy_inst_rx_enh_fifo_empty_bfm:sig_rx_enh_fifo_empty
	wire   [0:0] phy_inst_rx_enh_fifo_full_rx_enh_fifo_full;                           // Phy_inst:rx_enh_fifo_full -> Phy_inst_rx_enh_fifo_full_bfm:sig_rx_enh_fifo_full
	wire   [0:0] phy_inst_rx_enh_fifo_insert_rx_enh_fifo_insert;                       // Phy_inst:rx_enh_fifo_insert -> Phy_inst_rx_enh_fifo_insert_bfm:sig_rx_enh_fifo_insert
	wire   [0:0] phy_inst_rx_enh_highber_rx_enh_highber;                               // Phy_inst:rx_enh_highber -> Phy_inst_rx_enh_highber_bfm:sig_rx_enh_highber
	wire   [0:0] phy_inst_rx_is_lockedtodata_rx_is_lockedtodata;                       // Phy_inst:rx_is_lockedtodata -> Phy_inst_rx_is_lockedtodata_bfm:sig_rx_is_lockedtodata
	wire   [0:0] phy_inst_rx_is_lockedtoref_rx_is_lockedtoref;                         // Phy_inst:rx_is_lockedtoref -> Phy_inst_rx_is_lockedtoref_bfm:sig_rx_is_lockedtoref
	wire  [63:0] phy_inst_rx_parallel_data_rx_parallel_data;                           // Phy_inst:rx_parallel_data -> Phy_inst_rx_parallel_data_bfm:sig_rx_parallel_data
	wire   [0:0] phy_inst_rx_pma_div_clkout_clk;                                       // Phy_inst:rx_pma_div_clkout -> Phy_inst_rx_pma_div_clkout_bfm:sig_clk
	wire   [0:0] phy_inst_rx_serial_data_bfm_conduit_rx_serial_data;                   // Phy_inst_rx_serial_data_bfm:sig_rx_serial_data -> Phy_inst:rx_serial_data
	wire   [0:0] phy_inst_tx_analogreset_bfm_conduit_tx_analogreset;                   // Phy_inst_tx_analogreset_bfm:sig_tx_analogreset -> Phy_inst:tx_analogreset
	wire   [0:0] phy_inst_tx_cal_busy_tx_cal_busy;                                     // Phy_inst:tx_cal_busy -> Phy_inst_tx_cal_busy_bfm:sig_tx_cal_busy
	wire   [0:0] phy_inst_tx_clkout_clk;                                               // Phy_inst:tx_clkout -> Phy_inst_tx_clkout_bfm:sig_clk
	wire   [7:0] phy_inst_tx_control_bfm_conduit_tx_control;                           // Phy_inst_tx_control_bfm:sig_tx_control -> Phy_inst:tx_control
	wire   [0:0] phy_inst_tx_coreclkin_bfm_conduit_clk;                                // Phy_inst_tx_coreclkin_bfm:sig_clk -> Phy_inst:tx_coreclkin
	wire   [0:0] phy_inst_tx_digitalreset_bfm_conduit_tx_digitalreset;                 // Phy_inst_tx_digitalreset_bfm:sig_tx_digitalreset -> Phy_inst:tx_digitalreset
	wire   [0:0] phy_inst_tx_enh_data_valid_bfm_conduit_tx_enh_data_valid;             // Phy_inst_tx_enh_data_valid_bfm:sig_tx_enh_data_valid -> Phy_inst:tx_enh_data_valid
	wire   [0:0] phy_inst_tx_enh_fifo_empty_tx_enh_fifo_empty;                         // Phy_inst:tx_enh_fifo_empty -> Phy_inst_tx_enh_fifo_empty_bfm:sig_tx_enh_fifo_empty
	wire   [0:0] phy_inst_tx_enh_fifo_full_tx_enh_fifo_full;                           // Phy_inst:tx_enh_fifo_full -> Phy_inst_tx_enh_fifo_full_bfm:sig_tx_enh_fifo_full
	wire   [0:0] phy_inst_tx_enh_fifo_pempty_tx_enh_fifo_pempty;                       // Phy_inst:tx_enh_fifo_pempty -> Phy_inst_tx_enh_fifo_pempty_bfm:sig_tx_enh_fifo_pempty
	wire   [0:0] phy_inst_tx_enh_fifo_pfull_tx_enh_fifo_pfull;                         // Phy_inst:tx_enh_fifo_pfull -> Phy_inst_tx_enh_fifo_pfull_bfm:sig_tx_enh_fifo_pfull
	wire   [0:0] phy_inst_tx_err_ins_bfm_conduit_tx_err_ins;                           // Phy_inst_tx_err_ins_bfm:sig_tx_err_ins -> Phy_inst:tx_err_ins
	wire  [63:0] phy_inst_tx_parallel_data_bfm_conduit_tx_parallel_data;               // Phy_inst_tx_parallel_data_bfm:sig_tx_parallel_data -> Phy_inst:tx_parallel_data
	wire   [0:0] phy_inst_tx_pma_div_clkout_clk;                                       // Phy_inst:tx_pma_div_clkout -> Phy_inst_tx_pma_div_clkout_bfm:sig_clk
	wire   [0:0] phy_inst_tx_serial_clk0_bfm_conduit_clk;                              // Phy_inst_tx_serial_clk0_bfm:sig_clk -> Phy_inst:tx_serial_clk0
	wire   [0:0] phy_inst_tx_serial_data_tx_serial_data;                               // Phy_inst:tx_serial_data -> Phy_inst_tx_serial_data_bfm:sig_tx_serial_data
	wire  [11:0] phy_inst_unused_rx_control_unused_rx_control;                         // Phy_inst:unused_rx_control -> Phy_inst_unused_rx_control_bfm:sig_unused_rx_control
	wire  [63:0] phy_inst_unused_rx_parallel_data_unused_rx_parallel_data;             // Phy_inst:unused_rx_parallel_data -> Phy_inst_unused_rx_parallel_data_bfm:sig_unused_rx_parallel_data
	wire   [8:0] phy_inst_unused_tx_control_bfm_conduit_unused_tx_control;             // Phy_inst_unused_tx_control_bfm:sig_unused_tx_control -> Phy_inst:unused_tx_control
	wire  [63:0] phy_inst_unused_tx_parallel_data_bfm_conduit_unused_tx_parallel_data; // Phy_inst_unused_tx_parallel_data_bfm:sig_unused_tx_parallel_data -> Phy_inst:unused_tx_parallel_data

	Phy phy_inst (
		.reconfig_write          (phy_inst_reconfig_avmm_bfm_conduit_write),                             //   input,   width = 1,           reconfig_avmm.write
		.reconfig_read           (phy_inst_reconfig_avmm_bfm_conduit_read),                              //   input,   width = 1,                        .read
		.reconfig_address        (phy_inst_reconfig_avmm_bfm_conduit_address),                           //   input,  width = 10,                        .address
		.reconfig_writedata      (phy_inst_reconfig_avmm_bfm_conduit_writedata),                         //   input,  width = 32,                        .writedata
		.reconfig_readdata       (phy_inst_reconfig_avmm_readdata),                                      //  output,  width = 32,                        .readdata
		.reconfig_waitrequest    (phy_inst_reconfig_avmm_waitrequest),                                   //  output,   width = 1,                        .waitrequest
		.reconfig_clk            (phy_inst_reconfig_clk_bfm_conduit_clk),                                //   input,   width = 1,            reconfig_clk.clk
		.reconfig_reset          (phy_inst_reconfig_reset_bfm_conduit_reset),                            //   input,   width = 1,          reconfig_reset.reset
		.rx_analogreset          (phy_inst_rx_analogreset_bfm_conduit_rx_analogreset),                   //   input,   width = 1,          rx_analogreset.rx_analogreset
		.rx_cal_busy             (phy_inst_rx_cal_busy_rx_cal_busy),                                     //  output,   width = 1,             rx_cal_busy.rx_cal_busy
		.rx_cdr_refclk0          (phy_inst_rx_cdr_refclk0_bfm_conduit_clk),                              //   input,   width = 1,          rx_cdr_refclk0.clk
		.rx_clkout               (phy_inst_rx_clkout_clk),                                               //  output,   width = 1,               rx_clkout.clk
		.rx_control              (phy_inst_rx_control_rx_control),                                       //  output,   width = 8,              rx_control.rx_control
		.rx_coreclkin            (phy_inst_rx_coreclkin_bfm_conduit_clk),                                //   input,   width = 1,            rx_coreclkin.clk
		.rx_digitalreset         (phy_inst_rx_digitalreset_bfm_conduit_rx_digitalreset),                 //   input,   width = 1,         rx_digitalreset.rx_digitalreset
		.rx_enh_blk_lock         (phy_inst_rx_enh_blk_lock_rx_enh_blk_lock),                             //  output,   width = 1,         rx_enh_blk_lock.rx_enh_blk_lock
		.rx_enh_data_valid       (phy_inst_rx_enh_data_valid_rx_enh_data_valid),                         //  output,   width = 1,       rx_enh_data_valid.rx_enh_data_valid
		.rx_enh_fifo_del         (phy_inst_rx_enh_fifo_del_rx_enh_fifo_del),                             //  output,   width = 1,         rx_enh_fifo_del.rx_enh_fifo_del
		.rx_enh_fifo_empty       (phy_inst_rx_enh_fifo_empty_rx_enh_fifo_empty),                         //  output,   width = 1,       rx_enh_fifo_empty.rx_enh_fifo_empty
		.rx_enh_fifo_full        (phy_inst_rx_enh_fifo_full_rx_enh_fifo_full),                           //  output,   width = 1,        rx_enh_fifo_full.rx_enh_fifo_full
		.rx_enh_fifo_insert      (phy_inst_rx_enh_fifo_insert_rx_enh_fifo_insert),                       //  output,   width = 1,      rx_enh_fifo_insert.rx_enh_fifo_insert
		.rx_enh_highber          (phy_inst_rx_enh_highber_rx_enh_highber),                               //  output,   width = 1,          rx_enh_highber.rx_enh_highber
		.rx_is_lockedtodata      (phy_inst_rx_is_lockedtodata_rx_is_lockedtodata),                       //  output,   width = 1,      rx_is_lockedtodata.rx_is_lockedtodata
		.rx_is_lockedtoref       (phy_inst_rx_is_lockedtoref_rx_is_lockedtoref),                         //  output,   width = 1,       rx_is_lockedtoref.rx_is_lockedtoref
		.rx_parallel_data        (phy_inst_rx_parallel_data_rx_parallel_data),                           //  output,  width = 64,        rx_parallel_data.rx_parallel_data
		.rx_pma_div_clkout       (phy_inst_rx_pma_div_clkout_clk),                                       //  output,   width = 1,       rx_pma_div_clkout.clk
		.rx_serial_data          (phy_inst_rx_serial_data_bfm_conduit_rx_serial_data),                   //   input,   width = 1,          rx_serial_data.rx_serial_data
		.tx_analogreset          (phy_inst_tx_analogreset_bfm_conduit_tx_analogreset),                   //   input,   width = 1,          tx_analogreset.tx_analogreset
		.tx_cal_busy             (phy_inst_tx_cal_busy_tx_cal_busy),                                     //  output,   width = 1,             tx_cal_busy.tx_cal_busy
		.tx_clkout               (phy_inst_tx_clkout_clk),                                               //  output,   width = 1,               tx_clkout.clk
		.tx_control              (phy_inst_tx_control_bfm_conduit_tx_control),                           //   input,   width = 8,              tx_control.tx_control
		.tx_coreclkin            (phy_inst_tx_coreclkin_bfm_conduit_clk),                                //   input,   width = 1,            tx_coreclkin.clk
		.tx_digitalreset         (phy_inst_tx_digitalreset_bfm_conduit_tx_digitalreset),                 //   input,   width = 1,         tx_digitalreset.tx_digitalreset
		.tx_enh_data_valid       (phy_inst_tx_enh_data_valid_bfm_conduit_tx_enh_data_valid),             //   input,   width = 1,       tx_enh_data_valid.tx_enh_data_valid
		.tx_enh_fifo_empty       (phy_inst_tx_enh_fifo_empty_tx_enh_fifo_empty),                         //  output,   width = 1,       tx_enh_fifo_empty.tx_enh_fifo_empty
		.tx_enh_fifo_full        (phy_inst_tx_enh_fifo_full_tx_enh_fifo_full),                           //  output,   width = 1,        tx_enh_fifo_full.tx_enh_fifo_full
		.tx_enh_fifo_pempty      (phy_inst_tx_enh_fifo_pempty_tx_enh_fifo_pempty),                       //  output,   width = 1,      tx_enh_fifo_pempty.tx_enh_fifo_pempty
		.tx_enh_fifo_pfull       (phy_inst_tx_enh_fifo_pfull_tx_enh_fifo_pfull),                         //  output,   width = 1,       tx_enh_fifo_pfull.tx_enh_fifo_pfull
		.tx_err_ins              (phy_inst_tx_err_ins_bfm_conduit_tx_err_ins),                           //   input,   width = 1,              tx_err_ins.tx_err_ins
		.tx_parallel_data        (phy_inst_tx_parallel_data_bfm_conduit_tx_parallel_data),               //   input,  width = 64,        tx_parallel_data.tx_parallel_data
		.tx_pma_div_clkout       (phy_inst_tx_pma_div_clkout_clk),                                       //  output,   width = 1,       tx_pma_div_clkout.clk
		.tx_serial_clk0          (phy_inst_tx_serial_clk0_bfm_conduit_clk),                              //   input,   width = 1,          tx_serial_clk0.clk
		.tx_serial_data          (phy_inst_tx_serial_data_tx_serial_data),                               //  output,   width = 1,          tx_serial_data.tx_serial_data
		.unused_rx_control       (phy_inst_unused_rx_control_unused_rx_control),                         //  output,  width = 12,       unused_rx_control.unused_rx_control
		.unused_rx_parallel_data (phy_inst_unused_rx_parallel_data_unused_rx_parallel_data),             //  output,  width = 64, unused_rx_parallel_data.unused_rx_parallel_data
		.unused_tx_control       (phy_inst_unused_tx_control_bfm_conduit_unused_tx_control),             //   input,   width = 9,       unused_tx_control.unused_tx_control
		.unused_tx_parallel_data (phy_inst_unused_tx_parallel_data_bfm_conduit_unused_tx_parallel_data)  //   input,  width = 64, unused_tx_parallel_data.unused_tx_parallel_data
	);

	Phy_inst_reconfig_avmm_bfm_ip phy_inst_reconfig_avmm_bfm (
		.sig_address     (phy_inst_reconfig_avmm_bfm_conduit_address),   //  output,  width = 10, conduit.address
		.sig_read        (phy_inst_reconfig_avmm_bfm_conduit_read),      //  output,   width = 1,        .read
		.sig_readdata    (phy_inst_reconfig_avmm_readdata),              //   input,  width = 32,        .readdata
		.sig_waitrequest (phy_inst_reconfig_avmm_waitrequest),           //   input,   width = 1,        .waitrequest
		.sig_write       (phy_inst_reconfig_avmm_bfm_conduit_write),     //  output,   width = 1,        .write
		.sig_writedata   (phy_inst_reconfig_avmm_bfm_conduit_writedata)  //  output,  width = 32,        .writedata
	);

	Phy_inst_reconfig_clk_bfm_ip phy_inst_reconfig_clk_bfm (
		.sig_clk (phy_inst_reconfig_clk_bfm_conduit_clk)  //  output,  width = 1, conduit.clk
	);

	Phy_inst_reconfig_reset_bfm_ip phy_inst_reconfig_reset_bfm (
		.sig_reset (phy_inst_reconfig_reset_bfm_conduit_reset)  //  output,  width = 1, conduit.reset
	);

	Phy_inst_rx_analogreset_bfm_ip phy_inst_rx_analogreset_bfm (
		.sig_rx_analogreset (phy_inst_rx_analogreset_bfm_conduit_rx_analogreset)  //  output,  width = 1, conduit.rx_analogreset
	);

	Phy_inst_rx_cal_busy_bfm_ip phy_inst_rx_cal_busy_bfm (
		.sig_rx_cal_busy (phy_inst_rx_cal_busy_rx_cal_busy)  //   input,  width = 1, conduit.rx_cal_busy
	);

	Phy_inst_rx_cdr_refclk0_bfm_ip phy_inst_rx_cdr_refclk0_bfm (
		.sig_clk (phy_inst_rx_cdr_refclk0_bfm_conduit_clk)  //  output,  width = 1, conduit.clk
	);

	Phy_inst_rx_clkout_bfm_ip phy_inst_rx_clkout_bfm (
		.sig_clk (phy_inst_rx_clkout_clk)  //   input,  width = 1, conduit.clk
	);

	Phy_inst_rx_control_bfm_ip phy_inst_rx_control_bfm (
		.sig_rx_control (phy_inst_rx_control_rx_control)  //   input,  width = 8, conduit.rx_control
	);

	Phy_inst_rx_coreclkin_bfm_ip phy_inst_rx_coreclkin_bfm (
		.sig_clk (phy_inst_rx_coreclkin_bfm_conduit_clk)  //  output,  width = 1, conduit.clk
	);

	Phy_inst_rx_digitalreset_bfm_ip phy_inst_rx_digitalreset_bfm (
		.sig_rx_digitalreset (phy_inst_rx_digitalreset_bfm_conduit_rx_digitalreset)  //  output,  width = 1, conduit.rx_digitalreset
	);

	Phy_inst_rx_enh_blk_lock_bfm_ip phy_inst_rx_enh_blk_lock_bfm (
		.sig_rx_enh_blk_lock (phy_inst_rx_enh_blk_lock_rx_enh_blk_lock)  //   input,  width = 1, conduit.rx_enh_blk_lock
	);

	Phy_inst_rx_enh_data_valid_bfm_ip phy_inst_rx_enh_data_valid_bfm (
		.sig_rx_enh_data_valid (phy_inst_rx_enh_data_valid_rx_enh_data_valid)  //   input,  width = 1, conduit.rx_enh_data_valid
	);

	Phy_inst_rx_enh_fifo_del_bfm_ip phy_inst_rx_enh_fifo_del_bfm (
		.sig_rx_enh_fifo_del (phy_inst_rx_enh_fifo_del_rx_enh_fifo_del)  //   input,  width = 1, conduit.rx_enh_fifo_del
	);

	Phy_inst_rx_enh_fifo_empty_bfm_ip phy_inst_rx_enh_fifo_empty_bfm (
		.sig_rx_enh_fifo_empty (phy_inst_rx_enh_fifo_empty_rx_enh_fifo_empty)  //   input,  width = 1, conduit.rx_enh_fifo_empty
	);

	Phy_inst_rx_enh_fifo_full_bfm_ip phy_inst_rx_enh_fifo_full_bfm (
		.sig_rx_enh_fifo_full (phy_inst_rx_enh_fifo_full_rx_enh_fifo_full)  //   input,  width = 1, conduit.rx_enh_fifo_full
	);

	Phy_inst_rx_enh_fifo_insert_bfm_ip phy_inst_rx_enh_fifo_insert_bfm (
		.sig_rx_enh_fifo_insert (phy_inst_rx_enh_fifo_insert_rx_enh_fifo_insert)  //   input,  width = 1, conduit.rx_enh_fifo_insert
	);

	Phy_inst_rx_enh_highber_bfm_ip phy_inst_rx_enh_highber_bfm (
		.sig_rx_enh_highber (phy_inst_rx_enh_highber_rx_enh_highber)  //   input,  width = 1, conduit.rx_enh_highber
	);

	Phy_inst_rx_is_lockedtodata_bfm_ip phy_inst_rx_is_lockedtodata_bfm (
		.sig_rx_is_lockedtodata (phy_inst_rx_is_lockedtodata_rx_is_lockedtodata)  //   input,  width = 1, conduit.rx_is_lockedtodata
	);

	Phy_inst_rx_is_lockedtoref_bfm_ip phy_inst_rx_is_lockedtoref_bfm (
		.sig_rx_is_lockedtoref (phy_inst_rx_is_lockedtoref_rx_is_lockedtoref)  //   input,  width = 1, conduit.rx_is_lockedtoref
	);

	Phy_inst_rx_parallel_data_bfm_ip phy_inst_rx_parallel_data_bfm (
		.sig_rx_parallel_data (phy_inst_rx_parallel_data_rx_parallel_data)  //   input,  width = 64, conduit.rx_parallel_data
	);

	Phy_inst_rx_pma_div_clkout_bfm_ip phy_inst_rx_pma_div_clkout_bfm (
		.sig_clk (phy_inst_rx_pma_div_clkout_clk)  //   input,  width = 1, conduit.clk
	);

	Phy_inst_rx_serial_data_bfm_ip phy_inst_rx_serial_data_bfm (
		.sig_rx_serial_data (phy_inst_rx_serial_data_bfm_conduit_rx_serial_data)  //  output,  width = 1, conduit.rx_serial_data
	);

	Phy_inst_tx_analogreset_bfm_ip phy_inst_tx_analogreset_bfm (
		.sig_tx_analogreset (phy_inst_tx_analogreset_bfm_conduit_tx_analogreset)  //  output,  width = 1, conduit.tx_analogreset
	);

	Phy_inst_tx_cal_busy_bfm_ip phy_inst_tx_cal_busy_bfm (
		.sig_tx_cal_busy (phy_inst_tx_cal_busy_tx_cal_busy)  //   input,  width = 1, conduit.tx_cal_busy
	);

	Phy_inst_tx_clkout_bfm_ip phy_inst_tx_clkout_bfm (
		.sig_clk (phy_inst_tx_clkout_clk)  //   input,  width = 1, conduit.clk
	);

	Phy_inst_tx_control_bfm_ip phy_inst_tx_control_bfm (
		.sig_tx_control (phy_inst_tx_control_bfm_conduit_tx_control)  //  output,  width = 8, conduit.tx_control
	);

	Phy_inst_tx_coreclkin_bfm_ip phy_inst_tx_coreclkin_bfm (
		.sig_clk (phy_inst_tx_coreclkin_bfm_conduit_clk)  //  output,  width = 1, conduit.clk
	);

	Phy_inst_tx_digitalreset_bfm_ip phy_inst_tx_digitalreset_bfm (
		.sig_tx_digitalreset (phy_inst_tx_digitalreset_bfm_conduit_tx_digitalreset)  //  output,  width = 1, conduit.tx_digitalreset
	);

	Phy_inst_tx_enh_data_valid_bfm_ip phy_inst_tx_enh_data_valid_bfm (
		.sig_tx_enh_data_valid (phy_inst_tx_enh_data_valid_bfm_conduit_tx_enh_data_valid)  //  output,  width = 1, conduit.tx_enh_data_valid
	);

	Phy_inst_tx_enh_fifo_empty_bfm_ip phy_inst_tx_enh_fifo_empty_bfm (
		.sig_tx_enh_fifo_empty (phy_inst_tx_enh_fifo_empty_tx_enh_fifo_empty)  //   input,  width = 1, conduit.tx_enh_fifo_empty
	);

	Phy_inst_tx_enh_fifo_full_bfm_ip phy_inst_tx_enh_fifo_full_bfm (
		.sig_tx_enh_fifo_full (phy_inst_tx_enh_fifo_full_tx_enh_fifo_full)  //   input,  width = 1, conduit.tx_enh_fifo_full
	);

	Phy_inst_tx_enh_fifo_pempty_bfm_ip phy_inst_tx_enh_fifo_pempty_bfm (
		.sig_tx_enh_fifo_pempty (phy_inst_tx_enh_fifo_pempty_tx_enh_fifo_pempty)  //   input,  width = 1, conduit.tx_enh_fifo_pempty
	);

	Phy_inst_tx_enh_fifo_pfull_bfm_ip phy_inst_tx_enh_fifo_pfull_bfm (
		.sig_tx_enh_fifo_pfull (phy_inst_tx_enh_fifo_pfull_tx_enh_fifo_pfull)  //   input,  width = 1, conduit.tx_enh_fifo_pfull
	);

	Phy_inst_tx_err_ins_bfm_ip phy_inst_tx_err_ins_bfm (
		.sig_tx_err_ins (phy_inst_tx_err_ins_bfm_conduit_tx_err_ins)  //  output,  width = 1, conduit.tx_err_ins
	);

	Phy_inst_tx_parallel_data_bfm_ip phy_inst_tx_parallel_data_bfm (
		.sig_tx_parallel_data (phy_inst_tx_parallel_data_bfm_conduit_tx_parallel_data)  //  output,  width = 64, conduit.tx_parallel_data
	);

	Phy_inst_tx_pma_div_clkout_bfm_ip phy_inst_tx_pma_div_clkout_bfm (
		.sig_clk (phy_inst_tx_pma_div_clkout_clk)  //   input,  width = 1, conduit.clk
	);

	Phy_inst_tx_serial_clk0_bfm_ip phy_inst_tx_serial_clk0_bfm (
		.sig_clk (phy_inst_tx_serial_clk0_bfm_conduit_clk)  //  output,  width = 1, conduit.clk
	);

	Phy_inst_tx_serial_data_bfm_ip phy_inst_tx_serial_data_bfm (
		.sig_tx_serial_data (phy_inst_tx_serial_data_tx_serial_data)  //   input,  width = 1, conduit.tx_serial_data
	);

	Phy_inst_unused_rx_control_bfm_ip phy_inst_unused_rx_control_bfm (
		.sig_unused_rx_control (phy_inst_unused_rx_control_unused_rx_control)  //   input,  width = 12, conduit.unused_rx_control
	);

	Phy_inst_unused_rx_parallel_data_bfm_ip phy_inst_unused_rx_parallel_data_bfm (
		.sig_unused_rx_parallel_data (phy_inst_unused_rx_parallel_data_unused_rx_parallel_data)  //   input,  width = 64, conduit.unused_rx_parallel_data
	);

	Phy_inst_unused_tx_control_bfm_ip phy_inst_unused_tx_control_bfm (
		.sig_unused_tx_control (phy_inst_unused_tx_control_bfm_conduit_unused_tx_control)  //  output,  width = 9, conduit.unused_tx_control
	);

	Phy_inst_unused_tx_parallel_data_bfm_ip phy_inst_unused_tx_parallel_data_bfm (
		.sig_unused_tx_parallel_data (phy_inst_unused_tx_parallel_data_bfm_conduit_unused_tx_parallel_data)  //  output,  width = 64, conduit.unused_tx_parallel_data
	);

endmodule
