`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n8bQ9Uwx74lkZU/RLMpFJvL67MR6yMDyhUTpvw5UBC3Fle6VhxJb92Lbxa7sgSOs
d6oEvOaDQYj9PypwTkrCYJ2o9gHXCvS5DC6eCFAPu4qB31AJIlGZso2M13pDdkIZ
jbqXa+eHpjq6OZPxNpVvcAUVUn/4csC0Fz/EuxmWiJ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
ryE0QC0Y/PmN92vU3lRl5qz/Mpm8GwoqrctHal2CogQUJA6b+MxumyAPop1Qk5qr
kbm3FeJy6RtgpieRY+EdgTZ2Hk6NzyDsi7+5X12vp8VFRW/4IVVjBR82G21HAV6z
8VDQjF5Z6Vd7CKyidIb/0Vwm9oB96U9CV00TWjzrsK5tWiL6JnhevvVCipaz9GD1
ouI+I/VoJy9HT3fX3rKdtYo5h40J72kvbGtJiIb0Gx/bCjDrEi8gXPixHeU5mE6Q
s3QB1zb1pZBOfidkQ6q+1KiaARYLQCT2NIYnn+rFCLgETWbd3iIK+Ko+fqzNsrN6
fizrLpLs1VIDOwoLRS5lnuFwRUscsXlQi4enxAV+CVP6CxpVtEq6VOH3cTkoOPdh
dOM4sDjVW4iq3uD4JGdD5aWqbcl+Op3A1vSzNOv4VEw2sPvCKzATuIu8BSad6ZhJ
PUlB4Hm3em3C/wa03oYrrBTtGjo6IPBjIOtw22yhe0qrdz8pxSZXgRJbv9Tk/6/H
C2bu/rBOP9l3B2/S502j/2RPEVslY9o/YLFJgzkFJoIcdkNhAdORQIHOUhCjacB/
ebxVQhY5ForR/+TxsB4NH8fEnvUI0kJAxbwLqN+ZbplqIPSr5GnzQ9fOQTH5L/UB
I2Bdl/53zuuudT1wnSADXth+7kYDPypnr37lcOxP5vADJ+iKWkylBunB0pMLyJ02
PMAlB5WszoVPQESzlz0j0TtHg0DvqBc6efq3yKqabyp95nrleBUIfk3DkcZeni6n
yRXtBFHLYJFteAf4odb+oRgnWeeobnuM5Cds4pQXXTT7DyuRkGiEsDXC0CSdU2HZ
4WWBY7t69/aaPzxDM/ih66w9D5oAw+aqG3m38USO8MvYgo/8K+qWTr3q/Q1zbLMB
VLKRugQ3OMxTbyueCgwpIuAM3BjBcHz9G4O+dk8EMeqr7gCqxu2VxFpHEKf+Fgn+
+48h/Rp7iqyff8mdznLZfuTPMLwR+9LUdvmr4CDy8vc3miBQtsQOERDuMFEwDRP7
8KWT6glbCgPGtrMJOwyWuNnc7B8kXKPNnOKSCVZlDa+jjbdnbEt5xfiumtL+IVwe
B0KBGHD47LUfNNnQhO6F5y5JvRya83im/216ZIHaNt02SgpCMwuHd0eD/a+fTV2x
O9MzKzoXQv2SoNFMFI6J+Z/qn+5rU5VFY4A8sdYNKit9ZQNt1t63PZdIKBlidMnE
6MhCfy/VtyJG9CBL3Wu9o2bACWD0X28jFRyP02sYSazt/cdOY9I7+kEi1wpefQ6K
6LkTW7MukJ588jFDCLlRLr7nY61AMzb/l8UciziXcPhd+lkxKFmSOpdHfdO46AjD
fuULezv2TzC/RWKBJx+atGrJHEUn9bqBIYoYDewABRGt8VQu6nXPtEMpyB3NZSTZ
iFTz8+BxF6kBE2QQMqW70eA7ItFiK2CCBrtFD40jDkNnG0e5rzIYeDjrKCG5pk6K
LZb8nBDmGig6+FBlWgFZIP1cyxQ8sTKcEMwq7CnitOJeB5czjcAHuEDknGLcAGgn
U6eo1kim++/OGSrHVGPqbufpkjLZ+7O3lBNKyy49o9eLOmilWd/3WiSRILiunry2
4mnC4KgoSMF2mdZZ4BdoQEua7I644i4LJGuqkztP5QXkM10geHEriHr/N5YG8rEY
lddfcbY0JmMluMiDaxnj+8NVAlo7OyfOMtgJMH0qeahDZOvcgQ+QB/TR6lObdfP0
GSIv560XxUbGp5PDVYGyZIBW2c5fBO9C+BoGa75AKnbgHqdwhxCLDWgkDd0Fquwh
brjTqwnGIa0YG9+uEqnyxrxPXyl3YqKXOWNcxWHY1zN+RXVeHuHeuu3O9e5ePZiK
Nb0uuP+0ktUjZ/55SDqefUMIcZLRlUFwaZZDz/8Y7KPXGkxbnZnuTRD1/ZLtiy43
BRf9EUYwoWHtHNnV8vG9z9wsd3eW3xF5i0LwzvJpLwYnUBC9M4ed56wKxepU4EzB
7AERaV2R0AgkKCfkZvkmtiG/eVOnOprKgxgesNGMz6KKUK/3Kl9X69ubT6Ecn3nL
RU5cWnK0gtrwDCMHbjTmr3H7BL2Fw7+7+4YuuV3J7V1Lr/BOazGd4oWlfXsLxtBC
jxBPSXWFby6Ib40ceM85W6opO49gEf7vTfyFYVNX3p10awJuLD5O1MdcUQ7lUA6Q
kGhbCRli4oGENM12CjF0SekLa8PcYJ5kON5FDALrS6b092L78HS1XB+R8hZvdwbw
/P4Fhdpo5WXeNSDsK8+mg0OUE8c+bMu1hVEw6Bl6HbF8mL25i+qMwoNtWXKo7NL9
y9MnodNYetehlyH6e9VhEfI9Z65cMobxplSY+pBK77LGafbIOhNhXY/vEpXVqB5r
aaYM2zZL8azPx+aLjC+tL1RTeJdlqH2KNfApAu5munt6sqiIV46zdqOGyG3iU2dg
k1J/N0avlOU2x11aA6501HGFW4rmyJ3s8BjHDIyfcOLFrsiPKR3Q6gc/HzP5bN+W
nqGOWKpo/PJK92QowC7eHE4ltfIP+GyTvATZS96mJC+A8BD+iSraQXWRlnebCdM2
LNtHYpRaFqzjqBUnHsu0YX5DEFtNHahyNEmwEusXmuRgbzqYiVNgxa+14MLMn1+L
ATPAf07qvf23bAOmQjCNAjBfrHmqUrARLDyRTu5ItQDqZrm3ttI3veqKLbYjj4bY
wu9eglABKyL2dQTy4L2vu8DM6KwJ+baU3kx/y2rlgJ9mxX3FXWXdqsW7jcYymhdv
naAIdrNBEwDXql0jxbOY6EaEl3VF/936pjhZS7S2U83KsqtNOoqNd/b9DwNNqsoy
ijzohycbwrPuauZX0RyTnZ7aKkMqnZILGJMAk8MFoL3OhdhVLFZggnSQOa6xRF2y
3oTLUU5cwQ13r/bty2HChRrODFWQs4Q3FhssggsVv53Bb2J/w4GB0UDCmHLIxUK9
RG1toNf+REFkf+U/wZUOrRum4eRZ5bFb80H/TazvYcb79HQkUAJTpGxTnQkw7y3M
fvKsA5IZ/6lN/JZdxS0hlfn9te0lyfsOI0leyyKtcRP9t1zhH8ovkKz6m75frKK+
1VgrwLU2/3N0rvrqiZp+VF4yjNXHeZceJdSoaOv/fK0xGLkkErfmBHHFzBTgOuaj
dxS96sU0rWPy0faqyvHZtNweSn8pXzob7LC1F6Ybr5JTDUNf9h9v0aXzcTRl7pHp
HhA+upFb1hWyX1TXh+dBTFusValVaWszR1o3f9riwnVlqNrEWI9KurZwS6W2h6By
EYO8c/+M5j5utOheJs+m9qlmyr3cIUWjNPQv7dwDBmUgymvVKWzljVU+waxQtUa6
pGLnVUYLCT+HL6/e/Vnjwogh4hAo+JLvL5it/WMX8Nvrv0qlOCErrWAHQL4zY5QU
XaRn3ufPaLXVKEQj6J+JeZUWCiuqaKkzbTtGbCRsW8bu5WySuepnORU19e/Q8qhd
N6Sxms6pMdIlLjIgACTht4+Hb8IF6HhJCiua5bwVE+tHsLAMhbT2kD4hrJLQcb+b
wmFcMSBMhPv0EDFMtqw5dw49yd1BuniSKO9bfHZt7TBZZJK1tplxdLoQSr1Qiz3i
KIU+NoIegiPkUF9TdK1VD6KBX0WQRq/MNxq+qb84+xBWiOK9IJTX1tcjJN/LB6ca
AxcuF1E8dIyUrq+zpUG39uhI2O2TTbHzr+cef0fqpbMkttrHTQZWY7DTCwrsgCHX
Yo+6Ofvmdysh+pjcA68FbsTLe3PHJtH+gIMFabtNlpuUHqieQxhlnCPX6pb/icKj
3rAxgFxqmzpvBmT28DJEFts3NIKl4TYMjuTJsX9//Mu3P9Ha2gTCnYV4MK56uflN
4H9o8enWPpAjEpwIAIqabjJUHyAAz/6+Pwepa1ToKhlFtuWue9do6VuRjISQQjiU
YTJjSdhzSO+neqghq8FLIbIwGn2A1+hfoUEieW+1R0DqEJN3OCv1ligDXB1+s4nh
1ial7xwE8stypNynBGtjhQ==
`pragma protect end_protected
