// pll.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module pll (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1, // outclk1.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);

	pll_altera_iopll_171_ejgq7kq iopll_0 (
		.rst      (rst),      //   input,  width = 1,   reset.reset
		.refclk   (refclk),   //   input,  width = 1,  refclk.clk
		.locked   (locked),   //  output,  width = 1,  locked.export
		.outclk_0 (outclk_0), //  output,  width = 1, outclk0.clk
		.outclk_1 (outclk_1)  //  output,  width = 1, outclk1.clk
	);

endmodule
