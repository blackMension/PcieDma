`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tMGwzOmsUY+TSOw7aqAV++kL7VMjUWUI3Yflb3a6viQhXVu962tS8AV6/YFMfO2Q
yFU/t5IDwDKUC1GadR29FmGNIwztmRI79ZFUCVGkBAXhKVSAiHo4J0WvtB7Ys5Ac
1BDEU/jCVgMWPQOUXk3gF1jkiYRtCOfcC+MeYmn+qbA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749616)
YWRwnR4gqfCeEtK1pYrgwwvFZ0YejC2TAg7J0VvxbfPgfnlTkHt4Hckw/eifURxC
kNZCwqSDsKOH2ODPtClKsfplxZ5iPHBlICyxYypECWjt8OT72RG5CrB+IzlZmKk2
0jTrEcC0ge3GfuD2w5bu+9/EWxidi+Ikno/hXUZmjrrqur3JAL4AfZhH7dRelGlH
ch7TU5q58C/xbk2cytPzkTe1oBjXhp2hp5TFsBpCfOtUXBtuISwkr/W8iecRId72
XGLVwsAV+6PijlIt9Q4M1Lt3hjC+pe3Z6NZIh5gSqcTddvfY2CAgySd72TuaHGf2
eORBJZS+VQ90a1u4q0cQJ7ijC2QkUw2FpCXvo3l6lhRcdrkVJGFLHPzeHE0ZrfLf
Tjg63UanqBwGe4k/Ob0R2plsq7/LoMTW0WANWMv9e9rYteXs8N7FcA5066KQcisF
/dcuY8gL6fTGPu+GydlIeOsFo3M8mKNXP1MewEuR4dyrDRM+s5WvGrnRz4o+3GaJ
nhA+o/QAe032ZA3A1B/RwvBnwHnoAPYZwsWBlqvYn3HamqwTNHPq0eV5r6B2xa3Q
psZw/CCVRWKShJUtDBT5cOqa9JE/owofQNzzbE1ur2UWqTscN52RQPg1zXDtMr59
LdXDoFKnVOuS9c2/zocM7i29Tkh33bm6RW8165Q5lq6FL5s7dmdI2wjaNmnYSnOQ
TExLaAWKEVd7ldGVnHHU3LMFgCc7l/TMpn/jNR2E04KVIQ6v92VKTzTYQmB+rte6
GsQjkHopYCnaucYvaNOuPb/3H45HH3dQXGGjgLYgZoVO9WhiCdkUmvPO0phPiIU1
Y6enRGCO19gUhIlRAdpj824SeTX0toFZTdZ2SjfDYpUJBTYQjGNqQMLTf27kP4Pg
3p/6lbYYmYVkt3pH1/ZR4xXb8n/lHOqa6c4o9V4s+Hhr+KO3VIaVDUSDiwmHK8gO
5O7uBvdgl2fevVgkO9uCwF6XJTamVI/nctq/PpaXQtP2v8ciV6jytftJOqYXhNYb
GKmOMUACijj+yLhwXpBUUIla7TEW2MeAoDEv2sNAWe7foUZBop3v2PUmMDYzXJ0U
+nV4uLRq3eQ8pOx2A0EqtrD9Rlw4Z6Pst1g1wjvvR/xHO93BBCbbrSAveLiEAfjg
hznVk5tfpG5fpNTiE8y4Lvrk4DzNnTEBZEwvI2Wz0xBKfmdP0I5xO8zno+wx9mGn
31aUylQvjUMIWht/rj9X3K18/c78sQ1bmllshv+ompvns8MQu09M7EIIaXmnI6kd
sViE0rSSV/OTu+swl3qhYM+q2YxecFZfnU0X9Ilf7bjFpO8UwH1w80nfa/gv0/RA
0Y30OqtYZUjm8U+OAUd2cQHIAi6sR+HSSmpbgYIU4IvZTn6zTjnKcCF/sxiemm6L
YQcSybT1O/k+l4iL9WbVlZDo80b4gHVc2sQu99IuTlqnZmZUikvlqkkmn3pkOihx
AzMQ4otTIOIDVW1kdWY6YCziQ6SJWmKHCm0Hox5FlFAo7jZKtmU9vJm8sSUWoRqG
5QI7upd9DJxLrLzWsEf2+SQk0ioirADmC9NiT7H7VV9f2i5xerbgWcsm4//pjxJv
QN+C28VnbyzaXuhVivWgjqvCM3ECCz1eW4hig+gZ6nPV8xfKL09nO9h7zcLzH/Un
4yN3/KVk1f/f2OhVEA/fNuWD+x5o6kU4bzQWFsUSeT9YmfG75QRp/e6Hyd6rymaZ
C2Rk/wtiHJMbkp7XpI0hJrLhaqTLfmTTmB/05XDqBupwBIjZ6X0+x99XocctYn7x
Xgrs1++Mn/jtaGpLg64HLd6mVV755gP8jYCXwAM1JZWNkdCU/ji4Jq7NTPQYs3cj
dR2fEn7t0sWztLQySfnpJ7MH/aozd2WOJ3UcjnyfIDp+hF5OBm0cmD9v64RmX6Tt
FZflufo+eh07QlM/S1GyKgS80aBKr5hO3aVJH0322xyV71k2GN2QJX+aR2XrVL4L
lMUO9ZNmJ4oHDomCqdpj8l6dqnpZtRbR3J7r8OKXwlnFyMpBK+uhzKXQhzbtNS5V
yu71xcO6neoPBf7Aalsle83zGraUWuO6duRGujzEOgk563CH1A6cwdcoGYZVXCWv
fEtCcgToDKP5/ZutbkcOokkpESkPt8usYsRowJ5/XRv//Fnpfa1+Wp1nFykVVHad
+OCiWzNBM72i2Yz7O3qRqWuo7E0ZPL9b9YCWW5jKpfVOsnnjYx19U93kW6RddD96
z9pY957cP0Lhi5/AlCQOsEfIPtEq7yqi4IhmgNHczn9gPUeDR8tHE3FLPxUpGJmg
XV3ePxtfqDuiWXNJ/oM1xhciAolRpyQMkb4GzGC8S2qjZkJqwJvMO7vTem0U6Hez
fJTO3SzCPh1Swf+JYjltL8a2DANs1I3A7VSCXE2U5YzMC8SlbtSDQ5MWxLBskzvy
WnvHRrDT7lrHXfqkzquCmyB55I6gl7oRLD3SPTkJGaAuBd+OYdMK4f8iYRUclhUz
qdOkZiaP8fm7xM5ZQkcFoF/VAKP/gzMslsR/X14p4kw9B4FdMBAi6PIfFJJKNofb
3aNCA8QxBLVXS/Vqm7WbQy2vDiqueC7YTT5kEuOtipOlkTRqcK4eXXh/rnvPhWi6
wf8rsxSPvKKhOyKyYbuFTZlI4zluOafAAtRz163guEuYw7xEgHqe11dHgfZB5x5C
+ZOiKTOVq9j/DhPE9vHzCHt8xuhwdV85oShd2dpvI8Azv28I5gOiNuccwyAFF01a
B6sIQXaR4CwtLhtk9coVTJu5uzQKMCg038NL77tCMvpMMC+k3tGO0sub2C5rOcxQ
ir0cNGNO+WVgt6aqqUOTOyYg8YD4nftCCgb9g7iVzDXnb2ipo87sLruGMJfBDBvJ
ZVqTzCIbpffAQjqbMGp1aPFd0iZsiJ6IJfOdwi3Z0p+bQWaj323D1H0OnjG1Um16
tatFcg3nXAyXJT+GOCZR7uN1A2uw4W/tZbCC37vMjnr/KTUkAgwM/eXEx8PArX2U
ttIsbyttzTwngs2BO4fUE6huNZEHwAueKVqEiWPeG7cgPa6i+mVAes/6634yjnqD
TqiG83QvNTCjgNnyN0/qa7G0RTbqparHiWWL9OmPk7P03GgX/TTg4VsMQf7mcF3b
ZpqKW0ts75O/O9EqAiyc+fAXoY8DWx4R9Kbci6LBJ1Tmo1KCv6shGqQ4u99Lajwu
BgmUYYxcI/Px2AU3eZjzx1ThoPJoS3W1rOnGI4sjLeLkWLHBEhs6FwydJOOEpA+c
GMRS7IEMz2UCHCT4rRYU/0KGEIzqFnSDMPJhOsBqf70z+H5nm09LyjIfSmitNfae
Jq5JvOZgaHOE/QAcPb++rSzKHJnLoLLaASDkIVnUZKEPu6sLsJPXQKmBm9cOHAm8
1mhUoEt0pZNHaQyCyO5jhHGw68Qp5IJ4ozM1RrrulMjXXIsoLcpyDcae5A6utCJr
WFZuLhHcTHZPKTHeF+3iau19EDwvSRY8H3uZmuObLEyUcV1qGGrjEDRQat0C0eDc
iD5Z1iyINsQPPfRzKZQWi5Ml4UfCe2yMxO1sqiN1MJNO9NYyK3MF132p6OUl8Fti
iQjiM8SbOvX6IyRqzM+Upr30WjwukLXddd+JckJvhbQcv+tLHF7wACMJCUkg7wXD
uj4gLdpGgntpyMQJuDRn/5lJT0CON0KWD0KjD7jbQ6I2t+wuDzR9hmC3Tp/OWm9K
18tDPbEKhShPDunmnZLjYXSSGmI99Gadce+bwfYGhjbzykXAT8Y6ouifowkENDYT
Ud6UK7SNZkLNUQWxcmL6tXn+5W8Gb1EZQ3Wbugin//obD+a03QPxnUSN2Pytk25e
/9cojIRPftNz+nsov9zn4LI0bHJT5dj8Jc6ryKRrX3DTkhlttHjlDGFBvOYbZQPT
iq8KEXf/L5m7ZiV7lfTqWm+aWWB5yP/ZdV59pfLSdfo1mipWBFqdPY8CiKUBvRzQ
H9jUfXmVa5qtFTR/SJ3cHzEhP0URbHKnEh/Da6dOu0ictOGPSWJhEZ88fy7OFeX4
qtddjAjx4J+BJ9aQt1eN60zhOfmCXSF17u85VZhdRv8DmC6tVqAjoJ4hwGZcN4NR
VK8tw+6R/5eSiFW5BMrrGQ17hWdiQmUJOFNsG1CyfPiiz1V4FhWGgzGt4DMZMHY0
uxxPzWkj2Q7J2YmQ5GS3OvyXfAaNaBTqlbnlUONlHBtRDdxIrL3SsgMNFwPx8SQV
xpfIFBGUowVHOFcKtVyO6yZdoYY8dFueo3iP39qPWq/V3NzZFKXsXqrljhbI8LDk
oNBKaA5zROQLjnf61QB7QBd/YFOsQPwaLczy76jVn+SPIYl/aYBzYyYuxvz02oz/
VsfUAmVtatXctps4Jcdj3UZ5YzPFJ0zN8PMW2Q5WxNVn5fpW1pncI4wScpJdIeY7
55M5GHelJDwCqNusJhxCFKEJ9BZy2BBSdW6z7H7PxnmmqO8dh8DRI8rc4RBcdmnk
Zbrwrx2bFEUxrwkjIKufhBZc1e/KyBuf5dQvDmTxc+5gDIrw/OYohsnkT79CQFBC
WFzts0B/wA+Jamcw+qqX20AIfyFLO4YHxu32fHiIR4w2pTuespAJ0O7AzhHxbhfI
WEPF8TmOa2nvoaN7LD3j1eK/lXeHXa7HYCwxMXWe0QeKhSSeuNesGbTKprw2o3Ll
oxb218FZvg7rKQYj2cwMj8hyHVhDkhJQrOcOJ+IKOPY44zRaw7O7qVAgPYzXiDAx
wJioumU87/AZVFkssIRCfHeL4wRI3ZFffqxHWHCTvZ8qMgiusbJDqL3Snq2q3tCG
dbku/HntnAkFhyDiCmtLczItbtTXVLJDMdltXcv5eIT1N2LpgFAMaYyc4fDEKfiC
pLbpiLW8jns/25Mk7SridGPwoPG/7ZtIN1qoq3EMz7arHB/oB1RlF4UAkKrC70AV
DWVXexxuYGrCuipLWBTa+PC9hGMPy1yG6cPj6hfXL0ko2za4zA25R0+AbpQj9rfu
owRfYuSikpp8bWovvKxerfqhX0KRKBY59z7iv3KB+48iDWPDOq30mHrYGPOIgM+T
EnLbEDFiei8xVBg54ItYpKH/tucYwFL2n28Z3YYE/z26SXn5tIiucKJXUREcvcS1
OBpyxiBwykQK2322OXRyuH8Vmb11Qc67G3dvuU3SAuRVOEIBIaNJ9noyS2zrFdBL
8KUk7aM/pl/DUb/UNjl3Tke2NYcKHMdVcZTFXYuAlMjRb9XhJ+9gZgFl6LASzrGs
PjPdfF566Us5lWEKwNiqVeNrNRXBsKHFmAQS7Ci5HPs3KlVhFZQVpT73xQhZKzGx
GnFAkmz8NDBrJfSsMql0t92hqQqbxgjNOQ54FW5q/CQgXydtJ2oBDj+HsrC//XSp
yX5uUwTb1Od96BbD4+5TQggkB1PJQqV6QshThQUWmZUh2Puel08fHIg4xQpHnvo9
IFBfbBIIle/M/Ir9Fx6KM9prVxpECn+gzBQ+EyQcAXLpuN/d0v5tUiDb7BM0F058
EuimhtpMiSy3akmU47dXQ1LjK+Rwxak5+9gI4TIHyctDOkCp7NHAXTH8e0+8j6Ea
L4s51JlSpgxmjrU4t5muLffIaPLJlc3TRIVcjF6XfRhZqBS6ZWUy/7VW5UbPyHYy
OGEnvAkXkVc1hI//QqYvtgumNHYvIkESsCXfO5WsnfqF7Rcn+MKdxOlF6PfaGAi5
2+jINbhMAwom8ukqPGM4AktyDPBU01RrFiK9q+eo8qYUfykwLnen9z9Gn7j3tZbF
tzAnCD18ZnHgpC80Rc5ws7w9WXxON+XJTqF+YJX8nPlX8M3cSTmAZ+O17mB9Uu8O
2xTrVfDGJjiWt2n/eLo8695g9zwOuIxMjVqfeWh4kGpF76uZcxKs2dUGdQ2AwnAH
U5f0fW3fzRDN8vFcuOgSw0Li+Cq3/KUvwp3X4vxK99NmK/WHyjGzP0unZK8m/+Uw
g8a29E95MON6ZDIz4nkbiWJh5qZJJGpIWXwMufimtzd3dc5hqly5oCtAyXFkdX3r
KOl4PBtQdEDOeScNlm0Argr4DtILjQzveVC83OBfhehYTgRihKOO5cteo6eeYciw
YhO19o8KBKEKNCtDeWftJCKKO8IGsPr+eBWClkUF5y/bNBeUEskg7ixo5arbjijz
/Pi9VYeGolaIJjgI/LcjQi7ZOm3V1IK0kIifqMUnjQ9aLG8mWV4LxJTiR1RvuWEs
LS0WQ8I9H/dY5rqq8UMwa2cxL9PSlkLcQd8C+jvMhUHufOgd/+7R5ZKoOHaFTBIZ
2K2IkA4kBQ2D8nrYIXSzPae5E8X5LHK7hd1Wb6kRAAS0pRAsTrgqqKtEOiMgKD/x
THyAgPdMHgl9su+P9aXDiAThv7RE6rD9aklx0O3crJY3fB61BVA5V4YlWzgKqayy
jc2pLJ10b1WR9SIibT0qLCY277BNzXEs3f7vCz+krdTcjKNjsxXweVY+QC+KYWyf
XwGFh9uB8OpKINxlLbAGkm1eXBySritC1NHD2NMXwVGrswe3A0GRh8yomcPCB6hP
LX7WaOGhyy1uzyvZSNwgLFSWlnhfpID9Gp7uMd0C1x26WBX/CvCPa4mQMlRBt+sl
cWdRy0SC2RpQw8SHcLpWXYs3WkQuLHuGeYkzcYh2Xle4V7gVFu0B+wh/XcbjeiLD
eKnaivu2oAzy5DubGG3L658m/zw5Rj6+ZWLHSml6xUV8G3i1QmIQMBH6IzJL5ks4
8oyAtbYju/T1cw0ZGvNCpnDaSXHyf1xqpjovFnBwRw1DteRWiCKT5o1W9u/x9Em9
1ECvQuRDe1iLxjFnkpngPuqAssGM6bR3CkYTgk14jQoMH9UaBVL/DO06FkHu3Wlm
vKJ2PcNKiLuL2/XeTIAlIQw+UzaVI95anoveS+loK1+L6J/ftaWMXDUN5vnfhlZT
2kdQr66LZ/EnNQMKCoPcQXY+e28gB5yfJQ0otL1xV8Lw1QL2ZZPn9YK8Gbq2i+C+
Da4fEa/mR17C6AWGmbng8lIdExzgZ+Ub4is1kvnAfZYRSmrj09dy4qG+FhUO6JWl
/tWv6z4faacou/kRj1bEsyZZr5XiGDMAPDtDRUufh38ik7ePcalgka2GZBCzlMJe
hqJTbA18Omzko4TbycfYakGuj+iRjciVwexuUfVhXsChZJQzcn6DqGinLNix4NDb
pC4BwAA81LYsd3shRJ9u8mK6U5zpYqa6YP4lsqE39mdeIerpuT5jfxhAxpX4C6Ah
YFDMgLMiLWn2W4NuOb0ZaI3FlJPyYy694Ugiwab4/xApmZgj427buS20rujs4EhD
ruHOtCcMwOYqq3KVE1KfR5523qsTaxvjaTYEb+X9ALYmgN2xNnQlMB/lej3hTUJ5
hzUz96yDTpmzofKygft4c0yiGpY04hJCE1oMt8lthjCB0lhAazP1OIiPYek+ODED
54Inp6gGUn0Gsytu96Ws7o9K0f0F2iEqNwC4jn1o/M7Q8X1bNQLrd1VtZNNgCMx2
0SBsk7tRJ9QEV0x4qQOEkQKPFmDz9Fj+iYpAWDdGeneDxrehzqI8d9NlqeviKDlS
rS1a3yF+wmqAnb2NlIkfmSUxZW1buUa5rmNze1qgI4PMTOT8pEzr1uj8qIDRM0d9
gvTI8xU5pmzgb3O9vGQC6iRKPJR5Iid6B/6+ea3rTGk04vsopoUhJG6IrzXqxMVp
dQiLPKFIL+TVP9NaLQDFRxMMLiEqAau5pD+JxUowAXJ8i6W9sPuSAmsbQJL138Bx
E8WGZ/Nhr8EujFZlECMfvFBAkin9CkYnilCoxwtuwVeaSRSaEsH1lnDUo1b66+lf
H1I3lG5wcEs3ab3Pd7lZrRSPqimBbAH7qqsLNt5PnkBS6p8RuyumHGrMzsA79Woj
o8P8FfdrDDrbc0Ll5a+uhvigzzRhnm18pzGYpex77OUNigPUQmgpscMAPz3sIAqc
cok9w5c4hC4bnJJPXFvZ8YPWsTiY+wfODlFKgSpTXeJvRaThFHe/K9K1NPwR1kpn
/CTPd8ARgsQuF6GvWVITXRlbiRGVGhjwk7+r5Cu7eXvvhz+eaLfYjZWIKbTceQ6f
MEQWDaEHuWqNGCFFLWfO4mSO0MfEyh1k/HHtCKaOE5TSryOym4mSe58s5GtUmtMd
PI+osc/438NOYwx4251ZEh2ITk2P2+ATIbYPygOK8hvXbdg0I1svCTWo6KWSsJ8X
VC32NOZKDVxcRRwp4G8dHdu3EcNyjk33KlUn5B0Uv7MFzra389v/WKf+8UDdrnTv
fTa52YnxKEmcKO1x9MPVBcgGgsb/IGwiTRpjhpcGKYd8NRPe4jL7vFCG4CWg2eLa
2LZ7oc5tCLCIsvPAd6eDNfklXz+vmQ6/pXTdvLp0yE6KMy27Bj2boGEZKw1q7NlM
rfjnS1Wi8lkTdM6eJDDP1aCboBP4f3JSDsS5Tr8GcXe2eMDq7+3yIyE1SGVVlpRm
9aHi2t06Qqs7REd4FPhDMqAnNmVQilvmwnVcAx3BPZP0CpV5cQgrsTHw7VrUlZDY
QcxA+KP0ldZl3bz0LArOcf1JEBm8G4gaG1jzL6sOA0qnK27i5+hC9GAaTUbAujhn
GtdAYxpYdE6GnPWv0G99BRKAbEcFuQ6ObTVVfBRhskp1qZg+sOt3sj00zSa2NRpt
8NgYxgUl7u7a6wBD4WsYEo6WFpumwzd3Hmr+Aw/bI/bo2uOci6IJ31Thi3ZbfUT7
3NhoQZQmcr2Pc4LE7/YlqTC6eJayvIIv0ar++ISD8IJbkGCvbsHGKg3dDrwf6hqb
31kUbyXWqTczG01pxyPL6JMhj8eWBIdwAOmdTlL/nDdAS+wNEhSGBdD4tFI/HjYe
DjoIbXsajSXxb3mXIztcqFCgjj4HiDTXueasjA4zNr6OiE9cMsfNPoxv2tJmwgvQ
R+dU7NWVQc6UDOGu+H9WGuZImXgg1+JuNoZHTVHiONC1Op3gbR+B4TcJlEAaszim
gykHnFofAmGCUdCF8qfAXuG47hG/oEqPi+ryiO7TbDis2IU7RR8OgJEIjQMdCr/I
vc3X84t+ZgQ9igJR1+HPbcWpLvplo+bJv36UGUm38qqBSedgqC3HzUf7pRUWu4kJ
BOlBmTAGak7EswpZKtqZWUJ2XDC9F8AfSn2ivLwmhsBVFMbRolZjcGLDvEQ1yfuQ
KzOlwP9Aos35XEUegIWRi5bJqcfjchiKTQ9LdmVV4wITR1zmGD/Z+zWC4Q/ackF0
KVGo8S5t+hMT3qwIBc80DLBjKEAISiEPpu6gNDkZ/c5BEVRxrKnFNJD2M3UzSas5
Pt684pilQWydHvjmeQDsIejNv4q8d9FgT0qbzhutrFOftJz4X5g2MHSzAPS1yUU3
mMs1SnIU9NOyhiSfOm6Jk0Of9XdOBkzscQTs/CfwEjka9vR0+hJfB/Uqit9++fJs
RLRlnwCmn5BmEl2tPEOZsTPrBk99SJ9+l9oxho27YPlnhJYo2fIewJxfmGIZGDcs
U3TgLxRvu7DGz4eXeRIJ+NVTACg4Om8ozZQpvWPqJvr1+Qucw+2cDJG5YGvufvAv
/kiJgh7odoEWCqfgVC/snXYuvQqbvs0ICytmgUhh7Ry0hwZAYp/HX4+nz0d0JMX6
aNosebAFewiBaGgfefBejBFxfBMjuShxC8Sp2Du/K+GFORZUDbmmDQrXBrPiNkWv
3N2oVNxBnszlan8Kk37IworOQwUYiJyUFa+waWRCZa4Dxuz7/LoZnXxzs4kmsJmg
xkqGzqnZhXJ2G0NYqgXrMfjXyXbu6eB6OmR1P5ndcHGEvmTEBubHSPxaykzTpSQZ
hpH1nrmFqWCGHMzkdyJKGXs99fItoCXRkUBB8smb8juwfraoSqU9Vd09nv7PDETc
qOBSGyOm6gNNS1VaCK3Ck5xnVmoIq7aC61LT311BhjRCazOMqnmQNGKTCUFwfuNP
E9j0QfF+1QoTtdpwOeLzJzJ9cumg1f7kNHXwNyLIooLWuVv82xRk+TPR2Voa3Tx8
30wW14P6YKpnz2tVEZDQmkWDkxY+SFsY2zn/BoIImhObpEv9gI7dpxz3QyZ1hahA
KCOPdY3ijyXV9oTZitHGl4vFXunmp8hqhpDQOa9UNKvFzjiiMTtOzuRoDZEyD3H0
fTc91gyx6mWmHNBUppefpYm9n6+rhl+vm9LnMUf4CpN01V0QSb16eCQvIFlSovKe
nyyuPdLQlcd+gR6JHWM9BNeGYNjuH/Tc31MKC/YtMu8s39vwIGdmikDD7TFQ5aFm
1v3fEF5T/Kj/LzL3ch12013MYqjFkr+FLDGwyr4Or3n7kqS1LMGf5wOF5UXuFjSx
zceuq3kArTgohmOaFUJzSctvx/kihrNdsIuGctTgczNJv092n95i7KY6tVYMS4zW
jLgA6ElvARfRw0NHdkg9VVOenQ4QytnZ9CxOpKb1H2S2MZ4zr1a/gUrebby7cPI5
Mo6btfu4xl8OWtu94aqplwyTGFKl5S3NKN9YztvBktUP7UHs/5mC/QUSm0R4RDO4
KPLxuamyjit1DITT5aVACDqXkIYl1rRht4nWNsviXDmIu0JmuN49LdgfzkgkMwt1
RHF67aAzj0Nh7Usxqr+BsVQL19rYeccMNW+g1tgDA5p6oUl6KgYKi3X7ShM1L/Lj
pZmS9jK+vKBTrS0NUgT7MC6X0YQ1cIMyJv9dPoKz7Kh/uzQANBky3+2Ao9y5P6S1
hTf1bH6SQeUo3POqUGuocCMj/wSUxmK1cbr9Zq3VbJIOxFSItvU8IgdwX0mU9mn4
xmtlu7PuF9FkW0aVcSE56fue+K5PuZDOICU/W05B7AB+YXJrv2xtoAMcVnWMDEa8
z1/di9RNu1X5vgHK8euQm/Dp6yrwe/jg8WnyjmCMzQOZ35dBnK13vhyeP7fDxDo/
EgrDIMil0RPKeWZ6W3QLfWvoBBf+K3S2KhEmMB0108KElr3ESYa5LhNu1K1+ok5Y
QIOk9PQYVCRR3ZL8bJlHVqRq4NSbKJtMnh80Ngc16mGYi1TR//At4Mwe9TuCvXOt
5d/8+KCqK8w/2ZxYbo1YjVT/WW3+7gAkupECFSzpvHXS6J5Q9uX389LOgXEQcI/r
3/goumHzrrDOL3GpF7A46ccNADXz4p954Btx2uVDoKLTk1R0mL0W2hHwqw6Ou4sm
HiGvydjy8ViQB0gWbPm5MEau/xla/VD4Zzt91XZjxV8sZyY8u7+Xdi3sMn06I9GQ
lZiztac2iBOyh/oIINRinz4nIDUubedWD8RChqRgvhTsqLrU917MeirAc+/ERr6d
/pUxNmKmvmM95azoqO4SEOGdcZjII2Yr+j518/AionmRB5C+6PL56ISnzKWHj+Tj
Sdd/k3bUVWvowjGb568kJEA+mF/TQxmlHWw1z3QGDoxmdz9+kd4o+EUTkQ+DsmR6
r+L2qETPR+anBVBRlBbrprId83mayvdqoYQlr2qPljnhsaLEEglZ5vyrz8ditf5t
qgJi4JZaJZKdpAvnMQ7FHDoB7Q6fWvmGBDqRWv3YNIORLCMOdGcYOiXnrK7dNBmj
UI4XmKL5lNO+8xZ9Dh0ZzpoFW9qp8Pmh7lCS+2x5W+t0J6NAgG0dOYUxxC+w27nJ
lcNz+wdTyyvz9KVmdSRGAgWuUwr3YV+1fMKx7Q3GxstkMqb+dCcJptokzBcsC2JX
JyePiTuct7IZ7GgdKlMSFeKmpOko/v//OcckwCOftTdUy+AOy/p/qCyApVvjQD4C
+HLbzuJ+n7yRvyNttMIs4LHMDSld6HYMeXsJlW7ygMPBeec1Ju6WFvlGzRDaGs99
5WyhzBK3/W9A3rvV6J6Qoc09IjIu4demnpjooKhILq9roTuOx14fhr8o0R8BZS+Z
mdoOVWV0SFQoHwCsb9tpMdXdPXqtohdwpkYL6RnGWnccfYX3I8gkul4F44wwPzDd
SBdHl4xVlzVakUhk8OOylKSw5AVOvE1dcVaHt9nDHNVHVJOEpCt5ieFwDfvu+hah
CuT0Nn2JnbPexMXVDf2kExXcGr6EtMdW3wqMmxSZC7tDBA0aMvFb3JgH2ULZKvtN
66jejS9jadc3Hi4xLmcBIHOFqREcfsmFMJGfHcpNDbFVGbplMmTS2flxd9AgYtig
2gI7jMWWAcEFhcJWpShgD/WGqZ13IUrXCf5JY/z8uhA2XRtv+dWhtAytmYDXwNJ8
Ko48P4UXMcAS5c+yPws+0n38AWfItf1Oac/g41FAAm54k+bOy0HZ23ZBUaKyVxe+
CSse4sOYKDHsl2xVEOK8OmBXbcB3wxQRl1N+2LLHOUI52EwWHVd3f/doPqJMr3xC
FakUT7rwbsRhf/r0zDYR0h06HB/xifbrNABmXHaJRvTnN++3i7apoOtBmnY/5ron
EdJHFy6DviYkbLlWF98jbjvZgzYHDWqqz/ptZl7WV74otKh1tWhK8Nahn6GJMAg3
l1G2zX319ZmOAspuS7x3Gul5X7vqnm9qqBijR/+e+8znRkq6Oslg+D71u65AkZy7
avCLu5IWtHO7KdDCk98Pm2Tl/9luNF41g1ISej39n4F8taPL0Dc9AMOi07IWSsQW
6XpI0J1GH6sA7x3GluNWaxmt0dozXv01jiZHEgp+52sqsGUymo+FQ+N//KqleLTZ
ShdI1dskJqdkyQ2s6y3iW9vDHLWpG/xjyHaUEBeKrvnsG8NPPE5RgrRPCalBPLvu
014z2LrAFRMBB8Guy3Rzo5ClQyFG0Mk3IxrsbOhjfcY3KlEChQ3JBBuD7kYgbTju
6ItRwUcFUAudGykHJoOYy7n8P/yqZWplHaLsLdRT93IseKpWB1QDaneklNLOy1aF
xXjUE0tyByq6G29/365fB+dE4h9Ih88KZqxxhpFajTEj6FclSFyYOsu0WVGtLmYA
g98Oiv6db+tsSlAUOhV2LTC2QUXSeYwgSfxv06Tcg25X42YPwPFwVFC8n/tZmI6h
+wae2CepGFwcl3n2OmyWRRJ/Pi2sCuwZ5y1T+Xw7rbtJTdffXS9YpXYqHFD/a96K
l7htFhBq/lt5LufpFztHuBpxIetSv2rd35t0txVkdzQE4qEnf4qUMmiUCRQL1/Nt
ZFoPJndbB4rE4R4tZFYQyMJIIXEiGs14AF3dOeSxx0lrQ2KrhemKPyS0msoBGEP5
LM+82gM7hEqctvSJHLPvqpvgzUO5SA3946jE6Xh20YjQazzcfFS8EdICek8yty33
TpKs9pKEypjN7iIonVUP8Elh2dixLd7U/12eGmzexwy3HSciSMNGKAwLm3DKOVC+
ArHcjvopYT9dbNr6SmjZAFSYhWesoVTZUhlwH/g8jM+BDh4eEc3ZtSJk/uWvj8yt
oloz/+8u/mI+ze+Lscq5Cx10OsvTwAzmbWHRdhZ+qyWSqVPfsyVZyCjKm1pLeOO1
kQkCzfQvCgMtElJW6hkyhoVF9s+0pQRFbwsZFnNjHYx6g7/v94/dMNvsnskSKQqa
rMiCwftqofxvhUJXGgu2lISCGQogTSQr82lTcRWYI2NAchH+Nr1FACPiIKWqhOj3
IKwirtu+0iaLyF4VEE6uqa7kepAB2k97w7wfA48UYBqBf8Sb7GQTqsdwwqIl4Prh
p8YC2d3hwPlF1ANYMedladQEMLp8Xho+7nqLUARXmc06PwxwAcsjmB4/lwWtqW1X
yyEM6D6M6g4MIlDnVaLXlCfWN+aBh5FWutgaQ+XF4dsyBYEMHwdSUsubg2qwlZYL
VWenrEbq3WGsDa+VL4k+Fy1bByIg4GkB27HAI9TtIsMouJfATITQidb1zorKyYxC
3goIh2TjyugJrQ0Em7esKkR9qlcymDAYWEcApuMjr4qGv+zCupnt+/vTwOKbIn8l
+mfZzwrJg8pICUyevvg1O7dzEwm/g/YXIJPPt1X9EsKJBrJyJsbhE4BW4WNFXm9+
lS+HKYUlag3tDKZ/3KYXZJX+qHbWHXRde1qJiGj3n0v6jkKO53NhluEvxFfODWOV
w80P9jHU3JcbX4Duv76xMH6sur7f6NQPZUcg19S+JPvKJxyg6rqca3H09bMp5lT2
9qMHywhpRSDwmY+z0JBqRBKevQ29RF48BmXsFTkYlJULSsZS8hZmNLCss6FAG48v
MQXYuC2a29ACVIoIoKj6rDA9D2Tsvz4geB8ljfOKj2PoEm/b+jEHsO1nrSfQ7QPt
utXY9W2O++bB8Gs4VOw8VqGlm1IzvOWKIRmrHoi8C7hxskqdGoaPJjZ7TCrRefJy
RSeY4eFC8fnximkBirH/Yd4jwgFfXIvpn5wJeEdmGKEdRr/383PfLQcR113cPNhm
v4nQdkrfAU/+QLczdEHvFSWsARWCJriyHdIUgrekhqNQ868RVMQXEZXZMRnHSomO
fkLljsTdPZfuIahj9PX0go54ixGR5dkhhotyEiiMuG3xtfoT2XruQuJfqE/o6lx8
BWJMpQ3l+m4aAE/Sj4DWutHZ/4oa1mOUMWgwYtrJ6Govn6iwmNMRTLX8Pdx6MCfx
YyEJZHXk5CNWWQMabYMPEr44pv1jFKRZs+i/nuzcYyr2XtIj75R2l+SI4Z5F3jTk
w6SOm+gy4C6YBdBfAOWGVs6siQDKAq3HRnk0M/myli5esgQo88zfsvjJJsCda/uB
iIDrVd2Vhzcrvv2CYY6+7NsS7+7+E2ozAvyUJKNvAaoGyHigzH8+lT2EiTCzX858
NEWwiKpDfVoiDk1A8V3FIELWLL5kgFqTXKst3XkNoaScJofWwkS41xaqRq7BtQYy
jJyKDervuEnHJQc0kWJcIRwZDrnEPUVnq/wbKHVe6ys4mKQQ06eQCZGUglLbFNzv
+SgAuhYzVzc13ioSVn+iurlLxRy4JN0Q7az81A/Y695zeutnS/tYqtp7Pp2Rwpyy
T9mIPGo3d297WFCWsH3REj6xEx9GdSDVnPtdv6KuHCx45EUqM4U5z0roRNqclpQ1
2u2IQP3XDHe7kNB7N5RCeNQzrJ48nSopxbjW7JUyhLqtAaVfj3WXizvv/Z2gOgTD
c78zRUxnau94n9brUJr4F54D29gQNLMmKPdruXQ8hoqDSxcJSTomoz73XXGNDwbf
mLnG4sk3zDdaz+Tz5C0+PKp4MKHfgIGu983tH50KmQGaBvFwBZ+iuYPRnjjrM5jI
pw38hZJ3BAejp88pytIUTUI9NuuQLysaOOib8+oJd4hXKjNDtdOXCfBCZfjBJARj
gXA9zJZtMhV4qG43oxS2tu4N656aHGk1f3C60gf3PntPXQTq0jEwunRAqWrATRE8
/gsJLgChu1kWt5iRxkQrtjtUoT9skQHBhvPYzUJJ0qg/OmYPykld4YIM9B6lVViD
3b7mxOTQpV5TEz/OtacP8g/8z7MqODXmUSHqxUFBB5ZkZ9nzsngJKDSE3wGEM+/r
cVo17gB6N2poAJ7IGPgFa3aIod/WXk9Tp1JC6kyKPC6pFWPL3hq0difuUNck2tUh
ZrbPSAOiUs4p7jlmuCH6jX/CnqGdFKmB3peXsidu7UZk36uYA+uviQi0KRWMmtGX
tX3IKbkSAPPp66p4T2u3bgZHAM2UVT8WtfUixsoIyMQKEDTF3zYmc1iWszjklscX
2tSkksf9z9qFLGVgizLLif24SM07ZBMs0pOVL21uvjTTdsZscI8Frj1kgwznuanU
7cm0MjeewvJqSc6HpX+jRZ9YRl6xFYpEocNecoNx/I1yQzwSa7N6UQVFZkkB8QKH
979jlzIFen4OmCfeizAqF6e+E9OqVeaKPguwl9inZyKHdYHbJtYoHMOUW3TF30NN
1zpj7KsDVFCctYKhc0nnqfVY4Un+XipRej9ZAjf1iS9qoG7AjF8xC4VdDT+OYcHh
uQFBfl97NNk0c8FmS28jkggz++DaY5sBKBJvulGNBX0sLZaujgMQ+m5/BhStpR6u
WuGRenmywYNhKxN42PrRjpswhnTupUMR+vsYY8SQTFo8GsxryqgWzNRRKpZrm5+1
/P3uCFTuxLOaX9nPX/R2E28tzIlrhwr3fK/W/KJcEklMtvD26GISwZZFp7EYGZPy
kduSILEHoEr8fEZKXcvzVRKjg0IZl0zHK8NReKEzuajPwzhsJJqQqWYdopsR2byj
mECXfco63hx7YdfBaUb4j5RgVPAX+hJuAaF33mzaSmJ36p4ZAJfgAOmJbW8OgTP4
FmfNe8hl69FfXcjWuntpJeAWPZOF1dL928BF+KgdYeiEiF87b/PrbNIU23vX+zRf
CKxWBkBm7fBURL/E5ttsCu9u0xgwgBaD9RHsSLgPvNvmbvu8CneZB+qR0UW00QdE
QuLrJ7bObwQA9tiAOnMjwQHdT23hokpig8BocU33DcTeMwL9jq3BotFTVJhLz3A1
GXO9Eyxr/Y1SsDx4T/MqpYr2cp2Hn3pRRN7v5hDaT32WfPuWaz5dOFNQja34/aU+
dSdS77PDkWTI3KeyQsE0wfC7Ufw391s2aS5i9JgOplvWXQiIWpeH5rc5nQEriScO
cMAmM7tf5YXePCttVVfgHHLRUEY5hCYRWWQJwZHw/+Ww6OSfDxQEs+kLhmcBseDd
vw184ea3rtZFXdKo9VGtCqT0Pdvibr0FvnLp4e1f6r+pqX6RyZlvUbWVQkwvelI7
Hkz2O8nPAra7CDTvmFXNsZ2btbIQJ1NYK+hQwPyejMziahC/h+6J9f/HlzS2Fah3
3Gx95JgfCP9Z/B2RPCpQ4dBdnoaknZGERBO5uWuVnbof9iA069F80yXgALGn5CLy
mKImutnIVebJ710z7SeAF/4afn/5UCNnz0+NcYZlDsL4R94giylFQ/zEhZ84tbal
/xOS8gRWrxnrHOvF/c8QATXxhVIfbe5wf6rU9SmTjBiv1G4ZKam00x+KqBOM8CNy
VaXWH1vLVCkOxMbbOTMEZmgsAgI+b+VSPzb0K0P1+TXrT+jhX6uAgSDF1VDHOnSv
Jie+AeEYlqp6haz8ngNwYg2KQAtaM7whBeSGKakoCN8tsf/8scRBcekemd6VSkUX
ePfRdST+7Vnab+1AYJUW/bNJnXeNZu+e/l4VjZhZyhKktjmGaDwSJya5hFs9S9hd
HQMw8beE3GUCY3dMHGtmrq9q1ZyjwA8Op0g+MFD/P/G4m4ksefR/RK9DH5/Q3LzS
m4m0pLbrQtmRlUUPUSn74RhcwQQ6aKyE9ONKIg5+kP6N+yQb1n77xZP/3yyTpvrh
/aWGlGYszJEBHVW3ccwUDJf7c+87ydWWn6S66Hytb+CsjFow40M/sJx36ZAegTXs
56qs5XsVC+OUCO+iLZhdhom48XaSGvbgSa5yOKz1CuQ9jpTYFt3HVZyvxkeBY3Fm
/JbhO6EFUWu6AzV1ZY+g8MHjy0wUkjIEzl5ddsIqwN02nYuAPbJgE2F0isj/xquS
mHFcfj907/0nycwNHz45TgNgGz+Sf2oKhgEnQ4WvhOm/2GVMTZ9ygBLhqgFTjKqy
mx+UW6ih3ZZTqSvHZ6cYoaPx8O0+r5CXsvR5Tzuc24c5jX9PaPMITHlcjjzk25I2
waZUMD1117vgXeoAmjNZh4CFLMv5mwYaGGu29a5ryATf9ZpRfwMFe8sDbGf4pzhC
ZXEAbT04+fqsCWsmjt3eWriJ0lvaFw/1Eieb3z9htUWWOmYfRSkUEgyK5MMGux3i
o4Kdyh3JUjurtVuDiWtX6684rD3UUuY+IZdNe6JqWeokV/HW3XhEe2FzCn1n6KTE
JxGvmPQZ4+j/Q1hy7MUAPRw1mjQisdxm1gxuGbicTHBdYJqLVYuCcgWugbU5Xvqf
p+S9xZqb+oxxLpiaXGJm1sDbSwbvN53VYqMVJqvF5WRtBBM/aRZKRLCOfm/wN0Rg
5mQWAvE+jNMpog/8Uz3msuj5M2EyMFuTLqbSesmM6CS0n3vAbN6JeUtFsXLxDYho
Cw52Bk8bguDVBwz/g1bsnW66GNFoOjO1MpWmQ4TzTg3h5w4AvSR9sj+atC7cMf+W
U8niZIBUvNRvs0jG0+qlbUa7PjQIz7uNYyjEhJRSjlhzGyL6kmdR/+xUsk3ChiGi
3wwz+2zQPuE6UbVn6ezUtmKRfcKOIG+NzPLfc2quDv7m0u4kaUSeiAD5uYSdwXHD
g0f9rWceFR0lE1VCEQfaQBl86EtK2L7muawlfj/WaqwHv4Z+O5zVrrVZNX2DkDQw
M/iVfDgO7HoTfcZnyVgyAiEILBM/fj2DM4l74OKafoXVW63avfBNQ7PAZYl1HqxJ
DiEIs6cMy/vS12P7HcVWb/5/wclisgjs9vROlpazVAUa5BdWhdwRGorMvPHWWx32
hlLdWJKXGB2WXlElnfcviFJqZULQxk5u8tKP91rMey5MccpsjhBIlxQVXIgTyqPh
Yb6CqTeFbUfvW/6swRaoS9YJUXNk48ZboYP6ymMYB3dCtrJKI09xAnt7BnCAcXhO
hjaIzkJg0FQO92fwsuDopbE0Jk2Lz89UdB/smMgChHoTxtqJXNP2Uc3D4159uQbP
MqThCAoEKS/NAECgxG8Y3Gt4lvUPrGPZhJTf5gA9Ua6MwH2aKXp9VdtZuzNn3Wl1
15i16kXxs8eHES73w0SjV7w9Xwtbjim5bDIBmraZQARawGK/S6pWX0+WDOyQX2z5
1x8RQgNxUt+67sLOErepEve1NGcSdTyjESnFb4fAUu8wllu/aUjT/8nHrBipUUw7
6V0rAdFjxTviomMXP7k2+eaZNLGg5L+BRDtwdQE1Ajgxvwy4cYy0NhXsuwjjOsRu
2eMH2HGn7+0zDL8fpNk/WKT31q/sqARzJXQrfSLX0YptLcnQNcL2ZIMG5gV5Njj0
hdmrz6OOYeWFYNWwU+9Hj1Ok5UDfND2ZC27uC3zJd69mvbOctIX28f4Bh35GdeL/
9bcvTk56TeG8PbIGytTU9v06NJfuWuOlaIJ/PsYjcJ88Oi136me4vhw6QKdOF6q4
QvqQeL9mA7OHUrfc/1JIMSvEx5QKkCBABfh7DgEJvkLrxNL6Zb5jZhvjoVmp9ZTm
dl+xpKMsi+zQXvZ9NO9w7jSBP69qJ0sStfAOTCU3hS+cvLLjYlpp6dCLM87Bu2VF
tqG/T6OsrSLFpPCNuxGkKOosqM1g3cY1WjPxtF/QMPzddb41VvbI4GXE1cRF2P1e
sySkdPa3WadWMcSNavXmrmyC6OMaeBn9bDVzhpThrCEaxK9YRSrM/5TQkKwwdsA9
mgwGFURwbzjYws6tcACYB8EaaxjaKw2niQBS+VNJ/uiTSjtvtwy/OcNw0rchwZae
ADJWNu62Az21rVy+bW8v37BU0kvab1LayqwlkWkDH5SJytsCoTG08Xi8HLIPHRCP
dpSH2yT//9v3gdlirswT5E521DyQFzSUXY1CkxS9rfT9fVaTip6uC5+JueddfZHj
W7qiORYTqqyjJfkrARKW4LB6x2TaZ+0q1SeI5+6laj88UwCcX/zodbcY1wJloXtG
WymhPPOijplw+QjnZ+dvqCBOIn+hRZ2myBtp+BYPUX7MTLQArh+PH3uMinhllt+3
+qT/Qthp1ibNI7zBff3Is4KFcIUFqx+KSjgsZlBLQcDkCej5YvTD+bKUfvZoPceZ
/dcEE61GEjmxpN+kmfInBOp0PA0wo+n7NM5OB6Z825KNyaI1z7ZCM5bsNldrK/Zf
RfwovvRlDFoqUnbfoJpIt2T3nGSIwmk6ATEDcFvwv4ACYgEKkdhm2xA7fytiM9LN
BkdiWZxGR50/DCfLW5xZoRRt7tDsgjua+hBQ5j2dIEW+cEPXD3y1F+wsrTo5LVtC
ujjfgDlnAqPgHAaGkI7UhrG8+8nfh+IZaa8o/3E2OAh2LllJysjqDEgcEFFexLGM
CBGGO3uDdo37PIBFdn6HUFAD0A1UQJbHruP+i2mz/urCf7TeMb9ku9f4o32FeZZe
fD4rH1O95cigCqNnC2twKZsKYuCQ6LbyzNsxS6xibSDUe2lMIDVi3wMk/R7CWgCG
hRnTaTiOqCm9LkSKa844/JF1ZCD4OCrL73u4HClEseG+v8ME1bxg4Bg0VZe1Pjfg
epnoAR9CSghSqKyRoqeKYl09AoNjJcQCqtULgrRvUB6r5fY8pQ5oT68nbWkWXPwu
jYFWoGimYO/fnxe7yLiaCAlwf/2pdmX/OZ9L19OrIG93vUvsIis0QarSKmSZ4BWC
zSyC0nj1VtiDe07TNLCCd9L/NKhXz+Oio1cmiLHjcPj9NpbTynXTXkIA9iPX9CTa
qU9MWUIYltDGHIn5K7Fz/tnm4CXPgzKp2KCd/fAnHzFUpRFfQhhQf6bj8XqGfzaX
bFfO3VTHVnRRFtCMbcLnzLFzhz5+lPIV/g4G4s6n5URPgdtTlRQilqIWuq0Y84p0
rQXsSpjw0l2N3+yxvWhNhwf0mczXh+7eZm4rTQUKc0nhS1gQExcltXgaWL53mZMj
XGpAYyfNj2aN68mm08xGWAzPrvcCFTgdWw/5ApQ+XffsuYIIAYCDu6KrMvOXk5fG
dInosd6CsG1siZ2NXZYNDz2hSOhr5C4ikmAIb3EYUA5IJm1oq8YBFs8vAGvXlL30
LsiPN7xIjqp3EUCU1oksqlvz2oF1a+J/JvqIbzDoZ2pbiIFiP0QsQ79/3CJKQbU5
i+v+uJNYTbO9MUYw3ALoR9ybJSnRbVw/xhJE6R/Oo1gWCHl8urSKCXeN5KpLqCD6
MIZxqn41hC6WIdQBSbDwZOL9aa7ZM9Z/FKHow9XH81fjZpCtsuiEAfdYilwvFzV8
iip6zPZ/X0h04Ru6NR0Qa4A4ghBRoFH1jWAbiHYajOvCqQMgOpIAMh+9yNyHBTrO
2WtyPGDdzJqXaq3W41HQhMwhRCWQWuchPakUzWWcL34WdoiBQb8Ul+c8mrZibxcb
PIEstpEBPTFrx2l/M6iHG+04gojzZ70TGhS6NodBp9/YLn0cORuxIDRanJ/Yz6b1
aTUDKBSdekTzNxkc8f3O43d2T2vhSSsF7xih5aG3VG5h/JDcfJNvx0OvIQTOcMa7
7WZxqxhwRJFJs4fq+GQCgracnSPRDIhv0fQtI2ghCseozHTWr1OGTM5L1t57RXJa
HsqnF3nT+RzDhdemyOi0iOjcMQIzCKs0ILmqnGvRWkdTNxZsUizZZbngBts4vOLx
LcZIAmlKwrydlk+LMYiomMbEakL0UMZMr68WhBr9StSbknxhH1I6/qY1myOL7N+W
0ve7R6o0vInjGNn04rTPjTlzR3BPkv8P597Vs+Ceq1DA2TBIhmV6oO9B/odQoygu
ca61qRUttJzgS1h6lFAlyUe23xT3Is/hY0/8WdDzaSYNIuJ7Vxz4XJWLpANabMN2
e6Ltecr7BWDu4rzwsEWETfy792qeQbhItVfLSNwPx5Er9g2q8fq1uYEd9ZZHVp4G
T5VzdY1MShXP4uKQyWZLIURV/oMGKocjJtG/LhIOBvUq2tB+cYw47ACVZlR2Aq7I
gnBY10f4oovcBuNriOLk/g0RBffQrSttjPRlYZoYM2kIN8VV/DaVmovGI6ZNfKAD
8p9Xavdk6e2lWOWkwse1qE2lxzrFNBq4sZgg0Hxic17Q4VUyZnZM5AsOrI4CCZzc
5KwE7zxcmAG617xzknBfv5XSF9Cq/amw0LZSDdng13ZjftdAemDdazuZe4ajQxI0
ciOladQXDARJERdrdtEyaD0Q4H/YnNsNvryzwenEf1aidyjcIt+G/dnIfhnZtUQk
FTHahQzln2XzSVAkh0rT6Kge3vyUpwOne8W09R3Eg5yziDIvY8+/9Jd16SLhnTHb
mVzpk/ikBZkLKWBNLycuLVxi290y5wplOIX+InX10OvOrIGuM53WSTKisfey0fVf
CbbqZ14bvMbAxH/tZOW0mbqOWl3S8secPWliRE6tsJICpp7qTo9BkJuuZILJhk3b
eSfErJpxUjJg0IdCvrOqoSX6BZ9wfR9YZLYkuPmGI8DqQHQGDu2wsp0avMXUKBHT
iuvBqvaBeb8XL5TwemS7iwZJ4uAycxePzEsiWY/I2T8qVo3FWnMJcJTsWANd7UOo
AHpbPG7VcuqDAxl1oyYss9OpRc4be4z0yoYP/HwrzE8EiYkFlL5t+iqWNnjo7nVA
xZRCAVLdYtzgZpWKaxv+TN3jQj6DnrT/WTsycNH0EyVvlJNPVCleGlBEJ4zFo3oe
/fr9HU93S8RvzCu2v74t6D4ehOoCL6FRPfPH9zEyNyF1o7j8aVzw12OcE+ERX4FU
UotHEOsv/bfnkc9Uso1YO5pVKBaWPxPT2p0dniHXtgz8VetTE4DcSNlFEF1IP25X
4nHCB/1xsLWeaeubGY8nyVET86kMiOYTPieZCWe4oRx5NbzFO6NhaLWXUWYUdDLA
09k9OedWQ33jigg31XPtAvV/mCs4eK/faPtLKVt4nnax9e4Ra5Z9Oe4BS/u2sVfZ
w1B/18UHlMUCXEF2lZZUhxehQMscG9oiOB1K6Dyu7GoCpI9Z1Ynk8pI/bvHPIiaW
uDNl9nLvVqeArhdHJG0DmTepP9ZZ+UiF8I4/JsDvKXpmr4ASLAx5oA45GVkZJmXq
Aj8x941kchfFnH/u5C6qgKlu/S5T2jIxn4oassDbwVYWY4qSQ5IgfvRbeEsHdJyq
shdIn6vE0dELErO8SC5PFi69RihTUxxOS6Lmtq3h09ZJVQxa4cLptvqLjzecYko8
t7rYQbhuQnJrUfD3Bx1sfwWuNEjxlsBa7F2JjH3zWg68I1AmuJ8IVAkbNOFTKBlz
MxQQGPMQF2k1NMcBuW/YTvMErYXEaeGpXY6/garVvApS7TPjNXUqjSS3r1DPTs7l
ifu/viZCdtDWrnl+ix9zG01CHbCE6wkKEYei6DEkt8SiP0kY06WOeJ6Ri9hADx1f
kGCWLZ86EXOD0nQFmzL62gUdU/UiOqrHj21+kHI9qHOYhHdOPj40UW2BCW+SuQPg
MnijNHJWt/Y7XphkjGEStYiGNjgVvOxyHYYzXfL02kj4Ba3DsztFOlbKv87FOuFf
zPoqSiR7YqxxvXNqxszpThfaIs/3ya0YCn/3RCW9h1cPtuxQmMirmn99KxtOM7Bo
J+RA6vxnZtd6Pjzw1YV1mnvMs+hyb8gfTX32GMLFyJzqajIc8JX8uAxAgfNmRkEk
fa/4BSltj6KBxed5ZUSQPElZ/HkJLs2fVGfgFIEoU0HQcWQYIUFhRkY90JNBUS7X
vI3wLobfggJxHzsPEkPhPSxOYIshhnQ9XFoyKH+4riUSH2hsVe9mO43CtZ6bTz7V
//1ADVnW/iJb+OT37N+/8o3Pfo25pWtI0luovpBqGEHeT7qyL/275VXJtFzh7K1R
JW2eTYXNSrce3MymQy6C6QHwu227WGi94erI8Dg1BSsxazvY8Q0jtBVbYKsL9Yf1
3Pv02DqFuic7BH9GjxePKs8eqGPvzLT8pMTh7jSgX2ZbnY3lRk+RGIA9Ufiodc7C
haXmxCzX0Lqsbzw1pGR2qr35bcF8sL00nArMsWFBqbM1s2U7058AnIq5QW7T1wBJ
9EU0Uy7tJHf1SPhC2shy1ssBoCaqFw7YI9F4KpWk2JNXQPHPgQnuNnb7zwmeC52X
g53CHgBC29X6TGx2A6yQ1Ja/T0v56k38TJYV0tsyvJiZilzigwBFmWilrUS6B0kF
INmQV2jtl/wf7xZXhjJwwyS/x2sHiCHyZEuztRwQhf1QsqLdMmnIemlfNTbdullI
YrIaSadMFyUXlmIN2XbPN3MDDnjLX3DHaaLPWEZwy0hyKZ9VjSkTL1VHclbMxowo
QyYuXOsTvMB6DBVL9Lfqg448XmcCWCktLMlARpTBTBOMjA7Ak0GOLZ5yGyElY2C1
Q5OpvQUP3cTiNOrIWVSMkUzhLo9F1ypDL+z+nYbctWkKxx+DARr3iHB7rCKHNBTH
pubClgoaBjR6jb1xviFwlEGMVX1qJ1oAXnzXwxB3neb8W9eYmGpsnQSy5f36h9cc
C1v6qjrANa206wtOFm7Q5vsT461Z+BwnlGpKrFEpxI9SC0toArlYEX8fh1AdgmiR
DgNcZow99UfgeU4g2a6Nv0RYtGaNixF9XpmoxbLf0XrWmuWy4Wt1ub+o5b6wJ41T
5/pxderyY8C+MZNdGDdRXP45kM9+4TjGREp/vUkWwVkenbug5plyxpxGgFF0yhst
+GrHCk90R9DGMtaTVcsbnewzPWdNikzbYUS8/QvluwpUuan0x9xsyqVZ0X3p/gvZ
z3L+TdRPbMlbwNZd4GU2KBLYCEj3bgtm6UitJoP8fAW6MCXvRSlVHs7dz9mMQ93C
28wQBGFAlk5okgaO0hIk0jZTnG3arDOzvRB2Lw4279gDlm3YNUZiD/jus7iqQPxW
aQeNgRJBhiWMhMTHyveUMDeR/86riM/nE/svc98akZZHfmv92+n4miHJyk6g2G+P
8VnEd02BYDc3XaGSgu0L5xoLmm7Qy5qQwmlxfDpM6fjXWe8q/mp9no3lwsYc7gdX
q4cxHK7EodN9nXzQOjjqLl3GeZ0ezs1IaGWuan55XfaxfRvkh+CrcqpjAXnduWXp
pGVpIsqT7ZS9YtwX1NDPshxXhx0TDtWU4suZT1SFatExw9H3Vfhe+brMqKNCoGVa
+5f8O0fUqaRxSTcruReVBOnABXqblbg5j6DKNRcnhT36LX+/53cogJ19lgebMZIt
t89/a9NJMRwG0GVPXtgSLuDL5+CeUbCQro/8bqOqKgePJcMAtOSbMDHCTi/Pw8zT
qN3bK+GFWEEOFfqN9nwSZL3Ve9TtgROLnOZI25zHVTylbeJV7XjNWJKuWULwKu1o
FtE/90DH5evFYcqYvQI9dYDr5yngJSIZFchptT2MA2HEs50fzjevQIwAhRES9ebN
5cX27G8wEc9ptKQNsaW5Y+eysiVPsqtgxayPKSnlUbih3eMKDTsYaYeoG4W0lf0k
RfCxk3HQyWjps/Mg3J4mBirFPelKTll3RvXR3Y6wYzjhDSciZ5k+z2ntQQg49O0V
TSmfN4xev6HLxyGbWBg7Gk6f7E7Ly3AolXljACSAelCNiSJUzvIsKXOQpL3FcU03
8m4LBQG3dObSvj8VTjMjVJe8LGmcMulPu0RSjFK3epmbUdLGr0XAPB5NqxPHsrDj
s+qOA9ZW6lWCh6j/0JPbcJJiuZQGlUmtx3z88a49+KZzDQGbI8ZiS//k13Pr5o+l
5IrA72nJmtTe6nAD+0yFT+cHjWCOaCKmnjW3pFH38ic4BoQOblDzDH1OZPvSKXK9
fcmmhTAnDZdQ64i+ibUTmc5K8hYwcAzcZTW6kjthJO7f901tHsu8wUy0AU777+eK
fkZD3E5UIfnS3VuRejVJbBbq8kUgH3vw91eZd4J+IKYZzeaIX8G3LwpURrbbp0L/
mU7E6EWPx4thW/WQJmUx7N7bSAyz1KNXVqPof0v2+pr5qauw+Xm/oPoi2WjZe96k
hsY2jnvOq2jjTqOZDJj/k1mY+ZJsC6olG3AIcfdJKoTZHjI4Q7pCxYpsE5bg2lUM
DZmppbzmjNwb3HMOmZm14qXbEqpHghmQGrbGGB2RVfzF93bMmuUo9FLo5kcN5jh7
8mM1Jm5EySlCCYKI68+qJihhXr7hgIGEveXvOYH3rSBQ24VppGvb2Vak94/XICRL
BAKs5yumtTvidvonIDRdPSWIx7u3cqIl4V1yNyX5+nFYkuEhhKFHQDKHQ4O8ujpd
Uz4A4II2nxbIRS1x1riN6npxu2PMa9LHRAQ0zvwSnaUtJ7MpfKIDn2tInXEELbZv
ZVM3LdaJEVf6CQfknJ6p12/XXcvlF5sb74zz3scInnmeg7jf9ZZyEue2N0UpPJvt
LKOrHfPBeIfpI1koksd1PBTNc9cwijTTjvQsxmGPu/TcZEfimOBNMaEgyYxf47fJ
zD2bEpmRr7fySZNdBEGmN83lJeGEkjMhDahILcFysGmgORnbWRVJueTNcZNjuE4W
0/R2ejOKbiVTTNoOHQphpiIoDOmAGntpTg/zN60GVWH7IxvRwKzvKXoIVvZr/OBd
jyaeJ6rth7DNBYXIhtcJ9iKZplVFoyPR52UyBNynIqZ2sgun0UiaeYbPArjR6TuY
JLHTx5SU2KFGS1Z3E3lAb3DMdjjWoAxlPagTJgibm5p2odC7CmalFPBXrSqw75vB
M3jJ1DFPMrQguuaWrURoEgsY55JHqIPO701/av+Jfu7fegFKT8pziWYu/liMKAJo
bnPwzvZdM46LVSyr4mWLumc10fMX6/ZH4zutBqWFj/ENpWzBdzaoPgFEX/fUyRqf
qzu6vhGvk1l36/HS+94mJfzRshl1tshqSmllKfO0MvEmMzuuUg4UjpgbQNfGdD+j
6EA2KdSuxBYxoHccC3vtuul9gcNjeUNV+2wMaXXhw6xeVDwmCpHaIdHe08IOCyuG
k+JyYaY3Gv9OlC6rzYrAyJ9wr2FqlVec2LGW3l6BvT9Did/Mpl6BVp8wNkg8c+Se
d44SHy9x2GwRHkGCAB3Zu66Tx4xW5kEvpKe7hZEe00ZItaFY01aCTWp/wrAsB9LH
tDRYA7+1uBxg04l2Z4NW+UmGj5YnmbWkNibxidegp7pUqhepbvKM9E99VtOn+AhR
tHhmcJzKbF8K7yPqw7yDAaCbWxsP9rzrWeKGGpSIEFBPb9aFZY2ZedFBh5pYiKIy
xwT+9sRn1sE2bsdg2BUk88LwyqnTQubBZg2nkfsAaT2P8z4BWV0qqkUUosK/77yO
Oe6iynNMHkr2KKW8z+NZWeydtvZ6/6ec6HisbTSBHG9Em2npcXRo6RefULJCdGb9
8XypSBSD5GpUWnN3enU/Of5lPv3SpFctLo5Bz81oE5wuXSo1xfFHCKobphc0PoPh
WiXQemROXMkSyiD8IiDiXxbdw1sT4Rn3moJseWF5fURYu3a08UiAtspiAnQt1trj
lQ5Vgs3nqpBWXgbgLLhYX5o6bX/OQy4OwhlH4MpagFCAb2xkbQm3q20sJrGwCnfy
9DCHXRgihPATQtIAdzTKw5yN/UE7S+xcJoVbUrVb9n+rgyJUBH6dlq49japbXucE
ooJc3F2fvgGol6U3ouv1+Fgr1Tr/VaM270T3tT10nb6VtYW/9xp7JFQdPi4eCJxX
NWwDqOAM97uhSKKjs/S0fFZakbnbOMICv/k7SMkuoXCKfPHz//ZFwgIqX8zOJt8u
fGxgAzehgRQUkBxlkmqgqf+gfEYN5Fz8BdBbsHHGYiTjQUBzG3DP+KNkCQah8j91
ixlsBJiKeipU8wlcEO/3rSM7qHLsFnkzwcOEtT+Xv6VD1F+7fzAA979ZWkTarGNU
k8vN4sOzoCG1DSeAz2r1d+oWjbOv++JPH7BLQpOzhC8VjIL9TSchbKUgh5WHMYEO
CfzSHxSahid0EEmuUPWu6HifLG3SBZM0yk7y7BtongOMjmu2xlBMWQ25RpbZGTPS
B8OqE9ctZ7jm6NRL/cv8yS8ffunVrvd9flf0hM5hQrulf01SVL2TGuYhAPRYW+0l
c/AxRRgYCaXhFw41E9pLhgTawWIpb82pyNefM9vtTOV4Pk30t7bAxUzM+Trr6fc+
4XAI2XWSbJsYdahudHfagj5E/lsLgbOH3ibpVgL8tASWqWyXF/g3JEr4x38EiGV8
CmFt09RH/mjnjwIqxEYOeE6En6hRkDZ1Di6tc/nbEWzH27tfPZQaubB766p3gto0
QbFAFOd3wvYinSvtDTPA2aT1apspuSFR91r2OskfpKrmoKjz0YHbPdWk8GnF/BSK
wMXamiu7zEJElvatz5e8WL39XxsFGyICjSHInobzIuRgeU5Jr0zeH9/hdNRwKGPK
rHos78WV92milE6M+h+YnUTLxFLtUjQ7Pzq+jFgO5f+KFsyYxnplqWGQLKmA6FiR
7rxzXpEqFGpfYyxqREDdUaFjUEZqHXqWkiFlAN/LZdW6h9aKPzp7bMcb0s48ysJZ
kob1HCtKE1aUWdET6eac64FrqCxAqRyjBC7rY2xnTV4eGWIZeXooyNlWKXxHH+gJ
uOOZgiZ592jygnDigAmCm+RbaFYPwJaHSyv9L/YlTeijj25pp0mwVJoDxUO32aRA
Cr8zr0y8WMEBoE62K1b9H1mAL0O03iLEO5CtrNmfjgN1WI+5j2B9nDQEnF2vPnGV
cR32FsSPmBPuSoibkLTy0gd5IXDIHVbQjdJE0RDIMZFfv3gRYc+EzOwcnJfrVTpr
+B0UvQcBgOlG73pD5H2m2w8Qn5Uh6mL+9v0TQn5Cik1p1QGrtbaaCLGTYqq3T8BX
a26TCREMRKTOHhMtT2uwvToCxDaLHixTXwZmbuEb/M8q6TMF4d7YFZ9UkvvZ/vl6
kEfu0ehjIMPFAa+BRCdQD746AeMZc8GYrYPAn60JnzODpIzdoLQ2fxjT/kcLqZI5
SqpljIG6zULmMn0WvuKFsWhxFb0KEBq0y4I2AmDIC6bnvt1UjmvEyhHYtg9TYIVg
5PdtkoMzQvVn0bfW0l9wFIzFcyU3rfSbEBTFzxanWCPSil2NpU6WwNH443NNQNii
n/HjwjhzOc9oXvaCohe1dknHz75zZNBN1yTVE27lhQcncNOJL4M7l08RqhouUDCj
EoSYfYdkBIx3S4qU3zJRdSRP1Dn0m7DrCmE1fceb9EfpCuMmKXX53K4YI9S+AsQY
+vMbeJXai9CehTmCCcogMf9ZOFJ6Rs19NAsxRAvkXYWXlcpC7RC7efs4FBH8AKt+
8jfrXx+7zRLu6wO3vYNwWxb56m10e6veiZowSqonGGftTJWVhw1EXRtcowLX4MoF
qEYKQj/gYLBGUUIWJGfKKsQBqadkw2hWM/isbdE0NUo/02qYMrmrP63Wbbm2wrPC
LsJmvhWMg5HsTQEy5sqHww9VBe8NHLJoo+GGgLvfeddhqTHSebLYX6ySUyCbu/PE
phYpBvJFPncNY0N1AKH66jaN6bWao3w16nnLsVrKJ1/PV7kDopZck1JIUUrAr4PH
xO23wEC/sB/Jqqc8Ksy+uOwykxEHdJztoYCI4zYX37CSPkzvEbKj+anP1ClKJ5yM
skAie7iV+kXh55AKYM5pPBkTIpv0EjdnCUVR09oOKZpkmA37hNLQqiTf4VfREEtd
dOPo5LUbvDDkD10E4eL4mTSVoEtCj0CvcuPFN9Wgkh302lGb8kopBQFcIYX0DBvA
sEeXJgBkl8/BiiwwhpMwM5UQ6yMpJkmna8ud/0jX9LxY7zUM7ELWT6B5gdpF+hnt
UzrYF2tAgWHW5MU4rj9bRkXCaEMwapenSwzExA7SKqqXrJfxwdjUkyEYTOlAGKF5
xa020zhQFdFfofUu6N0va6dlvXWUk96SMa3skpWRA73qa85sIuIn+ZnkuuGYgKws
ua1USLgnajIRFL1iB0E7XhMqZu7REIgU97RuqWJwFs+Sr0kO6IllDvNaOck6+L7r
ZW5bQove//dPtn0E+z+fiqojwl1V8Eh2Qr+p254KyQR8bBDCfsKKyM15A6tHAgxt
oIXM/2eJplCHCG7tU1KxTHyYYtbdGsS/mtHZx/GjeD+739k4xPTGBTwWw3LCmUho
cedpRY7sQSjpELbr3Rnd/Mkv+vD8piMdpVyTFEeyrbE9hOVfetUEtyzHcu31lL5k
dUYnofHnhsx1GuHnvj9yHAKP/NihWxUAAp0xvFCVleJ+KRgKZsW4ektUqNQYd9Br
yPGQcVbE7FlvcVvCYL1ZIhzoZ0DIHFd4SG6FA4I9RGYmWZPp/S4KxBRutwtG/lWD
Lg/O0ifAridtfGtZt9PiKV7WYRcjuLHK1heqC+ADmUU9fKheMU0tHU1lCcPIU/3r
++IBqsS8kfsm2DSlhQZJF+qsIkjtNuhsiJx0ZXENbXwt/E7Zo9lBgn4t8iprAwgU
ntA/UXyvlvdpil3zj6hoRPxSJ2efLIPV0aFm19RyGkEQ4y+6lWbV5x9IGOiV6GmZ
G0qfzhnOKPs3WYNilvPMXs9EQpG4nYQiuPb+qSgmkEE996kG4faVitwMxoto+mlU
4nZ0n0C7G6CGOxuSoF6pSleaytGgwzNQApUcpL8PbldQJ+cr0aE8GBtulwP+8pnB
J9P/aHm4l0h7HBdVOXVZPbj0fzZ5cC96JEvRiNSD9gx5G6q8zkjF32fufblg9QvM
Z6UoYVulv4npug/Zi3ZD6UKrgLukjvzYkPx5FUCV+gzhw+g28TJW9C95dDNr/tj8
GLEaliI7UpfxRveEIyrSqKVhVBGzRuVfzXQTQ1A1dDBechV1cy4bROXIGiW2Rhx2
3KBysLJpHiJX28VAKr8DOot+BF+Ov/02efgcCmE+jWVeipEaD47Tr5ZV9QYiwE/Y
UyFe8pulD8TQSRb25iG8zM0DmsY2R38GW9IQwRLwef7i61Ii9psdWpNfXPEKGHES
+03GXFh9w6sSbA0MnYVDua0ZIxfVCCWC3+Gchxo2Cn9h6AZ7nFGdYSa6iPeLgAsa
FnaycyFPRkEBXuS8SsP0mw42O71yD/qcnH3THSQj6AZWLHT1UEVyIhQTtLouMGAd
JhD4/w1X+93eXw+AjMgOFboYVNWZ3ayvgmOwOvih3BytXqvj+HILkOoZ5H15+MwU
K+Qyb74lucUOgy6GMzh8YTYrblLmti5qrAfj4Y4AKFNgjvD1tBXdfuoYyILxtxqA
npZjowOBvkmdX72O0mYrH7ccHiDCdJYPor2m5V2FoDpNnkuztwnOPzE1p9Ouc7l8
55/b1MscDKs0fu6ogGzJkqY/9T3ZXwJ0llbqST42c2pHjcFMxsv2FBDE1en4wYOS
wP57zqnr8Y8+QiMJ0DcEZnL/oMzDOYgqB4z+TBWuzif6nmSsGvtH01ifd829bcFM
k9ll2l06/udtomNNT/FVdTMVdWnC/Lw8mL31eiq3uGHIgc2o8yEZ+HsIEOk6qoA6
glPrsLD0wt25N1T3lY0NBdvJBVaYVV5fxS95R54CnmWf23YrfqLalk1rkKJmsVwC
3pxOM/ngcZfO/VidYHFFhrXTrZ9nuLy0WcnLuGk2GQXih2/pz+r+BaZBKt738syL
VtW6C29F6k5M+1rgSHxNYR+G1Aus/E8tUKQ250qoXtPZteIRwEGI0JmNr+8wChI0
zgZVXqXkddB+w0aOm7BWKKBNXZOkBDkvRbCLY8dECIfS2UQwSi3EJJOoHEqE8Ccp
IdC/XD8eV3S3X/S32sGxxPVmh3EDj3PMzWmsWQ2XZnQ+s8Ir57LHHmTysTPqj2ZW
wiTfPA9LygQAXThl4uarIdKBlArUdjWF0FqBRA3hgJPfPESpGop9mrpWW5Cou6rm
Umey7WZ6YFkT9SRrcu/raxsboG/caxzsAxdeJkv/vZMBV7S6IGbjyKCGzEikQhOG
7f0dFMC7AoFzADb0y4ru6gsL5KS5/LBlFT0CfHzPdOZoaenrItA2L1Tb7ntVyMea
P8rRoKdyhDH+XHCByQ42PiW2dQT//gQcP68vF5/Kl09tQyQ47cUsgO9A2XkFiqWP
cXyvrk1OPPVw+wUVYcGwSufbpO5mLGqTndhsnLVV8e+/hgMMW+QO86frHNx1yABg
ud9cd3iSFemD6DDEuCOTemnxxWLkN/gUfY5SGlAOktfO0/sKqx2Qkd3p0Ta798Ge
/B78+r6Rkcm4Zp+tAPg+dw+InUVHIOos5hHxBZOyRg/aZYUhDrRw0IOO4cXJyq9w
MUpLD2IC2vJ/E1a9qcwOH+xeGFQmmp5MJ5oG0SdjJD2Afx3WYIqsVwl2iMQYwNBH
XOsTzpjrcoVR8JKF6vQAbML65aiNqB1GKM43+TNdlCNfpkD7g3mTXGYJ1WterG/W
Nwui3tH4dIhzM0D0ZIyV2z11mxtCnIeQ152ujm0oLUarkYPqdCDU0kpK2jXC4hwp
ed5eAX+u9jPofQXrBPjFhvUHmde8JKtjeJuXAkjQqF5QnU6k0oJIaKnuaYtBSFOI
qb9Nb5QS0HKcWk8RzcrKU85WyTaOHBqg6Z8k4QLc3D265wXtvtvfrBIB97qHDn/Z
JF3hQeR2uupTCekfcd1f7iT+u+p3ZdjPDGikSTMKdboJrK3NB+20kv7NrBglTLAc
76UQ7tPDJYTwBWQPMRsdwamWJSpeoVTYFw+hMkVc/VuCEE8MPYqrvsCReqY5GkI7
pdQyeGjqm/TjdEoVQz96G6oioZodzzAqIWfvTMJQg/UMCV2aM4/T0WrLt2U7+irF
zyyu7iThdfdZRSrCB+v2Eor70cMQXBLbxJo5HtedNfkO19jSg3VNKfNPKx8iH94Z
gczo3aPY2KTL/mQM1aQqdlW8YG5g7sywPnQ1lhISTHnwdeCkBNG7fMU5qj/YkOj/
Bc7pNsgm9E+8gCcwWhDm0kUuhW3a5s5goqCijkRMRHiJhfmrh+IJYBX6f4R8XCuX
4DnPd+49cQz8v6fE7tR6MsA+nulXZ+WevW1GuNUVvSAoIzVPDjP+iMeoTHxECtxf
RZguQ4DvjsPcQOSDXkpKmDsjYrho4hs00EtW/E+e+fKtocDq/dezqttu6Oqw/LG9
YbAb4qY3uTt0Fa7VXN65ydQYJDU8+a5T6yrqEjg9SFn/FD4/fn8+npS+kM8NuDQC
P3dKQVK+Vgu+C52NOytfYYxXwKK7MTyPU8gjjaVqj9YC/ptYmyEwO5oj6WmuVBr/
zcpGJYS4h720LibiGKAwXu2K4kz8/oUQqBP4G7mWGc5jFUsGtU/1VvhdoPovjjSW
0frzYcGbDM0W8CWkrD0DUOChiSt7q1dM5c3+Bkm+sRFlZqjALdYfF7W89ikhZocr
87jmNNTLtCfy7fYXZFtQJMDnFS/uvQwADk68lBtwkucBDSfq8gvgUw2hG6TfIx6J
CzC6zGbVvfjNFi0VKUl8aPmStzCpMMZ/DUlQZDyfvyjLIt8uTFpl+ki9mqd+pwqs
874g6JOAjmq9N/PIylzC5W397Fc7sWPb07T1mdedGkeCRAX1iKc4LtdIJnA25U29
i7rJmXDhXQJdP/7sIgdvIyWsboeMdEBMqpgWVAWkq+xJndiwslABW1fSVfB+tjbo
MSIB/n8vcSmnP+Dl3Ti/hRnPIu7SwM0TVQts+0gLM4ew/U77nt7VdlvQD4+RWgbh
VTVZr/32wE6koBbM2KOGotIav5Wz+eweB/TD2irsdfwwf4g4LRr7U7cll/rzZMBL
PZZY015e7RvuaIX2XzeFLKcaXloc7ZwdRh3M2N021aiJfYWc+dbuUYrun6JdoPfE
Dg8ZScQOhBjoUA+0Zi7sya42vXlRx6ferAdDLBJEq3W8vbLOUvSSZpwopPDJyWEO
u4E1V28eU83JIrfaURpgueg5lvxJDh9L4FG59V+E1Nn3Kr9o8Y0rAvUt9y3KzRaP
Rf2VM5CIla8/SB2/BeZdnazCgQYNpE0ia+kHNOulmfXk5O4wzOm9EojzUYFlW4hV
yv6gYoN4v8HFumzXFJm+9wOBFTgcH7+CO7M7UcaeL1/iJwoFDk+dU+RYfdLegEO2
O8PefhZA/BDKLWlT5K6NZDzcS6PqeJ5NmdMKNJTDnELAEnETx1eO32G1j5v/Kc6Y
tH5IFO4omlerpr1VmbhxgDLBDwtab61bNlny5Djn6VWYKpaGc6DyNE1ZnI5cec7Q
8l36k1QuNac30AfLgctl5aR6rpmQs0Mj5tPW+6+FTMKa9d4z8eMRXTKckS+I4ENv
WqIPA5nMzaBesdMXm7GZIBkw5JDvMpoJjYzWHL0WwLxzaZIC+CDczKm72ViQqQ4e
1PYmUzwpMIHhWuztHvFg6FQ+NftYDmjDcg8J515qK89fHWrNtSpmthd3RFMwjMGP
YdsraHaEnHsN7z0IGEZ84/rOTMAQf59/OhoyCHloTFZDv33ea4sx2G7nx3Co1Ulv
NwYw68dVIStTytLomm8qqpwgs5U3uWnlkvENev2FzZ3ClBxZfEIydopSKNFFrW7B
8tSc01B1gkBABBC0Irvh8JnMmsvIKJNfjIicuVz5aE2iU02R5k7gIOEyNasxAu+R
nwnciXNaWRJ7M7jHwfXyHDqFRtS3ct6/dIsJ1bk5HaCJyxHjRa7+ZugBTovQeEfP
eX+VSdaB492InBgH/9pyyJFlwGTej1HWF49dbpElGGJQ6Hq/C32u6aZNVlkKdluD
ajkY/y6G4q2DmzwgXfozpnAToBGTtjyMVr3hT1caUqj+VwxN6g7LQuUBwYXQmAnO
41s4XxsixJuPfz3xadZIWiLMCQ90VdHGmukcHYTEpTrLXmu76Xk0CSkd8MfZuc0I
w+8lECIUfG6yU8y2ep8mbA5pU9lMifFMRjgJTItSPiWALmyfcSv+Q2GUwqSv1Upl
ifgMVXXkiwSRXN1OghY+rEdjxgX9XdpY8b7Y1UkoF66vX5QjerOFo6fHwq+fib0I
O0jHpxkpm00rqqMzOA7Wy+tXRUy+VbCTc1qPAEL95ZpZEbSkCx5YK3nSUvckixBq
PbuK1pjEr8iyX1Q0RdzsvzmB9+rOwZvh6a7NarWdz1ZijVrNaSgCsRQAGQ9l1fyK
APyFQJnTkY3U3jqaMlF+TjwcVS2kfxGYFuAoqxdZjxlgxQl7WJZOdT7Lki+Bvv6X
bH6gh0qep/VyXRMcPcKU+JhCmpDnfJNTf6IpbYwdx2WSscg3zFhwTvD7jnOBINFP
uPCMOaCPCIJKzRJVqGzq36FBNFlaQNY21tjERXDo0kLGoFp9Eq3uTxUBBmhwoGjb
awV0kVWRzBE1mIFdCvNsmOMMHiiz4PVhANeZgGEoLU21P9aHQ7lFDoupSEovEU/J
XHBKhXYxnacQNNkoWxMXwVBLoP3bfvLkRWUHx09Ycs+Ka7iIAvMtyCDPYHGiFSKA
k/uG7kOV1CFuL8GzP20DEGkDzRFcn+Oww+Gl/DPRQfV/aUv3EkEcxPGaQKjwOMNb
jGKS2JEqYL39MI11716j+Y843tzYlxrAX1uHei9syViRhDV/G78qJ+FQbu1ReFtW
B+JQj1U+/8HN43tuTtDYPp3vkI+zCLwlhKCB5GuZWmtDinFSvHnKT7Jkza6LLXAI
p3u1nZTeAKnASU1/jkPugwF9Dzn8KsmNN1+KCebscIcVE+RE4OZn6sTkpdFEifgr
imb4oXA4gL6a4pP2kGCvK553pQcIUaJqe8r5UasoScabsrW2vhOA0zauLqI96ZkZ
fAOY5RQzJ/A0gWeeKw2iqMNFppSdHj5ZluLyPyFfq/irZoTUCtIaMsreTyqcsap8
gdBfRGajluAhZ1JDXh7LD4W9IE3Hm8ZSCsI0mAF79tFjrxj7abLz7y/Psselt1Rh
dnIOIOx10dg8EVMVmnSqH19GqhAsTmQys4HWBmvJzsiHrz5vOTrfbK4yeoMehn6u
cXVGbi/VMCPjwvBP7kmfLCL7mHhsFRcrhgij1/PWYNZMR/9evKNjy00aSwITub7Y
YkIO3z8u+VoDcQn0MpNCyzYZYNNe79J+89kT32VsFvzD7wQFPJveVRiuksdx8KxM
PkuZC52jEWd8T3LIM/mkLuqWM7WUD6SOznLYK0Hk7hqSG4WTv99dYy/sq81SB+MQ
ABWGXBZPdTVhdF62GX6MNh53MyuiSQXmHDllc5cvP1uJZfjvVqW3CAX+UwJYA9+T
fuqrZb5Zrxej9+JiDyINyqQUPBAiC0nOZ+qmHx5lKxPm4/HPxFQpVardZ5faWJlL
4T1JRraRDJ3Y1Lep1TEE/s7YrAs6CS9Z88uaBxbNyyU/20thITR3xKFsXTgdMmQy
qcPYrJXBGN3JtyUBL9YNGCV52Hi2ey/yv03iAoVJwn2udq+5MJ5q2G7J42Omegs1
UzJMYBVTbi0wuNddXb+VFu3ShkOKd4lwSAGv0eEt7pzIO7SHIh4++YSCgTtXFE1A
xWNHKE+R22hN1GOx7CrPyNFcqrOe36seeUSLsCsAJZeTAedFw7OCQHIE8asriInC
W7XB3FXeDwsTZz2eha3CysxPY1bPXZY/BNOJWzcdU5tcP0sogq0gFOSEZE3Cpqn9
JAXBh4rQWgHscZ2y1+V+jifYvGRwu5JolSG9Jh46VCty5yrFNCrDGGjkg5E+YmFb
E+GtyY8u2nCtZfThdYFV5Fa795mqlUT0a5e7Ko3i0GzhX8+RzBoiwJPyVvzZBp36
HOlSKzVktb5WWl2Hm8+WkEfwMWZSrkH/XdDavfFzIw7SzgygvhTfdlncENjFOfYb
vcCdkWlHl8deAdSovlPKHh8fAK9Y2qoveQBmszCafLnv7yZGRGrejv6ZOjMMRS2S
ONuXhhr3WoNxMOJYmGEKwA4HdiA/+7/YuLD3DVjaODF9kYLdnGw/xIKH5eNKJYGu
MexU1wC267SfVGoZcRVJkdHSCSSWAI5MMKzxccWhrNIUYjjLFrzbrr24S9ivx7SR
9G3GO6lDGWoGKj6IBNgBxjfgztT7tKbdPWzz8eu1qFc9DupMf2M1Tcz8yE7mg/Qr
vOxgqRiG8tAvzcJyCs0t7MegFeVDrHVT3sY7L4J0aJkUGjGm1j7VmCiWxBKwyon9
GPxgKWVgPpxVV3ao2Vgj7BcijroU1yiz+0LYtuI6AwfLOvMfZ6w2NbMME2mVa14+
a6/QeHn+wq2XosJsZ+cV0zEkdun0lspKHVOWGYqwAuylDNsYhBNJb9hfHZTJ/eZQ
fpi1e9E8SN1rTY9FQH0RArLeSDyB4v9VVxa852JfkaJSvdEtUUoRYvix0KodfSg/
U55mphguTL2r76Zj04s4a7ZHiTY71vZmGiijJcBnQS77hzI1f+I/45nqqt0dhMAv
ChifTr6xIyNwgRRIkx59yBzEmRadFB3VXotmkYk7KhRaqC0fsqutndDwrWIo42LP
HmqJxtAQOtkZRZ2YtVPHxrOVu0KeJReayQU+xeh+0aw7GpfOzCf8VWZ3xfy4ScJw
5T2HT0E2mpa9v1uUGRs1ZnN0IHIJv6OmP877Z/xEAyCik/+zYEqHavTwz00r4I/1
MUynkNMdiwJeil38v2midg8OxLkUppS2ONNIntl2plS4k6W6nE6rEoKo4ZizGhqa
J7maljkm1kT7eMz2Yhq8P4qd/gMoQomFqNXKJXFP23ILZEDizI9lZUO3t+HP42kn
6AXyCBz8/8qbvG7I5ro+CPnYjKWKiTmbYdQl93ODmPISow+JPi7VY/B29IlyfIhe
Ilh5q76SwKzxE/PKRIB/nip1ZBm4IkxCyg9DAmYsiKJleyvFVPimKaOpDiR7wZhX
m3geJgJTxVPXqW2kfPAajFRZYDGTdfW3B2a1+KkMFGipswJYRwE1k/Q7Ciz2cGi6
fcQZN4cvtI7QhS/+KmIX9nMxzgdh2H8KRrSPmSJI+FhXolaLKewarZW2+cO5SO1s
nXS8f0d8JG7v7Hi9EDWPXfYxx+qcl/0JuAtf/fhzCnRAnXEHYQn0VYpUH//2Ipvx
cfz0F6ShHuhE4GdPUNDRnEcgn8l1+Wre0iGYnKlvhdBOoxRBhzj1joHhN652JWTa
Z8usr8kvQiv416zIreFYmWFZ19/SJLzR6WY61AJ5N3E3FripBx3QwfVCqXGLKzQs
t6AlRKWWZB5ofG2Sn29ST8GGNCdxto+4dfeVUZHWPymTUTLuU3AWXDt8GTBFeeea
d7/eSMwNObEvp8UdbntxHysFll/IRpHaxbaXX3DVTNe1+GBfLqf6J/IZihG+b2Hu
bbOm/HwRjZZBKcbylrkowgpKJJoPika8f2JHCrFFStiErk7VqtxrRhhsvW2sZPRi
at5gn/PzP8+G1bPmmHKl3Ky/WFRcKc/xQy+JGGUer4aLBPDV92Uyja1QsbS482P7
trBwxGQgdbdD9umrCQzlc/1rFpixVh1Czacrx8duzLI8xL3Seki5HjW/NUOTRS52
CL+/NbMNjHL2JpFuqqYqXeTHrC0+LwDWy6CExonwpu1FYZ8n/k+LwzJM700CsX3Q
hAFEgsrJ9LqRENwLRPtiTIowf3xEirkzXjUKtDrZcoUGFgJkvONwRS68e7H9OOqX
5dbXGkYLTDnHtRwP8ouzmMtM/0HbEblVAPBxsJkHME5nPMQOwct334H7L2fokVEB
MAZUDhb7IBEmowEeFTEOXreOcf/HNWs/fcsE08M2gOJ66RcpJ42kVO1ko6oiDqgf
m+uh5TF8bJVu0pzilyuCF7Pn5pLNreLpH1XRF1ATd0Bq2SuP3lphuzzNzFHO5ML/
Cy9mFxyac7BgmhuCehOf4TOVCrL/VidpRqtt/VpsYlFm179UseyLsxRdp15ZF6US
wrDNzp1gjd0dXPfRI/lXDDHHDojdlGT+JEo++hAHiV0Xz1j2+h3YvU/2CvJ/yL+B
lP679RN7g3/owHifxCsVjF6OHI478m6e7P5ferRPszOHuLPTFR7bg+1n5QfNW5US
ELdRSFpuLaNgyuNqok8WhFndQgcxq8+L8STTGoRo5uITMoDGIu03wqEQ4lOl7r9v
hxfDyFFgXBX/9F2yvcLd6u+3bDdMERz3a/lbHq5gamK0uu+ZpNB/6k9kPY57skpK
nDbMP/IY9/4UHOpt4fg61UtYznh7DbRbZ9BiH7utaC8u/IXLsf3Yzau5bxkNYWku
oTrJp0xYk2tzbrs/80LFIKDUOnY3trli3iJfOTM6xhcyr9wVt4g9+/F7VuPW0wV0
LYdQwb467yXmzQ76Vdb95wEbM1T/tEj2quJHnm2MIU36oGrKGzeyBESnvujTlwXq
acDEwgu6MOvt+JxnaC16Oy7SziffpAVl7X7MASCaG9CqEzkEow1d+3YkRUlQAD0J
F11Xx05AhkCirteFp+JLKmHuXzOqoLfuwPT4m537wuI79Y/Ar2WE+CB+6IMepAbc
mf7OfTsaZX6NitQPlGr3bHVmSl6C1BS6HkT35/2OrlroT9AsdW66Ix7IqGKoauip
CyGWdmV5v/FccT0jwg+6jXbr3jLZt8dtde8uEff07T3+Oi1OpKsEFPhVG9Rkot8n
14XFieqpr1O3bggwu0X+OI+mrzW9OgcFmcUNw/LFqsRIs+WzOdKhHk1d55fnlUTH
7h+XPUT+bDiRohAuaa40aYlv8ZF+SRzXV+gd66EskewKgoR804D/c5/Wrg4+sVnL
4HkTaJkx3+oe3eLFFDWrdCXEtTq7zo+bf0SilfkW1B5HQr8PTUE79C/1rf8NdZwc
LJhVWzYp0DyFWGgm5mD/ArC/sjzFYgMnZAUHuNRM3wy3R+PcuVkF7DqKGthGd/Fc
o8ASW6f1ruPQttltXwVGA4oLVqpGlZoATXcYadNXnjFy/NEjGSM4MRjJHpKL0SOe
NgmL63UlTD1C1qYq9UNAADSu6HcCW48EIKTsL9JWfNnV5I6Rnd3DrlojkTRHP5fh
oHPjn/+y5x5T4AGOznsCLPh/AnT5jpVXQSirRZ0dTkzQ/YzwFKIghgLw+3z2Df/I
PTcUngmSi3K8cVE1wTASFj6ULwxjaxZQUxgW/irE5/7r+QhTLvvJhxWWaXnQxWZY
MNlmMi52jHSuPHHz2ey0drbuFjwC/S6meO3B7vlbwO7TIGzgsmvblY3IuTqOECZ4
xRYjfl6NFS3YHYCr7yImssLiksM4WXyq0EZ1sFqB5Rsf7/g7kW/5jHbqdQmcVPpR
IhuCUBPFJ4dO4v4JVIO1jvAKe/mmqlevuKQz9LDi38w8IoK6D6Nlvu461KsRPTvJ
d5VIuChGfh38BHa8lMzphHz0R3v11XZorfEK2R/QLDME/1ZUty8waUeVzXH5HBLH
ula1S3EnBW95i0WTc7pGcnMPAfnziZ3KUy7FSlDS5+jUxJfXxdJ+6ND9l8CrOjaG
6F9GL/CKbhBVB1YfuYbvG/zwQWeNB4HERo7g/ZBMXoCJOh9xjEdHsVsJB8UKebaM
7MoqFmECNHrKHYSoSIC2Y+D/TVprXIkrfP2BiNHRcvOKxQjPAXCia47gK7IK3loW
zVZz+rbMzilthjbd4QjyfvJGXuCC/J8GEr1XPBpr8JFjtzV//F0RaiFBB2Ovm1gZ
Qa9BrCHENTQ2cKJJg5pJgJPx4/ea4J4oSFNaLBHkoeYCr7aKi7/Vj0/tmwhTyDsj
VVpcuby7I/J79hEIuxz/6b8NJS2uL4EG+fn3ebdUPDQGBxJ6RizNjAPgGE9St/Rm
kXLyb/TTLhZmZhOr3GOFlIIv6BvddeEoBAb2n83tPJcqXMxgVbeJnv8PNiPTmdtQ
DFDuf5gcpcSAFjtBLIcYWtX9s4RWa/zOctaeEMNAvGzwjkoJ6aubbTFyeI6hNQ/J
5LrJ5EzQ+ta/EcWYCKaS1CVU43XmSzsSBH2DxywPlcmkec3SHJjDtPRJjZNrMU3O
l8TXaReAXv/1Iu8XzjenkrtIp4P5eiC3EoKm07o9fCmwkJiCuQ/27PVREWxHZfll
81XYw4Q/PAi37YjXiLptV4sbHGPQXFw74TRtVnxUcrrNzCBj+PKGxfd4859PtuPN
zcS8QNUMAcVMxGTnKySjZ6tvpG4pG/eHw4SHhgnomRZleDmMK9MtqEpUufASTyPR
GKks8KW1BqQ9wtKROZFsIqL5XJX3yNHRYzJ8tsJvstJQ0y1SRIGgrscQvy0fKDNS
C5YtQxz0q+Pvn3uNi61rfOtAPk2pDZt6O3MUAT8jsa9ryKocpQGOdqrWq9jtBjSX
BNcHbhoVpROn+OjjtEnbs889jc39i5wZh8DpdhB3T9FUWZh2nbCLtqE4Cz6sCyFh
7g/eCSejPMmPu47wFHiGYTIxUQtqw4/HFYSeI7ojWocAcQF7nmF1wogN0hmffABi
pEuLZi785DgaipHFE6tjfvg+De2ex0vX5JfYmB//U+40bdPvCUVuTKldh8mx/Uo/
YzfPE3mkvV58RctpHeqZjSbMQeoi0Uo85ITG5ZJoK+sPABFe6YIL6Z144RYfz+MR
4PHbjkAwx99RD6GxF/Ve0rYCWkkp3+SFo+QlDNS3kkvenMPizwqMatiFNJXBnBSV
LvBnDSlUyhqszFkzYG97nliEl/hUsY/eFyBFv55iVs/nMb/wCJ/HBW+A8BIEzb8a
CBZ1MYePW4SCyqFmrVV/EewJ0m5ZB2lGxtVk322hU4zFJcmrabD7zGg3lsxKRz/w
/cbvRxWSuEw/PUcYl3Hi+9lVP2QpTiU/cfCANC/CGS61GCDRCQPL0HyfhCdQFwNU
uNggCw4YdGd0gqaIeSGTuAixxraMcGi1IdXQFYF8IvPQd/y1WA3DqFT1+t2cYH/0
EXIRtjNICoaMlpf9fK4quRuozSY3uqV+VUiCNQXaCJm3k0M+/21THcoj3Rs4biTO
ZyaMAF5sF2TU4pxG//nOhOMcp+RFTPVs6bspVNjEjtEi8EEBuVXkPi0UGn3xiVM8
0uOfN+BEc3DkXuT5TGX77wfk4JCO0LYDDA0HqJ/IX3Pem4r+1+EV19KYgn5fpVqf
8Cdu93j0J9wWLItIyDN/4F0A4nufkPgTbnLgeKKscZWXmPOsh8W6px6gh0B17Wza
D0mB/AHjO7FJJwJ9OYDGMSRsq/lzk2QzXTaxUbNPTuq0YfmvE4+UCJdzV/z9T1Fp
n0HhV+J3ZuZAnvy65GZulWpAjmpf7QyucxFG72KKp0pu67ZToXddyw2xD4x5rSAp
FaQ5JBuEdoP31fCDAsU/PROB5T7PWq9pjJQXTUkTEjs681VWLyMpI6VLRsfLDUpQ
PjpokT7D57Bnq78UIWFlaTTO87p8zKPKb53f/Ke2zE5JH/7VSnY2ynHUYAICB4dA
vx5eZOy3SiWryFKVNA+SUISp577TOx+6yOfn43lJOsQgYZBBCaibfH0bfsrzfB6H
y5A0m8rhd/kzsSmNO7OVe4dDScQsLDsNhqsdF0A6LA8nfS6BSGQi2fX9mA0cEhE+
EklciOS77do1ONoWiOlDg+E8JqXDpoyyooA7LORRrNlV6JxuckOAzB29/Vdk2oWe
Brqsbmik1kAGRkVj7wua6VZ/pxAgcFcYFE8y9aKl+8cYE7p4LlN3FwVqagZBG4vG
Xt9BvkqaA4IxB+SoGJQSJf1frGr1w5++rMa7p3r19f7X3TYX/GdJtSqeacDLgYB5
rlzdoScSn+toDGQwMel9Bdq0fmLXunAXS0v7AzBagJccaRQ6UNXsJiMnvVF/3bvr
6l6QPj86Swt3/5oUHTuitek6p/SbIJaDd1z7xtASU7d4sie8dKXB7aCATNiQBUCz
s5WMFJPk3EoFrrbjrgiUYQPGIfop0v+M3SRxNrJtWSd3A6rORSmhvo4kQbk/SfI9
TxpIWVTP9ZYh7xnIvn20rP2RQgoOJXmHg0HRUclaCb6iYos26w01sbDmZWYIEY5I
KM15bzuSMVKfS9J8jM3wB7alQxMh7TrZEMvvfp3fF9tZCC7Bl5X4Ae0faO6Qw9GX
X3j2fcYXK2f+BbROr+mH7J7SOv6vB79Z3luvlNXMkBvSdvrdvce7TTfnBgkAyw2L
bCRhoKoFGCL751jfLSCnJ3ufZ34E6SgLWRTccKdm3vf1yF8Bn2O2G8bEx66g1eDK
gK3K+AwHCUmurjnq6wbniHqY5wZal8Eqf6j0KKtIMvW/cUl9dy6nz2YLOgm16JkB
Qn03Td/5yxw+HAtmf76QBlk7t1jDPUjx7qi1O4AswnNFwdyYZtx38nvj7HD0B/LC
kUTqtjFv6bSPe1wWYNC/OcW8yXfS3c19QBLJqLgAUZ6va5wVwdrSXxw2Tzr1AUuP
heRd2aUAYU+hto2yNQu7Q5xIH4ZSplrwqvpDdfffNqmKRZ8Xq6nUG7zgDiinEh7a
/TPO0SS3MgzUm02sRVt2KZSmd2kwzzdZWJkGSQz2L9wiLIemj/Nh1/8j00Ff+DAl
6TnRwppCodT5e6EH5PvRMnaw7OWKJklNa5MI45Pt+bhTj/r1i81ilcsYREr9vP/Z
bMpk1RoVgprTOqewnrWemNx+LolHUy72EQL6u3alIx+Kred81bMipOKK8OfxDu2v
m4uPaBZVedhf7kLJ1KStdtX9SpnQwcVJYfWCu2zj3SUp8QPbW7qgUcLaXheE/ioH
y+cDPS27tWU6WDa1ho0rgUTe1Ac4NyURZHW6ocE3c3Ix2nsocKlUncYvt7sSwM+5
VeUmlqcBLP5GrXYt/NsUOz5g+ZjgB8f6//E9jlfFNoNtptLmMNGA2myeM8e6b/Pb
IKEGqR4evNMkum2nh6iNDKOWY8mW/lZkTJkSa6DmrqkiXox9c4KdD0KhQt3RbzfX
Jb+4MwBnR+J/UFKvzX7vrV2m4l4HyF8TNxNaqFNdtAEiJlN5jO4q6aHwwbiCfHFN
ivbMTKG/IAVgfklCsIpe0mCW10uh6vP5v2BAc7nfBFSPJHFmYPoaApBKTeY5umJo
jEhqa/vcX26o22NIXkj74CnnKOz+dEAahC+qHyPLbFpm2meDLF6vrS3FoJtCHg7f
Mg+qY82TnsBNEcvPhwNaphWinaMnb1okZURkwAF0zaAcKQxkgJnYut8t4TLtB+ur
BWFv2JxT2B0aTNOKnh7I5gnsB/SwcaLBdUoorj/8cVnE1W8f8RlzpDouX8feVu2x
fDy+7OiChTY0IW10mVVbcjpCDb2xjiW0NR4C585TbK2IPnPdo8VOTvUU748wDOCA
4h9ktzWLhc2ipAwHgPSRiNADQ+ygxrqNDkbSU6c7BtkGn7RML424tV9Y5eQRgz8q
ooXqIabKV4giwMhSqNpnUTvizACpCTiXbLUJK64lilyajSx9Wx/7mQz+v2yLuEiU
lJ/PoLJ+eRiSzqVpMnSspMSdYz0EtX7VcjvPDiLQe5t4JB2dV+uccKLU4so1DpBe
u5NuXpn7YrKakNOnv0mJIowrdQ8bFe//fpgERtt5zr9VGlbEJvnSUYMMdSwgKqfL
pSWli4L58Z8UCe/KsT4SIMSDxM1YmTtz43sdjCAWeCtli8ekSO37K7K3ho8BrKVx
fGkyjFGsdyPvBIlOvJggD1Q5A9Dw7mQ0UkzJ/148Smbh1U5kajfWmFqto+e0yIwQ
PIZwv5tTp+gQhxt7zJGUUnsNJenPuoVu4XrJ9ARze2tW+ht0aeww6SL5WnMqPv+O
kaC2794SCmjVia+KxjFUdrXm2JbFM7nNmQqt3YEdxvLOnRFoHP2+DhMPQa4CjMEp
UvTXm+IpBZcLe6spOtVw9yhUDTEQnk1Ku1+KLRMVbEkckGMdeEHni9boteTWc+OV
9bL5IVOyohimwBckRVFN77u472+wa3ckgZXCjhBDee/x6doZNIcfaUKE6tMiPsXT
wPkuUaM3sNwnYQPhhZPF17UCEHb4O/fawPIfnhkBSKx8Etr7nZtXOZN7bgxkcgwa
rgoHhuFfqDJWqIByM5ilrmHLGstLfxvzLpMp5FmL1QVivicFu3Ozl0zd0lxmHMyt
19WlhYti7DKT6SAKuoD7PmJmYa2lBYuNvr0t7yhN+T/4AyM9p7DjrsnVKMaShi5j
TJ4ZfiSAcDVgWnD5yrPVqYP87AeNDFf4OcJdCo2371V2t87qYwBQnIOdl9e64F7Y
OC+IpgM5Q2anFKQJHBI39W9zm8LkP1B713GhgPNeBKi/pvd9AE1PHDfjVrkht2cq
Zhwo1bAUkgYuwWMAr9TJuRAkYZBRzGNya9UKgpKizy4P0O/bkPNdpwIhItXYcG1D
lWmgRGjtS9ye+xasBG5rory0HPiFX1IXgkG2nuXYSTXQx8KK6YIIwGsRuS4T1Wa8
NO2oUhLhRQw3youtXvrqjsgjLUVrgnTYP5UQw4g0IPpuUdI07fsEG8EzkjE7Wqno
0WhIxTsH1lOtLw+Cp3iBfyYGVJc+UwNT2DXxZT1GceSz8eGuFNjn4fn1h13iQNJx
2j1z6m0LIPF8ERfbkkJsRUAs5r+wT+hEELfaet6eEEb6x7CgG5AYqw2zyY97kRL+
Y2KF8UdFl3kaLoPyL9v+slaCzzvB31jv+nYS+hMi4R4zMvO87TWHCGSgeFhJ0jUd
4IuEJDsvLT6VNlZplySBggJFk/RolLqf4GSbjo0Zj9TfBkzJSn7mWxw0UpUFfvbY
tuDS4lc9AGfiIJd+ghmRpMUz3mQgkDOtRWKrcqsosRJ0ASeGD9brT3uz+nZ4pSA0
njVA10qBkh8hVooTigX5ucjYwY+qFYYgQMAIU66xPPfvyrwQoYbMOg3VfVj2DW7p
+BYcW6lyLAYO7VuLtEbEihpgV0tC8Tm9DD+nnNg76WjRpTTpjLHCXdgLeLo0Rzbq
ZXOFbTO+PJV6+TLnhXn8BZwtPATXk+ijk8Z5Z6Jv4Q84Ypcu0fxVYR32ewFAu+7Q
yJuSQTGmdzolawu4HQCEEYtGRm2xKYbMZ/Ka7htL+UiX50prYG5t0L2QXdHjMSbL
/1mGjD7ryQu9C4xs5eKztJXI+9DkBUe51INbHAjI7/ch0EWDR+WI/UaldXXs/y4F
SxMPd9OPXFY/fxRK8dGbZBl+e/UbzDTAoIIB/zv4ph+gbNPt8Q29Pkvv9hkqKTBx
vfzoXLKGyyXeQSSEptEZ8ECOvBWYrRcjP8H2w5pAYXnKHsTti3tDfs68G5I5/8oN
DMyk9RPoRdFWuBRsCgVJp6297d7yjnB9CbSvt31lDhw3tkFHQ+IZuciW8aJ41Fsf
nxfPtKhy2W1n72gay25t87lbm2DNQzSKB+ctNuTFmo6x0XrVA6VzT8EfRnF1U0WE
ek8JUl//WxsPsUKxQA23bJ9YXVGFuiwuwVuIxpdH5n1w+O9bfbsAU8QQw1jvkyE6
y1iBjnADlyDWk0bHkS5rtNpuwfrTRWN4bq+e3h63ZUXA1CH3jyFoC9eLXhpc7R0K
7ifu36IhOI3/9Rcexa3p7aSUFGSEuehKTIIGlbsW1jhB8fErIEZLjB2JxG/KrIWC
lfQS2jh4nZtPljJzOnQoZ04A2NzXUksxKmOZkqV3an1zurIiij3p71gxIP6d/9sm
Jl7ufO3OTKDFHewuV0Vj/rPQETE8/DBufL6qVYRtjNaiyiGkhUWt1egUXQi8PSov
dW1VrUQ83SQGs8z0Y4hXLU14+NHcUbsCy64bIGoHx+/1ktUIdafsl0sLUwpCrusL
FWjPpDacZsZ++Ywq5UK0NQooUOBFmlbtjInIDVMHZFLIrJUFuVFLbNzOC6Rdga6l
s88602DbyUbrCfaz6FPIVuxzg2/dGqh6Om2UNsSuKND9rKvtXhaqXTpgrgA40nl3
tgTPEbGKwqlb/rmBwDbB7I5wpD3+4JxeOM6hVQ+bDegq5IEVyjP1WdlLnV1CSLpJ
98OYHjm0t5K4RhuThjNYwoeCXkEo1SC6HQMwZ2SITz7l7aS4Xft5e/haf/gecb4J
r5tnWDwaFELAe4Yf2w4foiyofyOCzugVkBFJ8eZmGHwSHDI+FGkIYsXj5XUTLdqs
Zoi9R65iPpt86Q7TPrtv5szjAv3k2i6r7k5fSP4kRIvIHd/syAoZi12KLLRn/VgD
8ah5Z8GScEpda0UcfeIIVsdioUzHZFLtHTbgMajug2uXsj5zvF5q+DSgI0JJxp0Z
lRniaaLsK05PHQmytKZlnbKp0m+hRA3AmDC1waXTFEnjisxOmb5P/XnWpnxxqbNx
izraGGNLez+DzAkGO4Q5njq+u/xtak+ld8xPuTm4xvhVVjr+C9szog30K6jKHmKV
ZMGZT2eexV7o7o5qzEsxJPSvqfe+MKYuMt7qFr7UbMaCL3cu86FV7JGzRI0dBnmY
4sRFAC3bPoXqdf0V/0UBViUn/KkUOQGqrNxhxRxUrUUwylfxdFOXT79FBGrVJt83
VfTJhS0eBu57u5suQf9iMDdD82IQwDzv92KT2Ytzj4emiH9oOlwnLs1fAJttOcfm
lH4mmg7HnNQrpQ8R/kJawZYrp2hi7XuDBrc+69rVrW33hkcVZ+ufnFn5N3JIPwBf
cbE7JdY06tj84GkO4RYEMO99/FyUyRT8+JPG9si5XLZLKSudHP0kzbjObGsTv/ym
rMyCUDcQvLgQ+v8d4nG1p5XAs7MOUh/WEnuv3HvVitMHlppbeqymFJOSYVJitZrJ
xsb+JvnIyoqPFpIUyZXFjyWGqb5QjDKMQKcLvKkbGYmeZdSE6gY47S18Gn/5dxU9
53EXf+Lm0R/5QlkNcXWA9cFVt+PNC7loONK1DXE1KBq0HKzIGQcecEHvqrsTNYXj
Ncp4mlX517lvfBxPSGzRakFjpsozAsgG4KDQG52fskpulFCv4Z/fL2QW8d/YZDjx
qunOqQTPZCzBwPF9os59ndd2cwRlKM36/t1SWOXFBx+RjSXvUMkVUOG8pImcqAS5
gCMgocDYn1s9XslLULR8KEQR0cQHOx3jMeayLRuXJArEz8OHNfoimmYfcDE+JttV
HBjlTlYKz5dcrL5Aa0t7M/a5pscpsqb/al6Yn5oIgnmlDbL1mLk90qFOxjQBRAJZ
HMLwzCcW0YYjJMgsmhklO1qG3g0VY92/8ifgajVxil4zoW9m8fp1FEpowoN9Ngz3
pPltsq57cijQkt8AGWbKy3xFgCnlIsFm7ljxOLeDjk6n0xug75T4NOMx70jsOO2L
R7l66rZmR7pL/o4g1667/gml5aMFfyNsxKjTFix0loamZjAAsbOvaK43aPVHRrA5
8Ng1/cTBBLni0NpfLj6zZEfwtE5BdnpmZOE7+q5iUrsKRhnW96ZQhMkL+Fr68ERZ
7h0shfOcfpvCd2KzX9cd+Cs8fss/SsKRep891VXDz9d5O5Bvf/mA6diid2D0XhTt
kS9fTGJjSLez62flCI5L+fUj34gHZfKlhfQlQftymhMhv2PYwT9Nv29mn5i/pLXE
+oHKB2ro2FPni46AcmMyimv9gau9HSavN1h/TxlEMgBUNqi/WNKGnvdtxE9jkH/m
6odc/6iLSw+NQclaVFzu4XXfjC3T/bZ5HhxOQGOTQREUzYnR+N7B5tfd8F+h4pyw
W/0wGX4MX6DY8seJvaQzWKGpO8LhmZ9ZN1+Fzm0GAz5dwOeIIrYf9kwwnDY4eLHb
qu49ENIQHWXe1Zwjh/0prWdxnrM2lV4G2eaEDn/DIvzzDxorx1B8mebEvx5354y6
+tV8J+5hBN07UmCkEtIaP5nrmk9XcLyIQ3jtQZH+xsP/glRgFZqsC0vWrUDUlA45
bBI6q2fR8Y5r9G1556RfzAc0e4lFXHMQiPjVTTMX2IpPoe6HECVT3NwCnC/QQQ/a
3Oe0+c2zeTm1h0m/MxUfXSnLjV23agXZljdyq+R7Hs21BJzdXdAduf/lTgF3v63r
m3v5xYuwe/ks13dgfT/8ZXi/QO2Nq88SAAiJhpLdLr8r6UbvyukfuulauWADTyvU
qNBQj4gUHYpqYJ/Avm9HW6zzPv7gt0rLgn3SLz27L/A9TRGLHwrbv1iECCBZp8Jw
sIMPY1H/NkEVXfpbolL2lAv9c0Dcbx0N1Plyjd22UFNkGho3IiArRFrszZTSANft
XAE7+BNUm4Gs/gt9LwFXTzRor3LeWOOYg1Z4vnzDkfvQM7S6mqSzegf991Hr7h1M
zR1XXkNOZ47u5zQ4CPJv+p8qaEpdmEzfewuSMr0MEqOuibBGvRdsY0NVTu4CY1hW
W1tvbOOG6RUOPEWNigxfTuSOwCUyHEIyLDc8F2r6H45Y2fgGHgPTELAKWszrf1mr
MhWVOQU6sTKOmHoCIkeMqgoTPLmHHIYko6C1bNfwXrGmsZV+VBeRiFkwrJTfPtu3
74BKK989XJGmvR7gq9SO08SQwdsMwqyLrJH5ouAWxj/7bFQnU03nKuaGMC6lSDlC
2nPtud7YIiebIeN+eXGyz05FtH/fRSqYfkRSnJsW3EvxoRBoY0J9Kv1xu5WIrT/f
rKqGS9hDImvnyzaGBuKb/BABop9E9dQ1l3aIaP8wfnSrNtvdzgDHmKGGfw7ZQnHb
yMj0+iiYnY1326G45G83KLXdjjlZ27YOjECQ1KDksQZCtP+6yBNrDPUaklKeUQvN
YPT7C6OqoxoUzjrK12vKuKIN1EV+IahyUpb7qSf2XZUw7LmNWH2bEud7pMWAHRp9
awaW2sg8+slI+Jr4D38FYH/nKUBdHXC7FLCEv6ffhAsfpAx52hVueMztA+vV7OOe
+mMfajD70BWcKOZefxoHFp1ZDl+tVh5l1UUsCkAUzGc6JZLWF7CHfWSHsPWdA27a
SXlMgZCnEPIze5p0szvjVVFA7Li3RGNDYX5KEKIrpqzWiYfNFPJgR8CImLyedltJ
ZLNqySuC7/q7oHnRmV1daVmd++FPRck0fVWzJxHn2mQIhjIvbHCY0UlThN/QiUYG
HgtU4yATqFmKTwKJuSOp2Ki3W9fjqS+0g6CwWBBRBdEokzbQ9LeK9uzRSNAbKz0U
5hOlnN5seSCHb550DkKfdlb60/xTdE13NphuNI+/QuLo98QgZouiJrzgE849Od+I
U7rd9ABBojDeWfpJhwbYHcdEGBStFkwRP8gqaCTsvW/nbqcYCWBqwXw7NHLm2Fkk
swIf68tPhTZtsS2fqOTW2O7SKf089UNJr2IGZl6V6UPnwMvMtqLryxPxav/VLEWl
AxJX2LjwkXyOpVfJuYruTmc3/sPBUld4O4BROxb7sEzVHrfSnK5mpvGvNJJS0MSQ
ic1ZrnKqvDLM0dxitr/pQLjC1Nx/FGmWuWNvYxhTkwodeDOnA1hV7MNSbgYmJ/Oh
Vch+sSmS+hG5MQ1lMRzPwBWa6nxY/G53FG6aS+kxCcpu6SXnOj6pqYYfvJZXDpn8
bfIn2z+7l1QUXi5PpmSR9zQ6VFmcjlVKJ+vrvaTJFIiwrvt6yT1ABdIl9rIFTCZg
V9+3+X+hcd9bkrKMdOJWb5UrAQcc+N4Mp3x1OYsU7r7/qu92ZckHLIfzb6mJlOo9
TrIkpqV/kKptiW4/ddnws+oCmORNvQch01Sz30IxHjtTfPX9H1sccliZjYcF7psQ
FWaW7oyjcRfcgeqQK6ssh7utGoLlQ7aSOBB0RBRUkPypu5MexHcZhSoB2H1Yrr+4
+T3OGxxKpHdhJDVfzjeM2uY8yYyNkjHXzKIoJzbXfjyvtiLYbycMD0LwtJccX1fT
F/DcebpBgqDuqaKZFvjac1JGngsdVvhFbs/EZXp2Nw4r3fCwHMYyA2lpkEyv06Gz
duUQu9/4+xyH12hSCxzqm15XHAkdKyinzvNprCRRSsl+7D8AnfAty0miaXwz/Swp
v1KeIsYq2MGuKQ3Nbax7V4WUz5hHno+ir9YgsdCABQj6i0ILO5v6CPlqM+3cH4td
bd8u3guWgiO2z6tw4nujXyizOQi0gkPjfk+4pjTbmoyIurOgniMWuM58x7Cw1mRS
xChM03i6o9UYiOIQAjkf3pgiY0XhPYoqQKNKsjjmt8lmKkCl2rXm0HEq7e1M2PGQ
O2eIPczj0M18BsnqNep8f6iCc1ub7ulaeIft4fR+bhVU1hvkq1bu1j3ZhLYsHavt
TLAfET0HoZ6RWXKNw8o8nh8oZoyR55vkCfIqBXM1+E3l4kao7Dj/YDdHF7XcYxiz
rncpv0o9jvpOWGkIt2U39kH5e8LC9RQ4gL85jXYg0Nw6C4VUj2Sb0kuziDgoFc3+
YB1h0TAUvZcKgnn28jvoO2LBHS6q/pHAZl0UJXjf5UVEByMturQ0JJUYetxlSLhu
7FyHeDyjYbu+QiLdbjq5zQZenf02qdQ/YNVia7RLPRZouhsd/Sg7PLiqOkOYQyuW
+9BogqpRypZIQHTHY7QyasfzsZJ/0fg95b0h2O4P4d80VI+LI39nQI0FXvL6QTsj
p484T2Rkp5VnNySa5LgvXry2j1GtgtAZPwmBHwzmVzkhNQLH7AH/ETeJq3steULl
L2PLtvGATIz4l8TUS1UZa6F9+HEOGJyJyypwM9oL3TQxSsTrtBQzJ0d0w8W5t8em
y8NoHDCsP4cWGNxky5Ni/56j1vPK2fT/97BMhR0zmGIBezpAMlh65r9UwD0k1uoi
rVouAg/FAEPjjuIk0WXEaaJT8zDsqKpJ3jelyWj6laWxvw7K3iATtfeU/HOGfjI0
j9m0XXW7fvgLy+QQljMKaVPkg7AZUdoEtVgCdwxKdJtRe5qDAxGgMOeADjQMbSlC
m13VClKvpct75Y9ZC8/nPvoaSzrbBtaLWHgHPlqhkzjXAG853QofgHUHyyA5m//l
ByA6fJiB3zVaXPTgn3nI4VbpXvU0rfqmLQTfuR2A/BdoGhohk6WfbDj2fStVrByT
q2WiBl33X8+aLoxbPVe8TTJFTxPdWpLyGCOFgLmexVIKyk3oiXKVaGeRs6275ool
xQt0MXtROKPsYar0jpvZ86xfx4mJ4LjGq1wFSmPy/k1y/OK4Xpnuz2W+h3sK65vg
mRjiT5S2+vZItXjkx53/4ls4rYMFVfgysqf/y8RHqvdE2IWFHBal2Xs538WfBn4w
teNRutuNKu+ahB6pnCkXZO+teNE5Pn5Nxx4KDdvOdNqhqHljXGFk+SgSTh6V5sZn
/KDjsuPMooWxwKhOmV62lbVNIjrQzJUDkCgQ0X8WVVCLA7YAiCtN5gMQ7sqkAoMj
Y2PfIQ+fsyczxjR7VN83QZ+RgccJ6NwFfAE6oJRgaes6rBPS/T02cR4jzJcMsRtE
Ptcrmsha8so9WlqxmEgPuQ2hNcSjwUnRH9YLMK4pES2JzzgCzJV/OHfgbOj4nIQc
DdLYWvVD5BKKwKlKABXhny+Fh73wrRz0cRg2XAjN9rXIoUhz538bUfrVl2eRwWt5
pvBpSGMIH1hjRiA0eLeVnytXrailzw3VW+9/xEHlTV3CYHdyaNymGpdoKgRuuTBn
dom/aEw3i0yUkpxRIpluRzeXEOWaqiz015k1Qc2l7Qegh8xJdYptH1sbNcrxk8MM
7frb4sxrhZAAp90t6iuzjtYlrB2R8eaa5QPS16eY5rCiXnXF4hUvYOZjXl9PjKuf
WpYrl2mOSoidD5DiDbEjG8EklqEBP6FmpGYZ2AOFRY0s2z37US2FLlYbgxnX4QMa
bzY2H0rsmRJ/1R3Jom+AAKINimMY60zurFp0SZhIId7hmyFStTp0VQSwQd7l65YL
iGbu+LVuYcU/WcirrUyg6A34RFo0jNRNO2Lqn4rmAfzgih66sFUWeUXu+2QLQT7E
vrqWe+5jfA+6KNygRiJynhC1QazjyOSt6SRgGvEqQrWpQpPtNoZkfovq1nss/XE2
gfTAkUiJ5qXixQu56AX0kJojRFTEWcXzWVpyOt9JIQ8MN7Xohau7SntnMp/Zs/vs
p0QwETVuetzEi1XiHhCJgm9wBO1UW9+W7XgiAMpGjXlTz0WH41e4uaBEfv0C+lSZ
5kem//FRz5P7tNhG85qxEJM8YCodO8Mb1Dc2vdm8nEoAysndcElobJCLAdYorX1z
hqDf0HABFp/1E302uVDzsVPL/iDB8R1dOKioF1NthNMWz4kcX9F+VOtwQTRkGSm0
r1v4xT63zjDV7Fjm+z56nq7s/+VtsQBTwJODNIEdZLYkgnjYtt5m209lg8CAMIhb
tt8vQOxq/kEKdpK7lX+2ih51GC1ihZs0Gr17k55CR4gd0jr6yAfinsfV/1lncQlK
ydQrGKnepqJqrGC19zo1KMHrXz43C//nOjzLrZO2JosLSF/x1DQBaAtwwssjL9IM
8Yl9cZZLWaD5IxhbhAtbn8sX7th+9/BF91VYmbkTm+gP1fB4zbsmg6+QNqJGm2Pu
xRrkxtpYd4G/ArS3C0Pbgd15iTpn05d4kYb042GjF4RVcwKByR1I3sn4sO7bld0p
d6Vj2EJjc2yb1GYB6KSy5lQqA8M/BRW5DSiWXHqUk+Ur+9mAP4uMpObaxU1O9xPh
IXAbv9MWt0ZJOUEw5Em3nU0sG0jNylPvXtCOPBGTwpJjKh5SsB9249m//enQraCl
Q5Q+GMeRmgKhm3qUKJYb5iJaauI10rVtGRrZS7qrKUYCAnE//SyxX/1J2mRlZKjC
wT3sDkdrKS6Zlq4nBIhMl/AT6J07OJV59IMZf8H1B2vHK6FCnNYvzoDMmdqgQvT1
HRKcvv36qpLBNCPeC7VNGvOJa6osv1YbvmzPgURaI97i0yDYUOk9SWsT9U8qGBg1
252Qp2D/67RCbjSdNRVQMDRS8stItOoQlX4uj/dZdsObiC26NUMq3sd4ARw0wu8w
d1My/YVW+lO/Uc1S+LDJINVigIC1Ffn2WvTdJDsRNJQ2tvVMcYCSZMrr3+wvbXbn
ZchwFdvI7Wt6JiUxtZujmRfOdXzrCBzard1uaWsj44fwoZ3bTJo5PRvddo6VADpq
w2NV4Wlj3dr0RGt+MXjDuy6InNWyxHlMybk+nclt+k89mEMaAa9JFskKgqHGW6H0
vvIZ98g6nNLUaQ0NSEbvzgW3xLlH43FoqosQA3vG0/Nglig2Hrgaz2Zw3/IGzZPC
okOxciAUS+K2szQbGVYncF0fb8rswYxsCZD3so7cjB4MZS3Y+rErX0ijy2KNv60E
d44d+p3FvSUsJ29wvqD0otqfvwZLTrYI/qwunGVtgND0ZLoHvNfT5aWLS8FoH47n
gQcN1yioky7siyePJ/7nU6NNa58sCZ9XLGx10xUtg1YXrNt6VUpDfG5PGoIKNGK+
r96+Ha2RYMy06USCS/ZuHQRQRyhURe9RF7qC3ekkLLIUO3urCnvuC9jFmosKY4Cp
QKwD+sNO2v3V1zQlrV1jKtBGdEOZYDLi56WuGVZBpseLFPKaFS8NdksR1HRg1Y8z
B60RkYFz/cgvTS6lWi7xJS0ul5SYln5gQj2z+pKeIApNKGrpUCGSvlC0S50lZ8n3
deNN0jgZgn6x+OJihrpacP0RPO3fsP5KnHdLj0spXlyc6DFosYjnane62G98sbK+
oJAx1Y2NYgKjl8XgB7OCeHSRihJoMhUx01OB+wV36/dCSeej2C9pZ9n/TgKLQ9pG
FsaZmmOED0CLszy//8sRhN4byfcsdQI5UrBkEzP/nDkDR5i5wJF9xbInXG3olHr1
abks0Oki8491F5vB7NQblmhHcEv0fOl0I/wnrjCnBLn3ZYJwnsP6/mpzhljVMEUi
Sq+E+Uper+S6zJ+CspKLHxl6h5IRi0TqB3vASEpLc3nqGLfUNhabPc+lr5kgz/mF
XM6E7al4VnOik9CZYZl8WdIIUWF4jmw9uonTXvOvkzL4s9DE5h1lTvBiddPc6JFm
d3YfmBzg65oHNk7C5BwZ70na1BcF343oTSAqTko9YlK8D6oUQDDbXGNZSb4gssne
mV+NMfTq5KWc4Nf3lScSnTXdeETTcORZW5qisgzFu8WHdW+Ip5mytuk8gqalv8d6
Y5WtxGS9EUyhFMY5R3ERkSF4yZqMgD6Pd7H9WpuLRiiBG61mkCaxRlL2zteLRibU
3CmeaeIRi7oJE+itKrsrNTRP5BNW9MLf62g2ongUON+SqXfKdjOwyKX/VPw8lN1+
E1I5A8OHxgYlNH0khmMkwD5UwcCNncyaDB5PaAJt7eq+4va0FImvT2vRm5MgYRUC
uYZT34MjsUAS44fWUgF3DsyiYJTxYw5LoXALSGUstvea3HoPmM0LSQiifRDzeMlX
Q5ncNGBlniyJWWmarQl8bPMWl0fKp87s1tvnaN6NpVZ8EoBH5iwcsG6yMFf4P7K0
XQWu2Rl2Lr9hHHxtsxS5toASoiBP+RIYwnNHHs7e61cunpKe9WybWCteoxGK/IPC
wb5o1U/pKNWAOBEzdqwNIAw9AE30A0T122j3PW07McxI2NXaNhhqccd92xtTwqnp
/DG4PHLI1FqP+04nPy8zrcltZnDCBnV1ryPpbG6n30sxERwwSX7FlTWCJgoQuNr0
qmEGBBBIttg9dGhrVXINx+OpyZD7r2MuATIzxXO95kDbfKHxVjlTnjUiwIUIq4gr
U0l0Bpr+JkD5s63HJX9y8uPBTgYZ1E+JYfRcikz/MyK+mVK0D+X6XPlwawW+jNR7
SQah34DDb3YkueyP3oq6fTF8DpY19eaZTCx2D+ITMDeIG7Pe9dJgKxCw94343wJT
7WDzXF6VqbsLlg7JvqfFmslcCto3aV8wLw42Ht9iBumz8tZTxYNdTbFqDTTx+8U9
jBXGDa34Qdd5bGlnhA+cdkpBJXAn/gBEfHbNBX5YEWBdhgHPm5HZiBqU5dO2sIWu
Uicky345yvwHSXFUlxAAvQRRccVN7aJy3NUyx8+TiA5qWVaZ7YirW7Olruh6R7lm
IaY3d1gU/149aDbuAI1HjKERzwfXO+Jidvzj0BsQVPqn+uX5KnSc8dw+/OgyrX+w
mJ4ZqYm0JLpfDPvWLHuTCQr6frepXGaZErwnC5rtfArJ/BqRaDmcAJqjkG0QZ52I
vNciLpGuMcWYJJkZhcn/7j/KaAygxhET10Z0O+PA8owugcQ98sUi8gK27mV3ZLDG
i/yBXGkdSXjTyoBxqIfr6+rl03T09m3oU8bDwCvti1FM91EEPGXX32SnwrzumgDF
3j4PfQrqT4qowS5f54treUZclXKo5aA5z60yY5VFcnJArtgRg4Y5/rcdvkeEBCws
vp5qjJ7bY6azJOeNhMST+d816cOUceBxM04ewOe64vKHY86maI5NugbALAhKGMPn
AT8HWILcvCpaEKuqIWT1C2VBygFfjSuzZ/mkwpon0HHXAbWgj5E4uhM6U7ROjwYR
6qoaIGBva/Er5DX+YA7XMmkTXc2fbEWvXQMzAqhIxVbGnrk5vh4ERZnq40m0xmzH
Kv7hjXW1YYLhOGpQg8rlJrrpJGXN7s8wO1sbbksMrpBkHg/00T4dx6fzxZiv11Vk
Xo+Hfs7kGuCeNk9yKGtOt0QkeTCX+Zf2Cw5fhxEFqLjT1PNHbThWmCkg2e9BE+Gz
hEsffiFFq1wnvg8qNKlvjCDZE1g60lt+kGInSnKG65WXZULYsOPobB4CD1ijiJ2Q
3Kzfjq8IiX20tW/T6g1J+END8DLLLpg6WkJNLjVUso/VRR9HRZgeDeG/c5JPVbsz
YUyJIMCiy8DufS4MEvtYESvS5KWY/pyX0oT9yN+bwFMGWimn8ataXkuG7zLIcgb/
J47taEncKbTT02d/zlShfCCqF6kGz1Ec10CQrbMEqySxA3b3pzEr3WuSLSCvZup2
UjbW0an5y6bV3nvjccJ0RQ/yjLw2IKuEDClvCTrWEi++ZkQY9lDkhauMg2z4pFxl
McZEaLNdwRnBIGCfrJh1VLhCy1sv1WVXKddxDcAhQj9IO7f1+ut2XMkvimb/BRTS
C+Gy/DMLflCfGf9q3A9mEDsuWSkKUZkv0aohI3Ivb+u07tYwLJfk9t9vYRJyQj5F
unheVD8/GTA1SL5eXcuakb1TKUbvQyvznJjvkpnZhmQwTeXIBbYANmzTTHAx/fIE
VivdPkM0+zyKWu1Y2bekOQ4wn4PTSNzbyxKxsAPupR9jOnYl87/4lzw7bJagLMR/
VKR7G/lobjhCZYI/nZ7WmtAjJPhk4sXNJYyTPkjeM6u0UNcxR7NYp0d5l4rNEvsv
CvA4Ahm0vBJ00ErWrYRnpsnLJzva8eT1ENlK6fNfF0gvvMxPISl0OhyyuM7Rihe2
vTQgNQMRXPhoRQVJnGn0QOtzZSAUt63IcQHDhVpUluQrdfJQd8mLORH0VMKXrM3f
Z06c10/JdUFmlwxWX0XOkIZnfgGNUuf8eGRIVZRL0iDX4ob5xNjeJanWoAM96vGr
rkoiGyxsa5G6eemcaxWuHXk3QmjuM7KM8kIW3J4XR4F1AXP4QkgySxyXH3fgPjtx
XTPQ9HVObcBrpitjKkFyCjfEaXSJy6I3EuW0Jwyz7NbSSjyenUrs8K7vBKHwv2Ad
EZol5bbOF0HXOA2boK2I28y2e0VcNw1GA2s/5lWFZYA6Jl1YQIXjq0vP9EHhl2xy
Pv0rTJtOFY9Knc8SKG/wlxnQOhxD/RuUTs/o7oNAfXxIJE2HTfZPjRNbDbYOVxQd
+amDEB4hCO4p40xZiNBssQD23agyWbOT6VI+YJokhSHY+PgceCeWFWrhP2TfFjhG
qXRuVlPQ00/9mT96nBZlVmWRwC6H9Ud5FWOHJC7BRHe96cDQezq8IUD+F2rwPZyr
HjT8FTHsjiUdw08lYSQPydPpvhSWNRvIz3OXB5+RciaEiJy9ZdTlJz/RreUslXbu
e/G2iz8rD/E87pvqIo2bPLkaRdsnmb7VYolXMvftQN6NjloxXIVRi+yCKzbK667j
tpI1e1WDWENElBPzvQSp+WlpDkfCowIViXK+EA4s9b6hmadXjqq3Te7M+q6cm33L
vq2B+bWj1EqvmT3YIKEXYaMRYCO5PaFrvyHGs9ixG6qr0kO6Fazu3lghpMdNCtKU
lbr5TAp0KMFzG9vxhpeZbenMD5PPHt6BJESAN4GFsVZa2tjtwLiH4uVbb1bOS6Q0
1ADRRkrQgJSLtv7YicsUtNdTZ9vhTXvV+Otva6qd9ovRWjwvAbt/8gnuPyunUquB
iF/kqR/peHIBFkwsZxLLLJ9caCHTk3s3pijK15De1W/NrdO6H6YECKRM/Yy9p/Fe
ybRT8wE9IPjU4FdCXYeG2Q2Ex4GAC8lLeq8Pvou0chfOUiI9z1h1BWOf+4Oof8gn
f2QBv+fHwKUo3GhwVL7yzztWpWBnpteruuBXKyKSsTFlonOY4KM5F0SPjHCYK/Hi
/Tht9YIWL+J2ZogGTfszugKkjKJFPy6jjVJI+7p0Zh+lfUxOA0ZlTJRrV27TNWy8
IJABB2aBNba/9K9JKlMgXTgZS397pqUHngOZURQn8spiU2wXkB0YWqMcmG/1ht9E
IfOQg0LCJkPe/TrH8AUmx4/cN7HF8CG4jqgGHxarXyuy1NnZYBF4oMny8xE3txpv
DSp3dJU/FrGnn7E3pqu6jd9ae3mYwrbEp1gh7H+97WhlzH/Mhancfzjl624IC/ly
rHwifXY/gpfDNRaTPPv7pGrZBVN9OPsdNP9kfUoiK4Yh57JzMBxrwwMyQHExMmKn
W/nlzrvPEtTYkqHtH9uGNrnWvlNHdJIzpEewuiyAl7AlgqcR7y3Wvuf+ZLzqt0/j
ppjfKk4CcQd1tUP2+CUFjb8O5qPkkXH0DZ+JjtA4/BhGsfH5VzWOTs96Yjh9psIG
NEoR8EXsNOD7EPp4ABVEo8I1Us9R2AT1w6j/LXNjMNP66AKAUOtPmwuU9RdEbmhb
wj5QoHA3xZWI2tfYEBqglNL2FhfEfAafwPwNba6Hqb9eKtSdBf5b2MnlpJ3xIDQY
5xOU5GK+YC3tH3R+znDLNPKcqnU9efs+Qql3HRhCbscxqBHadUffXi4sLg7AHEFa
tFnwrhRQnWugD/YYdVt2LIbNIhsZLr+40EYBWUwvyI3WlVA9Wcp06qIx0akZewlx
YrCwocydFpkr7lA7cn2f6vUTnUN2hi4LHVm0QZ+jYs5vVkHsKc3MM/pN5g5HggNI
b54wwyGPZuGHx5EQBqz0HM+xb6v/YrVsQr4qEl4Z1oTu09gY3OXzaSycHyREpY0m
Wna369g6mMrZofllNuuVI8YcqLprebW6s1pBTR0a92RGMs5fNqXQxz8ffEplprAI
N73y3TKIMKLbRlm+oclGuCSOjBctSMfiA5FPyH9AksvPlt2eeDAA1nu8XpGgaEyp
z036qCXFJ9qCbx02UoZrYuQ0cVsONSODPgyn4ySnx7ahJ6AryFKu/MklSaG04Tag
hkJ4okl+H4BUeUaefTsgGcmGi23OW1Vi3dOmO27iNNObD2FHelI5wRV1BbcI6LVx
XKduvXhn3EmQszqNxc0zcopmlNcISM5GpgiK4Bq12bhROs/SvvoVl2X2Sd5YeH5s
hyQ2u+8oGaJoKlJGkmeYFvFrJhQNMjRLqxvViu+HZKOzjeuLoE21y+X5wh8uCmKL
aVMXv8mIseUhV0GdMfbcLVfPtlf0xthf8U4sNVUvX8Twl1S/6neCKMlzhZiWgq1D
edX9LhblzvfPit7sLj++xLNUOxZkzc1vis4+E7dl5VEL8GTl0foCYALXXmWUs2vz
8/jBQw3ywupi8o/FM0u+Ug2YtNKyn/EV5tzGdnjgoIv16PzDsQOUPDhYA03lfnDc
N/sdGP3YDrW4o+XxHFBYt8IldaCUVEJLE0HFrEMw6QU7WF8EjkObcSvAqW55WenH
wKqr1ONN8iIPYKJwcka9hJ+h1iOxmVvGOQkngA6S4k+rh8rQFu7PCrCpcCGsMyrv
pm7EyrjGu0SaPOskFrSEOIjmniFILHRkbIwB4xNesOHo1HbzHqRmG4x6HobGWkxT
8dvdsI/EHPfE1TjJP7dxLEUNnVr+u9ajcKXQeB7oIkfJVXJ7lufgOnTQV3wJY6Tt
dv9W1/otWDF1edlp4BMvCwXUrOZy1hSTSMF+7F+jq6TO8LmVRU5BvGFcwYnqchH7
JQSo9sbC6mIQ1iBSncNkJCOeIFJnjSRbmma2D+9CL489iMQGoiLnP/k4JBsdwUXA
dUlLQdc4H1aJx3nnnzcaFxjuoxhAZQ/lGwdsO3jLYdtYi1N3F545xo98AbqXNbnZ
fxdZGIL1wLo1UTEbm0f5Xna0ry9rY6gFBoqHPNnnF5fnoI0++jdQC9Gzlf7VnpZz
upl78tI693k4cxJjvtY6UNrLKE++TpQVyiwYWXBD1irB16F8pzXE+qnbU4ngwxbi
Q/numVAU06WeXhUvhOuhMGzcs6DRaf3VSYHsac82Un/g8i0ULkUXyfrCTBo2f0ex
GnRJhfuBdJpzg+UEvca56fuo5+Ic/miaUE2LSW0Snsh1iKkjpanFmmcx+Qo0Az/q
vAOpLc6y+pfp4tyOGJ82T3RY02UGkRdBmYK8dFL6VL5C/qq1Z29U/lOmw47xXLtS
3sZwB1BdNbz/i3Brd4U+0oT6iWVYobAadlJOnQ2/nawckV6IV2s+HpOtMdkRqcdM
8AsKIT9WWk6tnJngul839gdDzKggiED8sVyjATQ8uEG14X2/wE1SzZrzmAMxeiG+
JyJabM2v9J1Qd/B2qdgQ8SrjbjMQ1BIXi1fVsDLRTXlf76zvtzctdoSgAgLt0pTL
lDwgRFqxttZWy7WKQA4mUn8RCq+7mXs1IGoXpLSEVJpQ7pD2+dnXHpulMubKV99h
IfMiilGv8YvuzTlcpXdGZlBglNTIo3BWgQcvskhnBYkZ8pdErRUu/Fg5o9x75kR+
qjRYsZqrNeNxvJ34DaFB7oqQ9zvfaRp74PIkcqdPOVndd23g6Ziz2I3dye8AG29S
rl5o/RlXm1d6CItXe1Vvwc3roMYJVFNGg2rrFGr3wTxxhk8JYOVSoP57ixBoEYZ8
nyR4Ov1hYCwvlsOlBFE/F76gNHVu8he5XF5Ofu7ovGfd73PPf9/GciueCKiMdQ3E
46qk2KbHvFdJoJ7Bp9qGXvcUydmpWOrXZxLKdNZkfGxjk/lsuRhmWIy6ljyZy2gi
s1iqY4uipTixi+GZnzdUQjluwNvcGCL9ARvbIeBKMj8zRcrGWBI8u/838JKH8zif
UejvKRqNI5Z4nH1dNCa91NmFk1cSDPELC3aGX53sRz3CgGV3/4e+60+BAKzfq1ok
bwuQiYgXjUM9joCISc5BiXXJ53MVyTATaqC8536YSh9qGLDMzKfUuiTvBb0oGnwy
Ov6cw51BFzbKjpVPKZemPYEw/S98DylBqttdBv+npC+J/hXQQu/lpDX+PSUTXdAr
iaHBYuwyLN/rSiftjqn3hkPbpSlqesuPxTvdF3x3gZwTPspeFIYqPVCFlavrl1I9
vgf902Nxkhrdq9Oi5HnUuBR0xAbNAF2Y20jibsDb7oGs9WkR6rAB3eExAWjO8N/3
VuJthXwSEAdZi6uvX+RL/kELVBFHidJqS5f7Pw2sX4tUfnIoQ8mtHMzAJyMk/OvO
9eeBa8mPhlFB4CTdXDCUXGs4U8uCvBMx9V5IbRVNCUxLk8FqXx94UQcKkBcit0TO
bfmtFpWW79yHTxhU6pJIYllLkJwhm81peVCaZvB+wW8gvxAnAdvQTmLrP7XCRUrd
/n6rY4EI1zB7EbKcIgLW0XYADmNwPBQkKXpqkxrX9aWLwiQlwRYzqq804JJBE+zG
RoFkJA22tAff9q2UrKFMCol810BBjYKB2nx3BqEbZbwQ6P5MVhK23DSR/g2OfkOh
qkMrf944dlAANohrV+uZybiXLL9/va8DS7QOgoTBTy8VfMsuZn1nvglubXvvnelV
aRyw+mAJ4rFKF9A8xo1TRYOTVqge4PXmkLTJFssYtswA+WrIeBMYIYpnHRi+wYc7
2q7HeeKQf9RbqmDNlTxbUXCNZ88wWERV1nY/thSI2mE1907Gyf5t7UoSv3mRwJ6T
PmWJBGyHR3wIeotS7b4G58QKWDK3i0wiiNzF79oeuDHj0+h988/W6Nn9WjwlfeOB
2EDwWmuBMmsvSG5wsLFjwcc8xPOz02Huve0RfOaJfE4nQQokE0TBaNNiItBi6ITh
z2U7WxUf94tYlyku/H/K7rEb9BxqO9t9o7OTp2uHpKa6zvI+DhD9LxyzTQe4ML3H
iGxxFyS2ZzqSAKqBA2NzG1rhNEYqfsOVQlxQ6JP6mm0OxoAISaNKeKIyFsgC9mWi
UJhgnM0Epw4Lnhse4YF2mVQCbEIX9nyP7C4LeNZoxCSqFlOB6jPWRoAMKL0nGMTN
HlTTezOh9m71q9h10/Q0Pf4F5QP8i/QVHF2zmup3mLgblWyIlR34mQ4obAl/rjGA
bquM0CQHaBgpW5GQGgPjeQ2WnH0L7SW6xFu+AMCr3CPOrRv0hWcbdplYk0NTLx22
X4pO8HmFIbXiqTAO9f9OWml+ahNRI+pU83hdjpGAts49UrZZLWCnC2UwFvrF+6gZ
5uu8CPBnSoiRKVu4WxOx25le4imxX8aNUBQMEbUESPOL7JrqBVR28vUAL+XbjVzT
oAHjNnHAd4H8m95NI6dAI/FSWPfV9jFFRMahp0AaTjgrtIjTKYS2GGES3eGw4HsP
yOsmu5YWLzyBpQRCDUtP8lRmjz6pmfIPqxONc/P0gUbGCbP3HdQz82nWVQQlpDIW
vUwH48CGPu/luEWyMciEXs2zR0Syy74Y+T4twlXkkBX3wNfI9NXcqftk+nWrgCKP
R9agBHPG01rZLR+KezHni/Ga2RobMA1swziaM0txiJwq+Z1Z+xgsQpzVxvt9llU0
KTvVKd9TlybDqEgLtj7tkCcdfIWQaKqyATAjgA9jiQFIBevuErxIfyemvgHkONXE
Yl5jjWvQKcY2UdmAUNQNxq9rLEQbjhlG5kL6OuT6SSf7Js+Mzb18pX1PklU+KoTQ
Pdz3YpP6SfjpPOa6uAWUT20RkKciHc/AQrJxJycI2UyPHO5sCa2Y7deow7eVU/ee
K26+D9UZiylgEKk3EXcMw+CN9+Y6Jl+7aqpSjBt3EyZHmo4hwAnPzF4bG0jbRsf5
926PTVBb8U0/GELujc+fdxYBP+m/XhL7TIKJ2JZaK05sohuC1o4yUnSiBXmG4ZFw
63/iFM4FSyUZvGox1FLmCJqYiI7dJxZMmemBonBHJp1s4lXY3K9N1pfEP5pUKogT
4WFOs76ArLm/62yCeVUdWZVVltRGqMQA41w7pB2zUhC64diNI5Bbu+goQ49SYwS6
AmU1sDHtuf7S36Un1H0C+kCyhAfZP7SgFYQN+/C6DKvjrd/pN4p5DT9qspMaCrY0
6gKoYIwuj3k/S8vub+I7Gk7/NZrA3Ase74hvaVT4vAUwDkgMN1SNDNXXQyMn1/q1
Jh0RMkAY0yeMIJJDQ/IsRi1BmqUUff29nC3Ut7HkYo76aB6cMO0th8XoVWzweq23
Trf3OKN5IJDmeN2yocRWksN8pt+sogt3TVsgj24ygMa3R1eZ0S0lS4AffUri+1XD
rSr7UbDnKMW7ipnOqMm2yXG8OFV62oL0dV56rQCqfi55lSTwivClCRvj/bnaoCiQ
N0dyHQv+yRDhuacGx3Opr9IVGolYpMAKRkcY+1OgwBAV85pRwxl/uYJbsvX04SFf
aj1+elxmBI0hj1lL3M4fg28eRE/OI7XgNXZ3RQ1foK3AmCOz4WaqJcrYwMr4RcQC
ET0Imv6MiAElhDJMVjbLz9iej71EF31ZFOs0EVjbrpSkybfmBWiP8ouTOx/dAh7I
mGL9Obnys8lhnCuva7e+779DfiOPf8MMhTb5SLgfXHvjKMcCVawI2cY3PM7HQJSx
WXiKFDY9Ex6scXb5Izwv5T5JYopNTWo89uPoMzAtLTdaFK9JLjc5cVes1cyMKBYS
tHpCwvINKMA8C9t933Su3Zt2G3wYzqAv2wmyt3gK0Zt8mQWm+r2KBUTc2XBwo4MT
kbvtXT2NlYLQTsMwwBHFVYR9AKv3DLvGCsvejvtgwa+W2i0HTByd4sBQ/gynbd2r
fGP+aQidFoiOharYFz+z7JUTz/gcuOrHgmNqFa30R7uMWe7xXUILyIYw+jrzt0wk
chUocaegRvGdGK/jQCYWwdGerTRjY7aYgvvdLmFNwSFf1kkuvQKmWZ4W8WQH8/nZ
GlDmiHAG5V9/oR/60Kc4JtYxtpiLKcakFoIvEY3lhfJJ9g/f1lmZ/4Cxscr2Pjzs
IC6UPS4YcgOdYeUoHhNmjeFCANdurEo4G8GeTSVPjLaB/RDdyl2UpCqm7QlthnsT
r6SA7YgJIgnSObuePHMPrBv0uFhEMSMnMxNTU7gkCQ7yierPCZlAAuun+X8GDGIq
ohfRiTBXr6Z6iNA+eijkcXN20MK+zEidPt4duI8C7yJSvMVmDRgneihn2Ntr7IqB
FvEKC0BbHIBFRaUfedTf+y0yiuFLjLdraU4pATGqhVIbjbEjAuWXEzGx4fz8lVHw
xUV+ZXFlAAk+0mZ9nCjoL4/29BF1eMvuZEcETdrBQaXVVIMKLLxUM+0TLWcCEGc4
Q7k+a6lidjcx0uzyAkJYId782nf0tIb/F8NbpLkLL7ckas9H58EzpqzLpdchAmHI
ebXS8oFfB3GquJ/zLHItjQcX5p0hC7FkZB7jW2HSyfD+jmntcJY9sV0IE4iWYQLj
rx9HRG26ueSZ1Ov0ZYmtqMIybFSZxj569E8MolIKuxYlfCQNww2MzDwHQj4sSHbd
AxstYCjFzRVkNlHm9TMgAqtXJvTrF3Rgh1ZJ5X90I3zIvRTanDeyXB9SdJUleJXp
qShXuEuTy9AnI/rja28tGzN3JR31YO+XcAuh7GCssuwuXR0Rsd/uPjhGYrojjB7O
S9oILjgynlDriCwy0Q5Y/0PePu/i1sIeTIegW+KKtlezFB534cyCQwU/Lvz7gI30
yKVxQOK+Y2OPe6kWUdNtmpawrgcGUZD5t4AZBYo5EJ1W6R3dPykbikarioCokgQ1
8nyAnT78YJZRn28pazBcPkTt4PVxaKFj8L0tUuXGgmqAD3rIxhMHbsM2EDN+dJSV
6f8VAFG1TNWlsEMXURbe0MFgiMrGVU4YfrpcNWso3Kk3Gj48QljSmboMTs1ky1MN
yTdQKWurK1vzPFv1YReJlAec1mc1a+4rUDB3zp/CAUpeJwM023tUKRIF69+hLn71
udfo0YlktgBbfAvC6UeBi04mfhiW7qa6huZkLbzXmtPoKfDBfo+oJcwdN0z1SkvC
+v/P+mxHsM3k6I5s7AO5mkJjnWUQ0myuqeOYxuMejzaD4QjsXeSuSZq0rARY2ogA
MRbdwbf2zEdPHp+y284Ii0bYumV5PX7DdAFHDVFMTDcD4H6zfasgs4vEBwP5FxGC
fID6D312oKi2DthgqpKvosImhDD6+57wA0UcVbWRYxby0A/CHALqLZtawD1F4kmb
8FCb2rUQC+MMusNx2B1QEiaLVh6v+a0UcTN2Rcfxeei0ZXEZlHFHc7x9LjiPWaGi
6HjseeumMTf5DflE5afqh+vlNZepO18D3Biyt7ff9C5ym0C9590gzsm8L5ZdxWrm
1qGMiBRmgRgwR1u5UJ04Z9j1GWYApZLimXQ8zTYOSAgw3DOFQGcEYsk+4J+pyS71
0Gmld4efOdyUesQIw4KeQBIwvG45n66C7gXDfKDNmhzxFm3T0l8yckx4e7MYkzh4
qR2lS/BqnoNIDzwuYExP7I1l2CF0ZLmvvdpVzxoapx987ulP2xc6WqAZjR5diY7X
qDPCojFTS8YgpLWYfSMLcCBLS1Kq9EU+vGnuCIq3MUoB202ULKrfE2CfMwxNeDi4
5IrLc2IZdXm9HBoVj2HcA1db7/cNIo+99tdQ/c1Uxu9ElwinA4G7ByxS6ng5qqGu
Dx1YNr4Jn91MEcy1gNB+FLfNLOc4Ijef5F/rvTPJuCnsmNGyqBhWG5AVLKB2xsRr
iwoAbUN3Amt760I/v+FUKcGAA2Msm3X0Qvrv/PsgEht7FyAs9ZPA2lxbDjxWOsn7
ZJIJP+DQ+woQGR7+GU1g1GIjQJ1MJ4Wzt8hZbS7wrbZlWWhxtYj9W/kKufCjAKQD
85UfJE79KSBqv5L5k9y6qiHG98fosBsMheN8GSFnYvjbrE0IdSsrkIHT6+Jksod4
Hw6d3e/QTwcKKULgWnTmaTst3P2ggPBoqH4SEW5CD8rq/SIYB/QBagDMdznCQyVf
rWUpqGZrEa3HKl9KaBUf5QbhmogFdLPgVfcFZ3cEcetu58WVjGe/59nbobfS52yk
gHQN1Cc6vgwG3yvsDzhYuDYD/PrdicgbqSfmwnK41Sken5ry5otncuPRr63CtTmk
/pmls2YQZ3Jl+sFeaAesfHunTJ9aoyEklw02XL8blu/WVrY9JD9xQIIQgNrcANaJ
fSTZlpub8mwJ7p1Unb8l1Yl+hG/CeU+CILt9s6Chq0bhLJD38aktNCXZHAXGcC6M
0SU1iYehKX0L78jD3SU9Y44qDY2XXCNWPigFMQOHj39s6msgSiiCP67RG2FKxVU3
6UZCBChEHai+yRldMOgrPwSoIbJxOsJUmXEYx9g1PtlK9C0kr8QD6a7kbcnj3X9K
wmbBG7S7yL+KEd9oM2hyyhtkyffx4rU5mzUbmBTG4tVjb2+XHbyulMilc5+Nl9o8
2DTpJVShT3yxiLQ8/oTDel2LnOJReTVfC/DGLr5AZXUIEZ8DzMnFlJYaVDcFIl9F
b89PAj95s4R/NKWtVr5qIRl8WgXf1ma2amWyFJmDlA8MRLKFV0fyoMuYKTfVEa8S
9Brpyui5u1v3QWJB+w8MLVUhLfu+6XlKe52/lJQvKwvXA5PaV4Is5Un7+miiorhG
TR10opNaufDFE7sZ77TNQNLwYZonvp0IR90vitrX1CfjZSyzg3ri97/Bg8E0FNZT
K0nsXNSnT91bCuLGvJos712zO79RtwziciyczQqo10/XOaBBRd2QwPzL5m/TcMxW
b5gJOQkdpgnUfOTiR32g9akmErpwZpA1Z9BYJWIM/sfCKU/gkj5kZ9ibUuODIP8r
ZcCx9f5RKlBq0SYyFksfGhVTmDPcMTKocAKZmzYg6P+/Jp6P8/iUVvCVcK5Fb94D
UWK/gnMfH7orr583hJm2Sg8z/OtSmTptFiQaa0kM1W/3ABPCV/+T0IGFYZh3tnXh
dbDgPviAxQBFB0eISIgiJispPhfck4GWtvM+DsCctgdaIIemQ9MAyhthyl4YOUy9
JfDY+eKtd0txq8R6bsl1AdvqgENuPeLjlfGisUAqNxZG5+aL9n/tq8kJZTq/25zo
xQGTSewt6iwOVi0Bisrvmob5QbJAR600nXCYIAbdXfhe24PQQ3fy5ayGVWxPH5rn
qAyxOFVfTbELcVQm/gvOLv4e3HEOYnMKVttat89s+v6UWCu7O49M5ZAhSHVK56ZK
v9FG4ROmnPLd7prfZrBqcddsp/gze732DVfIF7NkxL82bw3Rut+y+RpK/ZayRpdt
yo+f1cSBd21ubaiUMMjB4MdevmNJNr5h+ImlN/zU84ch1exbbOdZRBgbdyrn5CVC
Pdt3WClykJLZmKnJ/Q88Jmi3jfxLxlVucOlf8qAR1vZt1txIhjjoa7EuZkz1Zy85
zf+Xzbr0x5WEsevVf0n2jGsLt4DwOKYNG88G7JZwS7U62mcsZQjggUFSkr5gsGPu
Ol07UV2BFEglAs+FYsOa16jKjpvxc2jBS739USkLX/rGIN0mHQwIiy036UJW7W+O
7RX0gD7mkMiidTul8RQdMtnR+5VwLPn10Mjrwf+ZYlBG7qe8Tk8jbYcdEpl4sQNG
TZR7uW23NX5O6xF6wBT3J0KHvPk0Z8VWfXEfw1vXh/wKkRBO6LglCw7LYMttiNYt
UlV9tJvyasogOYbfLlmaY9U5vlw+elUDislgGco9/VIS8FCn9YrzsD5raH4o9/r2
dhtod6Fy1IhWZdX65YXxUd6w0oQGomeNOjM7+PBRQgLe5DXRyDIAU4xTh9+scLZg
5Qtjp8Zj36dNB6UMsCzs3dgtTV35gBa1Wq64O/ce2FSHZt6fIbGUdSolV9DL2xFV
bemCyY1D+Hl+LNVxeoX1j51SA3CI7jTuvp6iOJWnWheX0FjrqrGqAWgHh45XvK0d
aM+Q2k+rOLH54yZQFtcUuDIgNGGtu4TYRjO8jCYt6F0GaoVx69OG9UiVV8QSHE37
clDBN02lDMk8+FziGz6OxfvWPrqtvxvvPpgumf/9COW2Q8WqobT3kbQRDp6hifII
a02RH9+EMYBz8cRNnwpPBRxyW/sARmaZ0UwC2Ug1yGAKxR7bIYJ7x6aFtVH7dQhy
fo82j/qLb+dlvbuCSMWRX8TH5CoQWgTaTaOL+FO9yrdMXztg/65eG7l48Dj+0a/j
Apyp462AE/tDDLP0MwN738BwLBeibstW1ZM00IBLPolueDCe4AZXk4i7CeWFmO3p
hMPAzuGiQOekcYYpay9/QJ7Zcvdcl2uJAlwVaU4nU6yGRZeHcN/zXEkXAiuqu8qt
lZUMFSj2ImayurlNfPPFYee4iG98VTjxD14oyavlKi10DVamXfoaUXY2HeV+b5HF
lWb99MxNfYpRfZHZEdpzfDpeEtGqOIJxMlUvUn4ihZ/6bN5CqmzoIyfQuIzChNvX
DX6BwNiC4UQLXwgcU0ieLLubxB9HolBxCvs7LNz1Qw4Tpboe37HehjA/CABEpG3X
hGDr3bWVbXLWDyFj1+GAny2iJQhCwuyl06+71ozpKqQpfZfhUamXBhjy6leAcads
eekJmcWU/19vIlDHDHHK6dDz1iO2g92s4HjV0UQL+myvxI1n9uBskTmkE+Zdgo1F
sZTJzrH19TERUXVzMo/hl+5pYYt2b6gnIFNip417fRMoIEeAbQfHeT4xz2mYq2n/
ZJDQ2b9H2GeVuyewo+altn+DaSIi/XAL8pdCHkQnnB29JUxBpFjy4q6XYrgw6ON8
VuUTrrYWFJld127N1a5/xNqomFzht8fbG5p4Y6IZOJS+dRuvc2nlRxzidCcpUyJ1
Jkdevga6ggv8WmHztpDHXLg4WT1lEI54JNr26m8aSdiOlSOVEA6jOiWlzXCl7SPY
YyaH+jMweeO+ISUn5nMmevWNV+E/Kv6kheh9IE+tqes7+gW85j7Tkw9PSAAF68Sk
SWoy8DwBUGb+5iOkbhTxPcGXJbV1jXWivYlVLRU3ASqD8ISogrXdtSDBHVYvoBsb
pL5Lys7K/TyJc/I+h1cUDigpwE8ugf1DGZ30cPlvftSyL8c4wwKt/0VUc5O/rmfE
uAocuvURyd8eGFDSjzcXS0arAeab9p+VakT+LE7wMxs70OBoHTG5uGSTmwcVfn9B
14NIYUQRRc1GxpXIMdz5KUKkQu+mF2WCJi8z7ke/3n/0bJNEIqQuxUbkRB+yw7G7
Qs3ON2mn7NFowocmJ41dOHttPP3Wm0kEPtNyrZzQ0Ilj+ksEFKAPHUfSZZRFPQrL
xotpejkIDSQOa4TN3756esxrWDgBmWYldnKUXvDzTW1vVlpbpICtn/HX0mPn6D7I
Cvbu7zn9Bb9CVUPQZTYwtsTpgXnu1u5algpfNcUetue1HiAWZ+nyf0yRX1ZCyl9A
3dnd14kKeM9UDpGpEecUd/D0GVT/Nd9E7zX2s26xzcHpbC0PuF/kZjZ+7NuJH/Hf
ZoRS2mD3QQt2/4+gtHYHwWvMYUQ45kfJXiI18DGvnFYH4EJ0sAICRoRtL4ceSkD3
b0AxhY17e3gIRfu1ERP6RQDa3GfGdEOHFmkzkQ93tLAcUnpyQ6Yd8t0RuXylJ63H
RPnHtniwdM6QuCosSb1o0Wfd3zOStWAmNSFQmG/rw20V+W5lwSWZdwmdGpS3+U0v
l9rYm87LX301M/34p71EcYzakjOnZ2jXJudwNRsrZ+GtFuIIB+znwEcqPobGhVOB
521sNeZE3WejyeIjI9rxmC7J7i4Qyl7XSyt2Xad3eQfux4yI8b3Gw1uNp4Rs7wGO
MBXeVYmxDuDmEv5HW9DCw7ohyi5mf1e2DK3DU2rJKSPEXX7E6pHKGfWfOGdKaG4E
67+js6h5o0ZWBiNwrOf0Kf3mWI6OJocqyCHKMdp65nzpmge+AY4OVQO/03u9P9OK
hGHB/XAuPIqGxqeMhBklp6QYBNJyilj96Hi2Z6MXXCUvfN5Md6GDluSV2hfeTf+i
zg//5cIbVNI8ephvMWu4ienNmV72CEgg9CwwH+asyoYMR1UFAVEBlnX4ovYdZONx
FFKWmi1E+xN5jiMavcOlLzWf9A6YQeQ5gm+8yzKDECDea/ZJiNZMCyCf69AUY2dJ
RdSQ6iaokzc9Gsci/H3A2M+Ka4IPKUODAeCnC/yYt4y7MIZu9aMYO4WhznYZpPTo
ETqN1JE7tNz8n2L6MTwpCVPYkNzC0LrAv1VtDuhaIVYhdubWztr54tgEK47Y3GMG
NCHGGHPqtYL/HPJ7k9FXhaY0ygC2IndcKbphNG1S3LDwWDcIxAQTZkrWL3eDT3a0
0qoxWRVtwJdd+/zFitBSQsB0lctuwQweIjSzVa5xBNbnF2v5PZkUcyq+JracoUeC
EwWiTiFKfySd3QYIbbGs2baQ75ufKmpXhCiUW8zw1aF6ySZlsqPJ1qMqd5RfDI82
RpBZtvQfYpPQ1wzw2fHOaaReOhaa5oyEOkZGfjU8w8reogRRvDqvuF01oLJAmpYh
9uZNSVMsCYHzf7Qy/W2XfU3MissH2/MAO974qAhrfH3d2WpcO+dTJlSnWYOAo8qw
xBmCDmvsKC75Q1gBJFLsexMbkvWqn+L8hcIuzuKAEFp4k9TJuIRFr9TEsiaQRXKW
p8J31bovHW1LnGUQRRA3I2ec1vbbkyH2xMtMjXHzQsz8dXxT/4BcDjOtovoZxl9n
0x68nCyJwYvWgbbRg+YzRUR7agV01IpVCLpoXJM6iW5ONX/8Cam+AzTXpZiFY8d6
EmieYkh+kgMMABs+VR83WxuYrRGETp2uDerS6NWCEihKdqm1p3IbsC+f2XF9r3NC
/Ngha0unSZKmUszG70cGqswbkMMuzpuNkXNaKVI3+z1ZTtU5gwS/BeqSOC4nKFwb
totig+7cwmZ7NbwRHA7aXn5uUSco8djNfZM7CG8HpxpTC6qbggOMMJJxRYsXVv+U
3XkYUDwZCVXU2WEYhwipV7I/+j+hmbG7QH7X2NP48gVIBUKwgRlKOrOQW2ZWHMWP
uiuROZXH0Y6WaKivdrAXMW9QZyKPG9ZwERrtIl+kmivmrrEXFYLvCPxKkX+us91o
4tJcF5t+4mWUxdnFvsv9OTzyrKG5r8NkeD4l9bptDXCaXWzmARUecZZ15EveNd40
/1pXVY6jGDFebZ+jXCrIEEFAMZa1xnRGdyJEVp/bisS3Hzt43Rf24RnRCMUJlPuZ
nWXp/FJ1D/rf69d9fa0XssSuTCcuSU7tSfSW1Q+3HgECpGFW+V+CEQTPIs0CXlUt
rrEurovt/p5gs6Ymb+qHAku1J4wfNh35HjAaiFR4uhEJfRtn4k+o19sapM86tI8N
fGYeU5hbRBtOPzCn2e8AHQRZYyfNagUCGNTTxoM50+bqisL0nGvKai2Ol+TR9134
2vX1VrKGr1B3kcRov9j5bQ0FJHdIcvbYVNJgYoFrxi39/w6qpVN/JUOkYFYDUebk
r6ECyQaLqtZyLURm+kI1nMVt+GNjxV/EO/WExTYKYICu3ERno2M5gzjHIRVh9sAg
KCvHXXUWBsAwARzPlr9F6rJ1/KgES8qPCJdNr+xOJN121goD/QNpiz8+ZVt8nyJZ
LxG2w5rEDhiH/Eb6V+MKg8+cQ8X7PPKDlJk8iFCz+O+CSNQR5DYz6l/1CX3Sx1Wd
XNvW5EiFphS3vxm2XC5AhtWXOQKIRcFIkNfwB8qoi70EAs7Toj3I/gK2I7cYhcN+
MQYQEMWS//MSLw9T1c6ISa9LtVObLwQu9lPQsTykfenNVu+h7B72FKNVAJXKmBit
x7FWlfB93suGkXgm/b62BkBXD1ugNbbx/ouNMA0Owg3kQJrAu64vnuO+bRV+KPBy
v7dfLr59qXuRaqcrE3Jjl3RsiBfxcitOO2uisbu0Du8yjNPW2S0Lv4JdBygljmqk
ALdNFHWRPWCKp34BQXMWibmR7HUB/00HMNaqRI/dcQhcOxvJ5wwXlDtfQDjt/wr6
2YJo2mlwH7j2Ls+U15PZbDhRasVOAb2Uh97gT3Zc19VKYdSWQHJyR+1UcScA+XVd
opPdNTm5tiMVEdJOv+nDhPsD+wmjAHc+dTDW0Jxlm7hk2KUnAaZLEtIvcfHiyQdp
NOWm83iFLeaDs/ybSzBDW7OeXAfEyH5jwx8BTW4ZtTTrnF81fDmDcBbZVXutaFms
mGEWVaj6xuF809Xi8pdp0otrRSkpRLU89kZtu4ap15cqmTr19Fp327ElAOydIGKd
zNdcxan98F1qb7raJkwBoocTE1g3gi9camsmqvDvo88iW6RJHTKOn+YwAnfUZoBu
qJmganPOotegVryMHj5f6Z1ik0PWYoDiid7vF0kB8o9In9jVDb9kGhLAWFNwF6sz
FDGdyBt6ewdZBqzHL2loQqWEieFOiMBcQAmMtcWMOsdTd4buLgyCFYtIbfshriNN
grpWxV9j5QtZR/NxyS03uCORptezG+tR+J+rXWZyx8XmZejFXUn+LLWRHQCu/VsI
hXcFnzto/P3prXbg+CEhLjjKQLPXnsWDkLvnI7Rd/KYDbdZOz7phZHgTKHKNu/hl
TrI/d9MJqaOod7tvBtv0kBebjjOMZco5FAskKPf66nPfnwRQxyMCky/rXJMp4Bed
ZALryR6UamHOg1/Tz8aaaxQwukbz9QTlGoayF4sq5LC2kevMOyzJfJ524laFlrsm
ziDA2zh68l1NupTZBKPVB30S06Jj90+KUkm1KmpjTZ4TT0JhRGFTTs3GtPtWyIWS
ACScpAOCvOjaXulldVnfy621YlfWbBh3u/9gTpQbhk8DWwJdX31i+Xcopo4Y3rks
qx8nHfRT52oofQ33K9g2C42ZBlBbUlVBZpZq1sOQ7fZAqw9KYT7ulqTrcTCBVkNG
YhNCZw7h5oPV3D+q9tQLQcUvyg2+1LebuVTFl+LxojIQd5JObe7ZEGxyPrvxs3g+
6KwifybYceN8Rl9NQVwTnl9zF6Z0LSk6fQjbOnyZQGaps+DCtnjV3v4LXwbbrZFP
ThAJ2NHBYiKoOBRqXoB14W761D7KHKSMteRjSZBMtTMWBIc83djTOSUeQc/NfBYc
LOYVRt3nj6QSDaEBb8DnlCT55c+6HPTWsprbjX4tqGTbw0rRc1m3ZEyR/OPe6FFV
50/0or6R3uckF1sFayzoyuHU5pjxk4WFYLortJiCyquJAH7Do/iJyFJxZ3cvYeyd
UKsWOKhjDCBXEGVptm/mwntPdYNX7Jyul424NeWwrOwelaA7IGYpD0rH/IzkvP3s
dhH4bwW+xqd4dBRaftXbWn8zt9Z3RhE2QwVSuZ1N08JERGaVOUJpUHlEht9q+AIT
j+qjGf1rtHBLuuzrJaNsDdJ1UzlkAniifEWxvwveMoLcw5/yxnCzwhpFy8v78H3m
0msNswFqjgunMciC2l9I3xBbypQwdWrGEVMDMz1VopkZsYbq9WwmXben50thvqwJ
NGzvGKLwMxMtmczUyW94h3CSF4D7PBImtQknkNQk+y7O00dxbfArxHN7TACJoaWj
HHV3CF+zAkbC60f1xAa9MKEOTPAedNG9CLMfd1hd9pjG86HV2DrP496gsyVHLi/N
IAX2Fqy2tdkASdNTQdW+douqKASm4pfE0I4ZqmxFLQ+234LZ+tF4Rmohejjbp68I
msYa9IHWXycqHYkU/vfvCnvDPHoPa+3FUnMgJxWUJkXqB/5jiPvB5tFW1oj/LD9G
3F9EkLuBK95wxJINznkqSKlc2iymmYvXEJql3Zgr5sbBZuVUkU9ty6sO2SLZfwSz
2c1JUDreHeMoCuMmNCX5S2bOlB3Df82xwLbyVlwquUyInW8K7rJL5fTGF9nwmC5L
FJJFa9oEW/TCr9FQG+NYCpabqbZfhktWFoGDsN4ecO3/MKNRU9mFdqX0Der4qlrN
4VDpLxK40cYTEnqlF21NnUjgf5z5qCOy9qn4YFy9u/paLXel7lXBBHX0MxQ+Eqrs
ih6yXLo4dvTSzAHS1ZcKMqdsqJR4LfBuKqxZRH94qqnqngjfb5tFqUXiPf++Ndl4
vMxUXfRRykMYbm/CUjfLdU6pVfuGJQLBcrtRkwiOQpULKEZyJxFCvGJWGXzbWp1c
0kYqCRHjUDRLFmFw7jA6np1IK0FWsbawhs6oV6zjOITCcc8zOVaVm8pVDfY4U18J
TN9yZ1oSN9TPO1w3UUN5Fb4GvAMHENGqgW7xgozKV+IxOMqVJ/lqEcWOGkttbyQG
sywUBEbXyvwyG2IkXzfcYMsOTm4qeR9hAFhRtniPxsag0q2fWAYoe+Ah0DokT63Z
5KKKVksJFKHLcubXUMl9uJN8E3UgUZ6dtvHuos6vJgpaG7YortP+cewF74xobm12
W353Qui7aIHR7jKXyLpst9szQFqTU23DW4DulYAdkI33of3r58gEg70QDOLdHPhn
PcnIY+mB1B3EtVe/uEGBJiQpCPH6NmzmoOB4f0HPOt+g9QcelKCoCfxMK5nNjN8H
h1NroKd+KgzmIOyW/qZv5rAJgcVoTg4Rj0uc1ZiVMWsTiDnj/ytQ9DWLhkJ9Tdue
d95E8Xh7sfaixswV7y7y0/8J9YHkCnWmE0J0109YeVj0vHqvlC/S5Wfjbk135AYy
sZW8VjFgJVYTQPtnDhxJHvTy4vQGtQdqHYXv5hM8lAinTXzZGtjEqv/wyalo9Ijl
FX7VYwoJeFbBaxQr2EHSqWf4RW653i8qyJhOId6noaM0O1J3xextgz71gB9wFsFv
ZmDxGqepQ4Sp56hlg5bD4rRjFdVinZByTzMtmN3I37Bjeg4tutpiAc4T0sGPQtUs
DbryhSjHTNAZK1+l0UyvkLuIE4ZUe9wdKdZ8rFy9EYDYDjiIlu5dVw8aOpFSFx8p
/39MNrS0shxIq/pyZn/jSaEYUZ98KPguD1QhbQCmd/YUXcA53wYGBE2IKleMbQKN
+VzxMkH+eEnydLhOoP6zs93JIAymmPm990TB66Yr6DWvI1lLIGkm3nDOlqHYmek7
2St2NKLxXDJdvkLQ25NGzWmOLbc4/Mv3iVDVY/xi3bicoMRerSdgLN/mkaEqcmHO
DgfqhzmGQE57VAGiGiM+zqNwxmfNokxBi5UJcXNXXFf7j33O5RktQe9OCTBl1zhW
kOgoNg9FXV4bg76/8v6KJERnuK+Dj/wUGmIticIZCb2PBo1VCuDegcmNJeN9uZno
zlx60nG4e3XASS/p38cKd1ij9ewA6KHWnupsx/GqTOlRvYxffUrE8sanKWe4qN0C
8XDXtFOK0gpJMcaZ772hZjERPMxpeKyEHHpkQXHh9muxkRHE+v37ImeeJ91kHmd6
weo9LjzTo9sU5wSHKnikktM9JuyYjhugMNodzQk5M8z5BosEGQcXXQ4RZu28AqBp
0ScWEen/RnhoZMyRGm7OErReSnmIeIUYN+/Jn7aFyE2sI1ZWmxkfw4vUGGEmNdON
z/FOGIO/vi+y16s5XRSzg3me2DYAE4dkTtoiGxJQ+dJRFp8RahQdoWu3dJpvnQBm
yBY/INc+X5C8nlO8GYHbDstqyxsMJzIqIGktR2SFJYEApzXXRMNLOjGPyv4nqsiC
zqasv9xB3U24YXUwtu8cZ8kqUXui9tAw5kKzwE54kSR9fajZB5KlM9iZWq37UnxG
OY8L/UQBSV726eDGQF4HyDe6jaFXtLBN9qZsxkxNGWybYGSNN2vUKZkUulGnJb7d
Jo7k7/W5YBWs0SVtLxdb2iMwC585zrTHRrz6uLoWnfVuD6n7eFRB4nvtgAsqabpX
H0eonuG+Z82wD8CUBaz5cJite60wZiX+XjSk1PTC4TuVcwX7/2U5aDjhUD6fOgqu
VA94Amk2gicA9mjHOLI9PVVPV1dQt5LKDsEzvHx8kwbJUvY3BYRE8LuzcdaJOFCI
YS0hg6YIAhEFd5Pb8UZzXXm3ClERlTF/MAcywokNclvMLPC3ZUNWbDvfwAmEONlh
qqo9coNZaybLk4IXnUQ50Ww9bSn3w5+TwsUWNcujOZcF5Qcpth5CdPIpRZtDilz5
YqtS9dYEeidhvkm/mXzn+P3A8WcIpcFAufb6F3qe8U2no/kFFlL4KZQebtaqKokb
ssx8C//K8uZXHmAUlvePUWwJPFXi4ho3rOHiNQp0+NSYJpACdrCqwPRyi3OAZucM
VOpNFrsXIJIEqfaMwuCD5N/eRb/g9Mw32TBBZQSiZHiKzHDQJflEQ6NXBe1ngUpu
rqPU92LfN+URofN4FXHtBAJQb6ulQZVHA0QPTdZHbeq7TIAP4urHw0oBa50I6RIU
UV84zzOUbXL7eL4waWN5fsPEpCslSvJ4uCNELbBb3lU1SicprZFNJVRQaoeftvnO
RhPp+ig1/1xWpng+FWxG/KZcNQnJFLdw5hOew8145igFjrFpROztQD+ASSEVy30p
RJCjYiWrFJXvqenQfL8pL6mSlzRqtkICOVEV6V0PxMSt870RJuz8QvgpweIyfMyp
ThniZaOTpfi7xFPtWLXvAwLmTVGrglooeFDYaYcJuWTlSi2flxsUTwT6FtiCHXwz
rWflED3IGxKFR4ZBBg6JVX3Y+/41y2TmiUIp28G5gf7FW2cSoLRiHJh2qRVvWtKd
rWDL9pyivT3tpVzyGBQpEOi5e3JFr9oRA78vIH8wv7r3NHc1Mx9wIOR2LUZ/r9X8
FxUZQgvrZ7PfJ7iGZEgu7eMTlT+F0RWiNRrQ9kBvMqzYLNg4t6f2rus1CP0JKhfC
WWkD7qsMpzOuU0BeqlTWJE3n3qzm3hQPca8z6cJKUfiQpXcOsXOWfONdL492VEAh
Q2POUsxqpAKrSAdQYnHAbavI7D/Yh8HXOoDdU1s4QLH+NnjoyHjrKn7ARl9ydZ1x
vnE4ZRtVrxN1xlNnfBvFZJX1gj8dUn3aHs5xHHu6563WaBj25IMCvj5MmTZJBaPl
JPoINyRsf6BDst+t3z5cIdzrbvTYGXnqQPLvMmYGyNMumKmuluPn5mLMeK181Ewy
cOa3fBfWLVRv6RKwMEt00NXWIWBkmxgBmsNM3GI2Hibw5IiLCFRuXK1JqvU+pkIY
Lrq9pt15s5MuLUwnyvvA1kDiJl+wIGE8ibcPRVDollsVOPAr8222E4PniyC2E0JN
33L9l4HdLpMSF6cVotRAic6w1Tv0+S4amD6DO802LUunupK6eoVfD9NH9/sdAOJ+
MGEN4bDLmdPqc/6n45yujetGsN4DsegduLZHwvGzGdIp1Sd3d2kra6T7wpad/f7B
mSZ7rOW9Wtm0J+eW6ayAE2Z/Oh1RMTbZ7h+4nUVlqfIEUBprrPf6Aq3nxMhwnTnF
Ky1YJkBnEYXKbtu/IeIR+TZ8mRuq5PiUkBZ1il2xJK9sTH70Nzs1Ih2HRwz/WGDP
EZawxVDoBg3DG9ttztChqP+0wzxUEjb/TbNXKCRuDp3jCPa+8yVzT8qUh505e/NA
cBOixWfsgC9du9wtDwb93uXw5przVwGwqDAsLws7aVyoUhiF3HY2Ta3z9Mwu2f2W
3cYq6OH60cyIkOLvI6/MTnp1/9B9guGiO3RJshjbDhF+1+CjuUpHo6a/T0+q9zY7
qdGzJaBcwA4NeAz28y+ll8W/nUR3gPd4wefe/lQ89eIVo9aqlDHjVDtjezk4W1cK
aqhT83zXBev60HOFIhFtrt+RiNyP6v8QcWIZdkgJ6Ncv3YtFHSC5TXn4vP0Gr2km
Gyg2sOPNS8JvzuzgXE8mIuII4khQ6sUPpKTHcWv5r1kniPGqFxell7Vv7WI89vq5
cvKAK104k4EnctSZZ6ywXmkJmROsjPp2tXmbq6cJFGVzp786UcNaOllvRDE+Qnca
eMchzWzY0zcTkTvJKYujxi2DIODBr+Y7C9SWwaLAq2LHZonGg/Q8SjuD7BC7COb7
HxuyX10qwyasQub0NpHuGjP0rAfiPnmLCAPVo6uXEfvYSDWPYyCetP8CuBvSVXmT
XaigsVkw9u3TefSBIp/8+2IgFE7UyMY/kl7vywZGNc+madYOcEJYnGLkZ0vX8uOI
yvGcnVSgfLSNPTscdodt+1bogQQkiBMjmncr0ucsy6UJXWouvIx/nSCPCz4IlTKn
IklTbZvo/jHhsSUSbyXInyQO8vZRQ5xHQu8iaw5XjO4niZRuUGlzGqa413caadpc
bVvn7DOc7tuKCqtDNEIEiyXCBRNLwgUAjEByWT+DaVZ7LZWLf6AX+bvknX/5mrko
HGyrOJ5BxFfnDmfBRmh1ld+EOzSbgV8fUpz1/eTbXcJGsJWnwfWD9vZcc7bXGTJG
6QLLRvhZsy8Iwfa2AnHso6yziXj0233ueqlzI1lbp/tV2oSgsMaF5V+Q/vTL3hlT
SiGkVPexpHKPloNUwrOFiht2NcuhizvRUmHzRmBeAKJnK8QfS+F7eYF7Xvy5CxUR
r/AI0gmWKVVVnNhwdVzOpwqknvAFzb98dRQCvVqz66ceukqDQQgP04JGxrNc0qBJ
nPR1swuLJWaUo7EymNvhQg2KJzz0c5meGYgveIPhrc6yzP4TbXQIIarquOSnHzVy
thd8zRwOcEXCSu6IsgJFo8oOaVmjN0/Mgsabx67SaE279RbQ6/LwL32exIqzffe/
TPspu5e9McAA7j8q9tq2RjWZisfOwQxuCOP2BHmNw2xi7+1ykGepDMwwKZZhqNd6
oRH9DoUi4yM7VDCG01LYyJFNM/pIP8/KPKJisKrCe0kyXL2Pe4/A2LqngnlhMbnG
4E1uqwE0PLKH6NUhgBE/Mj6ayFVAJ0xV5I7tLCzFuOke28k/nhoE+lrp4nEQcx9M
1E7ytRtB38dNyxnr/NL1wEe5GWk8t7eoGMoXyD1OocJzhBqY3UQElh60d0SQSxci
tyUVy6yyeOq0nPQOem2TpZDGNaRUEGea/H93SMYBqkSjQNvZ9qi8v0z7WNMTlkWP
41LbVOKSudCTf2uvvU64jCHwNGX0WPHj23SmKtsB3gZ5FGNenqT6Z2xCGytL71HT
2tasT5HcFsrO6HZzlpATmVrwY7zXkf+/ecYZ7B2p1nEmgOhLckYb77El37ZLNqnK
1WTYl+4RJlAzBZfhDQKeNFdhTvnOZEHdtbFNJ36HPpOrO7JSX6lPgNpX0VhNe6hU
ps0XffNpEcdE6sItK8a1s6iqRRryuI46F/L2eofBd3m2Zdvwi2NICJ0bJ2S+X6GK
AriYRA+NofVKWNPHShsV9ouZA+I+ZCLg9j+C+bpZDzFN7W06/9LHEa1KxIya9XUs
OAnghKgaljV9a/ok55axwX8hpRbNPW2/FknCu/Elxq1Op0Gpjw82cZEBfztwed1B
pR1akkSuxI9fCWT15FvthZOw/qlo0M/LPWvzW2A4eaSrLYHXKWC9ZUoFwl3c4Dz1
+vL9TGVYufW5zqn/rwvDy9Sal3ZKgWlE+Ayjzmjp744XyMNUHAVSLjHcn0uOm+hM
03zTLrBLP7HOpMtjnEGRpJ3i+gGnvxPScVSSlNU/wvPNdZSmcBckbxeK/1SffH8L
4UoY/IY0mm43OS0CGqlNvjbn2Ks1fEQtziJZg+41CEWN4j4W1vgmCg+wkYXDx4sj
RpWFOHcbWkKOY4ktYLP4EDwqdtDx+i7o57T1R9tddArZdqAjnc2eFS/NtN1PgsR0
pvflFndoifCHUYJCNabQyRjdZSbeqRLbUgeSzOBHruxbJVYHzNAGuee0Bdzav8GC
q4aKauiy25+ESU+zI/xreP5Ohd/svhE3v85kqrDv3eSJ0nxcnXnGFUBBUzRR4QRT
MDm19hZ8dEuKdKkw5vJ+Fp1VLgunRji19Tw3tec7EBw5A34YSXg9clEdk3BNO3Hc
X2VWKkx97Zll4CdUw1bIUcWPRBX/qjSokzkVwhAZ1fNsPiFEoH9is0lVBQSmgpED
gYdHe75dWN4hmLvWu6k8Bp1ellRqxmKDe6qPyiib6zxnVRLFwnWRnm9kPrGh5+1x
YIcdSozlJ9ijC6Vai9wE/WWIkwnNZ5Q5pP4FwfFQsut7yEKeGz9HMF0PYhcgUUaT
GAbkZfXAkLO/c6GeY/fleBQjEl5LpTDYiIIntGDO2mQ2TGP8iW3R6cKN3oDLKXdf
a4e1pvnkwEVp6Dn3KT5AazpOnAkYo9PC/1F3b/0rlC7GvlUzOEyRmWHH9tqbBNlZ
M5cVzNJtRhwO1aAAGcit+VsKb3oKv4SAe5ZqJrAbIGL+kTOZbvKX1FkO8SHmUz9R
E17z4O5vSvFhA7rsnS4wUxAQVXZwyDGrt4ilpKEyJpDdhYdFeWwZktZTf3dKS6Ih
5RIxeA9SS06zNvDIrCK6hawO2k4BtYhdk+IqAMViXXM9nZx0LxzaAqcNjyN09jKZ
QSmIjHBIUm1aF+AYtiDIBTaN/PK7O8Lg1L0f/YT68xEoORCDZYn3/GRSj34gT5AR
2c5MeGxhhj86DhsmsspDspsMxWVLF2rkcYFFbTho28AVJqjkpmxsuN5daB1n+6jZ
/HQv99xpaIJK9WTuKMw6KRyHFKMRjXFphz7omeH3BFz8oxb0gUdwTYruc31fC91b
ygaNVX5hkWA3gGz8r1I8q56vly+/xYiuHO9sld35DYXjxTOTD2+fTW+hiaXujloi
k9Ub+BFW7O0DoEW/1FNTCdbpLcGxmGdgCkjlhFj0ZdAupgHlSH7d3qlklxm0Pc9x
nlHMdoXLnJ8RENbjv2fizR2GiNPkD27ql+k4eJWf0sq0XenfKAokW+HAQLIMToHh
ZL78x1IaNJcY0vSmfYf8tgUw27Hlb+jrvCYJ9Fz4oH2zGCD3GlqAsvPLyYsbVMdi
vvexGgbnRqqugHxZEvAS+sh4HRuy22kHh1mNINKYw3PmVKL1k8Iq+7RFiBBXBwNn
TWdgXYlZZhTBpLVZvTdRVr6Y8ss0x2dN5lSGf12jVWcCg3YEJsrd8VFA96sjwI71
vMOmB8XqIFzvqymaiTUKb3KBC1OB7krPwoeeo0cK1tC+hYL9Yj67Eiot8BT+nbgK
CnTe91cTOq2k568+TG6zS1S7WsnP36CQEfixk8UifahpVqqBzdUQgSPHBL5C1kcZ
QuDB0xahAZPWusp0XRDCcRc9BSb8Wq8qFre4/iTz9Wqros6Yk6Yc3HO/5Dl7pDUn
Dm6Vuhz7DCFyUycGA3At7ikIKbF2JDVhhlIZlT6UTKRfcAtnTJu/Ej2EiLT97Lhp
oSEP/TAbjgsMnpYX5brQxOiiG7zIKYlEZJqF3PLcMsPYR/MfxG3b6dLltop6jNTX
uPa44W/YwNt6MAOjpFpWe7mISTZtIkJBik7SsMycwoVdLgHQqA0Pni04IU2Uvjku
f+ErXGE0OicZDy31de0qZbwsctoYNCBZAllwI4b044nR2yQaVTFmcp3+aU6XdyM0
/UIwdgpFy2duQmsWIIirpx6VuEJncJu7+ccaiZcr/hrzdqPJYJvrkhzY/bAg8rtL
uJRzxGKpU/efeCqA56pRI9uQxW8AgadYi1oq3qH3sNRbp3dakOsOgBKacfFrB1SY
2/tk2K28wdnIzJhM3jPnOE982qG11zH8dn+lVix0CKJM+ZWxRsPEqIR5uC6vq/KD
EIK5um59ivSD7ql4M1Q6t/+xEUE3MKse09GcGCCJ0qcHirncKMQKcoNoY+Ox+Hm4
4XOqux4VD1MlBUDIDdinrfrEdGeetkPsexK0BV7dUaaYItW/MFhX+khVCsKIwwAT
hw4m/s0AmTDItD5lpKIP47tOYF6jd+zD6FFJqPIeFoDZcR1qMH+V9oaAIQJ9pB4H
9JkCzUG1akalU+Ait9Yobdvl7nDO33kVqVp5SHeuoLlFO5WpoTgvzil8Hb3wmPzT
9r3i/wDUh1f8lzPUcNgM9IqYUoJiv3+yLpL82XspaNbgWCcn1OnVpKI3UHzEsWgE
Oy4AeAyYNpac7bU0MG0brMM3eGdRwBvFC3Eh0kC9Y/ms0TdkAhIi+sBK4MjlYM1D
L/jWIGpZgWjZsl2ggYilki/qsHDmqZbTb4SooWwO+KL8MyvPYlTwTtikRFpTgS6b
fpAgNbc2egrgNt6coY80LWPixBtMjM20vrA6dV2DAviSaXzqbgD1U17nxO80AKFF
PQ4Qbh7G5t8QDhBvFNCByr0NGrSFcR6td2dc6SfZ27LdxtKBObhYcEkj3VHiptdB
/wVztHruR6E8keEmXIJhiIcOL9sIojkk6ATNfUF9h201IL8rCfa3tQNtaaIhaK+A
AuDUFT19wshtWkE9gnymQfBT6QbeJaqRJxd5JDrYbYDYd/bUdJNawUOqdCvkBy4J
m5+th9sp+7rep0ZzwQep1d2vrTnwk8P5CG1uNct5eedjfS+tUJrcFqjuMfyJkKih
tiP/AglVopKIzDQZ8dtDTZ9HYG8cVRUK3A8dXymxraua7j3bII0pBmDSXzpSIxXC
CyEDS4XmxiPNgliGFCeQiUcOKxHBQA+xgqil4WFUarYWC/vZlI7jvFLm1LOtOMMZ
IfjuCM4VuOuvR/LFLt3RgyTlK1hT4TQ+CkF7t5ehwX06vwQQSUq+7FTasYEAj4ir
mLcBc+ejmKgc3TJeIF0Bi4kGLDEtNpRx6b+S75OnB+o3AiOnk3r3ry9V+z6UzHp2
iR2W9S4Avt6vadBvTmGFlmHPTKrXjTZi9sI3VBTWZHA34CVH7OyE5L3Awy9yedDk
YMoGgwV0Q9eNxh74c5peXW69/HrTLLBx96sBdgg6d/CXOjcxT5S8KjL70k6GzIVn
h7yE7r3Wd2OocyBetENDRPzOGjW5GiPmI3b2r4Xx6zoK89YeGxi4hEGf5DpEQsUF
bip2ERecn/Au7LrsesRPBKwlNCjtC2LgCiAg/v1AZfqbRGBbmyFUu1cYJ8RwMXMy
8ATwy7ftGghJ7Y9F/9twmUFLKdPgWIdbAcnLtuqUQYv67WeKsWqTFHojTLR6QMCN
62HbvyWxH+8RNOMpM/JotRFVxbtV58tuaHJyDfua8zkRwKWkToY9e0pt4UbNiCdg
QRimT+J8pxZZ8etpJkjLjVUoKG1PhbRqXgDKRSFAPvTy/SONsbqdVuDptDPl4RcE
5TQwrgq/v2p67xsaOa6XeH/doj+HZxOxS9XXLcuLLLV3Hq+4KmiRSZ5K2U562aGv
0m5SxFQjdI5U+6DLjxsj08pWWuPuqwY88EOSWvRU4Dp4Z+38ZtpP0hZsR3lJbXuj
q9HYgNLV+YoA/9f67QrxtxfRydLg69IVK6Q297XMv4F4ykOsus/mTod4fS5PmaSe
lotCL/OEFlVLs7KXj9rL+JhvaejQYLRr+RCkRPEs9ZYCebmh7LN586ZPIjJBPEOl
iTO0AnI3uDhWxwjA1wYr5QswxgooUsQpHMGJNHbov5EkbbbTCWKr3k652gLYm9OB
xTQVOK8ViE7AM15BKqFcL5dsQ6S8ZtJ1N42V7mrErcdiMnRg5n7vVkYx9mo1M91U
3kSu4gPAx1xrmay2pwFwAq9HqaA7vOezjULMM9E7y4NUgWHNUf+GpgJydx1w6Ch4
jRQRJsKSk3EjWSVGwvtR8qAE5b5rCuMQvINqK2YeELQqPPtLu6hltbOldbdNjgZN
ZBk2PTPI9pCNy5PA6Kf7Osd1vX2mCn8K2Jyj2esBTO1lpIYRgGL3eB7mGcWvtTvA
hoKgeWNctc2aOe/dktiR22IUvz8qSC+4gm3+AXYuD7i8jPwYEjS1DALtTX5475KT
nsOkHwmz5cfiXulx1fiTYMYUw1shPRQNQ9QOemRzg1gQUGm0L4jvkzEpM+e4NsHz
MQ5e2J/5LUf48N7j3gttJ82rUKH7wOpTcedyS6y6immS/PgUKuXFWN81NEy4Q8I4
W4cbxVx/8FwDF2ETm0Kn3YJVNF8dh4+dWbLzJN9tOIJyaW02F/pCW++tE43M8hMO
AK1WSnRnozgGwS1QRxOb1R5EPaveQ9btujVnS9oYaJnPQXMiAOx2hQCkZ/dDXhN1
oijv5r7q7Y9xYlP9Ary+jHN5HtByfcchzjHXOiZEUA/O0EGM1dCREB8lraKcM7EL
9hl1bqiepT5yoyRVk9+OCFOX7W1/c7G19TMkhn+REnN+bZ+3gkPWu0gNIEMr+Vwv
ySYP/FhBBLTkdEpzD+Hr/FvVxKdNpEeIQAWM4/mWLNMweR1ioV91i10BT/L07hww
uPTwIf+An+ipts0HNRH3qnTO1NyKUx223rhkCpLuzGEx1tMs2E7wGQjIspvlxHg5
NdYKEPT3xPv5ge8ucQIMT1M1yPL+X/DzdqmmSg/Q2FdKGbWaeBJA64xHVKjC8nP4
O6yrYpAAox5Mro7/K0kQTmXLycVYnzclxfDV5eiXQL59lFOKJoD5YpIm4ch6IVWR
STijXPW97nkwhGHvK5WHJWCkHzgQm4uTeCqfe5WpjPmVT1OqjFmyifUp30e4AE+F
1uNndf3YPqtZUQbfIn88qPiwoLkEmsU1biyd4FWhWkbf3ziDJLC/cyWSbYxp007J
IyCynOma0VrXmkoBSYxHkO1VQIGP3ZIdTZcvvP6JAEDCXl7UYEzFxzJ33fnoTvw8
TuPaGUgsQJuz5+SmPcTDqJ0RMieMf13hM1PStcRWxViV4xkdoceXzu5ipTaCb/FE
adHKps857g5qrxaqDew+WZwSQsEekjAibFZ208qG3FRM+0aOdxicua+gvfAWdtLx
xcoKBgzEnxXDKicZtmv63a+p372MnlGBULiCHNYXd5PpEf+dE4PqlwnmjbiwC6kc
mUaatYJzb4tITbOxHBzoniQx7p6Heys+hfdy6eoIAYRTj0qsdB536diNCj3HOWmm
ha5kPuN+RI1Ug0A1GyJtKt/O6JFnWD9P5Kt2rv9n+JYL8Bpv5tg8y7r6SL99GL27
uwGbb5oCe9JSsmE1C4ENufGl7H4BIJHuYV5CZYp5kITvRdgAnbAbgpWYHLcN8CSP
Ukh6DeiVr4w8Q0SBKEaRdns5qqN3+YKNEcuHIkn2rR2DGH0EN2g0jMQzcNZF9Q54
Mw4exjhioN1Co3s8G/zyblxIJ7e3X5ZF1LY6hXKNCpEJZ8noQ/tj2FBl2PFfxSm+
7rekRO/riX9hjKYxJaorP+i52BcH1dXosbMbI1I3sgXA2NEuT6XesxFClFSwIbYF
wOWl+YVL6hJwpBfZPpvlKAOY2jOtTmrpv3r1fP3BFkIWusb2TYBqvkx+KMJgWzJ9
u89XAUZl+Ai8uZLq0NHoil/ATCh5Gi6lbrJx5y7N+dY6d8yJIxx5YlaXW0uTkv0Q
/qwwLj65r86T7sZGR4liOv9169jV2X3mJH2fn5eJ71LVBfOZM/wbYe6oTYdHL7B1
/jPTD+ctwN+wOm8H3ceE7WJipbJHxnKmFBVaiIb5zF5UWdLLTxEEjqcDnKa1D/1w
81DHaFavKEQ8nmp05OGtBD6XMiWvIrRXq+SF8znAiBqoYTMgYRj11ZGa10CkyTgh
Pu2TB/tjgHMW/nqdkLZH3INSKpUIqvPotpLJcZ9XEF+izMIqW6zmGMTS/+JYhk/u
YWJlWmQbkoSflO38unvbOqB74RoDFyv+IwaBpAT7NxdIQL1ZaIKLlL5SBqqkISWp
XsS/PZBfh7MPOK4eD9tSMp12Ux85og2TNGhraHcEgPvLsCiSM6ySn2XQHbfs+OY8
rJ2zCBFH7naxK8CsdgAhXR2yi403Nq09tgVkCiCGJovTtaS0+gNhF0+Mq8CGOAL/
vuqiTdu1pIY8FY50qc73jtI8nQNcXjnbmNB1bmqSbNCcYJ0kQzRBEs58p1Hdp8aD
w6a+psctAXW0Gu9cedSE1HJdLnbOOB1WyfYaiDxPMCBjCAGinum69APzNyrH+hIa
sOAYVayT+K15W2jpB63osNZ0POOqJGQLv/MydG1iBZ93WHU61AlhT6+fAhdv0IUi
NShBj3Fa77VRg6InxlkPNhhzkqTXL0cPdVQr2OVCIaWawKDAFj4GzE/HNI+01WcH
RVWrHjIXmjnLNOV6N1Pf63wSJyh51x7weTY5x8TMYfNl0mKKfUaV3wP3arcB2ce6
jeP/IfHe2/03UH/HNf3r7kqXV2mp8G8cr89CiY8+lqwrO34yxan61mQwQ94hKe1O
UmUESU0lpcWjr4z3r2UAwTVah7Ao7GUKOyE05zna3fzCArpM4qd769iZmuowdN0D
CMStsmOp/ykyIJzxGcueFhQyL8oj1jXKLI+FHAwZQclXfo1tGA+lrrvuv4QddMIY
nGTodckZk1hRPqZyMwpkr4V9kvOlUFtqHzAwEUWDuENISCF3KDWvQIpqVptYNSbK
Tq97Q8RZ3wdTmOzpDPVluQ0S62J2O2DpTAt9ZwPhIt3fDZDQpM13oSYadqr4SZPG
8YrDPCrGQ+Cfq5JjWglXAWzs29Q2sUkZm0BwifQpmzFv3NIlRcwvZBMVyTwkeLpH
Zduyw2/ZOauqyDgU1KQRDdhi+WUsIH1J670IG74q0cul471gGltLdut0kLPv2QUX
93A6limzNiydGHN6n/nt/KX00BqoAr0HET4D5aXJGv+BO91H9K7maxs7oCbhvS1i
f0JK+/sVY8w3LTjC6rQYzt/u6vQjL0ZMF+MXYF4kqmlOj0cgDJDFuzbaYOP5nSX3
vRDWOwkKQVZnFUcc5oS/3Dcae4kNDd8UzgIr/NzZHXLptQqcxvbzoaZJMuqaLNMs
jYxfW3ETm02Me/Wttdq3RaSmDrhjoU/E9/GZXJe6ECXq6s+SJODk/++zoN8jnRb9
sEjTei39S/D6i3rcE1qO1seeNBHu3GyZP/fEnvWR4ahtZUJWcKp76yDnBfI7YspL
wk/ze8xQ0LHmZf4aUQRsgc8ykrH9q7AJWwperoB69RU/iS9pwc7UIhEd3VrA8udO
fvfjzXKGLrlQTz/mHvMrCnMCtTMlpFOqAHdFQACTOKgaurPsePFLv4HFuWiJV4Ud
jVGGru8WekH4gZXEWoe5dRmnsliCg7apBeuT/F4rjZH8nfXYb4CjftXrcwX6aQPN
10bVYSnnYxt2n07hWAIn/rnwDIdchdaYDHBnePaatxbZY1bQkTJCAp5x7cCmLD4D
uI5rgx/jXqU1bA6532IERAk5QXGvF9LErKT/1qosY1tQxki3h9hECWsPRQ3BcFLp
kDx7V7eVPRVzHdPrMfWgZniy9ANRann+GIEspYAM8ozEtCFfymy2WzIGr78HEqQT
GeAcb1t/fKUe6jsL9CNej1q9aMSo2JeclXkMc6o1/YZHssthblyOPn8lU4wpw6x4
dAissouLIA5y/JD2tBqwIFi6W8bjUB3XdUVar86uSJWZZK+o7AOi3JoUjB/E1362
PspwkJte43qwJDPFGsiZQjl20ZJJAFqXIpcwOMOZOxT/xptjR/AIBqvQ9GpdTMv8
YO28PfRZS4lBkYy1l+uqRiLXew09yyUbMosPvU0tsItxsIn7cDtX4hygEQxt8mNa
mnEbC0nbZWfgMpIz+hzlkB4hk3lvdOCTWkuWgLVYc5E+pLGOixQgzVwqs6c0j3UG
yjOWVn5JNjthmI+ey03zA95GDjcKy1YfJic74QOpdsku3A/DgCwlFx3eLRg3K0J1
8Bx4ZKKLQwCIRSwwL3lb1VfYkidCDXU+OWHVjNCGWnVgB1Neclb2FcDPLpftHA8c
hLxMZCDZtRSeUiOl+q+SQgN7jsNp1JeXJQXJaBMYOyCyPRZc5t67MmSdNk6sWI95
P6KRo694Uq1KZu5qZwuP6J2o9ceobwllw0HU9KIIJka8oqXIXQ/cYvqodFpVqSJI
ZDHGohQA6LSfvFUnPXWTlYtJtFZetZSHQA/RUtAYoyG1lc/rhT51tJ8h2Rm8q60S
lQqbodt7iamnVdj/9Y6j0iJhC0R9WM4XfPo/H8mQDnAKoQwtSWvviMbGQVc0/l0V
GV3QqDRgvB/ocWy2Jc6YEMWCie1x8XV1PIkTTP4OwUTItPXPZNn8800tXoctdPch
B83l6PYx6JGWFyVzltJ7dULfFkKI76COfW6r9ol1JkhYiknDcHjPu5jX6tyPm3Po
8Ish9ojO2ny/jhiQABwhOJJtFV7EcN/1cV/POMnzKKnMDhQzT2FBt666v4RIGmFL
q8U3jXtfdPyNMiOjT7wx3dckR2q52Pxl60aXYpF163rEgnK6v8dQwii6yBuTrUFT
tBFmIGvFIdtt60COW5Pb2yUJFU4LvLsC4DO9LAGwDgXPCom7rMhqKUbnnIGDqPgL
A9s26tnU27Q+BDQW0JLeqZ7c65UpWKJteqjMi2MKpjkrmLIWdwhZ+up3+/gKyEXV
htom9z0SWJwBi5AXBT5+UfSDqqQZiWPPvShaum+qWPO/LYGrALwyETTNwliwwXQ1
2bd+wiSfh3bvf7FEAQ44BrHgD+6d65k0BvvzDememvU8tlhClEcDDER6ptDfyE7P
jGIJPYbDY1PfvXVEJDbLDgNZNIviq0IccujGfY+Mn08yjIUJJSPsCqmhes7OCTnz
SEdmNmJB24kNCcPQ8jZ0erB++mdNr5uwld53PkElKkXPKA/pxngKnj1r841gp67B
vS5Wj9uOaYJebM/HSiJ6w44VtOo4HW3UUXuRoG4/AWrMpdndUSRO/IydGOqrXu+p
UStv1zcHFVXKNRv5tp9+OWU0D6CR5BDbK11WmJefLs+xTZdSmdgyj4RrVh/LTlxZ
4+/T6uvQHHB8l7+atRn9fOf2Q/7iegVf8DSDyuJ8aXBNs1S2M+Cf/Fk+p4n/iVF/
j2l7FZVYgV/hC2luWFTSVgsWFGw+64NVRMNBPOQm0mPVTVimB3yO+RuyZ3yg4SC+
XCmBxOahUs0PBxWpsEWtTh/DbAlzIT/7HvbdvZ8MHxODqEfi68jCaVvWAt5AzDbH
lsyuLkdSDuSQFurYrZ0wWUE1Om+N/dhlCCedZO9rUrzZkbhMx/v+NebxZCrVzE6l
tjdwxcoBiUU+NfIEH9IRspXSa7Nn5qYEzzqFPjkBRBZlVjOm3ocRn1Kx6G+X2zt+
i+bQXgH5rKlYBBBXyUtT2rSjQrSBnE+rqKHBN9f1YYlfXhH3My3qcpCBoRFLjK6q
+J6Ga84BS5cDBzoFfGkrpY9uYTUR6FjBqCeuMtJh1jpMfrXJcpMDd5oURjk02DAc
4yILD4DhcaTRd8umCJ7JkaPE/gmDo3IbRdYYcjmn0zG9PMeNFyvrMXDwv4g0x4QX
4oyKbyuVe86jTj2bbxBCgZxcpaHKQ3pbhpnFx87NICmt6atURYFPKV8wnLd8hFdu
BndEiSZFFWPSTWr6F5xhuxkcPyHwjyuVpWW4Ro8eWFsXj+2wFuUSB8Jq0lnTcpE1
tCdwLjvvjHvmcpxj+fK8P6dCAPfN1WKoJCDZE1rI5ny7R24l5zkbiMq2IM3Lk8P3
4NruVeMuDqM7/MxcJDPgUztEi2ROXZZUTyHJVhZUJSpMYjlafPwzYGeHVwQnYNj2
4HLMot5IjytFSdmnQ00TOYFcW39fnsg08AqatORhhAAJUw7FePgOiXNkdnNfIrwR
G500tAiNOgXSmMZlimgTIcSz7/IjSyeApRhT/Ol6R3cEoVPLfLAEqUQM/UjgxOEx
oR50ci4zI2ad2qsydLCpJ9SEmxfH8dwJED/xuE1kWnTCPnWCrIjjVnlSnWbTJ2gU
Is+UbiRqz7vdUNxEf9wNnIxmd+pYLhYZsK9ODWZ1ZdAJzfLXiKcgUL5gt4tvSDxp
npw4UFfkD9BV2zHBVI7bespaFBtz49V7aoHO5keadm4q4Xl4aGupcNIrHYQPPIXX
KTyRGkINznJSFtdEvTwiZpoo9RJvoZfh4B+zzr7Z4/dA/zEJyqiGEJBc9Cpmh6Ei
WgGD53lfj7sonttPYdRwR5YMieCgSipha4Dy4alqeeg3YiOvmT9WIJl3bZzsxigU
PN0YbqpsC3pb9T2s4B+5HTjta+1dk6u7dbJi63mwsczuJx3djX9poBSzOUhliob8
Nse81HsdUG5m43/2xArL95SJoXn/YhIir9qx1eh1dcVw75KRZY5gAguzbW5lFUsS
4BFJFDzhxhIDaBXpgRJDg8luGX0j6Q21Lx2+sppg6HYq0/nw8oppksZkPeXl/y0Y
e/w0m3DaFYajBgksdKHOYvOyOSvogY9YWBuxio7+HuqRnlFZ8IhFy5Tj1V67VHyC
w1d+dR92HoYxhMU37ab7VoehT4QCxbOpJhlyvJQc2ErRNVfzSX4KMV1yGf/Bg9AY
xwB31N7DZPbX68q4EKXEOzJjuZVlcDrWNofqWmi0zr/NYLpSCizhQeQPq3IvfFTn
/Rnyfgh8yE90w+E75F49k5NhNHR0DGWDhtk5LmoZWKpisc2JnJDzSn/JyMg/y4Pn
MoImKc+pA6mteDLOCnk0Mw7BQSIJBgCXDYugtcbiK/8/GwXPq0BqoQWzhEbjQYOd
Hh+efkuWARCIrmoDBVcpp66eAtzp4kX2LF8mzOcmUaWdGyc50cfK/1Usur3UmmW3
noS9zCF9VB0QamzAJv9NYGg0N7to8pNK313ltTO/OoKKne4YAQy35f+MWCSIeHse
eV0Xs06EGwTu9DcT0iaPuRGNtYLYFLoK1Sz1mdV4RKoPo8dFA56mgjFkdYweheW5
ZzAoGkNPdVypCdrC0HTaD7T7+4e0XhP+vRqhApbBJu5jL8bEUNX/58/GI2p5EOcX
AQddkwoUaaYVF0NK8hZ8XDHvZw8h1+ZC3VAIsJU8Ke5/x3QCRcG+NUstWXy7+flO
+0amzSVX4ejR6O28NMzxuLcqK7r76Ex0FCDSwzGnLsvZ1m92ZidzD0yah1e+W7v0
Wq1DONtG71ojmX9pNgO/zOGAeLvBQl2+dt2M2tr4ZNxysWSoFrYLXi+jyQR5dc+v
arMThU/o0beM4u+KpFk/R4iXMxhE4o4p+lSzl5/u+wqXFoStzPuWxMEo8u89hyLN
yQ/XkKXLLk+IJ3t6LqoZyQDE4R9e3vf6kvutJjXW3ANnQuAf3hQg/BB5JVgR629L
VHv9iFvZS1xsXXluevpijMnPjJ0XA3L6I5fhRENBKHwunbsYprYoEn+iVMPly03p
pkpEPdnVhEB2pkXByKoCARPA+RDVzXLEOQJKFBiJdJ/aVauthJ1Yv6r0uj/hicEj
rEHzKObOfDaSIFRm2NS/+HSHBtudw93y2eXgk3w2E06cppHn23vPeY/f+0V1/aFv
5SIMn0+FyRESVap6rL3H/pXHxNF9YMQj7dU4UWUd9uP3L57WpZqCuKuxBzmroDF+
ZMWlGqWFwWhnN43czWoT3Uo0RIgSeDTPKbcg6AWTv2Ix40SQ1405XsmLzACHgHPs
Fi6GmdWefWUWe1nxg/hO6fjQLTMIaIt8jcAA2ieql6FVCAtI5+ulQwtCg/FTEK1F
iPzJ7rBO/IcDJCOQQQOx0n4A5glAOs+amE1BxplHnBeeJdCyUcfvNfTUaa2HqeeX
nnK/6HJBPtCl8vMESC4qsfeCFZlI45rndydJWU6pm9NljnuPcT/Cxe6itGLwzTSc
k/LINq22Vw407/hKHP1uWCQ1HX83e8glfVgE3foq9V+XFgIVLlWfDZQ+4LYrZN4m
uvBw+AzQcNXDuhZNjJSALLmh6qMqBXPrR0e8JoqpLSDEGQZr0E/XuNb8V5W0SJMW
QaZMGgmFPoywzvuYgmpNjnSFAqf6PTR632f5ZodPkicyVWBgdlXAd0Axu/sersDM
oL+YJeFA7/MGku8kJK4lYYPoXD0zj+tuf2+bAYKLwiE60UHRU27tnJydvIGSbM9m
1y+fYsXlTak7qmSd3SbkjLOS4zH/vTg47L31FiKZl+biGLEj0ow7groMinPek5m6
3CWNSVmbnqglHpFturk3DTjQR1xP9RoNQQ1+l1byco4ITzanevqkBojasyCvV4cC
PuCvJLQY/hmrla3KUHt8wXbolyGTSkkMMn3Ym3ljyLzjW8DGGT60tw7GMKB0Vl23
ct0HJXbRMoKGX+fzXv8/A7EcTegLmjHMZJfyTs2TUg3Y6aNItai/ELmNRnvvxyL5
bEIOBQcq272B0zwGF2FrMV3cTpsC/5QJc5On21Azou7UGLzug567qdgjOuT07uvU
shkNfH4iquHmYbDi1eUZvUYP3wCXYhmIkpCVKn7V6xY1fZ1f3jcRNSJ40w+RS4HU
VjHMF7IRQvyYywaQrWEExM/XfQleo8KRFEiX+tK5gPoBJlPTLF6nheg8dQTq2Df8
HMXiE/3IjU4388H9BpP55KpFHsJ5mZ9iJQUrS8I/Wt+HsfVvcMP/PiDm0C3HuJTS
53QSF+kt/m3mYsej2dcW0QOy18q0YkIlP0B1kYjeeMVmA5wlLKpG62PzqgWP6q2N
Dzct7xiH0gceA5Tvxapj08RFZdokZMfA66jGZySXp4K7IEGHeCOwu7/90Etsw0Cj
vugxkdIsYW1hYrKHGcLiyxfKustx+l5yajxS7ok5Y+aZiFpFtwkzx1l/neAyrBvv
LK+Vo8CksioN5lBPTWq8/32zRNHQv9UBomiK1vgTk1EBOVDmoJhIh0OZZU8Uqqjf
JAEQs0Xc00Ui2Qcsx8X5NwzkyBX8Bgg3eIzejRZlsqQ5S7njHfsqmWCckOxO22LI
1Zr3iQUBWSe+OVGFakiMxylnonvSjYe4ugcfRbrJhP2eW86LAMM/dNAVSXnh6kUA
BM6sykMUSs0UtF9YIoMSI4e4gO4yjQ0Ex6RitquGWrpHmGVWUI9TaiyLy8of9Y99
XOuAmqV8q/ciXQYi7AkYz8MORUESnrcYklJi8Aam6VaY+z4IVu2robiAD5K1G25z
03HWc0aFw18DtcXDzBziPDCB+nhs7dDzYFs7kX/U4REtTv0szPkCuVym3/w2yPV2
nfGgDaFvcT8vxRf1u2ed4JPdMo5Url/npqiURCEeTSlqyVoHm+22DAgrJSkSZD6K
SXSXZ09wpncuaWVQQJKKHSg0X3Hk2GHHH8IG4DkFlEKoVq3L7JxgR0kGgn7KExYj
EaJMtFvDQovz6g1qJWvgabM8xCaem/Fjcm475WXQD7JAOnRJR+24+46mnMsO3Yt9
zrkoozhXZfxdbuAew/EbD1YB8whZDmtrQAlz/WDjrORA23ca9Imc0QCLlK2XuMxA
J2SD2VYnftkD53LEVhBGHvAxSGFyZkUeb4BpamOUSrERH9PnAwt8g41ZLJupEP9f
db6A58LKct45Q1Pqw7XpVQfKzQO/DAwG3p+tU6G8rJzJgorgMiKrnNwI6F06AI0i
ttxzocpk9xAC2pQeYjJLM1ATcYX8iLLPhON1+YxJO5xvRXLkiJqoO5KsHgAJL8ML
hmXOIFv217FP0HL+I+LJTvy95Zmz4/uJs/hiHSqP92qN1JxcGbGvlRYAi2+BmP3Q
iv6Gsnx6Q6821nqYEgKXbjlmJQTfiE6vT5vIHtrfLduGV/gC0sZY2GrL9Ovq0wuq
OUYr7/7kPIePyL6ErM/O/5qKyOnywACSS6q/0fBDNNWg7URSDw9AQGQBupLKRxar
A6ePgedQKPCWSOfd2ldhc7K5RjmU7r0pmqp1rLXbg279AzNlXaRNF5xwKSVh1CZ+
K9+snOiQ5ZYE26ZWfhhao8tGBhN0Xcq0Auauu8OepkniXXrKIFhvKLYE7omx2zvp
XVEJ7hmAiDFsY6zkD6210O58DYj9AAy+mbv2SWFjGKlUERJ/mK+kXNKDFc79rTcs
UIp+6wX10a05nuURgaUxYjkpfPbo0lmKuwZScp1AQ94r9abX5tY0OehFoCpfktIB
pM32VR6UwPc3pMYE8GUg1efl0Z6ljwWV7Cj57g5Db8UxLgLEEdVqnzQ0cJjAsKJ8
X31gobaD+G+0U547QodIMseJZD3EZMIVzXL2+KNjFEesD11bX94Nnpzi7CNelbOW
rNXdl+kA7tBeZTdeZRNYcKwc1/x0MiCr1oGWaVbI5Q/Vc6+TB9fqLI2YgnHUuFEN
1nCFTZ8wbjExIMxW5vGgB9K5IdsoWoyumAbv8AtG7roVF62dQtaapXkDGsyTi/cI
dYU0E60SQIZr2i6m1Mo4oLCraCxTSjftZAaECk9reNhAd7aH12PMK94FSAAF8cN2
pzq71bmFLfHemSQiY3Ki2hWbbHV9c69vn2OGP5kX6LeDM2NDiRqfRMrAeU+ZuTJ1
Z6lS+in0aQOnGZkm5+7jI9EY8em7HIMAz/qhMki8AWYCEvwXpnyNsJ7nOZ+2tLuq
9lWGWJYFCjprh9RXMMv7vKoBmTivNviOmC9wtTnhbtDVwxVWG68amwfV9W7eprAl
6nQLIlZSuOtzuzYjT8sSj0aIa/6XCzHtcrWJAWIqFZvkRKq9Uo15e7k3VTRtRq5C
zpeHIS5p6UYAodCKLZGwrbMbRdRmF2WLB4j7L4c+yJhgaqaO5AjDoXiV2wxMnmKm
oACfQ0p/kYMQfWOOSQsJKvDO4OJFRZDGv6OBClBbNdpjKrxdX98cNkGA3jkucGQO
qB8Jng9BFfavx2tjnuKw06DqAbA3uifnzzRU7F+eVFcEfsjC3me7RmbCaKyaccYG
kvicVxzqF+TopPGGPr8IeL4UTlQNrbku8uc5lTZ4dAoqYqHnDwLROooIHabaNQ8W
ebACbQrsgCMFFnNmfcpSBqux/q6bGrHtKYC76plttgSWY7KMKyMAz9Lwj6uCV0FR
Jcol+CmuzpXrAq2vlOeyP/oZZXtFkCUXKAqhwPyaVy+rlamDytjLdRtSTm1MOp9A
Xm+q84neMcYkoLxlZLQN94un0NL3aeClVIexYbDOj9rB+jZNKzFfT49DxyQBeJGz
ZRoHW+nOdBY/PyH5UF30jiE9HVa3RMQ/DVeEzReCY7PedkQEnppWJ3SuqatNztZ+
sSVm9lvA/hCD/IgWUGr2AzUszvfpGyrWfigE2nQIvXfopBRBT/a9CMOe47uga63w
FSfZByOztCH9KGtBXBUovq4OCHuZ0LIA91EmifGRfFKIdTlOL3NOyGgeGWgGR8PJ
dnO7fBeT1ziXaykqbYkObjiYa7K8dDh6xNcdhZgHDIX5iXrOwbrJ2PUF+v5zcB4U
FFDaPhsIMfzzTrqB1LC/SzAkl5W6ou9CEmhixI6ufY5VCYOirmrLvRx6u2hGvVik
FRvXTUiBbM7PK74f/EoksrIgph/44+Po+nJm2V/UlSbBXk3jX4Ic+uAfn4YKikYv
M3ZDQch7T0v9tozTvLtc8Jlwoq1VtDiFTyU+OKH/ltIi5+4GJhBb9oHkSy1YsRg1
q4p4UfRu7QawRJcDLjV3eHUpKcFxY/1o+Dir7VGdykAPE5o0OIFMSje+aaoaUaxJ
kiIe0Ccd9CZUfw9n2vM5DlXRFZ0GDcaXbsvI7fExb8GtaVDZy0iaLFvDDdvxFPYV
KewViGmQf1w0G84FZczc83U7aNMXjaNqcf2DpdiG480GY3b8implcqUseok3Ctc1
Uo6rXDJs4djD9U9KE68MZATThQEiCgGn81UwVhrzvRg3rGlfVh1uxhb85FackKWN
zZcfSTwKtRSoVQL/mLvxAjhSQsiGnwf6fSr0bPEBnguzn1XnwCQFr/xnp5KcoAXI
TcJm+MpiQ9+nAcefOlJQ1DIaM7pg96soV2r6Ce29ywBLMNzVP9A5JP70sDfwwpOK
fbUDhYiewPBt4Uu6gmxbFcVV+yWnCCqPYtm1N07/o2Xu/Lnje4/YCqeC8QEvIEZ+
jSZ6tB4zrySDn3xe4SPqi+uHRW1KpcGfTyWi+y23WMLMdeHBEWhuSvrGC7BiMxlW
CvXEdQZGBobwUrMXQeS4LIpVcpAS5qDzMD3oVYlGUiDvEgjCjPGkjlqlX+OXdiN6
zET0pIjT9O09GUdE+cDh53bN8VXAZWk/qVK1vdcNBCy0kyqX8ybaXU6ckYHZn67F
3HE1awsuZh2eKhSwrCGoPisj/tyFA1QxY/DznEmE5lKDd+gAjzicO+FueWCEvIaD
upFR0EgKsLoks2jG6c2bRVoHZgLW49EeFxeaeJEWH4OwSC+II3Ds4ymfUZOF0zuS
8rw2Yp/5rXzJsAgH5dC5QcKGG+e5+AnATICwla+1WLsf7JMYO0/eoRSu4lFjHy0N
SoPTqiWIeJEnRNWgcj2bjhOfAxLCQsmUV+PXH0BbbgTIxMBSjQwVUf4SjvMgo1T8
ESpVkd37HP/HxiukTI2TEUS+eIqrpktlMYKJnt/mXrT75WTqNtJXyh3YirTMaoS6
pjaCLas73OZDQWLBpbgkt7+0ZZk2EvxxrFC2BwfsJR5SRnphc10Th8jyElQi0lj2
gH9r8iMQ2UNGKYCj6mr1xmWDzUadAqpcFrnJiT4fb3X/TCMMqoQKr2w5FPnirU7r
/TlWMyCXNWS9ZSVljBnSLBD42RhuC6+iETppBmE9g1ScS22jltp5ZRSrKL0n/nz2
DHAN2bWhEvYyiLR/ifUqQLfrphhytuUAXp+Rp5Stgy+QNoYW11sICy7y3z7hR2lF
mtBE+aoElc7hu4MdBK9b6MnRIXi1DK9R+BYuiKgULxP/PGpDHe72OAKACq1o7wYF
tSa5CXe8uuWTdnzMcy372fy1eGVxOnTIS530lMEMND3wgypnBbL4HxkYYiE3QYio
Kh5J2b36C2oZs7KTZ+n8ghPfJn7OmHkmrRL9jwx5yGMRtk2z28AFK8dyXR80NLp/
xyMy0mMt9q09d3YZRlBsY4g+H9GsvgP9T19YtKm23JNmRXMyHHPwaxzw7EVb09HC
631jTy4JlfbuiSBotPzxTl9WEDPRRJ9Rm0KOIHfOGBOXLteOqkDdy0/Dfrx7RCH2
z3NDsAKsYkhW/cPUzYXcOsfYDDyxvov4cdsOKBHfaD+YqkLYq5xlyDVHJeky05gn
wJNI+wuD8G/6pZuHSV4T0Yf43dlGDNe0eWWz+ZtL0GKyfDBp1Th0VkTS6diLz6rv
FsPZWhfRA0oCRbZ0WXkSWlu/QIQq6t6JrT2t3PXX7d1gFDachs7+kgTWB4dw6xut
yEIuwUQNS1cpwZ28bNZsfuwKKtb1/9D3dPE8BuAzY9Bpzx1GB2hnWOxqI4+Pb29R
07iLCQLL1tJx3bgvMpuHjMaE0wvBeD1TLkXljX3qymOoF1YstMLEtgJcpha9ldj8
WlnW/4/pkXSccltZdtDze84oyYVvTizIFADoqcjVZZu9OPPVrQPIW5bzvfZ/TmU1
uI5K1cmJQ+Q2raokbXiMYShlV+VzovvqbGPo5Q1Mp5w0rhrhcz0ksio9Rh2qRQZ9
2TXTuRXMWcqzaS52PkWsQs8yQoIT5ioxPntgW5xImoz77GX5jOHkNdQrNLvsYGxd
Me3GeyPI4GNx3R/qH2wZngjwNdfpgUkMxVxmQpDNkYElI1vw3ypjo0JY5w12fpWI
QrJYBmvqF59wftIaVKul05zBCvjVF0pcAOvV6vlwnDKrOo/ZpnpbH1phsbhIImE0
PQznCUT0uznOfJ97/WW7FlMVJ24DqtCoG5fq52ZIH3RmVz0y3EPbd34eeiNik9ZM
op5tlHNjDSdy8DhwppJv47rrbBV2GT/Pl5I3SCJBmtes7o7bTudDVt606Zb9a2Xc
XoTIvGglr0DbznbE5sVmoTGjY9NBY4r/vacuHvq4aIjddzafa5lOlGF3WXS5bXvn
RnCK6brk1Yl3D5PzVW3yxwbvZ44QZwKLfKj0I63lNq2XYPfG6QcVcRQbErEHh/99
QfoGXJ6+qhNOMEeVByji8Is5x6aBDj6ss7MzJG7Ax2goIBzjkd+kZ3rvoZQGYhOQ
XbnO1dAnPv2cv5WZbljvP2nKYP5UYD5q7rOFDSRbtBD4mChT8HB4JkPcqWLQUGM7
KXbk+u39rKV8SReHPQRnvR7fTDu4kTyCwP9XR76+vBHkr+2bhVEAIj1jRfsal9Pp
Py83wrrbSUdmS/jhG0z4ooqC8rIBuwKXEGov+8UvBTBdayUpbPbmAg5IDm9NkaX4
qIJgBM9t7R35JZwgqPhbKypVSocFQdbL1ifj9er3E0wd2eyAm2OXUAdgyoNLU+en
E2YHPXCddQFfvBwg8osjqgO9v4THVLN5DEM4SgzPbJgrtmEPjfLoJh5Sj5DU3ss7
pApiHz6VsfLMmij6CGjo54peindYRh/CErKAzq07sdpqelAA6N2hh3P7JYuBSqgc
dJE0Y2yDX8c0LLO0APFuiD0JxJC0wvjLmzDUaZh60+NDYK+6KsnJbyuRDdEh3suL
lblasL6tB4hzwAbx/YsfI/r9clrHi+hNW6n24CbJicKTLPKvKcWNCP18STZE5uSD
T7KXGOqwajhllygIYpC0Il4v+GmFFJPfIZrBZHXY/k6GVcW2jyNfSHIk8ZBFJCp9
8nBT+hzL6o3ho6khxxVfGG+GWE1i6zbbwyOiMj3UY+beQ0PB1HLK7C9sBArX6WEf
U4VCAmlzVYcG270nHKRquLgs6pYe/vYjvLK6ooJf4SXkyhQOP4XkpE8psABX//CN
1zrI02vHkvm4UXwEXjKEIC0I7J8ApwiNSbAUphMxM8lO7/ATMTtXLnyRE37AuL8n
IaGHrLYt9Zjy1EbdKxV5p2sxN23WulaeNZG/Z57n8vhoUdhskPlKcqt49NjO6qe2
TtmCFxDcWam6+etT7PvAMhb0A2zGoCM+6Dfu3382JaOY2uy8vOm3nJTlgiY+WeM0
zsbarXKwRI1bEpuWDlQXp9IMlIKnidC0Y1QF2IUIP9GUIgmKC2loyYp2AFZVeyFR
fLwLArtT1fxeXpwZd5zMMo5JhypblnpHmrFm8bV/yPo0rorYw6Rv3SfUspeAYkg9
9YoE46VPcqHgAGJFnLzqH5mrW2LnnRpddlKU3YMMCE0+gArR2y47gj0mEFdUyF+6
apeHJ+sFL4X4XE+HlM46fy24ECWDxsBOcBITRiyaUhm5i0jBDPB9ts5ckw7T4MrQ
i37H9MIyj4aHga12TmFmnpdL6T9HqbBm43Z0T65EOxiROHlTacc/WOBR6Bew3lbs
9Vn2twiQSiiVnonVr55GXFqrUcj3NJSnC7w64WPm8hu5uymLhDIVpkr/rAN429Gv
V6FTxu2qUEshW9AGGHil59oihTsRUGgTkXd76Uu2NB9fQavTBbyyxUjrQPcIXSon
EpAb3Z52qckvv8tTyu72sdzqJwqYncgaf1kMWHbR1fuAtGKWsHN7AYHZPlCEBRA7
HyHVJq6Umk0MgiFnbj8KFl3f0YxHmH3sUEwW7LYW/Oji3v8+fTkZTJWninJrMV2t
yLg/gdHxxlyKVokNP4fqYAQ7B39t6dNeqjnkJhdT47qhK2lHWTYEWJmlD4iH8tMY
53ds7g5DSPaak3kQ9lpuAOAOeS7u4AQCUgnvwHNUH/7tXvulfjGr3GE8uT/jZoQH
LM/AmGQlJ6xSi/Bj2ZuB8LhMqOn0GCJoHqnAuuQ3DrqMEf9BGRa18DikzpfIUXpC
FI2cskRj4pu7GilAvdyxppIQv3JKL80O14HlhXmrP1Hhfz+9u++EoAHLue326628
3krzl/7qjC3EvEM2eZ1vz4S+R0dxX6iuUUDq6cxJyPonsOgRAiPzQnpmURtphFcY
BtKc2yM1wZKQHXHL+MpVNY4N68ayWygxTR6qgpyDcyg2gj8Rbheit4aEOoIfh2Qk
12++CfSfvyEciPiaf+/B+xwHy5aFZCrljF8Ccm27FViHLucJFDpbPZE6G9Oq0fQU
VOrmi9vMFraDtghMsFllrG4t2r6Cq3nzCOBxQiBkSiGSEfwvajwZwWBeCKf7N8EN
FPKsmZTx4kmSA11n1PAKIuoZf7b/oDTuNcQXobN1g3tbTkJrGNzuh+7d8aPs0c8c
dfyD/5bpdFvSnQnkInd54BQAoCy1p5qE+mTjFSiLvakZjTVkefhdnH1eUB34XVQa
ffCaq10sMjs93mJWupIi8D1x33/w810LZ+8svOUhcx65uPCRyrfkGGKXgA8dxQlr
570yEETR1L+ZEjPywnp19LJNTjr9jfjHDetA3cGgKcbXkqQWsEngb0X2nurT3/VO
QkyErcawy/tOXgkgNmswY2sGO7RqmOisGA82JtQF527u1LhcmdLaikB6ROB6MMfM
COiTKxMqH81HNitrZz449krl0CTjuQtAYmu5pg0FD6uxsFRefvcQv4cW93mjdHUJ
RVqSX/qCsSVa0qBGCpXz4g1Pwg5qWJ0W8Udau4DRZ0HEU/vl+Nsehc3XPwsbStTU
2cOxfJk3XmaKFdzKVhWt/2teU3V/sAkUnM0K2TONu96KycQLAezeHnIcuEFWpO1+
kEmtZd8Zw1HqN0awVLvVn5c9L3UIIK9tEXc1aoGiThgGYONfoxjkkzBPiQvH1gHA
3xYG2SQocAGxyHqQp6j0rXX1ZM3q44ud1cpY+NW+Gxf6ixoRm/vGBi+s7RLW79ng
6W3HjDzZvcvJ/kM3i3eMjr092T4Y6+FhrZxobOCfoFlg0e7K1VwWzUV8Kza7oWFH
puRL+NCBJhWWNWqe/3dcyPfAdaJ/AqsuBdz0wU66ZY3IK77WCAV4jgk2Fg006qfX
f5ge6VyQvs28PPMkLIevfew0qPYKONtp1ArvVVT0aZHnjwDEp6WrMWiqr6VNueDp
jhi9FlGk4I78LLPraR0TpW7AcESolY99uSBMlkbn9pO3J53inb/khjldYO4DvrD5
w/iyqFeul8xne6i1GBnVskj2j11pgPPe9J03GVTEwK+Wmu1Y3HvJRG2wnLEGtp7K
sUK9gRXPWypNNP+AfslfwAggo4uObZaSmkPbtIo4QMEJ0R7Cin3LVefxTKV1V6/X
j8DsZPUtRAHl9QCtS1g7hDHXh7hG/ICtjA3rTj+vmWJfrJ0NVKXENoLEiyy9FbNw
3UhBqlQfLX2uOntYeDVxuzYkixjCVf6YIZBYcmuQCZ4Ai5WuivN3SHOH28Vh01N6
IBGdQt+zY/MBy/K+OTMAt3QptOfJntrQfbiN8HA59v4kO2HEbH7uTheaqT+oeN7Z
D4zuVFY0clvLr0bDLSkE+5kNVsMW52GtctUSpLR7RfK8fmQ8tqrm/DGmqzt9n8WC
U6OBunIeVLUkjeZ21HDR8cg9CSKcs8mS18B4qe8mzzRlo3KtXyOs/mPE3s8Z1PRO
yTLHy05Q9HUBRfwofKvLY9WKHlg4zMTluNqm1ZF/4oa3NZYmXj4XSzWnl+OuWMgK
toFlu43sSwVgU8XnsDPcuda+IyVo3zNQDwj5ZeMEvfcbg6KvgLkTNMlkl4sdlB5p
MOlC5+aDubjFGIT+mDWwAqFEi6cqZbE+BO7yl2mPvojQLA8QTA2yHkDHDgP2ikbt
4jz1vM2Ya844gZZ9whdIkEAaMXh4uWUf+dkfdn+DsPNIvogb8WwC9JmHi5sSeUva
1rAAmjJrBYEMc2lCcesY+4NMIKY9E4MvCq5qNX/BHGdSQkPPQF5ecwh4KOez5r2e
2mD5RULp9aoYTe9n2J62sMui/s/84RBBqrlOq0KudTK4RVtB4bE/3gP3I5E63CWL
kEo+iJR6swFMFy47h1qxjq1365zQNwzDORxJOYxis/2RdiKWfzeIOCOPWjFRFLOJ
5NuqaROXV7rfmfxXrMnzuQPW2kR2dv811wTz3fcL4GY6fOVpg/oR6wf2dsKGEWLB
LuKpiwKH14DX9gNMcwOK9Mcwl0g18Duc5utWqbrVPeXn4OqE2EaolcOfQ/FG18FH
NGGi2mwXIS2OPVKzwy9BSk+zEqFhqCk3jZXAWVO507lCPhzpFIl3be2Pvy2gGyuL
ICVUQlSdQKsf7Zhv95inYZ11O1oinKV0eadt6FdF6WZpN9d0sOC5nU5ctQmijfKY
hVyiA9rB4d8XhbRpAIHaFx09hLhEY0h9P8gIFydyT5Ofz5o0tkWMIM66H6lC/GKB
vv6BTZjjTZMf49Z+NUbK53mtGbisFp+NDOr96RlJsgj7Y5gEMl2c7Kc3M9IyTegl
CI6fbxKAjeJFb4lA1RlXBHzAgSeP4+V9nWeSwqWCo3ucW3hLGUKd/aPILKeKfSKB
VOrnFiNHYSBzVVCTBFsrAqLv2hHSc58311Sj2sMVE6I8+nTYuGmPpQhiHxNRIrls
AoqlBqfVYuLVN9J6bvTe5B9CwSTEoEiLtvKbbG9Tsm0vx6EVRVsBNAg4WvnUrIrb
GMl9UGoMLLluua6DwYYPyOiD9tRKio2nt90Q+1J7sxpkM7+Qi7q4qIIM2ZP8suI4
vlyi1VWvU0kVQt2Mz1EjAs7EdoXHO7+Qmx5pJUHDFWzsc+YBkBWRuPlMeqQYenXt
UpwXq02CUw/h11KjYPuzLLwoujQOI7G72F2EvuezkSw5f8/KIaVtmZ0+AhS0nkw6
v0vfTjB1nNTyPI1+cnHDbg60RZeSNGkzbO2VUniV9qrowI+d0LCwy3Bg/PDo8HPb
Fdv3hxwM60Q7xwQAJcvNfZ8ZntzM1bc6Z6pP9VsryNEAgkGcW9T3vLGoqIvnCz2H
SYGUTbtWX4rpzufm94eTbVDjINOJDDyN7o9uTdFGJJUssXvuuo5srj7vboqmjYCT
f/JhnUq130+A5OIW3JMyuz/m+EhrNHd0LAi6eAZys5cdsUIleJyqbwcCvIYfP9V4
CnxoIVuD91MVKSPCDgDRTS+Aicepa7AEEg1GwRaxzvZn2qgyjlIzRhfcmWkHBNfw
/lXKaO70h8umhXVn0fztPoA3nrIqOCw9c1mIDJcGVsV+IHz0H973no1y/ObyuhMi
QKvXAJwEsKowkO49pUBdBZc+xTzBG4TxSAHqpdUcemSNNFGEx7nw0jID5KGNSUkf
PT2DFcJ/yhY1SsK4b7EYTtmQRL6TT5Qbev0my+Plw0UOrBKczzEuxtY458w1P7c9
qTVjWKJl1UbG4NEFKtmppu6VTJdSio4vc41JUVRHrB41OJU+uHKA+VuGHfvYbuYT
Jk4SwDojWV4mfOzWyiOwf41fxkZgXijQfA226G7e+/sy3dyS7GhTNM1R2Jo3YPTG
y1b9AMsrDvPpZWzA7XqrX2YEx1G9H/Go9zn3ATZp6JrIw08x8ND+PagwfTx9iRXW
5/Fbfdvd6oqa6TuKqIXZGOBZKIG5iEqz8P73B4LIRaGpqvHTgZdQo3pAnBlBePT6
++jOQ30EMzheIWafWu46ZwNos4EXO9xN9i9f8cVcmH/oq0UvQC67QQ5dZ7g8sXtk
CqkQDBUcxL1+/xN3mVpSGdy7ODCxVTFOJy5f570R5gvGuuU2FM05CEeUk9hje36s
ZWj1jn33Zju/jiOaBjrfnY8eOINrRiea5tH+oUDPO6GfgG11cs//xbp20W3Yle2O
wf6TdnK9Nb76zhQq6tz2Bn4VMynb7tfLqVYVg7q7VALzEGZALGXkVP2sQyMuLH35
41j5Zuo2xMjTklZKq8zgWieydM9rvlTkruIb81khABIW4gVv4GfHvNoO/LmXzF3q
Bzx75XPI5q4KjCPnCAy+/1IJVuV5MkQ1N1ErNO8oJ7JBY0An7WtH+d/Rhw7idSdw
aBhrX5a5RTc4ysYyHi50OHrWQjZnuxfU3s1Baok3sM0cpsQ5BBFy3O68wWQf4o9/
oWZH7GjCcGi/VUlKhxmaJs4Bi+iJ7M1uqtijdGWwH78QphRwm7dS91M3oftNCpbe
TlKBzPrFou1Y7G04zLHxswiL7tRwNI93vEWTviPqAAKn0vV1LK99DWywshho7upp
cJ/mCEWX43xZckEgiFzTXuG+KHvBZNa1b8CZhugOTCE1rGTYlZCkcL5NVnbPuY4r
nCOAhDnKB87V67mOgpGAizOnFu9mp1BNJV9Zjq9fOwU74BSiA/JQoda9CydqSQYH
jcQ18OEwecct3aMQ3cUNYCrpz9+UWtIbHP80GM2QDuUabZb80meysl7F63/vrmWi
MqhsIUYj00NNjKDgz0x0uGRUGK+o8o1rbFLmjYvoNcKaKZOU59vv5Fxk2RNmSBFx
5Hliaw1/CoBoh8v2qi5B3IPIRN02HMMYBpN4knvL83J3JyP/Oa79cxMwYqf+rfR1
wY9E6fnscwRYw/4ZcxrHyXYsDtskK4PiXlVS5rvomSR+cyxizRbucgcGgwG1Zwjm
AKww/lQDc5yES45FcFgB7tEjID2WvtuA12uaSojs6gLaoSY58dA/pzEEqcaB2SwI
gwiCOCRGpXcSH9zWbn6rC9ZqT0H/kCnJPnQoCu+PClbB2DEhUzvmPsduNUB3/Q3E
UUQTYucTs9FxwfdhMz2/dfWby0Df/JoCuDxo8bqu29W7yQpVd4aHs/vRzzyatPXg
duRukDdab8lkcQcatVGxOlpG748xzO7butxJyf5Jfzwzp5Obwk3ZcEk0KQZEuWq8
mhMARAQdaK84pbbB51aq98NEiHXHTFrFiU2pH4HeIhjD+9WTpmVesdYxxZv5Gb0A
d9R/Z7WAGbQog5edbS4Z+YlVhjY4zkjNIPwGu1PZbxg+hesSpV092ZQXtVmuE5z1
a6GFcT49m7WIcnK49qo22HyhG6O85gQuuq+gwakF0JLDFFsXPRPyLxXYgFUND6kD
joOP/bhtF22Myq53D4P7z7abU/i/UCh1iWXMOdfL3obavqtGCHc+X3dNaiqjcGRU
cQRkvtGjbM85GV/sTnBp1QUNcg1bIGl34efwBcT56XltG1C8ejEQkZ/hv+UunNta
AxjxCQDQTJDLyKb9d8irtAyDUNzZKFBwKT84UdIV9k7XccNN2eSQpGeBk1o2FlCA
GpiGylZQH5g+6xQGrNo43A6XI9jT4f9CPSpZYFXHMVGwcdAGtO1tyijNU+0BV05O
P5gVdFkGg9c+GAo1zUDnOpS6fZX/jtOxQkcGfNqV5TumcFWPV0XE8MpdfNNjVkJM
HdhQjHn8AewNDHc7qUWEefsg2h9BlXXZCfs8XY3P3qCD/efJ+PONGxOyXpkn7eS2
iqMTzr9c1bMIZ6PYx5AmfPAQTCDdw8e3umCrPUXJaoNLkAWRnclgw9ueZz9e/yzX
JPQ5yG/n132gvWghkO1NLwA6El+wt2zDcHbf7tg87fVf8+1n1bp5Nf6Vc6DlUCiT
mEQrhzlJffTh1MMkUTOBqJkG1IdwtUGtAxw0MUiCfMvZI6rplTF7ihdLsxYvUo8Q
5bbUK7rVPoDNeNgRlojP7lv0fpWd095A8axSIZx3YDNiYMfVW9Qr1gs/ZUzhaYE3
k10GRqy2n5f7mnQqO1qyANk/pVIh+GFaVQjlaA3je5TqMDG58u2+E9Pe/43QS9pM
4JxdqxYlYT4t7TE3Xk2xTdX2FPu232EyOTh8YmlzQ7SD53zYwZn3HlyLEWhy1y/Z
QSTIB8I19wxQt0xzyYhRHIaBx+Pk/FMw51VDgd1AxobJTmfTeIPVQqc8mK+BmTcF
LS9sphq1Q+a1bZljN6OZulg/u85R0CbIY840OQh+JlCz+S+16szFyIA55ycITlri
XNBw1y76SwJAT73D1LvORhyvKKYbfuardQuCum8oA+85kuI3F7c3Z3BNE+dq4owt
1mxfmbcbA/iwjTzU3w4XpV+9vHeW8TvrGn8oyRsxqmqFXNHcB6DnikPRIljUbbdg
Om0uahBW2NGoTQigFc2V/M+s6CuNk82NqXnRmG7MxQoQSI777DW9F+iyUkkP7Xah
n2QpIZ2RpI4ZB10yrAC731kzS1fxTq6Jv9qgDdB8wEMIQjse311S2eQftPq4WraR
KUXGcfudT8O5ejqOCKN9Qu6uHnlA/YGBhDxS4Em9Y+DfcV+51lnzSFRY4b9rmcUG
bs3qOSYPN49stWWhde1FopYjJqDq+hScttT3R7KDA4TJ90bl4sLS3/eavC1VGLVM
kdqH1AbzP4qF/jW6Ei4CaDWXj/TBapHyRig8I7UwyCw0wnbENXZtpUOI3CfSOmkh
tkZ+jUrZ7HIByo/KjRyHzImIxltsCeWQxW5aZ9GHuGfAziAB/9wzYfGLukEboCU8
bTGb8qQkuud31gcw3d2Y84WAiTx5or4GMz1TCCjU6t2W+FhuhVgfLImlEHku5Gsg
4UvoZeUf/EQrXWLHSatz7LQb166HHYtA8qCYj92biVQi4cJVN7IKKhDLpF5w1+jN
Put2amNmyF2ML2Sq+AFdgPepEaMRhSThBELa6uzkXkvmLtDVCRgVPHzmRCctc0bk
PRY4ILmBh7UNhiDZCB1fULLElJ6L9RsKy6oSwu6Tvj7hQxvtjZI+sXjGifq1eCBt
o2BF4cVsigDdNfd3gjROblq41o7iFXcaQP2c5X8YlvbrsCrkOsrtgmFvzZouk0vM
MUEZwRHL4bGip2hmC8Lz+6/AuoK3SKc+23qvm+AZ+NeOBfXW3SH2R7+9hPo3ELGz
NJBwOw7mcG9LW6dL218HeV6rjeTAK+sVUtuVYK8yJQsbno8GAZzKDAN4+RLuGb2G
hYgSWLy77GLeZrlI/nB+Cr8LJLyB5L1VNqSw6xmqv01SBYbKrQr66Qt/Fsc0DTUO
T/YXrptwWFaSAgFyOcNJPJ/cYP/FZXc3y4IM0ZBj1CXYFiqLrFd1db4eLfsGP4Ia
gXZ27zACb/sGkGKB72qBywEDKn2iXr6DOrqhXSnwRJZE2GgHe+c5SaYGUzt5XvGw
YUE1wxKOZPy5z1NdmW0rnGfWT7e32SFW6OXb1B6U7LqWrtLjpnuYJ2ymcqUWMZcr
hEJjXWNXwuvj2pXVsyVqgox2mOrjjU/OSr7sQEidHq2a0jFtEqvgBQhwHL5hFFiV
XN190fM28f/77XOoHGsRWFq/kxd5ZbUUdDnIYwqb9As5bwAJLCn32tI1BciPxoJB
WCSLETLkKrSvp8+QnrgpDVfSf3Kfnam2lREUVTNkLjKKubafHZ1BlfaKU9p+SHqR
US6J+fjwJHQug/eyh7aZJEpWDFyIl2xhOSjax44AT0ARtVBmdSR+u5+Qk0MFxPfI
9sAA1lmvCtAsTgFkwk8CLNRJ2hcWaUKKdOw5bPZsxJwFHnmju5h414MybolOvIU2
AUUeKa9jsAqP6G8m9Dbj538Vu4rCQ5vQPJtEmFSikEWxn+5Iy/W4K4VKwEgX6AR0
mWXRwLzWiWUrRjUV1Ee50TEKK8shdZD48ESDm80Hr2B2P/P7WbdDYsXq1O7HsyXT
t5wdRnCanfhQQoN+vNPiec8bbF2qv4Dt4RIr7JT+Zjy7AhkJa45DdydPG0WIKz2g
Snqp8b8GOziPGElgJEbwXikvW56KcVqBRmX1vT6UzYS5io3r0ciMo6TOXuzanDIY
PJrhW+nBR2+ORtet4KlsgCUoMxuJzfD/EhQnGmcILqH8sdEINtvjYSMl41W9V4C6
As3qP1y50HDcw/RytuPJDzjykAXywLJwgwsFRYHYl83JVbvQVCeLOmH4JzQpn8kb
tZL07MXlP0f2FZYqKoLBRk4mC2S/p99wotRIT8ADVtSMCGI38XXH2L3iJ4iV94u3
6hUgbOXzwqAOmJPza+YLJw9+xI5yX3trgUK3xdJo0a6h5oKOqVvUqh2R/bnlYwdy
x2bNIUzemNp9GPqk4hFrkRS7bHHcKbR1e6PcEXIaQUS5Zr45EwVh52zjg5kvfsxz
1uV+/4ni+wGTPjxaoLF0t0Ybam9LRD0JFHNrj8byPMfWKX4nhItC78mpR20fw4QW
hYSsiAoJYIVgJfqJ1n6kfodI7M7e2TQA1ZGErxD2OXhSyjlsg5Zf5eFftsDdB3Z0
aZI5+pebi+XtXUF1mdzOPmRmviFsvHe21vp6IOaT1s+oJo3nEFMxdIcmN06/l9gR
lBG0WaeJCw5AnUYJUOcTk4jLD1AMTZAArHoyVRWKccTfz5FlDE0BxFqnx8twthfm
RgcL9Yc/7pS5Rpw2h+zmNN93GIehhhSXWV8MV1WY0uVRnOdLVFc0/BOL8ErkqMbn
fxLvjfzqjBjCYE+/JXGb6MN7DXO9MfWxRBTLucVvaqJQFJPKVy8/KR/kXw4nDuy+
WISCgJKchTQErClMJKxV5eUyopiPtMKUKSBOYc4QMmcMwRIOlYOxIVnmTiwU+B/w
ZOaBGRATapCkEVQRKNHFnOvTu5c3V4i/mBQcVIIxrx69cqxsXjolRMT3dkZHxQBx
aCbhpnzpICAYHDLqer5T401Ed23QyVVoMCtdyI9HpHjV+bYIQm6ih/OHECuMhhcn
zlv5BA4z0KtBpaqYKQqKwWGO4f8svCY0mT5pvnACIufk/QpgYqR0/hrKq+Gu+Ecj
0/fFldAucr6bqeN+18PHz0FXkGo82p7AP1R5Xw6K+94fl5vhxG84vZv7tNeB3yhc
uPb11S19kXidWZ9wDR29alEYznAq+rpymorYvphL2VKrM2Idg0MTMXHzCVHY3viS
qbTsOFI9goAiSM8Vaondxjb3VUdqdlsu293cbvHkYOMGE864utaiAGrRGAxMGVv0
9nySOrGAzNn2qQci6yxeKEb7Iv/1Ky1tqt02YJ6iM9eW3aVzIqs7Mxh8MATvxPnS
J6HcLQdx+nAX5KaveMBf4NnpS+NbSCk7uq6U/uXqA3NBdlIseUARrrtG5Jawp7w6
9a9oSnwMlk8ZuAmeamQ5LQCbTvooj4iNWdP0i5yM1ONQqUrhSR3z2iPRKXcL74GU
rXPY48orGcnnK2chJ3xZGP3NI3hoEcjIvshKKD47tyVTsxSmwAvHehFjLXlyuQHj
8S2LUfFkNheY9g447pafgj8IaywM8xqjpZzDmZqfddSaDOrmJPc2O0Br+y7BbwlT
46I7la3H5VRBir5OgnFyb5U2BR60p1b1SZzJlAWbl1GVV+jvXfr64DvRUcsFyPxH
pkyFmAHjGX/Ju6rt1ney6TJyMCvLPmFX/Vc8RqCJnxLtQSLfWImseBWcb4ysQETD
oS8gEbF4tzSRfd8cpHwdjEsxJhYfsvX46/EusbT++3rnV376Rqu3+lTN//2NlkYm
088Luyu+PWB8LSeMOcCWsbSeZbi3uko578Sz/Rs0OeJjBykcbKO2jEfuP5cs4aC9
dv6nOPvMAMtyPgtG779HXyraXf+9jDqWH7QbQ0GJuHnMHPjHxBjAL0syIrWus6O9
Yvv6as7qX3esQ3BBFgKLVRqhmI1q2poL3VLnnJ6l1D8x7XkXVF75WI1kyZEh0CZ9
RlSutz2AEA8ZddgBJ4NVeEZlun1c5QXtuRrYcJTPGtINmrIEZn4OOPmEJZKEOqVX
70iB1uL4rUZ43t2LOa2qUMUHHedsJ3RdZBeJfy4fxLDmqil32m/dpZw/SktA5VUy
KsQ98uvySFj4L39O9RoeyXFaVAD9LeEY0VJxpXJENm4pmzSeWnqn/CV+KOg0pkEu
1dp8JJvtnVelqnVa85do6SLIFo6n1tq8YZxVdB0CD/u7crUOD57T2Wi1bj+d4qkN
CDDHXy6xW+BL3kOEbx0jC+x9cDtXRqtjvIMFdk/DOPcgsZoPWpdCRM53qfgiNww6
BKuCPOgKpH/5SaAdsXFBI1DuP3ESCcHcfokSfAUXVn46AHB9xN4/8MqAa9oMrKdM
agzCWS3yEzRQgjZg0IaGwmNIXurLAx7Z+j0Lhxq8sI3h88rj3CqCkT0JlRnUWEIs
zmVYBaWOt6lH7cLZmwBrSXRaEUr2PTh9e7W88PSN5jOYXI1UD0oYpkgQt88pICAu
LUuLtcWWw82X4KC1vc4nX2XnsWRmhf7I23HyrJ1Unt00pNWlyhVfhUUi2bz5SQRE
AnHGLwTRpxNVs+vYGLYYz3OmcDaD3vPX/3tHDQXrxUDWWs5P/NPwqKjMZ6Fw9Wsu
oYBRLdx7Ps4iCavaYxuNNbT7AjrlNyq+FRJ7Yn89sANKCVjHztzPb03S7sWksPed
7lE58KzDl3eSw6JR/pxA+SLBXcJvKG/Sibh/pAg0FLVPk6Fqs/RUm0JTU03JjA6k
HFPUmadY4OBGvYXu8ds00vWnPxdJr3Vn0ppEloXOVeHaJSSqqp8MR8b4kVTfO8g1
nJiJR3maZ9sPYJRqDZg0QDsWMXVqfNtVpuaOr01lzbeG9IxIT3vyIY2IxrEMfm/z
ln+SA/cKQNx0ItzPi61pE57skOG/7vxQFVNm0HN5FAYEexpAQjAl9EdHHwdgQ2oN
Z7ciLJcelniYUqmsaS8uYbMV3VXZQgx6qgynOwmBE1INf0ky/Zprlc6MXRVTZqnz
+KiR5bWL2K6JL48PRYpWKXERCbsjRwe5kFJsMq8GX2b+kMVsp4kDXR79ZR13pnXW
OfC3pSpxaBLLpCYR7N4UjZW+1296pdaAXSnGhVE5QmPNDlyThFmL89or3rHLtfIt
yNw1teFKdLzoM4hyWBmIWicxOXe10eUB3ydW2TxYpHmk1FhmMgEIdiK9QwXyNxcI
In5dIExHD4IxhcVWsVkldYYhPgcBskKYkhW4UDtQFY5GplZ7owZdRk6AfjuYPLoY
tJBG2mudWmD4/x0yQzomKGNgM7MRUDxQAPTOhd7fFGK6/oosfxIZ+/6sagDHTIDZ
/SFZrSEeHRjIlqUAXpObhMwnTaKaTMW15zIx+3PrDBK4IrfhSGwNQGB6D45srw1J
I6q6wE+MtsSALkdIJ6kLj+EfD0rnjHPBZJKmmuLYsiD1xatpCQoqy1/rXWVBRCaa
4G6dyZUIa32jRkoA07oGALYvZDhHxwW6bDk1GGkesfVfS1fsAURjulUIZgvhFzmV
cbUJ1Q0yRsLMQgGdORSWFH+pBFkrUGotckMv7BFDQpC51bfCAzwQA9kO7CvcZVk7
S28oYvjklK6EYX4FbDW0TZdVqEiA2jK0X4TXD0YhhCpPyQaSvpBUwVKmsBMNAzD6
t+nYelsm3fpGTulltQ9CDGUIBVIxmztUbWEdsYO9IJEaWuo9YpxCdZLPv4JZ9pv8
SX4U+LZj00i9V8WawO34MD4LUYWB6WAsNJ6VAmSNn2tdU5NF9fwPgvrN/ZUSDSW8
Ifw6bzI8mh4FDZf5HIb5S5R305b8lPfgaNJ+fFxmEQnTGhOM/zGGOclbqJma70gV
ntueffQUrdCJwjucyir9Ns51DZvHxIu+w/bU7WT19T1acmnPUCDhYygQ0Pdm8+1A
PFf4RWkVcnObCz4KppUNSsKID+LW4yjAbFkkd5k7qT+jn/alxEp94R6mBdFLp6Bc
YYd5zuSeVpXkoV5VxmWeYwUpMq9/CgNRBn2MyY3JcEFAeSR+VoV3zWp0ab8IVGjk
7W+T0K1ak/HMpXwMxlpE3INpQnQnddJqewS2bdox+tvyKJjp6tZ+ZHEy5hFecvsa
D32Qv2f5Bm2KmpwNZpeifl3X4f0Fz8Ii+mUe1R8zQ3j6bcd5Al48F64BlBkWecBr
epwfDBAXqPYnedJFm5/vheD1WMEOOgC91QQOOSk96TwdIH8KGd0GZa7ZP0724oAq
CBCLdJFigqCtkq7O8iRf0f9oYzVhdGrr69nUhL7OjAtyCGItVLdINqZNuCXpm01G
lZxY7O7thkrjEwtFA4uPdDgzPX58ZpjUqcvZJchmHWa7upnFNqVAdkw7olp5NEGp
mSNekK3X9b8xgKDYVnmvZjphyGgTVSNJ0uha1brZA6oQP0bhDtGjX2ojdWHGlpAL
EUdPADZHn+G77bLE/tvuXHYMMccFp9tKqKB+MtOKPKBeZ/99xU1QTgMIr+PhVlw7
LAjO41YCa19XE/7Aa8LMC+LSltqbQLVolzWDyjIumFHgpld6GCBk5cz8m0DDTVMD
2XWfRqO1GSO0jhzrH4gecTO086hL1mox7cH/a/Mk/IR1ZED5KjnADCPIt/KP2x+8
ykO5k8StEwcVUWBTpvA/wsWU+h5jwRSS+XWL2eXElznwJRYrAizGb/XRqTJ3AQ39
E2xiNL8vJ9LNSfA59qXwpWiaBz28G9JZ4+RjUYHSoQACeoePJZm62x/DB2SKdwRM
iVrORdj61QTeO7MOhvkvZ2PsA+cIK27c74th+nHDX5JLOUP7WIXdktKUT1vqh2iT
Ot2DY0Z0MxTZSQKhGVINkH4wsenLMR1dQtoxLuGRIclc19ug5B2dkI4x4VceFqrZ
S4by0Xj0LH/TYuEecNRmNdn1fLsi+9MiKvwVoIdKYNo8wwK7OQtH47S9fLy7QOiG
OOlJ8ktupuOTC/5cJe2FHikpSxuDtiQky3cz+GaV0PuvPBszwNpv52le3XmUoReB
zmkHpAlOHuobw8Jkzdv7j5ZqEyyw/TYhLZ355rGEERSV7Mv91hy8057w47E1vsny
FucN+n8vQG96k4gjsVAFwsIsaC2vlZhWQ6pgb7UASX13HVH7x0EwRm3EYfNiDhTc
lbv5xfx2XlWovMOcGwJjmhLHWrh7tB8/kk8glcUEuVoryd1Mgc/gX2wGTFxdBMS6
bc2gZiH40TfiHidqZGw8bw+JSaXr1KfJ8ZSStPOFOrmmCFNCE+qA1nYDfsUpS4/l
A0xCVniAC/ze/ZOmSkYGXCn0+0423pqX+6bWltdOv3MSzS7WAVSkg3qhDfLdp4sO
JO4slT678bk1hmpj0+XMnnNFgNjXAZfuoyv/uOvv52Cib4AoXmIk2JDWR4F92NqZ
weZTQ15PvPlfL2YEO0t2A5ae7JWuyEctvCXp7qC5DKSIsL3LIJhP00Dk5APChqK1
ALg+1ujedMl3+z32hRK4NIH/Ou+2t+MGZj+TMVYGkFkQRGteZbyl//Quou3E/NAN
W5oEaEKCuxjKmVJftlBmSgEfB3I4QK7f2JCf+lMWGAGjU5ZffdViJgyJRKtj4KN2
VwvbcFMdVoLq2IhTwmS5IEc4J2l/vH6RLcqgaAZyufOUCoZfCUY7E+z3rFXzjnh0
I0YBau7dUQ2beKpYg54sJkKFC61arMYM12cVjBJuw5in9JbOWSJED0aLMFCKVSOA
7blHjQxWP0NCoOj+5kF8GpvpawZXrAgXdQnWjkx477/uVT0XlXZWYU3ZQi6GFo9N
rwsNQO7MTKxjn31rLiogpeC2CvpJgx2cUfxH8HoXnCcDL+ihMwa2ZIM4VrjnpDig
BJ+YPmfV8qiPCbtQ/Oy7TdadubEfwFvakJYsI4bmkl0hKdbVjuKS9y5tCWCdilKR
sz0UeDS18Y6cgGY9nyf9arSBDH57rZjfiYUxQWmnOflJubveziqlh1bhrwr1iiUr
qet4yRbyb41I70gqC+YJt0y77ivuuOoRvmkb6qKR/viYd5l+SxpNxV11DiFsy6Pb
fKrkbEW6EENrbdMiaJHJkO8rWfTicm84DgmEy/jollwl0sCeKpVlrDmaMnOyWR8i
oWm3CYAsTnfYRtSDXy82KarUFdDFevtl97o2V7FnGZJvG+Dn/Dd5y3SA6KnJHiZm
kAftBViFF/Lc1GbxhXRMslrBISgaCm1bnr2JE+i4fkdl20+nqJ6h+uoz1XLfmKwj
kO0IJc6AzufpbXzuLXT6IzsJ0x4yAqjIHerGiDQcG0IspIR/I1o0yYCajjETZ+Fg
ySTjheyUHvk9Od2bMFQHCMrPJQRaIpYipq2C8is/ZuASKw7U+nWKA3RJvFY/wT6J
+ihMEGnuDgonFhRXtTEfsWo9j/x8Hfk6BOjTOCjGDbuLrmgjB6bbbthUD0np0eKa
HCWIpTc1HjORPp+6t+fABfUyB61/kmZNw9wZ3QGtMQg+cfrzcsaPES4QMLrjBgr0
swTVtO9UehrPXG9uy69659ATLNRA4UhpvcmhVUV0KDiqNrsji73mPLzSt3nsdNki
b+IeFMDmGAxkUxcbj0fWgTUQhxQaVrYuerflBEnIsmCWLo+yNBm3Re8QUzqCrsW0
cuEgx9puPDB7nEPRUJwu49Lya8o0UtphqYOqZXrNcT/NkiiRxOxChjbXye12swvW
BaxNo4m7i/EJ2rx2eBrW5MxmASP8EbXFUtJmNbghK9vDxujzxyA7JBX24bESWomb
QawaJuO/TeOFk2LNZ5tAc+cOShzk2MW+YSCwwt6bWlFcZxEhGMcEjO3+3Zv81aQa
2e9GoAOIZdZ0IdlzPpGXDVBCiBpQAXLZjB0EaQD2XjFaD035/bHOWkUBJ3ILH0nP
EJa003YTWXKeaxRxPNZZ8QIl7bLFlQLFSxWTo1gmgPVadFGv+RnoSBn54WP4ERDH
nEVwpXBrFSoFNGFlldLZ8g2bn2EqG/IP57jUMQD/FjMEKVTFXoy8M9F7O5KHLrzb
r2WPNcBIGwl93f9Xv1J6IUGU9qSJ1pr13fV7M3HeJEzogk5EBAUeNelqP3YSwwBY
gvtlsE9F6W6Qlv8kYiSDVK9chw+r/xpVG+v7NCCWI81f5cyXv0Cst2hEFQs4EaEM
N7iXWJhreer6VFn3ETxok7sVuAI4kaPNpfQBSDNuWbZJCYNGdUmeQZsHkvQ1VxWQ
Z76Hau50gXvWmEKVn+N8OKECV4om4BFqX8Xjsm5IG9CkuUhowWIlrpfLvq+nGfWm
/dxvXiDXxnmiVgADGJByI7cQHZuzzSibjsi8t8kIaK3xF0ZGFCBV0NerTpnftEk/
LqzXg9zuFc6a3S7aPOfozUvxVHWuBIaNYDoZabuJePus1oGZuNrRSBNKyJsssIpd
7Z6J5oGeL9GG7RPkOnzA/FQ372wExgyCCLErWfLXwphFqg1KVIVz9jtXsTZiJB3C
MFS5I7cSLOjV+PJLa5qxNE7yan1hSZemZ3ajpgapMZBaG8/kwzdB7Ue1+IWCbEzE
RtDzNkMh6JDyeG2SfUJiOcl3rYxYl2mfbh8tbJUquLtTdx/+csVY5/KzJYIrqLVa
DT5v3i8cZjZSEbesITfi/GlLg+YI5p5+jqZlrVj4RJuM8nHNOTwR3Qi3OBNd3i59
ubTEnucI59p0LiviKLD8SvdeTSIifEcQdfKzkv6g0E6GVVC/3T7FhFtuMRbB6r2D
q+lPQoXR01D5ntG79B3g/049X6rSEN1qkay7shekKiqeeND4oG6VvTu3TXabOA0d
duehK9cIoG/JXIghHnCvDOxzygDFWX4AmjgTlSYTtKHfWNzxLm8xtEp9Y58GaLcs
nhnV+1pX+P/t815IVKi7RIAFbVSUsZ/ZB2mTK3wJ+TSA0+8EnG4bHta0DWY+MmFU
MXv1JRvAdUUC5KFX42uWyKEYvTz6kWIRDORaBCNc9ak0DfjhBN+7eCxlm1vFO/dy
lnsR7CP9+ymEgc2U1wy6YHlYT2dMMj8iznX5lwDc2jov3eCVmVW+RlbrAFI1T0mk
bsgemUeXLHfV1WkVmco6ulQoowOA0GtBsvQEXGzJjMo3ZaBM+QEDXcDZ/Kfxnv1g
RWoiWaKkOGzJU0KJ1dMs602k6a/HbkAkLaDUm5T9llzNf3x5cXaShQJWvXXgJVrv
p6UvV7Js0qi1z2yN82l4eWdpUbazYr1DBVEDZETDXBLnqhAQFoL1cFtfKPnKP4Dk
SuDo3aOYxOv/vtudUhaWHGWXSkuR2m4blOb1HJD2LVoCKSFSbKeL2QVmih2kz06H
/WJrguIM0ojpNeAldfonob0sWZM3x66BPyv/HtHV7TLDOLcv6X5BdvHYC4+AjeKL
/uj1y+NJGm8hGW0rPSrFYnJ6ZHf6j26CaOoKKxRbNOdG0mTLw1MpTyeTJvM5MI5t
lYwuBgq+6uEXfx4oi06IB/2j4BxcHKXvNvFTylrFcxAWfWOLuSpvVr5h8f/lG41/
QfsCxlprT0a0Ylkm/21gy5SdT7L+H2kf+wHjN079bM6esYM5oTxqqAD9NclsdIMm
d7P3FVykW6Fw+3O/hFmKFQNP5JeEhxhh2VGRCwCR3a4Jm4q2+k3I3NFzWXWeokOx
DpLBWRREeO8WXy9+2gglAiO8EomkcyqlDJVYov/Pqj/0eav5nFIGDjw91X4TgSFs
yA8GgJ7O+ZbardefTX+bEIVh7QZtJUcaxAEtND6KYbwl6tYb3isY4XyHBvCJ01xj
P2n/YX9uRMwX8yPjPY1w+mYzIZNtwnhNKxOAlqNEoyPhZYj5aCvPbwewJANLxHTE
8NAF+oHnfd5ZoE7QiT3xPvm+mk2vVeER+a5gkMdtZxvCD8JRcjfIx8Gc60okVsOB
ZZa7aXIX15h6ylu1AAgWTw3KGXAtEZ2BPHnGyYkBlLBamQ1AfkhwzdZ3VAOPWuOw
6PMF3pooMIWiq4D11sVH3UmFvW8bA3Fy427B0Hlz7hhSF23Kn4tydrRH1wlbwrA0
/JXORe50+/15HuEe7KP+AR8WgdGu7TN/+GHDhMC34b56Q9mCQjsH4ormEsQudr4j
aoTgQzTqHUpgo13bMrIBi2zSobgBs2G12MQgI6iJHdSFaXo8XFWz5zNufM63EzaT
3fvMT9qB8xt+1DI/Ivsb5mCik1jLekhCxqPowsDMcq8mzWBFSp25ycPltoBHY4AZ
MbjhAEIuHfwkWkIhLy2BDASNynY/z5Okq0cW+gj+fzxIJtbO5ej5SB0LS9ptXTS4
choKjcEM0MAn3MCmTEmJLROzF67kPt1XiKpIaGeFACWxM7SWvGB6bE0/ohMFchet
JLUYrMgp47IhbU6EMbmwYcw6KaV9Q/um6HvX8uVTYwjgZ/R2Z53dNN5WzLZ+qvVG
DeaOMI60kBMKTlQhBdcQ8nVRdI4+tOfeMUvUutytrdykorj/Xvnlqwz17bpLqzgR
SkUwXVF1VxnQlojEDihd4lSGZmgtQjLjpvGPkE/kYsMPnD8y977EEqJmtatI7lC9
0VQXpi7FJvlwTJ2mtjjyqSskaqCZKo6vWhnjM6TQ9hkyefD2iFqc51QrK4V1Cat/
Lyj1V7rO/yS5csvWRzD/c/qlWMtJJuL/HSzzHkEcE7IW8RIlpIRNgrdWKVrNSnwk
tjZWraAuEJsvawqaGNusgodVPrNhxiE+xili1S7LUAFve8xw/PDhMl8rkOoQRMzS
MU5aDs/hIJCDWyMwdXq5iIIrqMEF8WN6krwf2YMkHJL+uNuOVFFe6pJe/aDxsU53
jOj9QH4d/9kA1xvxO7SuSaJmmGaBDif27D8w1m/Z0fSRl+gWo72ayjbVYpGhizAh
d4YaQAe+U81VbZeoe9rtQkDyb8xIFEwGSdCVG9mry1Kq7mC7OUALGnC87zvqZ21p
Z77IA/oBAcj2GoNqozGPDNe/8kpCxWfvioRu+BjQXUQaMmScWKSSIq6XogZBzoCf
dFHulbsI1tA7bq0ReV/dDgThGeLJGlED2Ux5A7THKlRuHIo6CUCreaFQ5JIspQUZ
v3GSIiM+5GSiTI++FAWGuZVbTBoCuHFWP2i0WosLZKXWHG0EyNtuks0CMiHnwzrv
qSm/RSSkggmQiMKnoNrZ/3OUOvUudoXA/z1PTTvajsIErd0Pt6cgz4R/licgG85N
k2yX/Bbxa6m1OM2hT8W8BQojrh1OOKJoJtZTZDxZxeDAqhsARic2NNxFjXkGnFIR
AU2M3n5l4ShEgEwLh36Ud3VXlvq7WNXB2PCYEB9RCKtPhhnU+xCgYXMLlr0dmcOe
TuhpZ54PAHvMEaQBv/uH9h5rirz834zgSi1wB/IVsR4qwsSDiyGI7V7Kw9G4zAUG
Gu16e2z42DhHUsPARSwt5j0hUaVARKBr6Yk35rEcuuHeDqD3ivHz63MasgHUqdI0
c6TL1uL8OfOm1NIIc7SLnKNlG4Q12r8FxECd4vgBq2bhxKhtzPRIALjmx3SXLlUz
eVychqczrYdsN1e6pePFVmPWZsJ1Pmxk6A4w0j931dhZxNjMhMt//ehkGG+FD1yF
jX5+2ah7FiSVm4QWo3X1VLRk2RsNpBdBcEQPxqEGAzzzc40j/xwbce2WffB7bk6K
aCgN4V5tez32gW+KY4Qq80B6MNc7Pesc1jzilxl3+SLscbfa7hXyCykNU3X3DuSB
jPlOTkZanlfpzdTnp3rFKfEBoikVVpCLi8Fns7S6HA+W6ghy5/liMoHjFWlfv+Lf
U6GRbQUuq/MqdddDGqEEzuG2qA8D7yGqDWeIB3A2fpAfl4pF2g4izxVm2VjfJhFj
IDF7TaGzW1Q1gP84/gDc82Plyo7CxoQCkFlPwTS8MpFPdvZbkAgIxVERye695nLC
4bd9n+jWdmVEmcF4F4ecIuzv+00pBnMuG/c8i0FchtnfAF30rnCTwpTX6V7BVPpt
39DUdzTV9Y8RDqN1Gw3EuU7R8LMcqCiqM/8iKpwpfxUb0CDPhexe9zXk+BQrVWN7
MA10//PhxFT+N5OodkRaCM6yBS2z5m87vIwZrEdv6OuqZqNRO1m24KZcsfMfyPlf
Jova9ehU9x9Sh/3JBwijTpomBkUbr2WQ33+LIUOh4VGaUrcSGOEkcx6BsGp/hWqN
TwlCZ9tFFsJvwqIBamXImUXh9lr/Kq89QaKr8meqZdzV1vN6SC19sEDzINqbOoXi
WK2fO84Us/CdJa4j5k3tq28ekH8o2ssm7VNo92D6bCqexHvcKeNSUtzCddJdCxTi
3TcP00r3gMe+IGVfGLylXcIHYBYYYaIh58/Ex3YOXIRYYR/ixkib+xpNxahDLxne
my/ZUe4Qopywzy2n4mAxmDByiK86JlwbAeWPU9Poq/xD4mt9EROcbCLtXVFOKw7Q
Us/0QFvov8/+iwL5UFNsEuG1R5QN69lVFAUexIaKRxbZDryhmtnC4NvbSzY28FFw
d5XJJbOOzAWvf5YgQFu2AJ9mIggJzvUyMdXndSgHv67lA3+B2RDEF2UM5WaJXkF1
5AN8epI/Bq9WU8drq+wUwrSeGAUXUIOak2/l2kGF/nA2WuFC/IsX64oWYsfo6HjC
+cXr5404/Oj/LAj75jMUzHg9eTInsIjERT0/BnN8z0gH6k70iXIqCdEjDF9hLr3y
8Vqf7f9cgy0y3LtjKTTKJwoY8KAn5+dHQ5VUxaUfxTc2VlN4wWL0xmRSISyGKbcI
3ydHt7mpMSGw3IWM1dIeGSMIbUElLm3p3aJsakn+OttLYBXaedDLNLDw1z/5iblo
IDESF13VXS2nkQz4qyzKVIOxBR2tBt+hTXwZaMXYH7OgjGXgjbESaYGxWitTDCiP
AelgAyGxEC9TUdEKWEYVRljDim1DJqQVMugDRQ90bWqkHClvFg6IXGJEyBHICHJx
O6wkFFEcRvUOvr947cv6/4RMsxcBnx3Q8wVspJlzgzqKNL2FQXHrEXq593z8S81m
U5bs26zbPh8VigdGKJeUEk1FQx04/O2ms1my+0VkkrMzUmrntU4es5M3TMSDTDjw
ZnZmBlK8+mRBvTPD+ZrqesUdCPmrFU6df8Gcisit8JG3jC5hKP+TIE8Lmaxez7JW
YxEoE48M95KoGmQUB1SJV+SR0KuUHJsl+DSnM1YuRomHCIOFOVO1iLEyD7GhpAtV
JwrtqiVNLsHYXxq8W/gl7ZUF9iiGeNBK41KZYdQXZzz9CdZyszsuIO0UpZpWZM4w
IAoeTT6ggO98QGaTm4lDovSF49i0lihDObOlXvM7kkPrcgySwS6UT8RHORDvTYp4
c6VubVWf+3eRJ4nvgkN0shEev+G51DscKXL0ipEO03BspqplJcDa7CbvhkfbN1h+
8GNY/mdNK9S+9SBHD67a2ck0kXmkpOIlqk852DfdRxvc1T2L1QJsiOs/JdODB1RA
c2P7DMttn+TZ5gnT4B06mQUH2RaS3rkKXBQzucII2Dp6urx23yo7FveyH6DnzvHO
kN1c9LWijVV2JO4lsuZkYyXc/x1qi40d0Fj6jDs4QNz/C7Venm1eygxtX9mTgsjT
xxXYI7YAH2o1Rtiyqz2hukIiCSUZs9ZXnajYMnHiBYq7HRA7T5hB3ZHeVJDrQzHG
f0grFM0w2kRw+NwOUxchuMWiP6/+C1jlWtt1biRK9UqA6V1xkxc8Cw+sREm9/Vq3
AffZYJlW+VvF9wQYf222LsMW95WEKAB6faPZOxEE9zwu8jVo6qc1v7M4+Wc40Gqg
uOsM8u+4ivctly3847KPwaU7l3jssKzAhohs+YVI0xdFllL9NgG15rXq0ePUPD51
3UB83a2ea1lRFD7tQcuAMWCpGEWDJGTzbt2aFTdlRbqxm/Q0S7tm+JIljQ3QFpPZ
GnyKOALIySdz3mEfBlcuW3elU7Jgx3Y9E53r5VnOrCp+7u7THmorDkoRYnHulCZx
bQbyfanJryJMlrG7lHDdkBDtozd8aAXztola9m8T0HzNT67LKNZjfqykt0P9DUn5
bnRt44y4j3W/f5JyI7em7sEFsNjmxisOhkkXgRmEgZrDj9CWKNN3VszlQaWUPdCl
azkO1cZvcbujEJjS3fXDlRGcOIUOt318wpWdtHRTco5ldxFJbuHvOm1zi8KqE9pB
rPCpnVoBMw+v/e8JxskBfsI5ETbqO06N3tIF5Rx1G/uv06LoQGM0VvxW5JeincE3
ptv4eomzaza/NPfA124m4OQsvB8nNiHR9wY7sQ/ym31nokDRP5ajMRz/9pOQRom5
vmTWBY/ccn/61okS7Fm1OvGoYCX7XmPHaRgEcmRxBhbqdlqPSEYDNGG/meuTi61F
ek0bs8IW4VqBQ5ylf4dm8ohRCQ7LOKFzDM90cDUUjGTiJjxaRksg4Tlw5sEREHIA
lLEHfhBnPobdcxoijaVh8AEMQWGC6Ndrs9iB8+kuoSNLn31g5kIN4FvERqIMOhIW
p2lfyoGp42279lYuIYpZFaQKHWfmvXCQHJn7QXWYcV5r/Cl5ETct5gd5AHccUmpi
aHcHmG5uivCVIv3mN5zVBnn9HxiDt673yMzPeSB2KwV1/JR64KtNa37TklDDYZy7
Z2sgXsAUk5dpgy8f7388iWF+EgP5NUtMd7sBn5rG+doAyzBZuxctVrVU/1W0y2wG
4z9WSU4lTN11NSG1yoZmekQ+Y6SZWT/h8Mb4r0l+bbH6f4ffftnIzgFf0wjZ1PsN
Z2ZKwJh9nTPugSyUv06lWsybU6gtPCQJgDm4bYQSCkYSM4UtnreGjy2F2o641XSH
fPKP5JjdV5e6sJkEx8iyb2JCg2W1z4peP91iWlY+tAmED9YuhB8JzqVr/3Gkoonr
rOYfCmQBq9TnuHrlQLlzcso3XtAyYCdHv2qhNkDp8GFwlYDTfztHWe5K4nnvtVl9
k3z/ybpAhMcUQgkW+hoNCHdAbMOyQ8+3Jjif+R98VBQhKPCszpMvgvEvgoRSmXXL
DYank8K9pJ3xdu6RHgvZ0GCY+GFXxiSayNbtHuDWp2gXRIEewxO5TLpaQP/Qsn6I
Pegw4dcgQwV9g+kpGg0QmyTTJQ+mcMUPgXqzwnVNJHGCwWOZVifP/stLZAKGGle4
Su0YoPqzyv0VbrnAFm2WVilvDEFyxIbU3bA7JChz4qw7URdf+2OCFpHOZOw4Kg2Q
zcMEVuCdnWi2yJvLk8cxa01ui8jyJbjjcxfdeuDPnH1O1GA2l3A7mMMAz8TermDt
Nn4k65ddtI34DRPMARnNHpHEz/Az/BUT1rk95CYl3CK3p5SIK1FWKTgbwElz5GKc
O6uXmzSXzhq5gpUiV3R2zkkQgUtOfT6NunDZymI4rg1y+JGkP8my6/rw+IcIJn5z
vw9dnuqfyFY5eQ195yvK30Rkos4I5LySsCILNwcLprHyjU+1OzVXvhDCFNWrahZN
GXx3JjQ4poxl4s3W/KOg0nsFkHQw5ox9pogafr7NAy9WRumpZ9sVJcs4kKGF/Vp/
dqnan1no2RaRM3iGikz5NheZS7P2EAKTksusOtXtWJ2LxukhOb4gPxIPt3q1VFDa
C3KXTpx+9DcHO+wyDWbxvkLA7FEx3uCH6VU7ocb4bEw6F+R/s+qpVjcETMqGmyDO
hr9k6ZNwphzSEaZdB88ZS5dX7GWPdafaf2Ia40fZsUQtiQLCpoGGse8IXUgx8Lji
huGkhUWeNfehmzUxhhNHg5u5WcNMKrCZ+0YRGRpzD1KkIQl86ZxS07+GlstPUssV
WLDZEgxKjmH+aHHogELCjKrm4CYVbkNJT2nMi/EHEXTs4sSVtkS+IvwU1AhNX5lH
eFjzmwXYvRlcRiCrllqaixHzxbKSZJCmcpx4bAnRRlinSnOwAUAIla+wMrnm/Q5g
0AqIQsBNVPKmLXidpoTnDkrpnYndxeMH9fmixpfqKQr2jmdCRgA4Eda1FWp6WAbq
sdIMuVNW9zeyBbdLiVt2cmZAl4yYJUdjUrLzZ30EBy6XXvzt6xhivnlTnv8dcCyn
Ky+Gimdsg5LoB6hW7eg3xhTJD/hMBKmBmDDdoezr5u6ftvz3ghfVstwoI5lnmCqU
lkneQlrJ+miSkB5wX/djL+yig004gyKbDLxbI6tjlPzW9EE78zd6YttQYxKym8L9
vYEJrtbi39CBQ2ntOYaigKg5FLX/JKuPSN6M7dYkucX36Zs34ymgQAZrzZqqJgXj
mfxXMM9Wm4jvx4KTZDvT44TK6IJxZgduxLphulgNDuza0wbRQobW9Md71GYcTxNS
Y+hyH0OMcJ5il4tZLX3aLT4oO6+euk5ucYa28xEdHfPQEhfcbiXV5LOLTRbe7BsF
Ij9YfTOSpsaLNEcIJmLLW3cn6LTB37s+CJEJXvMNueg9EyGa/WvtLrBWwMdSw3tk
eAWfeWz8o0q/sUITMGVLkM0+3GEPUyEVsyyBA/5bM0IuPm/x24J70gugc34iGGbA
dCnlYcTGXZcOB/Kc+tHqj0tmsRDxN8TmQTvOptLLsMpRgzBelUKvWHwk88D9Iyho
ibYgd47Wf7PCPbkYGbuf88VmcbrQ5Q7KIEdRXZBw3tQ+NsGhiwSZ7gJuxpZOvNeL
fDZMMJYL2EwdvMefeCqafxfP+6MXht2ZbuWucnA6tJeG99QJjPjN5WFU4cdg0dPI
mcewYIahHRuI6lyMzys9ZdvITkqCbxUE9tSsPxyNY3qZQQ/dZbl6sohPhD+5huu0
M3ZvP+UWTUu6UFvCpRa8vCQFZe2PphIgppVBzR8wjDpCkeDWVOTvsDtZ6H8bjUHw
U/D+guzBjxYT1R2/MG0JgZD2imnMkDHvf8Pab2KA1/mP0RVH4IA+XhIxHS+0AbDm
7XfHgEBHPCiEYqdkJZOdT5UA48CvLEBaKOpwFPlGru0rNwbVfimA9tdPPAbovi/x
oqnIKFw/2IrjjfLdSC7TI06WUpQN5TLpxqlufa8IiNTahd1iNXvdAzvje0elv0bb
bUdyL38tnIl19ZdDu86w6X+fg83vm95Jw9LESPCM3jO06aNUQnwVUnVD3j7QLlXs
Ql2qNspJMEEmy8FXwdb2XaRykWzdVZ/mZ1S17CixD5P3dCCB7yP0X/aBN9Yvk2UC
KP/EI2z86oV0ZM34hHjS7GjmWVBBtHueJluV16C/k88i5tUhX9Nb22sMXsULsJZv
Nlrp7gpBF02gUQTHS6yuXLFLpwmx1EjexIhqWkJ+53/5t3uA5VGGPgsWXd/Ar4hY
8PArPlUFI2grFCfj8yCVNdykeDY25MzUvZGmF3jUer7tAgLnTuLiGmxVx1Ea5Ori
42V8UhBmgcg/tEwlr8Qig4N0kYtaAUEuQQAwKg7n3oKsgzTuUeMYhOclq9eQu1/Z
bw6VeXo8zYEB5BIOhrBYOYJ0a3ERrjUAucZG04pAvwaZy5B4Lu/Uw1pwLPf8TkVt
XzXWI/BTMj8DUHAn4Gie217BCW5SfguJ+6x2n4KY9aJx+cvkonE4sivybXUcJCZB
1TQeG1UIxvJR3n/oZsA1nK/qSoynDMHcBHOID11Z6Wq21CTEP2HjuCk8Bub5gOfW
H9l4xkp86Kg1yga8ssPmbhx597DvKtgj4TFN7zjL0qszcqyuEx95HjLqJVOUi7My
/N8ljlbtp/PkUK5KxZ3sjTs3TWpkzgbQ3iXOIEGD3qIa/9fq47TP/A1dHlrprAUQ
mSRfE/bQ/5ppO8yg6nOZLqRNVmBNVIVzfqcvsVQEfkD7uxfTwEzkNS5no82sl5ky
iBivI5UT13CHQla8bFx137/AnOERxKX3RTE6ydC5/1+9W0tRVv1XciinAYOtnMiX
avu1ns02sQhePVQY1g0W9BYWV9u6hu3nH8NZPL3bVGIP1zic1FMHnX1ybD+rH1C1
S0bPE9HafxQ9vabi9YhDMQEiMVQF8o8+UAqC63DdMkPsnIHAgCICdpVft1DMorxU
tyHN8EkDBHFxtDwbj2ojvvoE8s/vIh7MhcjM5ksRaLFAK4BP/jvqAzh/vy2ugisg
pTnTBeyzAlFq1nzHT1JDRDCndB7KLrNphvt69oap3Zdrq/+/Xpg5vQ57isQWMh7I
ODd0p3kw+HKgAMIllEgSFiBCqyR7Q389pqlUNXAqg4BOhVC6n1tYZq5gz6CsCGRo
NGkyoJlKvMQRQBpHq7GwArPCJ0+A2XW5VdHeULFBkfgqJx8zxFDagZBhvfu8V1cp
wHszb0DvYbCBy/iaVMuNSdTCzl1+YgpbzHgb8q68WFw08JgGWcWd72FvO+JEl3aQ
ZdTQvxiHmclPWx0I5xJ1Y2xBm2vv/5b7i/VpVt7LPGK2ViecSvqgjFhH86KOByvw
t85DkhUyqJDqR98LDX5LtRKA9CdWx2wOTDiuEG25/5xY0DlaxRC7hMTRr4dEfJ8D
nCN+1srd7U1eDQt3Wh0hAEjmh5CwzWC812LY7dmgBEr+sJGxG7cxPZ27z2ocHXko
qHGua3ARTzhWC5vQuUmfGyblLcm4A0CbYDaqzpEZ7LGhQ27KnOZPyCsptl784zgL
Nt5ZZr0R5A1pIYS6RAuhjpS7ASd+2bILvq2dE4UkQhAYsNiD1td6EnyiL/mk94fD
K5hnWNBQrewgF9OOYfQgPq/CYQjH9tb02VtGLmu5/2NFooMD35KOOR22B/TKYYWu
I9XXlHilkDQU2ItXyA8Gn0r04Fh0DLqnNgQoNx5RhUv8S2n05MEiJZETJjTZaHyg
CGdddshNworGNVHXPK2xt9p7z+Y/mY2xX18QSQSBIR3U5lxDsrUN9Yl+9kMJ93RZ
sJnvhpaPeA8Va1T51KkVA/nqBa6MD+NyJ7hpuEAVjxm5BHq/wkM+EDVBDGoLZYnG
o4MpKEyhvueNQz6UaSpW/0tJxHUQGvQVRZL4B5Hg5KyE59ExLATajTNJIpAS4lZi
sPaQZvrYsKt2LdY/Rk88DUlMmwsnMTKBdJ2IaxZt8HdXwxs7KgMFLDfSy1XgX1rS
j9Jjg4DluGkSubkDkPKpKrR1EtexAJqrAGXYhDGpFoPdw26nEGoN8G+KJxGVYjaN
l1daNNDZMjWUxOrjqa3BH0SWMrxeGtPiEXjsjB07lJLrm/Ix6Yxi50XjPau5Y3ko
GQ9eZoVZuCqwHkOBMvsrb2C1K54c58p9FLvGAocimzkI3qsbn+MBw1cXsu0cfhj6
dWxL2bcTWNQCAED3eKBjPF8I/2HzfF8Cx8hoX7dRFuOXsZ1pyqYZB601sAQwX/Xh
WtfBUU+4zDwnkFpKYYQJ9aukY2n18Tl50FczwdyTDIb3hgBhcdKIwYui6N8oHIIm
RW4rZWXs99YpDlxt6d4xm/gDj92imxvvrZdld5BWAOzLG9BZiH/PXuvSzwN7c69G
4ML2zUVHxZ124hQIc4h0GSc6K9fvGxZ+ZJ/oArDCsNm1qZcx8DyyooXW1r/KQW7K
MrfxArJeWJRoHakxn3v142frw8esicdf2KzujxIGjPqnVMX3gI4vRoG2c6PRoGUn
XclMpol9nBAj0N82IdBpUrwZ2AhJZkRjEOYboG8Zc7QiA/SWWXLCFz64PwsIylST
SjAfDGB3Df7dxTBBm+C0zv7ZRdhfuTCOXotCpcI6Kr9mZM2XFI5gk+nKXjCnyD5J
xMg+C6pIukHNjcgzD/Q2YK90nHq3ORxYJsMGt5MaI7o2ARMozlcjKJj8B9ud984e
ndzyURm623321x5TuO79K11mBB0BTAXfXkXzOXukwCirBg37i/x6RL1MfndVwAQ/
JX5BNHZcCaAGEjQdEViP1NgUlbWZNWf7xLb8se637MwdqsyazuAcgP93xRNdOHnT
sBZAOK/yLonqiHXZ6mf75iqh+3ylTCvo0N75dGIbF4p2AmyU7HU9u0WaX1MPOpCd
kNc1ptoxxk1Ahx8+HCm8mBRmxaVcbM5Nrq0alVs1BiI4cjhQJMhREhvk6U7iQXRj
+GROiaI0reqqBkwrKvI8m49IRvyVFb7PIDO/9kdVfq9QtBvTIbDKkW7TaoMN1iOi
YS35IQLYeECvwKgAHJmSr+NH240Nouh3YA2fNVgt9Fg0nMcaxJ2rQThGMOzm1cmB
iudsE6sbuzgXtu4V7Sv+qpLAnUr3ZXXGMLnX5qWGM+yqQ8nJ6C5AQftXMu5nLmd2
+w3dyf4EgMdiDw4ztV2p9byivprBDEquOS+W/E+9/nHjbHYJXoyaL2D9feOsj5cL
1narir/fm45LgALc1jVOU2MVZOKO4mhgEcLtwHdY7xAovNXLqf0EEkvRtKT/U0b9
6h+MZMh/5kOFqHWypK85aM4QzhRWq8UvTmochYA/G6+f175x8feTkgML0cBzLQCM
3vQ9OTZiCTu39MsonBaYO6E602CyCsiOFXI9VXugJrc/gnVeM8IQfYmPAckjsOEY
+EJ616nrLG4U6BP4b170waowUdD81UyQAi81v29VvnDMI1NaR7Zwmb8OgmS7U0n7
V6Dxf+YvF1ISRNXC/+/HA5riVDQfiPn2bk0+ZvKy4oLkIFk8USyUs2J1lXALmJ1b
mhm/mVyufiewZBYi9Ws5DKyikyHqXFGANvJukENsUXYUufQPFTFdvWHDBy71DpKq
wQ1lwTARp/PxwWbCEv3nR5AbET7KAl8ua6lWCc2a9+G7kPS9+4BOceSGSyisvUj7
rRDAoU9Q+8NJ3a85VgZk2FdfgELY/hKc+J82UJoY52jmDBrGU2nC4K0HdcwtWS0R
gTlDVA+ujOTsBvJ29OM8fI8JE7Yi9X6xuFnKUzOpdhtGiueWXZlTHH1Tl2Ih5Gc2
pVGsNsgyuEDiUeppXMamEqDhM9NV1EfjE+gGvyAM+/PG4Lkui3yDbQz3MKC0iH2+
sGzlpg8dJtmZZ7FMMwBtpR3COkOyAWXtV7Po7kl1WvrAp/ojRR3CvKwwZqQFmIZY
qU0wrDwZZM3MFEA1Yi9J8OhBOTYStAy2plnm7HVqYEheOrgDEXxwyWur3zFSw+mT
QPf6MiO604jMnJqG5mcOcoK9sOIFV5IjiqQNY2fGjXb1/9957LuGLZ0occeDqleL
cH5YmbpNYTnKdihoXauNnFAJVuY7A4Puv7skI+SS9H+SsLNjql9tWsVagbkzpcrJ
3CDhcrlp1hP7IrWo0QgXLr/nOvm2n+5gyQvk3p4j+o/05Fb1ko0LKAZiXOKd7Z1R
3G4jDjUXqKW5eb3ujt9zrpfQL9/8A8nN85MXaKG6bkdgnXLm9Cf4LqiImWgud3af
8Jbi9RTigqfXMh2oP85tP7Qeqtht/laVkCjo76FO0g4L06hSeDrR7CZ0H+aX8HNf
OioA8q9wPNQU7+s8o0bOXjLgVtZuqE/C+g0wFdgXmO+CONWyjb9NptBlDWiWGJpy
6XYz7Shv6tYpKk53otAOayOSj/tUmyMyd2hn83eYuRsrgysNYitlQgGBiVEaHiGK
hu7O+atqxwuEy5bCgyprQFahXTwZO0EOYwPQSAEWo2x7+pfAu9cqUpxVHsnPw9jX
z2IJloWllKukRMUkPMxMlXarC4sJEmmwr8jpos+0izHwkRdw7VYhzO3dRy4uaaPR
AArXttOOMB/RrOhpYgRgjCy2t7IjM7wN28xwImDeueDD9g56qqGyaXpsbVVNh+gK
JXzkr0sBE6NFYL2EZygV9KLYM3i19mAtTu0iojMIrBQhx3Cce07UDQxDsm/gEiVg
a33EUECojsxumceEI7X5l+DVkyoNDR+mc705cky2W2ucuWdu4V8ci9Eea+xVdzzb
ptskHVfoZO2CgZJE/P1jvDa6Orzs2pBfjkWUi3cunfqlF1t1pO91I57zS2c0eGPN
JMM7U4Hfuelm0erx3vTpqzsbwa6ON1h9kZooisTYfqitoypCK7FtVqvlJ+azijyE
Dx5WyioFjfgtH7/aCSxo+l7ym5INmtObxX3YHVa91kAkEMRhmUr/IqKWHb5sticZ
HGacvtKkynYhYUNbsj0xrFY+8Id59N8xjE0MY5PzpPRabZrImAoyrQG1MbJ24bsi
jOESNwWSuq3646qFlQDIqwQOnSsWk0QEl3nrzNT7uoNM3BFI7Ij9uLb+rNW1X6an
wASZHXlbKGhwrGPAths4wEq/VZ5CwxZ1OYXfm947DpJnTOvT6jWZt/W8l3ZfOqLi
PbPdMJYgBulbCq4og2C9gSRD2Ng5aruxG7qKLp6FWsZGBb3vri7WgDX8Mv7JoUd/
TKyxJiynHGUseOweEIAhg4vWnkjBuXFl+STUZv9Kb8xL5NIloWTzM+GuSyMijCT+
r+X5q3cqA1FwvMOcHBqJJQGlL7ALambyfQ6njA7hvjiu7aQ1yydaG1YQ/sZUtNzk
Li0TEujxTU6YcGzIhxOjfoiumWa1NcbWsyUw18+XqQ0QLr+wtFiQU0HRJy1ME+13
FO4TyW1RbEhsMQgRLE9SXFvI0srmknUHccoDElSS7exbSKPxcbXKVfJBGk16qzr0
Jo2nT02OGrdzhzFP2gUC5sLbOT1MbfUuMv8Hhh4gbTEpP+wM73+K6GRFWznyDEy/
mGTn90O2/yHN3NV5brg46xQK5H2r2FTdlw8fHwdMq3X/U5p7bQ09p58gTe/oYSU5
yY6cCrn3BnDv/EgS/tR8od1P4jRVVANn37ErgS64OQ7Vs77blDS4/Aysl1vgsnAn
rq0FzEGuAPaH3VCdyntX6l95kbwEFqMhv8/ie0KvzhguUO0wq7OBkR3hc/bgMXAS
wiIHLQEkYHlNstMjhLeOQefXDbKoe+wLEOkGkm9RTp5dD071pDNl+eZQ5mBFO1Ch
07bmJWGe6lZskD4oTchqe/bqZUnlLK8IQiwsSzdJ3elR87kcGfNh0vK8KHFM1irx
HDoJIdcG4zFMDCtpHvy25m7aWodhm+8TLhS7zOoNMeYhrScpcoN1+vHLJR5dFf+C
RNDXY7yafou2PIT+W4tXHkdO4z0CX0lDDswRdR3dGptQnDJC3ku5qiSHvz8InvS7
7a7j1hbWJJVij1Ey3apMmxiradD1TyRkttJ2XyxwzIAugciV+/RWYmdfxV19P2pf
Tt7ePxt1dvrvsKjpSDwAihLmDEc/9zpWc3tynbDtFUKJ3z8Qu4ZluTtfMKSd88v/
CwaZLu7bwrmRFnsdpIor+QYAp+Bx6mpVsLM4u1sTvHEd5iqcQVsHL5OlEJ5HAXSt
AtendtvMq+JBlalDCJVUU6IUysuNtlyPvtyQeBGzypj1UMpLI/RLrzEiL4pWEHJS
dtOxC5LoVbjnAPcUh3KafzI3DkzfH2aMH5rvtY2uJtBjBSY9sqrNAj8I9oeRY6Sk
tpsrcXtLLKL6KQUMRgVdv2UT2rSTuQYW2jT4QCS1BaJ3IOj9m/cGmUv05uWN4gQI
8gOE6kDqcnX4P1jMX/jPVldxT9hIxFddw99pAI1KH2T22UC0TsvgcIcCV1M3TTZB
HCym0AraHPSAlSoLFUzmNE47XIN7Ckjnvki9ltJEiHp78MXRJn3RESc7UlI4FHMa
IBzKkDEYVMIuiPgMJGpOpbLbLuhl0NdpJyqwnvWGy9iq0eXqvaStoaViT+Zf/b2z
UZMZO9laE5qvXEXGx+kkS6nMSqp7p+ixS3oKvt40+8dvaq/SADnCbtIGLuXWMYwv
gdHKGrgaeJonEajpGst9FkRGsbKgjpucA6P+kxIAhGjQysJo8J4Y5aN/N2RkHGmx
9WufUxt6ovMX050Oo9aMOHfOLE2bET/3EQMwzedQ1VouXgtoHFr4Q5gnGOOEYoap
ycaP4Q51WKQ6POpTXgtUmZz9zzv6rMCULmASmhVWy0vkLYDCwlxJxo0+ZSPAV4uW
n1XuLARDzpaiGSbmj0lyFiq+xzVub9jgy15Dl2IKkS0XAQNgRqFkdHv+xpDCMgjT
dST99CguJY++j7uv2YxP0Z6Q6pR8yzjur/ZN+wWdIv57KFALEiCaDfM+3HOHuGji
gxSZr2k3Fd0Hd0T61whyi5h7inM1/IsJQmZYZRxLxU7wPP8nf5NwdlsxIq6d+h8D
xd3d/+20cxxH3vw14qrInSXKXIwVaiHR4Yen0srRahY2rlcN3PytRng64yfTDizW
s71pQGd1M2x9ZKFRKsL82Sw18Ulx9BJTp6GSJheEOC443CgXuZsk/aiVbUIWZuqt
Q7b5wBrC0kYs/uX+RW1Y/RrXlky5Ldw8zvZoFocc/89JAVHtiXnvvAV0Tjmylmcl
LFZGRlyRGDkOoyxyYgSlEgeQqwcH2ADsPVjm11g4PqJM+3ZX9ZkkO+xYDEQPpBqR
C2N+wA7PkrG1QKmRTqeE4/yxdzpsV+5Wi9OYzseZKVtzZg0drX5Q3TNNxztDOwXx
l8izhgOdCdyVzLOtJlT0/+RDu73lKt6Lb3OL5uqN+I0gK4Do2wmJaczl1ImIYWji
MzCWcJN1+cv9sfivElDHGGpV7HVvMH9ntzPmGVrPQuPpsbCLRTjDj6bbr4eEhBXN
ECMOKNP6bHn1zHh/aZfldBTTikpsU4LZVeApKglpaeUzWdYiZN99PH2tA5zzlJuc
b3Vt1t+JIZyr54t7K2ICQb345p2DPn1/11kd4t/D6SCaTfB4ZeI/k9JK5PfR2mit
DbolEvUzwEJ4knYE89ilLwNMjbLXymP7n28SJJ8JX+YclMy/Exd18/Xjr1281RnU
BtXvU2idsJzBOkgyqzKwlQKaxTRpS1vXF0pteZJk9FIaUvrdjLS2jyjt94Ue5USp
QYy+IEEU+wd9/Gu4hhORyrgudPYSToA8nB5ZdtZjFTZjHGGWrndR3ZlfeupYd5LE
uxgO2wsL3HXraNpfGr3P2ri3znQ6pnyjfKW1A2xj41+kS5ugbqcqnQdoa35+s/p6
AyK5NWNYfjEaEf6ONEY0whXJNrLkhpgUIFm+sg4ctw1fliWOVzeKYfJNVADwMYEc
2LPEz15MKrLxqdG/gkE5Y9smOUyxMUcfDYZk+G4xTD5ywpaqOwd5dereJl+uf6fZ
FUm28BXbQQIpiIVZUWFxTSYEamm9D9sl9Zq76SknMs5pTBMsJFJbT/3Z7ybHCaGp
L+usNpt3xrW3pIkh34LU3rXCZtBpsl6Fb4yYyUp4f2/1IDZ5+1VctAj0VcdpqPEf
yiG3v1rKvBBCY6GPGMxO5zNMNvqESgM+TLrj+We+6ru8nW6cZoTkNRoZq+XxuvTC
eFXOPvl/A+Q0JH3xCFkB5bXT4DYdmcjsVGBWCg1xGxkETM7pAF9Gca1rXLlpZY9z
3XaLDlZIxf43vu11uiJyasOcXTbN8KkJy+7R3h1L9e6WgfEHDSFW4gzDwAIg2b7k
j974rt+nWjEQdwqZGZesUM8coc6stVH5M/rJbdqeU8xNjiAjAFogWq52/rObJQPm
O5FgjY54UDoJ4lw8O75QR2iT/jKIUgAPr2gt106nzV3TAYyKwwoM0ptiEMhN/xaV
8DNJ7y+ZLxn1N4oiVZTjKnmTdeD5CHcig5ABjMWtW7h88CTDuWsMhHRBrIvKgl+n
75I0CkppdRsuilN6PdaL49dRJCee9szna07FhK+LED6wQ/Nt/+dmZVqPLMWKurBq
jYO8jSOEexZqv2oZ6XJwC8ixAVKqfzH7VXHiTeQmH0Xymi1nhKYV0/E5hXqnuiL9
0HPzaxjNJ7750vbp6I1xGGOZUculDtA9tyIOmAVhwquWf8r0UGKAGPfXCSSfNI55
F2/KOPn5flsxqGueg7kI5bLHpsUjTyt0/xqqaLyO6W36o6HiTEBwPOmM/yKzN5k7
PMLidzoK29H21FTmgfewG5v9ttL3zhRDXKa9T9Fp0ume3VyOi/AldLQgGQIcsdZG
bUHEuqEzuSg823mP3Ujbb+JnZm5d7+bjAZdggcv+HfSe3q0Y7W7LcZLLHwNnM9hM
FpJr+F5Gf7LH+sE3Y7ACTfQATvNdV75aIr0EsrMBYpBVaojb0xWU4VSjZgU+JSlo
K4CZv4MugnGqdTu9GWCJi1k59yAxerXZPdUIxGw98tNeLMKlQcMetDllBlyjGsYl
G0GqX23DHNVYUbPuFDIuTSljBgX4MgrdeWI24++gT798X/ujk/5Y5pg1G0RVgy0F
M4hhbABKZrbxo0w66uAPhLTFdQTEYh7uA3WEWTJtR8shD8OMjocP7GXr+VthRzyb
0UAD7jjeAaJLBaDlp3rTiObVsWA8BSvNynlijFmzIBB3b92GNz+ZKjCb/MRn8wbl
i1zdwImIABrzO6d52WpVeQTWAss8rQ2pRnUQsLM04bfVDFB+fBF6e4nPcMKBjb3T
JdhK3ZIyMoPgVWfuGqnO+ahJ1JfD+oqhUMEsXD/ZOfBkNaXF73uWNrL3ed4N0Vm0
52zdPboJ1yLnu1BH6PVBMRRT6i3hbHclhkyy93FkhweepVNeR67/6UAxivdt+czf
Cn2rwqC4XLRidPQlDrWrX5Z/rJKIbKZULcfsiY6tstdfvPO0XwWsYyh0h8eWKg/b
4DzWnCQlwqp3SAEOEMnmKZuw+f7VihGG/0mEUz4uQ1LtkSssdFih1bKSMNLcB5Yz
WtHoYPI2OcLKWWoXG2sZkowFt/BdQmexIzfA27kcqNoPdod+YuDlEAD8u6GOifQK
a/BuPTjCncyf6dNgBlkff2chqPJNcKB+uwtl/wEEyEAAZdAu4v6ul5HuEsE0nv8S
5nVGIgF354MPs0HmJ84fu9v3aA9ToONC/vn8dzViX16BVaOPEsrRCYC3uigdHjrb
RQnP+t6rFoNgqWdKM5vZGcYlnM+IfVQZBVbCPWP97ZY58LQPQD2gk7+ii26+AX6X
/fPd9j8Y0cIXXgQV9nydD++w7MfH/Viy3AKRspv7E5Kv4egFWgjdwrjd2sNYUFSy
zSc/z/6mOfVilHR64oPiOH/2Cvj9CCeqZPPSHIrxLzejKQ1MyxPWhnburtbRr/Mo
P0rzcU9eMgKDxvA8NIvW8Jua8+t0BTk+yyCPpZJopDG3D9GCB283CAQK2kpqGCpR
TR3nrSUvqUhvR/0Nj35PdZz0KyL2rg/Nl2oSINuYNlH8276XGhjVe6cl2QBBGnPV
nfvkFB1iTUFoIi+Lz9JJfsqCPEoHr96midahBzY4rueiuTNby4irVWFzdtDGJv9W
2PXlk1v21kpEkpeZQ8ffjxYQz/x+Rejrw+/1uEjz5699zNkNK6w8WykgO3Y3O+Wq
pC4/jn/RjXRbLXSuxOEag1DJcOGOYMuz85zvvMMdLXeKu6GSnpNg6VbkmVyz2qkZ
x/L9OpHEuh7oqOrPshgZQcVSrl4Ub4kxS9UTFI2/Qpcw/UHRvneF0bTHadf/JWWK
o1cFdRIpdLutXx28roswGIL8y7bYMKmf7Lsq27sjaFHl5Fz2k8ZNK6gdIeIYVyU0
scxdH83PCCJXNX4/fkPViL+jKEaCF+tzqw7d0rO2rulGnuBJj+4/80LKk/3fhJ2i
/naHXKQ27/50CrE83gRFefSEdDmGEwdRbYzDNJM4bhEFIkGkC28TJdomEhrMc7J9
dTi+MIY7ovmRdMXS+K8aB+rfczZxSLP5bpLevGrtZQTtUBbkhHL36w6ByHr8hjOc
3HSNPnxZNSzkQ/6F34L3XdbSv8nxbfLG8PqXFP7D9W6r0Zrzd4K+rmImrTPn00lA
js+iaKGpR1agl8q1J/5y7+G0i1gT07EiZu5/AUR0kvsPvdZUkhXWDOMQsPpR4H0H
pUIxLloMKRfvXmWj1OJGoKjgW9/wzOHsZdmLs6/XOVAKWbQ7U4NC5KlZ8grXbWJb
sTCTJ0W07w8qQiN2gaXo2WKDBFXruOJxfEk9WP22qh9B8CPw7jbFUrPf6Oc6Ug3X
oVwTuT4Z4/EP5cEJqa7UVN5DPOAndt8d0yq+tPJje3dlaFtdi1VXJ+qRAN6z9dci
SbYEUNoSBj/Z34IAaoUPGOLn0NQ3b+jar7TgsgA9087XFX5fXZxyvM3ByOI9sKmz
sqGSpYQ0VUhpBviDuC0Q2DLfsrbNr5KV1vH82mlTapsPI3TNlxb25DVZcCcX7Y9A
7e/LgeEiaOOjkzW7jLgs/jMwEG30r0oJWpFN+4IJxNmIZd3WnpNU9TBjLnMvgU7O
WKsFTTDo9FGXq8HyWm8S8632/58nbhIyvh6T+90QYlpUepxPmfYv1sJ9f/mrLNsx
YfIE/jsrTfxO96Qnxa6Y8ADK6nJjnNXfqqqmlRK4b+DrdY1BSIJjxvRYt5dS4CDB
3rr/sT0XUq+fKvR9PbvomTfUIN09NSeZ893NXfX/Qqdc8DbAFDmpIdINw2F6nFjk
SCxJqm45ImtuOqF6PwxtZmiTHV5ngGyCT/O2CI+puUM/IOvaq066G4yim3USKZsy
GkF3z/Z79XwInq0nCsYQG9OlZ1Bkilv7b5Y/Yl+3NFA8yGmQFggAx/UURjD/6CiL
PQFVSGwB+EVavJ2IgXpJ1gXR2fnAF7zgmXGo1qWSzIVfZT7XrgKra71FTgH4KPCO
MGVJVkMpPru3NbCu5NV2xDQR7H1C2VwkJwcGAtWj27S65Mt4fmO5fCnuMqOZc48b
dyQOr2NxIqJnDuEELI61TgTfD1xqL+9BeO7nIb3pMQJYJD49ca7/qOQoJpxmHa6W
Ccv5cvfV0hxB81Re+O96n3TuSaYX8gX0wDwj60wlsmqGUpZ82nScf1iBmgrnVfXS
UwEl0ziLSmouF0WPlZyNVlLpKoQzhwDQSD3XEX7/UMUE/yyvmwqyewFUOiyaXOS3
Wcy/NiNOwcZjve5W81NdSmxk5LS1wizbiARqqYROhF6NsYn7nP/hJRaF1awgaxXW
ECYGJuHtjAvpPPvD5cmklOCq1z9TOowu6XWalCe5qDrjdMWdQ8KgL36W65+3ts8V
FlbhzNdKefBt3X+5BLfw5mop4XGor9X9lfWzTHV2EWrqwiwSU4YgwcBwkhfnOd3x
tLPJyqOuX2/Tz+s9rHjl3DBCRADS2OU04KZPwlXV4ceycbUGY8Io1ic/MAUry55G
HZ4Yr9Uq5IBjxTbYcTkm3+Sab948qiFjpOCG3TwohuBh8k/KPMdPUsEfP5hBIHq3
7/jmks8pqV5AjxJQ3zDw+uF1fh4AlmeajMH/C7B6HGK/DBRUc92obTP2U+wMcbu5
d6H2Svqn0Jnr6S/4QniHPwacj0MMOG5iao+1CDEF8Ot947N/5ZPZZ2hUXvnx3Ych
yzLbCwWWeWiVkBZTSwfx3r38nZWM3+JeOY3GcT3cNwgkXv9URVdG7e+xssVe7FDb
2nWaEDpUOo9us0fxb6dhholiShfluvYhvVy3g579zeJYFfnPJVtqLX/oZJ2C3E7u
gtlZK2ZrVUq3yXbBLS1m3ZG7NNneUsK1byb/AAjGY9DTSHbxUvXWsM4vuV1I9kGv
4TmpQnPREbk2kwXxcs4unBldbGOpj1GvXWAZqJJ5zlsUnf4IvzUlaQ+hOEU76hBo
TBdnD8hfoiSmu3JDAN+FE8SBRMD4k4nYR/LrfRucDIhCsgN/JJxljPP0OJOlbgK5
Rzg9MRlrZO70ECiCf/slY+4AoluV0XG0C9vwZ9YHuHDnzd1OnIw80LTKkZqsPft3
kxZCiy4G4wy5E39d5TwsR/FWwvvTLTxdOl6vKJDw1lD58Z3nR90Ot8MxiZJpDctZ
Hy5wXzwjOpvqPfatC3bUlXCteP5PqKCytv+iVRO3p9b1EHjOClLQPAhFrjZmDyf2
b9A4pbptknQyFLVVYn9IGWpE8Mphw0C6rLwtMUg4w4Yohv++BrJujHiStkdXRJGF
UR5NdlgmpRsrjFUV5RuUGnr9IhG6G+AwuhqmVVVb6UnEfdLZCYmxjDg+6oBaLwBq
AQdu5qFCqFRnNCjV/LCDP22PwEuijbCSWJzMuXW14A9/Ngc6AbJVDBgwAoWnYpub
6+QqDkb/HQzbiIdv5Mw85leFuhvIejIr3umOXz0qoPfh9syAQoF/QC+DNhELWJib
LRxuW1iNuXhTPpUDV8JtwvFSBAC6uNAeR6rfxEcBCX0L02j2Z7beZmBa32nGHWtf
FvKugV4eSn7N/OZQcn2QiugdF/XQdlpUPNpaG56/QFldE5h8GjPwmFdAiS5KAfTg
lD0UDm/zFKDQOcwBScocfW3NR5MXDtyU0qqiCYwnoW4RSge05cK6k4x+Hfthk1N+
KBZ8lWxwWJFsYRk8Yc400YAEZ3Q3uV1A9Knj/4btG3DCFMo77J8mJsyrtdm2Rzez
uJlcOAmYymQ+4f1NTN0n6Rhs1guYVWclr5fP3UUByhTX8A6Io3ivgplBM9PqDP/1
R/KQuteHNcldn8fsbudZ2g51MmudDYBWv+FZw+yM3smJRtfTc3FZAoXP9tl7Rtp5
MGg3T3DhjmauzVLlaV2kwx3txuZd3Ytp6uD+xG2TbnfBddPhrAdXG13hr60nO/xL
UtVI26KaWh90hoR0uQfelmYvMOEl2gMDjtDyHpY6L6CkrMmGfhmYmW+3aZtiqNd0
h5uoPkLiW8qkcS+wIxd7Kc+4tlgsuEnYuvNG+Ty2nLeCVrfRlHohRV2xDZrEjfFL
4lqApeZd9e5/YxRwBY0gBgiCvLplLB4hEtKG1hQEeVihEMU+mT6tDI0lZFP/ZD/W
W43ra8MMZW6QqRZP7AdghBmRIBed419lx7t4mDUolLXDIe/JJGCbzAYnt7GH0Jix
q+DlGMlxCb78+Da0RSf7aHJ7egXTkS+WflHFp3CxYjaSxqlpq4lnd50pCe+8zIGw
wtxM4l0g1fG6DKb3VhZhcuTjMt+KAwuVXMrnYhjOUdGxmI5joupz3PXAqAvgsLQX
q2hEKZ0uoU3PRgbQhVb+ECwnV7Q8YnLzxT6ad79poE9MtFrPyZXSBqNPYFEyqzXv
8gAa4V3YQE4rk8VnytAGJF2tNEi7N6NplUKON8m77nDoDAMO6lBQ2Xd4lrndsk3c
T9JWx7yoiSUj6GMnJzh8g4RVaonn8ywXTmDJtFQBbVkFEMlw117SgRS5UxUngc68
xT3hzRi8kzU9G7lunqhFY4rGKcKelkRA2Ki2fM8xlV2dLaQi8bGIBzSfevUSLcb/
nqP+IGbaZXfXc82GB9pfsd/qOfbbLoL3V/RNuNllmcpT0MQJuY9Lr+GypjP5jddP
jPP63SjfSW2ygIMwIePAxpGnlxXSw7QoL2Q4RgkYc8ygC2Oj9Oy6Ktee3l3o/oXI
563RTVQu+4H7eU6nb7kwA4uD5YA45itBrISfcwla0/ExNFzIAG5uLO7mYJ9q5xxE
tuDw1i34dTTmwJ7b0RgP0bsii2DT2wE33wsE1jax4/I1kZeemIilE1j2ATAvAf6H
66mqEf5n7RjlYLVPj1W2/JixFz+XqTNzT7UyAdTpAlLcJvLUmbVMYaEfLts87Znl
PIuvE3q004JAyeFyIroJKCpWJt5c4z97Tp5Q9XKyeYNISORLHsafs5Mp7dMjzBBP
eL6umEsJBYR8QAZrA5AwlktMXTOzTjSTsTP1RtJ078jDfMJY/gK7d9DNQ35SxMvv
Xf2d+ImNvm6zaJ8NTl4ASA3jopZX1i9I6m4j+Xp8SOm5szB848xj3QPWfroX3e8W
N6BzCoBIE4VaIIev2qiiv7LjKue4vqCSrmra7YxpXVd/mld/s5LD7JYxvV08+vGO
GPQUga4HY2EoxiCWewg5hb+MBsU+e73C4/eOB2GACIky0BoD9NmHQND9ibEyCOYv
Y2eo4cCbonXGjihz/8zn5waHbmUCzScQ5ywRCr59FwPlTVewyqDdZnTwYC5Suaco
oSviiu7O7UFwZciPNX+qEsus/JIH14+7LvQuxV2sWfa7+Rjeeaz672iPqfyasdPX
HT364EB3caEhhQbsHQXcggvy63/xFWEOFOR5/uTQh4N8jcle7NM9MWVJSMlFukG8
OBaUc7m1n7c6+u+rd0qhuEWizWfnibEZAjLurHAgTEqgJM4bTBJ2vsaHaCRVA1gn
Xrc3rKk08ouWWfoYXtUxmBsVywtDdLoojicspZ8Hfflyg7/2r8QHk66FJ9vdQH82
5Rn3+WZ7DyIcgM39UZfoaBYTSypYh0cHRXeUv6IFf4QJ6udWKZka/T1Gas/Ymz8o
0E8JsCIwzSt2Rzy4d0Iyv9XKDqnJ6KiZL8ETlTJ7wySqKJbqVuzaVNnWkJFSPPhG
S4HSVeOkngW+1AzOST7zRFhHaFdKpXCUorpwTDcp7woYYmxA1u1Zg643wRBKlHDY
hsWmhMyW0fBCI7R/jNcbJ+LoRMyt5ba7g4W2XjIXeWHTe7VO0S1He7z8PkClfLSx
P6l+jTPtNAsaR3nwNORMJuyrT9VNvgSJrYLP4bC9mT1AwYUwPmo3vjPSelizt2h5
wt0fGpQOHj23L60dlgHLDWcKLK4Th/5jMZg124SakRx+Y5zfgwZs3jmUhNYOM+Ka
3peB26qC8WdeZ9dvhFDxrzLjaniFqmyr6zfkC1EGZTQgLOrXWQlX3kUd/vLpm5qG
wVs5HxCW2IgSmw11duAfW7/NB44gpJx8pMMRncskQmJE7vZa7zJyaV9xOktoNlvb
VcPjICyuZ9SYq9rsfwmHRucR+c5S37pvDW2Rd6epknfmoo18/Y0+eCAMw8YMhQW+
jtQOFqSfOdBHQ6Ukj6Ritn89j+ZjRUc+7WcoT+U18P4F52qk95IOMxQVhDJ02hVA
/Ru+6fgiV8OpBwDC9dJ+XNQX7zZYiG1wXblR53FLXNWg05zx1JDK0iVJyJQvPojh
teLXjrxozP9BadNoPfB1EW2ldAi/KE+Yyf1Li/cTZPYkkKTcSXPIck0YUx1yLNnc
wfAmkWygIgYeQNT/PgxYAZR6Duz3AZvFmK9V8aZYiftOs2xBaCY+dCSpJA3y59zh
ApMMvreGExPQMOCg0McKREJwf95qVqF0nzAdh5DVYe4R/E36W5ndn71jrlRXGrKr
nLQ8e3JWxUc+hNSCVgfzJ2ZrEoiOfqr2zDnLBcRijPA30bfOyLOuDuHzn52hlmMn
4nRa+7xIbjFKwueoHkU34xphaMpHLCPtX+KhLchdaajdKlzD0F95HBSgj/fWJp0o
wsYIynykfnhnNraCdbEuLQjbLQhgTOB7Vrrxv32iHjbmIOBFIRh8Ey+7Y3ghY59i
LkxnGpytSPBigiXNGqTajP0G89solBQqp03d8Bd1P7bS3bR1xil4uTO9FfmlY9U4
LOBpYLco2ZC+U+E3pcdTTgyyl/ELCE2G9iRH4XpLLc9i/z46SG0/9gTgjtVENSoI
nrw6meCdBqGs6X8dV+XH/25uiiOEPgJs5xPAKSmJoaLoq8jeC7gROFzmhBH7tjNA
yPrYl9erDjkiugTYD0ztOFYFEo87MZy9frAmgyVgvXuzTr+4+RfnB+CYY2vxCGsk
WoVGMI1rEpamrh9NZ71aQEO4gH28ZdD4T1/1BSdBDY+ztzcPG6mXPzvXWlobIn7I
i+suoyjy3jtiSNaBdwhuBqm+P4usQRuikMjHz6WJ8wo4VBkutw51kRnn8pyB5FlC
s8pFLqmZj4sL7LyT3vpIy9Cm/R+2dfaIum+Gmbz3xj1Mi5hWf+WuWsvG7yCg0le/
4zfdOhqEdqwOEMlgboPuwNaI3NZy0R3z7ocmuMjz58C0nu7i1C5h79MLUWF49KtZ
W2BM6Db8JkEXHaqFtbIDJOcULhTDdZP1FOdAgT1HysZjKjjyxqxnVIiptNsIaZkT
5ESq7Vj2vKK5JTYSl1foP/u5TgTCKRiuoFEZ0wWK9tsIbRT2bSxLvXL+alcaX5Z7
v79R4eqRxQlDyZp4HlBaBXBiV3+vu6o7ZRZm0R8rhyB6jg44P/6u/H96bAjREchY
3m4TOHW3avoBDC9on+SsHwuGeBOD5IYL/fkwDIJ2+rTbl1uJ6EsL/s1deh9AKzUy
gO55PxxO/b+8pAf6YD+lu9JY/4ni6+BL8D5g/QHnEobhefuX11DFLeh6ynhZ/ycs
mgNLcJkoY2x+L8bbNzbNrozeLM3Mz08IbDJO/eX77WLQoAbjH1AcSQclRCeDm2XV
Ir178oLEWqhs7FE80N7rWjSpu9TlNQcMvL/EJwu58tmlvSMUkQBvehA0DIwkdkyg
+I9wH92Slh5NxaGSI1O+opoRysvC2aKaqN8zT5jvtdRRTwkFi6YrZ4nB1l3pWMqm
LWESxCTCctuboSNXt53mw2kV6NNaDVo0dC3/JTW4TE+RYSiLJeQtysBAMBcCy6fW
ZciGO8uiI1614g5E16T37OrJQCY94zZSeKCF9knSp4bjCT4kfvWZYJboiuJcOSID
ZAKZ6Nj8p5pUYr/pJ7Qi2r7iU8VDAE1h1mCzd0N7hMUN269OouU1awEowNzAeOUY
O6Vm3JSIu/E5KMriv7Rv1AwIMx72UuKRU54Toy88qj+pYAjAONI18MSL3WgkoaIf
hfZrXlJK1FA36TpYyQ5cfAWcjbn5IjqG+AYXURDi7asVoZpDifX77AUUHEtIwcmI
ZPqT8mePf4dpcy3N/eh94jPtgLdji2q/sduDFnAtPm9Q8zpevXlxL/Ly+SxbejK6
9tkqF4712DeeMOR3JdK2fvZDMZuaF3Co4UIFrd04hqMHoCdEShq5GlKLhCfyNLLR
AsvSfKSLcPRkyzz2CDrmmpDs0l8rY35sD2uW7T+hiO/TcgKhfCaxUBrlOY/5pD3g
NWmCDK8sQtzUankxBHKWzjToJRSCYvBB+b8oZUkGRDtv0HBZ2MdCuL+OzoC2UORL
2B8Yj1ySo4bD1r56tiwqKyJhSZxQR8tjlXwe/3PUkfrWr9ltMWGqj7dR0KNJ2ZvO
qapl7mkvzmRlA9oLaXwZL86PA0Cqh+sxKNa7yJ18NA8PJRP8mIvyeop1JmrUNXZ3
ONMa44NIqPRu0rzRQfM5onVNP+GxFmpfeRIM5YYR+UimASUg1tC7l6eiHhxxBYtW
jMi/arjrI2hFDcYET6t2VuH1JIMl67qzQJIn84l/xFd7GbQwfAXw2JREE3mDuHwT
tQuYbPZNTlEbLiAeh/It3UQT6sdHYAOh/7is4GrzBHbWu+NMDkG1vvGBkG/46I/u
TbDuzXN/gTIeEJcjIhIzS9PMlk1Y/3Vda9B3tY/ig9h7CCKsovlAiHQ0UvKj6LNj
mvrLLnW7p13yhBjv36RSgE8PP6PkchGlmOjA9fierejBgN5hQtrW9FTxb67uPmbP
EmeWsD3ZvvbZ/D3ebN+6PCTAvulLhtOU2D54CejPvT2sdlu5H5Yen8mbpjarqhpr
+GDctqMxbFquSYG2hFtMlium9YgtqRYKDXyhHaZJLkrsuci5F1ZchpOJJmxPUA8L
Y7BqFjrDCKnFtWIZWf2KwLSDytJdfk00TEuufVyyd/pjOuc9A4l9tNvTg8nDY7cQ
1BS/BOk5iudXXlPzZuFZnqvZIrdUZhP/pk5/+aZpSVdB0CUDvkKihhDGrwGo2wY+
nCga/dku+9ceRIe2OYOTNISnRJfrbhsT7QJXk5erRtMnUVdsAIShvWzaW+PZZEwS
vixGuuS3K5tJMEk0fYYDGtXHdmNLLW/63cOWw3Do/NWBZP8vUEc3Id9p9RTsmTvP
z/JI77pVHkp6TXLZhQ5v/iJXGrs7WPUvtIZxSB1mqeG0MkSKshWomkkOrR324VL1
deQvQqWJjhfY54NcOJQ25KUtpE9/7XUMekBSuFnwAnbtBszcatrDfKQdP/fKfAq9
fFPJ6IAeZod2WglvGlgb91/WyDoLk6kC8FPqbrtqOrrkEs+P7xzEUP4pj55QMwvO
a36YRbUHVuiGbMTpRUVwMgZSMWrKVTdPPoks0pRW8EYMNGfT5n3VcLWd6kU2YMxy
fhHbfxGR6sJZNqWzyXaDMIES36Br/sERX01k0yLjWdL6phlrncN7dkP86pWJQ6R/
YaBL5Qec9jB6HL7s9oRSeWDvCuWuhjEL6cwlTwD0qLTOiirj2oONhcw+M1E7hceG
iy7qBz4FzWZOL3mQ3J0xPi88QblueWB307G+hXw9QwFeirHlN2HkHfg7FbZ4Dg4i
WljLdMMqyFbtTEU+TBZ57kBso75lzxGhta+VmcHCP2ZoDkdmhI65i6EiBNDcwkYi
0IyxVLNML0yZNWAlIKF7Xn8b5WoW8+JjLVWTVyq54Tx3slQG7TWiPY0rTL91Oert
K28hazF3Pjp9Xwp1/Cm7Dfn4BkoqRVijzULDnRIYRCYBdRZ4vGpGAdkOviAWXymS
GRzEmAIx45oTOTElfLw/zr5VH4VB1DdUfUXNEuNnjxzsUJ9keZ0E9mBozkq1AbWM
zk8as1R5hAal3SYHFOHulIuxjsToFFqrnHw35ERRBM3B5j4fq19mQP4KO/5a9EYz
QnT3lMjBXmp1tFoD32zZFHdfdPaAsOoG3pit85i89VqHOlALP8CgRD/BDcfgZumc
44QQNerf32ZvWPp0ozaB7u/j17ifj6UfjA16S96b2rr+ifhX0shHpH4e08hE96VG
SI6bm/0kHXRxR9csEXpkHO7WW0yiLIukot+JE6ZUlyP0UOChyWgQMf+qLLyIFa9h
gRnMSLwgD28Yi4v11INWS9fpcbilg1d145d7SkE0JX+ZFbI580MVCUcqc8Y6by55
HQB+e4MM/FecJGosG9j+Xvj5y+hNxjARP4sCepEu3mpHULZzawuilRz+LAI+Sf1g
1YgjxktDH8CjFFo4Cy+nKjBg/A4lf2hgONsIsYF17ieQ08i4j4IMrfxnr6xmWJZP
xWXIJ49V7zMJXpEwQUG2LkGILMn9fEKXjfNyC6HKdlPhGsCg9maVk8q8S2k6Fyu4
oRRtss9pWZH4pI+Y6HP7SlGerkveH2CkSCtRVUzBxcPA4Gg5FWOPsldOhLoWeSeZ
yLQGHu9ZOvS+80K31PwyGVl80Y41T9Bb8mEeJaUrIixQEKgCcC1/5rGzs4SPe1MG
tuwTbez6CcJNooDHyqX1hF5XyKjQ05JXxh6Z+mnOiWTqCbkpttK/zvoq0lj/V0Y5
mrCQO0I95WObqdQ+f/xcTC6OaivwOJdli3DjXd6RWrWMBMBEq0SBK8ZVKsuynblh
Xo/gog09YvEeBLEo3LsP0O7UyX9BrW9lRmCKnaz3jmFUSBmkcXiiJBBOxAvWaZAm
wFPsWxv+/ExHVjYbtckd9avHw5ARe2m0TEme4c61dS2aI/kN2vio/D1fXwHxBdKm
zn9Y9qnHU9LGOsCIV7TTKqWPBCuJz1JQ1fOmdqxrqP72EWUOOGAyH7oujgiECfdq
Nqd7FgUISOuLlrn9NnYIVp8/sHlNe7w4djcNG76Q3O7hNL+pmJU0moat7L1rnpAp
kFt/7Jl0ktIZSYQBdeslUw6JaHPUCDc/GVAXzTuWpHCZj1VNETvyHfKl2BiCMm3r
n4SsK6wg9EYIXuPBBr25ohn2XvwgiNkKJXRxvU811SynD053ZpflPnAxW5w5lJHO
EKXI+oabvEwfhkmhNe58r4PZOMNF/Dp7MKQYYWZ30or04++Cru86sXTXuf8R4vQ3
7OEFNBE7AHtX8IilNUgoStehikL/rNklZyOKIyX6T7WTTxN1TJefODk9wf1LL/8l
hkQ01QsCFPBtZR0pMJIg3r0abzN5H4s3phv42tBL3EWTovapkDYRC4I2Vk/Sg6bY
Zd5sqyC2CV91FoqGYFLuJst8t32uEFUeLvkSBtKrKKzqSTnYAXRf52nsMwXE41Ft
OaIjbcilE1IgI8PUimJBD4MYYqNqF+yArhKa9sRsQbo8Eze5ylqBPfj1EwodMaVw
LfG4Aw5+NSs5GHLGdcoSKXAK3zrxM+Eb81AGcCUvW+EzB+uNtg0BCKPcgQOf5DhJ
bnQ+E2EHEVzifya1HJcnrgdrCzQrjePwCRIsyKxNyxO8gLAYDuWlO0nVuc4PFQGR
/xLJwLnTbM0VcK0Iy5Bmq/2nOyeF7WW8QCLUwVZ+HnPOvJwTL+LYcSL0+m+Nb57B
ysO6SK7B5xCkzMB2ez1jhmhX5RBkLuOLHJ8dnGE5IFB1P6t2ZqxX73Gr3ROa15aE
h25RSCtfEnbLQvcyYjSTx1QYWoT/s/DscudU4SAUlOIQ9YzLu4PUCJPzaM0oFtdg
IP9MBMsf611z8GqTENY6aKjCVtnH1QSllkb6S/kWbOCfcuieTjLKAvkQWy3nVDpc
XvmMVngWP/WH7pQ+6SHxqg4snz+LW5gS1IWdXVVy7yEFGrA5cBqViWMbytBFbApT
rqlKLtctlLnMkIVTfd+LFSxzA+V7p/hNNuarN4b8bZ8tbAiqF+I6/prASEKxzB8C
z6hMCP8NLq93Pqa6xeJSMRxldk1uD5TNzREsncD4A2eRP2UCckHPcYej7Kdhcnlk
LJ+DWgWuZo9iWuF08vkzAeFWCPfYIFZVZ4hZdlQfADPsZ9nanD0oZVRfhKbxj9V5
zzSim70GvAANa/ZD0uodib/Gf6jKg94FbEoTfRlBVaf2D7kvminqlyb/GQ/quGYY
yNENM6qf2ptta19KGpSkBTeifNNfDu2t3IZMeqxRPbScFLvIMBy1HfHbbY5NsbEt
epg13nTywJ1nUbPuLrXtt3bQxUEIC6cLI7z48/A/7wZ5p8F84Ff6lGYbm6LNRXx9
XS/xBHIhLCwvW1XReKmc5Rg4S3V7LAW2pflKOgS5+MZLiDJKU+dqglWMw7rh58Zs
txHid2d43Som+5zT3HyfhFaQI2b603vuU4+xFmqsh6FqqbHxF9F/EP1sOSSm6m8z
P1IqJbmYXAHy6Sv06e2nKNJW3Qmzyctoyke1jmB4FejWSNrnnaDBsL8ihPsscAVX
CowrV/ZHVU1pdqaD1wCQaL0pZ/I34Ohvra+ea4cgvvCPo6HFVUOCUxlCsYNDuVjd
IOrwE6CgGjCZtAk8G8qAy8ssVp7GE5gFpceHfT0EuAV++pj/dlO3Qplmb3TgGpo5
wWYkW3OH/Q0PdXmQw+wiGXBmonyYEQkYrc1XJpPWb67rYxaaraWwpYkF5Z8VMgQH
KJBJ5pqAeF4T6yVHM7lfhBZHQcM+SAUiz60wY/b2B462gZM9+AonCAdRElabV3xQ
6wzSO31V4nr+ajxPMoVgFYwYjfXVfZL8qgGWP0CtCW79HQQbOjrRNT/I/BoLsOOH
YrFEzWVC0fK/NkmcKGNk9A1bEnv80BQorQVXhB5SqCRDYUXK7eT244w8d98/bvOA
A0M4rABMqpbO6NRSXWQkRUNCUlqH5nt7EbQbrtf3hJFk9JUCORZ/iCwGueWG07/U
9S3z2uW5goiv5VZCEJhb7vITwSfz3vxbliJ/pPD7eHhXvZLGHiOmbBkbedCMb1g6
uR8jtjVGUA4a7IveYaHq8Wg1tdl5KG6PtnWy3tLz87ExpzS3aztmBie+LIoFC1Ao
8Z69qqVgmwRfhgiDLGBvkkGBXvx/QUk3T9yMlhMZbyAbycBC5we39BU1zV7rU7nY
7zw/8XE5PhsFKDB0Pgc8UXD77l7cmt6j0W0QExKp1rVmByXV2VYWSyvyeWJhF/p1
MyOx72NjAN2pgiCG0wVDlp0rqsqpW9WXwPYdC9p8NCLS9N7/E0CzOLzEEFeI7EYE
9t74cMBwfanEv88PKlQnHLs1BmCg4AO9Jkystngp/Pp5ArqqGv1AdYxsv6QEmYAe
w58s4bbjXDkTg788/nzRsNut/FwNa4S11/IeMUv30pZ0ixeT4Jy497K1hCINxqYm
mpPkoVWalmAGPUPhEhlqF6dXwHyIkQZVCwzpdKwoOda2icJITmJ3mafZJkFaGQFI
vlAHpnscM9fWJrnt8sFjjZUW96LlH11i49g9cmjO5F5Ya1mpZlGZOZsCB8mK+ZqD
R3f7UwcbWueFQ08zNtGcJc+YkbmRYVNlndtD2FVK9goun5pQkZ7hlugg2iqSV7Sb
Hq19gZZvn+NMNLews2k77wIMOPD2j+Xt0GaJD7OL9s9CCTBGV6ZeLfCP4cpfoYhP
RasBKnMYh++ao1yJGAYi/XfIzsVXLsZgCuDEb/HgTSbH3R0fC2GGtdWUKFwx4Rdp
R4wqkKTPzoXePtzNHNEaOPjC2P+am77e2khtOB2mWVi7zeD/N70cQyiJB8OLzV8z
Qjz6X6CtX7BNCtZPd6EW9+rmq3OkjtkRPIpnRnByfajmXEVn/WjPlvo6T6PxFj95
mjuOnMhC97zfrp0P+exfHHsnEkDBhm7TuGfApPhz1Liuyvjbg/VWMA1TmguSxStT
PBZhalDmCHvbAklqpVH4NX9QZFODc4uHt63Sgeg/ccCLg3otOtlW0FUjxoPi+iqL
Pv/5SUrFfzZSYAo9EPq8FquDS6rnnCwvvNptBHLZJ7mDQju9d5cgMF2bEMviCOKv
1ObZEb2SQGP3ljdFLT4Ai6SZUsvoi2KUc64YTCrW1UGFxqpYKYkxCCsHKD9HRyLl
zHd+F1IQk4kMaG5xQZjglCAeQhq2iqLHehNgehU8budxVjQCfn72AW73a524TjbI
GDRdAd14tjWINHJOzIDDCyeKAhlIxjFsxKDTYeIZPchIbG4XHtpwIDCIhVoKRvBe
iqVe1xRFb74DnzfOA8sCG6bLDxFf/1wgoyH5KAthOTky+bnwe0Ez2bz2tkoUSuaB
IM9yuSTOPHuErESiElbVFydHXSTNE1besmSXzKBqT5jP+FqzSQKVMvkmvnJI8es3
Lnb+CExThOXEtJIp06tiRogrshGrdD6TAbKKCPDe1/dmcCGF0riNAwKcPj3u0U6K
7lQkU377IrJCeK9bk8K/dWKea3LkHoe7laKjxr3feC7TNIWN3/IV1gFc6v9tHm2G
sH5skRoKNDJWapC8dtobqLZyhpsmnOH7NAPVpDhIP5yTiKHoSwyO1Gda6ktpNJi2
5PB6YwZLR8UjnFDTs4huraiV2jlln3A+7MUE9rLjPMTxE2sE5eh0yYKxvW6EmSvW
pKSPShwLu7cLSPVAj7HsC+wtx2Ng44ZeLUW8V0vKjTKi41GkwNgYCiO65sA9lHhH
7YzJMYuq+/ICi0gsaB41/rasOiKOxiD9rs+zg0xTQxNqewWckWgtVqKM6P9rgIJp
n3dfmfpxlkjb6ClYphWOyTnHk7bZwzZv8kuiQsXHUDwsrmW92KRTzX5B8LXZqxtD
fLv3dNulR/zsm8CqH2qe/4/NGywsE42zD5Hr8wgqTSNB0Mk7j6/LKBqtTAj5b+Rc
DL7aKyDYTSA1YTt9VFJasoVDMw7zjcnIHEF9GgIS9T+oVDhN8u+AVf3r1wWV+MjT
aawNGtsXeJh9he/zTPRoX0vjhX2TdDPIj+rVvrBI/MkABqHHA1YJRt0zR/U7IAOX
FbJDK2WyPYHPVjrcU3/Tnd6C8GBiMNda1PxV99wADW2x/iDp2mP4BVsL0q2fsIpy
/awAAjNShW4kqr9uYsoL/vEAZyTG+owIG/8dY43i6Ovoy1vt1ddU1Og7rueUubfv
1mD4vmr3jFYzsxoOeVO3cfVN1PvyPiT4QfEZRqk7cdLB9Of1JptLRcl2PzUoXnRG
T1oIjA9jIPmGSB6R9+vwDg6kzYkkkPAv7StxUDIAZ6XL+6tLCMT4cBhSukjMjy3v
//4KkkpG9BrkrBEA7BIEsvhbSwoFJznGPSn9JfTsNOXf7iSPtPkF805Es//5MpCZ
C3VvyHDUS2OFeg5CTR2uboGs3e6tC9M7VykRhVKz2PpfHVBelxBsCV+NfNwtiR4C
eRcL5D/CqePPKejHkaa+7tY1Od9WdDniIK1TmP5cnk9avnKTDhzxSP8yiIGZMuUE
ak55b0etmOaGpnOraGfgSBRwOh4k5Chuq+yfUcP/ThPNgJpfkG+47hxhjl/PLHzZ
1o2i3NPNJ7X2lCgTN0zVBjlrLuQ7+TaswkGkpbhrd+ynbajaoOunV2rSg15+/TYA
rTT2t5hrtVNsDq0cDbw86xe3mmhmQtM+H168zM6MGWwc/cfAn0010iSh7etLjgro
pn5JVdnmvQQEuGklTCzOg7Rh7znjD+Ez8N7wvDH8NcoQoP7UuIyJBS2thYJ0tUTL
rMOUxmRSny+pXRNuVP2TBy+1XfCJOrnpJjhHbnnyuNhjLW728aOiu3xlxykHsdS9
KReyXicixObK6b5BH46o/pD9C4keHqobplcFcSiVYYGDRovnaA6m4+grf/Z2+u9J
BLtdIblXaTNsPT8VAlSIr9bdwJ3SK5tDqPlX9kuYcvm8cr4eHqgKNZUggD/MmiL/
kWf2Gduhtqf451JXCVmPiB1HUbsK6WGVz+W39vt/RbQjm7s/5ox8H/kRbHoL84DU
D8931Yy+koYPHGohkV593EMQKI1FBGYhsWNBZ9NIr6/HLL+6cZA3BRAsryRRNaBS
+r8KoAvEmCtIV+I21HRkbeDFmWDuwXGc+nZDNiyAbm8KRj962o4FjWDqxRyunGS6
pd+wXUo5bGqWNfsNcqYeu/nOpWVtZgk7T53JDzTV3zwirw/m6aLdOdXAoYyKIlr2
RVQkxdOfPSsw10j1oFUhtGY7nMAy4F6Nou4GHyLvVVqGTT6LmiiE3hHjvlbk74v/
GzjbyMjRwQqcbreaszUPlDEBFIaCGaXhAtagLQNBSMTaaLRvy1xr5Ig+Kpw2SCC8
rwxUjpxGMyc+pbn6NL916GmpVkBXTdOXJAaeIAPZPebNX9HFtbAmGvlTUOxQQ6zH
diKL5JD+UtQtAPpFhflQJMz+8bXsJAGeV4yEoAezUwpVJ+WA0yasK1c4VqMcpnMH
swXMa0ZL6aTVXSdeyt1+CBGJ0dlx9pN+ETzYtq9PBY+8qeWOrvohY7AL00w50m1F
KEcDJBF0el8GQRf0mH/f06pusvFiCgEhTOHWeQrC/1eXe82u7AmWB09q3sIiAn/N
6Eo8bR8UXQPKSNzpKO31wjDWTYYzzEqD6gvAR7lL065JjhltS1YXe86TGGVlRqU6
OClne4m5EXLOi80mVd5f4HcgSVD4nqbFpFdRvwwTLAx5Cs2RuX39OUjh1gNuyH3V
sr5MIhVxVG1XMt36YpcRG3TnvXsMMgbh7QlSQiC/S9MF2YopFzAERqQ3AvLxykOr
hboMisya0k/exn/hWfW9jAIAmOJlgKift2Ip56OHbveiGiESaBSNv8deFUXWtFnD
iXWCc8WzkmaETZH+Ma7doPdbkkp4eJIlhRQAlpOdhMFy5xOXQ3pq4IZQfDWi/uA/
8J8j+G5s5iKYEP8msqye0sp88ZlWHVTHpNUJd7Co1/FRnRyBwt5cjB2iR5m6X8/M
IlYcRlE/cFWo/dFaK9/2vdruaRWLX6WAYvoGmy6Fyzc/S9GSCS1BALzTteGyh8GU
PUyTD4oAdb1VWbAEF5bGLP/w82Upj4C/lj7A9gnAovfGcitatN4snV06JPXK6adj
DUKmQWQojjdEz8aUxr6WQmzxtHQQ9BIqZmq/iJZI73t4V9TBXIIGNHw88aAvvtCE
vZOOEBHNUohM+Yu0bjC027ZzSQ7VztFlV/myvrZisowVn670x8BeZ8QN2R35BBG9
5wgFvnElumbqUXdwlT1wtFBLeeLF7GNoRegpS6vJnL87SkDgEiQyc3Bj7Td7ba+o
NGInnWcIz4W0oMvnLTVzTP1KbweDTfmfElthmjii+FJYL3RrHO67xZ/cX2aCC2pv
Qv357mucMkBynov6VCTw86HmQXwrCKJ1K0Bc5Q8LVeb28RkAJeG97EE5XJvX4FxR
vvvf5W8EvYoR+iB9Rm9itEPCPLf1SWHLXrvO0HmQ8BF0XJdB4iquUKMxX6DVvncl
SHGLDlQNA3UfJOYnbH90QKphKse6oK00LEWmAp+aDY8Pu+GgVNMJuRQHt6ODPRbg
45Ll//EKfLhcU1ruEss2grMoPmoL/+bXGY67GXfmJBG1u1XG3qmvVS8uEsz3eQD1
xuirv40uznbSaOVtmFS5SFoDxctyJW8vF9ynE0Oekjv1UEEgRNeI3PdfL5NPBFkZ
DrcCbawfe0D2FM3GiTyGXo2FCy/5noOG22x8n7L6lgOl4qw6CIHa9yGhmf4mE4R9
wSxya39eFtiqSk0BetpzI46sPKFvM4E3kaxaZSRFaXSv8I6c5h2yBaxhlPMvOPwd
+zgzko22J5AkBUSgu/b4UAcI6OW5lMFjQSXZvTbY4FyPl797Vv846NDFxYuT83Xr
/tnlWdQNWT1HtY001CYF0a+neC/tqjAAsrhyXgxLuIVahTZY3HhWtDc3b0GK1Nb1
dhYraC/tsQeRCZ6gTm+vIbpYcRXXJxylCQFD8a9UHL4C2JyC5FzRw0skRo6v5esf
QV5k7ubaRmNO9zzL7DyjIAYjQNCPISfsgKPNCG8T36KPwnaJxqez4hS6xvNqnJ5R
KaxfiwLYWsPox1Yc4D0VcSZAT0bj4qSrzqBUX63VCK/B+GmgqokWogNlfFnW8HTj
9tEDw5E7PFpGizmU8YlaXFKQ7n3Qr+fL7XNn9Lx7VYhqRQV9IKJUljSuxmZEXWfM
j4NzrLBDeZwt72xolcZY0fGGHyBbZnR26ygY5w44V7irh3qWG6mFNp8GRTrWkmPz
xyXPo10DrIz5s6FsFzcj89ju33xpZ1H6boHjUwfIfyFBqlTVqEoWbt8JFQTggMgg
iCOn2ckGCGtm2uixmoGHqD8nxzJZ1XY4XyQ+5ANPrpQ32dvUc8SJy1dVS546kL9k
0Vzinf6T00eR8bXy9RHWzcsw1OPFR1KuHYUlNA5WRCWUfe5gV/YkgUuFydN0UxrF
Ij6J61a84CWCvGhWqaoDyAqRI3aIpLcl/5/6BzhOMOaHA3nUaY4ynyQ23PX9uLOu
f0TD9Ud0P1neAK7UkrDhaBtw3Ya3yOEgTPkmJeurvP4YZjbAcE7TT4QGNlN1iS7o
rNH9yN7e8XHd3WcP6QZPpbuLxswb8IjbNhVJZA/aUilaTFlFcM9jZ9kUJJI1dTUs
zx6Ff3TAUQPC55IKDXeWCv18azu7fvZUx9oiQ8n08rUhPkQNHhfRHmrvZqfgz2I1
V0NfP0Blrbm1zgVVuqcqK/UddC4YwJbKKSvmbbm6r2LXUwYyIEUpItQRllxkBm1E
CNi6GyMr+8dfO+Os870fWUlqClhxWxPXkYc+Akq2+J1seElxOd3z+Rkqw4uimfzQ
1ex0HB7pWsqIVt8XRnFtMjco3YAka6WIgOoK54pFPRBAL8gKBstaeFla5cxpDmd5
j/SsmOwaN7DwVlIuYVGnSjfpPWZphxDQ+VXhZSjuBaD0ggTrfLunfvcxAwhmT2Y3
5TjItPmzj+8Atd1KEMxLqoRFE6dyIRaxM4/tIPYecq4DM4+MqZ5VbcuQzVTlEi/w
kBh3cTbAv6lCZwohQMfxDP5s1e+jZduOE8dt0C4Jlt2j5asyqw6XsP/FzIyOsDc3
hgX4hRyd9PDlT0AGjCj2Tlh6/3uN4uDhNBtW5JOSrcqTBHtiGaofTVlIW6Se7aAq
f1wodZKMa+CNgMhBkrjQfK5aJ94KEIHi2MohTM19ixuWISRKODXoGuizlvfe6RZh
7C2N+aNcGNW5dUzksvce2J1x4EHylosbFL+GICXCpPrIixQcHqLVIx0BRDKzkN9X
XkDwwqvhaRW1j5bDDCyDmYdyE+RUepSf4TQ5Qc3wxotTstPzYjku02dE2ty3VBhR
wLHoGoVf4d2t/2ctwTqlEAGLkZsZZE+rKUO4ALgvZIoklwRE3KoeXjkyooESTUTb
BZapAUG/mjSOI36bq5t5GZjQE3flnSUEM0Y4QYZP8ilSXa6VynxykMTy5j1B8VaU
ON8Jl0UtBsRI+mRGPEyGOUswoRaJzeq7eQV3fxMgRdjOz2qn9y6jdQfPrdppupi7
mgbmiKJ45VTGG9hqCImmafbY1wbbOn4UM4Z+TAbTTinAZogB1uFuNK0Ko8oqozku
2Z3tMOwjmqMqjzuHAIMNgJylXrNNfUpt+Nf3S+grjljW3/49SG1rz5JxCrBS92kC
JgysL9FWV+VMnz3mNkYn6fN5ZomR0EmAXsyDdhZxkpKnJQr2Pa5KW2uQ62XFDhID
jYyOFLAVRDDe2eOOkCz6A9ptajc2Jr3X1ViCsrBWvDwGJsdEf1roKLk+HxnqQuhw
Pdi7Z7oqQgCaI/6ojVOHIJnzHWfKrBHxEqcK12jUtJxxeXvy8wOkkCNr5ZWX8j2H
YoEOSoEqhsboXE6a7klodAPNlVCcPBsXsntF9hdr9KLzmUknQg79YXS3av2VgbhA
WW+x1Dvvf3kDdomGlh/o7LcDvSDwHDDhwBnNPLMcD+0c2ZHnEvbqcjWBxfJmCF9U
c8z4X74P88/tcKb6N3zTLp3YA/fIG0sH7m1lQy9DhVLuDXsWgepnAWk8G9+TZKfY
k9byPIK2tvRSINT4qcKDT16yvYk122S6hxNgvju8LSeGQQY2QzILxMR1aDJo9oW3
a7j7YhEV1uPmLpUAIrPRdcivELrf5Rn6k9W/eQz0UaK8TB2H30/t+kEzk5Pwtgmm
OcaFC4IeinyESwQTCzadjsrgotXsNdhooYbSs1MkVPxncfMOm+D359nnjHmoh+jl
2p+EaDbi4KZQy8SmDVDLrTL79JGxgcYEJ0OLe3Hqr391WfzZgjNy9o3bgZrQ6t0m
8jVhABYCL7QKmWgc/5N1x4JklHZ83RWnjV94tGgvpvHQJi0reKesxOkzFW+5d42f
QH5npKU2atKACOxYWSq2/yKrl4HKsPhmTh7bRWQip4SGBzBzeajNSAbxdrOhwXH9
W9Gtw5gbyfuhyCMNiCjCwxF0ACLd26RsEG6pVtEPhRQdwulKKoM7rwUfCenubsi9
JBwe3n3TwIsDgeRyS9YHhiMu8uvti7XqN74Yct0f980ohoJ5wgKj4tkfDdFbVgLA
VtjKbtJsbndcrcbD81HokLbdnNGmiUvbc6F6eM0TGP5yb+8BRmVqnO5Xl8ZfkpBE
aZpTrWh8wGZE93K+CVcIhDyOBI0Ka2RItPpA8M4/GDkwOzXBYkNJsWMvnDsGE9AA
K/XPeJmsPE4k6MIZGf5+Gzyccrk+l+It8jMeuWKRInpQgSf3U+zGPJKQHWEDdWTw
1bGittus2AUtlLumk+Bhfu08WPUmwSSYfWwRm+g/RyqIm1BR6XjZFxcSsiOiodkk
yfMeSmKPYjYdlKyDM87mAP4fS6TZ/M3STQop4W9jXKlAqBgoElrbAMJE0lM8ZndJ
ZukP38por5llnuWXubJ+8hV/WLR84evrE5Z2GeDBTNU7RHLBTAUjDISMmyH6y4Ju
VH/rDvkMjc/umA46gEh+plIFGophsiNmGSKNvrIBZvPjW9lSlGz6AcTRsYb1lKX8
z8DTTvu9am5xYAn6GbfDUE2FCySRVThQ1X6qwLJ7GShvamsRHfA5YAiRU62N6pXz
XczKPmAvcNY/gGHhZG3NFKAJvJm97EkYue8x+o+VBxqTl7R1NZPhHT2E53+Mn5qE
EMEpC7xww5eDetWmEDpeXkMEfZ7ipQZQV//0DIBFCh9H+F9amRgi2sX4/TuwBleu
UDL5qsdoxKqvr8A1HYie0A+0sBOXF5pXcrZ1TBkFuykKF47nwYNxigRpAIpjtPHb
LBWBltfwfZNKP4PqeHQ6gQl6bg/B6rudPdC75JjGPE+JcgSd82BbxGX0w036+awz
PP01Wq0DAdPzBzzpeGvu9r/jKnckCFvsx0PXwRknRGItyOHeDZHoRW9vsnEFogrw
l+YRbZ/oMkDy+R8hR1agK1j746+1K5csXWN1RvFl7QzFK6lK1bkKNmaiAE43wUgT
IMHn+RX7zzd9d1FdB9SUl6iGtXiJX+XlEsysIE/fFlyruKZrfi8d6lenGh/YvfvN
2D1Xgj0hiSBx1Kd0HvG4Ivis+OcrzIAqZCL1WRZxKHgD1QsoSZvCkkXJJ9Nm4AZL
fbBbGGpx77WCx/+KgIrib3CUgt3nod65v6Qsvkj5AaaVh9XQ9auwMp01bb5vZK8H
i3Or/Kd5x3zLpjgTTJpELIaoXeLKe7Q8X029zV+xa2VeAywVtgYdzV7nHNmUQbFy
3Xs/gg3ofFCBRD/o+RWqbsl4gVG4+MiAY5TWGZmTlVd7nQuoJdK30GdCEqIvnB7I
WzelLdyCDRLLXPkavrYE9H5J/o+ZRiDt0z5fWb1cqGPQX3PhMXSIeipxiB2g2Sf8
3TNtM5H5lL4pjmVF7KVejpVg84vM/3CgJmsqDDzxjXpaz4qlhLjMpElzVWcbsAGN
C59ToFLMBVre7SFXY/JiZKJaYN1nC7HCMZujZ50U3z4k7VlwOKM170uhKnVGP3W8
a6oTtMFZ4LdYr/kpcQXoXDsPOe+pryqhXxbkkuh2Isa3VhHAC5nQvN6aXJK2ooC9
RgAsiwMquRrqZ9hW0H+5B/ghhIsTN8xkkOXg9wUXfKxaqFw5fJGAkX+LfMo1uPCX
5znxylcFQBu5Wd6xTwBO2oQCPSi/xR+pp59Q5nxdBLUbVfDc/6KpExFqdAlwOwL7
pM4b8pFpZaP5/Z7HvWVo7STbGo5YMCGi13Hz2WMMEVsqv400UZsX2Bm9mM1RW6L3
jo/8EHvtKFoxjtBd0EJ0BK7KB5DqyH2bGTQmjaGRkDe2+UehCMcGwQEsMItmYwsj
L9Ced7+3/Z56rpDVhexuzxuf/QSAPkLlT4P8z1x9hDwK537G8qy872ngOkZId9uq
LYHvYECfmLNY57BXrxhbP1Myi4jJD6eAGn1xhQdZb9cByMRgw10G8zs2vWCp4jyv
7GGTc9Bd3+IQiFZHXef3jIF/1+T9Xu2ovvt633jgtp9EsuOY1G1oIQCHCm9UOuiT
ZIor9wBKcP/sV6wXTEmEBV3Zwh3Y60aQlXzySQYEjaIz7CKIHaISd69KLtIabwe6
sL67gD1SrjJXtEXebso5yWwCmf8LKJBZ4s4Iqdyj88vqSCGg1NXyOHknA7mN3xNm
gLSUffY2dEAU75cpLQENaeRjThNZcqCLcFnxUQHV7Kfn77WsYRh1PqMpP2lndIl3
DvPelAl6LqguWPsMJTjp0yPnyt5lLQq7stzCLHYsimKOIdHl09fGvTzQz0ILZ0E7
vTxzuHO5xL93ihlK6kFY9dLYWuWB6bNxgBKFHoIHJYs7MyR3XKs7d7YgtzZ/P+SN
L9J/R/VdBRNn3XdlMGrotnDKBge+AI9MKUJmNANJTmnwYS6ooNm8gk5RvNFygI/T
eupkb4Vh+mGfbjlE/yC2QgKE1RLddDhB5yutkLMcNohalmI50zmkOv+aLIwYM/6/
R+WjdRUYroiWnoxtibt0ycF7jXaKtLG/7EiGypncNLAUlu7SFxNNQzNdSLbHrHhv
X2BPZIcEpgU3AzAVs3DAjPgZ4liu2sZ2V9tfZG6SU7K0dT9hXjevjkVA63xK709g
E6Npgi09JXg/ykWB9rq7ghzwhZWhS0S3oZCdrLMGw2bTU08BnfnVQeu3T2L/JW1E
IntS87yv4VrrtpIEp2mN2chl0sj/gRdnBc5h7Y2uCl04wpIZRbGUDz9I4EQ8e9S1
X4DQ3WTJUWPGfsP8uHuSuMddZD8M7Q9sziPq6h8FlvsoshrD0ZQo44NV+MWWMZBH
NmWfaNFEwAVEj8Ub99FU21OgF+p/iNTTSyk7RjDSxu4CFMAiUWwwErP6XzBPnI/W
jRyY0JJFiFN0owlTNopNlI+XbC67L0F9BtGcTgi5tl6dDuoSgm2WynW7Fxd9Vr80
Tw1ts0U9L4D4h/23BxPgn0BNxoUkzKutXfA2SlK9ToXsdQ3KApI0ITp/jZvT5S2x
Z3n2QE4vGlaUD72G3oIU2tgpltsz0UA0bQU8b+qqKKhn4auVfnj3FEpjVTn5ZDF3
kqOLwGl2I5gKXCcqjuDBAdb1Se2TUzqF5iiqvKW9SbR2+toJyg2lXgMkEcUToZbj
x3El/QyoqDxN1CkVsrFZ024H/+aRGIzobtu5ZqT6f3bsFjdlM7uBNW33vTEwofVn
U3FoV3YojCgvak6M75WLzkPu9EyVzoxNxNlth1No/OCXvb2eCul2YJQrXeCbognA
Cx5c3whUVFGwYRkBH9wkCpefFWSoyCb0p3vhHqIeaOSxO3RkrcybAT4lYfqrBCi6
QXKdnMAJheLqggzTB/GNSWrvGEO2IvXs9KOP051WOBt5/CHtqH0WBvB8/dIm9mAN
ffR1Z5xbuZMWC5WBfybfzeZcqeXwSzutWwK1wmGIJyfNvWKbtZQKWV8vyZR10dqC
zSpQYLLyxewZyv5mrHipJpJL/lbGjBa68DkxIbKRYWsClQF38yrPsDum5P8uR3Xb
SsXtvmKeDtTxJ/c5PhDO/c0cUSNAz3IsSmfV2kY/PuCtlbV/fwXyDISgWYraoI5v
2LZOHKmGH/jm3BG9iBTwnoz8jvRAtoPb7nAvgIruh/+Xc+ktcD/Isy7uZBFgt4gH
MbaEB3ipzhrVWj+kzvbrmXptLUscgoQieAlKA0y4zG/Wu+8TWwAXkT2WgapCmny2
yQ6qhdwnGSgC8ijCnEFCSAE9xSaWb8wTyoThblksWnY3YJLYjDIHaykBFAvgF6zN
aBIr/HjBZHMcj3nvaH65GYeCC4VVnLZZP3aJp+0u3m6cdDYjLaH/HWbYue1ei+8w
DzpbOTpqKdNQPWaxNAtOJ3LKs56lQpxKdBDg7H8vMIwpum7sxxGHbTTkIf6GrYeb
4NqwbEL4IX/BM1lpU8Leg86N6b+aKtlLSgRIjsWy0Dpx8CUqN4TsI10UEQu4CrHu
uZulUdIvIcT54v7zb/KrBUMKBKeydNmGswICq8jx6T8KQmFH4FGBYjnALVGtKaT4
INaUt39BJ6YAMhA6LQz3W6OtN8OwUgW2aNovPxYQuDP50GTZSwFAFYkERDQveoVW
o5ZEUU6xM5BRD92v9LsO0CbyMURiVYkG0rTxQxO5pNe8AkoB8gsB7nq58kO5OEPh
mAHkqmyqkbcau2Xt2guyZK5q4s2u9bFpZ/4rcrSR3IpIzCzp2OxM118tguzsT/Gh
0WnoUjXAyMA1XnJI0eO8wYA98+cMxVak23ZJzmihEW+jGqsxyi10wREkwEfDFezX
yVbV03QPDQaLV2cK5QcTJQCZKycANSJfImSutSMwP9cJr6GvwvLnRGDp7jorO116
RFK3HLNvQ7mSX9nKApFqHX1kC9sp6+LS1wL+ohZ9UT+XXoVDRwR8PgvqXT4hfxWr
BcvZle7aa8m5O/5ssIpc2WIWvAy1b/1i8cZJTH0ihUG743FkuNU2cLHxwILWU8/7
PL8DGHwnVyT6sUENiGximyQTEm6vxLm5vkbjzjJWWB0cFoM74hd2rOoRXEYwSOgf
BjlAtmOHUricq41Cw2RbSBPjgKNCrWEM8tRqHp2zaIgQ63/HYBfrs142MQi1P9Dw
HyisM1r8mJJ61XsRFx3gfD1/mfm+Y39RDhCMmJvUGyoeGMpvqv+uAm0SsMljuHpC
QyqUKopYVlU/3ui31djMII9qbHdK0FLd1N4u5cXw8t4igEaUM6mA4nQJcWBTjARy
LgXQtvddvS0J68Qpho4TuFA5etW++KkrRO8+JYEj8B1YdwJVbHUDAmV8KWn2fJrw
p+D5QL1sre278GB8E8S3o1zWa8SJEeIClH7CGCNoBCcyRx55cvRucrCaPWFzFfG+
bJOzyyRyYnvu7lm3e+isZrG77MkWX0NjurdrdS5oFLrZMQsV8QUdq6JVorv2H0SW
a26yGUkeAlz/iqXGAnmQ5l3fjjTccxezY5DqheNppwnqpqLdQJAq8d1SCH8OLfdO
0fgfQBH80q64chJQ0IK752Ozo+4cNtOz6de0bD3ucphsQrABEToUKVrQbeizOGwK
KeNBEXAQQD9Lo9/S8IeSsCDGU+YiBMKBMl3X/7geyOI7SQvUPyD2+sASQQ1rLmS5
uwuPblKb400rQcv0G72Jab/fKg/KivzeNWn0fnd9SzEsPsUTEM7xYqAAvf5G2r7g
DP6koHxbFnC067ey42ze2RqiAXH4i3sjl5eBp3XPUJskJUq9IlrCTiQBmeSOJOxU
EQbQHD1V19n2d4FLVh1O21Mp9rtBXPgH+srwFDL+vAtYtMM6DkGQQ3GpnGjBzpie
OxX7wEQo3PvTUsutWECnQItuC+rFKeers+NBiStrdilFij8JfiBIdcRRGsZCM85a
c5T6BrwF0WKEOnRPSvCFI1R3GLvBo0mwHSgqk6+F0Q6EJ/Czn32471ZMXx2B3FNF
FYDzgol2taaIGQVb+ckb2sm3zMbzb/alEh4tl2oLuH1+9HhRmvwbjGsI5iU9oVcS
GUiv9k7C8CGMzGaQ+PRnrKX1Ab+9mMhN3wBsyuF9Ah6Ml/ucaV+ipXWDqVc7d/NU
H0ZMCD7vMRRse9YvhlDH4FPvdbfhKId5aSdu5+LaGDnILC6KsZh4zUmtr+U8fHCr
tagibuasqFDOib3bcdI2lWVqyDFtEkhRs4RDkJMPrwN64tBHQ/B8tbihY6nRxB32
h29W9TC+fWnJoZuysNg9J+I/j2ZYK2TlzqZj96POE5iMuIQF2xszyz4OLF60w/XM
RbGIiBFGNq989Z8gy08l+TspaAg2+Ex8v/nsMrGx3qqjS9EUDzNUpW89JSfhLftC
bu4w/v6eoCdgTdnGfhoH7FjfkZwdcle1DYbEA/qBOl+FVZNAVTeBRmLOwp8hrUHr
4ek9KP3ZD0uMCaAwn7+UugC0AElIocxGea594APyW2gmOVlrAJUcZ6Qohd+EjC9Q
nVEefjUQES3HAslZBIo586rB02OViqFCi431aIcNqWhXyd8H6LvFqXvr971YrNn/
tLGxb2eIoAtwodwRppT24L8EC8MZlOfvNvH5fzdbHdKA2xnEuTk2d1n3HoF47Wr/
0/lx8dD2o09ueZ1h+bRFTCuVTW30BRwvWbdCjVQWG1VgQaTGOSf4RvBAr6Zb2XJp
qEHHi5WyLUv7RpjzhaUddYr9bH2sQBviGQswM6p3VlLRhdZceR4U0DzxnDAQB6gF
h7somtRMjzF12aImRW1hu22O3fNO43f3ZnJkb8JNXM6buTjbrAN4Rz8st6EO5r9M
SeOeQVFPB1ehXpGaa9a1SJaR5ojvGv4pRfgFkiB5ppB5DXZ/3m7oyoegffVrpYCb
8oBAQOGqpZDxEjBlbu1LA094dGe/WqxM7msHlCOr/NQYawIdiDkILxNRIIRlt9Lq
E3tixCVvWyDxIhz4QZRzTahgwcmkAbmFkyHBC3aBQAGGqGeFAkN+Gzv56eHz8Eeb
t6hfwivhNOy6TNEemt3YSts40u0gFsRiw+ZCOynuXQGc0CPKGcR0fN3s/bvlDAyC
xrErGOdBjkP0YVuBoPDaDWX/UdUBISMWwn29mYSxTFuSCrvZ6ojmgLerfeDQ03Ja
P669We836W21zhFgn/iksS6olSp9gcWkTm1kGwkQ3H87LgsuH2viLSqWMMijeq4e
CtRmgkt7i9jApxT0tnmxdjdhcMSOpRloCyjC4KPe7YNwt0AuROm4NKOucPqRK7lm
Dc6sPHVLWjTm5GKUEjW5//BFUWP3KdQgthhll0P/DS7iOFuZ1mPMRzBjLndDUnAt
WVYdIR32so8CiC8CKZ9A/JSQfmHYMBq7GPR6D3vpYFz2OCuTUJoJjzkTs9Nfu0vV
CeQ+BztGrimTe5BtvY/rdtiWtiR4x8UAKmeUND3uNWpxsS0eyUgLgr/YCc+NDCME
lvE3KL0N7hsh+bqgukBlOA4jMBRowUDqpOHEu+xnbhgwLCNbZ/nAqPjnZJvtXQ/d
RBVyVUk2Upyii+05tAU+Ka8QrejgS+UY2nlc1DwRbKR4wtwiYFgZnHnTvv+y5+Ee
h2T9WrjdKBH227D29rx64E9yZTff/2ZGIEorJTxFdd3DtSJua7dlfFQclZOW4Ij0
qF8IsxYj89XrwpHsI3RKlBTYo2AVtx/EuwZ7AXmn58UMWiOT8T8j6mJ3lQV6zM4/
hrqLePp2XlOoTjLk4nw29GuPUNUjja4UWrLJd8hxSJa4zajaq7Qq4Y8Zl4XhkhG3
Ge54gyLukpXgq/6CcIutuwuPvsw/M3/0ku9cq40sW31gUWVCcWvFa9pVf4aKrPTy
MZKZWpBj00VBSRLA9ALtfxA+XJPXjzetygEls7q91SuOqxXExQ6xg1HoHYaOR+6K
o/Lbwk1hitlmRDAoka31rj4dAMEmVL8QFHJyAgeuKFXya83DwbYiDrcfKmlFSJ0Q
EZrN/CyHbeEGM2V7SYgkQKYiDgOSG3VnZLLqTZMfR9SwV0owPGCP+IWw7XX2JOBK
w9qyxT8DvethbtNikjwVH5tuP+LYuNBk1Yxzkhylxdp9i1ph2R4X/lz4yy18FzWo
awm9rZPBD0t1gAHGWz/8P5E+gluMxYoVeXUulKGKAQoHA+/ENdsN8XpGnwoY/xvx
Q57iin3doJI7tzRjXr7oSIqAwq+CSWHoPNsa6Vpj7pbonvjuLivqElkJ/fBzAaf3
R2SFgIZ8nB7hmSnSI3xB3sUnSW2AS2KM7nQ/ROQBAjX/Kl4T08Nope8FVYNmfaUe
4XuPq1KYGnQa23pawRUYlSvhcQwKe1rkIYo4r+nWIgwXeD1zItw1E/hxhZ2t+Iop
9qb61qDBbMp/WP4IrABEYUcnUqiZ25DyFX9l5/w5mu3vTC5F7xPv1z+XU/tvqmnh
/74zuIBfMKWTkeZywOmxkPi2jGNY2j+lKrjTlh1/PSQSaBVbyOTg4LTTnLwrPPUr
N1/itcjw2rs3Rxr5SHBmepiWDOD07yL/7AbdUS/7ms5uGgGsJD/qipUBLsC56GG7
BuMRGRX+lrY+3SmpIivfBBsTaHz5Eo11QjK0D4yyG1qYhJyqG57n2Z88hlLOVeQK
kCzgW715IgtBONddVabhtpDVJ/1aSnoV5wvPhYyWqd2dxf6go6CiOryePzw4zXqc
axox2xNNH1s9CoCwtVuRwRVe1zfdKo5h1UtAUHLMAXz9Uywh4LMbz4AgyBe0O535
LbA7tZU7iyk/H/LKSjxXr7iNNcDniL+riBDJByV7zo8ImCh9yoM/r6hGHseRaudx
rnek2F3JO3F0RRgCH/rnAy+uZ+2beCKBSpyYxXTOPc0esj9QguNj3Qw/BWaOjGKQ
ZIXp5wWdflNE/cHwv6bbx+bkLfzZvVBIzA5nGGqoNVQoQ/vcGI/JzpKsaTMIGrf7
h0WA3jrPVRTyClG+BAcfb8LxKssbzsIx6nD8ZlsVgmHu6ezAaBJbT2IVciweUJT/
a5jYOjk4WEHNzT6awy77WTnr2xb46C27cfXX0N4an0aontSWhLeNWl4G1Rv0WYgG
+bs3Qw15tjBiNl6EWnNFyImdrgqVPDs+473LsrnZSr47HgikugwVVmERU8jMNjU+
MruU6N4ys28VZlnJTAT+mG+t9TIkcXPGYZExoOr/Z7mj+KnuGJnHAtPWRlMj3jXp
RL0BVZ8y4vCo0+YxthgVNd1+ZKbskIuFVZ3ZhwaWqFfHRGD01D6DVr55tug7Oss2
NypKnp78G9bmT/4ipzyiS3p/WsAnD34dX8ZWhbaU538NpyKLWjReTHi5GM7w3/Wr
+JepfS5xF+hGYDIMsq4Ep8CL/v5lhl06yyBirvoh14Ro8Bf8QnEiJkeQQP0HLHSD
Wz/HYM8cGJWfgeE1miaVEYyKd2HgQdX2NuIuZvrWt7B1Cr4mD/SoKhywOk6vNxLc
O7Ea0GyYwQC+xr2FFbsffYOnfOsMxXj5h206BlwiX9bNpRnn9t08+WACU+BH2pkJ
RmLYqiF9QbodqLN+s69RkMloiHAKNfKPKJd4sxgmpBp2py2EJJa6+Jx4pM/HE3R1
lZD9iB7GVxGgFiUOjXe9CUlF5/dgeux5e3IJmZaVGBQKW2r3rmFSsDLNUVO1hTTn
+FXkbJ5DT+3gz0ZlfQqWy/5Rc3FJA80d9prFC3XwMFiTGyVYuq+JFinZi1o3FQ08
l2PFJwatMrmf4KjeduPTh29ty0RWkoUxp7yS49qwPIlCYhbmWBJbOYYS/m7aPkg0
u238tTZfaDg58ZHcHER4kseH1n1OYVO4naHGP7b3Bcxe9jZDKrsMvNDaQiRAVick
Zw6aj4MbsXStHYm5i/0znBLj/DCkvb8p3jll8ynW3N7v7ppy5QhcSL+6t/F/Va7q
/hxhy+RztyJIYEsCs6rP3CXdulNjrBk7c3E3uLFS9It6tx8hAf3zqkHe3lTcYFdi
pKRiwQYn8hUGKyvOxIEYXTTcTRG+m+zM9pAhDi5ekEmoO8BHe8Ft1FJjukGV06xv
Mqg4jLh+cLlkxC7MSAdeoR+jLr5/ju66iLWXkXVlwUpfQsda9V0IdSM4Q5EM27Yw
ZaKVMDHLN2OP/CcoaLYy+jGlcGds9+55mNvZL5nfHbcgb0fthafu+3yjgmvccYlf
a4u3gOXG4sgyzhCrxizhvnRuyoVEO1QQbP4W9wf8lV9jzCuRupZd8j+fZj372onL
yxUe7BhxuLxORD/zGSld0S5UD6KJFTKBE1PIivDvvZT6QHabzs8xpRhkvAGpO1kx
KTNY0wBMT2vqT6Bj+U9LgF5rR5ro2PsC36bryvTG3eDFlV5W0MElQO97BYsAAo8y
uKmIzvrtLp4vUbktrURCOhpTDokmNPE5R+ArftFWrkALW0BFxbIts9BpjXO2rRwL
eJcUIalfyEkvfAfNXs2K5RCwHhgd1Y0vgtXTRLojNElvLuRo94kLsBbI3Xa9XFUe
H+fioglCfEWbJHcwBpY9jcxWC+8pGvimn1NiyNRFIcJ49sTj08QudWkBQjZJ6MVA
kBjKvytL9kLW7LGyITIDz41jzsM1oem0b44pqsyuwYRgN0+g6JVb49LOfEcCkII0
4UOdvE+p5pfZRmmCH7Epr00+X34/8M5KPQ1B9FxPuGxtsswK/SCtK++HhFtRTaui
DLQvY81Gw3Wh6wv60di/xw5t8G/8Aas4OfOMcQon/kJHYZHWjTU/qb7Dh5ZuJeEC
rB8Pu3xaVNy3UMVaYuzK/vtnQR/SAZeflnylI/MW0fzl/cVgJvwrenEtWRGbrqbO
nTHZGtoLwAnm+k/QrK+tY8Cpoyb3W1dV8K4TRy7/6ZljWRQjntq04IJLWc+Hgb4Y
fDjVVPBLrSSnRUPJ+yZUIH9yh//3dBwFsI6sR5Frahxf51ISu8pP5nW20+8Qfylq
PzD7zLkWWinh1VNVHfuNEGyGrcKhuZCZzT5pG0PvY3c5X/8129RhY2+fufGHJKsZ
N5JA+C6jkcQB/Bx1LFW/SYFI67TS9/MVAnax6OsAlECmei6oFAcHOO6sFnnBuc3T
9NEp7rxw8E68RNcP2Kw3MtIxkAlF8LWuDLa0Tm56hTE/Rp/Pl3LRmANk4A7oYg4h
zs+2qeryEyZLeBOe7PokzRXNdpccB8Kn7XZIh1UCLCZobQLcd0zxPMpOAek6TSlz
+/S9CKC6L6plxJ9ZAjZpPJ3uD5/U2NLtvyUms+SWedjlBP1G+r0BYZS4rm2W0Khg
hy06qRqIXuWFmrIO/7ic0OJST6u02CTh+xTB86TpsZHnTi+1D+cz9E9L53+Sf6XA
b5mFGyYuMQGAqbiSWnNpy+mZIPYKMLwASAXG916AR5OfbfQ5uLa1xv56650zMXtX
3b2TfLTBJ5gvUWPOYH6CF+zdfjWFaUoeEMY2pYev6Sp46XVnF/1DiFkADR+P8MZO
ByYfXcyKr4xuYraUKshrsOVKCrI7dVWDZPrcvZY5nqC4n3vV4Jt8TPiuBaLLLFqB
jUzDjJ9ztAELN3kfbkuAacanj3/Kr+I6wf4EWoddibBuduSJuHcdQOy8OLHMtAGK
9rCNkgTKXKYpr0uPQYT822Jwd/3/4TnoAmfMZAecddtaC7TslPWS56DZ2fbxicWf
sioS2kyeloH3/CvGN5dNhX+bMX98kg36/FNFoci2LzjQ1zrsqj2lTnApScYWqeZH
EOsPgRes62DaKChq0kKPJ+/J4/MsHwNsMxZx1pdv54H+j82IcSHNz6dPTJ3vnDOc
1nFk1NBz+ZNiJzMDJ0Fdk+vsXUhRh5Ztwcb/ecldcbYtcbjapPK9I8goXJXrBZRo
fYWRTpbnNwryfIQwy5FGyNuOUpDrxZBCLLwemrmKBeMgU1eH1UtFRri+03yraE1W
XocgHkYK5HC3F6rkyuWSERvtcOlv0htm77TgykCXrmvwDZO2scYF43xrUEbbp2iu
t6Q327sL+deaayWf/c7cM4ezrXeCeT4TdnEAYmyVoTFGTIbGFGDArJrdvCjEvbsx
iiJGKIKtuO+JpIlRIFzcJJYyw+CH0UcgVb/A9LZoVx98WN4xBn4LOT09+yk5N26o
42uCBnVT/uhVz3ExHRl2M7LiWKHuLL4G/vbaUVuXL7M+nsrJDSzjdqthYUF/N3Wa
kqbsj6iXyrS4+9F8ujGVABMM1g/kDH9HS4ZSyrvvBhfsDu1oCso1dc9gIBSTDOTy
uqiItGmj3MoTKnUcckMD3gtJ6MiAYEpPUXFB7MHM25ZgmF6l3HzdnJFwZwt1IftX
XJ0yt40keZNGrMT2rgb9J0+N1+qtLtlfORT9jrei/gvJ3v0tV6466AjVQk5GJ/Gu
Xq+QU8F06hHo1VzjQ8dY3jFvwyljv8q89Pll95/J29YNjtoxx23zaQBmeIBwn/nn
XFF/iwK8c2dZVV2CbeO9GuCLvKtSBfgutUE3pNIEqSLixEsB8TE6L8eOuZd3E6+0
5nFNF8Eg3kVSoLEqzJ2lCwHd4DBiShq/v6+9hmVFTUeX61kjopbnTvDy5/iKNSwm
ObrdrxKP+c5U+3ybTvhAHK/2bTFlv9er3IEVuj6WTwhcxoBGOn/V/vcVd0mntTQV
qyiC8xzd+fxUC2MhcA/9KNQHdxrnzoAEeDgbe4Hy+ee3ZDCiSY5RSm9jJNZKPhFh
m6z7zfdxgYeLoks8cmfUpt882kYy+09Ttb9emeWHGjYDlDqie/vk/uA1bwpb6xmK
keQ9QtGrWZtaA/oAxgfNGNTnfuiIUYgBG82kB0X5G/rRp8/KvMDFsiar80I7j+8k
Q7mluHFy33AFzDnv5V/7SfCPYApud8QT3EotfKqxJiCi5qSCZlH6BYR/HIOB1Gqk
M08UB9igDlMbg2l3bsaVvOBvlChSP+gyTs5MA9B3oAFowx8vEGxSxKLTSYvvFQy3
iv7+1HlhKJZDo/VYmpnH9YIrqSxzK2uDZWL2KfwCX1RoE3DC4+4hE+4m6BKETND2
bE/jLGP2a2XXPKiUH6EfAKgBiwkT0OecBbpGqFqZUBSrfr1bP36pOKB1N/5SWBUa
Ic7b/spX8evZKUdn011PwGXlK6zlqcMIEQw6cdT277VEezkAKOb7KFLODPbQhLdr
u4sZem1Qm9ir/n2BSL0laCB4iFU3rzZZvk8PxeIsTK+IDExhSly4SZGxFDCUteB+
3jvf74QeD3TC9yM07JUDXfC/njgX9nfOefdqjOdUii4M+NiV9C4WPysiu3o7nphX
wQ7irNTofdZnmWCx5pdthc9Sp2YonjB9aC/l/LvQHPAYrHxe9W7QFrTRf0RhkgFl
1qm3eF9xYyNpWTp+swKUxGV5r8cfNAEvK4+290vRg72kfjsw2PWPvlpiy72KXnzF
G28v+BgcwR+2rv2r6/JfNj5gHzyWKsUh/L7+cH2tzSdt8ILfL4no78WykfbLDA5M
ZsIaxtc8FleJ5LrSz40HBrgFVXlHjcCcao4TKUVlVP7iSmIviw7Bf+TmyY6H+Gj7
f25gRFsWP8/hbOrE+OkQgWUDOma1aD9gEXv5ALrTFkCL7/U3gHNTZBqXdNqLpr/w
9abjvJZbiReNoSF0KSfaty8TrzVdeITV0m6UOTH+jZJ9e0o9mIN7y2vheHy8s3Wg
az1qKeaRVdUn0gzdLa6kswmt1L5OqMrbTrpZA0qiL/v2bT4T9vp4GlsaClQ1ee1w
Q5SLWm2oVKAnN7QZwOcLYOrtfi61IgMBVf7pxmYRfgeoeXminswzoUyfdJvqVCqL
vo3MTL358meDFcb6wvnv2hvDelZf+iyt/gU5SPx6SnLc15IXRs2rb9GgqzmkCHJ/
gYbVXzXczFMR+J/NCo5UlXl/8sxIn5UbktTFc/52s0g0Pme0jjwdjUge7AZ9P4m6
HF9ndjPmvTI2WsoobD1yBmrkYZ5qYiutrxijBNtXzKxo+VM/HL6XZhokqq/4/XKG
UFro2lt2DtFnqMV/AeLHAitLjvZQOQSbnhj5MiOQhfDf8435rDcOyoHBylJBBsR3
m1dK24n2Bc9A6wxtyN5slQSlY390DlJuBTBLm+z6DCB/1QzUgEJ4E11GafeDEIPV
2pkJoozIK/x2OHtu1WAVQeT2Q2fpKRKgbyn7yEz6Hyi6dcfM27+mx4dW3Ueu8GzG
UP95smv2I0zJEVk2gvgPWif18vV0t8Tb2VKg7aZbOFwJoDo5wgDrlktgFCl9gMIQ
2PWeH8mny7r2vsQWrfThwT9HDsY3i3zM48Nfq7nIRR1O592BAcs5jdj5jpgIHMun
8T409wYV6vbQyuLLVmnJoI4C/aPjMGclGpmaB7Av83nnGOHLpxCiEB1xS7BAKCOM
Mvw5P/ZKrcvpOdnaBrNBcHdLQp9suMhmkjIsSdfS3Ej39ZCjHjpvELgNQdIHfxWv
zYK0oDxwWW+HBbjEKTCL/ZbrNwHE2JLOpHv0KATxS9WyKNHKgQBPztqC0YtB5Q7O
kLSjEEF4wrN9cXqHKM55WOa+ylu/iyER+BdEYma+hzNricyfeqAsn3TvaYAG99lr
wPQ9Rl5bY4/2XJP4SMoWdkliN7oxzFpifQ5p0A9ALoGD83rituLv6g/gBsx0H40s
DgpMDlGJrBAWiA/xQ5z7NJYx9v98rnT0+KNcqLCBjQkoYGqFEv8aqqI0+IIDPOA9
caxJ1weOd9pRxTf09lC2WL/36E7ez6uVQcrRmhWgD8+aT7MBfP25CQl7QbSvJNCw
3uu9UnLQM/AC5LVyZNE1Hfy9QGbfpCMVLU61t7eImblz7BeZhphE+leZWwUQhZ9n
OMOitJCQc/rGFOD5vQ0EtCo+9tuSRyIWAv/u2fYcgr7PdvQIw55J7TdEIGF6Pytr
4LcD0wok+nS678bpJE5phXwY8kiPY01JCRexieEYSX8GsUUpsMIaD35dyRO76SVl
MVm2DmyDLfBICLoaSVfB6dcDtI51goVCuU/vStin4qVn0jueU7KYRv+sQ/QfnZmT
BeKo4tQj4Hmd4ficHV4d7s8bktdVDqh/LgZ35+BbKJJfs4B7gYAV08/PEzwzCCqO
/adNG4+63z6YVsaO/BPSrU/Hb/ffJOseYrlxEqSutJWDPjz34UM3zQaFE2NY0qY1
ZQ5vz7PRKqN+xjZOolpGmasiQfcjKdAiwjd6iDgFE8PQR9olUGEBVsLz/Kn5WrBg
3fU+InMFKsJBf3SN5j/gC/bLdvohRYDNVP2W0y3tUZ7ai0AFklfmGXuneI5LCQFg
Bm3EDYCfiuaOY+5tZRPvGpISH6KcesSp6zoDh6ieFV9pestXm8Wy43Wy9w0iK/X4
AdOAhFrBSI5ZaxuFM7FtZ7QiZzoGlvyUJQcsoC7jK2JjPo2WyxFGPZjiyCJ+O+pz
31T0g7juJM314HTLBKS1JJ6WwobOSROmJcPMdcZ7KkvxfhfLhRh0zl6uqjHmezCA
k6cZYVgN59u73pQp2UOIlgDFbFwokZx9i9c9MQmA74UlFL89Wty/v+7SdgPhoa99
oykd2OI3RXRgNMbL+TUKYexXvi7lZzc4k7yQW+Dh+G/yBNtho2NTpTu0RcejS+xv
yQr8RU2+zdN0gAZnW1JepYGR8/75jeo3SMKxdgEuBOiLmxFzvR28xjFqXnyUk2eD
2qRndcsgfgGpPh5XVQOeWvb1EMSlzCWY2lBkO3vVteGYqhYQrIcx0uakfRyJ1PJ2
JVCk/yObPjDQ/N+3U5QPDnaGBp44vaZTUAMAkeKksYO4zE0tSfW9IGNYF7uEKgyR
5Trt6xZz6craXAHsy5ca/Rhs0L/GTd6d7A4zvmWejawsEjItdaog0fqUSAe8Lbin
x/jMOkfw9qnv7nmIzGklRNRPjNM8bICA4SjyAoYrqASV/z3wA8Udk5q9ufFHRR5e
NsJvgRyLxDJa6c4U6pRvjAAGjmlndKa0b2SqPMER3y8T3zqgoB/FxSRY7DtlFtSa
yGp6DsG8OHj8M5Ny8KMWio5Gtb4A3U4xiQ7R7rZAoOKEK8P9m38jY2owcc3/nlV3
SwyzRKGu6SIAm8VxVUv7GoZUq5q7cob/bv9xkcVhnl3UdmryMRh7opjYJ2wvBc2Q
a4DwwqLUNkRNQlKC893+IX7QE4bbl1NaP3Rppw3HrgbCY8Kvbm4esCWbd95Q1xrH
Vw1kGQwH9RN3dmg8tm90ZAnqrGaOMnwGzJ0QYuelur5htHPP4GGIS68ty96JW0UU
q5o9MkhyuLlXF2Bub5m2fK6MZoymPuuIIxkOaqY3dc2w4aaHiwcDhvXUliwALnFk
038qeqVjALixFPbD6aw3oA3Yf542BvK6VPbO7M4hKILU8aS8hT80woir4cj3jbaw
6CIyTcSndMMqXQQA+x/3Lzz5Fu4jay9KRoYGK43pae8lb1juFTLTae+TjjVbLb6p
fOm0n/krViAm5few5LCWxznaYYOvnIDzrvDaP27ap1c1yk1i6VAGV6Ej28Z/z0b7
ftFIJOmZFzGRgAk3W/Z0RzAGm0LiGJj26rb2WkRZkJ0tpDUtQF6+o9Rp1UDgadt4
nAM7RO/oBh6ys469+j04RecsObNL/D73ueH+X5UjqqxSZSMgObRktAfM70AH8Poh
kqj16EkXzxXlqqsUwtAu6LsJbHMoNUvO4E3t+EMcJydpoTJTF6RkXiDCqIpBIWWZ
bEKL9oZoSpduDFN4ny3XiSLyHsmi3b3zUHNd7jHp/5hDdykVQDNMtLyDNYtTj3DU
mYpsaHS+vGsdCeeMd8ursVUjSsxlNtDnPiZ6UnbKsyDSKkVNWYU3HbZCeCeK5Hsg
cEs/NFqnZu3Nt0/z8/epyqP+VkDVNLGA2ETKGlQHeUSMYnjJ0gKglfcqeMW2F7Ex
LcfWETk7JHbGUb5KgTh8cXrxQ6dmdPoYbEgvrUBsBL+5MC3sGLE/mdOu++HwnspZ
rFeANzvB9R9G+e4keiBKVINQjfONDQXDEtay//KVPgxHiuinkNEsvE0Gz2xWjNAA
Sb4vVsASUuRcX5nP5Tn7AO2IM9JBFGy/QpjNMSzdXvyhbDWCUoOiFV2Yll9ANtNX
lN7C8xP657RL+92Ymo2sp54WQypfbMpnTkU0T3NnnzGFgkIT/Q4KyIncKSfrVQMv
qWgmwQWH/FrkcM5T2mVYZupcvcIYHvZ59ddAUp9XiV74CKstZXipb/RQ4tlEOy8e
QcY/ZFb9geBvHcBChU5mC7nFAA0caxCsDZ0nlK40sjETXWmmMGt7mnruKTivHqsG
0beEuT7MZOHkW/kcNfVVsZG6DToQeIUA5NSTkSKAsXtKJfwnMeg+fYKphzjvNudA
Ki6q15t8t1izvwkZDounAeMgUzGQ0eY/9f9Q7sGkiqeeE6m2c6RjoiiuFvG7O2EC
fy+g17Kz5qED2G2AgcTeZcy3H//3TTa79mJ0JOWuBAfB7OdRjba5MUi1tOs/Cl0f
CPfxQXHcF99Hw/g6vx2y1rwiuAx3edOCYdzQTr1mjhEwRM7STyGT0gw2mAbqB2ei
ObLdHTtbcjj8k+G2z3TKg7D5gtzNKCCaWPnnTFCjzvKRO6jc1fxIfoUAveHBSBtH
u5aLw/ALtefRsv7Fn2jcCWPPZRTxowPm5xYbgaAYJoqbHncEm6RwnltLjSkVNmX2
KNLjPrykAjhXNfrNpnF8QS0gXEMzvdTfA+kw34lqgaX/aNfdF3l+CKX0MUc0nUyZ
A2jrJWYj6/QQBFDSMttrdvbEFLRrAWaF4eENwAXyi0eESoX5hiR4Z0dZP0Yru3wT
BKSruenlNjQUQKG9i/t6fzwZibbqcbfYsD6/V08L5hMTA9lcsGygF6V7o1k1c0ur
sCQSGr59Zvi30MgY0Cokkb5xoWckBYaUzN+grOrvQ4YTEWe11+7osAiaB1Q159q7
fPepPfER5PCzoDNowS1gm66Kjp5fITr2y1Gkt7oyDE9cHs98X9T2AAWxYJFjE2g+
drFgqQS1/FHyjHsduHG3h6pYtyY3a8UI6TH2WeQfhl1N5/8qgaf29qYyKSuoSC4v
n7xiTmksAJg5vOTapIgh4JQ7LUqmB50FHCd3G7pzTSyUtRqCpWl01f9FVXnv4MNX
a5vi2VCDr+ODLE9uCVE7/j/uCGWoj+tMZqUwDxtY3w5ZPF5zimwXiyiz4tEI3s1q
JYGCRUK4lF+xexS0Y44WEcmxTAbhfIJvLqWJdnofBD3UylDi+jaKGns4L/KqiArl
CK6EFButPuqVynk+SgdU7bQfGcWKLUjKER5C34Lc67OgNBMTrj0WEb2N+TTUqLac
n2FpCs2y185z6kLMFyNg7XkbKj6jj2ocCFB/0NzJ07hGxMP5mLSSZC7BOk+ADtT5
DCighiGzojooGOwnT4SlEl0WMPDZppZVReoQQHP4pjlHnFZ+lCtIkbzgB7ZAAd1a
+k18y+rIGgb2hCqaVvpGVCdA/IdhM6Ihq0J7KqHsGgpNrd5wT1epdRBG5EVguDBC
GvZlM0hVVtDkI3cLhOLDhXec3z5M2U3BMFDNl9wIsRHaicHlFoz2TrvNFtLDU4pt
Gn6UOKiboLG3L6I0H991G4EhcFLl4eug9xxOjA2X8W6bh3rMUOOkbnaWsN7ebK/T
IhFwlaSQZ/xEp3ndt5ZGiiYECVqCyuHLA8xuSphgFUlgfiYw5YxOlI3q5lyTl3P5
UNmvMyZG3BAkGQ/FZsHbMO5hSiA4JG7uBJJjS1p7ExUEZHGJRfHgq3gOlw+uEOtp
TuSN8J3xpIxmxHB4rBhL3umcaIW3sQ/5BQk5568ZCT9veI/9z6ytRbuuoEN6JZ1R
0vLPsYd4cqCLTkDUai2Azxk6agLg5yxsZrDNM/V4JP9ej0UUiaQCS8CH9zJ/GqZK
40z+zFThWZPP68NH9E3S9AaEB0O5matIXocc5Ky59jYTr+U11OneQzUaewQEsLzy
uJuO3HSqEdSSCsEMV7OjDBERpWgH3yl4tX+1aJmzbRCVWwvWtGGphA0Zh2hrbj+8
VEVV2TtXHxfk6Zg2R6Cs/2r4mhUBeMHcPvSh7mlc+2tJWyeEFbKVOxtrv62ZU/so
/7BhLyvC22FS7zEg7zA+s+D35XRmuh+FmXl8MPmK+Ph7F83m8uXDRbquqHdQgxa5
Ps8dcQZkPWb92KAj9g9wvuLfD5JsEj4IebDvdT42NZ60CkOyrLVXyPxrH1vSdiV8
zHU7FPiWtojWRSdD5ZvFcIaEltWl62rxzoA1jkNzntqNNxUMLgCZbjdcMSNVipwM
Emm+XvkhzGlgHD2z4HO4ZazQJh/y/ZqG/fe6TthY/0+YdsjLFcInveh3sRV01cS9
Ypi8f/x7eQRvZ3n7UsI2MpCcS9NJFbTYMUdlVNm7ZR1OrKETVEzkNAuFnBQQ8420
p7keQZQBBxdTpn45waY8/552+xe6A4KtxiXQYkzL4vWQTvBqYHl6S6V8WFLEZ/p8
BJb11GGtHp2pwhVjlZmS3ujq9e8RqwZBwZOS+vY1tDggKzH8950DsqLI2Cq0dGXU
Aa+EzJ+qDbj3IW/dcj0yBhDrtCwii2zQrrpiSvzmQN0PBFZslc43TdZ1Plgmgd0v
8jdmGmelABn2e+E9hIHnkkQ84dymUOurQdb2tiP/KKzXPWAiE7A6KKXpCO8BNS6n
Q0IW3gMmOJNZHsIF7oB5D1azJz3kRlM/H57RuLD23Gt4ak4/msz3jKGdmJlvIwOo
HqLFGtkJLiB/6/OBmwPNBXYq2KF6boBQXA+lo4iTbyPmyymmuxzWFbYZzpQ04pkJ
i+VJIaPQlHzCkkKeZRno6wjNnD5QDyVyjx4N7D5NbEMy/O9PT4Oil4uvkYXSXhYN
1z4UQAfWhDmSz8QCSZ+we3AQDZHJmgYLAWFy8DJU9hO7NHlKf/Z5q3V/ndm6tevb
NLrm/bIExc/JxGmOkod5SSy4lJkNhZg/z2zhH7RYALtkj5esjPBfK03Bz0R0dGTT
486IChn69Gkghci65vskvUwMCzJPxQ+1N1IgoqR+hjRxOWNTFV/Hqt2XUAW5HDA4
9lydX/ChdEaqmnqSw5A6Mm94YqlkEUEW0v+YpvRQiTb7pBuktCF6gD78BkfmGocY
+shXsmlXjTj2cLk/YFUR+vIUifIERcsjITIGfN1sO6EM2o0NHEQbrfEUt2uRTFgH
hpmCdnSm2NPbVffAkx1FE3azmnT5M6EDm3YV26AXGHbYL+LZtPQXfHoawNe5vp8I
2xZrbFXXIn7UGzZGeooFUFm+lccKAF0FVJc1aYweJjLOogYj9MJWiUCIt22/Y3F0
a7YGO1ca1AKCWGx33LI44ig0WDGNqCtaBLXBSwFa40f+17Ohx4FctqGkjBMcyrap
j6ZFkcWOQLZEIEx9NWjSh7VTITXpdmQI6R0/sAl7sC4VsVAcAKGxnRsH22sBc6fe
lOagf2ayTny2zdOKYbO0/Anreemq38e6vjLUWbeWOezG1eWdhtDZf0oLDD13kV5j
R0ikKMKueq9dXRJofH6jWVwAXdUsIBWw4YEdUFdYUZjF/nRHh6kheVL3m4mZTbTH
0jndnM4FsIsr++PRpNY3A/amcsCwGcHdIiyxsdAZQK1SRGU40m4icox3LMLkv9rz
9n/a98524UZQh4N0iDiEcmnRyjgF2sHgN3Ob+S6pQUdkme+YxE/n+UYnl8CRzlJV
Q3flxMbO4IY8ZN64itLsGinqBqCLBKyChotqW9gkTKLebQq7L7AiqdE7ipF5dpn/
ob1/70SERkzPdFb3WrRUu8qG/Td8d55a8he9fjCq5tPC9hTH2T5TIYzqHu9TIEfr
y5Sc0hTQQQ6K8Ts/YqoGgBA3nCFr4C0dWfK1Zl8qrjyNhyXxf9PGu5QIT8AdsEHL
kL2pK7GDUOoyjLUhRV40jTV0R9RIFYZlYzTvBhmx5A4KkKu7I0r3jXS3SuMzk9S6
Kw39zrBv/XUw0PXxES1ntcv4/7tBI6UVhV93OuivCwtRmRPJbtQg0tUyE/p6W/4D
2zoWzDat1JskyNf3pczWgBgeLdSRvT1uNm1OmXkWSPTZKIHKRSvjoCx2W4W991aE
0kNOXb0k8UjqzOVrBTHr1YFPcPpPdoW2OtkOCEg7GwAtbnjklRdYVlH477VmMOod
hdatXX59uvg7qRRZplkrgSzIcrL7bPfg2+nED4P2sm8PnIjKyspzFCngMW8C/aB3
mQOgBTQeXJYmIhPMBl3ecHT5mt/OnpwuCnDoEcKSJUE34BZQQDaV0wWGU5B4yD2W
pmUT6f54D8NxWvXhYhThbe7goPCvt+nIbF8K1mF+CDzzaSJ6OCynGuh3/gE06hqg
xJrSTPo0xQgBG/NobEvaDyKIn3Xf+nhZR0c5kp3B4VrXSUHlVK+n0ukpAfUlazNa
kwfveEoR/adwXkr6MAA+SnWZWpur/KUFv6md3qCIta7EjzBf/daKeeFbBE6rspRQ
ls18KlShBew1XKQp4RShlP1+hUwXdx598NuZ4VxtIvUIfUlDAp4GIdPZABflUUjH
4CgJFnA8qPOJkuTD+yePlUMBWJEnfTV63M7ccOVL/M8rtTiDs2HGIrjsAQPVvDnL
jYAMrcjs5mIOb4whcbBXOUu7mWz0AArYhUksvAltOpjP38vctl0j3hugbMpxy/7g
YIRlq0wnYQCu0nQ4e3OaKQGmZK2euFQuGtkgVWakxklNuCbsWFR28jfLo/+O47Qa
kvejVUciMQmYLmH891J6hazpSAW9lY4u3Vzz/wTvwuiFURtWrKNTK0u2vSSjAi1Q
/7gaj8+FE6u3gxKdIdEnbxdMgL2idlWQ1vLXG7vr+n1wX+fC7gb3cGWUCp9h2c8s
OyaXlDEf6/UI0q8DjvoI6LcSESqTtl72mYRyjmyMFo5Y8grymW4FEvTGXHNCSBai
U1ilsVoVj77vpi2bdtN0JvZuqd8J5Lcu1ynR+QZMmHOTUQp3YIwTLKj9WIKcaaGd
EyRx8nvL6IjD89QSqRkPws+YUccPfxdHKwzwZZqLyXnmuGJSoqC4sZFR6SPtKLyg
ao3V5L+g0lRb1MNNFQCX6GlkmcmS7a2zgix4S3HtKvHfSrht3WgEJSioLVgSgaXB
T8/Y9wcr7Me9WcJMBR2TEQQYIRMn2o3q/RHlcd1ZXa4NOyLwDcK8I76WLl0CZmdX
U8wA9WACWGJSkk9dNb05ibdr6agzf+2lIsZYY45wC3GOy/pGIvwE/HaHqt+HPvMq
fPabopmlX8Xigc8SGmbxGnuCugQJt01ghays+D0XlVBB4v0YR4ndznNvG4ccga2e
hrBciHdZ5+4scLKrUiEI9v/EUZNuOu4qn5lNmG9LUfjl1MuYIdnLawBE0OELNzWa
xLMIkdgxx3AIIDJpKJ2pvujFyC9Jlo5eVLKk6ARVWpnL4+VV55I4YeN4N4jl6PXN
4L37aakmROw8q1TJzUWd9FX0E/p/BWC8Wxsui9UBVYInFJFgeDqCstimj09l69q8
JxIrpQKI/rzXYp09ClKcI+8TcXDyPvqWKeUWoEk5sUzzeCXC7EdJe6knN2pxd4sC
QsjzXlJtgHxTyTxzWFZQf30l90I9q3d0tP85orLJx4krNCJ2bjbwNsecT7fzdtQA
8qo+3iOh8cadLr5JxCX+yhN6ijo+2VeUY6zW2jBLZgu0POEviC2OLsqx/fZyJtKV
NfcInGXPcWnFiXefjhthJko5/NHMBPY0x0kd8zaA1y3iCnDyz6pXmh4g7YZPA0nk
QwwSz3ujGXcZvXhrznF7WlJY2x6ZxN6Lf6Ky5V+LMb/BEzZSW0ALs4YzkiXJsSE4
KlTFMp7LlTVbAfn7gSUCak0VdiMjf/DKghAhOZB/mLLNk5MMHXs3kt8rOqsFOde2
wpUCZY371U4mIYYwaSC7TNK+NQ1H9TTCJnlWLXYR23USKsng4Wnx+KAS1Db17g56
XsSrtukeDK8cnQSvhX57V1Q5eKH08GayhoDr4elzV99MkTUwxAamUnqmpmqUqEpS
NcwM4VWmwMwbY0t976AZVq07bKGv5wITOmwI669jb0s8MyVoMsqOt2pRZSEfUES3
6cvC+Wl5hKExuqdCUivg3T8Dy1lF7Kq1l4OKPBQT3n1keSab9IVosr0P5HqGNeH3
3MNSQIrspUAJUyg73WI247T7FB6uCyxncFdX/EVnGmZuSh9n/MsnLOjP+KpXvWrh
ulkOb9LFFQ8PYXFv57RlLYafgflgWIaC4LG11qqyJvoovEVHk0GXhlXimhWXo4ak
2aZv3dbpa3lo3JFjxETZbYiRu9H6CMDgjHDIsa20H6DUcJEF+pudXeJrVCUe7QyP
+CsOC+zJsKEYN+UgQqkIn4SRjAhGVdgzzmhJfAv/xWNVxb3OqqDtxhDrhdhVRI+b
phCqS/GBOGlXvX/XhBbsBZFg7icC3lPzWHhdkST4j4nsuLmriIYSmWOnvbynVKDe
se78593LUKDb3OdtyUL5dqvs94BM3L0YUuDaEH5zK/HyO9bPICCVqx/aOVT7NImA
B30N/FvKLCp82DHrxQHKEcE1UZdJHKhDSJDcPI5tCCng0ZfeaCx7AwKw5zKO9fJO
ic+IfhXuKfFONv81ndj/t1OLirCEOFGoMMkXgompEi1Umx19prwqUV+thOIjjO6G
ibOjq9LlsELDc31lDkAXBsnK3IkahX7woavdsBDhS9q68veoXdm+5pBOWS1uZihe
FV72AHNY15gKefVCyOkdBP6KISjn2GDR6egsUwoVaAKtur774RFitVASd1TfkSBY
pp5NiM1MgG4re7aq/OyqUH25nVqEmF6l+RstNOB5mxOwR+jpVFwBWzUyfLjfz7Sm
xu11aYB1O7JGJhUr6wfwumj2CPnsNyLyBEuBFd9qjbJICfvNmCuZrjTamAwOj8rn
ee5vIuWCl7zwBJvdSkM4omHwBsHoXhwc+5AkfL3UJLZ0cRw35l7Hr9c4P9IcFG49
zEscYa+NIwn1/h7XIdXHh30BA527ODURaOrtJi5lKbRoUkIJd/MOd4s2P+kZCEy0
pgLKk8CLh3XKp21N9ZnjMT9gXOV6yQnnP1uoJRLa4Kkp1uJcYXH4wScVh84SjmNr
3VIl7KB9fyry690kfyTw5iCooIMxpPO6siLznZ1AtlVp+79DdruUI+71yVEgL3ex
sUHmO1BLGzVxJmmXITRBCKhHpzlQCFXscPEUpNFdS9ZmX+edSov3yeroT6hmsLXT
Hr13h4dR1+86LQNwHmd4L5TYf0JZq1RuAFMOX7UncO0dbuCePrYWci4nBh4ciUzV
WMubNr3DFIl/AfxjpO5O9hbRY2SyhAmw61KX4zpmEAipj82u5v27C6eC43f6J0Pd
afw8DZC0EE3PFPmfDwH5Ywu3viR9oHgRCwNJT/CMAXF5UAnhepbXyD74RU3RBVkl
8da+5VbbhNFyRfoEFr8aiveC6DwfHEzxgMPg5zl4aBh2cMIUKeTdqVwJ2XwoEI/L
0fuRnHBdaCTwf72kcUU68e8WCAGdzQCnokvrL+863kMCODP8q3NNOKYrl7xtU5i9
xgiNiR3+DNCgaAXWirMAPIe+GhaX5iAf6sI745DTblOXCLziC0PHouqYf6uKbPNb
c43SF1I2yCd34eU9nBFsx14xHpYvXtukbIg7qrC2V+gd23tJzbkJ9c+xtpWtyyt7
rVhbTs3izY76pGowvICRCKt6hl8ddb8JFlFo6aNsgZ26UudCy02t53jRYWs2XU15
KwD/eu8qLRRzgB7urZyN7rJvoRMsR/GXrQwqLnwEMMkYsiFzjvz2o9QB68qh8ShQ
xNJLLah2ciBYEkyo9uXZ+4skHU4Cq2wl4P4v2+o6EJax1HtGrtL+QDMrgKXNe5Qt
GyNxAMprW95ZwH7EFvCXflV51wJobRv0RgZWNzOx/UvidKWCDxNSlnQi72H53mR3
DGBt5m6qNLAG+iSRM51sCNElFaYSkLl3ElIUGyyJ2zrriTIi+3eeSnQqcWIxo2CP
ngT7oII7wPuh2wzaYbKdMAfW9sMwIr42Iib/nfApI4GS2QYvlGLBNtf7dflaO+GV
e2ibV29XWVDpkl8pwdxKjKqG/EI7F10h66BkfDnlhHnQt5q0MtsB6ox3EHShfYwP
K7fVEreFI/KfOEgmpzH1hPXJQSMo2dqGYOAZSA5WiaZNSDr0qkZ9RguJiS8FyUVF
0OgvNQz+DD7q1SzSPHleUIDrnHdPG6Oh0PKsJ+UZ65YqomAZgJ+CF+zgxWheddac
X9+tbMe81lqLKRDL+mn06xZAwlT0Zwd6PUVi88O6Cve8GSqDvRLdj+i5bjsa6WII
SrmN1+zV9MomgA4cUH+6ui2t6CmnsvgY8Gu+qx/LQK50oVMHa7K03Sg45Ze2e1c/
dyKtZVCALccL9GwWbyvlKh89fl17nLa5DtO2fSaGPxFXFVP9lyEgv0ga/jhm1ZMM
uPsvGevr5gmvILlXkRma8pXUNVHWnuy56eO9IapsmX2oITPK2fx/1pXFhOzNUAAv
ciMnjSdkI2rwPStOYUbp/jAOxJaE1RYneE6mV7xkH2bcMWd1gOH6RpAv6kd60rX0
9wJ36NgKjdfGrPRQ8Qhoj3K3bnNkQvvUQ5bmqogk5dmQWX0LTBncby+nQvkGHMde
Lu9XpgIuLhV93RdeJCdAFK0UGfPJ9npLeD5KDS7n5lCet4Vxk10fP/zPbLxjwWcV
2RQsgP8v740tN1uZ5kOKcOAQ21VKqNvgpAK9XLouUJQLuwirFVzkQdSyK2euh2XG
d6Ry1fXXJBB3vW5b/Qfk3g2d/glI76/eioAJgDgISwNcjySMtQXiwqqZhJmJA7OX
TSkqXwiAfV4m43cExOUDGTmpcxZ3TQVk+MKb76kRjhUZHJajfbI+LTd9WjBMJTaS
yv5w1vqSf8j9k0EaRB/9G/hq9fPoGf0HWWKNgp6sDvt4LfiYwyrSOjOyXKK8csmg
b1IwXfCUM12Ai4K75VKscXvxZqpm3MDVWCDXbhe0n3TvHkCfG1aPVYeqrQkChxB/
XhlEKv+QDdn2+Qc/HICNJ64G2HLnKG3FcMVpMEWByn7ZCNl7X+K4rZlktfPr64ux
q6jCxgNY2cWjpfysIT+SZ6a1jE7SziGFAHOcvR9EPyqiJFWRHVt9sXNYCMy8eTi7
nSNf9HjvE40N+dsDvu05fpRBqo/Sdt5y7ShaCA+MGtcBCzFhAqFFhBnPCJT4BpmT
1GW0Ztgy5RynQepPrWEV0g0Rby3oFp86QLfZoOTNZcGvtHWMsUR1S3hidVotVJhB
7W5A4G1gNCFJgG5QDcR7/ouGGCuG+ijHkCIv0oXdKPMj0O4LxAJm6A+WpP70IDnB
ZVCAs09oCpW3vZlwT19jLtX9p4Md68u0oPvGnbmtnR4ynFbrThRjIZs78G+BvX6S
nQGsnW76SMsrx0Z7w8QjfHYEqjhNl7vZzKMgWK4muyQSJ556Su0daHvStdPfNA/4
SJaQWZ3aUYLzvdeISbVbE5+JZGb6cN+3C4iQy2r3hePmrlg/L9j3WqrnYVzF95rT
0zpzLNLE8i8XMH7zxEA6PZwlgwEuiyjiLf4fNeYiky1EZS/0ZRFLbC5nDVnx2MnN
XpXbPB1gCV5kFc4NgYO7I3J2GgyKMcpLOBoJ31Y/n79EbTQhcO2TvBYpk0fBB0dK
0omxfDntahHSNeGGeNhKbLWK/S1QzeIBjw6jpYRU/H4kSBq2rPuq/dg7/lOnNnFF
w1OYHlZMrZPmokb8oelyovQWcuvZuL4lNR/4PMODwNL0cyIZJnj3FR98PNYhXxRi
1vi2JZlaazLb95chAXg+g9XKsSpByUN3ioZq0GTBSWIxnjotnmXYpvWkGBREkKhl
T2TMynXnTSYu9kxJFkKqpH9a67eegCFXHx+sauJKZMU38tfytF7bDUjK5YmOU3r+
3Y0q9IzYmbln9GaVoyr6cQbZximuqSCoerhjPN+XzpcKfdaLhhOPbDTyHf2mlz4g
V5Tk1R10hTz07/esXcJjO9Hm798EYAzBICtVjkTGZHNXRM3veHvPVhbE8RCZizh8
eFgyyopVMe3r7rBlx0jshyF/g3At64iNuIBl+Yqd3pvZpt4hKyFpPKb1ZbybZX2F
ODbpypWMGTJrMrmXOq9L4qgW5QSlUPCmJC+8yJZ+14nV/VlUp7Z2tMVfdguKukuQ
1Z3bWTc78ruLS3BLoPu7bIlc7LPtlqGFqwYY0qB1YN7WXgq7LSbbu7Hmq0+737Au
8jX0Z2xayPvBXV+iB3MYHHRRLMTMNEOTWHg7/MuH1DC3OSU73xFXtgRc6XM8XUsi
J9fy9M0Oa+Zl19q0nXCfdQy09hhlsB+cCG8c1znsmaIATjIEAybUkjOVB/GQC7k2
/zXAttB4/Ay44959yYEzJWdS8hhRctTzfwZFxpWbe3xLNcPjvPElib7kuYk8cMAA
9QCpLJqLcoZQeQ/A0PvFvrD5BIMLwN74KQXPgsslOIqkdODtfPU2wfqCvtIpuIa+
Zn1FRkT1vNnHFEpod54wgKQIcvThGJmzPIAyibWB+bYVTgyyQYWn1LZEzx8a94Bk
xW/FBasAl7RMnyRmRaTvhlNFdR1uTESB+1oMlLC2zDinEuPuQWhvnETRy4XOwGle
bm6erVGpg3Dl5+2ITo4FnIxWq8696yKA7cylcxJP666Isb5So2g27HsUbDh+pcJt
VUxv9Aq9K3QymBoCKX1uKTj3nRlXaiEDPdHQEow02ZKKiCEPlNvmBBw6A6NfSYzm
llWi4RJX7rHkiPq8I47YEapSnRuLzAkKjrksTAtcrXXAm/1JWN5IZopAgvF25aZ/
4ZL2PpHFr6kZrD8LzVA1McTKS6snkn1XciWogXEnB2YX4HvsSs7p1PEwTDgnsNLp
va7mEX6sYkmYWnvvLqJJ7LdZM+36hJGdFExnCezZ4yVIlCo2oXBKCvnuPa8NHd+O
MWNaG18umAZ7O9uq6rY5qjCO1kntz2y+NSE7bMklyIjg+IxdbTMn7yztALh5UrxW
0/+sTdJJRnATXMEANqCusA4c5R1wYPkWEjT7PyClSgvxtBz7BfIm+Gfg9reqT0il
LLRcEysPz7UqFc7Oim3x3xWT1noBUu6GyYAq6LEyHMByt1LWElvxoTSWjCL/su+y
eSVivSzbMDx3jludBGSbdBtZRAxOCr+aa7yyCqLC8zsO8XT/BAWmMdXrn3P6liWV
dnF+JtuBi9mj5+wrg6KUPiY9SSvQmNmUSuBZtaWMaZIOEXFH34Zw2dZkwihhgzzI
pTSvYqRcOSB4KXV5VCD2Xcfv4yCu6tyhA7jWYg0N5OYDbnS+qjsLc4rCAOhUaVxx
z75gi5lu017O90iV1J6ZYcqmaNMw6ANwFfTqJtu2v3n0rcNJBa3o6nbEEylZpUfc
IWDLXITxLGt7ZFt2XndMp1sPPAzXP1INX07xbB79GST1Rax3x6AC5FDdtqFq+oSH
FDCMrdeLYMTTMV1c88bbT8KSUP/vnoLvEbfJb/yJO1k4/Dof6n/u9BvONs2vUxfx
zo5fxb75MVLg8kBP97zpGN//pQqlOgVDOYpNpx7lw3Puq+4PVXQBWbvFfdNRmi8H
dyKwBJpSw/Zo2ntfDiSIY/t8YibQaHf5k9iivTZOy0NNgM7LPfALISbMW5nuUhgU
W/uQLgoVV+zDIMqeXC8f5URPmMwS4Bs8MV3hmCnpKTlvVoHq76y01XGDyZCTpjmX
cYqXKM0oOglb08te7CYy0c2gHbfS4Xtg+Ii/VFRq2vvCXEuuEGhCtJxzKQ3HC1xF
OCH15TdP7WCKJ8CugPgQNO5A9sh03QU4YwkSNAJtAKY86jdKNMzSXSpdqM9YJd8b
s600u6ybQPjIr5kCLwVLoxSESnefiNmckkPMM2pOEGHjrCxnYgI10Lrjk5aDNvXS
gJdJqb6ChjHG6L3ib5cp82z9aRpoKSM+V0wUkKznWm6rLFuwjA4nq8/yq6hAVTcU
OMeE8Rc9d1WNFEP7ZeDzsSwMXOSwRKXwXD8gVGCwYOAcnAD+vfDpIyv/1u5Rfalh
0EIlP93OqsqrwFtu7PHzwbqorNWmZPOgiqyqwtBgn9ExnwzznhDKhZ+H03pNFJnR
/kOU9S0bwy0F27tEJPRdvGhfg1jTYjjDDJjUHyJfn+mBw/k1EbJ+caHd+r4wAlj0
9LYOdD7ATEpQXlgdjX07FOK+7646uXLe5/lrBgO60MMbxq5G+yzZT3nXU70eg9mh
eQH8je22ZEUXUeHbRaxI77H2w0yW0Ozh3wSEarrJaOpSZdbC3WcjVTehJA7qFixD
HoTK/bOXvVGchImM8DT2huaB8sqFklAAAEtYAJ21/gHQw0nDsLqcOdYef35OinHg
/oBE1rwGkWHcwdVsh5cuMU0Me8AxxOlnMy1q4f4YwWdV3O6Yv46Hzm/Bj63WSAOD
5xARqMpaBIA+CxwG6r3oTTFt513z3onidi+md6IrWA0CFnttW4bXVaUfEquNHMD7
MAKWvlOzuryA6yg46W6mPEOPevptjUScvqJ+7zXQTd4PmrueroHvLaDm6yl6Mc1v
kABemncMBgCuulecf6aAk0CyNzh1iUvpwOmebTx8p28lSWrlOvlrMCD/HXh6PC7V
SYaKVzr7+XrKhhtObJf2wInRnzCc1S+QPqYoXPFHYH7RD/Ig6DpSoni8K1gQE503
CY8bvSNGYEhK81FFSOsY9srcC5Oqywwx3DVA1hdWz6xzUSXjtjYPPQ2L7GbYX/kC
pWGUbDi6WdvQjDdtMB3jm1/yX9dD/r43JClsASuGTO2qYgEgYUJrcOgUq4pscCMq
CSjkobRgQ5bK0F3SluqqSVO851KKmOG2cx9AuSxydgcnil0Ixzd39cRFKN2z53Af
qqPd2sMJ49wFkFU7UCuCTgYYrI2ZqJi+ABwxIIPvFowxlT7LTa2kTuOydJ/YrFT7
zE0a8M8KXWkq0EUgAQmubpi+xKNV/BqQetXQjrtZwXvVSwALrFVi251Q7omL9ABO
F7tkkIApK3D4xoz5VIXEvjzztc+Z/gJddUm/v5YG8k04KrQGbRWHojLG33rxtuhF
Pa1pM1LFyJ/6h+X3pJ74jjo0MkM5FE2USZpwFPM8puKN06138pnas1WsbwVF40KX
+UzQy9p742rRtTJ1kh5iWc9BCcp+NE0i0UBIkt3JnGaM1htSqIJurNWcYPkFAdI0
T5/HlQlksjf33/dBxXpYn6NtNjSmGH6FXV0FuUVFNB8o3PT8kL7qJJnjnf9g9gCj
vaTI4YKRloVuI8+odTEAnCwbZNrPux0nUjGduEPYfBLeKXmuZtCg/ekgTZ6zCVHS
y0n5ARaO5XBB9+7HIuMX/pgiptaoz6xLvZxk2XW56PqEKxAOtDrtWYCE1fZv8Oy0
1bKMxZN7UjSmGu/ztA+Mn7HCJ1Lat51JIlXCeoEski2lEBqkYAdNBXaq1aONV4lG
zYH/wPnKwpl7eT7FT+aYaXKewV0riPR8wMxK0zMXmbty+807nYwZ+bXJeB7ZM4ku
f+56jbKnfGON5n85ZOi+wS4vms1EOw9v0JxiBNlX+kdJynh1YRpkv9eK4Jq95MN8
ksZX/fD7ZSdiApOO5Br2NQNi4K4MuzVI3Q177UgMZGpV6nlfR03wXyyf2t58b1UV
e+ylzlIxUZMYSxJRhJ5FGPzyA9YioKRgxgEWGuzFVeoZQ0guzDaW8lp6dAPQMrsM
d+eA4VGj6D6Aak2zhMRZP60OWDgS4MSyBNmqD8SAUSfP2G/OXQlwl/Bk/LcHV3JQ
cfHQ7cQgnUbvXavqyR3pGx/mVnKj5UivWK7rs4AREb5gFdD12gtKIP6YbbyUv0Fc
o1jr8AIp7eA4GK4XNbn5PK3YenpHjW94Pk8d0yyyYvmvQZMmp/G3/S3pg3qUTY/F
ixKWMv4np9Pfb/B9yyswQGTatzaEUEsEj8/O7BzzCM3qxSkQ5fqqMEtvLylmenWE
zNKGrHTJPxesIvcN8cOl2Pqi+Foc08SuRqaavopzofUveG6sdk3IGksz7S9jpfgo
lIMMnQa9s8FNrkvkNjYT1HBxmYvWfKujis2UetzKQh4Qn71O0M4Q6glhgK06kkSh
Lgyqjzj0Sh8ciGEw7y0j5LdNnFIU7kCxI4ipddc5H/yZ9SALK/SkzUeIJFDl0HDI
+UwTc82jnTC0slyFoHI8vAmNyy0PZYcMifPwdOBsnq91Gd9HtufDD642ha/v6koG
5yFJo32L+0ZfDugXNLHbOF3QDcys4RougPmSdz3SSusfww9aVxudc/cSloV7R1Z6
PYgTYG5q7uyAs+EpH+swWNUb3ZsYJjLkoYFEIhHxx/gFn3BYGiwCTnqjHxu8NG2O
Rnny5Qd4bSS+FdLGmxkRwgwOfvHxmhAi+TSXNqrqMgN+6n+/3t0j8fTXB5nmFa5Z
NfQ/+aSz058LJ7hub/yJfQakwxU4IE9LqwTwPNoFpYle5kibCFiIvExEoAtLJ080
jLFlBqTQmNhL8LI8+6Q4lYTpUicl25CKkNYL4Xt8CPcH1RWt7tPwrLKnzJsfej+X
YwrDDJUkT8Q3bxf7/dWWMOVWUTRJWy9cF+WaZqqvQEyab6xgqpkRB3ADIJb+fRqQ
HSrrEiSFEJ4Ah2gaK67aQnhERXiuD9SlMJEqpneGq8ePj7w0rCc1t3YumrfKjo0G
6NSkdkQWvJt9wE2gyc3UegfdGXDJpy7ddl1XQbTvAGPhaBO70Q46JqNdJqOv2zVK
TylNbQUBG0pQQWCPL3wpwysrW8PusJYY0KKtpFwR5cW7BNiYTjgP6ekK7EXOkJaC
xLRPRVRiO9NqgQuhW91r47jcUtfwThlhKYaGwuHEQsOD1r3/veuYFYkPRgiSBEH8
HC+ARGzbNc6tHYvUeOJ1Y3x5Z1h1v9iJQzshO8fYwnx6LqCTkq6bWZwRX0Nw2kd1
4KbFVm2mMK1SZAJ+ZTXx+6zDuG3CgK+HfDJNni5swFr6aAFtB/FY04zSXlKfKygu
ukRFx6Nmi0wgEq0+SpsqWcnVoNjdXy7t2/FahqbftycBwJXWLb2kH4csvExgtohA
rnLMG+BO1q5oz2InNmqgyJPILuUoQKttTKjkPte6uRJwYlhX76OcrWkio9EPQZvW
NJfpgDN+A37rtgetKl3Z2vRxZBhn/Sjl/t9IVWgBHvyrJCUds/ZrOGP6M38k2240
cQdKRF3haJTPysu3v+NnDL+Us4HuTHSsHbNOdxlaJoUaypfYn2z3yRXtXh0+eGDL
9r2NauaLIWC6OyFObj7s40d5rP6qdv9ytFo7yWFOk6mma5PM8GyJWfiRWkScqkjB
/tzkj1J4M1h4UQNPxFRznhRKhYN6fXwovZt8bkGwBepXPfy+GuxxP9+62PEjbRxY
+59kif3Czpzu/55k/drk3DYC3xt7Acx5F3Xj46vRdxhkhLpxdh4g8m34TehJQ261
pHrlAKwBZEiLP0/Fb1cgiwIPMpfyjYbdu9DcwOpRWk4mWqAP8x7fI4/qN5xTNIOU
XnIQ4X7EXdwWxFJSzu0rfZmw2r57gP+96V9uc3Sy++MzFmUFCXX/lGNQWgzTdubK
LwQ/xIuVKThcklgH1jqk0/fDeS0vA1x0jKEYSLLtweDaiS0uv25QABfdhokmp01d
7P/joDHl79ypeiks+zsUNS1UAXxrf70YVOZxGeUKC07m1AEDCZ6YPceaUpiV5UOz
s5I9mKHAKwKWLmFuZUa/XjdBayNEWpJnAFyuOYTTwEzuwySO4pqY+DC2tm92E0OC
05oYKfj7GIICHYbp6hpPKdCdquRj0GH4VuxM7dikCn7rDwTNQvjFH9a0vRgGfgkl
rCpTzaHBb7sSHSk8zdQ4ev2816xVWQmzitzecZm5uBC/cPIUiBkwrQ/l4WLGrv0b
ZS00I+ocqvbwP8PZSoCZ6vztfomUBC1ohlSdG5gAcHmhHYtcpWXBAyfHb45lZmHv
2Nlbgtn+sfWR5KSudOs30OLWZSUk72MOlUtUB5XLkgy5U0nkeytVjanZfsNAIx7b
fxOW5LHuEJ0jchz+ZqbhtuKIjaqrZyrHTy0Gl8FjfzOC3ZivNSnbd2oKFXvUsGbl
7fjwmlWFndopx39HTcMJIG8yL6rZaEWZeVJOl3M++JRE9nbvt1b9k3xesUOQBiEP
t5wG/VH6DMihbXzEs9y6n3pkJAcGeNpJkS5fjUAmHeeeDIS793anLQisC5aWHvuf
lJj+M15x3QPSmec5OTbRLb+9Y81z4f6xe2Am/dnhLL9yIjlSm3k70rtcdl6F8NEU
p+JCOBHISzgnkPBUMcfBrcdHS6EJ4o0aQHzfzPQYX8GNM8o3xo42TqMmg9GNydm7
PODDyeh6rQMOzbPPE8ZeD9tNuxHqtyjtrNQ/qx4JgNHHLbfexbMZMrYnY3wCgaAt
Vdx0f3nbKNM/RRcYlN7pF8jHYrCJVSoMqtqjjYDeRmEmxJuX2c8hUeCS0nHJiYqQ
i5MyI1kDuHA76cU+2z5McKGlPnRVY+2L6ohQYFo9wZMLhjxA9HeFggZHQRZZ8mCs
O7cC1JMkEZUTmFCGK35xfx/T4lND61npDKMv9eME36UVQLXNbBvqi/YX+5wIO2s7
lW2xU9LIIrqI0vceFtxhytz9rAS8xg5Q5eG3nN0xvSf08Wns3MAMvXqBgjSfrqOz
AaMCxvhvh6RCsLEiEMiJKeOTrhAmdZueSZ9QCQkfXs9339cGOOw9Qz6gxtmpen1p
GKF5V1+naedMcqsD1fDVTLhm+8n4dmZWDlwtdfLtXba0cIIbGiydmTuZVipx++/2
36cZsd3lLZ4w3zJEu/uglpaPmEHctM8c9iXv9cTPkuLJCb6sL9SUbNlhAM7ShUmP
cG1gg0Zqt8xuhBhuDlFLGOa0ZmVJJrW5lL5apF9TrEgQyOih7i2rOsh7cZTFtJxX
Z+6qGZnhpyIkCpLbUdff3AFvkVQ4rweUprnfFc3xsrdsEYF8Rnb6OjmnpeKRoCAT
YQG4arfQyZm7Z6ClVodg41hGtDgl6ldDvsP0PXwcy285iokUOqdidvsmWC5Uoe3Y
UjrYuZKtvshvU2qtj3GiX5aXfbu+LNomts1MSaS9wtdcJDt37yxQPpCPpGoq0qC7
bnBkVK1AsRgjIeSRJQ6dnoLhzJkiCNC8/dLoC0ecK+H/wDLe3PYgdjtUGskWEZp7
qRmN42mPPLkCo1qMA1ifHKPWxtHqj1G+ctR6oHmV8k85y4ElO5XecLmieJoOkPhU
/cYpTduROHjzOHcNJJrZq2BjZaZw0lsL+mZ+3KYkYjMIXqsVshxhrKpfdAujOfJU
aYuc6R3w+t9YzlQLHm2E5C+uw4A/T391u89MPDhueRCtSuW49Q2TcSnQdsFmsq2Z
GXZj3z/bYLCjTyQe+doRoDqwdkmq6cCG2jlaYer0P0NiTNA3bS+eDxq9JYoc9WEq
FtXvoGdnXKbgX69gsaC0LcuUnFXspNLMsWPKRLuxdynQV8WerCqNBnAkZfTQldUJ
bg7hAY7KdOUiemovWYNuTswvo2z2URuO1UVN+RurUeHjk/qp9widYtfKzgbfTVhv
wUN5NO1QsqtYp0UQIEmqTnTyd8i36JNk+fWmgqjMIcJsiAyO+owSnl9Cw0Rn3Qt2
5CDarSNKcM9xYI5bhayQbjUUox7iVvm6+s+xuY/1aarv6a0LOxPTAh38x2m96ai8
C54hCGioftCZ4pZ5vkAmpdmakRe6H0tw633DADvQyC898zxENIFiKaPQSXqXI1iN
5/JqQjM4NyFaN4G1ZoXpz32cNrBDc8ItmZntvfYjmkSJ17dqjHTAVRzjmEb/Oy0+
l8rjWXm98WnLD2uMQgNplqUY7cfUj88lwM0bzmYcOfwH/L3P1mN+BFojesWKcOmh
82/b1qPMEyt1jngrvQz1oqQ5zMReNMe3C4zqN4Z+hxI8EREaOie2ynoccjNRSOE+
5N35AqPWflfau65LCNGWPeOrTUksWDHQdFUsCnUzDJPWWMTvLjR/7DXQuKrp2qKh
Kq20V3+yUrs/W6T3Bk7tieqef6lRMUEt2ftyv3fTtub7AibmfPS3hHRqBO59aEBT
Yyzgm9XoWIPHzkBqYwR7ygXoqNt2VpP6QqrAdNqCduKtbAEA79EQ/4ZktqzI/Zz8
ZZoPldm3eb4/oO8jkbyFoMbOsLaQefFBBEwnkJMZPATb1QYYJA0D/4oCcN2SbAEm
8l44VKVdkw9wcSY9KNvrNZ/15I3cQIAKmm/WOfrBXstuTvjR75yQIYSyIUkA01pQ
1J3DHAxfA6TrBaLVlZ9N9p9qNvIfDE9h0bQr06aoFQ+51ypbKVw/HY60xkqktjkY
hNb29OB26Nc2F47d4TY6iQJIU6TkWxsEeYh4w0X7wz7ynmROc1j2ayUO82l5rJkx
7FLOCUYWvmsVRAo6pq/p+EmJCAx7xuwWxPCoDZninXwVbmak1OIizp4gTXGJX4uE
aspUb8Q/d1SUc+vgvq3IAVhSlRt5c7N43/L+eq4DZ/z205cOZ4CxpaMOsHe37B2F
EmJpaR0efKatvV7X//TbNenYiL0+VCO/8RVoOirjF/fmm05RvsUEfxRZtvepFZS+
h6iWEWclqrG2r4v3TIG92ypzdAw/1DiyuiaGTgUbg6lE/hqDl1b84IUVTZA9y1mX
HKbaMQp37LGa9RWS+M/mm7Co9Nd7myUD/bOXs3/LruZ95FBmSYp12tYInlphkYOX
ieeoqvLhZBQ3VK9CLKmuepIZdUbNvkJi5EalpygglWPTuqpP0rAZ2ha6qW0i0jW4
NB8xTdmDWkCNS2rT3b0I1wU7Do8VKwHDmj2KSGgrpB9hbAYYhJqJJPI9uo9FQ+HC
gcTEuAudgL3HmCG7jQnTS/7X27axW3oltak5NMQ0ADzvQ3cNFaI+2/rK+h5908ys
U0oKC7rT5wW+OCkRNqIX72kCSwkNNmqxIUpNVk3ahLwfWbvuTMMzUJypQ0qpd3QL
A0Bql/HkVytQ09zi9FOe8W9DV+Ti9mvpEfe4cJoQUl5zOEe7vCiy/+mj1pvhpW0Z
ZwE2+YPOKDpWnoBWOgkNTVehVzF1NnNHxdeHrSEt/hMtyP5VnKG9uZrfQEwWl5W7
XmzbXQVRQV4sz3o54WNSkbdhuvlI06pw1gpioMQ2NLMvOWQBgQefsIF+gjHTqftO
XE3g9g9ev7NzOW/9YfdLb5vH8hd8Bfl386xGJhUQ3HpofdbH9KhcwBbj4jQwPaeb
zvriVR59dePgOooOJiEUuCYkJV6cpHhUM/PDR+BIowjyXbAWj4RJfC7of7oFrz9x
K85MFGQIYY0D1jM1HvP4Vzch9MWA3xIybt/edz1l7eObyezY1bva+jBpY3lk83X0
RPfbFwjJ4+noKGToIReMnXz3IS77N+gROpQw8iRraQesdQlYmciYGJ30GVvuC1M7
C+yx+i6xk3wsTZHSkj76dVEyH8s18dvmpXbjOaww8nKVzDjVoJH9wkxM0WfIY1NI
kfrhgqbMklIzGYPmLfJdeC+ZAns7YFGVyeykmUlSYe4uY3+WwOqbbuZCAJxlsd7R
ge/kqEkMuv2Ep3nsjnKB7y9EMEweSbRmHnYqLXbWnrHAH0ovc+U5nUgH7BpbC5Mj
AmRy/9a13ACZZEbrLh346oRpYh1G3G7/pXzNa4SDf9p5RlrDZ4fToP0JQaTnXRYd
y75GVpy8XWyXSkP1/SlXyRIxZgSNS8AqypmFamt2QThnldLepTrr+D57fIJ3bPDQ
itSboZiCbdM21EyQMgv6KN4FUFYfuuocR8Ol63TKzi0RySrobuNEl9nkIdNLPCm7
GjWOq5KkM49Zf0hl8+AV0Aw3TL6k1u+W5IStngv/L1f7Dwq7fYDiKUN4TpH5N2o6
vG3nowM/hLWX60/bUStD/66Qn+HyI6QRhAHENxG6teD9BVgO4MEfu7VtG2K9KmrZ
Tn41dPnwhPEVd1cxsXGq/o26d4gCXumf1bK3D1DohqPBxvTWNGxhbuZZYg1gqH3P
3vyH4nzs3Tx2oqvD33Q/aG+lhvZ2K6mS5EVbKE+6oFyxG5WEmyxuXzAxJMNe+4Bi
Iecj5c7L21juUWSdrrvulP0OkiCf9FQyPcRVEgpS6vYie56TfavlLoPjRUyaG49u
DtpPJlhXjU+bE7YBEULcYQfteQjmDfGO0Q59QzBU1g+DPMvlZWn3EuMG+lEolwHN
k15iJ+d0RpUYJygJVHhpadZ0g0Jypb9fNZ/ZCBXILDmudEHZPyYYMsTB9rLbCJJT
zOVsbf9sdJ2kUpQio2A0F8VJqb4k4MvBn8zOT5dvBa8jduGUuTUJrxwBOkIbNVFy
rDx/lkGYDysQPsIj11pCdrjbAWK2lv/H5v/l6mKl8v4s0bX//IxkHEs6NInZuQB8
9NGw73yccvoGLAzFpPtkkAVu/0xyCKQBMUBNGXXj1WhsNGD2/ibyaWfCCPQf1jvY
q66NgFE3UU9otq9uOoC9P7CEVGOHtzuCD4786x1Y7JLYNsjAgpNJB0UTBigVQat7
A9tBrRPxjiB02tKeSlSzXzzIgLsmxeRkx/ARhPjmb7bs96nzVDxBCvkdLc9zLzU3
+C+33ZzDYi2o1JeXNOihbbOnTiwJqdFJkbYS3npjQB5z1N0fWP4YpMD/efaWHpzP
J3l25lvcx8zypRJk5/tKz/otsOrPQLTZQfIUCFj7rvS+8Qc9g9QoixQfA4LM9XDh
RMweEJahAXwPqrVjFCTpTawKkhmfcaoWMPtPCJE9vG81G/m96nxOKWch7qryhgMe
B893mKGVrzZySktK6Adt4yGzhYLXVvm1rNJsoYEj7tkRpkZOPehg3r0SdlGvtfRW
6to9vTbOUGSjmGMRdTaoz7CRmhwBcuqV9Un9fBev2G5MG6+8U7y1YWj8e9mXNgdk
GtC44JKofUVqhqRsrySMvg6uI9Y6TLmDqoRnEvVysQrtLl1X0P9YU/yxZ+gC2xVI
9XJA8esqowsbeG44MLg4Mhg8i2k7f99zgVsWTFrNxg5i+GWKiO/S/HgGOd2yEj06
K+zOfmB0PX3ubiboQGs+mgFqsmJ3n+HrP4lGjI5smQIZ496aY0GH/7oLTU3GoIAW
cJRy8TRRkJik1etmwWa5ErrSpPW4KAWftoCw/uN6KFUF/iFT6sbcebEg4+aLEg3h
BPRN+y9p0jiMGPPvgCEn171WDOSExUSXWB/SQzKq7KT7ghmrMHIRc0MEVsmjU+uc
CNh7bSISGGvETb0t8vZN+rjGAKcGiOENS0q1tu5uF6/nwDWULHH1L/kNreGEhdts
kJEY7MXP+zchpkQGc6+2sYmnHzIrlhmHPkVbXrE5KI4JdBCu67orFbcZnkN4m+hE
786DQIhwafHsEfLBkWeJOvgiapuIqDTyp8Ir1bQ0gNjtU4VV/KgRyT/mkZTokbns
c1+cWB83tKMrBAWNPoxKtO8GjZVjBPDaOyIaU4wypw/8SGpx9axUmGq+9frt49B0
yTMdh//xu1y2jVE+WQ/BgH36Owtz6/4qEdIE/zV9GQtt5BQQ9OxZZSPC3pIivJhb
IZZWvAHUFtjiKdc3oAxE1zH1Y3Tr3dnc0fbDEBmj4DAcjgoRUY3+rY3Jsz3M9PYA
rytGc+6XsT4DevGyUpc9lN09bbxqqAAZh+WblWmyGcuV+byehXkq7TKL5V/k0Hi6
xXSiEbvc7+TkWD8Bto2jD4P4Q+XJ+CeZsCBPzpgGKvZVesor9YutIGSCn7pYoQfi
YqARE2sC61j7q4iga8/0F9+hn+iuEeSpuCtTNn7abEz7nNRW+n3RvDaax8ZEBzMZ
Ei2j4O9EsLTPOa58riugR1S4pcZhK1VrVhXfiN5y1izHCtgJaq549AA+rMkpKYDx
e8Q6TomAySt5xBCjxfkj7rYgapyeINONhb41o57QzHviZ3aGp7c7LGiyWrSrOHwN
9Q2uu6sIgIHjeZseth/F0QWRC+dV4oojwKkIOQj/3XX/y6K14Z00W1voDxggF9PI
AhV1sJDAdRO1zNax6t6jicYx2dLomX6XUaKojTVpjF6N89vCQ9q+tUF7oUeFn89N
q8yJulxL03e1LCL9lnD13t+GXn+ZrAMyKimEXTUXqoT7jGMhcTb8407XXLLFxE4P
/zBGjSmunmYzixbmheAczjVJRKLHKsIhTFpYXrnSQEV7VHv48ciTLj7MdQIl9MBj
3D1Ed2kBT2ZoYc3IQn+SkjsNjaU2m57TWtY1XkZQ3NBAz4wotFOnuv0ogwhJujYw
DoCYyd0AA00Y1zKYIrtuL+22Rn88Mxnlhc0ZI4awgWsmhi6DtMvL46CnNj7xgxTF
CGr94MrPwm8H9nw8uNfBs1Z/aVQjJyDxnnjuyXZjeuAG4Ysurp6FxlLYwNO/S1lB
U3ieLK3NldvNqyKC/TUoKI7rjXbs38hpM/CGL5BPGptDjgXBdivX21qbFKajuTFM
8Wi5QPWCYkAif9bSERyummxy0nlVouGAl5EViYz30WoPxaDw5rZWasrAuPDNlyeY
s2nbBK/eYpmdcdfhUUvbvzoDu21hgNsZ0dLPaK1Yq3+kvRlgdpp/dgoqLmI2nUZV
gCCdhVQvwBzIcw16+MQMXTov8ndYx7+jVLO/6QVg+IUTX5YZcc2v4lfmSfCiItlo
8a7mBhZQvMZcqzv5oygD4jJz1c8iboGKOuB910i4GFoKWuSAqr1D8tpirkv0geed
mEhsTL3JtljPx3XTAe+irCjluWkOtRXrO4hzuuwr4ZSVq+Q4oPRcLNj0yQmFWmzX
HMFPTx99H5zUrEM6uXD4z+CgSGKYTLNMXQKXtfcipJES2qyyengf8t+ah2CiONE3
ACmZ+1RgAz3Bv8IT5ahp+Szw7ptHv78C09PTE73DyiODW7JrnkC9jahk//ugG97j
MRRm9/p7rH1ohsQVQm9v0lgMar7S6k8ylYw3aPi9RTXxmWzidMjCfFyBvfm410i0
MhwVXrPX3B+iqTu768yI7IRHeeRftKWg7okq8/igt5f1jd3jqveWb8NUtyGXftYq
zwo56uri/PSCnd5w/NT3VJgKwgfJbQywFBI7XiGR7nod5wkIF+PWHuBeYX/aOdTy
yiQKqjIGsuFCN+s9vbRb002Cd0oS4hl19M+WGm6Kai1hzmsWoXL4PDR1wyIwCnaM
r4k5KA9w4lYliuLneR7+GnvFavCP1ipgTRgQYFEXfTjsrbj4rFN6WvvQNl7krS9i
lXOq03B3R3HVq4sSfnCRiItOICaPs8kRGoW+/KQSdZ8CMPK+sxOI10MiQFAstScD
fzo9Y5GHKsuq2bj6m/YWrmdwLQDzwcOFghLFTOilSeNLvd1uy+8iqdAAXe6bDT1l
mjP4BMLAzx1RmzxgJf1KpgbJyKJzuPYNVmuvX+gs4Hl6ugr98uMaw0v7dofCws5g
etaD6Kq9L6Ot5Lju50LbXe0ATP//euW/8mLb6umeeheJNeFbeALupdowkE+P5g9H
7A/DpamErRbWPcvT+UqRTGEfpj+0jeE0KTmf+zoN5D9sH3/tr9RPTadf5narPQXj
5L/rWmMVRLRc4T1IbPGhDUdShrEdzg5eTTl+5oszIlozb0TpV9eoTLe6+IUYssOC
vbhAmXlZ0jE/c9m0bAEBOzD4Eoi+q2IrwttXxHkWRfLsJb6BD8Wm5cMC3WgXX/oS
0iL8CyfoapOaLd72xn54z1ZLPQRNNe7fg6A/2W0FF2QQnoz9D48M4o/F3tVkHaNF
KV7pOFcFyn41CGYm3U/LMlDCxE8NxC2st7/NxFW9o4iIFlqY4A5L9Y/NSyjYeYZt
LlLywYtv6+0ECXDQnXbVm5cM4DlOpqTB9AUsTdcUEQfwgLH92hxmjs5qIG0tXgfq
8pVQE2NARVaJWI/f1bYT0Fwm00T001rpSLKYLafN7xmyAErH+2P1Iplpb8YTjIEd
fh8kyryAdRcX48iXvPY9p7iarqxzku6h2BzulJhN2sHSalktA7ZrEUYHcjcjAX/G
CRGzcqkQYQ0jnxxZJJ5SJLKBQNnnEfAbBz0gOyjPKBXpatRFv1mE2+0oxub2KAmR
+eNbOz3a0fOnjWNtCX1TmszFMy+bUvbMw+f9mLDR2WI01oZaLzHSs5RZAgsnWE3G
Za5zFcVOqwSCpiIKzoLspaKO7aqNi4nrc6up2VmOaAC60eUI5M8uoi+n5OgWKcii
7ytPXHR+b799+H/eN5GUCCtghIX0pSvmjJa94ULUej9/PstOgN604LiVB+E2gVBO
uxNZW9gEdKedbuBY0plA66XD4aYs+ErNwrGB4EO0UaMpc9sCXxNSHz4qnxrfT4VO
/4OKEUrJwIWRoYFGdFcAoblZtaklbVyvVxpqk5x1ohxgwgfCkCWy9HcxoIGjGDpL
AfgVwlJ17bgVbiz1K1wcRd3c7FwaPKD8Ny3hHEy85Mfz73klgNR7j6KaXefAP6ts
gl4S5xzeQaUdMVMtvSyUD6U241kiGC7PvBekXiswsMOs1xbPGO/UGenGQmkLaI59
k1B45mYW/UZlt2ueN2T+8f7clDKy0a1Y6TRj5IsglzWJi6XgqpFH5rNB7bpMe7S0
ySW1tsY0EqBA9aWP3jxQ/SrWgP0/wpJ+i6u+WqEaYQaz1P5BC+41yYoT1nnzRExC
7q/xjdsgn4o5PF1qlPKCYoumi3tIteqhaZcpNs1KIaK2OKWljUYBxnlVUR/CsD/e
YHvNpl28G2jhsr96Id0x0PwJ27CtZS2LXSArIjyXUCV8U5WKEL+OS01McIqvxQDw
s67cYRPtvQPA6GgPs4l/7+A2KNnADl77C9eHvjGH6FV4l/ioZZmdsi7gu454w9Pz
5kTRzy7BT+WAMXQPcf7UXQBeLayUL84IM8k/bGQw3nmMbpOMv4oj8EUywKD8WusC
DXXtl/oUlAhmlZco9ULvdATHFRlKUhZQ8+r6dwYXldmR+Lo27cVGnOnIQB1qRNFN
JCpProlhhtrHFXHwjRWeJTATaJ/zcanNXMzV+SDb9RWsf2Fu8gP+zLtXRozKRaJ1
40EG48KltVxvbkomQ2aPjaoFbsjsCU3JbUKtuYcPFTfqKa7mNGd55P432T17VtWW
KV/KnYsQO6uxA3b203SQjeDOVWwQuDtFpiTp47D8gQLpmlkGbczs7be3zFo/GB4P
EqXjVoVKrQOLyFqQ/K/+JyCpl9LWgt2p7TLdB6Yx3BBPagX8NaJTMC9czREp3Y0I
oLAnAVqEnCHYL01tFZRVui/S40B2JrE3oJuEYYC+trMzHnk0Bvke9W86h3xMBYrQ
FEItdQmI/CGl7vqRVSTka71MR8egZ4K2dOP9DKlH0CsduJoYnhyyOBkVsGK0kiP5
B5MDaJAwVl4u3RBaD3j0O3hV0uyfaEJihpIP5VZxlESdy9dy3VqFsRO4G0G1bd8U
o592Dy6FG6A77aOWLPBdwJ1esUpY49VjVAgDmIGLfTjr43SeODUWyTfklaCbCLyS
DaeqfT5k+nzw2EEp14GwyGoylaSSBhhPAr4kXr4bEjnMGKL51hjZN+RdgDb/WJrY
/Wg15xJtOG1ZQ9A1a7+OWffIYUwfJz7lkfSIWlfZaVWf0iYH3rOsxjuzTv4jlCOi
/lyV3/RfEjAR+sBkrBZuYblpFR5qh1cIyILMIWjIIP1RDWCE1+Kf//7P33s8b93t
mAGeY7Gs3YznfIyUXx6rQJoW6b/aGHD8wRXOCv1nXM3UtSlBqbYVpr0h6hMnwLxr
JWOu3GKuEGm2hmAML0ZfG4eh+vxnaAg8NOpBxU57gXN0fen6033mT8+8QuBCJ3hP
xWMMLI5HE9Bv2bIYuG6cslFWEC+xh6hZc9cnEAUmiOlyvK09gKgbUHDA8DVteQpP
3z6iCbyLAZr7cJLegmUq6K9l7CVscs5qYlCbOOQU6Rv8FiBv5MaDDh+xW5hOhb1s
eP7fv2WcWqro7++ejzC70+T5ISAWBb29y9qJM7hlYCOttf+YTtJstNwP1RtKc8zg
lvGoJA+iB9VVv1BSAcgFrYuzExfQPNx2xdAVEy1g1hJyIRMwr55d2Bj4j8awQy8I
zqtRludwPpdyZANLsy0rjRnVt3lBodq6N1KFGXHp2D4tCXHE+fvIMr+xAWfFpRob
FopoX3Ax0iMNluhSrU3CuqmxNpyVAbg4hy6W2AG2Qp3HvjpTj2Q54RXHZAawHXt+
X9n6efCtmEY+6gI1Brz9ghDt2GNdMukXNnfCOe87j694m4BSWRxM7lPAUKQRBJja
7x8vEeL7s68G9F/z+JPdpPVnUGx7skPpE7F2/60bE5fjBHsbee9jayc/r0fQhnqK
o/CaVaEwYBzsHBW0YliiwtA53l+Mo/aLkFohxUMHrqXtbKOXuOgeJ9p9rZ6xwYtK
IxDlXbyP5MFAJdf8uqkShvl7JPJRJga0IZ5IzTJnMqd7wQI4FQCRVgEGtJb4VQ5T
AaA8VDI5nB6Lh7adUhO5rUvAlIcRC/fz70VO09LEBq6Rnx4snUv0Icvfi41mG96I
dT54AyCKW6j4W2mjftfWUKQbNJ+LjnMsv+UeERst3008g57c4tW+XwXED0z3+vqD
xBtQwLndjhb1S3lnP803V8TzCmj1Uaxn7UnelxnTA0Wy1LYUsxMRCz4Bhnj+sfbT
f/FUXAXEOQ0UESIIgTvyg/r+htbA7a62rZyeVQz9+CLIfRauFJLY+RLQnLa3Ba72
An1cDlOdINQHtUtcvzRu/xdiWoH/G1Dlv2dx47L1vfcopNktyeZOrcl+C0ux1C7v
Zo7CG9fpJt4ba2/8dguVeCcvKuwdML0PPJWSD4cB/JM4j1oI+RrV9qrz7poebzWu
tXNvkVFehidsurb7kmb7D8CHEVpdPg0WSePhlUhN64bGmhy54gfkde8vNQ1/ApJm
44UMGh0iAbyvCAWTcXyS+Zaj+OZn2Ck6tDqqQA6QHsZxgZcBhYTBucmBr1h6RfyF
gArVb0UtxXfWL8xoSnYRkRKIFO69rt21Jqe/456PTmXJuyaFllBiUXozqHtWpx2c
bEqpSfzITQVzUWYorOK+nUph3JZazVwSKocotnpNdOPSIdB6MP0VjXbZMINmqID5
7jzdobciH2uwMyzt8BhGZajvpF5Jbx38IBW4+XpPcIkK62eHLm3DEqn1+dl1uYhD
UKwdt/0mkGeKn4aQ0VvTzPDuk6lUz0Tt3pYEud7qz1Pdm3tqbqHeb/af9JAnM+mH
Auk8V4rK4iczA1OfH4PRhN0KV6SV3W+oYAAxIlxf5wSJyx1XmmH7DOjUwDPZI9AP
Z3eLX7uQ2wazDcRWg4TSYq/frN5waXeEEEo0hOldECRpvO4l15BMglTVKQfxClRH
FaURRdA5er6LYOejd2G1ximhiPUm3U2V2ZMKJtn5pevfUe3EByMHT9mtl+tF91+l
Uazilx3Ar7fFWZ5EPCMEy/p7SjxpQcCcT+bjk/cBcIZqZupVybKtpZNE5GazzOi4
IGY055Owqf+D9n7LLhkoT7lybf/cK3OiXcbiJCo+T6aKLbHOHTu8IYZJePstcxrE
XtTFtGVXNys2RAZ1vTq5Qm1k128bwAgErnEaI2+KFSF1XA+IUZFW0GzxdN0Yd/JE
To9umj0puZ4O6eNZxWG/CQZu0G1pF0QLEfJezSYoh6rz24/dertbOelTKpT4Bkcw
GjFKAZh1HzpnplqqxH1oaKYpNShotGTIo2sfQJvb0T16uxN9TqEpAAaVRD03JgZt
cQ4H7EHiknksyLMfgnc22sWivqiQ+f8QLB4DGA1Qb67LtROoReO+B83nbADni76D
VeHDcRv2dBE43G/L/yi5M29jyuGE9f7fRnntnriQc1e1GFPMV6L6cu2vpw0llQ6K
L9EoaigDdiUQ+ajlypqMP8JOZtK25Am0s6YzKhzXn2tJYTdDLNdZItX6px1q6K5G
gGwyXKdGAmhBYxiVBdii1sBsXXqmshVX6C1yeQ0Z6pvNFEsddIgKco5zws2sCZWk
4NQxlPFp7WKdslleWtOu4bJ0/c/DuO/WB3LStOSx6JZ3BDirroKWpiQCkr3UCdxj
laHwUjuUrO3gxFoQMHnspaOWqGAXBTizvNcIzQkxOP9JRoxfqSb8oZIx0aqmFDo9
/VU8UHUogvqCjdzZIkKvorjeoh2QncW33AlHxOn9xc/JFdoCI5cS7fBfmsk61NMP
kyxy2j/ZIsYLUHPK3IWvhxLGlzz28Dov3WAACLIxk0kaLor8SXDyRh2enLTiqG1M
rmYK1BvRWm1awgf34l4JVo2Iq+EIsmW1EJ6j6bH1BaajRFAMNwVoOBMNjMW1kAGZ
xP7X/ZcDraI4kaMO/s2MAWOMhvIGPDMXlr+Q+IK6BkrnZQpo/+pBYCP90oyqW2SI
uPjncdzO326KJSiFeI1tNAuhh5gk+VkCfRwWwE6RNiURgb3bNO3oLSuenmyOmaE4
DDdc8NZT7UMrxucIIgdygFKPITHKq8qlkdoogtXf5quU/lgY9gJcGsx8XzYHNvaW
euNVE9/tQc7rIod1QugZTxejfRQZyv/gew5px+J/UFanp2xmP7FTQD5RTyPklNyV
cRv1LodUB4qetxxYkye56hYfFKThwmB3qyzjiK4YqtCJR7JYiqHiaIWHcu5afB7+
n95BIlh0089NlPSH7oeHIceAWUBzytC7SiNnNQPCEsfV8P8B+6aUreEtaULlCZV0
iY0mgxsl0TAkUxsuv9SklJed1WPEX2Ju9SuO+Q35qG4p3wogKvj4+Hybn8/82ek+
RmKh1gA2lLilRLAEqL1QWUQ0+39/ciyUi3yvm0TyPQEBZgsXHY66r2oqoncKn+xw
IRw9c4kzabGIZ3Vi8Hif2RPndI3y59YdlJULBUtxQ8gNDvxK6VZ7cJEy4Xau9Wv/
pVv+l2mYeOCdPdpsD3uEjkZXrfjmPvFJca+ftC5tHcagViVXgQpuOk1/EaXWD/Vj
+BPUyjti8+1aNW90UlT7GUdsHHaktHztezDTqfd7SSPwL1by/fE/TvHRrX91AXrZ
gVoW7UhCKTHXLWE2tBZaRhg5JsXTxoFAFi2G01mS9ZSJRAIlL80sX/Tl2E3Z9JhW
7ejXPVA9HIad7fSYADpIl3B+HMfVeECzOAAp0Eu/wiVwd80Oc7l3stFGiB/RWvAD
PQuihgYU/EGZdTrY+0O+OG+uZwvbBe9sw13QJBWKwLN3/Ae8sxXWTp/TOsuesASM
Hydl1lG6v5hcQd/DIe9B6CnI4/Tti+twoHw8tRpPQWOj0Bs5tbJCj3RVETAb9SfV
9a2NGeuziUpj4rTXXPBPSFWTen2BefjcqMZP4gs2Q9cbABAQWAcX3ILrKiMAyTfj
Yc7lMXH0R71S9BJIxW1G9lgI8lyUO0sOJN+ly1FqpGwtJWJ4AkkMvr2bRGB/mMI1
Peds7u7ZnpEkXLaVq2ofAMuxom3RhOMowivJq0oOYZTKih91B4Er5jNJitA4wuFP
J0OyoZfDkwUez4R5DS9KrPlkI/VJouP9pceWjDOeskIVyiWRPYS6T2YYMh3OXTgL
hjX8UgUlVhM+KWJiGK84R6y6BOuBXF6cKSxJMLqkD3dwhay07Upuu6T4IVPKy/Az
GV5sp6jcdzBoq6IGcRhapRCns4GCDRxIUnHqoKDEjoDzLvdYQVIQuXUm/AbSWsAn
Bz9pK9/O2/NRerVHBQ+FqpKf8GaoT0KurC5iNkYc9uh53IEiBRzkKrNWHkKn9OtM
yS9VxLyxo5WQDyandE1woknT+2XC7g6k/rTEgCBKGeqvaIcnS09ItIfESY9EFN4U
Vi0PjduYo2KLWihGv6aWlALltaQruO3mzbGwW/sK1SsRtJdYSsqVMZqQNFYQxb7L
BaS7ydyoSai9WBzP6f9uJB1SkOxLIlqlOQaZXl8L2WAiuERAQDASmJVuERRbBYYy
8h7ZivKrS2Xi900qSd4dyZkXnySyps1gbwrNGPMnYNOYsOKgcaCEtB828JH7gNRB
GaMVDPX25hJpvdzefObPYQkcZK0a41Vjrpjw6ZVmpNznlyg5yV0fT3qj+jkN2gw6
R+NgBbsvPJCygnRyeXiptj2NHBi7cvmvKQViKGZ41k+U1h8VN9wnOHWWeLtTmddW
MohvtJx5b/4If0EpSG4DJAs7Nvh3u8zWV1roGOxb7UyGFdDmfDiil/J640N8xCun
mQntQOPreJqMvSa3fMr7ZqyDbj/9Ni5vBiiUbQm5nhv0eyeq4Mo04mtO3gWssOKR
M9JtJToGlHRt6MZQvibXOT6TYZvsg8FVlGrZUZ085j+XHdCBWi3Uca6wwtiCbfiK
KoQJdzj+f/N6OxxdlVSDh1SKbFID3mvrAuZHkE1jddj6A/QlsYPCstUk0Mu+BKjy
Ba0JK6kLRYg/trbxE9KHbngp48q4w4HcYvH1KVjxyjDrgQ3gkaBottzJbtBC2SHn
BqrQSFdBtQ99Vy108Y2/uf2GMF3uNZ9k8KM+c2KCuVyWZzk/yfaQ+9FZvM90UAJa
LKdIbOoaJj/FQAff7Negw8qo8arBQkrtd81eUNtbteaW1WX8SDweGvbgclFCrJ/w
6rIK7e+xB+XEB35AbGXaGKNuOY4DqnBNy+K7kYjiQFIGjti+55p7w0Bi4XMDVYbQ
6lXtBzoeJnC/oMwUkVqdayWfUk+cqRDk3W4pY0NY26e5vF5eJNJZzzQWBBpaXGQg
CIZbJtUg1jVjIHXfj/JFii4kA2IhK5mK76BM0WsEWbtNh2HaFOroDdtrorZT1Y05
KLVjm7H245QouGCMu04g2FEfFQWuXpM6bYvUaUYiMD5pTBFvA3E3K1Hp0diyXC/B
VgnBLEpPE8N9kreMFoOd/R6c437pgAAs0XNGC3eq3GrYPYcK0IJtce4MzeaIv3oc
bU6VrMkqceM9Nt4XauLm9oz4Jd2YVUaiqFp1pMFf6fPmwOQl24bLY1Fb7Hxa+5c7
yp6FWFED5t/QAB5U6UKmNROmqtZYGsE158MPT6Iaop/dB704eeJetbnLpui7tTzq
FmPoT6i9pD1X18T1Tu+pP/wN9SZGG/Rn1vTGgOxCS+5RgrMmxsZDsA8mBQ9ihMl6
pr4qjkM2+dYBzj78lnRx9L5zuf9rFu1M0fayZc4R4DJTxfOWTZ6N1BfJHZj2ydSF
Ps0T2J1J62UHO/S8YY7qXYJ0fI0VUwwP9k5+W4y/LsNSVd+CBmUx+t2s/H2+p77y
za1sj7yId+gSpvHlcaTuRnHh3Zx92fulUM+ZCB8j+IjIJ2AWr6UWi40SsCwQBYUe
7F7saFdB9fo8GPkrPwihbKOFRL++UppKi/5tU2dY+1oGISsGKBv2LclYzgFHU3Zj
MWrjiNo61iUW0LN4seNpaLzWqiqobD7WF8ABGU3orE/NM/EG1S1FzeaisLTwA5LB
CHlfaMhUovSkcAeFTiN701/I6ZGVyD+bdppTCb8x5SKk8xTu40GtkLe45zS2g1eJ
AaQ7XKMDZWiUL9txnDGMTlDciuAE1Cj7pgIwl4c1bLFIL6yIeBFo11WCInBZ1T1A
aQli2v7ewrMqtYodzs28a/CksM5dxeBk0jiqoZzU+km93pFjvytRSexhAk7oeEwH
hzVmFoTYvRuKqaI5wMKiwCIjd7DPyLAORTiGqJE0NVbtrYROVw6YkwyryjIGbBEs
SgAUG5WFQYBTy+VdbFp2LpoEu8CMqnjCi/rwz9Rip4LAww8/HvlKhT4T5AQQQdUP
vqkNgcPIyI5rF+BdF8CnpPH5w6ILyzgnaFmSrw6hs23BbJro0Y8g8xfkG8NpPxrr
l9ojNsNzhWge+o7Yh/DxffRmWwLK0wjaX9heXR9TddWuM/Fxa+syZxb+MCGHsD5C
XNGSyThr5rw0+dBPVnQO4H8P9MAC07WNslXqUCQgjATv/8TvqZDvHKCU5R+2/G1D
Z1UrBWSOPlEjoUqo0O+h5Ed0N0iVDAkBRvQt21Qa5QzwRH4aXGTzQnjhlspGVHEZ
qZviufDhy2KvGGKtmG4Gtlmqp0cMZ4zoOcRcTjKNfWy+2VtFOHTqFfTGt3+TFQ3k
+WKMdftGZI2kFbPklW75/W1ytxF9ocBOb+UncZ3H0qQ3RcKfXddg4nKGqWGf9mhP
foX4Kmn2TlZOMLqWHO2+omCHiUFGYSzGMDR8umubnjx+ibkzyyV/ywjvYnjf2m9i
7LGkrxNnsb4F9nJH02OgbC2e9wV7lXaz8GhAIqinPcCQUBfzuV439NAAoDRxWmje
Ft1yEpgVNKOjtbDVCfKjMcCIv8Ty/p3BGz6XuVqIU0V5Rgv1PbnY26L34IQmb6UO
qLhkogfEXl2XMJXp0Os1whVXmmgWWaSuJF0xKX6bJQ2jEh4ITMulPjM7asdo/AWu
QXeD4rtsTL/sgX3FiL6z2JfCck3xzQ2cpXyuO7DJO4Xxt5p6fkj0vsA/40nqvBDr
+QCgfWA8WX60MC7Smi/CXgA1UjRvc+eChFuV7e0m3Ww0suU8EktKCogJOPkGMyXZ
+7Pp6569FpfHq65qoey7HaXEz11KMEkcL+iDiNRCdUNSaHkgGKraLBxDy90LKH/8
FtznTUvmJfq/r0jwcVCbkXfDmGJFFwqLVQFaKSb1wiE4tjuNUerNLH7geivBXb6D
WK781uUIa3pwMIIDxFLRwxsK0gZ3+b/gV8M3spEY2BLS66UPcFXY6HOAR9JzlQhP
/Y0BxFHT35S7m6Fd9Fp8ucn4sCyi6ge1+sgGBkh6fVJ8U/YpN50zVmmSP7Se4YiT
L3yaOi/DfkQ2OAaQyMMrpqUMe9+6hnvc5Ej899sxVM1EmQEB+frkftyaBqHAhZVR
9br9n2Vu71ousGwLMZHSiWd9Hk3PTbzT68RY8SDqH8qWZrGBVWwh85tLuV0f6nYW
2NKU7gsaFPRSdID6c9ZmK+X0TZWLwQH9HT9oVZzhQ0rh8o4XX6A/LUmBlukRKG/B
OxUHpiMZAxNd6RkzSYYetciV3uz+EQWsxQs0cqyrmLDo0iUyznKZMeljUUJW77Qt
MHM4wjrMmyxJD7Zowj3cXbdtdiV4UKDNH976EywoGI+8aAEOkMv9kjQH/aKoukYK
C3nSLLnNTFZmf+v9l2UnBUxLKCZhvn47bgA+Z48pXewIBcvZ+T9wFdI5/ySJXpLJ
lGQYJWc8GeqZsYS+H6kaFnrQPWxqNwImg0QlcN2+KXZ0cyXcxIvB1JvxEf0LqmT8
DOPDR+COAk/TdzIaQ79KICmQyCUuN4ItHtCTk9XYo/GvMU8Lg12eZNNB7x/7KrrC
DX2WxO6aWSxKcHvVhKda7GgGajOudhKM5O93Kte4Mgyx8wY/obLV7OXVmF0Rov6K
smwattuFZ/4wW5JJisUlCHBC5cPrJ7uOf4jRWn76MPteKTEV03z8vqcd5N3Fs8Eg
wo+EwYqKiNKYqsGboyqRfZiyUEE9WnbwQthdRiSTJzW4JOPzBwyN6z3hX3ptnfFo
4i2GdsCSNS6+Q5SE5J7SlqdGufpIfSv/hQFDsy3Z4SyRd/UDlRWkf0AAp669t4DS
j2yokcgbpCMZVDgD/l8TmRP4yqOiALVJX1H/ohW93S+jLH6vR/CV/PGpvwNU+whQ
CvSGLAcmXn6SBQ0SghtpQwUXZn7u+l2uySGWYmuqm2xh3AAwVnCLCia7iYnnBI3n
TcNkVGu2AlSv/6suxvgQNVHZusSA03vUNZFTruXVAVEu/Ijl5WZmLSermR9J9shP
vxcdE169Q0Cbw8qhC9JGO3wAFJtIDYHcNdVVSkAJWGjQtszHpAaD4Pp1gedIRSoY
7mjB74wKsE9FT4HYYKBB6pqh79tPbKyiTN5F7UueASJOAgcamlc0gc+OlHwtIHLX
G3kZpNKKgNXah9K6ZlJdmOo8+maxkNuXewy+r1VdOPVK4CKNDuVKCScQG5266LFb
PcY13zYjayER0AMYTHJJ8Z61wF9Tx4RQo75M50empq90qq2fnDjJzhPslgj3SMbr
C+bhbM0MIEFLzY270NBsLaIJ3Krmeg9gIVgkVnWeZfdo9RDng0ROrajUoF2ZqlZY
GzYTKPWn0FcjG0OJDokQ8GErYZG8+198pgjY1bluzz1odpY6mi0PwU/SM3iL8/h7
eIH4fBGVJiIZJ552z88Z/XwtHsVs/hhczFkkAd44LB+zUC+ttbu6OcOiHehty62i
2ybbMwFgqRBSasW29HR+5Mqgw2PW5XwI1twZBjniLdfkdycLaFby/9o3lCqcyLRQ
S2BwiqJNhZ6vqI73sO3ryw+AVqP9TGb5Tie7dMnIRUePySMh0GkP6b5+aH0E2/yV
+n2AQlnoLzrRi5HsrxbrTr6JPE0Rsa3o7prgRt8bhmqCy5HvzeeyrzIqHcM8PWDD
7DUVgDpgpU4kxfsiIeBa8LRpKrIpkUXBbTlSUySfafqbWj16wIBxH1Zdgadncg8b
6mzK1em0JckCjolqd0mPJCvzEc5vtPyGnPfdk3rRBlpDHoA7uN0rJjJWU4uePKl8
/VZQ7H8aOBRGApuyVLiFiedJrwmAW4tHmDcUwyBQfQZRByz1utLPwpBL0C6gonyC
1eMDJg3tMebA6uywSZ53LPwNW9khhW8uU+p1UVVSAHWx5OzMoNQWkOHGvLeJ5Zec
baVL7D4A+2/ib5w5+oAjTtCf5sHU2L6dSDn/Z/1KoZhhXq4i2gX+zATAIinBEVJU
/aiPRhvOK/9ds4oMzwPvuqmyqzQ/th2+8e4nb5sS9RCrWOqlRLPuuL5TJSl6yAKX
NUFp8JRYnaPaKEj9mGkHTGPxcUwEy18UpQdJFiTt3ynFiKykPlqOfyM8QaZ7auUg
RSuc5nuXz4q0XO0kus+lXMKCFqBRCLUFcVpsVxs5BWUkwJhdS2tES9OsIEYNSAFh
0SFE6EJjWvTjAxv3z67q6/wEbrDR7+u074UmIyx2NadfCHPi/mAlf3egVNN7HWNX
9jNnk4ecfrsX8ZDV4UBDhGMLmjgp83DznLLc50sSmBCEU/I9+JEc+ZZyjG+ETFm3
kEgsF0kvRDDDIF0NdvMgASptGTSHPPEwSLAfjIt5mEl8cjP9ZoE6HK+tTj14vh+4
g+rJFcRvwUjsuvCfL7wtwggajv4tBDKH4r+yj46Mxns5e2+7zlxqCFo4popCF6Y8
2YxGIZ2YfmiaTEOAmFm46AUMcP4/ow3nYpdxlKezKjCE/hM/nlBq7D8XV3lhW/rq
0V8UWmAs5RL4je7SDSXyAn6UYc1rz24TxzRAsHYAG5M5J5R2/Jkt4UIz8o+Fh8/4
tLbSXYWq4/Q7y6ttxTYq4cCmYaLKloUhj3avtZvm8B+n4KGrF5GVlMuN50eDwl+T
/pFoI8wEcYyvS/nv/8dBz3+s7t/JVfze6r5U+iP94mU+DOGD1ZPWb8+RV43ZvQau
IGf7FbyXB9RVRT6ZcIRqlA8dw6wVH4btOAdYgCC65+DQie0GVL9KVNLYPMKeYVTU
E9nB+RsDYNEgft5G4/3ylBanEsVLaoxFhd2aPGFN0pF+IbvBYZ4DLzK32riFfimM
D1716ZvtVk1YyEGgpuxsdTeS9EgLySc4QMYUdrHaxSltrzOhRfLyCgnmHCVsshZB
UCQfyC3ar9X3WOPSP9pvgubq5IfvFoZUzEvo3XRscCbQiZ4oimPvBg9bL5R+LoT8
aa2NhF3s68auRG9Tkm09zt7c7uDOHk39iHuQP+otoSZwQPIzcPG/F2DUpM/i0seC
gxCRIFqCKOm5HtKklFH0EPyYAnCcz7OAjIfNatbKSEq5k/55Xjlx/r2BUqyTqlTD
8azociiIvZsFCyNIt765rtH01ueS+pETYXYM0VQmHuLootUZ6xrAzyw1+nZYNBl3
mIhnqYVmz0X8rkWPd+eY0fgoWiB7xoQUzteOjgOGgpYGglkmd5PC+VWgossGpghm
p5C6pfG0H4DAzn//69eMNGu7ND4kD01gLOzt2zm1qSrcUD55kS8xIdevJs6QBqSM
VT9CMBW+POsayVGnck2NhXip3wxFeoBcvTRGOQkb3YZM7ZWlIAj5ZHiqunvL91m3
/bxE1CDX8OamaOgKLHLx9KrosWcQEUDh5cGbz93SGCZg//piUFDhv0ZJ78H2CKhD
vbzZyMf2VBq+7614Pd+79Yjs4Qn+vedKJHQe/pr0lg+g9Sgh7CjJTjnL0uw1l9yZ
yAqOwMDjzMSHiq5DTwfvQ/O+nppAAHu+CUMX54yOhC2BUEv7gcjdfukkVWKY1FJQ
zLuiWsaoTyAQ1QE8SUS20grGAn51gQqOcicU0TjYH6xjn9CmIqgXgMMTvA1v5NcZ
p4P9Rpy4hwb5K6NuLDbzLXRgvMfDDPqnxvQcCaxGGLCyP8Y6P0UZ10Msf4Tb7cvB
Q9OpCwXb5OqFyl5GsnJnnyDFw9nO2p5RWh30W37eIbQgAJmjk4OQlLmNL60oUL6v
BsrjmeOQzvgnz17rKhz+TUOjNP9LRoLQTnYNrKBHbK1LXCnTB6+0mfaoDfaJOlcn
2LL9O451Xxg9Jdadj6/spoQaC9mGnTsCRWAK/L0UFYiGP2snLJre4W3D+b2eJgKH
Vh8SB0wtyzxPsGsEiaI0yadkyC6MnqNfN/Gnb1dCaXkMb/7paT12eAMgHrqw/MrK
6vEmZExnE0HNOYKl3mAb4ep+m8Zlohr0ckovkL4A21i6q6Zu1yh7tpdDsbh9p2i/
fZYpvSNBjlK+F0RbBhqOKzbNC2lphtOxLro6UG5RSohEH3th5MZQYWeih3CQhG+k
SlLrQmi4uelqCdVUmOpI/d14hRYeuTxryN4K/i2xic1+N6jMAg3FA8R1BH7d+WV4
uQH4DK45CLI5RlUrABzpsEj1pqJVPaAdJC+AAaxvmcM6c4eiAtLsxlV/OUyuYaXD
y0X1Kc3rn/3LQFF3Rl1cvxT/KQR11Hk+MQEsekPGRRnmWHAk+H9VDO5z83PH7BSX
ffAVaiQGIcRx6cJ7WvX8UQircSfLn4Y4vHj1NeyJr5USN5FUUA5DK9Hj2LSTwLrI
aLwoPFBv72r1xK3nhp9H6LdjIWmBBsw+YTWHWvR1j5PT78szPgSa5OXDTRN0b6bg
iwPJAtSJ7+k7fpVBoYi7kvcOqmguUVjk3PeXlYOZwUnxWmhqwlOXTrH96mI2jFCm
DlLGPKrU7YzkplWYkDGh0/suVJtsL125w1WnCBbYmVfQD9Nh1il5W1pUmGF30CAS
oychnMvLgy5YeehaRYoyi3gP/0ZhTMmpwL0ZG8n1X89dQYB6YzBOpdoC2ssVjynY
vUuMjv0o6KI/foeBc0sJgceUxWU13TpM37SEf2CrJWp5I2LEDf0iMh8L+MOTsk8q
RzLbhRqQaisUWOwl5Vuu9f6mUrCNXhBGofaO5EVGi34al8NenfTU0wfUNYsiYDSL
mPy7w0Kpd66GQUgFVCvrIYqI3c0czqe0HdLE91cw6DSr9aLiZsPyagiJttdhsUGM
hlRolCORRgmlX3xTupTIkdKYt3x3qpH2bpzN8CYTbhTSC0idi2pyGyLkMwNDIe81
zidKnZL6PgyKcXTXNuvJdxlS4tkRe9vdef5/Kgrm9Befe1fC3NerAroeqRJNnZXw
STs4zgix+/mIOUaS/TZ2kzjip2yaZRS2miWiBcg5Zm/RnZmfW0r37KQmA74oWWZW
kXZgEbSc/fENjlgHTBlMhW1GuWqxoihBxLcjtvgefBiWxvOzlUqFew/C8y2Qb6bB
LBWhl+xhbM+Vn68d5a5nwuKYl5IQZ0/3J6Ur8fL5aKTxhLv9Fph/5ytAOV6Wkubp
RTBkv9QH+1JiX41u4KeXnPvV1spWIvpjt/968M9sZ8+r47lH72CiK6qrVyXFWHi9
eDy55CurC8EOrzGdRtvNg6VcVXQ/rRlK6I00HQNLcm08X4j6+3Ssv83AUzkR+8a8
nvVYueOSMGpDsyGwKh+FXclz/5GYNR2ErzRa90RnPLkZpkNMw2oun6g3mKFmYny+
5j+1k8vsvSdkSxQJL1st2GdQnDIB1t82pnLcQd/abfeuRkOyaCR45y/nZuUruQp1
K7Rj+P38kfI1SXsgNmc8eSwSmTrhEFhpujvzJ7hIcuFhF+i3zUs/inG5Sxf1h4tF
Yy+McHxFA5knPkZCSvA+H2OSmUf+OhKSG3PUKX+zrlCo2/woDL/osj9ze/lFyhrj
norj9+0SlYNdiIQC898U4bekYAvCOW6PNq/5gdag/5tYJ1gb2lHmPs5lXTAKFcgE
3IMoLAUsx4dvexqHHEqBPbIo8au2ITRYP0SeVXmMr5KfmzUmDi33m9lppnlLb86P
DCHlm/v5dN6ff13dqUx8GKqzEWdHQLsey29P+yAU8AF8sMHX2eDvXYxHAxVk5LUN
byFhIRaaxmgus7+PwOtZ7cfcaBHUsBbpkeojabV85Pv4wM20/bEsfyCVNIIgNma5
yLQXuJa4NI/7vO25DP+ZchXFlq+CwBCqjVkXzZu+afdXhAS73R8vhW15pwtV4VKq
1evMZFgtO4MpDehZlOXihN/eWlRtFiCixMUkDJFrbYmTEapkclbT73bBiUtY2/QN
VcNIMNiBTpgYRtOhCaaS0F4JdkgCBm2RhEc7RAASWi1N/qXmQqn6TkN+tNPXFnmR
BCrR6ZhxQD3j9sLo+S3PFXy8/7sfP/C5BzmJ3zjIe0NvBzwfKYHMrsZZlLLz0ZwI
SJUcEOp1OHbJNK7JCT+WYvvwF8fGaDja1vQHvBM4aEX+FcE9pVl5SWYl5LbJkXCv
VOQtDk/6ewIla02lrLOMArJ0PKHXSYk38IuDMiV/xj0Ry22lnMIXvDPp2pUcGB5k
Bc3nVpg0AbjluVsqJScuU2DMZWYTUYweKYcU5/xzovzvbmvX6lauzD1r+U+IiNh/
Xalx6i2mqbs8sDU0ZKXtrUg0iezaE2UDScl9cd0iRz33fEA+iNiyabDEqADUm9r5
VL5jspGmp040iXxYVCV+Yl4NvJWzbBMvEogLd/g55CBlKCSGBq0dj2h2i6MYOjdf
E7az6T+1ak+glu7CCjFaMxI11vOi24I4WDnGDi/BKTCtZz3hTc0rzQuEfFOr0FDY
ptzvGcpV0EuAwRnKBE8K7D5u+zudk8N6Sn7lbv4U6IQGUySc6GhVlWaj2Lha4kE/
0j+i50PAf7plNpDJS5stESgZGWm52ArtqPeizb9VYRJCRNNAa7/wtBA+aykawMNr
nxibVnED6zf3VSitThsns9creJRUkoutUKE/Mve0zyQuNE3OFH1lxEc0KAy2HQF+
0FLSU5cpaLPXCPWq1S5sZzMk/qpa/85eEzd1Y8B0RPNTL88E1HcWpBFtJodjcugQ
FESOe7MjeUA/mKYKx13nESi/Vudv8Q78adP8aru1JRef11NZHKSgs9OMjwtT6XOe
Zl2QL2ZO3a248HQ6hQPQQXRMO0zyDytvgwcyDwkN2ai9thDUTpu5pratCGTqBfWm
FOnCT+g/Pf3huYD5rZ3lQMc44YOKBUmsXPQjT2flKIi8hkdSFLagMRySQ433+cV8
YBoOV/TY4zhREmQlGCugY3JVd9KgR9nUH4B7pOw/GnWRs8e70zJYtzziF8f+rnTq
Epi67Os32wRZt5tCyp6yjk4bzG/fuLHyOW/tKDjflOS4f/bzwLQLgL7d1gm2uMSO
YcgFL8/xaoiBubpNqKWRYycA0cq69qik4x25Jo5oTiVu7MryUcth/E2qikvbNOTg
jQzmCbBDzGMKUDGaakcRp+HJ6A5PQ8yRBULYtGg6QPtMU42lbKnItFqeVBUUUnA1
UDJkks+icO8TDKAQ437dW7Sc2VoOuZfHLpoBB2GHi6B7aUG8vCJ096xjukCUR4PW
G/6ILtqXBiMFJEKhnTPBSUEbxv2GziM102K7LcUINOlH5EoO98X22oZD/i8vXmyL
XNHjW9gDZSJquqyjHBC8TIhuyjqs2o93Q3gtg/wavm4XkrFOTYOxJa9NFIhhQm+/
1dDB1/iqD+BJ+/QaWhoToRu+eIA9XwsTuFwFQrJnI8nZ4REN9h8LHd6FV931Podj
WDPIAbVHVqi+bGusZFMy3HY4aoL5+EKs/9dWM56kuE2+aZx6MwNif+agforZUWyz
ANhiptyqAzNP8eiIMZKkFWoA+7ytveV00/0kCBAjWUaM5EMF0R9qhVTxPLi2tuFg
+M5FNy0rFPKd+jX6q9/HxMPxybDNGZCBmc096dxqd+2YfFfe7Qx+WFJbx81TRgUL
hAWRbCi+TmJemHsg1wkT2OT0jkxu+3eFyeUeDmc3dauVRGeOTbLnGdzZfUs+yrsN
uCpddIUdtziOCJ5LgJbTqy9qE4eWnUL4vHDsxvpR0dxSXT0RqeLigs8hn7Y+aswy
aWLkl+Se9J4BE6ajCYBlahGZmcYgh0laK3+/ziJEIrlI7n9dBEgAbPKnBZ62Dr2h
WTz9k0kjgW9GlJ92SgdUrVchFvPewVFtCEvqFz0FRTorPPVvdB7fuoPPrMGlYkzD
tvQ33aYEQcPanGBSQxgzXEFiXbGx8kf+BWYtkMnD7zWau1270kvBLHR2z8rGp146
1IWzlHEAVFwjLKvRhaixJe+/vg5quczBpVxOHNOzMmcXWI0hW0X4wXp/SmJYMxCp
9vD1T2JSNHeQik0+ynIuzR8PIPnfmBGuZy9xNuCBPGup+9jlSWSrpbnR2vo37wVD
WqT+2xdEoZpuGOksT70Jgm8QRJjkF4GxH3iI+PrH/Zd3nUpWIZuNaBPm28QR5BzT
4OhgCLg1LSaZ+Rq/lo0wcbeJNfAvSRQTJ4Ja2RjdlZdtCmmKFhlEKeabqZg39Wi+
1FVEfBWihyggLlpfFtIMcFkx0hToU90Z0ib1wkxcCTPjEd/YBNuRPGuTjVOP/dwu
ytLFv5vDFAWgO2pBKLHz+Y8vY8osYjy3B29+eI/d+lQG8c0OXdkRJ/HZ7i6s7KIe
6lRQEw2Q/0+bgTHmhF2TMQVe8SXt5XgZm/sqfON3WuZGPEOubvADShz4X5SuqHsN
FNiy9FYOs7ElYmWSBBwZlgmGJkYphR5dYFbfRKXMubIVtaecJi++hFx07TiO9mbh
zjm2n1PAvfafC/LYGFA5G7VHZ6og95shadiE+AURlF0MYQa83CWraIwpYQeVqDH5
0HEDpt63HxZ7LfvL2JMPu/3plKbCSz2OVXT50NamPQatDQ/VGWKG9DihJoKnoOLU
YpWi02HAF+qc1OUwqzvPeirH+TgaGiuWDvv2dFKKuJiJFp1lsjExC0/UAESStQh3
teBQ26m/Q7ljN77apV5MKzWWzZUZIWX6m/wFAujJwWm1aZmsCxgZGqp0Tswobeqq
jzGAKheOn/o8H/3bYVZUDiEUcq5YpVs2vxuNbS90TGVjNJ8mJbfqH7HbX1l9hCQo
R8THHnHQvfBU6kIWnjK1om2oEs+xJOSigM+KSzKgxhXOHtb6fzTadAucrpba9xny
n7VCfZ+aZbfa3QfxlV146sz14S8bNu/uGmHgUibe6R06OUrz2rDk2aOA4yktcgfW
LdWQ4ztoD1yaQzwMixzxV/uZqY/hFs3VjYRj88pf7D6jN/mCq03oTyNND4SN/UPX
yR6XAbmm/WFIty78LKPgEJf3p7ga+URToUro5VNoiQaW2O/0Kqc5PpQVh6Q6SEFl
gXpIjhP3mXKYZItV7LGIBp4Zcnqj85ZSfOHz2eIDCFUIvDyGpDlERiBSI+QJ6ZNg
+K2g+05qAGyLq7VTbxFShmLs7ZKOc9YVGPFbzKP62fc1B7jzsBwvJwG0JNY63tdl
WKK8MXxifpJldUIH0rfQS78rc/kN4UOAZNE1vvMtrXf/4fHjb5vl2BLHHbNMzraW
vKMwKww3aK1OVSz65pLlz1fDEU8VAofRpCb1tl7JjaLB+xAVxsQIxj4GXJIXMLek
XF9OOm5gsgMwTNHI7H1mS+z1T255Jdu88mNTrAPPWlqlr9YVU+k6o+msfxRV2Sse
ei9bL/VWEqIGLSD1BjZNiyFSwwphi0MMIByLbbSr93OHJXDMUCyGiCIdN4Q53gYU
/Jqu1eq3EMMcodzmr6tRKGNvwZQIWhao9N6hEPn40zhaCltPVEwj4p/y0jyrIn63
ldBLESIYp/eRI5ZCPIy4AW4shu6rO8KWJK1W0wN4du/oFCASDx6sPGxQ0hiZtoNL
D/WbKn+Fo2I4HdZreJsk8P1ej9KnwbBwiHMVlPh+yqRa03n+GnjcW12Pmq36BhmF
tyvaIXBZQLnr9aeFr2cXCQhMYV2kmG/rzBo/TwS01H2S2rIYEp2z6g0mGhBN9TVy
ZcWOL8dbmLtjbz7PT4JATyU45H3dJw3+bOhTBo7K9QHywF80NjRKgPZmYABPjPRT
hqBxYkEn99ftpfNj8C5RsO7Oeh6vV+TZMM4Txd5GsVmicR5/nlm5+aY/bXsTIoWD
VOIiqXbF4+wJXOh2jNvAm1C4j8yN31AUzaJl18urr+HVYYhaw+2llpofsGBwsfJh
KS01hoPLYASRJUQNY1Dayf3xEy0oS3hM24F21ktF+n51AWT5n/NvhhQdGm4D8I5k
r3L+rZbpYOEalraOGjzXod16eNWDPdZIu/FbHBTJEXMqsYdmBd+UTkluJGgCIVgj
l7Dd9i1H7Vwf6fRZUOmxdC8uvzs2AMXtUbZYgCORj/JyyPuuhEueTM1y7l0KWfZN
6P5RAFpRGtv5fmLu5j5zzsx/D/j0kmK5Slr0N0ucJYmEaXyx2smDjRCSG8Ef6AaV
gZ8Uu1vWITtUdpPL5R1zV0oT49XbiiAXUW4abbFLfzdUPp92lbQRwhHU64iK3Y2x
L2oCkSsfIdOdLd7S0m0pAz5+LJLo6zFj5ivREcNR6GcDMwodq194UuHk3Tg6YlIO
qcCclJ6obkHgNIFoDZl5+7hPEWYiOGzorwVpa7g5eZirm9nyZ6wUi3usStVpbafb
HJCueIk3RgmGzcrzs0UGDRNGC8Lh7ADAmOUCkgsk5ifwTYKPDTPJuN7sSmBqpqw9
nNBOBlBg+fUp/SWzoHpQPAtUHGdPfRiRdftdqFn7xnzjpAhVI65nWPZhtLKH9cD3
N+UhQJWypQLjXZghho7Goe2Z1Hqd+ZaZt6N1GV0OdIJRzq36Gk0mjGlLESet/NB3
ciy8Yt+bcMOtztEVGwVfXYAlRuCSUkGt3GvJYJDcjmlxVto8MH0qjoKKptxaf9Sm
L/k3w1qp6iwhooQ+U0cGJDnEAsXfY20jOrw46DT6t0Z7XlwOwYuqwT7P7q8t8+fl
2jCivShxL+OkXLGVpafZXvpd7r97yhmbs2LuEbvyeSbI83xN4841B8r9jj8spwQr
FpfKVwqH+6FOa3+MCuYqNcovxYBXqjq+42VoAQOpjPElH1VEAHxfRjrwobeRgKQi
Lj0TBs4fJ7FIxjfqFn0c64YdEFpcVg3tv8kb/5KhfmftcfSCWHUPMi6jK3M+eGcP
zqPNlKywkALLD9cAZMnb2lHw13fk4yB8e96f8FGp4KH5cdnlp6rj3KkPeU0rHMp0
UzHJl/UvyTpydr9wLiYr0LseLECYaliWnPB2KR6EJ4Oke/s69xZpo+xDesUOQtCQ
RgSGKirMaH09YH3Tazpc06qsT9HvQM13ob0SOllcxeaBlTpz8ZvAqWOd6PhWehFq
v+yqfeIDN/qQWfNqi8EuGlezruL+hj9xQ1oi2CnOZnBcECCJCgiKQxM7xU+3N2xl
l+dvcphoMPhQ6+ptNBElxIJPnu7NCTBB0dgu9pe0lE6mvjh/9p1Ytweb1Jkwegwr
otr6UD2YfVSb0ZUYfNipm+hBvPcdZf3GejswTQPNGonxCJMvoeeVHz6jMo4h3w8w
2tsnGi5btxQIzV+m/CQgfV3/5MJ4HESodnKKrBngKSvKeIwUQ7/LUpIEX5uC0KJM
vcaY7zB0WbwUcUyyOinmFFzthVa8YpKXapQTOk3l4hPG7y90iuxZb5jnm6S+uijK
NXz0nMZGxmpQpZuUNb1M44kHxCd5wwb6JDrbeO+aVsSZycvLAoCYXguXZ8RE5ARQ
cbsqiFSRzYrDBk5KAfwD6XVAOcNaCYNJ8CC2uLK2H/EZ5cQuS3cFMm3wB0rP3emI
W+bbpgRaegJADW1Y5NB0bnpmwyv5iAc03WPzAqRhLKAxGzdj8M10v1XDjLtZjKe3
UlN+Fnjexmra/WEYT7LBZnxP+UE7Rk6BYb3Qr+8i3TDCBla647Fx/SZSwSvGZmOl
lGFO871s6cOFNhBQbVzL9zaC1LUkOi02/Gt9WJWKotH3sN5cfJxE2RpfMNs/SL+B
33cGmgiIuyubVCgTl3tg/iybOgSSN1M1hy6qTW2Io2v/hBWeT6NJLdKpheODmMKE
64BBOvtBtifTZt1McNqOcuBC6MK9RIT43DJE/OqqMq+E/eHUmH/QLctNYAwdbMaT
ACLoJvP+BP2mvWjWQkB98OzQZUpJMrtI7EN6JdQk5oei6DX7DD2W9Xi8bTZ4DTvt
dDw97sW5JUt78kAIQvwsCOP5wIzX5/i3p3C6NXwSntQMALvkMXIP8ACRGt50z1+a
4YLgLIXkm/Mw7QqyfhFI+QUdcA5d4sHqtWm3acgsp2L7qFA22XkjGa8t/TyLlnPV
rz1IaNpgsoQW/wPpZGecUfR0FLzWRRokxEMiA8KQRiD6LhN6PEYCdRkNo1Zzd1Q6
RhGS2QTZJX0TAnHfNw2nSwMJbTUyuE1X2QGEbz+x0EZSWHodnMRoXtc22abc8alw
P06tQ7ymIXltsGdKDMg0J4aqq1bByoJjlQo1pX0/F+SJ8uyz4ZhGuDS9/l+oXseF
O7fHY9fsp7M/fjLB0mDky8YSaLxCLP/gwhbvQ/LhTQtdaOOk69HVSKSno5zwxiIb
7zJZ+zqBmSsVhk6Bv6ehi+rncMU4KWY/RV7wR77ElbZFgOR5no7U4bo3lcPZFMrk
vyrKiLvfd1Wfbu+j1nUJPGaI6VmReDg2glzqsZ6sU6UWt+3ApWd+fpJa0uackEyj
LzDXfrHyes0tqF82MepG+Upj6obZ8I9zcvde8cIRBYR3FqJa02LhwLXLeUGp8qHI
93KWVU9kuY6FC+fPhXI9gK2oEz4262hGl5yLoVK1Qkh8TfBHJi7YH6jUC7QAaQ+p
oySeTalmUk2Hry20wJ8jZhAjTfU9z1KAUYerbvXsWFzUl4gEiaqZM/euVfBFU7z7
xytqwuQ7xfS17slBQWbHNsD2PdzdBVp9nmbfd8OEc33DdeGMj1P2mZu9oE/l8PXZ
D/mdgCl6l97BLKfWQFO7FKiyNkamq0k1QoL9savFC9YK+h2MHCW3lOqITCYjU+Nk
M8mbxGq1x1nUBtsdlufaGmNwNlNRmIuHqemr2fIYwEga2L68+7Uo8xjnBfEmGyHg
MBw903Or4UhFQYW86yDlH04Ul+cDK29Gu3scEI3Jpl42dz9AxzhveIB/hqRr4ZNu
xVfVCY0SvoDkljMZlGjOnLv9i12nLiHpAt32WUTnroIWKMHTzE5Cl3MUZl/o9oaH
W8ZeRX10OonaakAEqf6pU++PNv9AIW6kDHcnDWjhR2s3ryZVPKQBlYsy63mneiop
xiUxcuRIhtSCp3v51Nta7CbWrwL7n2u81VgmvtYf+mgRK+A1XicChPYqVCTcL2qv
evBfqZxNjMnLddqszWmSmqB2p/7re2iEYWKnWYaiJDoJ0ffzrVc4rgpdaQ1BvDTv
I6WvvczIGEoqOeAkxl6MKeWSivGI1wehkAi/Iz44bLWdOLqAIZvkNLtnUO/iypih
BHM9VFD6E9fAXSGKth1lcqhNhLUINoQ4WxiKdFDO2dr9dKjDgKv3kO3inPKWj1v6
ibmaiSd91HOUmqEmpeGZAztvaKGiWjf1UqSwXfZTWeTFi3gA4RA+3u8jks6DHEcH
wHMoz6jioJBCmAB5oGbb0HGfh1zpaLDv5Kt2Op3OTFiVHsIEnN9t/XpnBjI/cx+Q
uK/8FUUjoFnl1XKmRZEeU/LQxgHsWTncCMC6N/+uj4NAgz9PmycBgd1NzT8dDUvi
tVzI9zwM7wbbrFvAZsxiIDp4vPLuHFUWCREYPfiacwXzf+y6Lsev3uiJ0Mwzb2or
8nSsa19MoXkZRGzOYCYbrRkrGh90/IeQSZrGcrknxYIkylf5HVaRoWG7KnkwSbAN
6YvEr3ExRZ3KvIsxvBCWmFF9WAuzFPmLZnmxFIxnNzYfdq43ezWMFo/RhGZv5iXv
Krudg6JYT6RkG12BrbGtiEN+BWRS41ybY7zB26w33Wmck/BkQ9Nvrt5fsrW2Yv6V
p1kZNAJtAMc3UQX+LdnDizfLLqMb9yN3yWJN+MUSUSgFtWflMwx6et2BIErxKAGa
Vkyud7QkX9LQjK57MZ9QIWwJRBvWpQ2LVlrwtKDWGITyWQRHfm1er671bRelkYWR
NJ3Xy/WuPbkU6tQfCGrHTI6oBSHAShe8AwBGFoKtVkQmgWSb/ay09tW+wrlKcotn
d87dq78yhZRDXzzrK9oHwcU0Lrn1wHNeAPbhOhQlGEgqVjJVNkhwdZjreqiRIIVP
e4Sc97RKfX5LBOqvRCcjKN9h2Y8uotKgdtHL956bMwIuaSh59JxphO5aufbXttjs
8Sq9hb6TJYLxR9rlN/6BeN6p9Q5lP8AVArqh88/aeb5hu3Ms17QhcV9BISnt13Zj
31gwAWsFGUSgTtowSKcy4/cQtAv37IuN5KFA5yfWYVqTwBLbZ9I0ddEJAtCTZs5Z
PJZH06scSTGm2ydZNnWxdjVoBYPYYYS/+zUN70PIiNSt8QgMOd5FkR3s4j11rqpl
old4pxCEOXQ/8wf1uGIG+kDUQgv6cc54x3dMYLAA0+GZnd9sjaVnH9PGFqbK8r9q
6y2TUu5FswB+XjDsSy2jEooOQ78bS82j1jubm5mUGiMGaTdjtWkgxsTsbV504a4L
MTH2I7YEz8TvpOoK21Mt0LIlynDnshd8xWEwC/sg52lPTEPidPJdXBz5aa0nZwFX
gPPdeAFN2AxyiVJk+tLPiHrgFFIB4giw5J2cdppFC4K35E6BSg+ejErKrumPaDSX
kGmF3NWliiGduyri4m1KlTx+4RzZCdnmjDuWpqO/MpBfaXOriZQCZ2740eEnUrvG
AxxaQkWW0IXkzFZDwlv+LOMi0eHh4wSkcoO1ulcZh4B7016we4Pg1R1w//NH9txg
0z3G7TMjJgAPMcYRDez8drpSBtwS2GsORb7XvGd5F70vOd6O3Z6DQItykcOoccKm
0afkfkWCx+ULHwLl0PL+aZafYTwOIng/JP24WwW/xCpPYZyFxlpHXl3OLCGw+bsp
oNiW1cejI8y8tlwuVCSpfs8OtuUftFSLhIx3toqVOCyr/O62Lx3DASm/2+AbKdZt
ByKo9i2iT4W3AXDHRJDkZvM8p14/aP8qlJnC5JiuE26GY7Pp715Ai8baOM//TEG9
PdQ2/hj+77OfqlFdKJ6s3jpv+fl/m7L/VqQri5gYURxSLl/jg09OEn718zy6yNob
K/x4l7zrIlQt2nqWvdyJxklQ2Ko0aW16jfCq3SuHYo8hEaurQRDPXsmKSRE7kieD
kbo+M5tghxgodvP4hOZVHhfhvgGAN56uvo2+dfd+lYI4xZvywrICLH9F0rXZDZsr
aGeFCtgOfREYJUjf/W5hKhQNLbWhOJ7BhNRMEkoC4W7AxX2wCrDkUiSCvpeZ3jzS
DCen2A4bC7m3E5DQb1ZsMZevgAGHXEQBiQHujkoe6yE86jUVlCDLaaYrOU7pqORE
7tqHcxYyeFbI/EkhwPtk8+UgZWFXHE5RfCjaZ5vzu638MfzKkFz1wJ1HJ1+updNH
0HDpEV9fyw0FQzIiTzHUbTgKZeB6oGUQ3zgB6BZt7VOnZj7XRLsV5boixlQpuXUb
IPop3dVsmAlgpQKq/s5hvRC7vBtwKZqg+5ZPZ23knN5nwo0/Yw7cTTmWkU/qmPff
Li8bLkyLOmwSsdZpRxqgkQ2Kw+TlzptpUikoS9vN2jpUkBfYmUTlNfAilyJ4pIDw
GV2GP+ySbOv9TICT5YozYuEch8TDuCCzJjNYxx1dLP7BQcpxJO+LjIjLYDpkno36
IVJj1rTizr2J3+Y/zWecfARCtAdwaz2PZesdcaHdsZoTzOMo8eelRQD14ANH2KsX
i/8FQYlMVYyI3ymovad1NrufYEY/mh7nUIerI1Zar7coyz+6GHBDjsREHyJlZhLJ
aViGmHbcAFPizocABvlVeZex1Aq1JQiGXeb3sUhiWAgwp9QrbLYgC+0Wy7KpsoSB
pRYDWeDLsxwn8ouCDPc5UFrM4mmOwisF8MXbd5fAkE2jgpZeoE1qx/bvUphRYVWl
6X4G69jJGDa6SgciOrSatBZzcDpKeZ1sWT8clmwf3xe8S/C+2s3YDfBbNDv49gZ2
wCq+Tp+uNTLZmPDrAWrdDsGDBNeswwSVHeb67VHz0GOk1LlQkGu4S+H6jPQTiU7H
+68ZuTBX/ydmR9huRa3p7ktkok4txlDs0pAdWflv0D1s8kUSC34zDL9vc9T2qaYC
PCJMrBeJ1wVtogDbpnYF5Y8Y4jPfHQ7mrmWP/W9+4TfJe8qSQjT9ur/ZfzuWntu1
Gfw81wvcagb5d6hASamNqqlohj9FAjY6iC0XMahCk03S0vr5VuDjgoOKyUO2AqYh
5eHY/GqQXWfYrN5r1yZYZSeRPZnlp8by2N+2ZeaW3cEkP74HKaG9RxiB+BhSUT3E
W6uHL08ufT7HA2+gC8CZJifleR1l+noGEnGOSFyy675BMeYE9Yg2YUaq1YnhIxlN
aW3HN4REG2k0ErQFoSjKmKIJ9vxt1FiGbrd2thCq0uRKOYktJLETKXXD13uk9e1k
Q7sQJ5aaDIRVMcl/obPBUmcqJOSdhigPa7XITLuS61e2X0xZzVhiYkwu4QgsZaqJ
8SosQcMq/nTKj43VYyBNZROWt5wB3ZLc7t9DOkS3Hp5rRvfGuxiZ8oHcp2n2Nljo
htF/KOmsxCGCUqqzY5bh3b/nToEMBsAm2GWf7PBsi7ovM9GszcUxNq2DUWwJnlad
DLbJ1VO4e+TK+wodhAcpSFCfjL6WbGv819I0l+ZDHZf0NOYMpkAcQTGZRB5jwxwL
CVWOhfoE4Ggqpuxl3cEUJmktK5iyvFULFwZqLeX/I9d2aDVQ2We3ZxNLWqaUQ7cX
kfUnfAp4jMQq4fBQ62kBfB4X+FbKrMIgFYw7PHg/t1Y/uwJneLtPU4zU0hAYm6Zl
032ewv/6fwGt1wsVp1Xdtf9XOdRbj8zw40KCmnnPtZ9YKhAb8bqMZN57ClmFGhIQ
nZdL0dI7he6uh1uewuG/mOeDyjRcxAf9QN6RNzujrgs5qxA/j1U5q7LW/ou8y2HG
12ciklpnd2Pq6KZsBSEmbpRJHsx1Hy6BBibN3z3gctSRgFYv0FFBw/mDDI3KP/vp
us96U5vEKzFoRTrHY2ksxm6e/jHld+R3plRK54vFmnZErynex0x8Fl10elwjLRAC
NewbN4jrt8vfWZa6DHjQqR5gxLFWUHcVU4gerFmsTY7qhLcvnBGOHcalJ84IJ/BA
g1SmM2J/zd4qKyi10q74wj1eYObSKO75uj6VPov3I7ZO1NB8AATBg5tD6amRcd1H
QWOqw+ce4vvS2Q6DDr3PGoMjvH0i++94H1CTSkvU+G+P60HdNX5ZmkL00aKLGF5t
mKA7ZO/B9clFu2PMW+bPqpDlMjBauDZAozTmr4cJXbhv+YjScXCfZi2UFC1XlaAb
NkOdVD7DqqzHhKZlVo+TexJVmSJUGg4u77/PdPZDQBq/hTn61fZLh3VirNEtlSY/
58xs/vodLVPsLthsqsTRBwiJ8dZErUn/x+SRIkDNIyyyPWxZnRJK86ajEUsW3Ebr
eu31sgwmiltGtSyO5BddW1XqD+AxqhqIamCKflGQhymyvb8FRTKweJY5r4s39B63
mhocm3v6mjeMCArbEz2vxLNgckwcdM7xsLPrfoiWTYf2YvzFZ4xlYDFz/iA4Fo77
9rtSBfaELvUo/PALt5YKUgKCS75+yAdLD+f4EHlqM6zQt4hU9ASjA2jkgRhUo6kO
NEDO9hXmP1cbbBCtBOLyfEfmjAVCHu03Y1rJzl63sgOG7TRIgR39BSpCuj9727Xl
EeDlGQVX0PlOuGOnifZYM5qH+WTvWBEMi+XhzHtXJKXXOe6W2gOw8oJjgAkvu8pQ
HloqsBNq4trC+TJ52kewbpwy1EkBDa5RiYNBpa4g29CQMRE5YkHknQNTKgvsAxPH
0MNoJl76wkk5e762CPZLvAK0oQLKq46ppIlVUOfpJp6Fr71jtWOBg8KkpKY6eXtr
rccWYzrJzQby81HtN03a5m7yAigvBfQveKxJxep1Iiwt7DrmxPkIpsNnmjVqXabV
vcJ1F1eztHgCT29ul1z6Emt7osruw/8HeiMetJP+hUEbZ1auqN7uKZaRyQjhMqc8
jp5APBxc90pb9E7cyAU1AvJq8A8vyHGW4/jyzQQj/HgklYY3eJEynXH3QMIya/wI
gR59WkGde2MAcW9fM/NphbB5nGG4wAGaW5scikvzBd1JgkujyuTcexHJ922FZi9n
C2jopm25pUdqeAxYqnTRw9JtgUAnvlYsTBZtG3nKZTq2DRTpiZ3MOeAJaDFVKKLz
unC4/ORfCHlHYm1KXTWE/yHTGB1PxUAHivxRimaVVqMmXW+o/k3ZMtLX3RdJ0qnH
6sNA9m6qBrL1zlosz24HwYOjTWI2lwv/RS2zY5YewgzY81hpHXKr08D3ZFkE18DW
asqENYOg4ae4KYkl12cQVDWYYvYIHTbMJTT/HhwDHeINdfQFDxdcuUqPDzBeDMVf
8oiyGojxeYxtiZ1GO3tswSETFEaaQ1wQfd5X9GZMgB1nCY2wFbs4UNqxsfaQc9gs
Zn1S1Haz9nSyclrxeR8lM4qoZGen8/bzxk1DETqoYiPDMPO6haNL0C//YJ3rjyla
BueZBOoEeP/MYFYV02Ax3JSW1VrNphq+3eP3PRYIyVtRyp5tBESX9RwHnnF8IDLH
9MqdPq44170uTyzL2Z6/hEUooq+WQ8IEG2eBIccndCyQ6QyM/gJUbp11p/d9eKt3
nzLFtGOPhq8Nf6pu7ymPZfBQbHNgQqmFlz7jcmhyV7xLnNNEuj5xF28qV4rUmck7
3Q/ZPWmaU6yX+LnIJR3SQUlnFb88ZSRIqzMw3PSW1GsHTiiQnIymc4aodftsE9o0
+CD0RByejx9VAwtKvRX2W8mD4Y/s5y2TpTKuNZEylQs4tnZ+7CFMM6acZQubyYbu
cUrgs9MH5YyxR1ScbjFO9g6nlITJWOKYjY1Lkm1Eg0aYW2cDtA9CH0MPRNJ/4d2W
jBEVdUQo1kl1cST2Qzpe1FIQMcEdx2ZVMkHWtZy+GkO1BlJjKWaxR46uBfxhun0A
A5Ehcxu/ED6TIBJmIwHS5we9tH1dYFUXm+3ULHUsgETHYnoasxBsXjtfmd5J/kod
QzPYb3zvEpfMJ0LwRhdaG/mT7U3PZa9hYx8lQFnJNvydKwXQ9CvObMKNKsdCWPSH
2uvIWBffeySYT5e06CdcWw8PbmplpZ/EAA6IKIiCLZls3S5ynzL+nkSnVNnybV0Y
p3Z5Adxcj2hdN09q5H2KFQPBkOx4u8mGcCfZergEfJj1nO0KZ8/W90nrKqXVWFBs
XUf/mq5CcfHXIsguU4brvAplupjMnKoo8yH7+CrECZyS9i9k4q6swe7eAJnmqbgq
sSf0fBo62grjJSsOR5YZyDp8ZmPc+8TtMGOtQ93YBfYu8fsyT78wKKgeOyAWsu4Y
VIHPdR1tDflj+PFekB8JyojVsOwA1emorBCiGaJcpUKLLwqpjGv3+8bjWE9hL0UH
G79zR9iAs2Az2we2F0qdq+fbLePAhvSl6tUPdqsIYt06VVerY8KYZJmtbpHxJ2yJ
CYJnc7aLs1ZP6GwT00eXWToqGk1HHw9CehjT3dlG2BcWEmjzJdYP0fUSmdohQ4gt
X6dyQewZUIDW1PeQiTZ/aAJ+e3+NICWIYYIdiesvxQnWVL/5dm/QYk/xPu7Mask5
u4R8Sl7P0evYk0Ka317FSYlwxB+BjMlrSEiie7uoMMnsZrzJOtsposLYB10iyt0L
pB7Hk4Qm60N9IWMN7OCCaf7e/O2gOWFp++bGeVnhZmk460ZMQtLfnZDk+btakWNk
nM5VnDjZ7Sb+ovRYl/AubMKYW6AriPDsbyGYLilXOta/od27rhWa929+0Jfdi8cE
YEtj9lAKAXZ9/83w7l17PkBP2nEv3cno28inONBEdiANZYnjUIwMg5oEcZOqYXPv
1WTkgpOzlBBcILZetS0/4x4ndDnN0bnznPUlZC5L1tltC7MnPMm1+1/dKTMoWH32
IbgQXO3FZTfTAQJbjqQwhED1qPzJn66zx8RliuL1v7ICMJM+mogabigc0PNTSl6A
WNaXHFyrTZEecoM9P1PuQyFxt35JvhcQuzCUAeCYsetVOybV1pLgLSIh6sCR6x/q
hPt4NNapRptM3WjqJX6s7kQn45qErYN7JDlQVg5qvLKKl3fSqnuffrW3Ii3SEuGk
9dzxHQyT1cL9WLCJ86TfIg3JFff2PtnT9ECRQPKHl32A4rwaq+uh9wD38cReY8tM
lrFztfCI5uElhotMbKtHBcMC+XvKpNl6BGK37vtt3zTaaSwb4Nm2WUCrdP1zW/g4
K0ctvSs5tBNBqxVqSXF2R637bVKw02ixZ2dNyV8GEQRcNLnyEu/ynwfcCvp0HwZy
UqDqNPy/CNUYYDRGwI6U1b8wDOtop2efmlkBbcTul7vn5IKoZpPJhLj67rkmXCQU
jhnMUyA4Tt98AzqiJLHbNq88zgjnZroIxoBk3Y2MJbtCWXMgaiAIov/1voDYQtbN
JC0qA8hoT/SRHkVLVzhB9UB11xeLeboi39RrPgo8P80Th5B8Sb+/obk4DD3nU20f
Qed5obCp4VNQaRl5N3vUUgTUirCgcn5oY4jvWtw6tQx7HGQsyfYpfPjtZvvrFD9r
Rc3gJEX4byP2sRdgGtELIiYud7e6p31HoCrrFiwWYyCLmRVAXmRpYM0O8T0GCKOT
z9yaIM1mIzgFn0EfG6EaVN3WJNguKsqDEWD8v+opWs2PSXC9i+tluObfqFkqKC2q
4SgGrfyAhHpbc2vcZylnckIJTzh5r85WwGaqmVr+55Uf4JelhIuieBIhD5BDcdH3
5CQNhCLUrhD7n12nhHx6LPqVefA5vK2sY2bSiiyZ6yV9yEMs9SvNzhD3EG906pht
bDmGvuT99yxmIk6z3TTan+LOAHvjSrRRDyOExrDifbUvm15oSmTOA+4zEerGyQ3x
GjY6Llr5HWsc4+U2QNFAiZ7oUUeTFjfmWcfLfOJ0AktDq2mo48xZF3oVmBuhzPky
DiGcsKjVtrwEbGQrpC+/DWw8DCNwQP4JjJlqzL/YI0PxaQCW+lQrszCCAt1C/v+e
3deXOyaR1f5NWDXLT+EnPU3VxzAgWcX2ppMdz7YjIfMVJCpA466Sq3+28NgC3ZMb
EV0hhjsQQSiJH7b2ahDym4fCD5FL8Z+TuzDc0pYktM5tKIqKYgYCP8heois7sUNj
3f6TxwLimLzBAsrzgp0aWbD60t8nW53LzMsBk5PlmtXecbR4uoVP2nOKP21UIrZA
i/C/dYf1cIlfQyiNfel/B/tlIWoQeYLWnqC9IvkOepbgCEFjcSu5DW7TM05cSG4U
pdVoL0V6Aj7TxCsFwO9a/Vtb524P6k+zmFzYAXvz/py1sq8nm1SPCsb5oEZjX6L2
UAWxAYeAp6ahFl4o9n0XhyVkYsIDvb/FWlvSys9f5ZVxGzUpcQlSi5W/1w5pR7jb
u/CiJV8gusuexiZBn+hcAKwnF6mj9VDHdtCFT9V4Q0ciB+Fm3hBabRQwKBw/V30z
k8cudc9HIHyfGPAotxw6mRAfY/8m1DXzmmSWeQ6fpC7WshRCE7md3vRGLSfc1fVr
+XJCB9S/t2C/ge26JXer/kKnS3dLqQdhwA48FsshS2NgNtX3VWL9ZZkxj+idcU3F
ojMHORFaHhyUsuONK93HYs+P/zlSjnGZRsokyGDEzRjvEzrbBXfr11BWgtJ5Mv6F
jrLmrZj03uupYE4TxosweqV4uDaVIcpWGKlJjq5uUSLkHNTlAYtwZKEXWRz/QUJh
Sq3QNC4v8XhevJATAhfuNrNAE/3WtBsgVoGlosrquhzaxe2qYfJ+Zt9nWZK0pOuh
PcQwKPxy7j4CnKMbQUb4GaC39LvDz4Wp8hcEONOR30Su07Anrn1+youL9uh83fta
OnfXps7ueZFLISzi2Ffygs3RraRXMcYTdMPUpSw4ur55cWA3m1yPugrhyuVzVTBe
X2rctrlVG0xk9D7gDkfcRHhNtMs6X93moYE77vMWozgiexeLd0mAC11aVaIKDJNZ
ZeQX5DvTDl1jmnv+ZCM/P4p0wV7rfSlfK7kR9/JKYsnrbpFZoqH2wnzUxWhcR46j
OugC+DJADWKBAhOFfIf/ap0VRbIlZtKEMRTFi8ERTnmPRe0SZhnPBoSiRS1m3C5/
De1UDVZdGKbJdjqc/oLEfNFArn770fiFwmePdByDYU1ZWhWlGVtdDwZOsQVnP2b0
pu5KANnnRYHcZ+waGakuHAn2TkPd/1Dkcw1mS8Sndpc0H8K0KkPm18oJB2VC6Z29
R3fmUB2iaRoRn4qs2DL8A6XEnU4xP/DfBCwkuf++ZvY7GUDxEtkUiyIFB9rORuOo
0oQjFbbcuiWFgd/Ib/1CyIoAhbNnUeB7A++xestrUChG4D8YfKhAK0QcOUO2rNqV
ApM1m5X0UyoChHox457GgRFupHnA0xn//TEX0rphDbw1uLG3BlSxLTLxUZfwGA4P
LiPDmetOON3HUbAiLy+ANKtdmJ5mhaYsCbNYs/OnTIFs48MfEUBjFosP5cgNdzfQ
fu9LQFlc4wKfqhvTT9AfQMkfB3HmN8eSrbCKqPwt9rO8SM1UM8XMF1qkA5voUMl9
Fy4Aniiea4pPpcquTuigtoHHjy39hmcbC5qch4/qGuRvcIO1Jz/Ma93wIXAiV5Mw
0KDbsZWtMmgEtfKw7hhePU5lmPrpDmlrlAIKsAgOea+DgA1HjEsnNEqmhOGH2TGI
mukE9wzL2woWlwNpgjXd6hBRoVvtxokamQ7qoIW55wlVTnRJrWJhpgAi/2T3COAE
rIBXs9vJ/i+FqWECvJuQytX/iL+kY/xh/byJm3XDz+fz8tRQImrsZsqMNr8Vab3H
1EgDcDGAiJpTwA4JYZBSKtCspCh/iAsVPfo9dwtUQ/ov+hJWYtSgbKwhZMKfSbw9
xScdhlaXJ28gDNHRGdZkr8ldsfb9nXGQvLAbiTHP8piCafEVY4M3HlXMZlpMjWoV
2QsMkyhFo6Mf0hzbV+rNgBywsTWEjHutbvSghoitLNtgDzh8QcwaJqenoB94zxjz
vaXXOYtqsHEVWrYJ9mRMFfpcmFNvTGGNjs8OdH3ljw3pZ1RmWO8bfJ21CkcbKAJY
11u/sRutlT6jzt1WVeTPZGoLAfnR0QJSjmopNZdnw1o8AquIDJ7Nhscv4FYMPNw1
ddApNi1CVgG2M0zFMSzdpGw5Kd1PrmAWk4lcFx/Z66zIC67dpby+1DPUTQuwbzAC
gap8J1ePMFgY3o84OpNFkarU9M0Sx0M/sSWuJdOpZR2M8YmMcuN/JuZr00vmiFbc
yfXJAKIoAnp9hr2WjDElTb7cxKJ5Roz5EAX476uslXfisEpF5N/xBpwZCCt5QOO6
87e8k4FUPNmuSN6cDv2m1HCs9J+L1O72RWCZqLQLo8pYxrQBJm5YaiEUQ1S8CKu+
76t3CHoIP2xJPjxsPgZHfxiFlADdPohjM4nZcGJQs84nK+aQOeDz44WyTXZRKU03
94BgAYCJcCJgMUjO/yqhyK9s2LURIs8Bj+4jCn1uRKuQKWwBHTXIuB+bJyYnvfo6
QwYJDU7ImX6kThTPCeeBP5vpR/H10GX7fT43JJZg+pOokLl0LlVcOX9myyYT6wxq
W3d2wP1wchStIoj9xKpu1VvgsBdKYFu5xLqaBJw7I0ZI7t5FevVKActVJDhAJNtt
6F8Kflh4N8AApS7IeQUx7wkjmOgvVIMRt2zTS3YClx3+XPlJf0KSohOz3qyDHYOu
PL10VbxhkDVNh84jCNjMHUv4F0ArB5MHa4cGt3VLn9lk1gxcvOR5eqfI2N52GpKR
b+2g6fzbxr8XKvarlcRLxMuhS9s7drokLRyczwEDi3rBqLuAVmNzsDjzYKQ3f5Fe
rBD0nH0x3r8cSIXe/LJMA85Ed6s1Zb2j/teAuDO0Y0HrmjB2uHvpVKKVwLRhNvBD
rv3dYgy8nPUbCizqqTaKBNPtR6xn8bFNYG2gryOuv/d1nBLMU77AAISfcpnPp1m3
PEgcuiTqzzZrWtCaZEP8mNrx+N28KcN+2w9wkD4AqEEJGmDmlvEXyOQYXLBDLQU2
ptpXbABzd2B7TWyzsjToyFpFfpze5kWXj0kxJA9I4nNm/dZrrQsFyHd06PhTxLli
KfOxfUJwL1UeYR9i+0yah/FZ/+c3rmj4AfOXyjI1JGvjKxdrmeHYuVBkToZzE2zN
+yWJ91hZ1kdip3XIuU1NHAnC4Ta5tjggxPMOhVIYF1jEvySq7jGVECPptniVa2Gj
zzxVhHhAohLqDFqS8LPUIbTuHFdIrE29Ur64ZN/+tyOqjnQ6XeEQqUqGVqv11FGs
uuYh0u9mIXNwe3rmCxlWK2htjB1+TYOUmyjTYHRPN3mI/KwxEl+JK+pB3gCnHTiY
EmAawWzs+HS8ycqs+yxVL7Sqyvsv8tKl33m2PkL90qspjrMMWIYcEr2DmY4Xp2aQ
to+E2Ciza0Bbz2StQEweQGZexh5z2FAoVsUmoHSb6HdS/62/dtjMY00EHflfz4Mp
e2Wps3QNpfJq15tL+lc7UVLykEyDijjYLln+erzXNB+jGqfSM1jsbooEtiG748og
nbUZGkdMGl/XMQpMmLWJ9cE3NzPXhjqfEQ8AzsA7QwlkW7dpIuy4rjtc5WMo7FYj
Un3ByrVwmnIVbVF4a9dzam5J0my0qFKy8XPsH0+eJpKUPqy828yS/396Gof+ZcWT
g1Fc0p8Z7/tXHWok+eH8dKqoYPxfnm9VhwKjhWVzmVdJtSSBJjTBdvpLv8rGYwRv
Rt38EOM+50Tv0VYOTG8vx5CsTNeD1y0iGf66q5cVkGNANkmCSdq646HhUO9GJ3lx
UpLmzyjLiRTw6pRNiiJBp83OzQfWcyMyuBckYt5ZzT13OcaRNDLPIxVreT4NYEYp
NI17QF2N5/LO7aDixhdPxdxwdlSh4NCG1W+4grj9veSmjIqGL/7qhB+TmXtAuhW7
gNVZt0yN94R812J0rT1IxMV6BE1vwsOsU8Lf5O3KEv4RhO6Vlnd47hfKsZnRD5nF
NvIGGCAPYoFKkjQ3CEwVhUf96z5MsxOTVefmUfJTDKnayDLe4m2D1UXYmaXLp46S
ITNtW5qyKmcIzflwOYjaJLpDOFUBQX4fO7Qoi9j3K8VRREdSleWSg7nmUzbarYh+
Yy6070LNnX9nGdQrUCzEWlVd+O9rsIHYVoA/PWYCXKbstCLCqXdPfRe8fZbmYwWz
DpItR7oD9a+BOzz/KMx8XhLRaEdy5bVvKcGnCMnT6SWUjmbgKS0x+tFCRXywvpQS
nnIGsicXED68tZtjz4dCrmZWYFte4uoYZ/tj0L+ISXEEyw/xt2sryLbBi7UKjkZa
hBJdhIWBLuh1c6u9qUtwT1iDlc9VK9WM64UQiC4L/XFCTFJ0DEQy2UjM0VQqPS9g
BVACF8/3TBwm6XcfZvcU0Aa+pOR5AKt4dOQTCxR1tAhmfFZesdVjvrtIAJDf2k5l
SsSh6AoavhTu1ifuj8aVsoyIeOZrXd2NaikmXL0qzm0dRM9GEMCTsTtB5XbpZm+A
Sv3ICy9R9xB9Qa5FEqCAe0oy4weErIizR+B8ud/iylrEB/lAzQ6GKCE7pgiVMVEP
bCxKPZzJXsAwq9iqRP0I1NL/lxnexwg9E4XTklshciJ1+YhPZ1yiqW/hOsKa6CAt
K/K//JOUwwxAlDH5gScu5qqoswPgHpLJLMtEupZ6/WgjchMFBOz8Zm6Z8esU5kez
BbkwnAS6FdUCQLPsNfsnfcR7HBhF+M6EmFgWVGoc4duRWaXFPKYeDdPgcvlGuGR2
H54nUxscB/4FGhnHWD1Fdv8StdeuFvb2JmMIB3RqxX64mtszNdB6QZqLzVhBLL7G
IucIElpFtefnbZRInQbZt6MnqcsTSX1EvSo5EVw8ESHMDFQkox3ZUNbClsk6FmaJ
5fp9uBc16JqaqfPyRlYApzH3z9oNzYOB0AHCOIUbHxmzFKDa73xg0IsSd3NJoZHn
aIrtariFKzFwGKHgKicndCZfQ3X1fxX3CyE6EnxV1/oRuBD4qQYl5SfEhheWOkAi
7wmwsMEOd1vZQqzvKtH8XoaixP7PoCmpM2nOdXhi9yFw+wHCRIHz8oYxh19JwlzD
jw4E/OIVrSKe3gsL4sRTIz5CEwCa9Em9LGxeAPNj7Dk0xdMgcDc7SDoG3a1ka+z/
JHjb4UavjPrdrAbuCYUrDDhRKRqr4M3mea/lOgl6ZgH8W6ONUJaA2QPFr7AqCttT
kdnF/JjO/xAMpqTfJ+Dullgd4/n6xGqfiJz9lf/wkdOwcLfsPMafLoWermeHJ+1E
JYZExgLrxvsp0IV8B9L4BUtQ4rfSKljeU4IHdH0zVEdeamqdTYey+ZykhPAKaVG4
JK5ya9+cPWeVYefX/CjmSKRNBBNn6vWsot0WX6qkLMTwVciligxX8B8CEzcG7s35
p6LE0Ys3lrEtlDNBQ0Ezw7rXEuS+ePMXT/WH4UC+emV9+tCbDCY6UhCK5bH0yR5f
qzVQ2qNlUmINeQmpADR+aH0Tc6WkHoKVQbe0afmje85+GGFkPhWwXVd5RhO3+nCD
tjkem/3FxVz+KlNjMvfstbaz1bAu/ohNY2AEZ9SRjBo4Xwl9tMyTFnJTgw//DSBa
I0+fpAsfm8QdURjiUCkibLmkMEeY6YrVVDh8YIxnvT2No0QbNR9qz0OCe7O/eqrU
8tPYRve02+KwY4qTOp887OI8fyUlUZgly1xNBzfoNPC0XG79FLmyFaZ4yDQ4n/rT
pzSsN+R2lwNZ0dPSM0L6tmX0iWZ97jraDdjntejB0d52fN9zOAV2qvsvCU6IpNGI
iM0SHHhNbK7JJQlO5TfHLhjcUyxKG/qDc+ZxFCRwyhsZLRV3WFC/PClktZoW8XrZ
T8NtkHxS313M5t6wr4sQJ9y5h0xK8iRC6eFD/pBzHkkSgfMWJ0R4FR/V27jwdHXZ
R9GJrAXlaqIF4exTZZj60nY9tL0PNb3Rg0pvZz3zupgoFQnWUD5Siq9mSZTQ5beC
vb9Pz8U2XshoYuxQQSb9B8BqOvqMCakAGhlQaptq6dnofnC0uTv67XRBolGLDv0S
CA0jrDrmjI83mCIpiv45enGOgUmGK722jbj6dZCQs9eWBDrMAffB8ZYjhDgUfW1N
GX2eRS3k2Lshmua0R0yAi4VUwK6PxPrPpENrCCL1qehFPP1wGE2O+ZRB3OzQpfMo
r1GIj4HKY7RUO5ZXbOa6GU07IgG2jvlzw5HTz8/QklIk4ShjCNHry0zKSgS4jSGe
ZZbav22aN4X4ZPMtG+4ULr9+drB/Rt52cmUPG5bagBja+9hs08k1KXBwqWG32Vn2
2dEcQnPQrE8g0Ya20NDuAjrW88bDfJxN+jCDl+XtaQNUAlo3QnyYCXyEgps2VznK
uzQAlhYjIzKfV2J/AWzC4iSDL+hcAjEi7y7PzusCSGnB0ZR8W7ItGD19VmULGVbS
J40FZsCDnMcbV0g0OxPpPF8ptGweupGgMg7V9RmTXdSAl3f0KQHT2U5lR5mqyi3A
BDONmDG2pXN5iE+VsdGPa/J/RFICu8aiFyhoQMRAIllttevde458OarBPbmOYMqM
pyM16Tq12VOlkB9t7qOWPq+NbmWoW03kx3wCGKk0ZU9bRjY6q6pMOrnCEAhRHBE1
B0pzQhR+HNRuusrtDdcTTfMTnGBlhXGZscMwDJlu4Nm0DjesZQaEHtWzTiSDJOwi
izGcv7TllBcnPWno+7Qq2aNVLhwGE7VgIbxdbvDQmdmd93gJ8aPtz3oWAK+nPY0F
N3ZKY1ZtN4JONGWLi4y9rKKQ/ybrOYPj8DTKF2aNKwlRbLbp9IdSQONrX3a0SBXf
Ashr8iboZ0ctOlyEfCIiZYmr4BeaaOVn8QTpX2EYJWt0WnpITBpa8pdgyll9zqQ+
VlH2Siqz1PN9h0g+jYnmEha0fYT+x3KL5WeD2LTkUy+08UGFgm85X4woz+Q097d2
g9jlSSW+g0utJhna2vbwxdtiXLva2JjN4caO+Ce2NKRawZsE2j6aIl6dRX4Nwop5
dmpyKh+djpyMJpX7Mr3WEvBad3ov71qBl2a0WpELx/NUElXwrfsjQQ1i9m4XhY8O
EhKy4MB8xPIHnvW6Ez7Thmg7K/bqWrNPSFyW1u+psx24LAODFBWm5yCFJvgiC2jT
flLt15KTn/gjDD3VystPGSglWXAk+n+zgNrOsXDW6fFj7vbo6sOueDXuhtzWMshA
9krSPccbnJdw7gIhwgSlzleInvmZNjB2B3EzmZG2v55MY+Tzjh96iQx/P4SQJoT5
PP66E0GloOQKaq5ApWFqpScMo5gxoNGxQr0WQM/PsnLoWIGTxYy408cip/lMaris
yBYJ9A4LO9+J7EB8Grh3QnoK2zdcjU3EZ16Ed4jfRpzjkUAu3vQHplTOPgoPSYnO
8egBQpvLpLNsPwgfhWtwY4QU+d9wRiMvB6Ys30rcsuJCY8jSuqAAYHwHKUbGX+uY
Dw9JUggz27gPE3qe0c27YMAVpeetubqDUwhXonUJ0U011dynngg69ksJzd7rvzMz
zOguotoAeerqJCzsAP+zIcpP3WT9e4T/vyE2+IjX2z4EGTVPH87hkEUXgTvy8H7W
PJbsAZTNfmOOuwq+PXiG350lAdu+r071FHl/ZBmigiOIdxUUTonWAp9oIrx1yTz+
lQVbg71cxvu0nAMQ7flwteLJ2EsmH5sr9s6R6uT8JWF5bPLqS2RlaeoRBGZvmecX
rams10rF5QcevS3QQfeoK0/6BlOOxm3ah5Swdy0TYtpy0Lu1z/nEiBxTc5RVdqpo
l+QoQ+WSKy2CHrYQKqOMLTm7ldbG6IBQLmr5Rku8EVqCdcg5+gMBhfabtlkTKekT
1nWNGgobFoO2gUadQIqgS//1V+owiHVTk8pp1nOOli6RL27F+0sge5jon25XlTI/
CE+4gy1ALR0YcaRRnDJHVCqj4hME/jmtS4wi7z71qMRzWR0OYD7qGtpg+J8lrNUQ
i7UuDtrk/XgCvlgiWynDpOKfMALYp8ElxNCM7UeY44xhuwSuMWjbC9Fazog7477S
IA8txLxjfBGjAvdtLb6iNbaS76cmZfVaJ8fNeRRPCD9rG2pidKtMFwmHi6iA5+7P
g0G2dFXkAo81odxKaJedtMlb0F+SWyDCISqt4TlyZyB27WEgXIuRnJ6RLxNnIN/T
byzjPKxVT1Y6Y4GXcT4TRAdL5bjWFvsUcr8UWbe/ZZXDN1U4uXgb0HqAHNw7cW2Y
6HiouIypbEG6It7JGefjJrO1izJDxsr7eEzMBRe6myyCPa0HF2Cq9sVzYMTaj3Xm
tGd0uL0XUalvcx+HO480I3L0pIiQM3SVJcH5ydGVZBTX5Urkaca6HK+c9h0PU4P1
GYP9sslLVkrW3HsxOP1se9YRU2Qhj5BUlVIwLUiGCyMUvVcRfYAby6bTVLPkeuAs
vCAoGtX8+Tt0MZU9yO+xRwFXI8Bv+IgfROiUUynAy8Uql0RL6WRgol/elec8Flyw
t7xAYav6J6CjedwY8YvT5duBgpz8HCZqUyOxkvVzg1T5jNEpzwKeqx4wxeE35MGl
+UO+RmPxjX+g6mn7EP8x99uqP3o9zfOTE5jogotyfGrViKE46qEGFzdtea6Y8TOA
zOl3nAqUVLtJyzCv8QtJPMJZUxReby64oKzbWdkNyHGjJSZxF/4+4qZiYllB0tTA
ItwvP5PyPkeYe5Qr8kTuVrlGBwMw42OeKDuOk3iPzrtSRnN7G+TavvXzByuIPwzS
vUppIKw3ouqzivVuCIAssVqyaEDDLJgwXkj0yTK5ZM3O79RdkzSVU77boBolmS2h
Z30hu+rcN8B6YAECa5CEf+hg2BPrXOXGkWtzYKHeLCFQm0jbNl7tYeaU0eaIHeTh
OCgFY5oGCS+SpQ94+WEKRB6r4arf2coCC1xsxoEmDtgA9i/F2MMRGxIyvuHHWCVk
/Y4f3KoYm9vMXgxX5xq5wl0DREVOf7AwV7b/9IzI1ogAMlQN9JKRXo5bVCg6FSIb
ch56q7QVv8GXWFsGZ2YhsDeHZgIQBkKdHXHtHSTaehuAamubsNyLoR5BpqBj+FiK
5Er3B4QYVuc9QIW+FXj4Tu8cOFTeyC+OP7TYVT2GTZQDQupTwVqCY+HubMvENqk4
Gl1UXG33p7GG9RCunaK6C6yAdPP8OhUk4ZM2dNAI8arTSWQGg2i8P43LI0yMRXzV
MreAwLzvT5tK8KEaTuLrlbFVJ0g0cM4zPmIMYYwIRLP0ejspACOj+onKPTRHS0ue
b0rTJm+DbIsQXyI4eAwlsaHAK3MxOZuGlnX56exWlHNGSGaLt6AodnAaK1770TNT
9HwOEbtdJYn9S5fAng/cR9q7xB/wnbr98eCBadhZo9bNAi+Yphw+ZIh4ghYxVxfK
f/m6R7rW7o4rv0RkWH582KxEhGZMxMf2d0UyANdOgHuFKmAAbC3hEPA0JAnh35mK
YxTd6NXPZaleKgfz0ugE87KJ1NXLEpecjFOx9ln9lNTpqlqJf5fOKXzD14cHfyzz
1UNfhXgTI/xNwM/U9ETgyPpqTyJWB2COZLb3dYZC1rqA8iuYmSIpJFss766U3ocS
CKhqws7ZsPrvrGzfMZpdGJXMQGYXpAp74yGtjNcrZ0zF2LPN+Hu4BonzdnV5JTCJ
/Y+CQs9UixFi4Va3uH2qIvMoIcQhUK9db0Z64NF4tjEsDSZMTGDCn/tjNZTpprQP
CvUiDDoIAGbfdUjePMNLVd+QbCtXhqKkaonFAzz3ZXKhTvRxhFtHGO5x0cw7d3Jt
2wLypWfIhNyg3bPqsKHnH4eJD1yIpODzE7ilSZ5bFN7b6VS7VCCoBZMX+s8vCiHl
i11aac6v5AtWXtP0c8IUoiudd6vJH507+Xtrm2kyngqQMWVu43aY7Q+lxt5l0cNq
iZYVu7kwkhkg0udhffBlWyUzhKq0vglrs4U9/i2CClp0tHcdZCn9lZdU5PC3iKZg
aKZU2NAK/xx8eb37l4XDUNXHn81pyXPcSKCAxgnJ1szCVMWCRKMu0DnFghDwBsge
NCxdi7gwl4ITAX9V6XTYv6lfpkQFKCLp/mSSbawR5f3FPdquJP35l8JImHZqnZZr
C8/IJlzkZQXTFaw7jgQyZJRytV1HQa09T7rcssgrBz5IFAxgMwVtknDcsrp09r6z
RgC9cKco73ojiAYdjs4mEELAs5zd3YZEcU4wb7XV4AQ34LptCO2dbiuNTCELpvkb
L+3mBdObqbdKKkSWLzPnHjtaH0pLb3uQ85yFXlR9rQVb2z6+gHOPvKBsPmlW4ptM
jQRUbbgBK1vY9q6NWO1o/MIqORdRPX/3nBbsu8W1EdjRImIVqR9ZUwwazD6yD8EL
yEQOK++GHNe1pmGF+3CoO74tyk+KQMbrn6xO/GeaV/Q7L0lEDU/FFE6M2t1+Q8cX
nxsduCLas2xnDt8UAaWNlkgq8eb4wUi7BLTuUmJznMcicO+AlEzWDs8rb4oBaHwa
Zzdax81kCsSx9MpU2NBH0hC3Ot6femv9IWTryiIkulSS910I2lqvy5pHSfXXkpix
AvCQWqnV+GrAQOuDYA2Lb0TjMATBUjIYXy9u3SoViT3wlly+hnrnitD5N3vLpsyf
SMFW4JGxc8gqibTCsIONUertDPWOY/m4GEsLoyvaWB3kiZQzay2PdUp666Sp2tsC
W0ZYcoSusWRNAq6L2jZEtPHZVQKtG9qic2ExfJzQOMLagGiyflmgbPkCt88ioCXY
bHzr2c5jggT4DZYnRODI0WCVC/ra/w6PH+DNFJ0P7aCZ6UE3Ejv09T90a88uwwaA
eK7FsGg34DNfISeoxP/K/j65jGlRWpTh3OuvZUbS1Ca0d8Dds1/gF41zauVkn5uA
PR61sQ9DXjtI3ogNWhj+h44y1WypwXg5JkKvagVK3YG/W+Sv4KNgvT8K/fc8/v/E
FtV4/KC9dPPKnkv4Nnmwhjkf7ldTT20WZ+PFECmGRe+/LTT6T2YAsO87HqxPqyfR
9Kcj6IzfB8pLPWCUuUrE47LhnMIpwqpmimBtEs2WgDnxJL5xdOYPmbRYS5Anp+ju
EWGP82/Q0d7oWnQphfD26NX4O4Dm+3+VzvWQqFu8TtsZbQMhOB9c6LONzetiJtnf
kJJN5t0gRktkJkj5uB/BW/8IYp63R7hfhqbYG9nCtD2sgFt85LPrDEd5itwd17ja
eSYY+fhFnTbM+RCp0oP48HlS9WnQgKj2piZILzD4HUM4eoMH4LhkoW/Uei4acvvF
r2c/SAGrc2RoApSFPH++908ofvH+oAbCqLerIy52hv3cK5YsQ+oykNAYin71jIY6
B5MF3M7CqE5YhYy9ckUyItaKAfKDOSFbchMCy9v3lDkee4dJYCbIhYZVX5y20wZV
QF9YUDOPdjfqJHROobnV5dndo1OBxM6sLZ8CcjsJ0izcn3ORRNLd+f9wCd1U7s2m
jeXHUQmiUsfWPxuhL6f0pwxWsueBeZmnm31likGOjA4LKw+UNNRH0fK3pxsKj+uV
B8/tD5a7k02dzqymShpkVY1q45Goqb9CdeiOux+vRjGKkk6nAJAjKQWyH5J+ORAZ
N1ugfZR2y6qaGC/TQX8mP63+v90nbIaPVI75LesRyCyzf4346P9GUzm65Bq0VG+k
7pF2UsWzGsD+Skl8Jz3FP8ukH9LWdc8aKI5EzyU9alEWQwG9ObijGOEGmDocK8ch
H4riB1Fz2PSBwWENP68uHCA9CXYqZh/giyPBcJfU8eIJPmGU2URSkM7WWPj9SoTr
VpAQ6KSbHeGYXCRP8HgZRVWiNz2VxSSa/7poGH1AkkK93oNJRfWyvNvgbYsDm6KW
EfcxKKnh8NhsYAEviPHo5UgZmynFG4CxP2ovjqhieWAHy/VbalBkSWN5G0cGtvjU
ZW+jt9MNW6aflKjri0I3SZNCtl3OpR7z1ZmnZnO8Uq6g054ODTHDEpvJKVsPW+I2
Oix+ODdlHS6wx9wq1RN4vko/W4xgrIh3G/4iFiDJPIbL8c69gsWuv8PgNw/zaCcp
O+moOan2rzNmO0dbP20AXs7h7joRPdpLc9i7afMiAfVSPI7+KUnVSYS+l/F114uk
YLZ7gvZoJVl4Ao16dITwBfTck58h6bo2uoK5EZ/SJn6Z6HqNr+tFvKTEJQ2tCsdd
o5KazJ45iT1yLYy9Y8t/I+7f5czCf2+MS47rHkokqkixCRmOcTXQU0f92ewcjV2m
HOBBtbYeWlFJztBwrpJFMFUK6EurmlCd7XXN1bGC123s09apIGDyrPUAjMZ7G4hG
ETthc67+jp3wnYn81DH9LJ1IhazoACdBDwyj2bbpjFw89qdYC9WqntHHCgRehVRR
43TxW/HWM1eqIOHg9pkkAYRjIou5QXay4DcQj1Q0ZY+XkqJ2nJt3RZh/onlrdOEp
qBqjehwZiaO+KMo6gnMMp9M2cqxlcIklZDKnmSZw/JzBFVpLe+MheN1F+oDSmT1Y
LHVnCwgq7O8PKC1ZKlpfIg9A3D2LmEPrRrYEmbjfEAQrQshDtVHZ2L/jcZAQnDVm
jOWOlCwFFdKUHjk0Y2khYjas/LtNrxGRH/BUFHcV3Tuycqrqkc71a5mdhbuEQ2OX
fh3+ipgKnb90x5RbmsnAR+fhdNXZ8VrOs3jrvI8DXaNpuSZ12Sga4RsvFHpDHUjI
JDsx/6VICRZX/IpgppLTOiE/6IwFdXvq0TLoDrM/Ud7gjpnnx2bIaiPrSizaa8za
CNH1Cshmftjj6Ebq1GInaRu9D5TSK1N233IW7c2OFHnufwsJjP2tt/SWFbwQDSi+
eFmtH+LAXacFEViX7CzJ7Q3wuiF8T3zEImBGYZY/5f4jWshvAdO07PO0KQu5mk7g
YfQx7gv0aNVaKztC3JNY1xanrjR91YzA4eyKPhXr/I5SRq6xTWlGzMDFI64AQfw4
ZhgGlCcy+qxzeWgHScJu4X5m0QnV1E7GPKAiKcG2bDOL/CdZqtqCQwBYOYxIKhJ5
BUIdKNEUJO5WmClQOy6CmsqbPdRP0CBgZu3PpKMR//nWrAUbKSHUS6O6TJfvTcKq
K3DH9NO3PFjD4/IHphk7ROz6ynMqt2KfL4Y4JbhIeW4YPWMALN9lIRiE1+g/a4LH
QhAW3aQu6jgY8yH+atK6mVTyKH3OJ1YzdQv/JTVTj1YSxpTbdEzUMsdI/u3qrfph
9mVAqtKaTXMauDIWN2Z+rFgZKFzaBm5z9BB0tMtzp0ET0aruj+P38mdEpWC4i8BG
SdBUW/5UYr9/UmGTUGMUtwk7BS27Jiu8HbfDH19DNV7tNueAy8hrJTmZRcz8lEi0
APHCM5cCfNn689ggIyMCQ3sEH5Vij/4glLMXst4QCXyO91oq7peuCDDmLMXhS9hi
Qa+xgLjjODwFt0vTenkXXCXViwS0Q9XlzNZ3bb+C4FTuoXoMa3vkFhaFnTeLgMwv
te4Feq2OMuq0w32hJ+bBvbupKLQTR0WETgzGu/BfEGAZI9NI9d4NrUn/xhBQhDqg
uFN0+D56n7uYLv9blCRuNosTa+zNwPTHt6QIC1VEt9K9hi8btCugKdCdKt64XlKC
J0oieZvPYzjtdZwJEmuA2gz9sl9KpViWozpZtjTzt1rLj/QABSuGRVGVWmMjw6Qs
+2HVdrtFxK0s8EX+UeDxJCY64OhXg00rPxpUnE2Wp0i0D8TVv5xWvkwFqaoxPbOd
w3kIHpO+A/whEbDBCL/qBUlimfiVblFw1ew4yzIoQuAaeVa3jfosobD+IrvdjmYj
xPnH4bD24Xjc4TTwm1lAUM05AUSgrbUQsP8DU0WN91YYcw8L8ttnSMvANFD5WsGn
f/7tdGwPkIdjaUKGnP26axgQIqsmhXAIi+hdZVN532dDu5+gSMfwkDw0t4YJpVqZ
4/lYInCgFvMRzhbCpt5fCzYRh2joapTRxt1xs9sOjzuefkt+vgsgPupsWjx4Muu5
t759gW3oPmQh8tQzP5BMqprx4/GTbmKpQimjJkVdmwXuTokminr+3wKC0t/qz6YX
AXr5mOTN/iSF2PSMJ8mM47Am2nTR9vxWjO9Qmk9CgKGTwvQuugfnku9nJOAXC4bG
kCHGTKqqc1eRRALj8q1pdC80vg9n6OdlZgTtZSE/zDqNK/MeKNZP2aAYnygUTIZd
4os9BRygcO1HfVfbA7JqKVZmrswcsN+1ulk9536MJT8ir/kXol0CH37/I9yC7cSa
Tipdod8/upAw9rONE3QpohcwojiuOWg5SVnbYDGA3puWsY+/Iya4zLASwr2BI9hY
Bc4GcV2ALyV47hq4adebupi1Ky4TJsTZJnyEb+jAs4zrUq348Ja6Q20swMCup59m
yH4SUjsVxh+k3bp+LO015c/ZblIfX+rnJvZOp4HS9gXjpNUqohDDekknlhqk7uZc
zzKCpF2HZzt+W5b/Dq1V7E15DPewNHVIrFlEFAJrBJEVWmcO6VtfOqY2r2ptLyBU
xQAyppK1RYK/8s1TuGFUHzy7H6UpHRJFUtEeitLQEioW1oCOhx3b9pY5DSKyEfyP
DNcfrCHXW63hk1nShyqQ8JmuWa+Z/KVPJlvqvrCRX2m3Yhg+co+3tjQ6nrWAFdGI
9DTJdx5RlFvbHi4AQer/VHY7NFSPgV/ofTvtSD/OuXl5FImCh29tvAFoXRu5ULL7
ZzvEY0exhyuYVjVHxAonc3uVgLxUPkyRya/j22A+M7R4Q2rJ+kTaejYdHK02R2GV
CaFn4d82ZVZEjQhuhJz0E5BJ49gL5vfYtrhiC83vSq3V/lPTW8pj7DfXpxM5kc/p
jAy5VNyRbBCZkCEISFFX+zCv/zkPl5VYd5j04J76uz5Ph8wtfZePw2YUTsm5SDkk
eQikbkz/AGgAl0mqnirRzaVz0pFREzWo+h+/140oQG9nFQhCQe5fh+KBYd3+G+54
+8AMUzMjoV3KKaHQqc9DLc2RLxUeJ+OQ2DMO/G71kNkR5Y+V/VGT9V/66pnghr4p
VRAUAtqqL+tONorYH0cQwyEgOJD+UniY8KaESniqX1qNjZa0nkQCT1mMNmG45w9i
G3eAh6hQSYQeh/WCThC/hoCgqweCzJe8DdNE0kGEbjjhsT1VTbDL+3lYLOGPuP1t
U1vlAqbw9xEbMFwUNNSJazGkx5AHrfxgGraqZQqLed9lhT0MuiqF43yLaTyautKr
Jqll0tdfmmB3jgQAEiRE8OqF3nObg7ouLVa5xe4SIYj6JZbDXY+BmFAMJP5wTli1
sF+BCGQ2hcTM9HYq5HLApDoMxgNDCrtlS3wG4xj4LfYdUIkzDwBsaijbFpWriXml
DX5oyQ4lEfV9+5WXGM1G1ybuhObo5wZdkl+zaIt62bniHlZXgPApqPbiNW1KnXLh
C6jb6ZL0V0lo6EG3GU3GFzPNpvhHLGwgSjXpOA+f4mslYPosYjx8DUtbu9K268zr
XAXnpy31wcArqZJxEbTX0EssFAjDqLnf6KHARz7DkkfCqolZid8b9XPw2D68jw1b
Nty2e3BMKhfrzmM5ec8u+UYizhiOs363U1XTk4jZss5VpvraHMy5mdSc2ctPqGzq
nuQKrnrMYYHgzRzb+QFrmudqCzHp78NneFrfYzTzSp0XmXlBgKBAprTTdVOBxRjz
P5mf4AVkmJsCad6PZoZtYgdqSD0eqjCIbITkuCXjUTKak1PkHkFtrgz+Puk8BhqT
bmEHuInkW58I8M8xq7pV4Fm7gb0jS/tbdewBtWYS7dSZ75Hb1NwJI0mlttJPvWcR
Q6bMyxEODdJHiLfsdN/cO1Gm61nU2s6Mf95POO4jrsLjw7GkgE29yZa9ADY/Fmum
/Ngcoee3VA0evAYpVrFjldDsoCuekTeT+Rzlf5jVTVsoYclI48AYcm0LGAQuHsyf
93ydRxj8G6Vy7G/ugpAvY+Lk1ZsI7kvkK+CfbGsDy1zCpTWKXL0hrcye0Z88r2I+
LzMuRrhPc0QEzDpaPc6w4k8yRUR+HqzELqhg/argr/57E5shDWF7ERsuwyerbF1m
1GMu0bB6lA7+ePgqE19c10eM9UeHKqDIG1jwUqsp9iaJeFwTLos2yY07LJwi42SK
noImDo3ABZzyIuxNitBVw3qgPes1rVCq/1HX0RHGAqAeHN3nZF5Fwgppgc1wkW7/
sfaCCAB64H1jy2FL0smKvLcLmsxwniKa6Gt5bbCFKe0cM8JneuHhIyNvcQnvctUG
9sL4C9zR4g+LFOkceV3pYgq/bBqsU05VQAGXcPEk7I5vHDInBorDMWqyAeuMXwPY
/qrPDtG6QTTuCpxl72HgmiMbDrkxi59soJqH1OEIFvv8vLdf2WuZMgM06hLh0xuI
AgiMcoxcIzOULSvKbeCjS2kcJCCMs5zB9yEkRPGVVz1TOrZvXrfcn03eMLfgGAuS
uBecthqkUM/cyDsYS3HwLNziTScI7xkmpLBbdFPBF09L2MQToM2LFhX9RlQWb7If
+XzQ+cJ3UhfGutVUvv+iRVZdjHTeUjU+Cd2tdBKVX8ZQJcMWqNHAuGKnWOc7/zVh
DRQ/CPfxXFo3fNFYjWGmyfIsOP8nO3KCoFZAbc2eLr2Dz1sNA9frtCkAL0bWbZyk
WGkdk6PyGCHHGzk8WAwAGStG2/R+amgWRVi6kDjIS8p1QuD5fKBJknk7c9hJ04kd
EixE41wYehvOe1hTbEL79mSOxxjliA38ne4zFPIb1fkBTbkGfWUZ0MqfV4Fr+IGH
/qnzPmL406/MooBy2zG3GoIQxkUJWLDwsJ6+Q7rLHc3mKFs6NErGf46P8vHPsJco
pv4+OVmOyErBcV/PJomDz9eCyjfJiH/VlOtSf91c+Hq7PwXlWKTdH5kh9Pu17WWT
Teg/gS4wKym14vC78Mu3lac+vtxvNumbVwn4Oiy80n+0cvuMG18vHS71TMoHQRuF
pTD8+DBevB9gOYjjPAUiUryYr6MfYX+m6ufbl6ewltIlbdTJEFXgllrxIPdlrqS1
NTBVS43aPWnPPJjUy4aD9EeoMWDLNhgdmL0QgIm0Qe8dhTT7u6/M6i/uP1z3vUhc
hoJBkOS2NeszuAiq3LkwkE8LjuPJAgcnOhW4hHNI5UO4uFJ0DGh3/RuZW7WqZpAo
5DAGSY8zvEdVeblzrVF+CB50tnQZ0YKCvqRGjM97TmKaxBLg1Q2j3v57E1mChRAS
GHu40EtqOR4HsESWFxFvj/a1K/tOxGSNPwSb0Py1zlcioWjiYgRS1mHyvN6xYg1/
8xgLp4jjuj/i4Ls9fpPQoeFNChRMb8onRVyFx/tzXmLlV6O8h2VRHdQqCIUI8GJD
XZeJUtV8eP7RPwboulquVf6/i4Bvl1WjDo4CIbf7TGwSfbewCX7eYtbhmYoL/4t1
QQlbqPb6Xd9qLeCxFe1mJ7FyTYGWx5+iGMFIThiJDOy/CTstSefzBnrJX8wTCTn2
t68tb+yGJ6mT50v6eAQB7zCi2V/7fVWqm75UOtYZRlRal7JltRBGLTPgNnKgcd1U
V43x7yKeRU8y+bwpZROBhxR6d6OzOtUVSCDni4gszPccC1F3836e+wLsRJsZaGJg
CtQAENP1g3jHBzbTlFMGzPjzQtD8gWtxV/6oe8UutQ+xD7oa2ERr4EU4hToI9r1Y
YAiEeJHA/mA5eTTnqi0FMkLY4StVqC23uxC6Rs7PRnllQN5/CKoW/AfrP0jsNqyl
ISoaQYPMIB8IvwnREL2TBVFgDMTujhGrlM5IkN/kjs+RTyvZ/b86h8WvoKSk529T
gci7CCRnKzb+z08vdZtYhACWwAACDZg6Oh1lKHY/gU1tQfpPwQOFMP+RdfMYfg7X
K9HMmz0H+BXboqoY8RYu/zo40vRvtBUn7WMXYEx9Pm9HlPaXK7+AcSmGRyH5iSvQ
KHsfASVbCrK9SI7Ss4faO7Cnjc8jHDvYLADCTxHKgH+wzCWfqKiLcpzxxvWrErqM
hgKN0p8RIZQNMOGDVm6T47yeV+1mx7Yjkn4a4kk+W50Q7esiM+7Oi6Y7CxUQUj7g
kOOFeoQ+9EtWlGsBHYhuUW1zQPQfl2F6l2xtiqquoKQz0pYFDsFH//ovP46KfYyC
7ZGScvxlk/9IIWasVh1YxiK0HCtare5lGiX/Cl0FZdyfSuLWcsKjrPB4NCkAuC3h
DNs0+tcRd4WFwsSfyE7B2IoZJ5vRMhs8LslK3C71SOcU1deOwza3A2WgeIGnnUZF
RsXLG7ePTkAtilsmi9Bi2Xq2RdEJzSSjX3hhU9YcyBWdd4Gu6P08ZkjXmc3NXkRR
4CGBIWJ4USTTsy6RHQUMtqscgIz4FRLphkv8vn6VTuhLvD0Uo9yKNiDimcbABzZv
XTEd+d08eOYhJXzKd5+LdIoSP5wm3FB9eLvgBNxNYjFVyYFTLfKCH4AW7s6O1fmu
+AWt/QBV+dpjS8Tev1aHBwTjwDaUX92hNtS+d1OxCkFGuR0Yyw/yUMJQiXj6ptbO
FK64l/RBc3J4jHZgx6nqN27mVIUB7eVohapzPZ18PpiBYjW8I7A/PdGDyneNDL7e
aOd3nLUJAzNcUrn0e8JiYO9LDAgFwYpPaGIys/h8vlAqNlOgLsBDmel2wP0/jBh/
SzGYIjbSYzwDplGp0/9DsLi0Meljy+l+u4fnnLlrdVvAGPl4++AFvq8PwUT9MpYB
BOWwzXNFeHFNtI68TdQvI+if6OAy/H5yPSzvwBUIJl+wUaRUOlAgCblYl+yCLE6a
80Uf/wnnrwPVBR7GPz1cYLhDyw/VW0GY1stFC7pTkourL0khlMHFWMFi/XezyAvK
Ga5eD9YJFBLhP2jGg2htEXrLBwtxYPeR4qF3ZNLN+mM5VijZpWKdEWgCR50/Q33q
2nHgvY9Bj4BDuxG1hefnQybMZ3D6uNGrAZGEkEig1DGtlnbyFXNtdmHCrMkxPMIW
FPhhI49aYL69nJnLg7j+sZ5zvf/5xX+wzZ6cv/IuAiJfwvMy34CWaY4HzpsV/9AM
fyX/WpFWa4QyGPK9ceyIdrPUzgKTNCbKULb3xLG9i3KgjjtuRAT1+uj3bxNdoqfJ
/0XTIl+Oa8R/ARFxDek6RvUtF9nG3U1rlypJB8oLbCdP3pLrAZmH1nyek7Y/mFes
XZ+mzTSe87FXFVg2CqLTBbwKeNSpMsfQzaAuM00oBvB5H7/4gzj/nBBVWgj5A3ke
LzAX4Z89ps5VO8E1BsxkWqeSgk75mhL3OOEZLIQQG4GEnLjJxDm0N/ds/75uqujH
kUgjLyavcQBOpDJReU2lPPgaU4g4YCPZKhLczQvGijZbYu86GD7uD6CwxRmVqjYj
NS7rPQb3Ie2a2NppemKdfPCucGW6XTA8ibzI9SmtxJ4XQ9fnb1lCuZGI7DXM6C3C
hBpkhHg4LK7MFsYLknngkfilU09i/4DHz1SGI8LhZjC71zpmbAe9GUv0T/NHk19y
fgOvZ/6uatbL9TjeLyyGC8XZg2E5BKqw8vANv3PWjV9Zhn9q+IDYO2LztMT62Llv
AQkRXD6J5ZOqM9OTkEBvjAPzgx7qI4+Vzz3e6+DHVNIrit33n7bgOE6jvrlNmY76
nMlo7VbQ3WZElL5aPSJ0wcUfzzRfvKn2Jn+P/I5Tj9Xy+bhewCzl+SYYjv6SCidb
+okn04+GCsSIrXNDLQ5ghKXk8IGrRnKLB50I0Y/0FFxbhkHiKBhJn9AA9kUPCB6w
THnFHTU56BDzZAsmvxypV8gOuLNeFvj/FdT9qmE20PfVQWcT1co5Jb6x7uhGOLVH
AudYPR5t4ab+5jMqUxQK3xRMvnKTQ5/hu6dmfDTioyYPQnvDH5seTpTd03LLi5+y
8A5tEDkJ9QkVxT7VbRIeEdr5TTS+7C8d6wF/lPvYxeRrC2BOjtgQFTfP2E9VGBIN
dH28y5FGTjiweGRvCy3Wp12uY+GAVqc5smLFE8yYmQsFM5vi2RhCaUQpSyG9c01V
5/QSHzzXrOa5J9casN9jBuXVWEWaJpq6dJlrd3EvdHZRz8xj8eNNh0J/g2PLiyrN
WftUwRfwVrPZTlfjGkPPEfW3dRabcJDyR6zjLJjIDPo1RlnAya6QpGqfVSXs4Oqh
6gOKRwWVmIVdCUHaXyJb2KQofC/ILnZ6qWZedRTbcQqeO3tniYZNSlIIvSm1MnRr
ZQYnAT4rchvR+UFXGW2hS5j4PDHRyFSYmP+VJ6WS+6SQAQELoWemyMn3sOfLZfLj
yEW4n7KX/HdlGcCL//ynBXEtLYQ1pFVAafeGwReSM+5zXHgVLBKbg4LL/mhmSPox
R1mOsi0A3YVCto60K3bIGVWrj79Bjba+vcvebebdDEsiw1Oq/6nQPN5t/09tShfI
zSi17Ptw4ZJdy8DMP6vSpux776vDBYtoLGiBhuBS1WKwBiRbULLKjZ3n+Z0Qldqy
jD30Xpv1O7Hn2SiDA/CJpBo+5HHoYcS2GI3YuoWjrjpHfANlnRhQ3R4lfrUS7Ti+
RKw9rxoibiQI09SmIIOaH5Y1CkF6cTR7IPi4FD1vmXrmtzrmQMhEoIH4AsHsctlX
JduKAQc7a4m0c8ZurSDHH6gS19l4o64k4YQDKsjufaShR9FMUlZtwNM+4dHPPqtl
5r6HJ76b6WKwPRSjG+rFlQA7kqRlOqjqdmZScKAOR0qybkuWmZXPTkUaGT9gwFME
5bq/uJLDmjdgr/jf1sSQhcw7TBoW0sW7DJRf+w9EE+gzaaZEWaz/cUBoOua0eK2y
DuOjqStz8b8dgxpQeyFQKo+acLvOtBsx4ms0COe2EygCfh9GTWRH23X1WLfMfEu+
XYO/hHCBMnyMrlSgy6kNrEpOko8ljUxiApJobyyV8m/uhWc5H4ztC/kpZAswwTHb
IcJs0PWbmdEY2sAOkWtXikjxYBs00qcOC+dicNzCqsVhMQw8/T5gooLf1sP0iGJf
T+lrdUqLBSBBxMGA3w6RZsGpl/r/dcfosmHwhXbAjNaVFO3nIVHkBL+liCpWbUeE
PHsyob620r3K4SoMmqmU9Nn/OdV9A7vjpa1HfUYkrx0rmssWyV9Hcx+fMWsrbUKq
HaKozn44Py1rxk+n/HCUNl7LRb8cjcIqBUwk4CbA+7QsJkBJWg8VMXLakKe8dtOU
SCTLso8jRIVfmBfOAWgpZCr4WSyB/RYvgMIr75DZ6SnvhUDms6ROvEqPt8pWod8i
TB2L2k48uNV3TxqdU3Zbsp36NO2WluYaSlFdWbasLodzJAhBuJ2BXXrLbL/k/2+j
rgQ9ffw8i5C+XMtsbbJrJEsa9AMUU9omnWQQ2d3n1hn7/tDC2Ytn0eSd6CkFmVK/
CJW1qzA1C8HplOSUm32tezfowFXL7PeiKNN3p0A3eP3mlCAHgxYrde1sNGLDUB7r
xqoiByYZBEkezEIbDSMAPqWbSjNyM2kJ40WVa+Qzd0RZc/z24HMY41ASGmiQxZYg
ZRxLfudzmWOFSWMZrS3Tor5K665pBjmnP53TURKTXeTk9CxGa3j1BXWZyrmxYT59
9AaQ30hxVinypQc+Or5wsv8QnEmlIERmd0Tx8Y+F1SfCOuUw+cepOmlp2E265D3e
/Bi29uBSl5Yp9K94Su3ObqCgX3MezhrZLSlNjepbp3AyLYFRBzhxUOktIM1P9Hqu
fHsduiO6N+LMpSNreRAkHh/dRxcWGwg5qk1dzXgPucssR7KHebdsosce+LoXC1Bd
x3dsMDtPZmgST/pUzLpOSdi2bqrlqaK3dmrIa/UXCwG8YcG8x9Ep/JaGKnJoExx/
E8aZACY0D7jreazlROECI58/pX2vGWbuMBbEoZSvLFY0U8pNPgRVKhG8ro9Un2Di
TC3y+3+oBr7JhGlkBaneGlpddi/iv0DfZPfuzGFtaTxtSjxXF094wMAaMJCfFzyQ
vJJsUj6Rxv6fiyYaJuuwC4kjhJ2Se+TRcGCJ9jP+51KoWDhT5UyTC/Z5Fv9w/VGn
WSvVZ9m90GDN5dQY1aCyOmM8QwQl50NAcX0S4Kh8LmLkSq94P84BagTkwPCPMU3j
LMjV1kR4i179xj83a6v3RabJa8yEzGJPD06fsPjJXAjGYftcepFrZCGRjvQGf/V6
ZqmBtV5lQOD/fiPUkqAqYOShqUJMAfwzTGIYyn7CsRcix51u3M7DutIZ5odMUxNO
sbt+8vRMx9tgNoVYa1HjXhPj6vbldgW0cOCUZIf3pJEXDqRo3H0yn5I25pU6fuu6
ViO3H5gWT7k9h9lzil75A6SPCeZnIMWUTkm8s7heX2z3KmDiJ85sOzPLXEY/UJVN
0j+3s2WJxhOd70OP1MNuMoEx2cKjiO4nmdjHRCKdMpHoaWuUuLfqTNSN79OYwDcl
OcXEw4NeWSsLLp1UmILgKQypstLQ/O7/gDgWKD5D2a0+239KYRQm46kgid/0zHZd
tUzmm0/5GxQ5ZKJLfDKqZmxeUaVMQPf+vER2SSDTeWmg/J3ZLQg8zKNUW5dUNwxp
3uzb+0MW9UoSvhLDdzBvQHGxZUousbWjhNE54Rk1X+S1Aly3VGC0RDD1Tz7gaVP7
rZUe/50V2qTVlEBS7E4zj+zpzmkTzvQJ0i+U9DHmCHtrf43pTj3kaFx1d7h+5aBg
3JLxbgd8oH7069rh+zAg+YFflnxeuqNX96+uvh2NBwyScA7WiXIxs3h/I2TAlMW1
VConc2fW5aikgFqbhl67FsKmtRdfo0LyfopEoFjQkWxvGlcHbN5DBF1Tzqs4J5LX
taOTuGgomo64Zl50ySaCPZxZmH8LlUS26U5t0t60xzsp1R3l0LMmrpAEhLor3lBu
j7ydFZEjPQ2LAANL/jRDoMPSurxx3PLyUyy9IkLaTyUQzWg/aHjYlKQg+MftOE7X
pGK9IiAGNrnRSW+4w7oZ4hH5UBiS6DP9GQlWFU0rjCsGDzYcPZCddMIVzWZJampE
WmiaQzpTj+929GJMkQNYGfQuIlm65ekSdwMgMQjqYZEHWTRSFHK+OD8MHFnULELO
9QR0m5AcCLQLeTDwFTUtWKirR6Pi/cPwO2Y5aPdVBqAYcC0fWOf4ODUS6BkkgeYq
ujLdzflmen+PScR9F0y97N7uIG6Al8zXRwC5u2ljRgxHioS/zMwkjCpfiRVlqdC0
1GgdmnVcndoX6Oyx7Xn12+9BMCrnwTWTv+TkG7d7swegh3TNwnTMM0cMcKs8iiRJ
kMEsoecjhc0SZ6EF8UPBadrPgPczrG0jsD7SPTc4E3DOUxH4M4FfHrzfh4Nn4CzA
7b6d8vwMzw3f3b5hUk+Hy5JN7g2Cq5S6/UY9jWhy5rwGNy2SSc5o6GIgJCST+57K
CBliQQl7fgupnckGo5C2v8bDs0q6UgBrdyHk+L7WzXDHSDmuNz+FF99/PHTTtk6A
Mupp0qO/BKKlO4hqo+sF5zEqJki+svF9EJHmKVkH5ZnDZtVD+qpRpxxCbD3iiq69
Ba5588GXDtuzMQWwLVFC0wYzaUXn//m4paFr7o67bL39hpBZGOVZtu3JfVaZru1S
++NdqtvrhewupHHDIoAVtphvUWwx4ZAF4WhaFiFcbaRjTKgYnlx8mhwgZLd0Mdz4
qsZ13QwaUBRSz3pQiVBiXyZxvQN3mtJrBFj+KLMwL63IBGUESAgJtxbuPlTT5rRv
diwBFJRaTfbWINTGMY0XCecUOH/JEIgFBKXrIpUJWx0PF98z5JqBAfOU5/+Ad+R2
4ExjYhR8J3/f0jcUnlWkJHSU47HYi+m0/mmlFZ8hKGYWLHax72Ij3yohnpyrDb/Q
vfz+xQJIcuYPhunC0+tC2JCeS0vK/E/VCVhEud+PVyuD725XMuW+DN5w7Q7ScB58
VMqPmcqkhE4GWN4Kd8Cys9Mba4EsGUgdSXeOxRCZZzjzr+NL7RfKv/DWsT9bUa3/
ysqjG3+2PZtNqas3G4MYoMcrh/MjRAMiUaUbHrWL3v7+SV8dNX2on0boEw2TsoZW
un93SZndMXPVpedDeXLubXkT4NCk3NPhocx2cX42apPssNGnRK47RsZRiy0Hjnbn
/eXr+nIpYhxhdETLtb4AlpD84w/p1ncnr8mu7A/qvmRqPRjjf/uY7JKSq3THBogt
kjxm9MQEnly0AXeV2qOKZ9A19E9ucznozJWxYkXvUZORAnSuzAfXnh1qk6hfrug2
XNH6fXtRvAdAD/0nLvLhMbcGSaPpQDjWEj5Sl5yzYZ/UuYgZ4+qF/DctwLxXgg7U
gNxudLGeFAfY2UFFQHTmIzo8lskTzy6OEuRyh7gn18xhbn7gpxkZbpSxcnrgim4z
O5c3/X3Fy2ekYlfJ6VnsNZxhy5MtJpnqcrJwhDkjaDN9T85LE7hrIFtnRkoBJTXk
PvBFie1+tHaI/BAalkEufm1/CRv8TXiIGSbc1t/ouyHD8bba/eC6Ge2z4qQj58o+
b+/YNu103uAWZ1epMoSJvV6JIi2tFJsTYs1NzP0bEVdie36ODuEdGa09xeu8qiwv
ytN9wQoJYZ+hZjeIFjWgT5JUfmBS27osd5EXxDiEUkmxosn9V093l8a2lAhPZpy/
c9hc55dRtgn9RHJlP+CeuDhgr9V77l2Yuf6tOeAQa1Ao45gZAoaEx/fevsLxnW52
V0PQQnqQPhS8rWMqQ7Fqf/cOQSFI0gAX4q+EB7FhbXnXawTOF3FiWXJbp8R6ckDj
vF1Owd0bN3H1TwzEEeos0tcu9OnHo1V1NCrCCksb75D2iFhXFxKSz91M3Dq8fUgb
xyMCvdOfKEWnhtf2kU0o5h2utKb47Xd4yyfQI6di/AvN6IFwDYQLGH5huMZucQct
1PedQxCjmNIcNe5kCmMI2dfHRC7gGxEQxqKAJ1vbTZL/QDoAhQQlDcB5TnTHKtFI
gd+Z3sw7m3ERFF5TOctjRWWS8p/TAorNBM6otdWWzi5X+9+/Om9HEAqcjesVhJwU
/vWrho6rB6n06IIvy80GaQRVELl81yJZKCHv2zCQhDH3roY8+WyD93j64ICYKEhd
YLDr3OfMFP3JgGH/IbQ0pI8d1ElTu9Llxe2wgnb8+Ds4i3xN9nHMm1/6vUvbQlK1
VbF873Qhn7WQRSlvaonsqnX2UoedNJjz5i9dcmw5L0W/4U0UL0oC6NdeMFcwKF7T
3aiiVzMVgSCxyUal3k4RgJ32ff36ol3Qzer4SFsXslZ6TnRYYktR+BVp8xEwUm0p
SHu/TsC1mEAJxYGKVqDNYDcPcsW3NWa+I+FFUUX9bcJwIE2ZvUuLB3rSPGazlSH7
Xnwm40XWbbil9fHUxIT7tE5/h69yUz4oB+MVIMaAPueGweADKSw2p6JZgD+yRjEq
J/ZJqe/zzJmRWaDbYLygGce89SJjzvsFIbO5nbAJO5rUyoWGSss4XzONc2KUE2jL
/t5V+iCxydeCyWLwg1XWMpoJYC8/TUxABogGJUV32me5T9ttwKKk6oUIYuv9E5Xg
a023JzkOJyTCjFUs6si8n11A40mgUxVL1RzwojGHvEHIJ6lI6SC1uWTraUodzXEF
95eomwnLS8Hy0gk7ro3ddAcLaHS2cGFgwQ1kw1hj3oRat11JZkUoc3L+dz5DirSI
qyFeSHDcSPCKyhofIUHtjvM/T4wpp5VGs09eyZlPMZUsCELM2+CoqMUCsd47Xab5
7/5+2oxyPSL6EohMovAMnrmSzADyM+M/oWFHBd3byJM+nQJAuULnSNMMT5Hr/9Xx
fP2e18RtPfnlqa8SbsjcyecN3YNdhLl62bX4ZLL8x9zKzhdtn2kurVTHP/f1dko3
JX7UVkR2ItDEZMW8MtYV6oBSseTqPN70BwOUlvKCJZDyDOHfpvMa0YPyblEoSdWA
Cx9kJQF31/pYtNJbqSJfLh0LI4YDlnCIlWEJ8O7VRGE8RoFrnLqNE9ulFbIke9Qb
wkvUWMvagqrshlJ2B0Pm5wUwIn6I1IZ8T+upHzfdKa1yylnYDjZY7NhbEWuS8EkC
05Bja3VO/s+T4XqTfqak49gjtPo+/yXXxyNpWPwcxCTjoEEsvXZ9sOoYHIBWLwqs
ywCVdMrqCfkY+2zgRLIgmBQj2sm0wnQjU12zMTljPAzNrfZ2Jfx8H0l7mG4FsAPk
HzUIScxbsN+zTf6EKg9jMvazkoE06+UzDImSfsUmU/B27VhJ5f+ZdzgsGuwRQey/
3CaP/P1vwu2Y6KMvdD1jOMB1XZy5j8+lHwE5hydGgBhqLQW+15QntgwmLpBRa2a0
AJKcq7VLBWGQkJ/A+hAECxQHnOZ57e4dj3+lkZH1BftxeVCsnCgVCFGUYB2wy/oM
Ha9v+dqryjTQRJukzRiVrjm7j/O2sYUKAU3HBOQuFD7TNkOKREgMjimV1FijYX+h
q43p32r+mb3saNrw38TqFR1MfDD03wiJcfz8uxq/FSgr9ULTBoyzi4u2h5FNp/o5
rMTnCrYqB8Od4XrtfbCrJvSRPIhq4JGdwY0Imizytdvn/z0x8d+O3gpxHmjtsGBl
6024/3vSPXpKQM1PF7c5yawetscYihig92z5ZmU0EoGksto+ZMiYnUtfNMuiKdfE
BzjTpIL+mScnglrzeH52xbjH2l6OKT21tJcVqWwCuFNiNvhubE8b/UiD/oMpF6Cf
R5P84t4aR7Wd+uYEuENujKrLabN9yjmpq0EpxyOwDbKFyZPsFsA/T8kNBFGu8Q6/
1TTNdGUUwzW7bu5YdCAduP6rWU34UpydDdcRR/E/MizLh1jvrdx6N7gqz+Heu56E
LK9zMOiq8ptHfNQn2F1jkVqTuKsWl8Ov+ivvo2PgJb7uJl+GsESfK6kpv3anJ44r
AEXAU82DaIyO2A9zljBrBQmHSLLHQKnVcsFvP4mpxIXfmHzQPpU9Mfi9MZUMD1ae
5eFFvFg2ay6Gp1+nD6UpyyvZQSYvSJCQ4vqufafpjmfezOo/VoOL+TSaWkDJKkLB
VMLMVXmBUz+mBvS0cxzfLvowv91RhejASXXyWlq3iensDLYL4c4tBSNHY/rHSrA+
SwVfrmMctAcpB2XjjSqvBK4WBEeKOp9JzRRRuhoRiD/NShZvLNaQsLTzqAo3bxxr
Q1CgsGw2ecrYolJxlpoyJSd6nftzN52PPD5gnmh3IdQHsAYV80AsNwlZlbTOvn2Z
07LnxAfWGQjy4VoAlXZZ66q/oGcNSUWHhqdjMQuzdp+66q3I3Hxwmw/De4lAOk9C
allmYM8VKwlxemm2fT5rq4nk8P7mxMxi80AYEA2v52xGRizLpJHvM6lm4H3qu1V9
N91eY+G+ZAofMUj011AdmE7Y3GqB8ES7w7DYBqrpYKkc1upS7c9YcpZQ/WTuixsD
NO77UiHoKu/asUYR0EawmkYy5HMDL8OtrrHnCQ8edd7V/U0cRu7MUIfUOfiNhGbx
2jZ68ItvS7KO/KgN0iTlv4ebeCTBII1vs43i4PoFXac0z1Ku/9kmufgtt8xU4XHo
wb85yQ94VC/Q/tIeBPAxoRy4D8kpUKBNb1jQ7DVkv5OwC52kGEYbUkv5DoXAnlLW
0+W69nsgk118MC1dTL1YXwvnMO08WVql+wocZ4pVkspGLnFve25mkG5v4puC7K98
FSIOy1hkvyK6hCBtmSdXQ/2QDIkPYM7kZEJnGr+sZu6SmJ3PtC9EdXI/9dcCrPYg
oZVnMzkvnuAaGAGobYwczM1AeXqvP8vn4AJylnbxLfaEZXuuAZv2p7bjH35KodCB
rJuo4L/56oh5Qvyk1N3jSNm2Lyq1+il7cZVFwq6mmdQiAInzkGgv9WOZB9acYWFF
HAlA74ZTQYVN8bcuGnbR0HBmzieeKYy7H40Xt0QGKkxkPyQ9hhN14VS4J1I1lkZ4
JodeqZ2IrExfpoEZG5wOzQ3RM1xS7VjV6264AY6aLjn3jv+z9T0iZuG+u6MIHj5H
2540edbICBEQwEB8QC3fioO90uyxzFAbvYK9DivLUo/3fakan/TTr34OtT1QSoNU
coET7oAYFMdpMIRtE6i2TBM2x+e5cRzao3l7QKm9LQrhP/RJ4pRS+DcljGAnNBPN
auGB2DDbrtaq76eSu9nmLbDt6MhsQOQ5L5p8unMFcbdSL/gaOhkvWQ2GH1yR+wE8
OVhcH+sbTBKvMAYnpUIXYpXLJxL2x+rrCYuvkKV30HFrOa5tlqJjboKM6mhU6NAD
19ukiMVuW6WeqkSC1IPoE0WoK+Zux1aUawQdG3AEMnH5p61RCBhhJKEY7CeLa5yD
HpeoVDBHAU4H+NDUCI1zc0KtzpwecsTJoOrykpIm/u1j+9c2Ys2J2TfuYaVyotmN
tgX4K553VuWcM9Yh4RruZVMqulk26HyqzJKIAbo/k7XN7lRbhrcb9TEnVBxpJwNk
QvthlXmcL0CF4760FOYzDsMJg8kc/kG/6gPDXq2cBp3mCfz7TbK1ulWBV6Ijdgul
e++pWLFqmtWBfhu+4xgu6ph5fznGJxDrWUkutEopL8ovn3kBu6QcaZPA/QB8FLuV
VAuH+SbFgK5fKEt4GIy/Uj864398jOE6TcxeLbhej5k3H7ir/RqlpQras1pDv+xq
V6bDC4a84bTFMvcHyYh4ZY2pDjXNReCN7mvh61uQcxRmDK0lV8ZVGNqZ890rgICg
gVeZ2BrjmivJwbW21ZFlSvllz1wpgIRLFwK+7hGkPE4SV+y8Vsn6+Hsb3HKTKFJf
gO4ueQO6a9iujr4a0aQtL4Ws9LP0GN+nms1Q3to/8fesnVRAr1Jr32RwcuqhWoi1
xVT5KwONzSFobroZlSYbIbHuFzKEA9qZFcM7sO69cWAtyYeDRRSBgtqCRJSA1RJ8
Fq+9CM36/aI1ysiJcefuBn2eHkaU6GyJNFetY+yfMT3uMNXPF+WFzKbM1IEHTUWv
dEEdTPoENaVcj/s0I7beocmP9lF8tt0fBtva9P/KepSRM8zb+Prr5jp9TAyWlqrM
e/lEIJERzU5lmUbXEazlIMW4MFgpofn+jpRswBi8VxOPx80kozAy6U7cyQs7ofKn
QCdV8A+Ijqw4m18shyKP0Nhl6O4BrHDHMaRrNwFlZ+Jbs+5FmVrVBGA2MMaIPXnX
y1bgMyD6pzgWjIYEVe2nl47NScYB27YHWsHLvOtKRPhBVvxyLJCqLV1TVx01J6+Z
8hEZAVRgYjKq9g9vHpb/dKDiDJM8RML/1YhN2JGGdAFltiK+7wPj+QIfZJxn8lhg
umWvI9JKfyhNkLyzhD5JiF9O0nCPEUPrLHAu6BCeMUaDLzj17UcygXgRn3BPCBI/
Q+VArs0ScAbE80DZU8qKFj1JH4U3JaB4sshwhTrkZEXz+zYi6EtjEmSqSqHXUf27
7rZBivzczkAfs+6Ywn/3ZBUVhLbBYkvg03RMUoxs4F4Qcryu/dAcDnYvW/QMdIr7
vPi1NiQ9+/Qhx42yU0Hi9LfPHy6GRX04EET2i2DGgtgC58LFWaCuJrwkTcmv4k+x
d/xJV1Rfpf3++NX0QNs6rECkzH00BRiwZaNvYy/YTtruwCuovC6gRn4gB20mLJgp
vILB5dsBWyLjZIi8h+nKkKHawQFDvPuJrXGbHPBZgNC0IP/EV9+IP7LeJHS8XlOJ
Ky115PcJ9Nd+sIYWWCwR18J4B/EpzsQcvZkCYDWwmHTd8QigVmU1NombwMPZJSt9
9VVJX2L9zcLXtr/REB0mck7F4/cSQ7rMfRe70fELYppGTxcthCmIp1noGTPafsRB
PKzdKWdlh1HdzCIfADXZp4SpCcwttj/fJuysMeZiVOpdvQQP9AGGr1grlrKbtoIO
VladLcgGuKAZmV24v7+KKtecmAZaOVDk/JQgRsXnczgyB1z78uLhOZFSiebmyYgy
TXViSn03PhE/fav0pvhaumST9upF2OihtWudXnFpi5gErA4i3IzajBymdPXdXck1
W25MVfRmGuW9cIltJ/IPsR53TXzkPm0X8pSPQYm0BVZEpjjyozmnkm+oFg/vXi1s
CXekzdVKlp72Gp5ubAMlsWzZISILrFwrtFcenS1YSlgu6kAPp/GNoaw3Jq5+Pv7P
m+XXx+GPnmVGUN3IudMcic5TZHnqzTbmwfRJgIufmyYcTC3p7/H/zkm49bp3PPTO
JjBY15DVHWggN6reELtNMZkyMK9CKGsvAlCZrfXeXMVBDjGrLC1jarnRwOppv/5K
NT2Yt8CdF9apoGY5QyZy+uDIOVTnb+Cqh+Kndf49e2mgNp8EFQy+E2RhmrrmG1kB
3fbpUhwb8idUGHqc4vJMbItGGy9lAt9qrIS2CToNLjKtF87vuXMohZHNL0ibZ0Pz
E1/YHS9nZET166Ep6OUGfQYVNvERPPTuxBP+HRTPyUJDmqwvLBFG5ioMvzjxsZ1e
G+mGSvs8Woox79FtqI7dOsyc8V/qn41WgLZQkn2D+F+YoRc4x+uaOlkr986waNSQ
uVWRjXafshKlllDvH2593JSWeoKi4s0a9IktE2/ArVsl72YvmFBSPtwPGDEzQEGM
NtehND2g+njcIBFxlzAujJmxGT5/8OQUMbg1uzM+Ppf5iMlGbFOOKClhPSHv/v77
97A9kspjWzq8+qaCmbPuXC0IzniPGwrzV1sCIl4G/68KudSXWbuSdys0IFcRTzG1
aO7slFey/nsBNk0ZJhM6OLSChYKJ6c7q3hJYCjC0jKoSNDQ0FVE1I9Gsyw1kAZmK
iZoM0mHbKaxlAltIbRoFZY6cE93qFJaEtc4OrHKpFavu2KQDBZ6Mmto7az5oMU84
MtmSZ/MRxhj9ndLsaRHxHbBaVrSpKKob+Av48U9Zh0a6g9dyvqAo7sANTX42Z3cN
7DPg3h1c3uCKfGj4H0jgXIIehY7KetJULETmN+nLD+Sb3b4cs0mwOvkTVrhXQ2tY
9+3qWZdm2fE74Gh6t4VPvyqrfL7whvprW17a+G6KnRxYv9aYGanqvq2KUE048HMg
bk8XOYlFp3BRSfncRgFbeTBDyI8D2qAL/yvcHGD74KL1EmPaxhDWp1I9GGlkcPkm
B+CuSaquxJKoMjiWi3TOeUnNQ0cuJkEfWAe9jaPPjES4u1f7eQFjkQTWpck00St+
bZsCmF9MSpBIOHqzLc0c2jdNfUNoGC1nMsOWt1EVbLDFyafBiM4u3nDX5vs4CmJR
uC93TXisP4yLr9qFtR0LUV+mpbOFJFA4vEGcR13eCYgbSX7oD5iaDn1AIupfeBOa
+JVlUkfXndj7nyzpzn45izmPHqIk5THDZNZQheF2hTtJNwHgOniu2ilr2JJP/7qZ
CS+tqZvy42Kjc4gLdzuvOIkvandOQzEU6YRO8dTEiQhcI5/x0S/VnvbexzFesvyo
hYllbjRMPoIRyB1NX6ekT7zFCKo0WlwiZcGUMNIeKPXzAysT4iS51sgp+qo3HjDn
g2cxfsE+3exfEe/xO9h+zx+AduPPreSyUu/LbY97j6iMa/JjlEKKHAzTzbgBKuwr
3Sbt614FkZgFakL4bjemujLhTFD6FL6agYQWjTMtSijm6j9efZnHLhJ/o+ENJxn9
2y2v945knznLdjbIk47JHV4okpIkfnfhTskFRMqZnE0sKhbdx19VOttzR3V8Hf5U
QzLHPKTNo/nFzCqbseKcHuVTz9j8ngQMHF5hwVOEzup4Z+E0fvo8T/NQ7YVmcJry
rX2RyqoSlUsggWXXbtZK44msrJ/uVGCLOT7Wa6FVmKS/YrI/o2CJx5iAEeVaoY69
337uuxbTny7ssN3k0/+QmyC6Pirvm9453DMQkjw3vPTtdO6nflZ5JQqhBwOrCktl
wgayVlbzge95Edu2HLhrA5y8CV4LGWUxH7Ec1OEiAP7A8UvRnw3O4aeC8qGlzEaN
nQYZUvB+v5F9UXtyxThtm4JdtzCxTBQn1L6BjeesWsnqkduXjev6FjiJYU7ub2eh
OCzpwTkq+9RP8sHTDJFiTeX0fUK7C0TrqF+0qQ6DFIavpZIU9nVeG7tg+ViExfG4
knfoz8RtuHtscw2aXwWkMxmCHYhEyd05alvYzwNYXccvQdph5+g7KKMYJmB41XNl
hSfIJIpWITbwT50rbROahZW+/m4kQ6uhPaUYpFJh4smGIBcsJENkqf6h0wEATCzs
EDJ9DJtkN3xALN31D/ke7CmxVMBEMauTnceTuqhONH7vCFOszS6smWJr938Z5GFV
W7uSuWuLR4eVo+Y0DVPpQZmdVaBqn3UJCg7t8R3jSHtX9n+o3ZjSa21etWxV/asx
DEkkNDhMt6B/sk2/SOJ06l3O9aUX+M3Hw+XCfwn14ikHV3FofHlxIkDz/LtP+ulF
MwZI3JaeMg0k3mnz2buxNSwE01bUjEUHmhnddhgNDooO8hBsmq0pyrjCgiKVCUur
ILKTNjkzw05EAvUdWeDAl6+k4F6ZwP6BCPtaxbTD9HmFoT1mezpoCKxp3ZMqX6x3
YOjDkDkjEsf2oi2cFWaejTxLy6YX6iOaNGWrqTklSxxWiERvr2ehEBdSRXXD2XZg
+iSu9UQ5nO/28xfM9oMf6G+awVymfkPTsj6gsGH5qJJqv/ubhhJjQJ4bYJzurOUZ
s3e954I3MmeOMK6kDf0azd5vtXSLUIgIS2p5qjDnB5sjiZpjtirgTDoW9c+94jYh
AMlMDVZc7l3wuOvpfQ4UH/CG1/6BNnpsDujFc7xq0BE+xTXSUfbxfpVkWeLtbaMl
am/aeZ07EfwDdDfvT+DhWZ22pUg3DU+ZIALUWOW1MlvnEyTu3zi/wP7zmDCRMS8y
YQaGAK50VM8AekIKAMy4tbd4dBxPjv5sNKOqjqg7R32/WlV1p/40uSTEc7gqnlmk
26sPorWz774ihnlkFV6x5UFM98E9PhGTSM6jETkIjmbuZN5DDD2NgY257kLv8J0J
+dI4tp5axFcdLJmSGxWwZ3tgmDHp7iHvrjP/N860LLG+p17IhJhjI5GJls+2pdcG
WabreNymYwj+UD5LidCV9kY86Z1Aiqi0JxFIEBaMXO37HpkCDCmN+NlzC0J249hr
/sRiTeozFm6Hw/G7Gi78QVIdD2xPVESqUXDTU3+HzBWarixytGZ0Tkf1+AnxD04I
CYrPSWVqkD/12PrC8TsG7VqrAaBl3SIOgVvhVImE1r4yqwtfmLrf8FfK7U8JbhL/
o3HH/jtC3iKDzArhPa132av0cVFX3SuDhvEsnnK79+M5gi/kW4zADLEzfKoAWRLA
TUv/tVQoS+LiW4c5a5MjkoJhJ0khaOh87Dzoxy37/v+JKPJOvBKrfAaaSD2ukzaB
F5wBH7Hef5W+TnzecZzW2A1TQxHKp5+LWX3PDMpQVXV0CmDeZHW3Y99ToMg6ThFx
mMQLGfhJTHgclhTsU9636qdoceWaA2bp7qSlhlT3qoYqOacO9UDHW7C4BydIUX4i
hOGIlfzhbINmK4OVXpuxXTkTZ1MD6UdHmzSIJ4zqQPPAzP00ThlXRAwujYJHqRgj
40Fl3Q2fJcsAP1mU6dpBGVzQK3/qmtc5tHPBkJbFbtAei+Dohblv32hcB+IpdQza
SQF/6MXnXlC7Q9UIcHT8Uy/LEJh07JKGfiZ3bLKezYjtwwNlThToGTZMl2AhHRSG
qmFJ/Qnz+Otsv1DkO8LFslQQta4NH6Si5+f59226e1LGeRi2FH9iSVcGnMcTk1Xd
nAWc4LHmiLqzKvD77fmzKDpXFvJJWHOG2tiSL7IUbddSAwaMMwkoUFu1EHBplXom
jWoBfyFFQlfhaWq9AlEMy9+j1lJTBauGkexQ8tbRyuFrDHqVK41kihpksiTdTkq6
NTaY67UcX/z+JvjhuTxEw4coJvTNaa7XQp7Qa6P3awRVKBExC0eSd9ncAosUeweM
u7I6F7BNaXWi5YZnuu9DGbwL0YEKmXpQg6cobG1BCMsAgCwwR9tsM5TG36Md2n21
r2LUEeBrl6CpOiMQZiffuqqD+Gcw3RNfhSjkc9nalaJaVHQQaczCRZEtM+8S8kI0
/TwTHU4paHrvL3LuJvP/WqvKGDeqq6qe//8avct4k327AhskVH98UqfeZPKkzS6m
di238QLj54Ulbjtt56YrOWRm9xHQtYpSvOFSb/yeglBCUjmhyY6b1HaCCXzplyBL
7gYK0a1Hp5FRRFmSDI1VhUfE5v/Em22c1J8XQs058Pfs4+p0GkwgsOCWws43IQjG
g9S4dPuehfV5t8SVT6/R1L4dWW0PPc5T9YdpBKYdpLzN5FpAvUOZcZ8Qdkzim9/t
0/tQlCix/Fefa0WmuvvzOyMZONKTEceFQN8Bj4V/yETHUZWgyWssMbPP1CFGxSQZ
gVe/u+0MXKA9T+FZVbNLeNekSXrnm23bFrgxWgtHS8pxLC5ORa8EeLA1uIDdoIT5
8ykI0KLm/BvgPwkxkY0S9KrYmNqXuWJtwa4i38hYbbsa3vh3kYk0K4lbKTBXb5JV
IZoj9EXDKFtL4yz9H+DAsmtb0o0ZpUeFZEPS3EG2VOEx8S5aJpQVQCyRHrZOpqat
y9G/A7wJvnRt1If1N64nN61qB2yu0VOdAPX4iWG7tB0pW2l0iHZkjZbp8WB3Hx58
T6o8PqiuhFvmdG0lZLyLufTqP+uolxE0mZXKEOaL9s1qQa4swO72maKy10EYaKsb
IDiSLO20aK9r46fYkBumAHCSDDeYdFcxhZdvta5k7lzqA6DsrQGkmwKQDo4BUaOg
uJUxReM/1kB3K+OxpwBtl4VXvIl46hFgYI1xtmTWPebM/Bk6pIarMAHMCIEl0Izu
D0vLJO2zuDj/hzOP2FdGiw6bqjak+o7k2ulVcxsK8UGVtEC7jnSTCwhH+3Fktdov
KrvA/QmllKuRfGZWMwmnnmXvCuI8ooTmdvsi9ZBfz3VAGBpqAcg3ZkFw5T8jgpxV
js6KO0w2z+g+OPclYbAgOguZ8YFTP0srDTlKFBhD7McXvaLokdU/paE/YXYrfVQZ
tx5k1/QDo4sNpxAysqrjvwgjdyNYAcar/8uk2QtDLWTDKSHrDtO2tz+YjtydtOdI
UxKir1geobl5TovFIw7lS/TANlUQGjF8ykcNSDhCvTIDvThpKjguQ3hwX6m9wm7G
Bb+TM+w9BBRVBvIenRtcV03Xj3iG8XnDu/UuZLquxcUl4Z0LefDKgACh4suV2ZL6
EvyzRnwhe+6cLApbxTDQUMEhqjs9T5692sbZ7BGepEfrvgnHWIYy9vBTnJ2PLogL
miWVugLlmXv8ksCJeGHOxDQD8Gj+9OqgjqQMa3jjp0WJQOyDPCSvtLUoL7NFD5+2
8VLI04sJVn1yexnXnSVXg0uRokXMapv9To3G8zuTONdPU2kf1RaFva8kfqU0UnUu
GccogWscZX1FCQtvduMoc97v1YEjzq6KYvAIVp9GmAxknPeQC541BsYV28gOA9/a
MsiSg3/OQ6MZN8NSIyLdvqKA9OSLcn1YAgBP8E0hCk6Rem87l2m+JxlWnjuuTqb9
Fl4YzIVhqIK/wL5MvtN+2OpDtk6feucpZA+/QN3lM6jiMuJxWOQ044Cj0SmSiKT6
eqEktuMThNp43ECYMjzsmFBnGZSAwKU0iwppG5difPKV7xaQbjb+AmarMhrxEeHG
sq4DHDfThLLGr7fFhKUWNYrgkW71v6P0HF/gSDhQfAv+lfrLjYbuTI/POONzJft1
06Klyj4ge4DT5qvYOktc9hFHDr24zkpdO2O6GR1sLp375Th1gvatfX4Po9VQRDQZ
cbRhNL/uaIcVvbQpuWza5RVdU1ESDC6+ThtP3Ivk6tSQpEFY57JdIfllysi/z9Ef
B5kg4X14YF2a6gH0o7+N4ro8mIuUHEv2EUGA4WVdAJ5N4m1mkwE0Q4hVLGPw4psO
Dc1LnvJ5ey+yt7v0EeJVVJVi0NZNHxTZWqTKgmsHx0IBDV23R6UrD2vkyNV/BXPF
MCop8tRaNo8kR0IscG0r01ws4bvfHZV4x288JjVwKJgH9hZUrzebA3/m6GYSjF1A
qNq3AgwkCTONDgoEv6PtWpez3LSdkQazQ/7GV4Lfd+ScJx4NSsOEi9sIVTpdEB5h
mWEXBKbOhLGofBkE+QftCbuGKRnl4gLdjpm/Jr47rMhhlMv2PizxmL4cZmcsNQN3
Z65B2Bj/6ZUg6fRIlCyDUUXKgrsw6PuCxKSV/QI0fSGFSLh+kcqu3aZe2GWnVrYv
BeHEhcU5C6tjsFx0zXS6JkJqJWBC//3Y4MeDeawOS6yLaYvp69sf2b9rR423bRgu
3AkABXHIzEpowzEvDNrinUuSZcX91GK8Gj6cO1/qJ/YBdxiW1l3MQf8v1oQbEUF1
d67UGTFXlJRbOi9sdF45TQ2bG8UJDfHhXaisyQUJ0MPWr2neYrs2FvPPrbrFbDSu
fnmz6Zwm8k1CTFNBkCOQPZAT9CQ6rGQYmWuCZuuOdBRAblTsNWcrRd7LLCg9MkbX
zGwx9cuXteReZVWSAQVN1Kho+7pzoQbOFB8nP2jhJyQg8MgUKUwNCIfxHQa3ooXp
A2X1tLLDhkOiffIVjCU74wgXAr1EjzL2mjWzIvCVAilJB/ALGFja8VIQKyEm5GCa
RC5Zw9mG75gUwQcRHagObQr56nfOyKsFUArRccy5t6zCXln9RnmSkgcH8B5gd0nF
EIKVYMTWgRXjRppvNLTUZ2levDTaL7a6MQwxXuvwQM2nd71ruDpct1s1FqveNUwd
eLzZgjR9nMDmBzRptdJF7QTWtktehMeqyRBT6IlMjkdawp6lZG+Cq9ehA2QEeqix
uZIxTNLNFwPECi2WZBcXuQMW5akhPaWwXESEWqeWNQ+0qb9Ugr12m5x0RLWLRIOM
aqd//CYdSdYT1MUR+Sq4hC2MAUwq5oUz9dxzqDQ3a+xDqeykVaUQcAmem6qMP8zr
sj3fu6Kj+KMtpN2yZKdNGxbA0l+M6ycuWZYsghvj1YgAs5CJ5ojyWIMr6RHKWHhK
m2u2ePyYfy+uiF0JnCRgo+eizxJQzYDiAfC1fC+jkxuCJjuAa7f09QjpLPjVZ1S/
gHjogdzxWxDregMtBTT9q3cLyFdpZA4iuD1sgRxuuW5/4l5gnVp6oYYDKEPY7ETU
qOcSzKST6P7q0CJ98IcbkZXcJ44iJYzpmr+TSo8UIQvPwxnq5p+pJ2yIrhRNyP7i
ewJDaSydtWrM5s7uQ3lwKG3lcyUbJ53x+ucJTmcK/wOjMAoskUnxH7lcpQyhkhvA
28eh+hdJ6QUDDG9oDQOjojcCU1RCBWA0C5OV1TK+uXDTOIWVa8Q3izlWHsF1HXkT
3U95P/NhKf+dBWY2H0kYRFogUyBHYylGOyQavbs5zZzlI8ZgaaLJnvRnMl1wDeCG
YlFt3ZC+n3Hu6o/xgVAeYr+A0nS85xPi8QJft7RYomG2CerFDTz+NEc7Lwgqi3y8
OjuN19A074EiUL7I+S6099JZjKkYObnwDt//CXSOaFax414fd2LnU/FYiWhuSPAc
beA1TXm2ez3zIrGa/3xSgHaeZ/wpF8wyh2Zch+FZwXC40H1MOkIDXIDiAt+HrWrv
0RErO9PGQPW5JPGpxkCvG8WGrz72rheYwFxYvSPi0xaEdzypHq+QQKfJApoe8IsP
FgstfWbmm18/U2RQ2oSM4i8GfF2pOGwvaoMWeibbLX9j77Qb6YegvlbUcm2jiF0l
4i1vfTFEoSqlayCEXQe58QMRKdhrwG/4i33iQ5VPUYb5TRsSQPhhMcdfYg4oiee8
UcqpqBp8zQb+mUMt8z4+mtCj/qmLgNI7VcgGhHjd32Gn05Ll4URHhq6P94OGe1oz
51N/XpS3IsSNmTqDGmn/gIiUqRoqzSqlBcgH5PTg7W9eSX++F7vS2x7SABiqKDBd
4gyjqzEb9qnb5UBm89WLZ2oxKoKs2NiuFJ50YqHl19C/7nvYcs/IhJKlpZWw9AjD
IiPnVRiASwsVBeHkJj140iXcznUnpxmzRrePDDIyrKhy0EkUdP4uF3JX/rijeOor
nIjlaN/pAH5Ux6qq4yXaPG8FXiKzdI8oSlVjCgckmlRI75wCkYnnuhJREaLs6fSA
GRbslh+98Drcpe68npHufRV60HqeurG7XDQAt/qlb3QnQmIbZ4inKYLP7ktGAXxd
KOIvVIgedvggLPO1wDBzuoM5PXz/pQTMDJWiW9XVfAAG+sHlrRZo+L4A7vPvybwo
tIiAKiQou1e1nY561GeRhUJoH+E7KqARqZHaPqGgA1YYFTVt1IJHTUMY+EAm5DxW
yyXij2obhqJ5o1a4Yninh0Krxal5Pv6pYuqsC9M5TV5AydqBYul7Q6bFRXyjD+S5
i6zXUwdLlwF6rA5qSnS5AakarjyfcK88JYtvGQZeu5M8HIcyCUUgmY2uww83q2KM
c8ajWmt8l5Log0xe2Sw8+Xl+CV/TQcvx5xm05KUpP+DXX/6Oy6NV9TFjDThdmbPd
1ehTlI62pZR+Vb5kR0DUdM5y+5drSw1S74ccsTsIbT3N+hhs1sBwgB7VHEqYgYLW
I7LDqD5vUJodwLP7spYTcowbKRlYVLwAeOjLLeWUD2ofTyVS0lFdL/GtxjKrUklq
Oe43ctKdY01xK+Lit3oCN18hgt4QBpdCB6w20Hv4GQBEH7LNRffMe9dhAYpFswIT
jHCF3v+hsrO+KJ4KkSyXz3daLMsPuBOW2KZV8egUjBvEKdVZyBHs1azr5zyon0/M
264KnDy0CwxBgaqw30E70hYuA7jbLvVa1o/HrDB8Zc8EZ/sjW2rfv3j2HRpRzs08
DipaoUJB4kGLa4/hQHLytKk5uzb1XGbzrPAG1i+it+OS/RhMojRRfEPbyHiRMzEb
xBCTnAhtre3rNHvcVKTSxXCkVe7TZDE3g3UKvsLB+44qPNDsD2jcmLWFKlzGo4Ap
M1e9nIJx1ihiLkdElTDyvd3ffDdYJxWdzLsb4d1MFUTihXkdtBmi187UwlIJP1p4
MbOfdK76eptv8N9sYkUyERifJtR1Y3k/YAKh8R/ahpDCKaFQtRt+ShTN0eJXW+lv
NUO4UnxyzoLCkEevb1MECpMIVg+YhqvWU1y3gEhO3sqjCzThijzSaQ6id+qlWFSS
2SZU+XFMShwvmhieP31Iyl3DhUDVE8yGw1lxZTAOirwbXfgC648KS0n+r0rqmHJI
YHCQgMYzquO4Mov+kGNb+MOw8VH8wKri+97+IQ8/GN8E5CLQsMkVeBUCpD6T//5i
11V1qWA8MeMmlcm2DiPm/3+btYs+lpeuz3lFZJOWZTZrrtadLxkKv0MNeQbceHt/
8S6VLuceEsR8f2PYGIZMEMv/uaR4joSEXfMpju+obFYMB7aPpOHNw7tDHnd3vSZq
v8pgnV0oLQTCoxpoGsETCQRfYiN1QyCPnH97vY1qQL5sZaKyCdKTJ39SMA7d6jkg
FpSh2bk2O2AIUYh1AiNlSI6dCEEBKFuWr1QWhEXLuuL6BhsqfSKRvkMOf9DfloLf
XoGhvCNlTraOY+wbqWbdITx3ByfyQaWIdosK6w1jUlLfXHMyfQ44z6tgtLr+EgZ1
BR9F+fGfZNuOMnA/CeKl1/GBsa87M0LMVqnkdox++Fh8c3MuENK4B1BfZV28FrSD
JZrMkFUM/M1yuVaCUaowOq21WuIPJH/E3foJ79d7w4unn/HOi9RTUBcFFnGVX9kI
zwat9ozGAKN+TY5ttmM0R0iUiQ2t76ydBJbYmBNJC90SLCQHE5lmIUg272aFlrDK
3ts5SuvbisTOymtynE/0kRdslSrdekXvvxFhH4DDK2/Ro7sRkWl/6OEW4DKnFtKo
CbnsxUHj+HHGss9OSYUcdySx6PQqCDqsipVBlZxmSV7kcqVNjRWVniwXXvhLdJP8
/8ZDuPHLqEKRI1obOdfqNHkWch0fxbGWML8VhBOtX/qvhBD/hrgvh1aJOJVAnKeK
90XcG26Ca30HXxwRkEoGXkVAMu9GbQ4R9tPaJfIh9EkSZrTRuXlLCE+fsyD6usdb
L6JKUMtdrSZ9lM05Xa8FsExjpp8vtPO/pQFzLBtXXIW7/x1myUlKTWwlG95u1rAQ
3kwVJiOXMVeFGwTG6mVa7q1UlyJ4O5ZI2kUFlHbw/x1HQCEmyynyFEb414G4ad8Z
khIG9lTIstI9egsruLWRPa+KPeKeeHGxTbPtnWBSxlcTVhNRgbsVrFV8I/Ejw2Vw
RfeUP6a/SJTct+64Kzs80NJsZSeWPEmVg4NaGuv2TWttrjVCNiGJ589dS7L+zsFx
JvU3Jc6dTz05AEY2d4QSM206CTwErL4ERMIBQEExvLTO3jQjFuBynBh77rtwoYWb
wvy1QKDDuBVeX2z0OpQPmy25T/uAbsTVe2oiKLyQ0hElojilfHXLgscDtxA/bfUq
khtV/HajIJ76Qz4MBN8NHO2zaohDpT/UcCfUj9thhdvg9VD9dOJV2TS6H0pt1JuD
3l1DP0+IycjzlBNcwXZVw8oD0qyxxhfgAxIyaE1A6Uf4d18fIEsF3MgVY+jpkZuT
mIkX974EAIolVbO7dRkZtY3synr6zaF7VV80oFV3KXyRfvIR0X1x1CVQwstrgK4m
KIHBQZpLYPMZICjTr0jCrTAr0QWte/xMm40Uhf/YnCnbZo+XDJ57YIkRGEy9ZCG/
wYqvy2axMdQVhpU0XC8XR0oQaliJbM3GmUBbtxbUPTJrXfZpF1kyMfN8xkiFp3v8
krD0MycsHub7yyAFok41YHNN+sF7bZzmGMVCQ9KEQ0/Ttx2IiDXl43pczxiszGwq
REkuaqNFd/bYf1ya71jM+OkNevilfcbKc/OT6JVVKQUOmwN9coqtWbUGcZ9wXytv
8MyGp+qm+KHdUmGEilo3c0VPaUHy7xnXai3Wb25vcsjsRkS+1NiKGQfyKamLtjMh
+fq7RBlm8Elc4aC5rJD5ajd/BNw9TGwQaYJA3N7zYGN4mF8Lq+E/I3BcA4NN2gve
B4pX1pWl7pR+L4whh3t0bqGcm0IP8CXof0xcAw16LlsB2rtauSmskSX34x8Wm6Gi
k400Xb5MjjPADrfhJANKVIXO4O80Rnf4mjXQmk66iCw6K14yuY18fHKrrUn9u/hH
+G3/T6cUfHhNBCRBpi/GbIOl/ubZIzDZS+FTGB3Ssa4W2Jvrl50LOzY2cVqgYTPv
qmlE+eGqK9sN2t2+QBHRo+e2APSPqJzbkTtPII1AEcRq42gHejnvKIY4MKEukPgw
dQ4q91l+gWNBWk6gVaKBSFCFeO3usCojN+0+LDIudQxyw4KwwpWY7g2mka70oK03
6GC1IC0bCBYqC7ffX9wuqcyJ7tdNFfXKsadjzsClKwO1Ux6igXdwdxz3aprOLzno
We/bNT6OdPAW7Vm7jfsDe+Qlg7H2FMhUzOkAhOJ52tHMIbecyWcn0ci1wDWP7HRe
EZqaJVS8a/Zk/pkATt3I5ez8WrYAVmENC7idOf82T3xIVpno0NctKOCR1V7QhQZP
G4fv5WqDqKxSvtxvtHnqnGo5/wuEln6U71SoLQKTuPPkV9kZ9p7QGOaP4dumjK4e
+0Kqpwm2FUXYrN2zpT+OunBf2lGtQA5pSxGAIvPdkzwwPZ0+5F1LjNL+fHOLnPJP
8skR45IemihYK8/1rDQlgUrr/O6dHAq6iWk/1JWmuuAZipAHNORqm5CMieSch3MB
sxDoXBQ/PyXLwNLCst+Q/5qSt1Hn4IYKGVwOxRN7Z30clI5KGN+cxB+97CgeUtG+
ApoU6Alhgoc4UL4PE9C8w60ZF6pOTEz4gKcl9cH0l+d2ebzhT9KahujfpDRZXrhU
fSYX2/3NduaZiZIRmpZAUf2Bx1Fj/ID9Yvq/VONS5yPG37FaoLSWfFfNvG08ZfFr
Qb0K5J/wiDTnF4hG/TIVsm2dyF3BTq9v1c7Q8BLR9k6xFjl5+YPDea9YLJ3v5HXP
Y8+ox7ONYsYdaDhTa7cdiu5LD9NOHBI4JzaUxstoV6zM9cQ1adcI0Y17Ev5W6NwQ
LMWvEH3YvrgcRG4NnXVbZz554ktMi+d68OVKvWOapm/9+oS+h/msbKiOILpDwRrA
Uig/h4PeNYaNzUlB3HBOajxSgNDsL3DcX3lsOgucefj8vX1np1kTVjuGjtBF1L37
/ZN32ZxPPTqqyrXnK1FN43Qu/LIctzHtF4Bg94l95qIRxA5x+4BFS6EemH3KJtXE
rZ/x2Q5iXNCekvpc4Wgb70zF9y65rN0XNLv1nF+Y1ChkWC34VklKMmnN6jkQ+gYK
w1xj+hh7Ij58irgNbJ+k2PKsqd245PsCmJfJTVdnTEcQ/JIJaTu1BYZPFN8JwWO9
Q1KlloWJgim+WrLFcfAbSsMo1uPUWLs0UpBuwz+IYY4Gp4ygP8qyuS0WZfMlohid
wyuxqy1TMUoMQT/52oIagFoEqqtnAWo5aO7eQHUEvWNpIBGGKxvNJ4evYGCUYL4q
IFpYLiTFZY8q9mpS11GGdZhkVRCAzI8e8+YCUbVSRY2f3vtB6QUbbmHHpB0Jmm0J
Ls5YTjkrnYZC3a54pK1VHxd4mOPjZuA335n6QP8qhBAavU0ulRe0ZYVBpNxbJ4Sr
gteDXwhYuFrc/71rNaNOB6dr4/D49JFsHScLjPn/sTz3igqvnjur8nVr6glEpy1y
62i/g/y4dP6GcDV69DBDrW4Qzn+SFJjSngr5Ctq9UI/yHlYrpxUXv+OjYHgolf7o
3cCoEZ0eQadJ4itc0aVhNWBlZ5tnYZIkqs/HvVgY7C/Mu7a1XVfyuJkJNi4NqU06
yqvUxbidKCbDQUuArl7R4ZierkMBjrvdmg1yYTNLSzmJpSVyBrum6TnLNYlrk10V
YjG83w+9E9qeuUng1m+BxkPvDqwDcad2bGlpZIzEp9zhozFF9FiZ58A6D3Dwda8Q
NBMPBPrgnWsMrkgIEqgK+2VEtREl+jLKk27wdTFnMUMDtbvvCIAXdzBcFmALMV7a
tLVYANXi3bRqj5so4/FdebrjDKbRNO1g0gMjs7qyKW0e4F6TDsw4Jc8YxrfY/1rw
gzoyw7+bTlv1dpreL546KzHU9HyOgPPwdule28j7xuT7hTfe5LbCO2uuM+UHDnfX
pJkx4wdYQz8ftL0K1kiBQS5WN/+S7Ecpxf9FvtKJtFE084lmKuJQSRSA7Im85gRd
CAVC/GI+v+RvD0Gv4MphOR8gzbu7iyqzS6VXrWIxNM04G5JsJjFgFDn1tJYhkLPP
m6OH46+GsGUK7GpLwqsC/vzdsWcdhsQsi6efmCUjSBlvM0YiKwMiPWGmMPZzhl1v
uFhuGUOlmri7LS2iktY/Tis4KiF8yFjlMu2/6u/A9YK7IUyso3mjUPsydsmF2L5w
NIf4BxsLfpXJaGWnEiru49E7WrlJDJhhdYIwYDZAZmQ2YIJoAF2u67w94dadtp9r
rHPZcsVUgOEkkbiTFu74W1hKwRe25lRPuI6f7H8Sx1NSVArXTmD7I8rPrLtZAym8
rmWK23eZ1djt2yz/KMnd0PdOxAiAugXM+3lOPBjNig6O90HdDWZ5LelhkOiubUjs
DgNm4EHirU3U+I3kXt+u8uJQEFQOYuz1EpbzKn1hcda0hjEGPpN1JS1Ua84NDRnJ
lzDhMWSWdjaNnAPE6/caqOi64Ewzi6brgw4Jd2VvMvQwcuHUTOtzJqNfAaeawW3M
nivh/Vsdzq94UZiCF/V7GWdTfyymzVg2icMmzovhFYGGnUzJKH/zHd0POz03xjf2
ufS5D1/oW72dzI5QCD5pdds8uVUsdhT7FEClmVKmPI3KQHst83AisEPP0SLzUiZK
UXmO540voAaIlPSK3MAS4E7NpSDzA+JL76fZ8LWhG8mP7Na9hJ+pu7aX9cE6ZA5p
e/fbcYZOD9uA5JI9jTitcXI+m5w1p7OZH/YUuMT5nDdxZccGnk1J+tFo8LXE+IQA
37IThO3lZYIxFl0wz7cMOOCXZLKlQOgL7ng+D6xO9ba8mUsPMz8PWDAXR/lTG4mY
QWDpWNwXm+P/Rs1y/DO2q2NVNZnGBJeybC9xLhCDGaw2OSNn5hIszzXgMNj8G3ZT
nuUF2qySGi/rh8GD4iStMFldDioOsWdDa02TAOxGpmxxXiiKfkSJRnZR9QUapWlU
gYoy699GI0wANAV6eqtDOidkUtGzFylMioQWRA6ycazEKpQXYsh0lb1ZNi864khV
cMmCh19ZLo+jYd5B+Ru3eQzmBkJp5i2x7QdAP5Qb9Da2W1A3cFklrO0MRQub6+uF
PCnIWfLIbmhHoWwvcGsFyNsxPrLMnuHeBDDShR20z0yh3ZB+ivvP05eRGP7Ae/M/
EFbXvUsDNO1s0htzCCHSJonVao2Mgv+3Xc69W7wb4fe8Ea5I1HDo6PCu/Z3Ec0Sx
Ia8yT3Rs3tL5KiZsT9QtOXn9mt/kyJkaH4+uf1F0SVwrBqqH1rQ3dAqdIDtWe9dP
GZqdCIzPU8rv0OsrLF+JQEfOy1Qvg6c/7CNEHe1PZ8EReWC6dpvqikMRRY5PUOLN
J7L0oaoAtNyNZqXjrSsyIfh8IMlPpFjzui7ls5AlPsq85mlX8HiA6eIYEm1lUGgx
ral2JUh9R7GSncGiaT5zCsQkTP3CDmfSiXvWaquPy6KNP7Dv9xuV+kqWaZWxbx+N
QYabvtiBWXZfEw7+0RrVJGprlMQVVj3w0VXNOo92vGqEaXGzZOdV30D9WIoAvo/Y
x7uTVI4qz28o+WjQScJE5nUiXydqF93BoEdyk38HXVRY01XZte3csmnljy2Rgp9Q
OWWE4pqxG4xQNV8ECuSqX/WvUlGvc0l+ikbvDlvWeWzahhy8mTiiAbczK/I8nwEL
fnfYsMFYNF2+/z3RTqI67k/MfjPbIB1QJ9BzMzJNkv3Xrcl1wJ4RcUkhkYcDqm/8
XyVYSiGJekA2W0serOSdihYQA68PJYF2w98uZDkifNt+IdxR7llpeueikB+znUV/
O4NXKjbYdQ6yVvv8waG4Ffx3TZKYu1dcEd5xxEeE3vOf/unUk0d2MoXLWHtPpIPi
LVWWpG+guLcb9oa5vmsyCJ0qsqp3/QzHV8dtRurTWgQnaK+ktffB2VxJuMhgUW6T
dRPdrCI1U9cncyEiXgAQjElbxpTfIc/x7lLud0G/OZqdd/XHIpCZweiNWXTmAOIm
4rm9W5vxATEw4phWqBVkyJ2MY52+QydvVjGttH9rTL/xzz11/IFDvXEit/3fNnnU
rG5Xbg6br6yoh1RBgS+V24gDf0tsbj9uTgaG4K8tCyILAsmqmos1PpjHhuXsFtbl
zZ6uI/c2gg3CAzt08Gf3v86eJIARzTNvfB6Ei6x2dnb4os69iUufaZAsdaqlByNB
PL+ph1eq9LS1H9AoGgI2wr9tyV+mw5aQxVm+3wqjunwI6C0HCMcnUz/LHFOvQTst
+zuv/IQY2dG0XSLGwnIfeSdatvQliFCV9r3F5OJDOIqNN8zA0SvINwY3HuZMJ6Td
OEYFIl12R8DcoEhqy0FU984szEiDGD80i9jze+peMF+Kd7Hbhstb40vGzHqDkDkX
GTD//CfQucUDNk13ACL8GEsmixevg8KkDqx81tiC3p8jyDYEnQe/PK6amYkVnWWM
xdLWB3kL3M2ECoEleqbOv8OAiF2DRPnDBpJnvozVkREgX9Rh2RjuMuGljBCf7myu
CFFyfXm9HNnQkFXMf8EEdEGpgtOm5zZs9juw0j5e7O3zaXrkIjYAZbCUq8Ipz7uz
Zx6GbtvhrILML9HYyK9cQ5Lpgz8V8Les6V7JWSjVGM6P6JYC0cnP9456HYBftY1D
pU6c24Nt9gsyAQhvZsnb3E0a5HRmlN8VvsAXsOwlySwoea/yhYyL1C3ImsJm2oMj
/BIS2z1PSQ4YuqL+K/uRFJ2mZuXpYrDISIle5C2oOLX7WVeT5pp/0vIQWQ8kBqEy
jCLz2/Aysuk6qmYEjvnEpUGvgEYTolq43VWhnppy0iNzh9IXq78IphA9Mgi3DmVY
TaVm/AxW+uDzGzG13vjBACFr93TOaO5wqeOO3h75DjQ67bXnCWd/wgarENYx40Rv
0H0KYrHUbOeLkXc9Iy+BIycjtB35Ev8lMs8ypLOXh+Ygk42kqHiTBqUGK8uqjivR
7xGtl4yw77O7LDSIqR0yiYCLzsUIBfS7SMb6ua+aLabqESUS5oZha0lVHWx59J4J
VIFESkHuNc6Pagt7O8g0JOLB5pQQQ5GuT8W/CdqYVRdkPVO5Fzjziu2bP7wk5Jdq
TLD/dez5cM3NuXTQTDumH06ROOViY5MCCt9C7qkAfulRONHM+v79M/V/aGTPEGJI
skyRqFkpo3qpe1YGoFbEn/RFQ0BWva+RSUUBoG96B40aemfEXzW5o51WXgWnxVTp
gjuWn2gCjy7y/scOVG6X1hCD9QCCgaGMumjcB5ID8WFD+XJ1ysAwyqKNVElmK7y8
YbxiWGwaEnggdAdYTHZDChWnozFaPnO1uD89OTNy+63xsgqMfXwJ6wvu5Pt67mRl
XfevrqwVf5d7M942N1jSCh6k+028KiFRGK8jZ649kYP0/b51+lDrMW6/zxn059WJ
aYQs3Bs1Pv1xpxWNHr2x7HMV5n4ZmlNW0l2LD20n7FMyVSD+34IQm8kXeaoHIY4k
k53I7e6FjD+SFE2e7sX11Mrsr8ra16mv3xkpSFrUYEW3dOnKEzJVwTDFUiDEVBn5
GmsSZvXVzy2yrxVL8Tal4t3e7B1hPvLeziETeGmvY5TBiehtrje2aL0JIaEdF10U
rU8x9+0Agdyy1itf2MDvdBZNk3zs6Yf/eAI2BPmVeKiCU2DQjPZbkYBHFAuk1xUs
tJ3iI9/Syg6lkte4cJAqmnh0flixE1hYwY+at4PQexJIYQKqh55gB44wWHnhNdZx
7aUzevPwe5erlcSSh+OgZ+1Na4q/QiHEAUG7gTOIFkqEdGfx4LStzmC0wpxEbnzj
yXpbRYM9N8zeSMIH7K+5bSQvz5Bd2OWRGHGliqYwjXjf1l2u1zHWO4h+BvipDS8f
OCEHNkrlS2p4pcRcsfcx/BbN2n0RkeXCsk+msA7Xs/Tysx/ngLrFJoytnwF+yWiS
KFA0SrxOIwdW1MHRzD8uk0fsk1itD+5Mp5nR9DekayGF5YBAmlyffv4oaIbyw1Gb
xI3QsWIagNTzGKOe7n65IZvMOVSN2yTQOiTYZUvia4CEUAb4DPnhxWUq+OyG51/d
S3o2xI0sb4xKJQf2ZPH3kiv+w9zMgNg2ZhPp0FY+QVAq17LSfNezIMfxFeknsab/
Se9gVjaqw85bWvlCejtXXRNtQ/eaih1dHMrL/XMec1newG06r/QtBPvW2Xk0jaRG
r8H2f8Zuo64RjAsn+zjOEPnKnOCFy5CiIwpOkj17xV0lMZQA3L09ABHMhdCS5kCE
EjHivpuuCrTh2WHA4cAx+Y4skrTT3QT2Tj1QQDbytUBXjKIQj+NW+fezqI+Wbr/a
ZLLKE9Td3wp0yQGD35whYmhphhvbDLhFELJ8MrIuJC2Ky1tBRWn8+mV4ECRtdjrB
QTj8G3Ux4uLPVYYKu4NLBoDrzQz7Ds9xIKXPJsMj90aJrLdAddj2DhqTPMIiEzKr
V0FtCAaL/Lg6Q1ovy1+1uiqwlHKUG4OMYHRjZeWXgUqiSts/w869g0STJ1jDsvuL
6+k21kf6RoLMFYJT/48d4vT7PDp3fM1oxSJ4G9nvozc/e24tNnCYq/sHIHmwB67X
v7GMu+4iivKKFQ+3FU7FHwmrw/j3V77uu4nG2oZ0Je8ylyhOvIeA2utDhOT3q5Gd
5J9X8Osnc+eEIGcLG8BqIOGxOgMUuvhV3Z1M9XwZx4HI7a9diBQ/ICUsC3+O03jI
vbiIGoTPtNWfikvT7uYpUEyfPHudgEibm3GzM9au8GPgdcNdG/qGgEBbZKLAguGl
W/aGuRkyeL44c0GpbNVlFZXg4I6gklBnf33XUyouOD4j+8mO1cutoTqPTZi+/TQH
gwqbDHb2OqQFGa0g2fRzL5cYPsi3UIKri28P9et/MFB3/8S7wkTFViNvTWgKdxr7
OlsY0G1d0iENE3ePTDKKkPnsFYP0LLYVTAgt9FJhW7vz/x45Tscl1B/PZYpgvYOo
tjscrzJ409qu4LSuWfz3pUvliDFXBKt/xmRusuPnxaahKKtNHqbtu63s1dvyvEfY
2PFPJzsRvPCaUEFcFIdY0wzaa5u+prjKpph4iUXDRSpsi8W+wQ6EaTcdMeOtYfAP
FGQEgjwPo2w1WzUD4ajDAaQSumAFO68dOKuyy+Z4YyIza8xYT8RweIXqCebzhuWL
jWEfKlQbdrjMI+0PwV2uMamtg4TwAAPQ3d1RGXCLf5niBPfCb0LMDuEUtRYNXmj+
HrNtowMIXGxqm3riYgTGnJ9Vl//0cYSDkre8pdX9Jvcj0VdFYUJd8RgM2ePF1M3p
fl7ub0OQz2zRGpdC9Udw9MZMOKsAP7gg7NbFfv2H70/GkDju4SjhkogSd0TAVsjB
qHCWwTFfIRL0jW+OFM26DRF1tUYeZAX1LUM6untwD7jBFoxeVFlMaM9g/AJIBO1o
h0DzJUttl9FJH4vb2rxn/1xSinsnmqBP3j8KtK4ML1GM8aicT2CwiQosRJ4gurGQ
Y2EongGdziA7N9FWTORFgFvu3WbxS+UBjFuGLtwNTJGQKFYh58VB/hohZFY1ZpCU
PjqxhX98JS9+JeYnALtBr2zdOUnz2nMTRFLOaPowAB9BvGgChN2WGpiPti2XztCI
rlGNAFmwskCgjdJSlgK07L7drqlN1jt2gHuHcA1NNTGP2ae4b6/khO1OdPuT0MmQ
Kb2YHrW2vvIoLn/Pn8HHdI12Tsmb/7Qa78MvslQtaBs75a6Yv5qimnwtbqGoTbOn
hoScZdQfOFQo71M81nkD1ryWEEW0OmYo1BEvYD9L/Qch3bR7cgvypaNYxiDNgElu
ofEGZUZM+evYSAex3uVxU20dHEkuJ2y52OZ9X/FHiKXbBEmbRfOidnPUNX2RxJda
sZ1/U88XQM24ZLjHY++qsdlhHzNKXOF7e2jPSOVd28amoIRMGu83oeRQyCjz1Hm9
QticOJ+ux3/pky7eekbCij45wao4tbZLRg8lvNViqlpM+Hs5khEC7S98G8zmZHu3
dIzG6vO6X3dxfMoOeB0BMg8fbgUaiq5+LHWqmV5BSlBLxWCNzOSdqPO+vbC37sNy
NdJnT6wxr2jYqDUl5WBkZAO52RrqWabm67na2+Gni9/bnK3jbkIIKfcMUuF0guUL
u9CCWm/KVf6HqEHWvtGxofN9+wAp+PtlDn6ysMZlXDQxO1eXM3/LJ2z0e8SLpKcL
F+LRpIk+HPTS4DWpqPajv7anlIiPVOS8Ov5JOdOVNJczFep3lYHrHs24EpCt2GYF
eG3eKW9LlWr+ZqHkoN1xxlVM8Au46bMnK0k8kdsaC2oUfpV8SSbvL529y/8yd4WX
fOciAJxTylzfKCyIX68t1N/+ZXd0IFaX5zso7aSFmT6+QUX5LaHa2JITKQ8XuoNK
iyj85nKXRLJuCakskq4LWQvorH/9qIPFgNODsUFn2rkvFu8PUdCsEoYydpV78G+X
fEB2BKzDdqJUx3oOf9xVlXeRkUt9rqvfrHnsRj7DnbqGDzBjRgFkDzcP5gjlnhG8
sbSWZbYCw8JAsM8JH2ukmASofMaeunW2jjtYu7CItHP5v3iIvxVg+XnAZM9cLt+M
SggY/rNJNqDQVxcGYcXlVBN2vEAW5aro4nraTV+zxPJaH6yIU+kdwJVydzzhnDOi
dYopf8FhwI4/JU6zvLoBxZbJve6ezt0zS/J+RSxyljEZBbRYl3wXUi3aTkbRpt0I
z5BMvutACtOmOOk8qYXTyFDUtrA5Sm+XAA/uO0+7pEZn7jI+svTC8T2WmVz4H7Ct
E8ZoC5TxgQF1BD60kpW2looGYh/2tP1w+qIwVk6KdPU4o/armZetL/QsEa1UU4yX
nAPX0l5Pmtp5N5Sd6YAbcaTEZ5FYT3u6l2IAHCX1zTcY0O718ILt0tVFxzlUNTkb
Tbuk9EIoe2V5iGEGA7rdlIhJwQRepr6iqHmIYB2EY8v8NO5mE/QeZTOX6z5sN5CZ
dSB0eliYnOtJdh/2tI89QrqtpGkvNJvaUaHyKNrHQBJNjgu6Be4CzXKGpHitvfSJ
lp8d3DIbyGssA3v9Lno2sGsLCxPDEV1Z1t8Li+hooyw2Lwo5p4SAy6J9qELJ/QgU
W5K8SEJgjj60ZydgETVhxPzA/3uCpcx0FBdWPTr/lQJA1iTkxl9zZzgykM9yrXyp
RVYH8hV2SIjkVUwpn2Cr6b9G3kNAbv+uvE2s0oi3YKrfJFuidiGhxMM+ggZEaV+2
WNXlhDjgsF8eXuPYE+5JPWbLrZvidlwNmt+TYDk5ZlY7oZD4jlum0j9xoLzXgUqB
eAwy0JWWyk4rJRA84q2/Obe0xH5oX5VpDAA43RBDLHCCRf8OYX7b5VClf+GdCr1X
A+p/PxKoyxo1XUXzW92mKJmxf/gqT1R5Hob6nukVLOhJCae9oHtV/PAmWDC2iHw4
pptLougUcPqVQxvwbSNeOOSbZUMFK7yMbE1/aFPGq6UGyFxECmOsuxoZeIO4SCv2
JNGtZTfwtfr+Pf+dSz+U6dH/YvmmVFrEC//0XsNCk0eYDvIqbTlFzefEVNFOS+LX
ev+mXJlGnaAdDSGIrrmYZK1fd9whl7ga5GKUdlPZe7/bNue9CntLdfUz6aDM0ayv
SkyjTAC68b88iBX5MrXEGiLu93Qc1I43j45r9mbSDlXDAxYjglAJh78HLXJcWIYe
K+raIngBQf1Utbfwjmt6yWPFgx8FzIUTDOuk8bBU1qkiBLdmh+bBLg0IHmDRHnVi
SboRW4oVSTtTntsw8LuRVKOEX3oCaVvcOfEVJSm8PMMo9K1tu+7xbgiKdWRDoKxQ
AF2FWwBulDUgYASD90lr1yQ/JwHwYwssdqZnHZCTRK7PmOtGxJrlP99kX9U/BxSq
xwgT19vGeQ1nZiKRCeNRDt0ybvfJHoD/6jmNfQ9xXy0Ey6DnVESwDwIQv/d4lAWh
TiR3zz2WadMj/B8C/SMATsG1U1p8jxksc7uiMlDxRulbWWKEa7+EbfgykoD/P1/s
9zH3yXp1Tim07B0Y/IyGpUVSgDF9wzFM7OceTX4gpybs13CuTnsSBoAvxsP3sULr
RBOmsQXD7jjn7hWoLN3aQWBSmyB5em/WmRQMkLq48Rn93aHPw/8Tik9B90tQPaYS
rjSq2GCwERqBCOHv72QXm1HqZ7ZS5UOCPWa5IqlF/U2MesVbaoNGtmBVTEm5N2KR
RI/Wc7M7z2JyQLv6heTnwDq2ZoK+GtwP+wcTja0kA+5Slz4rCnPrZ4ayDJpa4A5G
iPqJUG1fI33PCyBCYbmODBxMx+1yVQFfnM+c5StoNa0Je9fgD1dTdGgzuhKdMkoh
LaN7grcnsoe21+vbDByaFg/OKlqj812EwhyyXGSyBlMyWpn0odPQOnfdBF7/pPFx
1xXQpO02nt5IpXP62t01TDiqRlZdxlHmIaiDZp0mxe21gRdZ2Uwf8BCU3IF20mwV
QKln+D2Ob4jVzjO8S5lE/hIhQFmx8A9Mkx1RsOcOx8JuyKRwtphPNyDCWt6G79sB
Ca4r19Emo43iDs5Hm9390OHHub7ktRaNt3+EXQ3DahNQ/jizVfkGSHwyrdHKskYS
UanSKEuoBv7YYD/rjMrm0Q+/b8XPZ+BBtNa6qBzwAY6pptpIV/x2dXW6ZSYuRiCH
o7lf9ADjsjrHaZHTEAaPaLpSjzNivbzx7C82ZlHhjD3ZlfvJBoRlY7fR+8lbve3S
N5nDqq5POGilB7YrGo2L62I4jc3TIY/DuXJ/qF/7sWBE0up0Xo15za8e4G5s36ZB
kwtKZrnHRm3CKHqnukit6t17fWTSePJRVQPp0eSM9ycL/1S3MCM+u3kQ8CGCJSjP
NMXLHvq506txRXlkxCfiDwCktAssoKeLqQPqKHDsqh/qOo5mkkhKU/eIsXJ6XuPu
U5kJVTa8EBUnZunJzq0jW4IGcXcvgXp4utQzO9PQqqcApUHGIC58dF1+buFgicsg
Onlnjy8FKindjU8yVk6txKGmuPiUSqxIKoLY6AJh1HUOv7d0O6LpolcZMKBg1Uav
Y+KMUeu5m+c9pEPkwgR9qNtbp+H/HU+UKdN24+7twO7oZNnxM1seYzMg5/elJdAy
kdYqexa1gqNEC5SWRfATxGRftDbZtr5BGcaYhwHj/SsvxdexDARdLrusbgKiG0yX
X6Uv1IGbR722mdEE20iNzkWeZY1bMItfSD1i6OsoZE54WCh2SVmoqreH4z28z949
Ti6DkCfByw/RVfa9frLPEYxAcq16cP3aYIID44b1pstjmuLp+KCB/h/kOFk3jy5G
8HQIOZkgSOeyAni1qCa600O3GtiuUfZUheh4E2OiIsdt9iqHDkO4VlSVfHTjpjFp
no5A7yBIRVgJU8pND4oMPTjmB9e7rOpoH2WJ45cO4nWluHmUNx6uO+l//bjXsCb+
GHBHiRueRs6Ae0g7gc6UnMvSoYq573tuQK53wvbdZZMUVpzGZ1J8vzYo0vlNGPB+
Q1PKuln/utgIuCnIMlTvd1NLuwAJhR9lTsozGH9UYSdhhgkyv3Db5hc2/NXzshUu
XYIdCaYS4igzGH7mK7pu4uCMqdg94sTob3m1lJF8C0dzcNb7iwJLynFWe4AxPvOp
8IPdPMujczs+Fq6bAOjRBgiH5b6dffYYMXJ16Kof1u9prHO+uKyAhWwaB+WTNFw3
Vd1DsnI6wfxPSiaC2KgMV733tYsfXMExlcLYjJu0bKMckosCZzlniUFPOcFKCl/v
yV3YQrXAa53b8e4NglxifCjaPAsd9tNUqF6FODmbeudkAKbJwFbhoI9hzgPt5L8s
VKQnSo2pAfO36RBm3Ks7y1hHwsptpkPOW+jKQkYtl0EScdYX0jI78nVY61cc/eWB
Ipy7adDryecJ+Pv5d0CHHIu+cdbXN9E2mWMezxgqb0rfinQW506T0KERShmhnuYM
gn2DiMo0Hi/wI/2UIkWxCZAO+86RgJ2JmWCQG2MtJTtPfVsGtxh5TX+i3OLMM7WH
NwD2ZZdEs2xI6Av9ZGu9E0SMrlRUvL1I9f3i7nATyXhJ21N06PJRsyKXE+XrumXR
m+bmMyVBjfMDOnQhoQTu15DEOL4/8IzjtD90RFiCzZgMmp4k4PgUNSlIKMQZOqFw
AcGQ1CiJm2GC0hDppr8zUYMhsLHKWHjGJx8XTVUq4r2+94NKIyhPQ8fXzsfd3SP8
wseY6BWSXovr7+0axvxD76Y4nrMNQVe9OK1FgPcnd6bifEjj6RU0Q7WOLGLFHA/j
d7TmK9GIb0xgtG/jj2DOmwV3qvcCK2xjUBPh4xTv9LKZeaiUn7/z1TO7o/YwJWYn
4J1gn/bKDdFtUMnksaBCtM24opWy48GPk4i4zSoKy9qfGzN4UKi8ciiJgODYU4SQ
t8+WFUwPh3g7e2qI/vyZgUB39xpCSdq6LQllHHJMO2NpGJfBagSme5qCqoB4XHk1
Fx6D4mM4YgCJs/IGc4M71q9PmMkPmjkyOAuox1uFK5/laaRonwQYWT+dWg/CG1Lq
DoXutlOtkLUb2BLMFwxmcvIpw7wdP3tct73YUe99BeyK5e7sfivx8aM1KOCnVFFo
8LnFCGrmnkWizocAm3IS8ytg1WDLaYN/IHdOLUPrlk9vltsM7t1K1sClP5DLrkOg
cB0QryYh6hGi8W1zWQXQKnZA5DaWBwqj3UVGsgFaXDJjre8FHxyy3lie/lHr1X/2
DSUXwP9PBEIPwypksJ6TqLgndOL/GMu4zQjk8KFG2OrG2ND+tXkiYIsr8Ot/SuH9
lFttKXK/SKjtbITgVWzmPdI07o1fx5Td8HegZsuHG5yqjmFFzVtUj36zDdk/uq6/
zzySt59NY32Sxmc1jGyi7rUDwAELmURX8hLaGr7jPENxgP/6vbi7nJL9tolCiUeH
GOYZ2vnEx+k6VXuwt1FFNiUlkDPbMlHeRuK5ccvV1fvj7u/yf76IQTNV4IayLIv1
h8Z2v/xRJcCoaQvNM/13j+DDDQXKGlDBiQ7IqP7uujC7tIBoe/BO4Qf29cgM+FZ7
HJ76Ik3UOYSZ96m7Yjvgrp/VtDIk0BD1mcubrVyKRkaavpWpy717Ip8Q+h0WfMgZ
HFG8G1746+/3Riqf9W1fgF5ymwKISH1UmF0l+EcQQcAQN8vDqQJXul89PsoNsocb
r9DOns+5r5X4aqxZVabwf9BB3XT1F8mn4DV/0fHW+RfTP62AFWhvXscQkdnYiT4s
LjRQRjsFVmBWP+LAZfnT1T/WZ9KJhp/SZ5fBBIeo90A91K10kEIoZRdbv/fO9+GM
vPd7MBIoqqNytRC6JCXEMX1LG6AmnEWhO7qJyo7a0Qwfjxl3G9OIDJBmYkbwnw0o
Kigv5IGv1aFYHj+v1HKuQ6npQhzrTpwnZEXWZpBes9KHA8RM+yALp2ib7pJ03yvA
j5dWkCr257I09XOiGogwnnsOj1QT9UE88Qb5V81W+gdi1Lgy6Na6gFUi5OTF9jse
hbx/jNj9OnygobNWKjZlS9KMP+YcKMEMZ+l0VlGcjyqMxMTlpO9zQ226I9LPwRwU
QL3s5Z5EnvRWgk7LYK5wpuOZE5WRn8xqDb3M28TPAk++3YranMLKeTq2UI/4kK6Y
FhnUpg17H3tL03cePoQ9v0wiZWEaZYdocl3frcZFJL6WY28el+o6PwmOBcoEmSJl
HwevZw3oqIDAOMK1VsfqgVcbguX/8FdWG4QoGmSI1HEdbVPZJ5DIs+a1i2hyz67k
QSGOwxOz8tRQtT9qlOdaH1F12535t4e3YHr//xQjGo2xzWJD5Y80wdzEgfKkiBiG
NotoOOCsis8iHEoIobnFs3onQXJ6Byn2gVjFZl92/tZ+LldaHsK0j4B7zrwISf1O
UxuFZlDZCD7/O5PmU+FBYfgcWJNAaNOpFp6D4CnSKrOHlMyofQXZfPx0JYVzHUTX
JoLKdprjdW+O3aK3NE/BvvPNTgghP7HTBHDWBvZrurHF0sZvte4e4kA4GO+kK1zu
ZzKh6t2xQlUFlH6b4U1Xd2gX1GHeYrFh2etH/FLand//DZPTZfjBAYe5iA+XAQxT
X89FTgiFXYHwCTqpUu3zaxo33LjEWTkEx3YdTvAv2kZR1bNSr4AeWK2CZkaz/QjM
oofFnQcDgaz1kGI0KaH/ZVemTx+yPY+0aGeHTmVFEmx87i4SLg11A6P/tC0r9ZWQ
hoyhQzRNgqW4JuqUUriyfVw6g4jhp+q4j/hh+1+v4QP2+Fyl1BtQhLAuUw4iUPTb
o8xQSUKtWRBwzVXyFKvXUbrudJV2dsCGTMJcbdLcfzXJRiXatPSQXtWcQz1GDxoi
tIcj4f0hO1uo0M7JH4UPTjRzzzEqluonZxxx8f/jhHfUhErXnry1FgfV1o8hX3xK
sDgX4tpdEyUbpyoL9okzCSWPUOcqutFqCeEjzi4esaS4f3hD4wgoBghWA0hHAxf1
ERuLWAN9FLRDJZgF0Sv/Kmiy84VaBK1DEeqVGGZue00IeY0Y577OhkMFWzn11F7P
URp/pV8xu/fRKEFT64a9+eJhN/7+/h5sC8/JH6p8eiKVyBMm6SqjHLalvz+5FMZ5
R0QzKhWyKzs06H4HS2k0GTzZtxUhT7zC0R7rxzMyynzSz+hOt+xdxw+y0J9/x+EJ
kGnFsk5DkKBr0AiOVjJoP+1gMrZQJ8tp3qSPMMkUvXBq1cWb3PhrNOsRRGHWIo4F
ekZr7EaPZC9IpHrbUGz8ajmSzjWACWHvQz/2AeDCTCGVZPaKVb9/RPDZnk1p/rLc
8uC5FKpGIUpo4VTssPvr2+oC5bbfziZoD/PFHGsFnaJhSEU9i8VWM9GlOFdZqjWS
SXWNMKLSWCqcCGGKmx/0AjE3J6pWz1VEdOOxzsOJ2ymhSCVNMmbLcPkQxUMqKiUU
5U8cUT+8Xkdk6ZH5tO8W2SxPG8VPKbPSZGbdnKa98WLLCH0qk0vm85v1wtKKlF3m
mvYs7dDiE+Ac3MHg4bMMk5h69WmCAjtNAfGT5EVHYeVDCHlI4kGTVlb1WqYfvhEw
0JWJ4vhgwVgP+hD8U7ftbm2BI7Aazg6LfTVcKVje8geN4dlgOxega9JXgi2dL87+
Su5pbmv87KSvfCNdYDQGaFp/opHkm6dLvlAPFsTleB2OnFuhn56oJ8G57bcxzK/E
ECVGGBTuu7++vtmW5TF8EA2UDyw2Lwf6Z4sPNwulD8pkvSAgelqHFxjGr2vB8AA4
Fuy/w0XigxqKNg51u/ZyfrNAxCVW6cbCtI7f7xXbPWxZ0zEu7Kw05GqoaF31ipsq
pobIdI2JRz+jJ4bTAeXsUxOi+8h6oyVZcq16iIU/h4ckHFpK5JRfB6B/NTPfMAO6
4Mx1aSFs6TEOImdVoDcqTNwKQ/1CbMotC+6GWWIIctCG2km6zwcy5FKBtvOb9vIs
atXOaNqoINzZLXwKF4mKZT4/FkKdt1A7O0a1AJ1+SC0elC6Pak123EgJMinYI6On
nre5Wu7/10vTXWVzq4xMk4jzqG0JSIHi6V3xHTmGttkakoZ5tyTouQYPuQ7YOQL5
4nqsIGGFbxCw7rVY4+GRig0JXLKUXtmxLmbm4ZpxzqKmV0syYx6ZkH6qaFVF8I1s
kQon978vyiy4Rq1MHNDvjjXn/k75GrXwNcjSLpU5WAB9LBxtM4E9vkITIopnLZvh
DRSVNgue0ELirBTbLU5W6NX4xGzuDnR/8Fo3qgLhFrzwNqPgmnCh3sjGz4Ga5emm
X9TqaRAiRGYzC7HyeAFanJYDwUu+l4d+KtgBCrYFVegrCvByP1LSljv3nEsXiEhK
EzFy95hOZSXE2PSgwhfMAC5/hm2HWgVzeFwzOFcUTvXyCha1o+paHsTtwNBlHesg
cn/DyOyWwvr4htKQuTjJR1k4kq3W19QLXAxdWbVSWcGud/0lWlvHJ6KDyI+3KHQw
3sw95Dy3U/uOzuhOQb+4k/By1bkKHVubrpvIWEgZf8z2z1Z9373qrXQIYOHTFCgv
b5QNL8qwqifmCr36dxYI8ne3m8FU8iekTLEy8jea/DG4Nu/AclCa+SP+w0nqomvZ
Gd1CnBionn/eAXZqNhXmXVT/ZC0CF+WWQmVRq4sFuyM59H5BHnJ9fb9jK7FmpUuZ
3Wkh4BqLIWwF2sEGyW9Psp5+lFn0GKmRzkBkrvg8eA8ShgrkuFKixkWc70GQMzeA
P82iFpms1rU3K2AyO3BO7Pdj6OUT05Odo1IgKAPoAx+S5B6fA/WKJaMp4NopjEDe
c7PYX03yPxNX8EYRCVEMrCCDFq64VAWks4BY04ECfI/Pqd99fd6eUcDHjwXpy9LP
xMAv2UT0Joz3bSD6QuRfA3l42IOdfzTKq4hidMOQg0Fwzy0D7T7ENg6bKccj31Zb
9TTcZlLlagQs/YyBZ3aHIux23U2bQwYqCNPBHKwpeyFvGQhg0fHxaK70aPYWf6ZP
GJsv1/ZrT5TbBglwnDV/OCAodmQQ5Tx7UrOyw0MjL8kt7g5Q7qy0iMDKYntqdlSQ
ZCD76YTCixo/vIep0JAdySHn+rN0Zmw9BU4jH+3x9bdwUHpOESNwrs6cMK78CD6f
SHIhXfgWATk93kNw3bx7vRbfm0PYElXr+ccCiczmY76o03RoDlNJ/4KifiRq09JF
dfAkHmHQNluvRS1rsN/XhY/mvJU8isrPVaU1i1YEJLL3T0VgddbPssyx4yLV9ixo
+etsUf5bNTYPDpyeycGVxbsQqr/69g+7NWr83HcJoSi0CO/sLLW8KKyN0+VZplOa
tgG+knKDiS+2mUnv6PXMZtFct728y0aHPyZvZjgWsRoBC4ft2iP9+/o8/SrPmT72
HjE/KK54ku+SG09zOfFGFnXCTYXwF2XlJ66hGzHzRZy/puJ5gXOxcEMBG9ER8Q5c
aJly3gelG+hneQYcUc6khIrIBryNpELLdz6TwXLp2OL0Cc65DXSTsrjDfsWLPL3/
OSXt6HB++BWlGcTl/Y0CGjysbdBZCRVdbUCxfPejZ6ncak38Vhjf/mFXNvuDOdfP
2HAgspR6hn9Y+1Heg3da+VGVqunAu5wWqXwtfKSqpSUmzsSsfwry8UCScJTNXyub
P1CV8mVtixed/Kj4t+8eb6XNSUo98A/Q+wBg34Pru/V58HuTgXlZ5Fu68lfK/FXh
V7Z2ynAJDD0iyJsdLTsZvlJ/EEMiSQlNOV5igcvDoQ/NANXM9InvqJfq0jEQ70Zl
2w42n0tOAm6DTaLg/hiJWKEnZSon+lkGCF3XZh8r+TAoxx0d2Bydor7D4sX/lyVg
iFUMPqgIy34DXBbQrX0Bz8e3NhAj5r3+qOl2zE70+Mr3gjz+T+OHIeUu/3jx+KYm
h2M80Ook441Gm55uwACIdBC1XJWetjydZXc1JP/XNEoHDFzbok1Z+a9NUWPDnCeT
iHVDuy0k0ukGd1XSDYMyd9fpaqjR+qfoU5gg2VnuL1rC5Q6izE79VfhMbhX++xlE
lcsBa37nGE2SJVdO3wnVAIgROt4P+qyeP8jSz94FR0kd9Mmah2QgLRqgVJSiLqnp
C7lwwDdlTQrgll2u1azvxmTg3uWar+OKledjl72RNYfLvjaeNEx679+3+QUg4sRh
jOockXXvUZD/DhKGYlS/1WI9gqLD8Zv6ksRndwmI/5jxquz6613uO4+uBngQtsUS
/ct5ePCPyjYhSg5wojKXrFClLvPVPLkQsQ8ijchQkxVbJK8tVrgEpXm9p3kurXXt
Bb2ZnbtOmYQ1hERiNvH5VPmCuGkdMmIYBGIRrttLfAe4puphLyPnsMbhqZh+SNzA
w+hC7hCVipM+YMkkB5147A2SM8swpQXHL2gG990Dd9X0dNMb3xCagrg/u2CQlHxY
Qus2aai8xATByuWutLONn/RQmfJHE83x2bquFpLhLMhlBzpKnVjGVsyGziBMjgYa
EYOYPe0rzh4sYdgqui2YdDFLaoC4GzfLyllPKimQ2DN06bzxVCwC7tF0iEI1y2Vj
5z7/ELhtn3cXx7sdXUzsX8IQ11AdbPu7pYiDxGJhB3Klv3F7hysx/DkdyKgcdAsA
Ucl16Sx2/mjdBbR8vVnfiqFLQfFTpc4nMExM08Du3S7JXegcD/x/y8mgWMa/yehc
zDl2vHO8bb0HMWMjG7M9xJUuETqPUPWHseyDi8MXId+oZXLhy6AAD2gEwiOpHygY
9GkZZ1Dm4r3FUFAt0ndFbQYIbxXNEQ59F+fUmqud+WQ7ZqxhNJbIyGXcIUQpvieZ
KZjSgcs1qrtRYyy3DHayDwDz0tweFwN2ABbXhUB0GC4xXHJtZr44/j161QSdCtKj
2C7GJSH/OCIPCT9pGtKS/YZwPkk+wLp4jZ3MaMnTU4cc2kLaykvPdU982dGBMRJ6
+pbXL8yCWb33DKqTDWivj4MJC9l7U8KrIuhNCNeniS+T3ZVsVQDG6L53bqRcxlfL
rtpJz3sNEgmSuKtQYljZ3IOVjG/238JBmtcbLc++azk7NhP8WsWcFTb9Y3Q9FBlh
qXVUf54HnS333//oc0fPYBbwNANshR5y/l2TgbqbdnSmVePqvfG4f6EYYrDC8UW1
ylhDNTOGmTyO1R4mySoyPZbb+4GluPwaGYNVoDe7BRwd+oqm2MpsETMS4wBifXKd
AuXIOKeDfnp3xFnFowd374Ci0ly2kV3KeleCyAR6ZcRj7zEOGB6EXVD+fIxn81RZ
ipNj2L8CghHuitituSCpCzsxmzxxCeN2h1LjYrLWRskSYFzoXh1M0lYUZRq9Y6T1
Y3Xb0WOZ3mj6NedwMdWvUT4iEhJsUPAAUnFtrGb7zM7K59WTfB5t+mDkpZd67IfU
VMXhJUxqf1WA63VerDzjGSLdwzvHKkLaHdav3ZqZYMC336S9Am+tu6Y7n1RnYbTA
e0HB0biCx3LbWjA6Z/Gebk7ryRSM2KKdE5KUzoId1fOOy6/a8WvfnU1vspTO3+Fh
r2k7WCQ6YJUiK2pJ79EawOuYTP0iweYWin5/7k2DpkfuGPdG8soJyAs3LW0KBkQl
BaoAap0GzaQLlMaQXI0EpFrfH2m4wZDpGHdPa1PfSdnZ19yu+SjzY50qXbHL8coZ
FOB3qJFH6yDtJkk02qlb04EeQGl+w8Rm1LAhd+nOXLbkcIZhHTU7HoCIbcHRbp9D
ky+NfMcPk7MfIzpjdT9V126m5ooU27pNBPwnLAJ0avOKM9Cww5TGuOLTe1IqVyrL
fh2SeXahvbzRW0gw5X9zThbiEImy8gAG2TmTEL/XjaZVJVxKulps/6IrGoKviYNi
OD+Cruj2aRgxDfQULzkT3Z7jiK2dTgyDiml3cpIQ/2RvI0CCOywVptNGaFuBZZrG
KVB0fnOhY9dUiODNnCcA8yxfYZ7XPqsjr+SuesVu/NyVAjv0kktb7EJL955Nu2Mb
Bs+IXR5fMZrxgPs9+aJhUghRe2OJxJx/ccJ4RA26Ccr3KOue5+gxVq2DCRrEiey2
z0GT6+myUK0+ZJ0daXuG7qS+wRU1WxxLpA1+VhuD4I6fpnE2Y0xuLfx1fVKPixmO
Wc+H7rxs5kI2GYrwwMvGKIWpe8HAz3CwRHr2yS84q+xw3nISYITno/GYc/SStbun
53wCqG5F4u5FmKAHOxtCFwzH44eH6+HnjgrxgWtk4HqIRgJ+1hnu/vwZDAJYf/hE
Xu40QdpUjluPw8IdbWiEQ1U5dJJsumSOB1UbzT4ScJGq2ejSY9RomEcTkzDZjRWP
hAlltjt44RtbjnaEhnoTFxb1Sp+faJ9+Jjrak3rZXw3RKiuwUH0YFEhBnamwnRfj
OtMfjkBd9Zu2oLR0KR/y6RtJAOjhUVkYNrKb47+nKaQMhWSuTeyuBd7KxZa6fOu1
txx8JdXc6ZcwsNDhrYdsxuordawmp8cQJSgOcZFGcKbpkhsZkadTPK3hzJikPFdx
I9DBratnP+/mHX1z5pjmN/1lWSo6pIAx8iimIunNH2Z0vOTCfMmlMgwqZ0Te9mWW
BjfmG/apmNpr9Pb06qxz0uAE8vXrdQaXXk41qw5PAKFd91/H2GeEhaqVYIB8ugj/
eiSpWZso31WkOUCZbHX7fHw4wf+8ab0FPbi09o7v0N3j9SnDYrpbkDHsGxtKp2pU
63J4NtNnhQPVIkLEEz6teU/VYxQNKaDLQ9MN8HKAKQ4E4X5lc1nb56lybYqu+mdb
EGa5NIxdyXsdI7zBrEmUILIAtQCBiP3Esos4vwnayoV73Rr9KMw9fRo1X3WtDoyN
o0yfgrI50ln51MI5/agi+SwB4ohCZn2AlFkVGebsRla+OOvaFJPKrJu3X032NuyK
OBm8iADEbrJSMf9Vb+kz8GRKdPyMdV6bV9BiW4V8vGoHGVYeELXUkS2wUVZfxXQy
BTdDTLMoL77zIBkIRDiWcJbT1Zdc46l7RYf0qwJ3JM3gz1x0/SZaB4jhPA486DfY
aDNmufGj/h7hmhudtTr5491dN2Pjp+4fXnGUWzRZqwAGQGm2nTlinxLngMP+moUl
ddqHcAdihYFMwG/bER6vH1GynPjyfxktCbSz/+QOBvRmYFuOroEFrmyvbiNaz8ka
4plDqQ1BXZ4k7Rcz18sxidL2nl8odtQU3O/XSMW/cOzRi1rUdKPst8yyiCq7awDQ
EJ7090Dr8ZmvcYrh0rEgwgZ4EWOb1rFBEH6JoapW6hhc3nD7L2ozBNUYNSq/dtpn
zarT8UOVqYDZFfnzxHnuUi4gQm0ZrxE2WQzsvUPX4kLIrHy6HqiaMrj3F0rvy74e
NbDcGpfoLgz6LqgcTmHYcA8mfZl/gXMTvghJGmgxi3R8dkpbdKreQFUxiE2ppzGq
8YSyryPyv1Trwl3n9anjs8zuPVDqlyZpENNmVtboPTsLfxX5gSFqC5pzvSZkRjDv
0H26Aq5ObRTrglz4uX3Lo1dgxNEYclriAYPrk+zSJcI1X5fdQI2SZOBwTzID2N9I
hn4AV/zkiU1KRPyTW1tpdXxU6ebC1H3IGsh2Lf3B1uZ2/VL1fmcCqT2I5RQpZdAF
IwawObZp9KVaK6UZr6B2F6MFffYgraEaKqSXbYehYJdCWhIgY02MdXtaaGaQxNlJ
stxj9wtryL42EjF0pgWdgKEHMokJcgFvpnD7T4G4fTx11A++iCPN2+yNjfSUDw19
9LWokMDcokoA0RIerHuok3l62kdcqkrPiQgSeKdPl8CCdLORmDiw/pSqULLiksW1
C3lPr9u4pZz86ca92M0r4OVWxw4wBejipCHlWMUWh7ZHRCg96G62HFSuJj297DaE
6a/2p93/1NoAUBVhOatQnDi9wGTbWJdxcXCxJjFDJ9BLi4U5j9/Bp+pNFK65gx2z
jRgHoc86XkegPqX2fZjIu1xDwnXvP0wMmTq64noROcDIeTC+RF6c9kJBbFnHkJNd
k0YavTb2K9v/w8FsuNkTjts3Qohhg+zJoL5oeqCcGFbUPRJLItB/8MQKgFjBN8cq
ZaRNvOExyuHCBQ9tlrjAs5ReoGKSwhRY2b6h7DVFXCB862uC0eVh8Wi8ZNh6DjEE
KiL58ZRVjXgfT5S084n9+ifC4fY1VUHtJfj0ZJVz2KJtosTAxMGe03G27zqCbVoM
rKCJLtD3o5hDacXxQniG2JsLyyQ+qrW6Ioyg+Eb1KCC+2n6bC2HV7TKXXgi9QN3a
4kOPg3CaBt0UGEO1bErqfEpCxxx8Rjy3Rl3YFt6jhkDbBxVBQEhnpG8MzF66Jzz1
DzVPiUqMW87vjRoqQgBzbJxix2QIRdj0fHnLKZY/teHF7/k9kQGvXiy7dsv6DQk0
ertMc7kO5S6X1vNrxklKR4OwpFxfT9ak1VL0frr5kv9wYohPvKUu0T9cMD+C1KP0
CdUAnriRdOeKvSYU8y92Gku4il/YmuSimc35WhM3VPsmvj65KB18Bxg4huVsAhsk
Of3BCHpag/LszO0/ZXrYsAx2JIFAOAoHHimYf9w0UmdFBq9bucg/3ILxotLIdHUQ
6pZMx4vP5WwMJWkvBZbNodLdJhKHIYRAqKPGd1QGobe5EkxYG2hZpTddSJ9XuKYX
Im3zh1xfEIYfDX3GCgl/ttSpYn0EwaP5YopGSsu3d+tWvVpgA97QZNVaxD+jlOm9
acvHPCWsFUjyeMBN181YmyoJUgGM085MVt6klZd6vgzW1oIBhxV+nduaHXOsHfQY
MUFvgv+ehr94DydIXSNcMhx8qNGEfOpI+ZkM79pdQbIxpOETL9S7CaxlHAko9Xc4
iUTbhRe5QRpGJ497IzjZfxExJxghgBX9+KU6+qyPnoAzRHtSs3+sYB3d0DjVAcGm
pjoM2Ae8fmqDbaZjydarjgBKOK9i3nzurR8hlwP7+D7isTAEZGNc1dms9JKX949h
1BBCDcG3H7du1zAc0n7qugNsncWmzHPb5ErDO0ao4YBAKsqlUBss6sfV7wjSy1g1
JhPRSmkOhtfZxKBejFqLfTL7ZxSiSmJA6oJ37omiBRAnbSwKbB9miXjzFBgyqQND
mOazW8uR3BSGCjdC1mflTTW2fUaj8QIwMCPJHRtlLd4Jfl6tYBHF81aVK7zIY16i
Qk6yrLcOmTZcUO1aCXk0ZA6cFHBvVH1H40ekf9w9VaQjx3rXBkRLXCy2UM2txQFh
v684OuXqvjAV5cQSHTBVJ/iHRW40bBlIQ9QTGe7S9aGzeQrcA/vl50Vs/dxUNC0U
g4clWkgjTh5Xgle8eunp7n3Q4gUf9xDZSj1zzjRr5/FN2BU0yeVLBqvMS4WTintV
IqUdWnTC8LTZURS3tf0ksFZA3YzKpseYHGm5VCbAkIOomiKfM4mTKoanB48BoBp/
W2KanaftCGJTKVt9MtLxfyrdZJFTTodESTvi275OVwS84lNr2JMMU14XtP0BJrvT
egx9HWVuF+6wIAdoUOGpS3jnPcA6JANp3VUqh1VX482LyECCA09EthRzEthBubA3
+N+LmH+C8DRrealt2l1f+W2eCSypxJC7wp1zLGHFfa0uhgT9LupUZlt0B0MtXMuv
TXS0Xs84WXuUn9yqpdAVJfK6WjNlsp0Q+9t5RNBi5BobDGQC99E8RIMZ/64dq2dk
yZPmziVQGCkMTMHZFES67qvDMmRhfwM/R8C0gqur5mJh3zTlvInZMl3FRfEGlJuy
SACT3DOfVBF2SAlJFzQsEFVS3KSYUjsVmkKH3rkLpYO67JxjfOmh7u6mtYl/rRDx
b4/hElAiUFiZoz7LwlEa9z1IMtS+iI3kwlhTMZxXgSO6v+XEAXJ9AGOyUxmNbFYZ
3japkBC+j7xuc/hu/zQ4CyghnJt3ngde4Zj+PMA6SEvB/Xu+8nb6K7PfDhPgGA5V
ONjvNBjIZTAWAhBAlyvcOkFj0newlj8zxdchzw+vFrYUDXGr6cJE8OI2f/v+Vw49
+4/CZYzqfZvsgUszQ4DlXxkG8tEVdZ67K8zNVkXeZE5GG0GBoxq/yv6mqrRjf53l
VKBDFyUySmrjXZQUNbgjnCOC/vdIWyUGV3sfjAvmABbEav5DFYKyuJoPRu61HPvo
zctzBHLGTbB/dabOo9w+N1ThBbgnFWbAycaiuKbl4rXhhWJdPGT39Ujc5ZZAT8dj
qsyWHs/Ikn5NvFsz/hiF+FMlnqHIU5xyT/4RG12accjchzNqkwMPKqShyGoIawDW
vgzBDnpeJEuxl9pG93J+diiXUVj15sgnV7j7CzNplUysPaYcS4boQmiNel1Mke/Q
0dr/+VlonzNERQ9L4yCRSc6XsrOe9QFWM/Zudvc38RzEAzjhdnlLRCHv41bseafS
pOUeGwdGxUPdabpFncR7US+6YKwJb6gFgUP1AXZ4DUVeVtY4ryFzuUQt7QkqQJ2d
ki7Lr0V3yYiPqjdLubVAKxFPTe0u7f0DT8LGKVaLc4qs6iKBk5GX4AP9ccnexDG8
8x85J9YmN29e/xnH08J0avr+eJDx7mr6oHUz3Gnd3kXbzJW1l555N7aVTquGS1RR
OBAShellioDbxJ3sasQDclihF/UlJ+BozbKLmm6yuM/ZoeGSVMq6NV7BIzMyPtBL
lUxq1bcIL6oZARPxnAGrAGsHok7IeWklZAGlUyw6LRJYmrcZ1x9pozaNwDuqmeX4
yIIM8VRfoCkxC41EYjEYuVq+J0+A2cgW6CTqdv0moaxb1T1d1VeWX8Z9TVplgPqA
+mboyITRuUOepyKVwMXklj6xKGQLkxrJJ34V/GifOJLlO5dXetwaV2B74NHy0xSB
RvYNTvCpfS+0QV3tYpbANMIqWyXe1zVuzzA9GgikU3bXLVHJaYzD7t3tVHPxRMfU
P+21C7PBdqcRBKhf0wqfvOEfbdSpgelTY4dk5OL+eRGDLb/NRpHSCV41U6Db7MA2
l99w879fzAyb9W9UHTpPe+ZLeZDH6awML0doQO+MDiX0mQtsWBtNfDHbbiPuu69P
1/6IIpzP6KYTALd6sUNaOXLwM4c5+KYWRYelGQ0BOZOKQ7gGi7ZfSb/vNgR2EkQB
pSwPoEu3gCxFPIzqDSTg6G5OAuBRyS1RWvOxRIDLn7gwOyWGTJGnpEIhtUydQQgP
RL9FKgLyjVbnbcXVlPeGvotN60Ub4idm8LSby3QnppxPmsKCdAtM03B0nNSOdwiC
vqkXLJjwaBK1kWpa+lBZ5Uatd5eRgWrOwsYpfL+uZNrkYfK3Cbh82Axxwtt5GB4n
t3SwddAH2/uATOL07lYYY/vAhBoU/JftLLMeCttLHwDu62D5EeLM8dWYJXZT7pSS
oAbD4NS0xYZhrOjYehqVSv9XC9hH5lWovhy6/SukpNH6Vww7pWCSfQYIp4dwOeUn
uJtnPOjR5lYi4z/Z55HjyXvYH6kZKCN8qPLB4S/mvSE8R/qMUK+1+Xz18RbaGqwU
JkC+txWlumlNE4iVavqJtdNY6uhAwolNF6xzxfZ8zNk8gT53VL4ZWs2hgC8xQoF2
JeO1RSIt+6mZN131TspmtTXGH02PM4Ckkmd2YcDZEtltaSS52hC5B/SET5dju6FH
rLpxO6MfaBDgvu8EiKbuGHsetc5C3hOcSgZCV1lQd0ULuIbArU0CBD93s+VImgTf
lenqSGT0D9RzF9MftmO9ktySFxUQEwlTBsUsgmX27qR3XmIzQYXVAhsS1gJ64FkV
2Mph5VisiPDTr3w3CaW8PGoKMl0w6h8C1hHuG/RU+CNyEJT5lKveea3HyTmuxV4k
bJVHLIFlx3+z7+E1RbiwPPvvUss4lNUyOVSLYA2Yr03IoednlZY2QjURq7TLFZii
LXiaKTiQ9Lg9JxQLB03vgvMfjntIXFmHFgCtynvceDLE9StaHMNOiIkzVs3RINC5
Wp159lSimIXNf8H8jiUl4CwFL+A6DZNvq5MjD/Pw7HomczcgPnAKrVQKYKZPLgSQ
gAA4MeK6ZV4npNo1uW4AXVIa1ONQjX8pAeAbdp9DNTXR9p0hpC6ZBK3TmmP9F3+a
dxKejwvyRVIXC4BVDBLbSlQ45LD0Q9c5R/Pv1G8uW5yZ4tWA8s47MP5KZsL8RDY/
c0IWt2724CGZS6Q+gBO8CgeHuviD2oysGHjUl0K8AF2l2r+aSb2WMvqQtCPE93R1
FYMhh2Rk6eXWSmEpkAbMQ4jHx7XsM4tpr4u9jvIIfK+KRoan1MouYuTzaK/SE9oR
OobkAsBeU1gvDhWeDcbF8UdL++4gTGNDc/QKie9QBbU5PvXfyQrifsNtSg19UPz5
G5NMFruxJq2WL6yhdgd+af7ZE03nNRpVubLh4XaxsjsvMBYXYkhQIFXJbJn37V7t
xvf6uckG+DY+/NlVEZMlupVYD4RiBEeoAaDv0JM69c4B2sM8PF1pfq32t4TnEZFT
KrX1Qw75o2+DP4qMHel9C5k60ZHXMLzfMmYQQLpyC/SE4nbRdob0WbHsLVC/Uao3
C653QlEVOrHwLP49OSrRsG8CAQjjgEqkeFJhm7RN547TDf6kn0oYBNKww9N9iD43
xAaVUudCxqpPJB4Ahvi2MyV3jiUhUZviEOZpBuy/bVVAJDkEGmiYu4LAjnJD+85a
oKZ4Kg6gTd+jEwLTMGtZkN211s+xbsfWWo1NTc2WXpilkcamxY+XY2cNiFRoLI/l
8a2e5/TU1ksj+3x4m7KAwff0IpYWcXH814KyBMPjFjJrxHYvS7Rk/zF23EGEhhwZ
IPJwNMeFdUQOhjnArAQsPPvF5Y3kFCOhj6mF4pe0b58uLysDZglQDwvbmkfT0Ubv
0WAC6VdZMLWB541tkcAW+moEvu+dVI3G7f7ajwuwnPfe7ouQn/BCVLF4XvB2O29/
Iz3SZkxV+R/eN28cTVQF2USr1tdkRA3DE3nFfP5X3QrtsZh2G2X2nqi31t+UWScq
Fta+RqnvtqFVggW4dsZtwE1EnIHJiR9Wj3dArWcAGnjiz+LDdX7rln7Jg5TBHQqY
Posdb82xlnVE/IHy3iB8WWmduXtmT0641vwy6zEdkRONeFAXBkkZ8T8TaXdGp73o
XBA17/37FVn0oMZuAF4Bfa8HVls0b+G9k0LjLTxUEFhQFntI8OnWQMitqUGlCE4a
bUSRzb4+RisU+ZelaJR01Ank/2c/Js8Ab6EE0OAdJPjuJJpNJYAaXKLV83dQEbYy
nnXh0fCU1lxMLe1JX0LvYZLug1MZSWjnPz+AdJ2liOOZ1ENZfB1kKWhg55RN16p2
PRxB4po5ZyYSSIhbfyxZicOSp825cqaKD4vG2lhj3bWEOvt0bxP/J548BBb+ws0C
SYZ5a1i7Y9U8iYjtS6letNrGdOAFeiS9g4cG4oWXFH7RQ2sTWQd8Ls1KfbndgxJn
X9q9f0aIvAqGIyi9jWcCVyyms5w4w5gGSFVgVuo2h+EKfhgjsaI4ZWNYIWyBlBqs
YYVhdjqB3QN35V5tfADJ+cocKIDOLBRC+NkZd+qcduvy2aqu8BFpfPgWbtLhoqzN
hTri2t+GY1dV/tS4eIwiPVWNJ9Xr5GnW6KdHo4yXcySUoFBmGq4ZHsHikLn83f9z
lovkBEbJQ2hlDWInCbojprV7jOHtoUkaKkV3lb6VQ4mwCPLs/5W7BpIwGedCsjhk
0ZxCBiVggSNk87I254p8BnNNsRzMDRMSFlBPfkWR3ZAazU1FA67vz618j07DgVq8
9s48yNr8cVWGI19oEtAvfRXsGBZGLEYYbxe6s6etRi++BBE3dWLt0s74bwhxq/8v
voaJ6+62lzgWQjdGHcNbd2/Ujod5sgRhsiolQHsUF0NCFKEgnYiEeJywXDDCKzuy
gZr1PxQCB3SRteEM9SoiPeCziakUFoK0hyFnuhelGl3FQfnx0zrOMv00/LA3NjmF
hM5ikysHvCeoRit4GPDfAPhwia6jJrZyfZJFYEQkobKoCSa9UQ/9piCX5JLoxPGe
Ly0046bIoIsJ3/TzdJVE5NIo6tVWTaRv7qf8REU1pbAu10WtIw8eZYu/fwPN6UKy
bbG4ycvyi61eTfL5dsMMD7D2Bb/a3INk7v0jskikqIkbkoN5sWywHrOJ2nAM1a/3
95fKmUl7RgWeysxR51Jd72+PQfGRFU4SsN1nrULtqXWg4NCENJR6Tm2icya1Ln47
PzplOKTKh6w1fQxAeu7WUtg+Gw8wAvdUzpplwbRdp1hxvzxrrH9wioPO9GFS4Ak6
cN9QpWEUYsT56OAEeOYRmfzu2DMMk8ciXrEWNVvKQ6w3pizQ2sMSPba66IKHNFKQ
q1TbxGoEe2nljioJ1jdiPfDTMfcOpZ7E4msicKELK06ZzRzrz/TydWGv0dShzMh3
GJ0zuiXWtjncyuJJAIttMDFQ1Ki34ZTjLP6eePka6GZJQu00J8/UUk2JCfHrCrlv
T9ITFTIUFnRQNWGMr5O2Wsy+OOPssU4f00Dm+nOopN8Qw0ZkIj2C655IAg0eL1fS
30f8olDpY0uVmWlwnzZPJ+i/x8c918NUriPKWaxCbynWeSpclQxB3sk4tm9VEWVl
+J18s4Raruix80LH3HW+WaRdQMHAT4c0Ya4o6p2vLXb65PWtKBK9MwRxssLmOn11
xHBvVNCYwL9qbEpHysSVVLX+UqsOemWXapFCN+E93a6LuIdQh4wdFXTLo8Q1MBZh
Upz65QXsbyzY+n/T91HxODE7zoZTbAd3a0fKdOYQ4hvobRWFBJDfFu2Wik2/na+x
W4/3owZxwvou7tZiIV53y55YuUu2tCuoRcBq2zH4vcPlkOQ1Nnfus54E2LpQ9GjF
sDT2J7cAgmXWAwSQKBfXfCWh97U8VrTGBxYaY2PacHCk13iAq1Dd4VsDTPDeFq77
kW2/lUGu6/2ti0F+wLfq7qnH9uOeooCoa8/AodNMPU+XxRpZJn/tXGoNriHsK3sr
jaHfzd/npvmsXjVeoNxUhJXZolxo5HklHRL+AJymeluahBNsmJZNiPkVFKPXKxyg
GI0EmKejyzE4GJ4huZEjTZOq/ec0Cqwgekn9Y4PkZZrpktTnZgW/3/3UWCZmAp1z
OOYM2eITSlSqA+WcOeMxuN7kCfd4E6fynbWcw+HUIZdDuv0ey83r8uowDG3f6BV5
e1lvH7wJORNI3FPutpbjyyNjNlpzP4JT0bqJxKJuM2VraRAFkUV3gcDTAfOYIH55
R/nOzvubc7W7iQupKE5ScTfqSa+FLJFVjpxZ0WT6j/GRx1EUCon5QfhbcXCzsZdw
KUWHhWn2GGZHRawGImNC51O7iYK3nsgG0TWozzOfMieFTFZr2/dFcCGgrAtXQT21
6Q4x6XwgIPj8sml7kB+/Ljua5I2e1V3l7+70jZHrNUNuxEOP8VtRQLL6QE6qrIKJ
i1R+DXRX5NaDlYYzKoDCPcRDV0YVBU7Q8s0ibZ2HFSA1xPXNyYg9wB91l1IupaGe
l4Lk78YldbJ4+dT+Tl8uJ5xWHaUg1PXXUn5BD3b6ryl7WnyOxAD8fpPZPD1yY14r
PEs8ZyJjm2Ci2E5QHKOmuiji4Z5MoUSeOhKAsWzolg1cyPF5KGj1ddjYEMOi9ScY
RNrT9r+4tpfoTcmOLQaB+x4jTVg/eAj82/MsyAFdN9j2r/gLaAPjmztTGQmniayW
/lVduY66wI1lsiZFk9gJKx4MI9e64jQ6R/nL7KVkZQWTdoqKidrNusf+Y6bCeqxn
2YyVMStpNggDP8XEOwHFvHQnP320phM8lOe3pVKldcTOvQaeCS8/RbUWKBmwTuka
bSqBvYi0qZD1CRlYne4JKP1iXfpjZHDmkwvm0X3YIarKYeoQtx3GTaeP3yjVUZC4
k0DZJ99nK+lC+gi5vNJA0RyNCQAIZ+n9mUWZuvh9plhsbEjOs7bJwwiAzlDXh4zI
bYCxjSftqKqy2er1h5iwiLRc35NZICLvRS5UZsT9lKYdNntmvUcdx/4baOGUJUn+
C3oyrKWw3MkK2SNqbcgQ8OagL0yC2nT4AURUYGn8/CW6kdPyMGhkSmCT5ro/rWZm
YcxwZ5Afth8ASlKcAvJYqw8aC/MBnEg+l+inLDoXWPbtw2ZrYFzO9VtezkAPhTFg
2SlMT37GWQFFmJN0+DjR02Dh+FxrXO/CWQT44PpMOEhaxpMdMl4B4chPISj3JIYC
+Y66HKbWGaWuqj1IDyKdswwL6DPlaT/ZPAryFZb8o9lOQ/j0216H3Qq0EUksijnt
QQR9nH4vydPEkhIJyG1SZDCKv4fyXzxU/8mmPWhUAIjlcVomWVOZ2N/iEC9dtSD4
ACkUyR4qtfEOVqqphnJxYyRi18nPLq8FXr4/Kk8mkIYSuJDKBHn/HfRR2UMN9pvy
X0Lf11ywoZ3v2qAeUT6RibogCyOxOqEdsrI9Fs/XOMFGwdvaswZ0l22PZ0S3PNuB
4Zo6nYd/qOP2aHpUzy7wP0jsqzToiRllnoe+NfQ5vDxDRz0dafwsRDpK+2DsJrED
IT36PnOxycVayoxNv4yaI7vZzBUD5jptE6PYnPfx5idwOXYwe2sBEGyVFoxWkP0T
nl6BQVDjXC8WAw+8n9HQJs4+C6bIj9rD6mUOnCAhmUEhddz89H1gmYBChTivYVm2
t/OTyVHuom8PsLj5cbFH2W0xG0msthjsFZNQW4uYnJb3/m6fjywHMZRpVx7EPiL7
kcbRojBd+DGKgGt9skeEAFF8ysr72TTg88DpH5SY9+r4pHJ+FHKxzeAgmHTyt+iK
43cel0aPzvHAF4zRpBXfLLdJENB01tk2eP2hR+w0LVk+iuS6t8PE9DigsdwR6c2M
1qZpljkYYqAjIO9t+0xRjYbv4jAhQTCyX2GZtWK5UgepNZ4MU8oLIK7iolNIQUPv
9STKEDat6/5SrfBBAh+SsTX+oTL+NmefrCZ0BzKi3zt+2WmWRhhq2wU6iC+3MKJx
7Yfui0oX8eDgG5TzLBcbgIMiTn367MvdeatC9Y3E9eCMco1bKZeg9+YcEVfACy/s
oZD166eOkTlh/A/d1rFlTq1M4MruHJ0NrSSnpyP9LrAeNdZ/qbQp50vHh9RRJDf7
hOcFXAoMGSk23L7+i7Yb/IvPSDk2Tv2isbbLWzN80gbT+yVj6QN0KbkTMaj13n6F
xxri16Q8Gfwv9F2PDNltksJk3//MrHfGA9lK9QFtWKtfHtefleJ9DWVSsII2esVq
uvoXRNxqU4f17pg4sioIb+yNlPz0q9UHzzYyzXVWu1SuGZHH9/7FhA3Sl2duffWa
1GcxGjc6NfLh4VKNYS2xjXrmJSGEh+O1iE3NLT46I68cJq2qnNW07HRxMfVtQNfP
rJfXUix+Dj5kLm59o6m3GPq8I1/FYRgaxtycZ7A0fLM3A9XcDxbsDWjOWCc+nVAM
4y/DSHotIwbMcgM64lP58qdJBhSB/7qmKqA21oVvL6XYLYfbbRNFnB+C6cXoHVto
BQpidJczB1IYRg6fPxTIlA/8W6vLm7iR4vuCvYAT9mwxZFXZFg5beH1mtAItjM6h
VpWxCNBdJXDDVCoUaRnjleppwjeqI+rLhnbu8pUE7wOosCbQtDJJ+yhDj1rBA7cG
hykuQYNAFbSZrt9D3PevTvi9MlzW/AjaWZ8j4WsFLUDN5sdpKZQsTlBhynpx6Nxf
NOlQC1ULwR2n/XVibOUGAePkM9JuyubvE1+QvdqjdzVyhqVTcIHtRoas8lAS2FMi
kQJ2RVk0z87ai330ty4wYFA1gmOSt7A9EUBU5t/+VRgpfV/f8raHGDAmlMJf9A+5
7nU1k0jDp3yZoAhinUF42AMQhhXF2vF3yuHxilhxVyw5v8XF+MP4BfTEJD0iVojg
uyba4PdzLTqS/cwzjNMQoWdWN+ueujwTQKbirFwlpsa1XA9EddwHbK7dpDMDe2h+
y9Nw3l13+7C7AhlJn0Tr4XIMG9EmgZ5yRuURPNFz/wCqdGvKccEC/Dgchc5RlUcd
84hQM2W/qxqK/C58wrkOdH8ciCcQjj6/Flx1aC+p5tDQZvjhARgDTLvLN0fO4aHm
qTT40YTSAilf7N+A3YMDd66tLFTqJee+JCTv+TWEHeuvQl+FAmjG7d8vndxh5aAt
iG9J9GT6xpoxUtiWewt4kX+UTwjA+RXErWUV9K6qcgI+fg7D3Wo2mI4Soid/lH1L
Li4Xd5ek68HzggYDrxaLal2U2EpetV2NAqml0pkGNubWN0OcJ5R1dfehx/fSgQdN
jRrUl9Eexp764+QpxUPgCwMw/C+/p5XaNdKzR09AHQ4PM81imfBZ9yOGVYV3aPYO
qSOy2hwxt29/Q1jwn+p4aAek0tOIgNG5NnnhMLdjHjdxETF/C39VgIr6DFzubQis
F13O4GGaJveXtsT4fA3CFgkIF/EXHaeRMXwCTGaKLNcFgoJ+HFShJmPxuf5CUrjI
03mOtyvHDYE8yBNk7H+2BSVW734p97XLQiKqOb3cnv6iIQB8HVS+PwRMGkIhyBij
WzXEZIVb/W4VtGzi8Qq3nNwX2wFtb599a7WV7TcHnOIMHbqIXiO4LvIZsIbC5+5q
uow6QyA+aMtBPWHv83/P3UYYqplQH01+LT7qeGF40YZD3HBvYhRhE6zuCXP/U6Pp
YxUhFaUddx6bY2eexOQBJOprtDx+HQaCsLbczH4WEcDc0Q2Rjq4VQGJco3uoLbmK
7/+Cdhjs4Zyd6hgKicbNCDc1e16AscyFE3HXRjFaZl9XY2LCGJ+3em61mgM3ZA2K
F/8fejPq0XFb/SKwVAESpZXMcpVJ66gA33C0Njn46qx8WbWzLB+H0HLQe1+drHqV
UdAQ5GjqO5rRbwbOLMX+a5hUZCDKZc9C0lmBz3BJpxyFwvwB/U6bnLYxGsPPLh8r
mZ1FxSD7CXgYRA7ytnJNUZ+830nFFw/JpUMa4GmlWWs6em2GzK9gGjS4oBvgt7bZ
+33I7b/aM3BiWeUYcMl/GMl4fJbA9f1R1zzfvKEwtYFKzzg8j+UeNtsOxwGUxYuE
s5wr3zsy/vq2OYfURKh9zQzwqN+7/V1Q5aNKtVjBq13ONoTQvf/ezEW2kpeLl4rh
b7nDCoi3lM5lufIKKlAPLCl153QWE7ROmK+UUx5EdstIGs4xBwN7ynprJFelkEt0
ARuIZAsNjZdQZj77Jc0bqNRTSmlTX+EwUs/s2jTKBsUoryyZnhoxy9Pz3of+r+X0
dIDCknm8jG4qq+6A1nsuvwv+dVP5Og9l+nGQuN6Ex5Ce6U4fyULsPjFCYPEvgk8R
Y0Ct7XzTM09Xa3MC56JKOd/tpx9MLqHb1MJRwnh+1Ew5Mje79PV5pDkI1cRJop0/
OTER+tJBzS32F5TgvZ2Fmhp5GA8NAEkU7ZTwC2SiTX0J1MiDdwKD6PlS6AJnFEIy
Dh1xjWSEZEiJIeUwuHRXn4VHWCuQzctUQ/u9VvZyZXXBuxcB4/PlTDmERF5cR0P3
5O4lE1Zk7W5d495N6m9Cxr/wgVC10fW4pjTxeh3xCWPSxmlYfRl9H84Vb76TaSUu
tYo/yYTdIakw5druWGOdUwMZflrCCoARTUPuBPJ3HripAXrZUT1+yPeMb4tuo/DL
2Gr5LcwlArOa0m8q6iPqbu2cumm7zbtyAIitTJL6mY5jF9BXbWU7/lLp5UX0DgO/
TiGuGsw8mUR5LuVDVRWMRD1hL6IG/7FeP4AH45VbXcSkuquWp8X1osnac0kpTUnF
1uMPPsY26NQOfaVPCGMlAo54qdv6gonzYfZvMR4T2vSUnythRzazZo9jP8kAvp9q
kWItAqKEemL+Z0IK82O2Ownu8arz7Suh635cGecBcwZyPJ44dSW3hu8gk5vZFO04
x5b9dLAG3nOXEAXOihmYVPCx9EEXVE+WNM8UTO4hcdsFYOR3PDLpqYn/efWgzGxO
gHELQO5jc1kLJ1FmhcvOq/RfbUzST7P4zRBq3TP3PhCQF0TwGdlccFzYMu3KJj9r
lm8MPiNovGSCjJVRZIfXf8sJTb8G1cL3mn09vGq/6vBM1N0koGTsf2F+NdzJUFB7
C/u5hnSGWwEQutaHHCfsNN5OaBs94QXv3X0tGmxFrCvFKZ7z6s6Z3XU9vRFH6k6V
tGEbRX8N6XAWeuRF0m/ohy9wiZVfECkIMLTZKN3Vg9XV6OlaAx9jck23QRhExABX
VkRO8nqxDnU/+2Y+Ivg5Jx8FvMXcn+U4ar3kOvZZBZId3yIYratTLVgv6Rrb0ab+
4u5rrNhZVQGsu/LXW0YOBbVei6U7kchHL7bW2g2sm1hKbIaESfPoWMP1IMy5jC45
/AYLzQOorrdRtJkgYAt+lSlTz4IRCsnRoZK8PzcbFDm7utG22QKMQ1zcdgaDS3KB
Xde6LgnSejtpwXkhCmFPF8BvyX1oHqiX+hjvBSfgZtq1hyiYMw7EzzpPbs2bswkU
Sw2iw/KISPZD5T0gcNKHT6TrWz7/q2BooZn+c421uvCWv6fV4fHh5SpMgVcUCffG
r9Y1MD2eC2tQzHaEV+lggVv+9KhDf9D6cStFn9bGuV2AOcp5guTF/k0Mrpj9G6Ck
N+2jStB9u8SZh9iFwi0hzSPflo+eJgOufz3ZF6Mo7NTx4TegMVsWRCfSkIII+EkM
78l0vnquFdkE3TetyJUT4pc1Lwdw8R+uHylM2QmIbQa9iBzrB9HRMXG+EESrv4Ig
O4lU+QYYo3C98rTO/LNjsvNd1wk/FVHtsghOjXcnRVX/EVDEXGnpVjbozop/nzB/
uTsUlz55vTkgnGRz0vOV2pJzmlmXumHHmMm6p0xGpU6u2JYMrwigdzlohqrddjlI
aA6YGHQ1ZvVwTc1oXPyghf2TkKK2CxSmxxD3GOSsWHhXg/FsbM05PCMU7zZw6YMF
mEsklBNq/Tg/W7PioClDel8YQI/tXWNhFl1ZzUem1LHB6jeGzuRBMOahW4CIdCMe
dEmud23hkxSoof5OXSyWP5AysdTUNT3xp7keWPZCiOZkjvEeLvc9uzUr97kZZkbx
7x8IVPZ8aEZsjjBJI9QmNpeMTcNJye0XpOc3c8IKuT6vLYX1vSnemaTWTko7ULAy
AgzhrKEOWw3ZoHv7WQkoG4vPI9PX/qjaNEJNTPcra9I7Ve4A6UsgsuL3iv62DEEf
b59HTJISVY3fZJAQ/CgvVubZmXpv7onf33TlvmtrOs8qyYM+Q/Dv0DDytqZo9GE/
7MNpFkiGFptRDSm7iBFU7SDN45GLvrAxApunq50/KAMrpU9RDFdK1X75T3Qb42Fd
SzFAd2ZM/mvvJNA+i3QTtPdkiuNWGMSFr5oIyLretXFjFbszrAY3op2VfNDhoZxd
7lExczwYflv36/IsEoyFysmn+JiKphBb0qkwMn+IkbB4rK9qkzv3w0g2643/h14q
MHGpyjKgyu76cvtoY4sSrDPMJ4LueUduH22yAllYh8p0ZfsbZdYSk4rdW4whrTf5
TxxgDEg5zO09lXfr63v78RzZqz+C0n58oRUZPJiDL4J4tqbRRIYz/xJ3vZwPrfPM
iBIShXubUvQYfh2RKOdIllhZCBGQOcTvt1SrQVDJ8ZH5rfVhWJLcKTafEkT6zA7I
vrEn6Y61Vpk3IVN7kkJwq2cBGFdVCBLVlJk2ERO45++Uno8ta8SzVba0Ckatdfqz
Z05XnATMnNzhCebZlBk0FOGoTRfBHrLuQH+Ywt0Am5B33kTe0jL+o5yaDxJp1zRz
q/rTEx8vAOyq8R8pwTtv/Qt6AasJf8JH1pd6kjs4voBLbXncv1aAzPzhkP7Efqw3
nY/K+tfkjcRTgo3IMot3TTyBh0JsZ1cqYYZCjoe6Op+dmPLivQXynG5FbQdgvLjg
UJGTu4FFLltZgGn3lMOcPzVJntmZwVq6m2J51DYHBET6Yj/9upI/1HS9KcFU8Iqs
we1jmz37Ea+TUugXXTPvdDtNIwSPIo9/VndgkvkCXv8EWLD41BNjHKWRF33pyIgJ
tH0MLExRYvuC9sK9ic/m75k94oH9paAjsnB7r65yWJRhPP7ovV7CS1HLhvvYqqq8
NXSTUbn88E+8NLZJjBLozB3D6GzN8U3hLwLnrjQnDhMtIpaiSgpgUjbY8kU8jGSN
Fel6vcflxKxp295JQC4pJgPoRyjz9fR+dOm7ocAAmuW4XtZjlf8cHD06Uaqtv/NT
dtuzBVitOnTg5CHacn8xMtlOXJaGkj9YBKw/gCDUENsj6yx5AY7veM2NCrrsi9f8
KpML+4u+6Tsb6pk4Avvt0Vz9hZzUKsoOe0YVyBSkpANXkZHknjKC0QaoSZHIeQqX
Bfv4QTMAggyVWpzaeYHEiCYcWjbPdEyw+svaHnI34oNmYyfRKZU42tty1Z8d1Hio
+JC5ogjxPpc4AQj889U+KHhxswM0KaZx45CHHHTddpWaATA+wB19TLxQEdZmZu2L
/suXUcynOR/yt6sanGp/k28phNISeZvIWYpLdcBQe60SXMyJ7KJzfJjjlOwSchq/
kdSbArD3Jpt+yLMIVpmzvNkb7SWcUQuTumSQ5O5p1Kr9e3bb9fehuQ0tB44InKtY
Uw8DNW/44NYbZTtUR7SYN516jWyF7xyPOR+8sseYdKRnhN2UneUhceqQHJ7jRZft
bhP6ORlNW+QTiw3jv2opuFyp+58enDmRy2jRIp5bjfEa87pkssyrFebgusWcmIIb
OMJ+xbl5wuRetsil81TYq30xS6F+/9BEw/rW6KzTYRsVqDG2sVEAZenfobpW57gT
SyQPSYFK8sUx6CDnDdyzGRTAXXn9fn/o9MeoHLhEqQ0YaEzAdfWGglYqmyjGHiGs
F/EwBvpyVULlM8am7Uun88Xw2ptMut2G6qiwlyRlOFUj2L0Eqhwj61DgfuVjneoj
5yDY81J+94GLH8xKpccunTYK8GGVD/p7U3ueNzp3hI8LRKHLVHAvMtDDZIjA9f+A
FVo9DHFSSUsmPSGWr2FeL+Vy9DzJJMplKl/X4Qa8GmWSEZ7TLY0vJjXifrHMl802
eh3+1TFGoCQLASYVQIHIAAr3dT5cbkCCWhu79aSkUAk9o4uEeF5j02mXMVJYG0Mg
oXd6WLJXoWsE4Q3NXtJ4C0kPeVQSJG/ryolqEssvKvgvoHir/6/nu7JMsStZO89O
h2It0dbG0R7074s4XrGrWlrFvvNfDf0F1OMVjLiCnQDWO/t0nyUSSaV8TryQouJa
8TCK98jQSlEda9PE+NEKJzbOKSfZeiOiZurQ9ZjKIeFjfp/bXHFqH1YyxtEsBCKP
BLH4SUTHe0GMZsi49pyv+UrmCvjphpOUgTMg9GpVnFF04d3ipk6S+gbs7ytyZwyD
qNlYQ5vmI6uj2nMNg+UV3G2RcJUAn3k1DvB7SIg66MZKEYDx8hXsSXk7RIT9rfr6
/GHGpuTXaYwAZtPyRoIY1mPNgkWcsEG6tL8QVJIrOV3OsWzoOThYIrdcCMMYRWRm
7z81YGC0r+Pol+jbQ3mV+g18n+FiLgxj9oNKPc3W7KgER0H/hzgH+Exx13NgYXt3
OrmRaEU9DcKHSFjwS3odx8bF0xY1PzMn3K6UsAzgOtpLyf+nrFX5FJELc0ia9Tj9
JYamz8AESslCFX5YAcqmrvP4iGjJ2atvfforZRU/11+5M0WKNJRqzhRzPvQzw/gL
jVS4SOBhW/8j86/sxK6gwiWlW8B7+DAKAARhnEksVi1FbUht0SRSD2jjJTRiOwt6
xigE3PI76lMxEYCclxmaqcJPZEl4kzaW8wgDkhNvM0BctMyRfRADCbO+ztpza+1+
1HiA5/YAJpRvtZFtWiqi5/2GeJN8FJjxgdQi8Nu1oDAhrAtZjITDXQDxVg10RzPJ
VNT8/jwIVRvVts+eb5kgB/4ry8zeM6cXkMbLQ+dEzyIrqVkIqo8KkDGG5UQ0vAcg
qLZE/G5y4BqcqQenEGeoykuwaDhz3asg1insxgVht2y6tQFxDhhXXoQxL0A3I3Yd
Xj+NZn+lFy3gSJsGO2gYzA+GDjW/ikm5TkuNrwgvb2oTpgWt9p9OSkzN0M9i9ZJ7
wCJtpseE7aUYvGCzt0JYBlsTkzC9dJmRvAHosZ9Bs4pDBzDRQ1NwV8RKH1vM9cl9
rhrEhFStFhgiiPX9g2ThKBhczeqOFpd0aRmGO+Ew6uuXB6B4BSXD61XLsVRPIox1
rnTc8EHUamWKffK326MG93B3TOpw+lsVTaX5+4AU091Spkj/vAPa08ZCU4ZS5W7d
wIR9YsYKpTnNchnv4FDQF5RzggZY+7TvJqi8H88tZ7yMHsmEjclRKY2FhA7tZAgE
KEk7S/Wknxa7CvfDEmR59OU1SUST5x/LfDaZOiQyV3XUpIvSkFtxqia6nUmJVOrF
/QvVncd5XO53mYCQ3U0/UA/KnkH7WJiPHGBRDhvK7Iob/wAPonAVnjsI1n4UlL8a
faAB77pvzZ/ejL0YDoqypdhCJOH94bb1OKhKUvoopngfWvsYqGBjqY1oe1edfG+g
l+1hUnn8IVtGPoQDg/rmM1x7iDl0oCW5Ri/D+2sjc2/1CmoAKVRxaTDEZvcQ2UG0
8wIMeuwnDL0B59UAqya/UiZ+N5QNWO1ZzngAeU2U/hl1sJxbTX0a6z+69GrhxfX+
f7W049VFnZoVkJ9XqRrZ0YF7DBkHiN5sdu5vKXPaA3Va7DCCPK/8HqGto2Qs7d8i
Jx3ExKTqVLgdO67qsb5dCRvB8K0wgdAD/N5fwMIm64PenjGxH+lSBJ8MkfOvmDNv
q23qOdb6Z9Nf3jaIC8XGIhA/C0Stl4sfderZvUZbGrXO1e4feLfQJP+tKCqQi3Bx
jeaJVvG6CITZg1J+OneQrcdmjEo9PCfBcvPJmYTsGDAaoOTqQVyoBcdvSnBUIfT6
sz6TcYKEmXjsp7iPg4YbY12MYBG8rBfJWh7IGl4ZDhm17Y+aBcOxoRI1tGre2hZ4
37Z2iRtOkMrU50v7njnnaaU5sIhL+wPsJP4abKvHE9oo0Xo/8PmwT5NGUsmq2QKg
UjuuDwTa9XNz8NuAyCIc5+bTv58RcyEYaj14AFCPZ14nZoQ9gN/XAGWxWId5+Isg
11DMn5PxHk0Sptksel9H/85cP2IQT/25g0XDi/oqnGnn8Glz5GMEV93P/q+Rj2Sa
E+fApTVi2aQbn6JJVLSJlMBqymRHTEjw0ddKHHkMQX9qQLFcHCTzpU12o82Q+sIx
U85UUG4oGa3wv7KokctnlyIPfj+HUV8eMgxGjY6YKhMmo5ldg9PTYSnCSBWHAs5v
mGA1waT98B7xZQtEL0qJs+rDK6y9BXsRfU6gkXUgiHk42TGe8+Ge/EDgtgoujYfi
OG2vm7a6YRo0SHC+1PXar1KuJnKKxFC5+KPto+pb3arcdzvYJZ45JJdiwRpwY3uX
VnsTO7ZxRXytRvZl3KgA/uiFZfmFAZdRHMebtj1rhlj52XNaDYYtzWmePsMydFGN
j8W7pFuSnV12k/aAguJEIkcP9mOvjR1ZMflTHwS6WyYPD5sorcQq4/dJgOrYmUOr
h3MAeD+lu2E+THMakxnuS71BwDVgEkdcJh+zbBFZo2IPBCeeqiv0/khloxt6fXXR
YHL04D4jtQSDemiywaySTxX+OUpjio1acEC2EqDa7k6aIScgW3KKn+Xr7Ah5YArV
EMqfvgBtjbi4CXo0mXMrjyz4Udt2z7LSUh++YYrR/m8WN1lm7uNB4oeGqXd8Bjov
Y4XGK6sniVPkncEP58I9cAVhY20MfhytC9IB0J7qnLb0Es8jvs4pPCt7L+Fr5Bqm
lEmaeZyOD/aRsCZ9LqDie8XbyVDH6wggAXPRB88Ebq3ZX4UR9qKwKx/6+PSuqiYk
b+jdZKB1rY782UFhTXGdpHykjOys/H0FLUOx4G/HpF33yqO6mjEDjAMEQEMNtmX+
ZzWLG6aj8/8fW/hCj5RgbVeCP/nY2yyk8qTex/NFL1lXTz25rxxtxbNLcQ4eijE7
z5qualdxdX2rfR9CO9D1QA9HyuOwKfFgvAc2cBdBsH6YICzPKCmEZq9DfQKUgn0W
oa6mUVGVK1JdL4mVa47ekb8Aew6b3RpfiS2/iLcydwpfmPkkxE49IrfsAudHVsNd
WFzjp7E1c5q/7kam8NX6KzQDI7nZfWNqASaiXpQlizmhBK3KJy6WDUtva2K3mh3K
kxUX6czVOzk5hZ+s4KvN3ZCm5R71NKaY3CNRk0ExT6ECPVCTeveoQOktOvgvluDD
TfPDfOw1dlGLnbnjYx3h0m8Meow7OX/weKs2gbSnWqRz74uWIT8kyGWK98mA8ol9
pNKFWa/trNVh/ITDFXwcpA4wI0cjhN0KhyQfThZ0/ldJLyYzL+Xja66UL4rqpCAo
MahOgdQllKHPSc3J3x8BRTzkt5V9TQtfscp/9XqFwomO9iBGyOEyA9RBFa/TM6st
WiavweV6jGEXw0jXcMroop+BKOhTNFfEjbKvPCDmvu2TWuY8/HJ7KADxubVX/HqB
10K1hOQzKHcsDaGrRFcgmcmLFGMM3ABWysMx/AXWayD4lCCFVpGNVht0yFbtQZSg
oHNbC8JPPB9zkrLD8PCRlcXGMFcifcSD5UGOzK1Az1EHwmSDCeJ6vqrQC5r78SIb
aXQZhjcBF3iM8f+OvNLKYcWXtl7Hun1Gk7YmJpd5AUFhkWpVHYrNYVl/pMIldQE9
9T9n1fNJFesVo6dU0H4z+wIUUvIv5dSz+QG6BjcEC1wHstnP7euLEp9Zkz0tAbqo
D8aKBQ9A5IsL1UaPGASMzPGC8SF67m8Fqp639BzMXtYQGS5XsW5mRVT1YAs2C0Ig
YrKf6+as+rO05UUes6R5NKhW51/j2I8FLAAw9GyL90pHFrsbDxoD7QqtBPW0yJdW
+I9w4xadxd+gsqPDHbm4TE88YKJLC0VfvVR5bTvfoAK/2tlnecbfcRzD9D9b+NH/
veqAkeBIze5UDv8z3OxvIEcVexVbLptwdmpevIEOe5DGYOdok0w+L6umG0z/r+TM
dhCjGfHeMJtYoDAK16FWStn08sNBfszx6wNfiUQ6y8VIWbrvMauqKzaEI0Fk+LHm
KNxKdfgZBYpVfT67lhYsjLjsrFKzLhs+uF6VmJNRVGycfASPrQj7B1xFMgJQblKw
8cLTaXNgGbg2BFfMxW2iSKycGUmXgwH1iZwxVf7o4yXU4egQs3N0iOrerrki4lkk
K2BLWG/ieh9NJqCEXD+ORX/z/hV9XT26wpqRodc21YCYt+avIuKK4Z+SC6bIqHc0
VSt4LE2VxPkejH5TQwyF/hQ1ccMkamggaDTyZayy1wFaxME2bNJjGgdlmA4Ub5n9
cLZFGvV0uOmVc7KkQ2zA0pr2zJ6AAPyJw0yUIsOCyJiq18z6NjohSb807HHKgxne
U443QqLzVKI+ocZmB8Nqpx9BKije4Hhzz69LPFsvZklsZ85fEeOUZxd5K6gO4PeD
7a2GqA/LfRH2WfVaQAyhcg8unvwYITJfgp666vRIUf0EZw2vTHuK9MECZUyZvOCd
neKYFBVwOOxxOsKbzJjG0dGEAMGDIZ3P9v84au81X2caTmfOE6GRe4jHXpb++YQO
OCUGXyiW/iuob/STOuUhZVUr1HMf3HDnltKyV71T7XfVP5fzhhvIWXvyCnYDGfiz
yBuf10NXjtZDxWFNHDsSfkP16FYSlRZLYlvx3aQnBAB5HdQcHUHcsktgcy/Hprw3
7nrzl3zBQVM71zs6oxj+eXMTfzu5TLniwITb+mq7V+UEiWRYhxYX7fSNlE3rCkHk
rtxhhtZvk0VOfNNWwFCKsTYGWqznJIgYvce0WFSd5R6hcp6vS4qP+LUA5eetoLz7
1qcc6310Aq+0QW97B5QQbZ5fvOSvoNG1IQNA80LGVknXY7zbjBwEEdMGMFGV0O9+
adFkrxYa7fc8pl4Z1JOoQj9ka0+BjEQIutARcww9eJgwL32cqIV/t1y969NVgBGc
CGQtoCWYmQSQHjfdLpx9qilw9lpBNvZwKu7S7PFuo8ytzv9aQUJj/bxiTnNHFyRP
udQFQlMPbOnrd3qjrSvvksTxR+LZ1BsApTOdN4uRf4Ptp52E6m/qTXdDdb7wpM7R
xMggC+kBmRnCBLV/rkFjEu56eAaq8Gjb+iaNjV+L8exzjU0QkhgeFatGfgsPk/w9
LkWR83PyGymEQxJ2Dje+DVUeW5+EzTRVF12NNrw3lvqr0YdiBLyfY71FmIpjA4kL
Y6u3k5ZDbxTUASdrVp3R5ZQw+IMa8kDMlSXTJ+0w+IBNw3MLd0DhMwy0pzkJ4WSy
EjipYGvRcBaBsJ1cfVI4FfIjeI5LfGpypgZsgdUXpMci4IlMSz37A+KpN3Bvu19r
FvS/oim4onaKD09he21ySlreskpMyyGxQNCMVQxN/Sbl/V8fIkkTBNC6SCtP59AG
bQtN5eLvqmVXTmlRCHzXXh6YenL/Me3+oX3nl8pvF6SFOjkDG2ijfLxFSSMoLqwX
9yAnLBOakoBAbKGVPswKOUUZ6ZFLsF/1ue3JC3az9B8XdaSVSNfJe6T4bi8itcYB
WR8qpmM5Q+OlWYmuvN9FpNvQW/EOUzBPdtjdel9DpNPpIymF4r3bIiVzHMYZZ5uz
ehkYluLPv1aRFZ471WjG5gqXPOfvqVJ3Ye6fgUDUMce5wHq5LB005XQ/ISIJKSDT
ewszkAxuynnSyI8Mb+rywfic+q/Byq61FJEHQZqcMsc/r4w3v1Q3dy5FN2uopFIm
nJUnc7WZhfQDipHoWEekfRnRCg2Lo3oQqaaZYaqwr305IYce+ITWmE0iXO937yy+
rN6985B5la/Pt73KT3dhO1adq6ac/gQxGymk+IRawVjgsJXu7F+3Rx9oEzicebAT
79cxlf/4NaG3pcfKhO9OyX9m2jUIBDHk9UUvHLwwY3hV6oRGF/nijbDuMzYeK7B0
oy+ENiiA0kp2ySTp2NxmExpkDqjhYdyIGPcWWRWEv7kZWRLh/hTYDyASj4GStn2P
fvy0SGcnSP+A7EKVpyL45Ft/l66QDLOQOscHj4NnKUhWNsUAHiispNPHqwOadLai
2x0llAZ5gD6w3B+zy49iH/AaauAuHtooAI62kmmAxxflJLxGDAWjC2pm+DQd3keP
o3LwBKe1bd3frpheAoc9Idpp8ENlhkpcWcVgClDsbQkE87WgxMfIy8BV4t9X9RLZ
uosmDAtA8XY2iw0b1NtEPNzj+l1l6QP4Z19+SNIlZn/uoRDjP5oZgdRURiz3x2a+
c4jb29noQUN14S4PWM++aug9gi54KRZLGtlRRHbJkFd7pkeunuyRHBg/pao4Z84E
hHKMu/+RjVBMcwKDWYsXLBUKM/A/s4MLpj8q+reJfyncdUmn3fcl1JXJY2soBGbm
6tIDUvgva7xfJfAZNQd7ENXOX+d90o+Y5w5L/E7anaZplEzMkGDbQIp18LImkN+1
V8oYjqKhJ40TrZ6aJrC0Zxc1QOJWKilPPbGJcExuTS3THyK19NbYslo5AUNexvMM
o0NZd8YU+WKMs36hAaFyjpvHONPc7fH1uj928Og6Z/gSa10cUXLd4Hkml/NciBzk
dUjcllpOVZ3Q9pDy2H7VAB3/2vjVYYlYaAZSPONTnNqLaSP57N6VvBbNw6O1jB+2
Rc57etS02F0ifPoxXFbLbJr5adqRXR8rQgx3Qp5UM4JhvsQZyiieXUuEcdbVr3+e
/5XKnTIpNGz4C7rtkmxJnlBaa5+ve+2EB3oRDlKD/wwfQI0imBZwe6Z2GGGv3xvt
mgPR8vMdodM+ykKb/iytncub55hDOgyzzcroA23wfIMOW2Mi2usm9TcPpUhEdCyM
RNqvGpF/ljOyHilWyKNV40hWevfcucPcXmOSD7jdy7G0xb0G/p26jRuRNWTcz8fJ
ANyPpSu7DDVR6CvXAYj6j1l3xYYjJoaCQCE7G79PGHDcLBLBuRLWfZdpo9Swvczp
KnoQfvKuk6rYgOVLdG7in4S/nxlVvqI9WBU9zSUeg9ZvNqbzTCRMl3e18tE9GPeG
4dWsS8tZCGjNaLKJCMSRNBTef14qNztu+adhcw09S88sfCjbw99Bdp5DdWrrLGi2
ZZKjVbE/nEOLjtooFfXJfdf8vfaGl2ayVd4R5MlZofByO7mblbocK5N/tb90hRSg
puwNaHRuQBVI1y7j09ZXW12fHDnskyCQgE1/GyLwbbRHsMT18w+rE48ZndVN2MuD
7gXtzZmHs9GDhzH7TNwhEVqbQxiE38KB6Bk1y951nhvCe1CK83F+bkpFQ7aDzqHN
10mO5AB6D5YQA/kfFocmsNcScAeoiDJzNTclg1ynWiqTHp41w3gher+hN5pvy3DK
CqIbFBBGQFaRM423Pvah8qwcnfmbVMfpxaPO7yiS4xOlQLWQTVtnhtXCtkY7rkxn
ApNXVK8U5fb6gcrQh1NFLHezKDZHrlc9VFn3b3G+0qapzCrAsqGyHCMc+vko8K6E
qyr5g4yDejKZrfeKYIl0KFqaajBuHmjQJcm0pzXF5hK42h4vVfTTCt2QEDYEBrAr
QoatUbWOo4P8kc0exA1phYt8Z79yron4vtEHiLyH1jup5JVMFBxcv7dadzORlIYX
604XLNMc4E8G3e8WUqS2QU0BtL2HKNFQ5HAu3VIyklmUKp02Fus29mXjyO7syH3H
NFv1d39o+31Sqbnhv1A9X3yT2nmf+60hp3d6ggofJka3csMgQwx1UB6SaS03pLhT
NfhmLyhf+ZcaDec5+XAz39VkVGQ2iS+1IsRJ1Cocx+nDvhLTFNDwr+WnAUy9wwLf
MVL3vFvig8bTul9R5sq1BUx2CUPIxxvMLqzsQRGt0Vwvf+f0RNiD613+YPUQo4xh
Li5uXvdW6qB6SvQzHLROc3c+dVES2uyQc3ofpIm2d43HgXuEt7eE+G/+JHtlcMmW
OFLWjIIPpqbMStgJFNvCwaWy+vgeXWt8T1dEPjoFY5S8+DMFKvNBPXs+Sx1k5gYo
7iFw9dMz3k68lL8iVtYrmCDMLe3zHNqkRxLoGx/vMzRC3f0gwjtF7S1bZKrvKEVF
ws8Gx/MuFCbBEwIoMloQ9s+VtfJ1bCV1kf1Dz2VMIqSMWi/7zPsCkKB77LlTG+Uh
APDQaErQeqmMiUvFyAOjAViYMDREYvPQKURvqJSYKVxEhDqXPJg2zSJY5nIqMZhp
yggVA8qB/WF7Dr1YdNWKs01mqngeCxIxnL5CFAzKLfAzRsYVtU4cv+3MkP2749Rr
MxuHuZ2PVfmFIpvz0bJJcb1Kf9CktuUnDWStgw4NCTXw43qjL/OJlDdITyftE0Ho
fDXHexPBM0eRRRb2N42YPnFZpI4/mQzO6+/8bBDFuWBkWQOCgzRqzp/sRnhwQGIS
JGpIaxkNIo+UZtu2L0jWqiw/Pr33vuRtfEwIbWvlvGHrM9SC9PpmADasOTupHkok
ofTkeMoOa+1HJ4+LG4w+mDbN0YOb8FDZHtLz6mRirajWiJBOtQy+E+q0BKFqhQsr
+SNYAg2+zEt58dDoEtwKxSs+ax/YrAI3rAgMtTgKELXvnIlw+BU72b1pP+AENnn3
zCkEgQEYdA2tGi9f1KCotP+5B7FPfw8RYbJy3Nh6t3U/XqzIzKkZ6bp1FKCAZOJa
5uviwiG5l66nDuuhwBwmqVbxWmUvCirm4Ny3h1/4kCFIPZ0Kp6CZoqMJeS/MbzZ9
BaI6XgAZ3d+FlvVSFb7HeTzVX0NTvNNQG8CN2neVYo9el7iLG8UYT85hkxFpsyWZ
od7scoFYfoEYZjvJjHNqCQFFVHbmDC+Z3/MTqU5UI6VW77COy2QCaU1FSSCYLhLd
rtAulXCysn11wBK2LA7vmOt0OZzxiaCLtBfjHtcL0UEePkfFS3BUYf82CjPM3rLF
VXA4QCHbggFDxSBfsuVb2aV4TpDV6ntDM/QupdEzI+3hCkQPvX4MDxetjCi3Bi56
MLYua8FYsFj5idzcxkzG83I/wbPBPyNJGx8i3AG8azisM1ejkGYTAlxcKKViLO97
8S5ngSuGvaIxpVCJ55oHD7q0+qxs9aQ1l7xMNv4WoNZj4vL2YDmrWjv1ksSnCIej
SxnRLIwc48MGOEFCV+/bq8rfzBgliBc1IDz3LXt64yFQR7FbYSuTsTSS6TpDjRyV
eZ25Y1Q2d1tGE1UyFI0DwtZ2wj3XrWg4ZX8xS0vDJhyJnTjZeBh90E6xPhK2Tpdd
ktF/3z2UDZYvdJTRaPexNO/12Gvqe5YGBHndtXWuLvsfqjcQVDIv7r9wt0e7YBog
LwKj3DQAc2dN0fTgvgWbAF9H5Dv0yOGB5VFDB11yH1vd/ioAsUTpbGts+7PelI+L
3DgbhT9f4gPrP8XQ9dgqAFI/anznWlq/x+9Rp2PYp21iw9XoHSS3fxLQNnQXwfff
GzCgT+wVbEo42/R2miRLByOjJVNTFOHD5pJaIJfc0UWpls+rKTkFbv9MwN9Lq16A
6c8fFPckznR629Z3f7qy8LDeyj6R6Nro5ShVoZEDx1couG/aVSOqqJj0GHxICcuL
LNd0X5upacfVy/JxDYbGF3bUFFN/gdE22V17X7kbdImKjY1mhp7zdOVhTs51o+Z2
q4kQPeRJ4xFyrodUsMjkykIt5fV6Xdvpuy7EyyL6FtVh5M4GYObyJzUChoLJB71c
9j9FsVwr/s+CnyXez4seyaxNnOz5tU3X9DuC3ObBemhP2BrQqyh0mqxIWlA+OUlW
DwSAUNz7BRvvyENA7mFMYpg+DMQasPFTFsOVjTaGngsRn9v5N9Y+hKSYoNn5i7kL
jG/wuLYD0GaXet10ChT2lHtpI/XEkc9OKryS0Za4tuBZ0zvmX1fUsx+MSB0Ez+2/
Lb2MvaKxTqTRSHLMg0Qe/9f8Zp2r8gRGjku94iaIh5vj5ZF0bBMfaEDVi9w2VQKd
+OlcQp2MNRqU8c/NYomJr7hrqWP5p37I9sFCbh7C0W4lC8CCT/89y4YwZwLgytiy
zMSH41KnFWguGinV9DOSKGBXvozGd4W0Ecr2Tnz6QF6ubsGxzV0IObqhDD6tYk+G
AqdRCsVYmIdGrp51Iwr/2VOEpjvySX7wGehzWfHdbS6Yz734qYi0mlj/498/edpt
1L5I/XowrAf1LeSWH6zFnYitH4iEh61Rysiql+YQSU6OzfIiFfcFsw+4VmBp8f35
IEpAGSKWnf45SUzeUQwgHbO9vsqT25Krgel28gGvryUvkBtO54x27G59hMvsi3pc
zQQHuZWv3IqPomGAD3KV5AzFzcKbKVOGVOrUED5q4PA2variVd+H6xa38WpHVuBb
VNGZq6Ud85WQ3hfGuGbK8l5JLTQlQaTFbWacz/tVOCPlEavr4ql/gQRwBbmx9w7z
FswtNWNhc5d9sOGfMl0nb2CyS5RH71VRfjzn49ryHx4WV4HOCP6suVl4B9MNvk3e
SbUtvC9aTWQKkGT41NQWXdDfA9rhLHlzO1K6JyH7Tf5Sbh7YWNxsl9ljUfN02H0j
S69+Maubn7PGNHozJ/OGmlD1hR+9tZyBNbI/secAa+vnqh6pWukWx1rDfPBkNcsx
XV6jCxp0Bsn2hWsAY95xqoCRd6tWcaXXDrsSeNBTdPSsJ+Q0Q21Sn8KrbYl9f/Zd
1+EZHQYWVWHClhbgB0PD/sJxIfHy8WPptDDeRNsR3fEf9mW+APeelAbdAvQ41/0C
564inlQ1Vmvz52mHJ1hopnepPK7o2dOU1rYBSN06KY+6uQO8EO91CLyZxzax+Wqk
06qwnC+QyQJBY7wiAdGGkJhrOOKpNg9SD0PEAfbygcwoGjFQMkNA4gVJzCnkfKBi
k7XV4Cl21fxCvxo9j87ziRWvwGc50IG9cmAc2PP+LlJY5fLlM0mAMJ31W1JRuS6D
jaGk4CyWmQN6DViECrGF6YKB/lBTNmbRjdq7HOSPNFbtRD8zylCv/TLwcQJtJTjL
TBucye+Y0PBL/YvCXdCZyOhffL7xIQ5CWC2B2PXWBwipOEMQi55VQ+jwEvCQHgQ5
umAREhjm/KlbdFDfdL/Bw8smlQGGn7IpS66YI92Q1H4K269nI5oYMLulMJxLrgh7
ob90I6GcmSWIOaV/srODWfOxupFDkz4BWGtkIn41o4GG/c3YscbudV/RL4BIIjm0
DJ3n9e68my41oApog8YDCS+fi/W42TabJBZxx7NFnML9qfLn44Kiy9Hy8aF/jlao
bXWbrYXs2UAEgcPIwuqQ2aQOhO0DI4Y3XlIS1ciEnv/Cp12AHMjLE+NYtHmO3izr
3TOVquIU+a9ERPcb/iXOnyJzOttUystLdhQvTcLHKeoqPdMUsn26OPo6R5Ew7Uzr
WhFTMSQjI385zLR+FZM6g5c+4/IPYydZF4P5Ef8+lvthuqFiX0Rb+YARxdKfFBak
p4vSBU/luxfLIa1G6FyZWE4g7HBv9idwCGTZD3UY2Tem2p/cTCI/CMGGEZojfP3j
zKc2xrW1/FAA6TWtsdfebJCyk3xr5MrDybkJJ8+rQy02Lujl5g7ybPhWinYqqRll
Q2wdGsr+rUyhlK0GjQDQcc4s+EJxrRtY69IaHKhOXKI8q35RjSSf1+rnVVHYCDgi
1NdPOolZGMIAsKVfGSNJ22HmeXhZTPEPZu5YGcWZ/hkmhQL1VwXdyTBAB94vUpy8
3EX97I3dXFmmKHMMp2SGbNgztT8ur2w90v4+PB+S3PAtVfjlUbxsp8ug8kc1MlNl
p5OjYUcVMEvR9N9nisP19z4jT+TCyMlujPjKBtJmf6r/6FkM3iHEHlB3lgG4vGTB
mR05PolD6/VJloA12LRlUkjNOyfnvNVEsH2jxLyIXPBQz64AvNxAld/fPuYx1t6m
ERsZ8jpFUDk8CzPEXt/Ko8yeSKxSIotZfQv0k1lJwfo1JJH9K7A/EzIMesWUa54B
ReBy6uAljojxbX3pfe3tyEE1f0MPEZm+MHtbz//cGFIj0s8yFNLoMFsaMvx5E97J
MG/zwI3HL4DEh0Y+j3TzWIPH7G3Es4VrlKJa6dNuXODZPkpVpucBXZ7AW1QyAVLj
M1OzGeFjme/2xzLwvGvo2If6RKJxP6JDHc6F+P6bTIpBQZJ0lyBBtE7l3/u6QpoT
ZdOn6sqcxVLUSXTsAexCnx83e8thFRhF+GoSpVZ7JCHafQVaKRop6TXA4gf/ssNg
8nHFHPdtT9osInBlTZAkDl2Qxked2pYyx/Ofk++Pz0rxYfpVVNKq5cMbBLbjJ3FK
gKrelyv6IGVixhQS4Q7dwBlPcWNAucqkfaABxEgxlMOT4NU8CtBUceulTK7qIWza
2dDnOX+6iyv5BXdqKJZnx654BRWX3lGX4IGzMhNuuYF4RQX3i/u7kDwRIk2S+Xv7
xv6mHKnkX3Y79dOhPMdZkeoXeawV3cAPI70bWt2yDrX11HFRWZ0Jupnd9qVw18UJ
Jyi9e+fgaBvtU3CaQ6Y14n8U5YUYDqkc35P3yz4Tn86R2sW8pZMoDlLzFCCRA7DE
jFkVtjtzCXbJv5P2aZJzpH1kVp3nPmSNh2jy63t31u7M3kFfPGYsWQMt9+eIJ8op
Wy/uTebiCBvBtstjFgwuoj0zu7njobnfZXVIhN3Q/iOTiRbUD/BiGMJfB2qUFNkD
mI/4AOMs8u8wUzhqcxbUvfSYLdy/PxZ8DV2UtvTnzkMUZkiJGlOLiBpTYQDpA45q
z9ani5s/JgocZ2LCA3k9Chsm/cTGpqjkF5NhOp+VsVtGqqu7uWIa9NN3dN+HsDbj
CilJdx2oOSy+8B3MOGF4Q0LtrfLOloy0gvRI6EGPW+bthtSyP9UpVzuNtietFNpm
sNZ8oqPxvSThmQGJcUwujHWdN1g161uIW/hOYvbjia/SmrR+tyEwBohoCsJhTCNu
3tKtMxxd+CBvKbqq38kaGMUmuZgc6Y0j8/z06BPgvUL/w+V+Y7rYvH1kJrcMx52y
J7DbOWA9kqgmgu8/mSXudij4FKogtdGErOwqye5LkA7tIwRYkex3B/T/MOBo/bYZ
p/xwORIkC1gPEOmgPzkx2VXsCE7DbHh64CYY3n48zJQeAAfWzpIeBO7EWNq339dz
umotMo0GR5jYteP3Ukh9Y0sT1CoFo90uM3dO/rYYdlNqLS1XEHCj3q56DsHPSLVQ
d76pD35bxxGHZjIORTS16+ejJYJ+NxlolYcTDeO9ikPUJZYmT/c7HLZkoc5bPswU
FcXKx7dWvwhzeG4fiEySrzkDnFG+1ngFh70AxFlseAsZfRwdt4n+cc39oFzh7X3A
g/9xxFywFmbuOfki9/SiTsTFMG2H4N5HPE71pg8qjOqVhcY0N9bEY/awPNowLxbH
aEchgWok7NtV7LZBebYgcMZz19ds6PvCZKetHmFKhmHGEHi5ZDYioLtP4jc+KOa1
i/0/WL7rSD3PdWOJcSp/ecxiXO78gFnd7xW6PAkxj0pp6mrXhZbREszZxBcVaMSB
HX+v3mgVwDvzH4Z9PhraaJAsl/VI0rpZI0d9ce+cHt/CAStgckKsJH91vzKdup3a
31Yx+Zp4kiO2CBQxjb9jQl1mkUz7TDE+kr6/LPZOKWIfTzqUW/fD2i2WaqRHLQoz
4MNcoH0X4bU+pc1gRGONLFXRRudThWfk8ZNpP2lee3VGg9QOPj0nj1fMCO+eG17x
iRXdMCt2hdbDdKhzNeKQgaEqmW0hDPuD0cAoHXlkOW7aOsf1oJ5Gu5L/W6tSJ14V
UKXOMk2kdUKgUalEhc+T+VpFAEbrU6y84DWo6Ihs9EHT/3pABHBKNP9Ra8nF0o7I
FDPYAI/5Z4bd9q2poOTyDOnNuwINPiwdX+P6DlGWuf85i4tjRvSc+3Un98ux+q/J
zn+xEYvVtVHyB2HdX415STlBuahjCd/kOt22FMa9NJFIa5vX+YqLVLj4bDkr/PDE
UcOCtfVJv+HSq/E2Z8/XBTagR4FajCS2Wfv7KiN70g2R9hTir1mjnqM3Qh+D1E3l
C2DrszSMN0GlTTZ9s3XD9jk6BiWuV66nfw4HxJWgasGenS9th0OwG7/Mo4YFsRkU
fWMxcuMaINTi/PgDsAYu5/EehIU5iWXBG5NxLIE79DjhkL8ncptlE9GepJxQ9ICW
E0auT4ip1kH1i8JbAOtJPhf5qS5K/dvRIp+Xc+yJZp4yGE7NSTWo3frNiiCge6pu
Cw1PCfsqmIZHx9EjNc35ow5+TReFalPcyqYO0CcbQqXhj4VlH96UDqF5syOB5scx
Axj8DDXfJq6SEpJrIPpxupwPw7db+nqOKAoawJ5S3ga//5eXIVLLFyjS1Xdq4goU
Cmc3ANWbWICKUEV8auaar5NtrA8Imhot0s9evx1Xhzsq4q9Ocgn+kAVlmF2Ettw+
X+9qrnk2yzruDQPtXQAS/Fao9fE8mE6lgoGl8sOwOmvhxsk3IMiNJ7f912jXSyFc
d/dlMaP1hZKKr0FIc34CHxlvpSzdnvl0+8hf8Z02iZCT0gBsiytavNpkzCBihWrj
iC/COqIbdVT5PLUMqQVFZ3PANhwOWfMaNtT5A5zrD/IdmpMZO8jPMuImVPUqn2KD
TcTb8cOjOzcJjU8YfOJaEbyXjWqeWYgW8tNYaLArLhk+LfReQsKjxU3XB+vqkk8g
VfM+ebO05bdp11MvgDryiw0M+qv9+MmhUhRJ3XJj1ner4AmvMBoSFB6EZIDVM8md
xP69v5Wpk0UVA7fcE9qM7+zfM/85VTNMWa3GzGk564nc9Ic9uQ0XQGYjh22QOxRo
MJhEoC5dLa173ADSMGpENC6MkK03zfm/b+4bqrvS8QTm/w1YwtySl5ohwbhSwU3V
ZFLAj0+FF8NyfJyrr1toaa9WyZ92DesjEwuWRhIsHPa9MBJHHhnhGGzdAfJ+xtPJ
2ZBQvJARzXg0H6RxZmiQqABkAA/eiWvaZ3TDgWdDfg5+wCeD0iJSyAK8+rleKk3I
NezW/SvBE+eBrvEevPMOh9rGFQSucJmMDHers9/rotVj0L4qmYFhp1TXl2ozkQJV
SQoiBctAI/5tmfU9S2M1B+75vjZX2rEwfXvHIFP2e+g/R9Bv5qq564witjYh7Ki5
ZeTwW/71vpkzniaFRzNwNqHGD2wUHw1XIcEDRnIlGWJHPH/ROnMi+zcVD9kFxKTn
g7cJK1Xc7EgrJXAUFIaHHe8L50A439RosQ9QHXyijYwXj8WO3EUjM8A6Axgm4Rz5
LUZBb1NfWUMCT+43Q+iwmfDSlmsG9h4B71BRcI5zQlDUT29Io6ScEbfjn3Swg7JI
/SRrJJyqwojIsMYXnDt/m7CvuRsRNeC56w4ubt6GSviGSqK/Zw21sJ1Wy9eskVei
pUl8PV3YKlw0yNmL/OI1gutkPWHHD3Ocho9f6+Bd1COS81bCQ7p1uNyk+EUZ3iGc
8POeRet45Gnq1lgTmtFKjewQaIE51Pb3FqgS+DCcK2KZK0sWQuTLiFuCBbl4xTDq
uxCeniFmCsxws1nrYHFkzs9PRQw+amU8gqKIMmGHWqaUGhuour5bvTiXaT9w05n3
z7ATJ+rpBTrW1/8Egl3hpWdJLx1BFcgsSydr4xgbO3d5l96pp6EE9vcXSH3Kz8tA
jZRZCYyIzaGsHiKm6fgFEIb5/4fp9yf0Gk2ctdNtL2wE7Md5a4QHclkEOvyf0YCA
zce2xMHPMNmnVx8c4p1/Ew/Z9rmcwaimFjxRWEYRe0gTGseMDhHcPnVBCCNa0izd
w/Nx8sgBz7Zr5BsSQsBlnZgDDaCL3G0WH+PKjc/xLuWIHu5J0zU0elGuiV0Cq4mW
B4G7/tggOyMoMSkBQaBGE/NnPJ9fy3HyWqOT+ShsUxIIjn+F4AMXRkfV6xaG/xx5
/b40mOIiP7gj54frTUn9L7qRboGBa/rHJltVktxdmWVU4Y69joVMWiWSzdexDP7M
QmbBlrVtcYfSa/ZJq7/XIi838ez3ejFJeaJE9ne+yOmFyOpgpFyj9E3QbqrZKamg
5Y4cJPk6KzvwNhX4UxtPLcPHNRAU+BfG0cf1/FSsHxLiUEqVrnaWllbx3DTSZhKd
7lEII3xj36yGNfOhtwhzUj9H1MzJmkAhHPK+Xr/jdzVqPd620EQfRqOcAzTyVh2/
vkdJ9vFdtS+tQjxRQ4Wc4txHmT1Sq1NUP7aEns4am/OBv+yuKzCkQ9V1mSwBceRi
XHuxSQg8Ow4Id9ybuQzDV89t7QdTTZGCO7OT1TQBvCfjh86uuRHG9DCWq7RTdVJA
BcLtIvpk+aazKtMTq1gouI5MbmFVuBlWMrZ2TMPb5XS/o3r3TRGUSaT/4onEVLNL
IjlGqyodXp8qKKu4tZ5wWnEWhMu5xEMzz004p/ldMcuwPQRagjd55TT4sKEAULl1
c7pRGCYZpXnGS5EVwcBnyTClV14d8b2zpaZYK5EZqgFV/sF+9j1oXHrllSdk5Kqs
6L1sSUP7TXOuGy6m8DtswThw0s9k5S5+69a1uZPIjanS9qj0vAB9NtUk+wv+vXsW
pPViVwvvJujaiSUBNJxHDLjn8Cgd5bT1nP7D8WydeU8xfHuL1oxl73JTvn8ZoDJw
gyYTXqkmZ7l/qBsbjnnwUHCxpNfgdTStpU8Pl7IP3b4VjY3zUDeHiTh31f+ZrQox
v8/VnEjIaw+rigPwDLr9OwlEWaK8P6Kqm8CYHfehzAQOILRENWSe+PI7fKOYSBVp
iSlb+Sq6JXkHw4fOrijse9H+0V63GeUd9+IPlz4zJqXTjXsKPpSD0RbFR0ZM5mJv
NfryBBUAIbIyRO3ebRREM7KbnjavTD94N4afTiP7/BxTBPjp4JeI3lTZeVhznYQB
gRrCTqulDY1Lf1rRgKVo7xlUxmfMPveRNTVMHvOROXc/o4Pi87O9Qsz+ds2EXuxg
UmknxSvmncwaF8tGjIj6pKnpIRdBHpq/0Dnw7gGr00Bf72xPsIjcw31CZvvV9cbD
dXLcs1oQGHbwIEYvA3PMOysLtwdDYO4drMw/notGunXKqNSNsL98VFNmUgHqocUh
SujQkmu53Hnm3W4icUKsk/ipSUL6EB9qniNVwY0ZuT14CvIPo8X559YIrg3+mY71
Jhw1DawsTHWQSh9cXIhQvLhFRThS+eU8XrjxKJes76XWbF86+97kw+3dRS950i/F
xWKwpEAQjFsRkjDi/bSNPZ1S76GJ6l4IHdC8jjScxhx23/saLWIsxoWk365lg4zP
LDOe7GXBjcrgMwFvZJ02h4AM9Q+3o0tX+TU0SZFGSAXvpdfrW31Q/l+RZhHoLVwq
37S0Pv7/Xn9knl/bPwjAwKIM6UOYtKuFC2PsxStk5kNccJYzIcSecPaeK872Ujp4
o8r+NDtSKPwa5uFfy0TN8SSUQsFmDSZ4md4AjHxMp5tVu19fvQ+FeSP4O7bNmwKf
KfiPxpEwxFe9tN6KzSQmDTodzYUvo80cZX3vh+EBV+yY9aQ53Lj+/HoeHjLJwEja
IHUv+0qiZ3oeaKiW+vsdpkdstrEMSXcAhBoenj33Fpjbb+O737Bcsl9cRDW3o19h
QWshMHHLNrbArwQW5Ds6NPBSfrOmBJuac2wHaMaPxn7jWuKn+aFB08RA61VSIkxN
3adhii+0X6zAXAIHJBgPS/rSQPEquMBkF6iHsN9JhUnPhQUvYEou4Fd0gegp3dg9
R7E+0dRoNzN5MaBYmgi0HdExutS2sElKKAF+Xlze8TZy+OTeE1GsdJza875ICw6v
6oTo6+djGG/zg+1i2J7BdiDkFI0e9eE49K9yWC8Pm93Wixwldp0YmWq7zW+dvjp/
ci3vdz0OuqgNvU7Ad91I1xX2RhnpWb5eWYQ3IvZIwVRJbOsCtlbEGIUsWr+inb/7
C+Sn2TY0FtC3bQV9khLe4cn4nlGJcbUTEdlKUIMo3zyrsC4fdbe6jyyoQKuKc1Li
7M1j3Re/eq/DKkIpzLRsY9bT1G3f8DZGVtKRBYUl9YvakMq7UnzgmJ2wQW7vJ9yt
P28/+OpujsFLZYHaCR7YOR6HimUKNJ5Vr47WOC4jLAeKak3dKljuLfI7It8smLF/
F8xnLyfoQnJar2tee/IdGjjvc0w/AAwumP6WyYK9XZBf5D/41wX6ZXvpF8BdsrWP
GjTy/r04Xg2oIn283utFt1TKZCxMtQcLSk4DHlWOwG+gOWXonBdRZyz+3pRnHaHR
QKFPQEwxHeuTy9acpgBhDLX0ti2dgjfiiq5Nr/3ck2dIebF+/cMawHO943b10bTP
SWt/1tr19P7/6xuXC8k0ARL72f6LdE7sOasaN6+3sUAfWtuIzqg5Yj1n0HoRmU97
x5IqjtzfU8ihqwqgQKojRFm/6SpNBNej07cZMCP+WlDZB43ce7U3usPx0spNmtTq
Tuws2TGcnA93WzAIOWaIChTUObLrtKCDyof4VyN0Nt7JyDhSKwIMbgfSUmhcKjKg
0f+c0wf52hbCG0RSMIfIxPPf3VBQgOEyk5DygIn8cM7briXKnLc+ouMrEgkK9Dvv
DjBBtVA7AVNer+2bhXicq3ZJOOZjPnFJSjFxfaUEcL4NA1oTdqZly9a46LQfzlNr
jGlEHqRsGJZmpnBAE3Qh0bDirWQUwuAWF9LOjEfBNrAFo979qTMer1ZyxXDMLyoV
M4GLKTFx0HlOZnLWV/FMpoqdJJLbMlqDx1Z5y9xMBpD65cJbPZUU4ExIEilnplST
V0Q0R4xjDT6GEtrZv2V3rRQuHrhxm/h0PsPYuTXLMN8iQtNwUasiuiNHmo7/gpN/
8YbueG1NF9KEa8zTlYIHWsMV2uH3xUl2UHybmiUQuwGlcBOUgcdZhXt0uA4lMgDI
8vNOcoaDYcqUQSNjY/79UcX0hAx6lJQe3Ca60aeIPGZnLRXUxuKCtQ7W6fuiMdM6
SlwglD4KVCA5eg4kFtmi4XYxsEaqnUIi69BFlamInv+nD4WeKGkg3fAjZYjoxtkx
VGR+B2jhqdWw3K7uX61o9zjXk1AsEDHEbDDO7XioHHw+ipiGHYMsxEeaqa2e23el
oS2Vrs/cd3lYwxc3Xiy+RjmeTJN5lAj8KflCh2m+ntZurClCZgAaPS/oiMNH8+pM
sPxwMQ37qBWRK/h65bKCtfVNFGTajwj4aZ/0d23LSMbvvpGiqZgDGzhzi1m3jBM6
O/8TRrPSkTPMLYSl2zeOvgfJXZShxJiwfySypY2HmvHeSiE84XMyAF0aUn6PBTPa
muK+NLZeBkJM1/1kppNiPAoxGlWYL/U9SZXqcAcTn11gCgWlzWfi2GoeR4tVqz8q
3C7cXmnhJs+TttaCWuG+FphJXxxJcr2XNGgwEtLfn78Tbj7401/9Eujkl03d7l0E
iFappvSkXnoxBptUQkzh63+9EarPw/I+JXyQsW9DEgJFQ46jbiPOT8gvpPC0VdqO
D5Ldx5hggUCfM/kp8XN/kgpxE1ni0fFX7gpFo+igcK58d/V/g2pM9Wi3X+GX3KVv
eH1m6/Ov7iSyQl0ICw5lsHmQrqm7iL+FAr90MFw5SIo1HyFR6F4RreY3O32kk4kP
0DSX/pjXzbfAzOs5+KDTIPCUIapT8vIiH33jCrkER2g8pw5Y8EEgiMLbPYypqvPp
EomGdmGvRu8cXA8mHccLZP4YqNULtPb4KOhO2kprkbCMzgKNf0bF0QRf9YjxE05q
5g07h0+UxGjN3MsG0SAZDvJAX5t5cYlTN3oYQdAlLy3zFNq9AjW8llW/F+14RUHH
IxNEwiLxl3UYEVKwmkY7bMv1kL1y7G3cVfi3FX+jBNImrrVZbPIh82Rmqn7nM8uy
FBHSgbVEWQRha94IYdu3V2GGSzdGMVIk3T6M1N3aowHag25AQPA5+P5s1YCN/erk
XMbRMmHadNrKoq8MxSAtLAmx3quQVT6CfKUX1Ln5TIXcxPctnhdWlwovxW11Z3hG
o2YPvvMjj4NCR9tBJqHKflKBXGEKeOxFsRERlw0YJ2jjEYFJBTCtIH70ZzBjIKjh
zjCeoS5Z7cQVdp9p+b2fSX5wV1CPmHjdvk16FJQ5BVLe8IXZxYX1rN9S87KsNlDm
b8gje5wE/ii2XSWEYoSG5jZXKlCUlbvlaMC15HG/Eoe/OixHzZIAUrOnYta4K3a5
+zzBusYIdl7vUn0HdEalW1cCFB0C020iKsnX/MAZu+4lgUkeKLQswZKc/wYEbqn9
fBBdh8gfusDsLZJZvYvCEuF3EMSoj1G4kcVtEXzvCF0kPjvG1HCYCxlhnwKFsvUd
MdSk+J0rMfrMk0OPX9/bSl7ychqr7fjd8+tmnWn1QX06Q7IDja//osMSmh8IfSQ6
1h1JD3JpgKLXQ5H9c/gKFW7NcPHpOkR8iu6D/1j3o99AtOBQAM7NtJYyoHSRlQ1h
RU2BG+VdhKc8I4xYv2Qc0SGaNS9kNmfCDYE4N0c9ZO2FxXtz9kY6dgTlbq3BGWMl
i1vJrYK+JrHV6dd2fQMPmRI0txdUR5HpZq3sqt6Ql3nCL1KlGJ7iHZFpousCNzm2
65z+arwpJPxD+xxC/H6qrsUNsbBjcvfrvNBNlATppoAUpUOJVAC31uPwuf3jsumv
HRx9qPB1a0xNKiJ3HkqLKo6pHCDH8QTuF+bz3/g4CqUE6FWWeWyMbDsibfnawShs
QH6SgoPMc5BQeKG1Q/EEo29W4jXr+IWMNRgPsfktuLHvllHVMq7EwSEfe5GbfBbt
azIPYJ3nPHKH0EVw1Qt6syCxwyRM9JnSNLPjNdvD4i3ECOsB5NcLie0Bri8TI/+V
nwkonLnMiYLpS0rNpmIoKpt9vrItWa8ocI6GuQqs1oTPHTBHH16DF3Q5UvMrTc3x
0igPwWmnqqlMmmIE++3ew+Xg6YTawsNN5YJp4+jJWQ+9nxlcJtkFjdqt3NHW9f9z
JgYRmBqq3Ca/1aKc5R7N+r+J9nIyjvBffPEGjk+AHugcOfXiN7m2c71//3P31+Ot
L1t6p1h/TMLevFWHuqgFGTwTnNxjkup184+X2njj9p4x6DnwNB6I6mLRVVfAVQ5c
+4O4lgQm7FhwQ6wiKby2aTGml5gdFOhXKWWMrujlaurJSBYFlMb5NBYiE70RbMLC
9zBfqwqenvtMkv96sJDBlr087Wak4IX8feBuCW/MopDq58/6KvEUDDmpuHtneQ9g
YrxEFmAjw9Kj81VWCEeaMJ0oaHdZnmRFfjMqnrEMvnD/GrY+GousbYGFMRYhlGFr
uV7ZWfA5OQ68d/OxtYRBPM4F4yGS/m8Ngg/fXupP8TAT1XpahveA7tYlAs93wu6i
Wgm7rpQdV5WOdiehG5dHlOpKYKp6EDLenylN5opLHO026mkSs2vVR0tVjPbRAcpn
estzeclqFEYsT9yxC4eUMyU3CaVPuE0Y9Ura+inAytWNIf4dCjQr7oPmNnlH4E97
KPOjNy0ykyUjrb6m2WV6CRHnnMqW9uZg73xiaOQAEbr9LnToSFgIqEocnQtOPBHZ
YA7rYooz/FwguMtRv+GDwq7c+8ouom65go58+8U7L0AR3O/Tfi00D5K5Z2SUscz6
Hu/LyvOTCW2HP6eNiHuJIN5c7aIR3KtI4QHWEXEhcnSqJKVNNuBdVQYXsz7+8jiE
dz2qB/9t6nhbjyLxoAGyh23EpGtt6KnBL0qmuaPRALCZTC0Fe1wglCY9iSJT6C5i
VhLpqj/PexcJ22qu4y/jMYjvYdTiWwx5pgNIY/hjIUAOxmdSpqlR8kqxnkTp6OAH
cf54vzjIg4ztIk91+YAr9200RyUJ3Eiy5Ez9sGyZHVp+Sgd3bQ8ip020wofs/Rkk
l3tzkIu/QhWQMYGir+nnYZM7yK/CdEiBV1ykaIFTZc640iWF0Kzab9tV6UJ8Nt0Y
D2RncxF/UoYS4n05z/kELCO+aVqc7xpq3oouNkg7lHmnbrrNyL9M4XUZmXB/PysR
ttSa9/krO1eK9QRmjmSRLOvM1G5nImvJKW/zGS/hKfbWz/u1hwvAWZ6aBjhuVDBH
4owpDkED4AGUbC4+myNnp7UZirLBe43e40OVj4c/qH1HfvDUJl/rMHyeK3vtXWVq
flxLmIt9SjZ71V4TlWCSgdSki/XHxoWG9lFD6WWQmSo8rnXWjVmKe/juMwqOqiIl
K1qFAO2mpEr0OdxCb+obid0B6cCmwn53h+f+NJBUzdbvQaT6bGA3VSwPLTwirVPE
jOgJyIh+m1cSB3a8QW/k0S1yAy66Q/Gq/YtaMdyf7J7i5eo2PFBGYOH+nww4e58c
5lmVBnYBtLoYRYgEtYjWi3J9MS1JWs7pkEEJNLsslndbtZzcvPzzXfjYUaxhM6ot
Dwmat1QwxnDePkuztupif81L0NYnsKPrwGK/yIjI9Q+HSUYIfLy48hZOntoHnh0w
nXQe3IJ6y4HI+zQzAj7UWyzpP6YwbNPTGU8iFKx40V40xAH/OfPSQfDeSKXgITu0
JjTAa7m8kQftqpf6bIoIkT5EicyBaXvxr0gpohPTRr5JN/mP/pSoeYvlS1l/Uo4f
Bv8kUe22YdOlPU3EFMo26mh6yMQAt/PMhINq391HAUaJ57GZAqPmHQvhQ4YYzpNx
4zQRAVd6o8/H05Z7u3SoopdcL8vKsXMtJAnjih4Asg5yVhF6rKp35VtmN8SSonxS
XwgEVNyn4wLg4rT2bTRwu07AKFc5QydtkhuR0spfOog2++bL6ye9390AUMSPbjCw
EG325zlXOUdqIMlEDRQLkUza75WBC0M9PHQCEVwI1Qctj+c1kjdEP5u00RClYjPN
HWVGw4QXn6qh1hV/rxVNta+6kCD8nyIxxec08zJKJBnyUw9J2lgpCFOWQkf3kJFE
VT7UtaSdX6ytPgRrHpip2RC3nyeovhD2/psJnCbWiWlbUQeNecLgHWjITyQjk0Jw
MtU+I+OUmhHXZbQMnSydsY/3IjyB+3frrLbqHKyxNc0o9ZJrf3STuVbwm4sUyE1J
qUY7s0jkQ2bsNrau5Z8XKgQ5hkMCF0YsvIuAn2HTHxHqxuuY9HVmivhaiZiEzpx3
2CBXYoNZ2fwysPMg8sZhuc6sIQgAa33fQOZWg5yr61sARE2OFPADlrOCspwN7nS8
XYWIdBS8VzeE3NjwCgEuMc6cxtjihYUA3uMJ66/5r4beyXSCk9t9VUTqoNocI9B/
KSBHP4ZhfsV14Tyq78I9fKsRl354cujVrOVgE4U90qppkkn778lk16q+dqsBj83W
shFtABaYQ5sAGhl82MguPCisaLiYuRmm/yYXoT63XdZX4HUQltsGRFVM8eOPF7d2
ms5j81WU1xP+x9TRwJKKyi0VBC6UamTZLFvHb1JLasOsfnaZmOdkDO1iCc/PQFLK
/pliHoT6xLGPIX2YrxQBgVBeYeHP0LLFZZ1fI93me3niUlRUz+6hJBJjcTE0JHZj
juH1H1jTX4E3kyfRKdLM2w15u/1o1H5naF82Q+2aQkVBJBbIzBPmiWFgeIeG4WWS
3pGU6LaWfz/dTzQY4Zp4pZDsJvSjmvNQOY+vd1fTBD6GqC9Bn0WpxDBvjsmwuU1O
0+4FZNGTlbPSqGpLWA7PbAyFv0qfl/pitbGiXlkXDPaVfDR7+CE+uS046O7VXGZc
x1kVkeP3zXOZKOzj0OQhEtYx6x97/O2sbkZq6llwi2XNEBQH8YArWtZ1Ov5Tmxx2
wfJFrJM3WJUjc7D8h/1lfRiDN1yupdCwHhX0nCGKD0TfJ5rNTqYwSdguVI0U6Aiq
nUxxUBoAxnpcFg9tVeD/IJgKLpTze850hxtfcSDcTHKVWnsaIhTXdJ++3iikN65F
PE5l31E7IopNQuht87Mat5j1/WbrAy3laPCf6xZqhbtHD91ZG3RyC+Aitg5un87y
eUBDtSnM91KZuOqU7aicSmm7S05u+k+1I8Fce48erN4HwAFvHoIyeZP0Uv4BysGL
n7JGFBBZIta5ilOTSbsWUjz8hj87ohBrAO2Yg322FPklzstrqhSD7muYq8u8oZAh
I3TAeHhL79u9HKegTepOp+bXrteJXg/4cViVFmL/XdHPa2+21QxBiGD7RXaRntIB
GlyrjNQUyRyWxSPOAlMUoQnjXiT+2hI5iYaE8Rp8M0A054qjnh+IYETkx9MPdEEb
xxue0b1HzG3fJhCM6fbJJVKtA0oRuZR+iujHTCQ8wRe3Q+7/STsn5sP747To2nXc
L1pEX95GCcPXyBSl96+GipMDjOjjdYeeGfyUxGheuukbk9LmIGvtdFXeV1ogWfpr
B/Di/51sCxnGxfdOxUuyW4Tjpr2zVjpAvqUfTI73V8kzJLzFEhkSR0fS5Hi5fhfb
7OLE8wlmuSZJmk9BDq7NwHmsyjXJOl92hF38wBOSEewePafZMn76qhd8IPin5Vzj
Ukdw9VhxI1kBN24hY5dPlXEyxe01+o+St/MDD26WtZyAWS0k+JIGYPB3WnaYGse3
B8EKX23i0frUdXZ66MhBed8oLRM4qfvmHIECoN4tmTTPAPZM/JUqPjJnJSmNfbZc
shD6/i1osKxf62ywzYxhY8Op7xtJvOb6ssIE70fKFtuJn6PZnvo6qyOJ0fECDP+S
Hho+W/I3FDPHGIzV0ADcvMsn/pKf01oZR+IQfDyqIUQ91eQJ2V7WrN3QbCe2i8Rm
RBkcRXRtacwAACOwX/eiSd+fmHO1aNHMzZTSNb5w6jwQaXwysjN8dfLXYyvzm2CN
HDd47nXqwg7LgA4VzRWdmiu7mafFrnzXnKRg7FWO7tlL23XJtuNZkLTVQMfJ6R4n
9Dl7Ol3hIwcrgaFcNEcnOnOZ523i2nP7Q1xjol0pLROB7TrwAnK2df4qPoAMxHm1
yVzd+KekAh9pX0QmKLa8wVzRllgTPrKY9wptCZLmD/2QAxd6FBp5FQYE59r4E0Pw
SCQyqvbVPl7HxuGr7YbMR/mQ7j02eHUFMvftrgaGbhWTJ2ftOA5OqlkfZgYx493H
rrecgfC0glL8D1kUU5grcvqsONzLHx7USpHv5HhkZ4r/nItiSMIiXxrZQp2tbRFj
r+UvpzoE1741TmTgjMPnuBS4djqrkeA/wEbLsuAKszqhqPCblxUHlqyaY8IvVNc+
YhiRNxPOYKLCNamiI6OX7BDzLvRn6ua4v2N6dcHNw0MIE+0cXZo7lzlrb7olyUUf
Nfx+Pg0rAaNL+FC5bQX5QhmWABSKdstNxkSsd/Q9BRVPkabrIGWixL6TWzLxQbZw
96PihoNpKE8DtS6YxdvrhpyHEKcJrWXNrMlreC9RmJBucWojgy4hX/qTX1mtn9O5
SHD3mJ/lNmZdyOi/ZEWu9LPOYQWFA8I9xP6PzEQSi21pLfjovZvdkYX0Pf32Oq4x
QGUpmyOsaTR3JZ5xy6jV2T1Yg7m3W7seGuzwi+YXDbKQb476uJ2PIsIN9Y6mwEHU
9PqNDENSfHeZxgoYBPtQuNxXlFz91vBdeujFCO7aW2kHbmZUDu7vb0Y+iDunBSvj
cfl5QhjPSwN6IETpLvYgU8NdlakrE3FjIgAL/vUe5CkpUoXBQLUkhxUgN+KgjBDf
eDs8V4UoRHfBx6fhqVzoq8mFV+L13a+K6Lhu1Wb4jnO0BXD8i+6FHjlaGl0Tst4q
pi+SXA8awwAKhBKx3jso5BrHqsQdKo+3sLD/Crt9trkEVkOcloPfOWXYyEbDX9f5
+VdcQGhnFLkwRLOlmnYfZnrHwDDAa5Ko/uhkxRwoVlHrhZyaXUCoiza74Y8qsAz5
f+Jt5g02IDyZGPKOLdrgo5mGKy/XRd84vH92fSFw6I581CS7AXtKWQVm1E6I59V7
dnTuER1vOpB0gfk5PTXi9iKPd8Nn2JnP9DPxu6S1NYWYEOWPkQU+Oj0EQTAepvto
EioIQJTbodVk8ChIH68FAsLXdHVeCXkHdhsVNUgtzZwqJ7QqKaAcTwNQveK8mUe5
XO+1SFs4LnWszbi7l1XIBo/euffBvMgMa6MotXLUG5aYqIYawR6L1l2O+Ol63xhY
ws6dXe/h1YKecABjY+VnyPMAT+RtRVAN/KdRfSmExCCMEjhkbK2cTL2YzDSGSqcX
unhx7wlkJ3xqi6o5N4Ir6858eDUF7EwUwHvvWqH+GveuSrp3FhGYnTvpDcsnZEgp
yIexY3XJIV1D6lN1/7h8h1kSW0EcFZ/TPYs2RuP2CONDttDfwgMveuRyl8g0ABQj
Pv9X02TdYLfznTCb1P2fT/UO3pe1U2v2rv4xrucToJ63tV3lEKH9d/9k5VFetNU7
uSh+v/TI5LEOg1PsVlD3nHv2XgFQdbb5ysvp6q3p0vW4/ERlD52Amxax1U/CrZ9Y
OesA5+MEE8diNKy+0GfZdXan9FUutf3oGoHAOs7jR4q61ZqanB1EHDhScEhzNvw5
CrZD1OYSfjOk+iGorD15YnpoMlurPLR0FBvVxgEcwshvhrS/2awTIitXW2KUs2Em
EsnTrsjsiAtKa6I4DEAfNghLPvrzfdYgtKwYYzrTA5//oi/LEu0izErupc4cfDep
mB6lgIsGV7RS4DkBg6GKdieE7T3CzFyQ6YSnz8doYe/Hvuo8RDq2+Sgs51o/i3kP
aTSWdkcGFBK5k6LhWMiZfC6iA6TdYNvGkiv5i4EHSxHzaXOnxNqunFPK+BgPwLWv
RLpuKS3UbV48kKBJMASOIvPeOUaBqk365g4GklS+C3wknq9mY9fW9krBiZbphvdb
jFwMobGgeY8NLuXxgFGJZWVGFkRZ3zk2lGlKN0g0eRk7hmxrkC0XAB6ndlW13FmQ
DoqJyTe5654N/hWbWhqiTD6sVmTCjYvZ0fuGOKOr4vc1/VDB87e5fEWw4gqlG014
uHv0gduGhc1TYasxGEkoJNmv1miAl9cCuHODYSqASdZorzKErOUKZ+tN5T3Hd5Gy
lC8sdjUsq7G6ifG84WKyqv5Sr0D0YipZeMBRS4gkHMiIpi/GKrt4yVTinGK2APXS
RceeVhwdikoPcnbOozDND+/NIj+cryxFOZhP0pgxAcewDbUmFVRz395PXeKZQsVE
+JVTJX/on71YMjz+Us2l9AhPlMKeo6M/10USPv75/DgVR0218wgQD80U0q3cbnwu
QI62AX2uhKgGGYG/sjNbHRlsFTVyw+zdm/602vDGv96b1vd3FrWLw1OnWNDWPFrI
fOeLlwZxGjrDJynEmgIn79v92xgK5icfmzQe2a1kzUmC83et7xZBwD4PGgc7zHdk
1Hxsx/ypoZN4EgIxOxHMz3Zr6Wtb/yajPYfUtMv1NvmQer12KVpzfN9nVp4iRnAI
3fNWsGBzr1odcAL14Z99iYG8tYXD/MjlrM53nZSJ2qg/FlWiHaJqMZlJfYtIK2q/
g1wx5aDkcvMspTkGP9VU4TNGlUU92ImQ2ni0yUphUNgcPdRp4FdtsxtucJfLR9zu
COoitgVy2QqfMsvZ/etr/SItTo/8KfCm5sDKaVUbjj05wkYvRfgnTzIhKP73AcuB
oSuldBnwRCiBti/iOp3KUCs0pahAcX5HCFU00IcKDEQ60AxOhC05HfogIDysOq9X
I+TPKd2/o3UUELXrp2S5oi+lkMBKE+AT5ihsoFraIup9XD6ToqhRLByiYByw9m56
xUXoilETGVhAOkfxCNuvXCFmUzUqLKa/hLQgtITMQ+3j1Ox5Vz+PfC+8OCa5y7ca
YvnpnTbto1tcWmDtgcFHVDN551a/KKPJ9MAMq+9kc8fBg4qytv2XBvXUoxwbGZ7G
J12jnFZyFP1OEWZgVEMwIptnra65wydJYGSYc8Ch5/D4DyJHOK1ChAfO0i4atKy5
dSo8iW+hjqKabhzk86mnp+/kbvJo31kzdJ7yy9h//z67KxtWKsERMa+JJOkto67K
WM0gwV2d8wPC3hkB4xirStV78STIOBXxw/OTPt5adYOTZ7F6r7tda32t1HNsWSLa
vmB8WUPqKjuzYHvq8M1Ii4c8jAAXd0GUq8xsXgv1DZJwDsZcxktjZEes3kQ79JMS
sJ5mXc++Esm0hiVOOYj4rRlMZ32SXsJoGQfdq1dZFrQ4cxgdrhujjVjymxXTN8sY
0Et7LfjglnFLaGPt3tAEmD7pky1W2nuHP905pR4ccbU5sLaftoJSCPLAm9Rz9rB2
PLM5xUYuTXfs3Zbja0FuZogpt7yY9I16DO5AignaYEghCaDxPrZkDOoj8mFfnuGT
0EtynysMDETb8LFDH4H5htDENjTLnXTgzrKQ4Hxo/GbIYMA9o/YdsGPDISmyThs1
Pjh8flR543ROQOltx6MkUr9mB//PrH4eEqdCPA8fdc13Q6q4VF9DJnn6jqL69rz5
+H/KlbEJhSlLlTcZ8ZZSzfNstFhbsoDGIq2Rexrp6FFCJHeelaWKsxyZCm2pkkn/
IZbXNGoTtVisU1o3ATevOJ7oBjIBB1y3GJQpDQA8pUz3s/2j+kZ/yssc9i2bG+rM
ASxkj3fjWwOpnf/9DVPjEGvYtiMLqA0SrFoKFoJofLQPL1yU7S3PD0oKkHsJiOPd
kGwwb2pKVGNXZyVzYbQ28Wm9CQzTzx7s1r2QPaaxwqZpH/sgRHyt9g5tb1FNDY1Q
CHDhnyLGdKLnA9gx39q21JtSaR5jafT8VUmTUd4Z2YHr1i39kn6EoMSyO01oKKv5
7amdQJvQ0W1RWJFkh5ZIWJbC+k8AlyKsHIWjttgS42qNAkUIDEwQlsNcqyfJxvBp
Q3NALvCNsUB1tF8XLWtXeKGHNptH4utiZhUr68I/s54IRSBFeJ1yrGza2ss0fshK
oouVP7u3lSQ9imBliLyw4JZDJig5i5YN8oNFZ2eoA/Q5IbIA/5lDmy7Zmujc9B5i
mQLcA3OnPR20vDpVQ8fDWh5hDcvWoBmvyqTVjEUi1YYl3JKV4cOHAX1CC1doTt7P
rLCMh1ICvTVIkapAO5SQ8pHJ8wy6q2JVYsPvGPIPygQeeqF/h3B5vLzOUvpu0oLx
aP1zY+Tix2tLjW9uVHLMNokUBMhBBJd4lhlyEztk0ujIVK1+joqxKN51tH2wAUuz
JjTVialEMtXSGot2seF7d9QS3q0jGvnmzN1KCDV3oSp8KmDswuPry/0lSyYXDNQk
vFUfuCx3zx6nnNPpau/mmuixZoNYWiTTPd/Vj88V2/Wa8ibk5gLv/j0NmFcMvw3Q
g6xQJ2FA2UhEY/hwkpHThsYmGJ9GcsVIBbB8N4GyKtnQuhRd2Ktoe4dnc7AjGCR5
/ug30D1KD5v3WNu/8mSHdj72EDkyU484af4QJ/DBziz8qpeVpYJK+M7KoOaKUlGb
d/+GecJmmHJxNIaTccC4edIHUo3HWl19oWMJnXUIo38P70jI0Ep06zBo6OspYP05
pdgqgLiu3pLXozYkOlw1iT6+zC5Dd699z12UJv0Dw3xpaUyjwDU4YB3ORe9AMhVa
m34HiJVJlxkYgUm65/HRP4hVqclNSPo+PefkMaNi0YhDxuABhFHaVu4tN0hJDJU2
HZe36DrmMzG4zmyVt848eCTgfENVnm7v6opYBSWFo0/TSRlE3bUZzD/0mtzTZuXz
yA46j6jgBjeGsE8VITGJpAfdFDAohD4riJMhor5RR2qkqihHhIaB0BJWdKN86e1h
8kX5lYLBIImoweVLsXRxhb8aRhWao61z43MfjJZAaghErcKXSsCazAezz+Lx2cY1
2B4qdz8UqeiUaPRCNPp+maUsOy9UMzY0Avv5SEqsh9Ecv/pMujJ0ryV8iKcpREBT
8N/1m401gNPj69dSd2YhVzbCpQapMFoo12IY432SUf9FehuZcaGoU+5rtDtlHx7Q
LTPVcZ8kZr2sKQat1XAl1QWLnz3Qntez4j7G5rtDFPsDVqBK3pYQmty94Pj3yAYx
PL9NLA6kwIws5U638rmr5knyCTB9GtjnjoidHwHqwSzT2rPOgFuqlDUVLwYsGWpY
YShR4D4ZMpMBIFzFiq/myzCdYXGBO+iJK6Vi12Fo3QSnDQACBLNSvDspR7cKFJuK
qY9n0CKDP8h6oTTc+DnW4SruDCJTJ7yNeXc+WHM/3PDaAnJLjRC8kmD+ZynDolE5
ZQZAI4SGRx5ur9v+dA4+zM/U0oYzZhj8dZodgzCZJ2gc6jWc3K+fG7YPSLcgtGJr
5ZH9BInK6a4SLYJepr2L88HZJBQu0sw165V5KPzi3yR6WJThYJkWzumZ1mAMSdYn
iMQyNOYvYOM6B4PRjOWKrRK9xPaOBXgAKBv9HG1k2yvCINgFELxhO7upQQFqACdn
URcXAQH0XLe5w1kE8siocnaLQxO5w1Ef3RGGsdCj5Mcmy5hacmMHigiWPLGmQ+YN
Fv6c25/IO9dLP1KH5gTm6wohV9kUgHpZyckYHTh9Qrg14OiOWTy0rM9/ibeAvFlC
UU9Uo6goqZ2yHH7VbYnEb3hdcc93EVDFffihaSVS6kwZOA0YgdElNg9vsQLrOibt
DGub1DIWoPD/1OoDNfUON6Y9JvgTExep+kOHKQLjLw1GafPK58ou3zW6Mb8dwFFc
Ja/36mQyyh3/VXPJ/8o0pV+xVwSSpFqvnhikaWHMNBcN7cmxi/vn0JydLzHfwBfP
VbFWtR3e5FhPPw6NGMNQWcFPT5FN2epEGz33hK0i8iJarYVDjk+j6raMQoWO46rL
R7yKmqa60f9ah26Lp/Tx9DlMA/G3gwO1X4IyKaZsG0ispCXNgbHBwxAmTx/MqEPX
6+6MhuN+eTWEPQe5O2DHpSYSB+if/Xyd7m2zV5BhDri4C/J+ruW5RIQXcmF3qxKL
Uz/cjbQ+ZT88COpxa6ih2/Hyn++fN9aTDkFUVxwx5JDT2LfySvZx5wy0KqYjus9M
Ke2y0AgPz0uRBJcGaNMTrXE+15K0RD1uz++UbVTcS4mrKyViCZRRr1Y7HoJr3ye/
namq3YdvkWecjcvVBkCtxSAKNqIt5LhdAh2oMvg08avG7uj11RepUcCZWDTvfHOx
0cqYwokLKh1Ge3T7dh2eDtaia10nlHx7+azDhsWoFhvLBX4Fj6EnZdv4OLLt00Ez
zhBvD3dqO+WCmOBJjpCrx+cwaPJHs3k32TChjChjD4FYByfazAgxEIfgQy4oPrcL
sOHdl180SvGvSby2pmy0VY5xTE2NT99FRvxG18HQ8zsk/iZavbyXlFTJ2LyG5qKc
2qPrNKBfnT15FbHxeYJJriaeBqzOjf9OEws/JoK5Vkm4FNRpNU4WfbvS4ATTozgH
dvDk9E3ZBMKsDy1YR/8QotXqdCsm21xtPGxVMHlRxLGEOqLGthDmrM3YGX9j3NbF
jlEjYVd2RVG8mB9mrpjegWoe7AY7yevWAd2yuWPNkatObAifrrI9dJT6EWahWKfa
CMPZOxT4djQUG8/TetJehiKr5mgIRIakz0/3o4CP/wPKJqCk/IIR0qXAbJnM1ZpH
Btr8o4Xwe49YXJoZH4u519oCKZ3I2xcya2uj3+ZJ5Qzdtsn2JSSGR4IQmbadfaLN
jlO7p5Gq5gT+nIo7LbyWoFs3Nf3hJJ1lKviHGI89tdnnKLUsde3q97quRqQUQKqU
lCvm+UFdfSwG5aWU6MWb+LUyjbeWzCQq/ZGq56+RdAzCq6JHAkF1IAlu50udZOow
K6RFmEicIga7lTQhER2NE2BRs7Bt50b36QQByjDEsRlPB1zrjTENFwfFdx2m7sTZ
Yi2QGrfmX524SFKS6XmTeHVftblImXPj1J1tcfGRwEHbrUHjUJhy2XWu0U2b77dj
A0x44pM9UVzOLdyOvgJtTelpvzb8hvG2fdfvESDqSWmPjzT0Fy/zJF9UdR0efxZm
EZiWrhmCXjGfnJcLuwlwGlZLx4rHhQ8Jhj+5c7hGDJRcK9vC4awiZ5lvbmYW/n1m
C1ocgpKDRPGbS4I8r7yg6Zw7jpJmvd0Oz7Ix/RXVxknWGDqUj8dfoUJcYESfLR6j
E+2z5HgvwwBP0uDGaAinymLbTgRk2ziAG3gMVuMIeigr8GaSI0vYKghmW23aKpFd
ntvzMSI6UhxOIx4SogDe11g3eW+Mj99CITmATLbN44yYIA+V9YqWyaviyNTas15/
RiSXnfiMwgUyybHOha4zME3cLU0Jega+5lq9lj34Yv/azy82wlzQTCUIInuyLNhv
cBou8EXtNHXZhdzTeBDbzEqArH0x2ClUbXWGezGTkO7d3+wubepFVSE66d6FHvWv
I6Adv9mgb80x2COZ8hBy3MCysn+jCRxiUTQxAc15ftR43stmU6YCIEx2FgtEliNg
tQtiywpMggBS7UlRf9POVqhgE+GmQFSBAifed/QdN/D/zE7uLAuKG9JczcTVKsOn
V9TFi223Kzg5AaBmL/zHb4Zfiq1l9DmEBrZe4tR3GSV61IBB5+F6lSStw5e+pnLI
qLcRS+ys+4ki1dfTVj0xT+EpGJ9INP8OEMiADc0OHtkw1+7Agj41YRg/t4rU0coh
RMtVlh8ZSrs5UOwSq/iphBHyck0witieXdp4yqvv3RjLRu1u/MLYVkz+wigiDkZx
M3P2T/+AqIzpRKD0J09+Zv99K6fKYDaRG1uAe7eUdLulfH/RWvhjGUhfEyygTD3w
owFBWP0c4ku0oLaElVTuqBFVK2Z7fGOCfDwdSkjNe5EHvLkwo5yyK1VzMUXonBFp
uTUwYWiIIGvo2HiEIt0PBxdUXm3a+AGuXaqfKXTQ0BtZYmsBxa5mpbfsgM94FTqZ
iV81QPgDjXz5X+bMISjWYGvM9QKRwf7dmOIULE1zRP0kQyvhA2ArVTQ/Pwylw8ur
uEhQKTNOna09QRMM4kCSGMSnXO11n5dlHYVcQoPyw22z3+ndrL5MpBbQDmd/t79A
OrEBLyUxDj/uiM74S0745LKu827NMJpiXLwiC4jrFoSZdYJJS/8o8nPUa7FbMu18
du+buO5qxSFL7Q+bmvltfhcREXbe+zVNi02W45KDG324utcuM+HZGKnF8oN51Xx9
MofNFjXr9xVmuaSdhSTPAF5T3ctKdYoo8Bfsj25lDhLXkXD8+kofdgR+ubG5rcP1
PHIzJkilnZ/0f49DRHogmKZExdNRpqvnT+aKArdMIvwKOD0ODhDBmwWVxo16T7R7
30m2Wk4mzFi/OGv2rbzpm3g0GAiqWDEv4FBgvKEwhPLbwD/XFUZ4LP/ZqJxx9tLf
SYccj7i2QuK59ePqS01yzygu0a6Nt5uElaKr8K3K7th8tBcU4BKyDBflVg5QshqO
AIA6f75kLeCIutL7kcJLO8VcC644QvIR8IM8Dvwt7yqIIFD8aslHwrc1s2nWQ8X5
Rp4GCMO18SpjuI4FPsJAYEBIfuUDg6dSYEoU6h9nOnfDX/+4nMkP8jcx5v3vcN4v
KJkINIvPmJFwe56EHuf0n64rvNJGtOx8SJWqexAa23Clb/AqmOSZ1UGGtl4p2wJs
I0rc4qJlYcllxIoi5cdYZjf2hgk3DXRnRHCAD6DjUuwyHbbsSQEGVMUvxddGRf3n
HhYppGqA+j91bwHVHA0dj7GOPsLEENXxw3trJN0um7iDeHEcMYjiPQqg2so9lXm0
nk/CsgtEG/VUtvZbWdp06YuX0Fd92ullkItTsSQ8BtETtB6EzhbTi0/73tCXdI4w
DVZk+NueB6LbeJA4cMjcB+/wIuutGnVQGDvsrnLSdzxFxQTFd10q6aRAC5XdsKKN
uCLdXP9X6OE/7qmf2KgvGnImWH7Zh/CSmQyvC78xhJxU1Ua2GFr2msi9QiLDdxAD
c+qzk/P/Tk+vIS04XxodG5kTYanFz1rJuGSIlYONaHICQTzziAU2wbOk1lM0owaj
QONJjKvdlK4q7JVLR4nDBQ/FazkidCbayKzwX5QZZjve8ZfSzgFrjrSHthfkTPig
9R/ATfUYv/CtjmVD+cpcwVopFi4qEmFD7eSXGNyE7xibqR4aTwaF1V9QCchwA61C
7nqsL18BGBR6bZQwkAPeSrKVO6CA4719gjUSJ+DJuTnUXgBA4RKErdgl/Jgq3x7X
D25rSg4TOSGWDzOxlqu68JM5f5dsw3yCTwuTU5zJrGnmHLrZzmsNGd8wODC6CddH
v2UPMR3qnTRFP9DZDxNiZU8hV8/Y6caUNmuYnAnmS/llw4stXM2yO8VC04GtduRP
UANXrNA2rKTaYFaEzKjScYlUSrMbnE3Qrw3+zgN/zVeOB57kCimVdpOR4JOdxxad
oqS05IeR7Gf47NAyPfHZ5BiltqdM2jOzDPLxaqzIR+f+jS2G3L+WwgxazEZgArcm
JEK7Mwa2h2m6ltLGve2EpRvZpgcdZRojc3SIePoZShhF5Td1iR3N8G+cpomTls0+
qA31lSN8mRjh471i4iXf+t57hJqVk4dJZV/cZyPu/nF9RlOuzuPvu02ckwYhj+37
wjg1oM4oyYYOz75BXi+MiHVSp3gRrTOrMHvfSKQ12r0wZHHVlJt53PlIs0LdGNEa
cECeC682ifRITny2xxpX8VF91N1imAmNdDcZ0Nb27fjYA8eyA2RqJyvyNFc0vs7R
CM6ZSkP7tt2qxwmQ5WrWq3PGAORkLiOk1ghHa0kZSwrjzsveBV8HQkUEuiMonMNB
FiVWYF65vPBg0v0Q7l9Hp0JkfXfVHD2gKdDgUk/olmPZ240xtoWW1jLQ+ywVTLD2
iId0YDkaoSfD+5YE1ThyNnpfcsCf1y3I9VYhXKRrdoK0/jVZLqQELajD8RKxuJV2
PD3sNahrxWJx8YoEcinXa6ezrtyO5oh0a7vPuWVwH1zysJcrUJRvtUZ6Zw/uE0HO
RZp8AtL9QSqbb06FJaq9Q/6eVOaHjBvtDSK0EDNvEf0YTZEk1bW5+RYFqfzEhSqZ
GwBOhOUkOrgdZOOSncSGJCx/vHT7HaNxceaAHzdJVp3rg4aLpINekF/2LaHw2g5V
B6UcoCszaLqHJY8PP2phU4ucZFItstuDtFSAVRJJgHkIzyn6yxsGS5AoxAr1500S
MtNODv+HTnfXCymfKi+hb6AD1tLv0Qv8f9THPJxo41ldQ5lr5EESvkjbZp3OeY5y
0BPQiT4A31V3bsJdAqmeetYmFtmfA8jrqWSaCf/R/RPa6WjfjLYMvZgfLDXSkuYi
XnSu0GkqulrF6pf0tvV7A78ppR0Ultb0A8kqYt4mn+HUQg+VKxeQsnGylLDkyzME
1+0OWfFIfR6BxoSWNuzYjUvhQwjcZcM6BN8wL/r0oTSYeIxEabRROYrOIEgkzlG1
s0jNdn4tkl0PySNTsl1Pxdr0VcJW4E2zky8Z3sum3gWgH6RYM98pdZgcqxwWers5
m5jLUj/tRwtdHjpC7GnHwfwc/MD2tcnGTS2B3qHWbQ/+FSJuwISIen3Eu/kpxm7X
kqjjcuF8l6nKRvG+3B5EGtWWU20Ikew8RHT+3d6FSisVudd7TB5djyDnTZUhASGa
vQU0gJq8KCvjl84r2GiMu/nfLYj9UzIcG2c5lIMUSVRzMFoPgDXQAdg3ppveXKPY
/TsDPbneZA0jY56xdbz4L2355DEmX0jhwSZ5fv6hkGEta/k5dq6tMghjwfqQCnfK
1T00/OciWIjUHzYhBOq1W6U14KGuJN3l6buPZUfQ7WLlDrxT50KvRbKLXd57W81n
/2dcWRT/GGl0wtLEyf4hNfnTHXWsrXwQ8xlvfdWCeD31wDcCsEuVNFfTXHJOu88v
+XOE3+AgSSDg3OQH6yMTXpsK3A4xdLUV5FhrHf+BMwY+NM9vlvKYNDAFZFix/dqf
wRxI94XWXcPkbhBZQFjktqNcYmHnTgWoWtDctnZuzOVYMQK2WagtbcdmZAFbQjtK
7PRZ6FqSz1gMB61EuqEmIs75+rJ3V+2s9em+UbdDILkrDYvvVPSMPrFGWNtyps7Y
hwxUo6cXmWFWSy/LE9F9TMgOrFV2H4oqqAm6r+Znef31yUqTI1YQcGn0PnOTm2u2
1FN9FsUCxuhhk0K50mBos397jQI7uQsnNXA4RaACqKtqcGVZyprSlShkjYM3QLbH
aXKcXZiVq6mVf+2O2qJ0nOTl/jXWXII/Av9jTziNTMDYIBu9yYaKHGaQIBvORL01
7Z6YPoAlu2kmiZb32eC4hZJdR6KBM+LhPCOQJ/nd1Btp990Gnb9RaTN/vKzOf1ME
1m8E1dorCB2s5eXm8FZWS3RH0rWiHT0juyIlSDNSXDtwP3gc15oPUHWgv7I8Vm0r
DFMyBoJ3XtLFXNkZFrnefmZR59Q6i5JZ3nplDn4PpiaZv+EmEtpS3AdN7Fr3fKVo
/mO8Hz9zSKszAPrhh6ARXAcRieJP3u5QeP6fTg1NmEleg0TmmzvbeZLvY4L8yVBl
mDxy9fULAb0L1bdY/l8Jnfjq6sOwtyWro9WMmr64oLJFK8bRJFir4vw2F9f0dkwX
Gv5dLSLB87/FE7BrMcLu5c2A4utk7a2wHTIOQDQAHohVcNbqtklUfEwjSnhGOP7D
TdhKKz6GJkwFVofgV/ElWVIYfTc3FocVm6KkhZCumnFpheiM+WE4bgDKpwjfNJwF
aelx2Wqn1vTp7/fvkHzH30H0aVLQ/iepXIiNuXZFFpEVeB2i2JE2fQxHjDIkSofJ
EfkDPRHWBaQj6263PSGg4MwAY4nBit4frZrlxkHjaycNCre+fi9UpPP+Im6zIWPx
6yHs6DziIiVvAdPfWmsQ8xVuj2YZ5iyeNuQ8I6UODvs8s+fq6GeKM0yVzcpnJFxV
MXKrxuTaSx+xS7MlzoJqKs7Rt7v9NBwo4dlESespGFXi4k0ecBieCTChD4u3LQEt
Ksb82GYEzKGSLPDhZKeacI9BPDS2WBTIJqZH+nPYBje5xdcIgltcb1wLUUozegJq
uvvaDPb+2yQHrROvGF03qObRfpYKvLH0kiYUWixjII/5T1b+OYNwzSiMh7HOrYcu
vxaL2xxDAjjQdumRNXkHADsOK5TQWVBbzVLatN0uXKl02Pjakk3zqNrhoic4yXXn
zIxkWWNUD/Sqdahif6pGf+m41/o2X2C9bydHpz+Q9/HIwYGewzuc7NQYQCiaOi/G
hnV9WZR7M8MNDjodv+mt0bMhK1L/z+sSOAFaY0CUg9zxR2JydqmA3KwRA5bCDrd2
o142Zd6Wd6U4CI+71Y++eqb6tdOdphFvb5owJ4V9xU7yroUpK2tf2cPnNBNftjCL
J1vngqWX33GmmL1txvhosl87V6RE61jLkenvOGbfRJGiAvqDBQrllh2ax8Y+b8Ke
MZqcQcFeUPO2BBX57UOhEyUrAx1emZeCvhjtVVUkwpiOIyl/XcskBCT5cJikpbgR
U/SEewl82Oeb4mE0DX+NapKD5ji1rM8hkXP1zaTEvbkOUppqW6XH0EGQsonGXDKy
olP+jdETFmSPfTwae1FD/7eh+oisSc7nWcoG2WXTkgvn5JytbirFnHTX5bxy2h4p
LC7oHt/2gKd3/DY/X4DIiMI7HhIsZkyx7sgzaEWc7oNUXgs9ibknYpxlogYmN9XC
taMWSKEgdO9RzUQMgBIE0CQS7tSeCFF7erBsqrPw0PAYeg5TaxAdtgc6DUxaqsgN
JAawYhlBj6lMMqC8QLlWugMbPpc/MvLV4HACDOFosD+wmpuXLVg776W3elu/0bs4
b2O7oF9/QpW1GMOfmvrqB/OiynA6Y/jWP15D02wuDlt1QapDhjne6kwQY5Qibdlw
WVN9zs9+ut7MoXAnF4Zpr0u1r+/LivDkwgij6e6kGqitwx3B7uVTfPURnO30L2do
RfmqdsiaTPeYZqsotxUrx+hbse5ZBZ3NRyez3rqqXgxqrHV3F0INI4F5JKh6vw9b
0api/4I82TeBZ9IYpi7uzYRnbKJ/o2OCoGCaGF0uDWg8VO85auZQx9kUWdQyW5+R
RKMQPrXLoLv1RL0+p6VDlt3ffmaNazcNtQV0N0NJUDyUzKwZfWKNQdVg4csUjTqA
blePLNRx2u0IIpop4M0NtQpPheUIKu7YqI5brGjvvjSleH9a+XvJbR/SWcsLUA3N
V3S/AJHlP7Lw9niJRZMRVQNln+oCuzizVKdQHHWU3kfuSDRwFWbcg0TsFXEwz1H+
VCrol3upYUAp3ecy75yHlUYpzOhGZxarfVo+rKF4TE67R/UGsqXp2OZ7cMExUqKs
xS30QWQZlZZYYzUbETHLAAL33J02g7a1KBilvQt+jtoHoRJmtrd3M8sLFsZ6aQxv
sOZHVP43NAB+pCzdrqx6EObZEyicxFPlBfXXhYlY2Zrd44bQ712T28aEEY6hBxaZ
NTrkbpDPEtvGdMxRRBMHAvIjPdBXnirZ4Nwfk7Pb8TDZpP1x9Czw6QYwrcC+lGD/
RA+/cvqCmU6bXvcl4EIoMjD5mH0Zdj1+0YnP2yzmkEwoqFy/qWvsNvVjHmuc8nQD
bXmua2G0dos4IteEbz1o3AmHRVQ/DIw0HkQi/FlFgtOyiOXZtDftsCtm9lqspgPw
dVn3ck/K5ZAG9NqXZUS1LEzXciuHCzyEgBkgzk0/YetS0V6/rRdiuMKxgh4LJCfX
ihSPand9MMXqCpHw1c6TxrDNgHI8SqWx+cWEGW8IjWrbuxSSoDakjEE14v29ZNAb
z62z0BnPGren29GKpWQsPOixdn3C9R/P8BPKTIcomtk8qpZHrWXPwXx3zr8esIKq
qaVKWYDkjHSDUwrGwbMl0iO3V+tCurQIULqLsCV+GR6so0tjuk54EkDE9C2m5a60
GSmZvTD5OHKq/WCtB83EAgO5Idnz5ZbW3qBMmWlqAKqVmu9JVJ9PsVZ4+9PvTOAG
f+XulZmym6oAdF39hBFBlrCxLnohfxu1gYCplHg/yjJtIjnetLT/hzmWDGFoBccZ
EUTMRZ2bTlE48Hx7vnTuTAJIcb/G/UN1Xy2oXV8rftydCCnQVvaiYBimjE4PFlq6
SnWZQ0hJ/x37fUtcWSuH9fSRIQ/X6e1QZfl7JvJy1x32PYZSry4l74EeYX+iMvkv
UF+mb3LAUbSUCQ9pI/Yr7fbugQ5P4QLAxgiTxA5/u6SKM/WF1zcfLDERV3EhBvrS
UeqU3nBNkOXh0jZvGgCYKJ3IaStgXFm51cUSCaa+AveiOYeKAa7dpTyHgBilcvHx
ld1in8Jp7hxtRRQLPOq373/IeEJfZ/5MuTxnYaYQJVwcGVqVMQu+wvgaF2D36/sA
41yhaz+ELQVAXAK8YhfoCMODKFQFSizfZqMbmuEyVQaq9Dbt8zx/Foq2vi/z9xdX
524PvTRXJWyb2sOGoGjW5Wm5WpbGqHxSSEei0vLBoHa5UVQwSBw+W2MsRVziaM/u
Xz40GZnbWqDoqJIICEbUtTyPuQQmK3cq6Z2zEOowbrypPiloE5xv6hdnMOgf9774
hz/37ow0seGui41Yj9KuXAXpkel2yuutDmjNHuf0nyw3A/7grya1AG9iCTadFfez
1LBkExPHlP/PJv8h6lmltbvgq1ltGyn/7zMDay9JSn4RUcD7BKjXhEVQmMtTOpU7
PlwzwjRAATIVBsn8xui3mPbJXQH3F+P8ccbxAUjcPglLIwl8Z0VCQe5UCrScs6vz
LifeBn+btMPH/7+sUfknH8H15l2P7iZOEG7XWI5zaqcpzF18rF/ZHZBy07nPQ9fQ
DKJfk1Qjl6uNcFnO/BGCzGrAcG0moc3fdDfkMP54CvU6GD7qFiZV8wybm3A7bzyE
pugr/f+9gDs7hJPyvyXxe9hsQ7mcBKZRryh0xSq/DttHjMAYi0Lao3L2SpqsD8Lw
IOw0pdnG+GsZel599w8xbo2ih+qo3ryeB+QBLpWZTTWWSTwznPgs206JAvSFro2H
NKpR7KJDFWWmVsIvh3XSZhP38a2jyt6x6NDvwS16nFOYrdg5ixbSjR6ePC/vF5Bx
W8YSiihmUEfJuegqJgyp/iwgJju2/Le7yH2PizkfC1Cry0hUrbfFLJ88rXK98xMG
6fBeuhPsn9+aylFuwwbelmCKpQl0wwBrobPJZAKu+spljk7tH//xE2GpJCxX7m8d
0try3PoYePlr30hGo8imVuCcnX9KaPE2MW4awsDwG7HwUu0xHOzNA8c9TfNV6TEK
px16XUuJljn1Xe0xV24TnNLiU9oK5XsIsyQEChvaFyf7qLonf4a1WOI+1YnUR/B3
hpHP07RV5hvl4OEHFyPlL3NDNCrm7iPnjIwUGMNfM1xJXaugZpIsfMxA9SLjB8Ht
00v4skN8RoLqx3M65dmq4JKgiGMahIXzI97kEX67qxGoavWlxlB9YWlO2LgMtfz1
3UN/vDX87MtSQFxkIPCzI5GtjRwFIY34lVdZd2SbgAS+ctT0mj/xunTDmMWv+ojm
qo5hih6MduGKLEr9GPoD5qlsPkdomWuiKn9/ZYdIeCIshtN8LqWbrUSTobbRF6Fc
t0qDdgl1euo09PoSu6xLPZhGrrcY1Z6ZHozRggQ1/5jTRU3iZfsV5J4VFA7eHFNh
AQKDwI8QVi0NHiV6+OXQtO6c610vuYdL821DSPzvEhels/6ytS+nR+/2tajB2pTv
uoBptmsDvmq4/YFaw+7MdyE8Mva3j3Yd9ZG4eLRmXkr0HxJtucAICQgsCiUES8je
qYNj4QLNVnSmdVCofltzlxUIiXhgkS9c/lKzHgp0sveu2cyx+Y2ZjJiz4mneL6UB
VgPfB4ojnIkHpyYQbkET6DF7n7q9sQAtZmIhomz/ApHAulGODyP3wXxg9t76qgUu
MQ1rRi5wkLt6ltaEsMEcosPyjFTjw42pGus/5xCGwIvxBIWLaoHM9xROyjotBmJ6
yhZIwEDgsmyg+GzteEe5E0o/IDDUSew9U4FxRxbJ+g/yjeiC+PSdRdqmuaMFb2aN
aVjH5D9/nDqIozWh/2opWgJ+VzmkS1nto0XvgOjnXYlR7ooX+CUlWNdqDtWAzFHT
q7UUuehprN8TsBY8OZRKAJtAo6HL4ZxQpfztzW8dgNKXhCJ2ug6TyMx3vLdzRF39
7Tm0kZgWPi48ampq9Ir6Le5y51xuVpPUB/83dnsF79TC9ByE4lJ0TL34kZSijbh5
zdJDP8mWeHyDJtwsi6qUi0xfQ6APn4wTZcurBaOwoKr/86CJOhnDfdqtQZIQQ3Dl
FoGmSyPufxAaR8IBWvGItIkc3N7tryup5ImmHrBsGCDAVp9hTx3SLnmbRUTqnx0J
fHp/PjPm5ydNyOgF4hvdVvc+dqZ4SE+0/22//I+swmCN5BEkHAVx3sfBr3jOB8nF
c3nYVfhijzT5TTKrz2Obf2TxTiX98X986nPJOfvayZjYFvc/qJ0Jq03gbUQDttxR
BSX91xCfSr/Xt5qKjlVuk1xSJqggeGedAIT5U/z7dA0E+1mzSogk1l07GKzGBgNu
Ee2bx4VFil+Cr46MK7tY5ywpaUGudcXPlx+N7rvQpafhPC6Fgx14vTV0RBaOF8gk
qQVoWgQiWEgrZ68zQ86iYO0oMzM586ZTXW0MoOSj8FZGVgwSi8tyTpRY7aiZMBgY
F19s/5/4/5pV6R89CcDsHgFRrzQpbEhVC/NWWvXFvoS5MKUa/Iq0lRX1wa6N4Cs3
eX17bV4p/AdzRave9rPJeT+0Bdy1EGu94ezGKk/MCdmuOmYs4UauxhajXlx8wdm9
S+vNicTfBjVU1MEkrT6VRXl04nmqVXEJp2N4tdPk4lXVvM09phEihtxsel9Xszx7
ICLKzwZEUedjRLyNfjPtAhhsz2pBfOuYwB0wexBI+3Gk4v1TGxnnF7C+MySgs5Re
39eerRKIXfI6q7Hg86DEpQcs7Q17noT2XnOCyQZko/dGUZtuarOeTTpleH7I7g8A
C4ry0cZW+N8/tOA7iO8DqkOydhTRt9zOZJUScmDDbtwcYq5dNwAHTxUMHGl9iki3
Yl1r3EAwBU8lLDkSrem2ELSv8ObgT+XzuKMd3Qu8Oma0iFBj2ngvTVE4lq7pm40V
y6UHVGM828QKIGjdwlvxIUmyRbyQT24LV5jwHpUtnkaVE2ZmZ6LY3PMNIwL+tMcE
nvUopL9CBqJQHMPmB+2ZEDEA7uq829pUp3r1sD0asJvcoc2MtKmYfQAsmwjSM2Sb
0DgPya1oX3drCbmMjmnoG//0sMoJVlTAz9rj7+tuDwOTjB5xqOe2MPJ4MeICAjy8
245UGP/5TARfuJ2O69LBJZKIUoWojFw+kMGvwBMmHCHdPgpeH1WLTs+DMnm2jOb8
ztcAeYTzGNOiiIdHVyZj43gfgYgiC4Gtd6JM4/cYKKmPlIRlFUMu5JqtIZWvYgnZ
I5AaarTEXVSGIEKHEh37W2htqq/mAgG3rOdVk2hEp/kpjuphIjcY7JofvGXSxmuS
UFOEcrZcEkWzwgHLj1ThpsiR2VPtIoxSqGfojV1MDALr5Y16asLSPSNzse7ytIC4
3JeZ/OenOSX0657tzCwroSCdF6WsbbaQeU9LdCnDiyHK01irmYzHC1M6PrCY3p+G
xEewz+evBSRjZILqh9v7jgZIAn9Be7S4SSKJcyV+fxJQVLrOJ4CgwXtuYYUGoB1L
A2hO+wu6FYDS4u3nsw7pWsIzPiBjJKJoUpb+aQUe5mrtb6wwi8oJPtvId+OLAKJM
wvz8xOUuQitQwVoKSXDnNkLYz6CiSV7Ji+/wNG0NDFTK7gVtp7EimbPfUqxZoWt6
3KffRpJYGvUf9WfyBl7cWS4CgWV4Xt6Nc+e1jC+KYc8fbeQ8vTIbfexzEg9Lq7b+
ctEHmH6YCISL/PgaKmVDYnOiZh4FqzACS2KlRGyRud0aBP9cH20tXuRMqF/6glxO
D+HVzyiQS4htcitXojAkGWM/g0UQQxFE11xuRyzBYY16kxLLOVCBwcIp7PbFa//5
TNvMDqT/vzd4kIbTQ8WIr+0PL9Rpr0+2rzhcg08dcZOY59Ryfa7hgjpFJj7Qwh6G
nYMYBXadDwtrcojOwuID3x/85xDYe0U34UgqjkwR0LyeO3qRe7Vv0sxdjVNqgRXu
7rWyYOx7Y6CYmpdG++CE+P/Emk9XYlPqqlxv0s7aa1rX4YpGpuIDWlm943QGUwta
WN1yUJ2bhvzAN/GZ/Q/VDfyIYCdn75FCIE0UO6C/P/+QhJn75fFJL6bSp/MOwKRd
YWMtqDHfARDkYLbIRUPg/KXfg84lhb3El1t7+PDYV35tEwNR9LSKbH5F+HDvdCmg
rBEcPClLG+jS31lpE3x4GgoEANdiqigMPNrz+TzZ7cFYg2zFX5sjuujIcO1V5vI2
Nbp/pSBxd+KVGGSrFAQoVPjAZ435Dr+79+C5eAKZ2sb6/+mrptBmz5qjrOr7g6y4
iGA8tzK5eRCxFWC77fWDQ5XDVDSNQH2KCtwPcYA6gq6348vKW3MwSpFn3CarwUGq
3Y75Fn2iMO0TyZE4czsocyH17kr7qfNPmh0Z1doqvzTRHG1j/4Ou55/XggwQ+2VE
ysP/6Ao4Vpu6bw8HtQMKEesz2T9r6q24qy97g5FXtQOChEpSu4w8EqimYlIr/441
1RYAGLi7w7ts0qGDUS/+IcCyjD48IlwAG2IqYihQQompeylUZxt1DdUc3boINKsf
ImZiSVAS8Bb5GWVDm38cBQ0BKwTKveEfcWMrZSKhd9Uq3pdeEzVeOGCPjpZ+lHyM
OPcDEFH3ar05getnyxMt+jLVrpqJ2wULYEp6JR0hUnabmv7tIfDTaRb+oN8M+zZd
m1GSaWcTslwdDkKj7ywxyNgZNpgCAwMe4tF9JWSYJyF2hA1KCMci3WVxsXEnS82I
7qRdZDGB0XWmRIOv9kcBWk2UHnqhYWbezehDDryu+jiLTlMWsJWXO1w+gQiFpYJb
C5MT2ywCxpLdenVenHqvYbXEKjNEpHQ9F9ZbhmDuy08dnbCLIKArotn0atDR6lMU
Ih/Oy4fJMRLPc5tE8DwQeGwJ3Qe6qz62VmU8Dk8yFy9trS4EbHKJhDbC5rbegbFH
RJyQIWkP5ej+PJHi0TauoXGJMfYBPh1N4uLcoqiMQj5tbXbuk/xN9uazdun2M+mx
N/lvYSrIfIEP36dRkclM6CIX8aM8IqE0mUR7jmQZ2pHNiBE2Jg/rYyAvDYFvIE38
xbFhL3t37BbqtgLCj8R1ocRQ+w1dr4i1IRbqo3C6DgUcVFfAd2NIIZWsMlTnWA1s
mFcREfbEM9jbvWfGvE3FojxD033CfeWV1hbW7WymC9K82nWhf6hFIsM5GXHHgmbr
DZ66UKFApOejxeLN5NCgWYIwv0082RefTntcCJTUIIqiWvITzg02My4WuQjUsqz+
nI0FgzHLmBYFcv3pA6fIx93AjBvKmouAJzppgBAW1uTV8dzfDRrqWaFm+rv/6WN0
oVcog9H8zbxEGo4ia9LkkR8ibHLlwn/fVTS7JqwtDJqB9xs6hQxEqCb3f9DP2JAD
IvniguAZRULYzJHoJFCmOv0kyKpJpEV6KuVbppgyAsblu8CWeKWLFgQcltBRoQb2
axLEUrUREtAvg75CArM0RcP2hssgRV2qxTjomvOrtvvXL+vGGc/hcbQFi84JaHkb
msBYkLB3V+14zSyGpCRT1MDajhIhFzsZ2E1V2efs+MT1R+9w5wD1n3mjn1v4sxaL
dRSEngdApduuzPGVBJ0gbWKyrlbgUVRVXvUdljXFL3MBmAffuyOOmtHSO34Qlnoj
lyb5Gz4k5u6yff2SsAlF7+t6XgRHZLsYv8LM6iq+dUSsUC6kjdoXADyPKaGMEa0d
kpeDpywnarAYEQcxu5oPMeE1I3LkuWvhDs2usF8WHoBlpNYhxu8cc9W91gdqVo+9
uRvkjOCe3qI9YqQvktRMgWdNTCf9bKm1WpCArsiSYyoJpRKtjPJqQ0xVMdwqf68l
sD5epXnN9wUxCLL7RGUW1cY4FGs6O8X/W+d8JzcZ6d2JZX4f8r83HgQfYQUHj9Ew
nEUhOuvw9a9BJFS9KooCeRI+o00HBnODm0+g0rRV+Euhs/ks2tqZb9C/nBz08wL5
mSpV4dgYBL0xbTRpMOEgMyv6vAwEskHMQa0Os+edBTwDmW0A+m08DLPZPyWkhv6H
YxTvZPe+1yb3OtKFHIOnCJC+jvIEwE0hg91wVOw9v5ENMYVbb4WX7CiPRA4xY59e
Tvk9PzIawLWLfTW5xlyzBsbcif3fGqvSm0rGKWrAC8xL1psOEWXPmvSjKbW6dF5m
EGm5+L1ZlYIEPsi3/HCAFkvVm7NU+dPn0rVGbTjIg1hQbc0RVF1E3EQKOEfqrrec
ksTQ2DznWdG2UdWQLTpWdehnryhX80/R+Qpl1Cg4ggq23N5YzCrEXAn+eYON55b2
u4sTL33XKlq3g7XhauFSDCNOB/BC/5j/A1I+FB874sejc8m8HOHa9ZPWIPMLTaT/
5+3Ncxf68tpvb1A2/FucUl5iXg8da84yMrF6MblBnNYSZXN0Q1+Q3oGOXj16J5sF
4VHhEwHb0kr5/jn680Axk6/ieaRpdht+9ETGXZQXXPElAn3vyNACIm53mkDqABXs
CcUXZCOgiEdPaGRBpkzVddESHWPquFlcKnOs+SW8aOJ1GRU8VU9raHVRvj4HU3Xf
9HbGEFGrw9dwqJ9Ehe7iXcwAh6Gk6QGWDcSHi/bfC2FL5Goq+yLXzQyoCzRqtTzW
RJKYiv7JyouW2IUXqel3cs16XeHusSQyl2FxuXlo80PJbFrTAgisUpXDNeBDMQEB
yZ/UyE9/6y4yQkzckBrNLNenbATMsm7eqU1aw9uRl2jfaimy08zpl77uRzskc4L6
M7lAuhwEATPuOrSbgCNtnl+g1Gm4zZ1TV+zVBaGFEUiU34FyqR4sSlaUv79la9la
TDG3OpsweKBqodrJCKV5K9dZHQ5qZA04hSawrYNjVSGzBQoziWPYh+/SaZmjYuGw
FH+75XVCK5w3t7LKnk2WG3HcpdLop+exZn5f9NJL2tb1iL9IwyeF/G4XqdK7EK36
zzr4t8+Ut+Wx8O0jtipTQrTgQF+KZr0uxTJv93V8NpfBvl9dJzz9pvTbsWId3O3G
M+u3LayRRBqwvKJUfbH0HJuFD59tA3CVJNT4LDvophnjtL82Xo4IGVwX29dXr1gR
GmkmsCE/ICbzZYMsJ/VHgFkOYA4nzI7zyPA56lpmULSpdDErjYJEKoewKgpmiEBf
mzKup1BTQiE5oEIzqpRptS/a7yv7kft7xvsudmVZlfehaVOl0Ea+t6lYdnwZHteV
Gxbi/LYbxtH6v2yguhdL6COyCDBrg5bg0TUAu4BE6T65v4yWd+mO1Pwmk4jE/KsO
T3WybSfZh4HpeWTuqFFccNHetlCO6+sLqnSJ6owwLnBRQccjUFbSfPplJhEaU7jR
Ow/DzZTdjXtSxjmkRc2a80Lte0nhDv/A0+xW6B8rnziBs5UXjDN+zIcBwNJeOVXQ
z5fhi5XN38vPMC1o/+ZTKQdOOAvGicvnOvQi6asus0+JMuPAgHZmbxuREFwz1RWT
AmColuihCjIiMa2vaFfWOo5D4sgJC3Y3yql+vk3vyv4DY2TwSl6vvzAZZ7eAM466
SUsq+U5lvB93M1MKxbhX7shz6Xybv1lvsgoOdYQ/wcUhqjx3TD/3NcC+lLS8BkCT
i8HMsQfKOknXy4omntd3x5SjZevt1I7oBOoZPfyE1tuYigROBrV7vrrNerhvoa4x
sZRiyYNx6tc3r/Ggec4YyzIF69w6UjnHfzGsismX0H+s0Mgwgv5afvgulmjuM22r
cHGrZM8UGMfuGAm8APYIOOmrQOKS31ahwC7VsKVKWqzp30gvIxjYZ20HjXMabnE7
8YjSkSowrBSKffQSG9XNjIiUsjDRwGbYtYFcF+c75wC5tA+h/4bu71X0xtwF/WXB
hT6TuNk6hNb9w0syGcIfRnpYnUJbDojlYdcCmznNA0JpY/WAy7N1MUtn6ZSWeX5j
zfROy3zwQ8EqfEO2n0TpdXL2+kXyzRTQiTae12vl6HX3R9kMQMhllG0YB+NgbWzZ
Abr70wDlcM8snr66lSPQlemDulcbQV8ZEqlbZOUtuwB7UHHn+My5MRED+0rYRYEI
4hDuj8HMM1mVmwCPupJGUvZflDMIiSEBtFneZTxuyXn26+20Y1cAHChSKruV2tKW
9akqOs5PP04s4HEekUxo53DhU2IzjtSCsc4edeSS1gDNEthfzUFwEnjRYvTMlfTN
WGo4tccDg+zhrtFyfyNbQeHo3+ekHOqn1qIBqzNFQ5+C+d267I9PVT+ECSn+ZnUD
3cF6Z3hAGUjNZP1ou+/0RHdyjgSfXuN11gz/1Q+CCObc3/h0Be6c/QIlyf6Y/pb3
xCNsquS2Vdaf7y8VEvbJD7VKsHCdSqlaDg6nX2k86vFmd7n+Fr/zTCdSI+sPyNBd
7PGTeB2QZZsTciOIZIR61GSRqCFZa3Fmw39tNFoelC/748/pl1LMx9/Ae5cKKyOY
Z0wv5W/DwX9ipjVAesKRH8oT+ycxie3udgYGietuRiSaIWaIFS3xFjiV111rsXng
m2J1iWtxfUrYIUfGlubNA9yTwBnycprKVF6QdnwHJLf03El0Jnfd6W95wzYVnYxT
0oGRPqHVZZK8Dxt1o1Eigm+qnNfSW/Rh2SO2ifVDeU7L+UtBbFb3hPpuJInE95Cm
mziC0X7hZQTeJKzN6kAio4bgyAuER8ccM9HicOxAWyB65tzDyuUw5tlPM7okk5ZR
8sIJyE4CONjOv5NQ364SY/8SiTKAjD4XxUrjvgqDWS+3D7+a/iXVgLlAE6JomURs
AacolM7nWxMrqs0MvOPQa1rZZD15eCSIwm+8OWYv987EThngHN6TH2P7hHypGgpz
9Fqf4tG7hEe+udym5UVCg4j3wcEJgC8NWqJxEpds6lJZg5RAx4P5kHR2oqdyH0Rp
hU23FXKTnpwW4bowODQeszzxHC4GtBL+n6178O2FEWvcwgI02oBfJm0zoWKzlee/
RkWydfmTIUO6cPrMsACuTRuqxNkYrKKEArSlS5cSXEEh9wzGBl2xAtA0WV5Xts21
NyEvGh4WwcLEFrGYwKIlBYpWKWsvAhEXlqWxZtXZb+wyzRtMZAf4AUxTz1bPrPnf
YbZZi9oV/TX/rmi1k1icETmgUzTy287e8IVoAq31xcNI7K0UySefE+griDEX+1YQ
gdWAfLyOj2ANgeZe3C1y2+qr++kAMyIKuO01g/90c6JbWS7Xi2ESuwfvjFc3oLHF
B+Aa8y0Lza4i43idCJD4eBRY9P+cXxQr0xFeo2EV+kHFAgpKDILsgfD5PiNYcfda
e9dlqjTIpk0fqkKidiAL4MUT86bYUkNbDFeHIcxBPB+KYZZw88eLZBrAh7etRW/L
eixEjwcmnzcN6MqEWBBTiNKBHyEUj29HO7nVpVkz+9ZDhoFj0yhl4rDxoKzDb0+L
4ZaNHe2cO9LzEFSbSAvexTFTxBEshixgZsqrpd1caySHENGXSB1pyKU1g+yutzFf
BuujUXHgvDoXqUothFQGBTwqyOBeAZfHYgL0Gp8W3o23RKJNEOUsInd9psowfBHK
OxSHJ/Mx/K6Lo8AawA9IdDdBn9ShG8z5aOp5x4b/92Nl2llXGFzHOBYaiS8+vatY
+Dk8vs1e+bITmRMiEXY9yxORbtobSeV5h3oIsNzP1q29b6dPUo4AzvVRMnJlYAXg
Eh9zdKfXmm/0PCC+nutLPpcbIdXpRTcJPzqv9Dgb1lCeyqcVsb43YL5TX2LvXnD6
l3WQh7he4vLWI2b2TSF5pHuv2rdr24Hd60K08mIYcfHjIKsc5nd/TICK0bBYmwEu
ZBL47anbLdtNL1URH6q534epCPzZfLBGhblPWVW2uEpGJxZFJR7D2581bZbM2uGl
QuhcSeVgMzBO5LdtuiMI24SZRG/NJ1m+CdDD4YWTgzNVB1Q/MpSG34BgPFt4qPiL
QVVCnAiG8OlSA0GAT5W5aAcspWt/V1LUTV9/5NLbdBdVP3m7X0TaJYkcM6pQM7wQ
E88AL740UggNXyYj4e3y0gc1OyUCqKZ70oR+IjZQD6hLmXZ+ou7aGE9e9IcmdRcZ
YJ/6aKb6tcOjOjpsZtb/MRQLQ8icLYYYFgL/LAF1uUu6RGgveafSKEw9ydbxttb0
3IHkS+PmHLutz/aj0sk2A4w7M+P78zY41lwFgK5asQp0RlNJV7Wi0dvOusGIl6t1
6AhS6OvO1Xm96rH5RX96ELZk5DF9EZabMbFxjU2cR/MWepLm4w3zjlY8yEJXYyGr
db8txf8mctZxC/wbjAeItGOPg/E5ET8j9fIh/upRoxQS1UsUmP+n600SyL0cuUh6
2HtlOoTC6Syhx4Z/5h3RuDfpzVQa/03oWvvheP172JGrBdnJZgaCXLybSzXlnzMO
odKjzhJ5a8tvJ8SWKBmpqbncVG4WSTCPjrkiIspH/vkIZ/Q0BXI+93S1Ej9DzOIt
+eJ9PDR0s9fJWGlx8YF1766lYJM0mkbuRgcVghYlrit2cCicdU2jOhCiOq7gIRg2
8lgNLC4zd8NCJ1ImCoCOfGjMHX1Sn1HlYn9v9Sjio4/pSn7QE5TSrjDPlzRt0MnJ
WeGxHc/yTOV97bMSaAorpaZzwmPxvOHH7SlGV1uSPhKrMbpWI4joAEHHMVTWB/vi
ipJaWbaRNX4rbERvB0iHGWJDgrhQ0GxaTEXfvLnA75s8Xzm9hHyDQxTMWg4/mnVI
aTbFMdzrqLlgXHeRcT/i+BegT1VLzbxjjY6JOd0kYT7gE6oSKo4G5x/NJ7IQO90e
cmYArCOQLsKmiWodIwdcm4uvBcJTtEXeeA6wo/1gvXkM4cT3kmeLOsmrq6RNMyig
FrMO9PKU7bbwgP1s1QfQSJRVuyIAeeNtOAlim/PCxeCADVlkn7KtKU5zA62vAM7Z
G8nb+zUOuPgcsW5rPLPAE4vPmpvV51fTH9t63pqbDilaMISF62c5T25nLXpUWKA4
YdKck4lPmNK4kMTXaxM04DftXjIAFOCbEOhk1DgO+SobL2GblMYnDMe8/1b8Ihon
/ItXp9AHiqXZGCCUCuxneJ4KD3hVzVpcc2a+Q2lpn9bBwM/dh8docefg77kCOOqk
CnKlAJt2YDHZrizD16E/fKC7qBY5zwj7OtuQYw79V45SnMm6UYQp8sjrW/iigtLd
OauUxCX0RFSTGgXtEqjnhyS1f7lI8ghwUb1FwXxvX7e7mc30+uenp0ihfxM6Cfux
uNKDMXF6eOg/Y2bJWhw14FSw4zInNESjAXrrnpUIa/aTPsaJSs++xcRgDOamtB+O
YNmcqR4VN2Z3YVKOMIGocJyCiodreLO0JM52PD2kjv8naA3U5OR/t/xMyCnDkwTL
waWsX4zp6eHeEWw0rH7bIgye8ETlvRB2NsO186iH/WMAyQy8b1EnQrZ9xIBDGT81
5hxEbpyH4LW2CDWlnjl5ba5M/SYBpNyxxkZ7nfRV/s/rjSyKq5yJrpqrutz5WEQH
AGToyavPDvpdM192+GcmWUd58+ara8IuXMa6BofuU9T6OE3OVhwN+RtCzD57c+Hg
hn6dZfqG00FMlgBsGeODN8pqw/AxDM9METkGRnze1wMy75FKzBz5J72lQcHdehkF
2IdCHCuPfmwYHiHOAdvgJWmzxEOKkxdoM3aI6Rv0/VKulnT/h3tH02w7vL8f39Ru
uazRzueaLKchuCDgU0b0qPlSRapnfhptJKMGpjbuoO+tlYDQBQLWaxeSl70EAiiI
g9hZnN/NhT5YOP+9HVFnkeZnG3hgAa4EqCo8FHg5xf2Wn98aZdGFcvr9l0LlMd0/
51dbRkuopR/p/VIaov55swonvYp8ptbInIOPdMvqRnOjebrOGDzjPXxEMbdP1L2M
P4LkORFDldqES/9UroJI5+EKNtKbJjt16McuqgWyFAKtRIzAmzys2pG4RxxO+xqO
AkZa8mQtgtagpKj+rqtotctpEKFBWEYivMELAso3cSmKqTPf6sxfK6vwlmA44LT5
NAQndXtxn2mdYuFX+2//cjw17r5R5WOc4oNrNA0gEtJszrhushRzKfK/BcOWZHa4
D9J4HC1b5og1rPQHb/c89sse1BrrZg1Ft58miom5kqemZcv+8DM9jV+pcdLp/xMz
Pv9Q58WZ7+w41BZkBplWiCQ71U/r9oy+DFp21O+BZDwTGkTw9iKH6KrqHbSi07r6
is/N2yXzAbzHtY6NvyISFzCtYqgwY9JgJSFvQxRvcTLFwHyCrdRrnSe50uiDg638
KnCYamPz+6OIHjdf6TbDYn4XtJl04nrYum/8bprWh7/2BTdXcqJI0zI/EOYyGEoq
uosdIsZOlDWWs/6NmNAZV7NGjSNJ7e1XMPBgzONm852ZG8S7up3pZ0HmYxiVlzLv
VEQu7x76Z5cr9lgXVV7peo6RwGkFo+XfnlL+gi9oIYSU53KDV6Uf9MrL1xgOO+ww
Z/Vqqxx6V9tTfBaFMWoSGZxEsC8BDXq49t18gvzCpn3Ad+AfGpflk4ZRAruBHMbi
lf6ncwEyEIscIkz+dkUuamBVE4MhrFqfp4Qu5uqRth9ueDPzh2kXUsye8V5kD676
IoaxMmzTR94BkM0x7Y9cSoyYUYENiNLO8u9qNZg9r45BcQT7ThY+u6LhXwQ7tS7z
nmYHq87brVR44Va6KuR9E6hI05N2A0PpSbcJBlzL1dVPlVssFfrPF4OSRl2I7t+f
E5I3hs/3ZJqzZEYD+H15pp8llI3W56CFTnzDku0xKCTWEzhWxuXAAsQYqsPOPy4L
JEHeHYUcYtJDIEqZvCVZYJuNlLHusssjWsP8tyXLv1fN0KnJQ+/OsAxvJn/zsgoK
gFh0rr9Ofx25dUyDFiXss4q4vxlDbJBVZt6omigAq+BfBsdHZQgAClNQLdFHFtCY
edczg2Mx3AT/dHVHrCfqFMDEF2JeO7+qZLzGfcMqSYpvpOAv862eHtTqpsqDt9GC
Je+0XW6FqbXgXjhdMLOu456uA0E1ZRA/vgvf4ia0GkINw3DnAs8DXxyBCWd7kjuW
aZSu/2poNMVt2R35JdWZDZ+uEHxesNnHEllsjYanV4Sin1yfn27fSXqMqD1c4M7Y
vuQnjjXJ5et/oC24iZr+r1WvDEtV1VlhBdpSWin6pTFwePPqU9FEIzpFRsiO2EYs
DX0R9jjsTVvFOdQ0ARiojsZFyxqrDtuMvoDhc75u/hCK9jZFp6aUCTaKS8dPFHIL
0n58/QoOdboFyix+fUjx+UVqBQRLTagjtcbfcN6zuHOu+j0/fvRk9Doh2O36NxUg
pNcWy6lfwuE7pAioG14V/waXb4SjzLG8cpLZctQxy/1A9E/ATN9yy9t/opb880i+
LrX3Jeo92cQgJAwr2C80hgwMi6r4Fv2f69LplcdzQ0nDqfFGGN6rlPJFrfZ8IHBO
3Zy/lWB/NK1sWekmj5wtCT28qvS0krju9vjJKXOb1yPx0x8Nr8qJtjZN0I7H8G/l
njP0rQYyIEnoHNz6t6pcuTujl6qRbNZJPa8Q9iixbJlA0BeDjesHQVmgeTIypwP5
Hum/kNbGsZZR/+lO7uoISYaVwntmNGoN6lryfTTCHat8KBmuzlr5hF7UxO3JPoyr
TtdEbVOidRTtPXrMt3VbTkiVWqzzRaZvvkx4r/CCYWOuZM8Y1VE3aznY+rJVmxUj
kEFrGyqPYUJklQM86MaMpwl6T81IrBT5jLkEEk5utptQC1OF7Oe1PJywpUVdszes
jDUVl/bfzRHIB2ceyNmN3iR3DJF61r8kB+0unwwlpMEVvTkjxWoxlODHunxFmg5t
D3tgXuYRCWN8JwaqyJQ0Y3hABcrWwmdMO+rS9zXu4vRQC3jovdfkL/ldNWiQWXno
u9rGNZI6ZchzP4do6qrtGFRR0l60qKtL2UNp/nsOGZVpJn9Bh+oIz0yY7ndJ11Mn
Az7tOaxQlvN440MRL2UpiV1qBxG+MR3bBZotxSnq3TH4CdAv0t+znpVeQHHH8OW2
USjcY5RrtDhJqhKaNF4r91F+jH9lwKtDGt9tAKwTDDRZBbDCbXgKwW7sdXS1DJgt
HQV1atC47tLTA1ZE3d7yqS9g5mFj/TRw05cZ0L34RoCHSUkbRghFBe8kWHsBlwTc
YX7IxEWwynLzgJqCP/VLXHuH9BeOObHtYXdb6Cns4fsCLj61LuwxqXYWi9XQHl/Z
LDNZUGZMzcgTJpTGLLa3WDNHmJK8S0xW/hpgnwnKCQE5tIerJOWvDOHQPvmoYTlf
tN7YZr9K5NA6vMlcdmY32ju0Ot7mjNkp0CF4w+G/8vq7bQ2XBRgrm1E4WvNiZuM1
o749G6Z7iTma4KWAU+oQzzaU2EfEMQLiyaBw1S6mvVFmPyA/hqWvOq8tmiavsPBn
QLC1YpAPhV4b24jmnZdJYOWa+R9g+vuT3kJ3H08h4Pr4Xy+Fpuv77B1KSvRpvAiZ
xePoSV7UuSYq0eOS6FnMSybhV/LItENo8ryZBureDwOrSSkASfQRMfEP1j6ShHWw
oB1j0OWFFoVobQGb+oK/pKSCfuRU1hX0U7X7vhtc1FHFrPcyomXuk5opqC1+iwSj
yHoPLCO5kMelMEonr1717HCHdYJaVTiDiMDQ4PJIJKCYgkIUmbCcxYunndx52gt2
Tra1NZeZxBwcBOPAdZ+u+CnGLdQvic37NTUXk10u+Z+YWKgaHjsfaTSv4+Yr9Alo
N9cMFETtYhm/ojnh2x7XwUO98a6y550OflRHIc7JM+YoY0ARXK7UT61bms3HFB0B
tNkEwO6pOMv55aa7NQaNVaI3baq/DFjeM642IzuIxflN0zDlxPsyv2gTjBR8Zew3
BEgOP36Nr5oILSXYvHqcHvakM4yP3E7whvCZ/dip31s/3hcPc9Yi75HM1D3r58gl
Aqi2WaxrM6FgkDTcgs1nyzpZqrahl+zQlTAfA9ijiEeY3s/AGV//pmvps9tvo6th
iyE57Ub2EjTuGOhXFCZF2Y55Gej+FU8BFbm7VKoHUaj43t15xiHqyrjuYQYiq2tZ
teO6nX4ECgx0oXXphr1KBJjQ0Oy2Oz+ZjyynsocdNeN3XUciAiL04TaldJe28FMw
6eg0Xk5RBvA3devl0pbX6MKvRenj1ZwOj+G1XqFTVV4G6PdgcycqYRXbd9hgqHPC
D9nvrbVrk/YkW44tlXQqD/IYAxw8ecT82D5+EXakP3pUdMOOvSyZuH5Q1wW2O9TD
aYrdRwjjnRsWHyCB5MwmpWl6L+s9CyXEV3rTyuj8Mcbr1DF88eLyov/YFvIR4Ldj
UtOdULGli+PeUsU5wIChYNK16hNb199Ei432jQbpR3MUdJ9RnWGPxYf2MFI2I1yf
/QhvjP/Jw9+fSQdDfABGY0wTJvu6/TAD2OeMyPWHtG57ZFXALejSckvFqSW5a75P
PNVn54DpGexS0MfnxZ8a0OWNsqTLLGiQBK+od7p8KI8FIPm4dgipp/7uwxTgwa5p
NbkiDWSo126t4CbWo5wpcxstSce8m/LlPgKDKmQetli2tgXk+fyLvBbyclzDseaQ
XBz+yK/qaXzHaMxX1vNUyRCMoxsbD/srl2QWzDGT8H5NVxIBtrEsiEMZmdK+1lAc
/JQOMEfHpTtkLMT0KE0ffQ9ShMr+d6/m5AkXlW33+/m3/Q6i6ICeRKT0AzoOXSGj
PPfptvdrt2YN4g2E1+X7RbgJI2iXhpsrxfOBzb/9211A+gbOshxXdjbBEbdzPHl1
R6/mwTLHSbB0IcH8S9lX9qYvaMD8Rd+xUQIfhsmLOROqS2ClH6rR3En3IOOY3YTj
TtY+5g9tCAxvW+dxwWD4Bmvp6qZnYyPtIOndz5F3lE8YBERd6JHcAJbkMS10kzQq
ICFQIvv5k9yS66iKCHhAhfah4/jumaKOeoMh5M9NkPqi1qobTt3h8BkojEQsSe9a
JIfyE7iioH4p8KAWFsdYIphDVl3kktD53c/3Om4rUCI1TvGae2VGJzGJ+qfbWAYR
IfWw1ob+euQmDTu2a4SJwgCYC+taXesYZR6GCXlbIzPtNBbu9YAyBMSA216yBapl
hAnoYv3Y0Hz6On7KdVzzBDl5S2r7YB96Tukq5bw5I4iD7X/jEBj5mPkovTa9YiKx
6FN1ROLAgmDeQrz7b603GGNm1qCCtxwJQKXqSYWNUEJNPoM2HWWKRQZbtE9Tp3nd
3Z36BwcmimfGhTPDTkZA9RyuXwOQaPs//Ymu7hL2ht/P93odXhc7Z88BsuFv12nO
xH4lozJkkvTGT325w1i4jutOCVGS5CHEh7SFc1lDh1KQvFDqUuS7QknWW/Oq/tmE
AWIQJpXpYm0OC9R6293W5fvooujaUcQmvMYq6pcgNRAZ87R4Z3cRacreUZ3bPaZ3
Hg9zM8MIsbkJmX9XSinqVZVUI7D6bsPJy9S6W6OHrO3rFogaEdgSIPU6D1yQ/+zA
8f/Wr67YPm2z1Xch3CR3Mg63db/YE/+szJs6OgxfAZXgoroH63v5ozIhrm3EoWVC
qKamuqQeCGw/9YlR4QcPOBJeu3h2f8vEgtANQ0TM2FpE0mvJJWmCvt81BSSZ6c5S
d4UuWYuqVnIABNlVUzaSQqul4PEjcdvmiYIIw+Nq/FCCn0Bf9Hgp51OiLFjv7zIp
Y2AfJxzVqCuCei09zds+aNYtEFFrpf/whkswCq7STa+NBO7dgbATELFyJQKVMVEq
QxIBEuO3vQvZJiow6HI3KUMb/6yLSC2jsWX3MwzlSjcNzeg64KTjOiZhKkWkJtKF
nvF5HI3KLuQ9r0HdZlQPsfwewAbOGTN17hEoN7w+/GY8TT+yTePoGQUxB6/Var0t
QmL/oNDvksNubrlLWmZ7Y4J7O1THdDm8vf8gPaO4zltsRq5t5ah2re3LyxvCLGnw
KZ6O/6nJwrVdcysyFXRwRGvNTShiRLwydSRMBGFIy8w9AUrmHAOlc/xTpOXYSi+J
c7I5KkIa+pRmUEjNTVKm3PPCuO0FobryT0fqOgGjEwwK1YvCEPmaiXFXDKmYYATg
R3YN8IOhhHMJBwWW4nkoD1//oxYOVN3neQN5UKv8ej0d0k97zImq9hG88ePA5rja
3tg0GwzPZU78lwnwKTpt3vj4CAEt/tYZUKySzQZrFa99AR6EnNy2lh74Fkpqia3b
Dyhj03pN1ACubROhWz44pE7fW6SAnFj2cHp5jEawd0BaTMtWataeVUMseWmDptZx
R19oC5X3TrwegiefVML5DylNDdM+vstb9jEDAOvGpQrcC4qj9RJKrmejosg0Lz2w
NSNOfqsJxSnzU1eOCE7fIB9uo5B41m7VtM1bRg+nuqRmGOC6vNG9sxi2J3NK2Got
ogIc98ZJCOCyIsCqqUi9ZyOq1Pp97/Mw1jrJqi28ZyXmu+7yZyyvkrrDHE/vAIAk
hcbtuTInLNfupxKnMqg9JYTbacI13YUeZ/SIgIaEo7XFWXSlA8tOIaXzk0bThaXs
uQoQE945NLVZiEmyoFJ1WuIORGAoOa+zTFargqXF1Jzq09USJ9mwudEogn8/Cifb
SSE26T3TcOqlND55LiqkiTBsi7KDu3bauLze/KN8n3hfIHaaaexXy8/XknVO6D8+
8Id02O5D1/X2tGH/61pOVL/2E+Z/ceowFMsRXEjWXaOAsW/hz/+Lr6opYrFGraPk
vhyMYLPvoq3F3jxrb9aCVIkynpAqrdT8Er8covQUVlrXFhIyTnSYuYnCP1JQPZBI
2dnrieBSkOWaBXCFWskFVhvEr97O1E6t6aK+lpu4xdtXRaxK6V4GphxIfYnWINK3
aaJIY3yo1v+dEZzwF2fGiakQ6JCZ27kcO38P8Q4hPFaGGWFXXftj2eqk5hTOAGmu
AIuIztmWLyd3GVdNgbRsykSmRx+5TkFjFmEFLi22LiHC4PLLDXH7oVBl6b0ocRpu
sEWeLJcOOEHqPMxODdKG5DiSAESvyMPYs0+HmI/x5n2jSdtPXpaj7ODV7/Sjlo5X
xYeRO+AM/KrTREqAr6frC5yEN7rzHCWfPBqtSXpJEiIFKkSRLFSHfxjZVWVyjXAC
/V/UIWPGBZHx19cNXoJ97oylzkQukRZZEDkL4FGKdcm8WRYXyTdm5644dB9jpb90
T/bk0SPlu5RKoi2wjRsZxLPXUDjamK7TTT/6u8RkoGw94Rsr8bMktnK0ZJYWRRKe
tyyebsXqERqZk6XwcP9c7GMK2zzoPUBoS7No8zsXeqttqP5XZlzA6oXP0VIMNLB5
cX+vnqbxKpqX6XtMtgDK0SnsGXKZ1139yL4bsi79ccOvaafwebHLdBktiOqnZCtv
YNFZHAMs5E9hfMrkctuaecW5cjEFKb2SWlSoaCCDq/xe/SN+CzWAF2TMucxmZGQY
55HZ3OaXj+YAQc3whJt5unVW1X1CJXkDvffv/7SVDtFxDXFDwcFPjmFFbcnkT8eH
xCQ28gYhPjYv7n6tjtY1XEJ65CD7uXVAYHV/AxuyQCtrmpiRX2FLbn8/S9E5ot8W
x11ZIuwm2MRiKe7qEpk/CX74fiEZWDE1lXoupfOc2d1COj1rZLUxx0VWtwVx4zAG
EJgCAXUnnbLthiB5476JrOVmZsp1y0yrjp0VVX5GJllv9L14mjEMUDXBXOhLxOad
i/29Pg67ZB0zqFcDMBB7MRJyf6f0Lrrqiw4JHrrIV+LZUmprtZJ1l+FzbD+03GsT
Hkmh+EFc0g0a4vGwnUO1yVO21TrS6JMnnVO2WEYorQSyJ+9tT8O8B6BvSccBhHsj
XHcql/wexn73hwoULu3DHMaamqpyoSoOdeax/Q+997pqQqI/IxTzVPU6Rlq7oeov
NMF4HOrBONHntu38Qly+mZMZBw2+uchxZhLBC6fVH+/EcYPJ60txPkVeiV6DpdA0
7YuZEsE5xopD9cn2Y2ojVsU3deuyewvOrfZ61Vc+TjHLRkLZVg/VVdsunqxYDrFd
PBGHuFXIrug0MHFSs8ulhXr7lCviL5kMrg5cNSZu81EF4Ht/jXDkpSxgn7TcJ8n3
TOPLydmNqxam3464v76TB11QQPLYYHJQkgDpHu1v1Y8gVN5ifDHeSseosf4Akcrb
PQGkDD0exUlmJvmNr/8nfykBZTvdlBQ3z6NsyNysKYVgRhJgVP1rrQZ5ngT5QcRY
d++WNrV+IRh6Ko3DKxQfpHsXv+BzzoJOkEN7k1RE0DWT7V+2WJw+WPd+fdYpcJ0Z
P4o5kLORwh8ihtMuH0/gRuQldAEaPWBBqMNK3TUz/BF73o+0uoYxaSp8hx5WeD7e
xOCfLB+72BR/Crvis62h59Ua+uqnziUf4dgObNPcOUGra8FD99s7mx+knGV0K4Cr
FYoV4jzpfwk9utvyFtNylmwXbF6xdWaJfQ+wW9cpLscexINBji1Qum4APxK4BLzG
6+BN032O+L1MVMHR3tdH+FlJEaLDy5B5ybQmPdO+4iH2CElR5Lwl7H1w/pKvq27p
9g9iAq73h9GXd9OhSV4h6QkExViPNR9YinEeebqbqdMN9aT4OY5Z6aPAtM3dDOk8
rIT0SwPb0rgrtLG30dfm9tgxw/xV12R0iLRpmEg+PTs7Mj0D+7/OVjcMqUpUnuzx
EF2zt1fmTOw+n0KfN7m0EpkPYXAdq3Vf7uBL0PgV+/7AwkzuS2Qb6ATEWIvGPIL3
OyNMRBxD6UgE2sF3FE7Wi4iKrJnaO+EPF5g2CDRICejqN9B/bEo90uw96iV/LjBx
y4Rc3vvnYtt6qBXa+9lSTe53czLbDNll2AwvF9B36CtPM+tzGrTkDlYTAHur4Umr
QmY3WuJMVbT2p6SZLIF6/m4eqDWTz50mms1/i0ZR9AWcgids1GST4BFbhEOqKAi3
ybTtswlS4O5mIAh2s+s9HCwSmljdToVFAS8LRNSoOcuoRmA5qexvvQZ+a9oPx8Gk
JpzDI1NY7z0nT3icdbQihVwd1KWYs7Chc3659UZJZsyTt+oZgzVqBjp4p1CkLaKE
bLiexB0QR/pq0AbI4b9yeNGcbZ/hHvtjKPMlbCMh+TSNkSW7boeByw55NAuztyYm
ea31NNAiQsCzd0yHCAQJC+/k2Doyqb6unMkUjjF5VP7KDx6kjAHfW/NjtzhgOBKx
eaS9ZUYeV7wFsRdfLTT+T7KjNDSbH1n4761exVqstfYzNAVRhRC2fWed5UxznxxQ
ZoY2Z3jU2B7WlmddhrnRKPbIskIER47m5HbLszWp5Vt9viCxK2JoMk6VZZlozY5D
byvVbEXyRk79VBBAEWBNsgqYN7xtoqbHw6e4gnXvscT6yGJ2Jz6ESa8pC6PtRj++
0myYnS9c+pPkdSldvhrz+5AuWucWfviBUp89otcXbCS2+KZ0+zC5gYaP70GiBXR8
PXv8LcKPGT66VsgEouPF//oFpG5DJoWODQnVhN/CPRov8NMgzlY/84xDAeksH7lg
muAettsVF4ToYLFCuVO3EDWrszO4F/BvOFFGN/ubDG+9rvxyT/tKjN6B6abr37Uh
ei08djUA0wGiTtWc8qyaDnDBeBxp1L5m4ViuvlLFwHw2J8swmv+xLg5kQO9n62Ol
3/bjeys7mjxjToUdE4IZopcyp3BksDkSCZTG2GcaZbGLudzd31X1yTo+wQuGm4sb
JZ3Bh965SmDMuHb5sSmZl1EnJmJeIPLY7mFLDFaGLzWEoaB0MoMQMKpBaffnzzgS
RUWiM8UVupuHWw0gfXrADE3S7uytAX+7XTahIeLsi6mtHuY5z+bwDLmtAJANKYbA
5pvmHr3QdBzZFmm5N32OpqvYHj6m2xB8sEWAbl75UjL+nXj0+jsDWEv24/hxWBgN
tqHl88JFO4e8lUF3C2HXaEMnhW/bqyijPG21Rgj3GohNGteA7FDtrI9G7uv3rXTc
d5ve8EP5zgV8gFXS6wI1VPJWKWyjrF9vbAoM/tNmnko2Avs008jwlr2QJqoYmeV2
wJeeonEFpMKNw+6WvGaPVtEiRD9C9gFLcoVIyiHwJ+XN8w8JE6RafTW5LxHNsTey
zpKyznI6enoRXJkh15Us3matrm610qzAr22vOeS8Q9CzHGwWHhpS/D1bYMnyMJJc
k1t6c7jqkyCiWMKnL96C42a2Gb4LFh6l7I2Mb8hwFR2gIPXWohokIVQraXRhCOyp
QtavfIM3vCgOO7eTMzpBTQ2T6BRVrOLwf6i1VcgUIU0PGyde5WXCutzJh8EBARPJ
pTj779HdIsSsPXTwy7o15cDztYm0rnOm7W+in0A/+YbDxODiZx/UGa0TBow8P94b
xDaPaA0nLpIrnCwIijA3NzQtVu0D8uG0DP7sutjttXzdD/Op2VKWEt3FDaOYv3wv
nFBxTQ1A5HW+ENFqMWl7H1JWnX8677X00NNszhDqKWiiLAtzX7OlKghhj5y0/Umc
Secw8oVUGWyzkwtnc3Pq8SJdAod4RCylM5gDyAJFDIB3y4ngu77edRn9rDQXdL0Y
vviP0k8Aeq78iLc3TW1DoaHuICa0wrmFonWzRz0UUJPZ0O97FLPdMBv1yJoxlqQJ
82LeA+ERR/G9miVVwBRjmAQYvX7MlcUIKW/H+9suX4sF72NzR7Ela5l07vw52LiE
OXoBbb0qAM4ZJyxE+1YqyyWAVcvWYxTLHVq10hw/knGqUAmoA6/0eVgWCxFGECjz
+VxsuY+4A/1uba1OAWN6U7+ca9BzD5Ab0HRqGZ2RKSKzNER7DVEROLwvnd1gyGNA
pkYHvLZbDSxX8DQd4p8Yen7NKvvzSddQqzCNm1gjDE3n+dIFRanaQZ4OwzbMzmxn
uqbsZBXNN4lzIRzr3VJwIfcEM7zuGa3PVGVxt4F6dI5PDW/Kt4ObOS61L73eBxec
iiVndPk5jRgZvssIbm7eyyHavCuKmead5hwTKuklVBSRI4MBKeYb8GSIBZ4PeE4a
iSqRJG+EE6wgH6I8zOdnL19q5TZ15LCoL40oB/p/9/KeoZK0FP45s21NPqIhDcEA
jqw+xrpo8gXOI5ixXEQheQq+QhhN/YSXYhOd6MyIKzTi+EvBf6A1HAJf5aNCYUEX
WgslhdvQHq3Q/VqvoPjFqsrgE0y+vNRQVgqr4sfG9b6K4iGtbXx2N+YMH9lek5O5
tWYBa7UHUaJ5ttf2yweZTttmeX4gK2XX6K9qVVV555gfrzat8HVkUoPxrPgg2JmX
duqg69PTOIzQzix9Te/5iKjVP/Cp29UbQBr+UJRZokOhzB0faIezjYPLWZOcrlLP
3hpJH5BQ+MAqxiqKHIyfxHNgizmamgmUvjZTFd6gJA7KRcDm7b/ypSmeEOhcOGZk
nvV9bBT0ldLgzhjZUlSG65DKHP9UVLmUUkQwrj5qMBIFVXCOuqKsXkcEhbnnbR+Y
A5nzIr9Z+e+jkN0icd+nJ6UhyE0gFbjRpCvMwRsyWfgRbkZ4P4+6Qt5cCLuaaK6G
lkCidtfgPAWu+FYcwG+tJ4mZuXQOfOCG79PKiO74EWkz0Z6Ayq5NCrGOUG6+Of6Y
kK2G36pqhksl2OoBB14CcAvZXCDfiGbIlJy4DxL/937KkJL4zG5Cl+GSUGF8KfHt
MNGGfrUwiMcc11L3Z11VygSsblfOwI/NLqHbjW3Ss83Rz5CrHIPoFUb7wr3GNRxi
+08yz6uzYn4D9YoIFngq5LlWZGFyDcO8sZ9xgwGozXsJFF8SOH5hssl5tNdodrCo
aK9FE+NnoVNilFEEGksrM08hxIO6FPZqTDBBCWI5nSBG5+wF49GF5W4ZGD3L0BWf
iEG87bYBsy3ru5/P9IIGrgpuZ3DqooTca6I38lB4P38cS6coyGrwkmm1dJig2GMl
MgTcyDq0XKz/31x7PfWkVgQxLuPVFs3m9SQ0Z6K5L52jPtlAx1yNOCGGy29WdLXj
9sImOUq5CvDqW6hj00GPgcb5mDsZ6n+mKitk9E1M8bmVHyTyprpXUBDSO60g5fdj
w6nqSFcEXti0vJxYrMWdpfu2bT14R6c4Na8WzzNYw88WZOx1HystDco6cbP0IuvE
7YROxQkuYjpI/LJKmmW1Eq2+zQsCbL/g30TtPILREXYvxWeE19ixgq9J52RMgvxi
nCdLWh4JSLnYdgTnLcZ8xRRv5aAv3di06o9Yc7DTz0+qvXAcv41I0grBLL3w12or
TrYnSATBcMkwb0RbDAtdlZhXKR6d3UgnpkOgbOtHx8mno9AUUjG7/fOndOFmrbfV
K6I3Qd3UmLhQCxlrIyc1DWuXjSvAwlZYdgaj8c3RJaw3Jf+6N0eMtOjnof97UUV2
VdlvG2nhM5S0KM+zXGKirT2zWQlxZCxOLMS6SozvD9lhPaGs7solFgD84g/aPu2C
uFtRjgM+omJWAzL43Tx8CRmNHBXXUT4xyCk3rNPS0NkcqDGOTU4leJE61tmFaXhu
Z3kLvqVBmzbEp9YKs2oU4NiJU9/hOcWAlH3yPR+lfdlXkh8AybQCSYeLvTXKeD6y
//q4At3APl3WBsjie22dhLp7a2FNzJV+cBmPxYmMFZHONCqxs0jNXTlxSr26/y4e
5bQcMZJBIglXOHonR5y6nZQygLtWzH68ucE3PXV1p9dDvzOS+vJZfcTUtzg3eQsK
ufiunaAm88cTOOxE7fNJPRfeHowEHLL/ji8k8n8Tk75ViN7EoAkBXjjGMJ1KOB+v
NmqZfyu7v4KsHdkwKSqwf6DPS5h0vNN7MB6Mid1gwiy9DjuLPG3euJtNnXV1WeCj
YXWYVhD8Em18WiM+f3BayfA3B/jZsHd/EhC8aLSxZjqN1jS9kSBnYm5QJEf9rpBo
44BACKWBqZlKmglsBangYIPubWwcPJXUlr0b/XSD7TbM5g5JBJhzrKqcwNnu7eBS
gaZkmkZKV5fqPwSkdwMEslrC2WblGeqcdSxb9UjEVR2Ods7bLn5KW2aOxwGedH1Y
azefjdLJNANgz2oiUjovp+6g+JQAWdyk3VUHDq/loSApCj5W/nQYjHoUxLmIkpUA
cArgC1wDQdiaEySEAmNgD8dShJJJ8n7IUg+DRNPqSCGr1Sb+dSALLyVhDm6lSmma
hkeo7Z/6uL+8CWboTcEeflS+sgHUJSpU6fVWR8z9k/mXv776xuSLF68Oad+pHJU/
PMlzq6Ra/w6fQ5u1YBUdAs5kJ2A8uPHb5thaom9tchM9cTuwYwSiwoQyp6+WDa+q
QMkXpfv1+mN8AMJQCgUU+2ilVzKba5vV7CDbdGGOF/WF4WQL1HEDXWL/Q/aQMdY4
iJfAYweb01YTOQHsxuW+kcTUZe9i/Dckd21O3q83QTZ4gAz/QtqauQD3we0pe2yu
NXcx8SqP2sVnAD38Q87NdNMA1ZqUFxWqTzo3wQVKTDypaLxAhbWobmOljXw613nz
ZT5SUBHOWJeRnb69IuI5fi4bHMpjpjuk40yxPXMvAnCRi4OHcLkAxNCj6hy6tiuH
SMYFM4j21lSusTSM6VW3QOXMy871pjzm5qAZbtUmLx7r6YYHtTfdNN/S7IrmQcBs
5c+SS6ZO9YgGVaqQKdYu8NiMnyqcoeGso7a7A1IbxZ5d4e9xEJhRLL1zq7xCx4j3
R+EaQB2KG2qdkmenox/4LQfitEP74H2w15lhHt+FXCt4cXoPkY6Q/Vbqelxwwbdd
IR1g4auW6F7bdrJx0PQ4ZMuV7mhBLWOX6edssjmHlTL/nrmtbzrrHoQA1c0zWMIh
LHkpPHH8fp+n27d7dPvdAnxaMvIGyQhqVx90G7UFhHz2Q20xmRyZnOv37xecWP/H
P5R2m64FDTwWH0DR9g77I78qVN+PMwYta9m505SzQFxe6Wh03zI0qT6cps/3lKaH
0kEcc5Ol1BMHPI2vmCHJGDH5/OsyZuSq5P+yYVSvljV0lUPImYfIaEJEy6tZtRww
/m8Lti7GoG5ia/He9eFjKH4dFZgLFenJ129OarAsTPu1NL3zs8DqUprZ53QWOVDh
ZxqJe+BtobS9BCIyR++1ZZIUJSnSW92BlV2LtiVDFP8rVQZvF6hF0QFSwwAu6NHu
5Pp1OIuNZPPlYgGMQ+Z4CMsNYm4rOLefqO6hQRfj0nvRahGZ2E9CRbLFPg2rLrrB
kebI69b7LWLrRSb6Q+FvW23R/K1keVsTO9R9R3vIDid306nh3FGGs7pvYrYt4eiu
kNXyPz0FUB4nkCiD0AyIfJVLQqVKqtpZOJUf010TAwxQ73ExiTrnUROdTZwW/WXg
RwsjOsUCUjgIAyZl6VJtBvXwEmJ7MrXASwgHNEeqJX86lzLOa5jiMm1CU1bsL47e
zKLLWWyYCSoiHEO/pdVj5ZYBOPtawSxMZzsovhaF51ZuOT49rZn+o6bfpTb/RxTd
MYjBVE1lyAAeUSp+NvQ64MHg8ld1fTSw7UfLscwv/xW4+l3+o1IbmwTiCSdz9SkV
TsT5HL+fKrW8484qTr7s9vY5fzN8hlKsUZ1ti1xKsPAn37XhJQeJoZ4TQGk0cmvf
uEv9OAoLViV8Y+g7c6yegp+srn3+1K2My4tmdxEqF4mmqTk0i6WflQAw48jp5N6g
a04dQXA4B8T3dxTe7s7Qp5CS+1VHPCxwJHh15OKCdDFwshKOGCzf1OtCuIswTmXF
Xi90Y9Ah7CZdDro91oU8sHZfROrhmLSvjHXtl9txJJNGQAXxQ/L9gU/U4RCLuCnv
ShKSNydBU7RbAaYdOhCl5Ij2TR8zmtx4diaUnHj5oNIu1mVWLIazf+IwaDh0MAMR
Rm6tiOG7QONBdd+I7wZrWp8B/k4Fu0U2N89nuRQpAlzbaYjBc+/FZUeL94OO0PIx
XxNXMrMIQWtyQReCkWUmO7+jQwc6lziOVOrMrw58aYvadp4LQDj/7DvoXDW+8aM3
JcEaqHqydsyZY0ahhRVivQdi2bNmRWRUv3DPojIWaEMyulMyJtJ3Lwr4aVGp0W4m
/K3UiCMjmH5uv5DGbxQbx7bevtYVT7LrFDNDLywy/luzQEoDGB5GzxKr8xTUYPoc
3ZXEbBg+Oqx/VouEJD5Wu16s5g98XSGayJCcSB7fLmS/YODPQErDiDrrYn0kObYm
U7BW+a93708mrAzZGLHwkY1MIJCuZ/FHVY2CfTyXRRyRdjdDP1vIQVVRq18ncZ06
eJHJmH0WtqJKQoWCjFVHFvYt+5uB0xlCzcit2JtNl2SD4lmpXv+deyewjoHa0FoN
/0EN37YkHD/7NNUsuAW0rzFJI1lqtQ6XRK73QfYqhs7GKN32n57ekvE0Uo7Rw8GP
lkiC176OwOplYQgA4FN29Gvvizua4oANwsQzJOyM8BLzcHeSybEoRNi0Ep6e6qEx
OWqsophMnIS/6b7qe0e1AxP+lBRlWSQUkV85PQZVCkUndPyDEH4TbsrY32nJ8Sby
nQuA6Z7OuILSJLqv8zLijfqCST0BpR2de8RNLOpXAj6KB9PkMmN+X69Z2illlBgK
VMG9TIO5bzTiM2ciqxWwnLSgEMCeRY6lkpoSY7SGpH82EpZQdfOFBndcwBWN58zf
VEzYObiAAdGerMjwavaD7YhEnMyQ3pUkgsBCNP6PZHUY6YriBHmXW5oJBA0yAeOG
0xffLGNdLk/UbGogT++9+2K8Aks3cU5VmXctqJ25N91hzBc2lbNmLO8GjIpnNYN8
PgZ/a8yAAMUN/VTbIG+p2UgLVe9JceQwfRk/daIVx3blkVnGBIvHvPsIIfhcg0Rt
FPttplcaMji50kvvzkPUY9zVNSmVVW0C9PZQ4gT4tJqZRpVTZDRd9tfh3Cs7qNO0
5IvqurEcQIejQ9sTMGT9lQWMlUVtBonZH8oI5LZTE+mMYUiMmqAXnOSZ/BKAT3MZ
iVnQp8HJpWwq2TQwKLGaUhGSa9FZD2uFfFtv807/n5sA5FrVbWv+TvEj3R7G+7CN
ZGh9yuCllzLe79yWB9AZBFut7k3sLctgvRKkABc88rlIfLP6P30cf8FVCjK+qtyy
+GfUJSHIcFxsm5USHxXGIpqtc8HUW9ykB6S//FgZEjzM6dAc7JcDfYYOca5qT1CC
9r0nntipQCKHqgzEqpoT3n7HKWjNyhvCl/J84DOHKZ4vp9V3M6pzrfv69LKFSNiT
c2w8SiqHqjXLlDJ723uoD5OGpOlYpQ5jXnU2VV/gbggvFnQ3Jvlmep5NVcgOmi2u
f2oyxjT0fMS0Uh/YzR+NxL0ukVSERC4ENBMKxk+9p6LdkFfNLC4hWpyPWbBlqMqP
iRiKjGaGNhq7Jv2fJu+MEo4GZSlQg5iZIMTdlpdhZMjsvWzvr8RGQOz/YQbJuaB/
efiYKuaTOLYFCE/o8Fx1IwVcg4jsYiVko2zHa2AfQOXC8tx7Q2kCsYHoA6tJo3UQ
Y2ryW1EDQk7RshwwIc5EVI5ACJVFIzMuyfijgDBe6s1YXh3zP6Jjj+lYBgqFJ3Z6
z7+jBSFCwtt6a6ndSWCL6QRd0xw9WnvUXslL27t0bb676C2Jft/aDo60tKfkrs8u
9mucYDvSroo3k23xUJ+4prV5NytBGrQr5jqT/+rEWLK+qirtohdq9CudOLKhomS8
/Wvshp7Atv5UeeaGLlxV/D0LeY82YCe1kGzvQOTTbx5/ydFhZNGEebeXSotMzeIv
9Pfke5Rd70Yt3PHS1KduWaxnkx5mGVb87E8ypWaADBT59hEiucdVFxY0wlJ7xpVT
8gYPpXJ9VSXPRLWWz1Z5LDGg1XngRIEeguOy5VPiHW5Dtme+ANfUFqEn+AqOSdC6
05mCPGplPtNArj1QT8KOjoyN4Xlw/74mti876v5s0bkzzlsKZpnRZ4awdQwh40bm
VqtrZwkioprHI9US5XlqE2dD3Fu5Pbz/f1mn1yvWJH++mSH9MihOo0mh/XKU484z
N3zzvTrwEke1keI9nca5ZIoeULLWDGWbQgzumoiVEU1SyhcMLQT/mXtFDj+3nFBB
+MtSFuhUguRs5ft2DqjMJRTpeqmUTvFcOD2VxAgCCmS5/Vk8gPlHp4kzV1uapRyR
qTJ01XfizYlltG5OToO1X/Z2Z1oTIT+OYgSEOlkmCFCGnzPvMzlC6gDikJykf/ZE
v7mcfYxLHTDrIdCrSnU8Jsngcdouyu4fG2Sjrh656VrmiF0BwOUcki0RLoS14/GR
BJPkE2be/3BFl+FjLeble/VYSZ9DitNFKsT38JF6IBnauYTSqMEUnaVhROeMHlsZ
+kiwTSRcD3ZwIjr3bK87VTYK4gC3Sc1+PzjPToh2bkuVCp8cj+wwNr/s/MsszsYz
xpCfYS2hK2uCJYJoX97MscpHeqkf3QEkNCUZskBtVuQjBEAdMLPGgQCrtP5pPoEU
K2y8eq+Rwqa8MJ0dkzZwVBlR48kP4YtM91FB7TGr2xC1GAKIDxLERpF7AfzB0nmJ
k/wt7xMZ1dL9+tauBW6EZfM0kePES4TQDpjT+WTh6F4bIxx69kx8AQAlZ2taDmvp
r8XtvNBfI1HxqGmM5ppG5ERJYf1iVqFIlHqsqGmKH8D8RLynAbKTNSdJt/W2UQ/h
/AkFAyS8YrHXuCfg8myh4NvVF0yN5JdhZwjiGi4EPzS6lRl4wDX8Iz7GdLUUq6x9
lXQTlzzYNnN4oGOzDe8YseSrBwmiRzSNVtidtneWzNJT8y7CQvyJqhYKymGNbvZV
zPtpvFMGS9OIyhAF9DM4vPD2toQc2CSJzNBH3jUJwc/UPvRmOl+kMhEM2T50578B
lDLaZuYnY9k24kWLs5LIWspuR90Yq/EKOiqUlAA+cMvrcYFyiWtkn4ybXDJAmjOQ
lsQpY+OVkYaOi40WW5DRoMgLoS4mwOT7D7UrpB9HmF8YHFsm3QgGq3lNrJmiJOhw
Xpnz4VtF4U7MjrIO/JtiCc7ESOYwIsOLMvRHhNBdyLpbCk1bqji5jpYft3KXVD3/
b/2V7Yf+nmrmURI4gIk7zds7qh1CCB+U7Zl86jYcANgZE8dBdRz+tgh/QBoR3mkF
5LL1AYLXSp/r4ePvOTw5uaKBQJNIUNS29G9OlSMVTYAodC1T4Bl9RzqEaEFQ15HK
BthcO/k1N8jQcXAgej/PW76A5Llq++EFUzJK/x+OR0t8xQbgtK51nWIdD3Z6cIg3
MCNx4e7k3Nh5VTmfmGhiFe3BK67H4N+afsvB/mdXl/gE64vvtck81Dv3WrZYyf4j
ui9fekXVDdSxpJ9DOl9diZtWUOdHBfEK8vNWdJ2kOVfr9C9WT3449sTArz/B2oVI
O9Uqy83aWTKRrbIC4PB/RJpyDPYLzjANhm/fmtufIKEe9lVJkgKjt5ywSiMUQhwl
hDlIcLz/Ht+E9h99gGawHaTL5JDX12wWnwKm8aplLVh6Us9EcmHHDtNMC8MuvukB
nxHDWEyWHii2Diy+569ppR4bmjkqRl/xY9nmBjye3QqfYI9vhS/8G645DPA9cFSf
yaprAQw5Q5eIl1UI2/fr2sXZdNauv8CecdLLXivFBY5mEiV3sCliRVMhYdJXtYPm
/j+oXx0p7fuXoxP7rMbLu/LvkkTvIs5jE+upSBCzF3/A/CdB3QpcA5UQQwMn13Kt
/Wt8AvQFF0luFChbDskacEaMTwQmWJggZ4ErWN6puwnphQPHvNlJexA94fT6veW5
QRxoBV/nG4twHW43eXZ1GQPFv6EZhQVZwBB9C+aTZ48a+oy4tFS0rX3xPhmBl4Ka
+qTZbTxbc9j2ZAOU0uATkZhcFWEjb86AL9WminqHvNOoqGjGBoHJsmJkXZdiu8N8
gkUOBpxAoxZnEbDezdNBXVad54tAezUAk6HBuu6BSqTqrBf53VATlmtsB1jU8AEz
K+IxUuMKu5lVCaC2/T+E0j0Ne0U6eKnhLr1EyS95qogjRByICes20SJssS87tFVd
jpRd7STiMkVOfh+y0YoeP4CiK6w5DRAcdsmp9oCFkbYJZ13GTSSVC8acXJgbD+oT
NopgBQnRSctzhL8+2mUZt+AkBNX9PxvYkTj2e7VcxJWM6xtGEp/2qTbI4P4fey1G
Tg5dOf4hskc+cp9OVHB92eusVEesH6HDl+3gsT7B+3s+9gqTe+zyvmJhavoouzvd
Z7se8hPZ1DugO1cfFMLmz0xZJVvnJ93jJCSU6OA6Kk98O328SbI4o9mRJMUxOnH6
hVwbq1fa8EHVCKZ4OX0gz9UMuZ96mzYHN6qwaV5pgVlk6nnO5ObIkGNuwwD2C8eL
/FcDirIlvhzNyiTYdZbQAVhIAApYBQKMZqENrljAhOmYBHQM8ETchAbFUqe3dpm+
TRSXe1WcANYVZqvh9AUgF9XaLX+xQWfuX6r9TA/26rb7uutLtPeqojfcOMPJSfrq
WrOmbFVdSK1ZyKLwbX6xrb0S3chDw8XmaAj7hmpNePivPQFewjBsSZZvyJON8yu2
5GUUkyJFunqcUUx5fdKPQ7UWWT/AoMN82oW4AHGI0p0SBL1VxIZnMi9OOghY7Cc6
cGAhvThkCwVtqC+tp+spO51iyzIG+9UeEeE2OTpQZL2ymu6XgiQgs2zBzpigKFba
JRF/PX0CEKd8IMQoe3z8WQrJXGZe1X5pqo2Ub2jxLd1LhCS0RMBVLLPaCaHQgGZh
wF8mDT2E/UPBzF9nhXvlfuvGVGvp3xnH0CcrC/AaGGHh0MF05urGngu5mWpAY1t0
CrcEY+cu9E9TXui4Abjmd/S7DZ6pgOVwdijbTgxWXwS3422DlhlRqFTOJI47YD4H
VlGX1ys1yAG1mxtVr2ecubqyTrmrjcQFi+yJSkKcDgqER9ry8SVV99rF4XTJTy2V
qRlmD1F25q2sNmXC/bdcdydn2+axJktNIa5yyNKrxlqDbA7iKwOPO9g+ZXhljm94
SICBAEF3tmc038rQeEK8kjCme+Oa+G/NX3gZWPwvTUvu5Oca994I3rXk02YYnO0K
Y9Fuk5A3NLrFh+vMHglhu1TYp23+ftC7tPHGKMdTIxt/tHhI9oudgHJ4vlRUV4bk
P3e5NlOeHG+kynKklDaJONdzwufh3qeFOigRaEwoWVMKFrhZonBzl8j/QpsiOA7F
oeQjSGA+kRbR8uDujjSnAVxOmsCY+zCdCPxsy7fa6c3gLoKudqBg6tIhufsg7Ojs
yav/PmvvOBJ9Ee7Ii6E6bBF55lcK3KiqFpe+9Yt9eEkXzeE0g541eOrEb7GHPTyh
zqba8WBMT9o5tx1FN6M6l7BUgQCdzXGT+jsLEW9zQKIYcTAUF/nCtgAaUQ2A44CH
six2mEvUwO0WZ0IKLP8R+t2H8mHUpsX/tyBk4GeUYhhQq8fi+na3tgcrdD6FEkZw
MvNLvUzCO8IetLzIWHvffpMTNZvD/iXS2c/WJ+VgBZLhBsrhVGrz7GCp7v85T2SO
zZbYL+EocL0LfVuodQjuuAaeT20D2vsKpuLnJJbsZuqFSircg0KrrNOfBbeYm1iK
kY3EZBtj6aC2JKUVSKDjgc+rKHpXzdEWdPCMnOMaZ5rG2f7ixtGePqL2gq3vNr5X
5yvQaPckdLTMWusekx5kJgydAaynDLtlLIkNZpjXmuciS3rbN/7S9FZwYXlj5aJj
+7ve+cLqDS5eKAtsr8Zr7pgVOtp2wbvIwFemS4Y5lrv0RmBua1vZXvT9NxLTt8FF
9AXejKn8eW1H+P0SuYMygxSjDBBZk+KudFReI9urJBZigNMzbtXNluuoToZg2Q5/
dgZXUIObCeKtflUYMtxzVFTtItzhnbitDfugDaYUy5jmAGrznnCHcs/jaKCof+D7
E2ZRn1wGjrHOy6PepRPo/ir5iqc7xNwbPxgwr2xd7rH0K/dYWX+8BBrj9PscHnAN
N4g8+Bkx3MSjt9iup8TgfS+UkoLBIsWVQQ+ATPIFgtv/qUMCYv/+jjLznZqWTZrF
GNG6JcnliN3WK7IkTLIOjlR+YPreq7mEMheEqSKfvcm/fI0RnDQozl8hpLaceJGM
xHy9tV99XizHk7F3HnQhkjk6lRtBPeG3CYCYmom5Cth2oqszfdGrjDZ82KG+GrHB
dasRtHXmKBUX4BiJpoJSNFvC9nHDOx4wfLTtu/2S/RbAikE1tB455K1VTGvqWjyb
Ybd9EMliBe0C6/Lc9yZbHo2UHN7mYZsN6Pj8M9UnOEdxpZzLW9T3pT5rqb3yQvL7
RiqXdeh34dZ8m9l4skwyjEt87J4pvpId6hDK2R3Tp8Gv/wM00jbiX23PjdxmeXu1
mxBjlKcW8lKTW2hqZPI5kZrnBLzsvK7j2HVMMGmoYSHK/jgY/aUAosrTvtjQOd9H
6WiUa81GbLxd/P9XORAQWsg16N2RTKB3oBY8o71IcPU/rFlORZY+nPhROlZD8bDh
3hrb/9J6rKDQdJZwq7IhK5TeXLjqVQd9tJsXF+lJosdjPxk3M+YrTo7WAVhv7e8l
CVAyLAD00b8z4Hj4fYLA8doCvFiZZXLAsy02bRFEQQVMj/XEEG1Bk0dm0QrxBZLX
+aReqmJNS9dBtx95PzAhBjLI9unmOwKjgLt8tcw4ejMJGG0jVcFskHnZjMRE7JKs
mQqSh6A9WQRLMzRoJlzk02ebI2VJzHJKeQJbnNbgvMyG3h5FGDw4XEqKawtJNgEd
lafqhDIBh7kjdxlNJ6K5SIho7fVca0702cH3t8o7VyhPQiWi9+lDCAhtRCB+9cv0
JNNi6OaFDWgCfzXO/U75aF88uwuZOtit2ZD7xUjGqE9xDVa6peGn7Uz/mCH7NnlE
fn6/0s7LQofzcox3pR0rHdO+dgticqGOCJ7yu58K4FETHatGm/HhAAcnh/IhhFsf
//wujlQ4fCOHcCsvl4DjnIhMWWA8/arbiEbrqo/r4mz4yFfHq+e+xgSoVrvhAOyv
uabYWWbt/2WI50KXsilKUFu/Ki5ytSv4fXOGVzJXDU5kt5AANeqHfsv1wbCZouK+
20ZZQzi93nrV+WJQHKqESlMCJ+HOpNVm8zz8JEhzQrTZoOjltV4gr+3GosQeKHRH
xG0ngZlFmlj5oQGtefvCPeaiSbVxjAcONhz5rBwH6vgTqViK5v5caf9k/EFCUQoW
kNhRDZ5aPQmVIqq1ZHKTzdkxWAlwwKk67ErKsYN2sxXUsMpKT49oUUDw8fBGtaes
fhAMMIH92wQTZD1SVSB0q9wLNhaFg4utzH4uLQTiXt8zfUulOj9yGW4NAPR3JB0C
5yvAUGzdad6SbmOhaMh8979Nbtdxcv/meLcj8mG00HzRPqTqbmcH/TUIPpez9B7A
z/4NQYYzmWNVxDIw1aiVuRX4WhsbapKHi9T2zGyqyg6CLEvpr9HtZqeRtj6Ob392
nJkUjqSu1D6FC5UCQVtnlm9ZJYOrprQurLsluYoJx9YEHheAc2w0t38etGrwpgXG
l6KGRYTjcZwd8Sfp9gLTjTAQrz91mgQKhH+rrnjWDrOlgPY6yHfoydugJSBjru5f
bnwhJPzOuIXkxQzUpf1YcB29dbhvt97kondVTKbQyWsx8zbHFKCrzQc7FRY9FKu4
VjGhqqq0gpcbAYRN/2tZ4Ufq15GzV39WV8x8/co4ul1JZg4vv1L+hmMil/Vvf0/+
62gq100D7Ufb0oQJPWuPK+98uBnD5YNNyzeSYWASFIYZHehs1YcMgjBEHHYxtBUD
roE5VOmLGUqr7BAqZPbR8UsSgS+yfegYOTZ6BQ1o7GoWjmSCX1urlBz715+0Ad3t
mUYGmbq7LtymAEopqh6RHLnZ8Lh2gWB7pi8ICe2tS55m3PzElGgTRaw8zxk0xW0L
BGVEHh6Fd6NF7/AJgNjRyaK9FcxCmckl/YqvgysfAdUmmcBBvFv5D8a+1Bt61C7v
ZJdUAxx6kJzCiNEI2OIDzPMWssnhMDtJFvOeaA21bf88E4azDCi6U8zNmTuJYsfK
iq3txoyIz6dRvjCNTIbMV5/Wbo8UzyW8w3Ncx1PiiriNLMebekUNQfy7VzFdYWlt
FjQUKyCKVIMgpfRHVxX0qm78gmGhD1mO9hCdLm7/2XulIQJZNGD9vXesuiQgssW0
4CXGKTIW0anAXk63BgIGy4aKHM21KplN7ONxRiW7jVn2WBp4bt8PI77shp57tBWR
VaVDg7bdIribSltpFjKKK6aXjUtnVH+hXR7Ee6Zsc580Z41pL9qTOJkUTVwxGI1g
Gf3GKpHpKZQlviKdTO2fV9WpnB+EkqdC3tQX4Pw4jRz82XtjYkwgJ01vcJl4JSCW
R7pe+ne8w/0xiR9XJKKiIF1CguGkFsREy2EBw2CX65z3rBjwxE93aFEpETVb21Xk
9Loe1tQJFB+xmMB4yGiVVX7sIUz1M+71aUr30MzydRB5N3ACnNtm7kHApAG07E1M
7mPLJzaikCbSZNFlyQtUkNXgx0cbNQcABemZcYkQQHUXFDwWzSXG494CeiShzFYi
de3qzcZkyWqkTad/rWnDM3T8+s7HF8PIUndnmqtwESMW9lG6pJpUgbkl9roifxsd
NVY9nJLQEsXPg+dpzO8gA5p3R3c4TyU2h8KFUvr1CzxOwLUitrO8I2nX/W4kHeZW
fUFNL+ErKg1sbkZFCeZBL0pyUnluMifh6dnQtAixIJFusbmV2JieCdTP8HZLun4U
NPAByGy3nlu43GOtuZzb+ufovU7ZE3kvn6enAglJrcy+8fkRhXWqo6d0W7lXVy2+
udhw2VADCKv3LT1w8UFbWOP6Y+KVQNfez3Fq0v/ec7v4eopSu+2MZuGGBLbgrQIj
s6Y7x3eN8rvMdFTZ/ssk1MCBc90so935ldfBMoneK3nA6p3/SChE34DrdU56YgQz
EtZKBosMGodg+baOVz9/8iHSn27rJgCJMEj7xNJNbuCeG+gyvTej1XITr6nbWIQw
lMzFFI8NX0nGQy1SYy+6JPOccT+vqxzQYG2IndFZfhSuREg71qOINJ5pFKS3Ou+i
mj4rZozB71QlfbvBw/jMfdSSDwD+GvxZid842dIcM7bEZY1FmcEoyeAt4cwzKJv/
NkKGjnO3h2e+GC2ZgVFMMv9mxckLa9VAkvN3iJaLPnMxyaHx1O6u/kfhnCCYKjyY
wFY2/ZOPTNHcFDOnwRDcD1B/kKu56VqwUcPvBVUYfnsofgPAMiGZpmT2C1kE/yIh
er3sPmyI+mE8NdfG4D6uP9QOQRwuijaNiaf/qnauBPytmLRQzQgCsaQ26rilO0gG
FIUpvgjgp4tlZlE8UUyLgSPvmiO776RcZj/RjPxaE0DjG8jk1INlZyCfiGRH64/8
ZZhMfS88VhToVoC8kA64M6plP38JmbEsnngOWuGGVo00BEG37hzeQqrJUDL9sZff
rCpnhO/GGAqEDuAOLRH84zYHEjq2p4Ollz0PEEuoAjUK0D/qCRWBsQoL7tjGxlLo
2VhleDCYZhkOe/ifZO5dYiyPZAtiPTX80LzxdhzcZp9gQeKQYgygqxiCMR+ceqiY
MN8R+DXGk80UQKNgTsa7dm+TdFSwxYYcfIZJjQQYCjEK0L969dk5EoKOV5/hyPcN
GrDPJhKoPoTK3FX9VUqKOcCJkaq8lvNlghgyn9B1laVNw4xYD3ETwFTUcgpR+JHo
UCe6/O2RpmpqmzWeqLkIYpGEehNOQt90ZG7erxB6p2qdAoqZe+90AEgQcIsg6bkp
p/rwZrxSPRtZsAWVEkVGARHapblUx7CugAIY3XsQs7yQgyUZC00vj2NeGRGGSwWv
qVQ1deDyq9hYZaawP5A9bMqx9itK9+WtIIMAaoxFnIE6MrsN76HsW3s7SzUfR0ie
b14oc89ooJotQTzwac7G632G9FJ0xf0ftnOgB+UbyoN/cyoeBVYMRdobeBqU552w
c5dHUnQdH+redq0dKPHOWjqCixJXalNx0PANX2IWUV4k/fIbkDN/4nhsRpqQCDX9
3xPW/Jvb/vfNmlcaYmf8MAdcfAFHOAINoO+uO8oycOK0XRlljRpe74MM8UE7ibIn
VKoUgDMMv4wCUfwgiHB+AN1kiTb2cad9enT7A9FzDMQYm8et1Efd9FFnwmD43zbP
A1I07IzYKpCvLw5GFa/t8f2oZe8g8nyhZhKWdIy8j7B2SLKy0edMajsN6Jd7oBAq
UqYOKx2lY9Bs2c2BgvtTMB/K2VRoIHNfIo9IetPZJc/qgn6eG6xf97+/SvgXT7ID
PYQCDvJwi2LurA24/ZB3+KZebWU7BP+Kwu/5aDNp4yLqcQoeYBK5NNrlfpPqOdf0
rw3Ih6MGpTcRfLsPBnhDVt6LuhXsV0QqPF9gVJi1QpN7OPFwoDQjI/2m0ZrCnu8J
osFsb5FPbqzBA+fgjFrsNbTiOLMJe3GTSXl5kQZvMPLRhCxatKR+SV2onvPCOAhF
288dED+UuXl6euxYUqx/HOjwgIXpzPclrN8aQsTySA/o79LkWzET0JdCJzt6KUen
PtVwswPrkL+1PEkDQA0eYCdcCSGtgiLy3Lr57skUR1uiFIfoyqwvqtPXicxYjnKn
vFRIFB3nkWglRlcFL+0le2NkrjDXw9QX6bWNcJ8WtWYD3Ii6yz/3pVYKiRrWAy+z
Hk5uqOR979HqncCKAYf/fTnzh0yKg6gfJMMdV+I5Jw3eBSv1L9KxK6rscrz6k61q
KLo9pmBDo7XcS+SgHXUHsVTK1sd6x2VJSSc0zzOjteI8Ub+/1s8zshPHakY8FgIV
JRE/vK5OaB72PpT9cXFX0tiVYiGB8GPCj9TTRPY76xjxq/2PINqIEZSN0Vx0aMrE
WvbU4ky4wgpAthKQCbcyppgOYNqRIkSwEI/YbfwUSiwZxAZaXkqfAomSWPPTqZEU
WFXFtOTKsSMLDpA84hMkJAGBL9sgzPlTbi9OBNagzPmBSqEFBrNODCwciVGOfWe0
OzgNcKdtdjSEuiIA9XTN8mK2QDYuyYSxejuUVnX6Aq0NVuvoCAD3DDNvgSvSQ51l
nlEjAnfPC9fxdPixL1TtriWhN6L0yaRqPQB7PS76Y51TyaF5XHdPM+lZy85hDe2i
tZVoJrZCL0Za3tCchJvQHb3tnoBAyCFOTeaZnGG/xpA9JSaRxqZ7KLVrwY/Cqgb4
ki2Ma4vgWEPYd5gZdfqjSQNZa6+H8I/IsKqADMStk0vftRpCwph8yN6JZymfgm0E
q5UfOe+c790tEx3fh+qPoqIIksMUI6FDqFSwtf7zzxy17jyTQ86Q8UVECCdAKCpi
2VnHRPRAWlztPtLbcgEeKbGvWVYKKU2YzzTx+ADbpx7vs38p06eDCD79lVG43yXD
ueO8Ir0TQTDu0CnoQcpk+5/6+T+RhnoWuRje6y4RbNB8CQc2TYP6ab8KaZfOIz1E
UCzJtFaw78YX2ZDIAlV91pe5SSV8vYczX+vruW/AP8HShpkDs5IbEeiBQtdpZp5s
k7Wo+tHRs7p08OQTdRlRfU4BGczIZnE/+4DbxVSZhCzA2sNaV4wXvkoVEai011D9
35VWc9E/TCLv9CC2E5EP3V1dvVH/RUpWfS2o1NJgspvGnwy3tLk1jbGZChDkpQzW
LiNsr3EIZFKmx36930F+1N6D15us++cwkcp0GtzsaiFGvCM2wD/uX8BrN6oZdqlA
Iow9c2wPtGDGla7r2f9tBBuvGg7RRsuVFhKJiKqoMkpRQgQUGPFZaN2S7ircSq3c
xrBjn2WH3/vF80HA/Z51X6ItlTJT8o01z4pQcOuy4QnABUfrSusx8optyKfkpNAz
6yYCee167+Us6rchRvUBrPQcVRiWV6NeizCbCDt61kDwWAeNQmP2XVH1MuH0Gdrc
44N5sPjukA9ztvtNuPEKAN+Msj2+QXDBa8DdAoNcskaUsMzezx+COfQmkRNKxZJg
Prg7I/GG3GadHFY2oOiUOzZS9blTGF7n1PqBAnxngU12ZfvtlCDd7qvoVLnhK9/H
jzOVfTkyKZViSyzWQu0MWfK0APNDker/QFUWHKrgwKzVrRYADZPHaWLEdlJE2xOo
5wVz27pzGUQQ7xi7fHWvxOanyig+9p52OqlAZHASrGtMnnUytZ1HpM7lrWLfbwvK
Cjj0Ue8QBr5yUQRqnnlCpHNPp4LZMTPxWubw+bJ71hHSiVNmiIxm+DYBNyeNmaGg
FKlHbnOk61O/kDtrKXuoZk0YfDBdGtlBc+M7TDe6jQ0fjXEkkslE02DbmAPbbUEW
oIvI7dIvLKqgJsmwHK4gChlX4NzGsr+UIQdt2+lJPc+zToCMJ1RMCbi7RD92/3TS
uoZp0DaP/Xw/vNpaTqlkDRzu4svMzCEBbD5Hv3iyUQAL8E/jWQ+zPNE2OPnquSsT
qgANkJ+msvJrdIkeWUnbfCWVF+5mjAHOMkikpbPyPXSKZU+miFoA79q2J4nyQ01I
Z6Mhw5ywKeMHg9oDqnHtGGU2aXMdCl3st0Tq/XGK78SH4ObXJ3hpAV3X4Y0enD1a
qR1ej3tVQs6zKQ+SirulrE+RyHw9czs058ceEEBBFjSAhGghtmwUNWgBsQnY68dZ
wmyQAVkDRdB0rJH6xLdVzUwgwPI3uE6a/WLavlwdktQWnISZMp+o1VH45GpJruOB
9o9wXqr3cJOpnH3KOAzCQraXaqYyYFzXLdWITpeOYSevImYwHYVVKmb66e4m+3Jw
TldAzUAxog0XpXZKk0CsYdmK5E+7pL+rOfdQ7xAF0AoCi2D6t47+Q2zhi6twPla5
vqsQbeGQTXhv9Ujn40DxoAUWgqnobQwKgtXYWFFsA5UV9AZXZiX8AgMy8v1ED/4r
AABAegEDYv/XTvK98GMbjTbcrg8L9tD6aV14gC75AU9r5pY5Qt7sJ+m5D1/uNvte
CYmfea7YR/dYNtOCuM3uYzGhH1rBasVDmkvzxkdQ9HqzuqXM6QAMwNlzOYtR3xGe
z8vAI3jp7AWh//KTDjS6T/q8BeTNt8AnkY5mNopIY6amtT1JcwrRIUo/Te1OOykJ
miGPZ0xf2ilRIwGP03sOaTvFuVlCk7ftMrKFdt5P5SZlcJjytuJXAW9KA91OXxBz
16Aw8zHiTFWK8X1XQGZ4Oa/1DMkYWnq9Y74kPwtpu7aXmNvu0auUN7B2zHK6GzCK
YR9NpTZAKgGMtpjIjbSIECL8Bkr9W7DwbEGvRUluJHNeHfKTZ8kmryI/0OiO4Tns
1bKBwaG8R2o+D1nHrClmuE3mdnKz9a6PgQ3MqaL281R1phwBOL2CY7Kq89AAV8Rh
Y5gRNDyl7su4rCtmBgy8/X9zAsvbQaB21yhtDui2AMTQMTs09nny02ZyasAx0lta
eGJ9R5xZznQM+2bx+lgDCnVzUGcFRfsmYhESaSdPONfBHdaaafdPBckMko4Wx4TR
AYh46SQVkwIwBLfqrIhft4K8gyrIiEQ3eR4xbUkDmftKp+9z2x2Kkw97mg8MrVVp
HFyGC+FR5FKfAGAA7VHiIvdQvgs2pkr0whtTs9s85kDWA7j+XjxdaCVNknwUNNL7
JLWhJx7h6rpLw9D3OPV/4+SOvSPk8oVhT/X0duALvv4Z2snFgleqk1c0+TkRsqrM
rrAfnNMUekrSBENnadtPrShrCorMqjGMxbV+aD0lyekJq9kAbcDcS6gIa/AAncMz
dpWP4yccK3cxKeRzZjYeyrJgYa93SxnbXESr/0XbI1Jdca+EWF6C6DO3cfYoXqJo
MqY2PZrmnv2lxqJBp+4fpJ20gNl63Qa1gjbmMGa+l+EorqvHpcSoRpFZzDtj+ou/
gt6ZcdvSyCyC/EKUp1YFWuccdH5Hnt3LRB4aAzxO+euHQWA2iOWeqXzZqx5QCduS
CMVPaiizsXQaoUnempyYWlmtiMvEnti2Ger6ot9WtQw57VQllL8elGFVSxfimloE
yMdCZ5ipnLiKJeXMWu691CA5YcdmS2bEhDIhBpz/f68xgh9BfYIVcIusaE/giPRz
JRfNJUVcxZEt3m2G8wVgEOgji8FZExf/KhC7SXJC6mwpTQ+adIn7fApNGIa91rVF
UsMWNnE5lOtrE/hDjjsev1v8MdQWXCQxVNlbmVyD6cX0D4iK9iuqmHJUKI1rszt8
Eu+eptHd6cV56gfwD5nL5M5bhP2w9ZxSGbBNXlz6/fJ0pLrIrdIzeLxUsdMKyxdI
PxcXqE4Lf7QeIrJTWmAjnCfjZXE0TSDLeLjuppWBkkoEy/SDWeC/VFLJGtQ5J1Cv
eu9IhFZ7ZczVcvoTRJVVisOvEh7yfmSMA2OT/gC1fW7bm9dosrV+7gX9+wMnLPDk
Jf01fK5LK70zvVmsW8A6R/Jc6Giw0Y8D+8yBj9NEzwf9sCOSqKyoqcb6nqZJLFGG
6bLLf8Sv5EK5vUx+WaqLKKVhgJI2Hxsa+qWpz4WkbOaaLpmOXUZkX1oJE6LCqhl6
v2S1Tbfr0y9a1PFEQ8QYmw5wYqP5n9uDHFWVqKzbheOZ+nCXqxB5XV13dmwBAoQa
tsN2Hu/lweENh2KUnoLzskFhPuvfqBHd5P86IbOEWJCGKK2QZQCDEFjQ7QQBdTwb
KJMfoGDNnPy15CzKgFDuCqdO28GVpfMgV3wfxZFXjoIDoqypX6oJQPQwURvBdQ+5
P+enBdCmUrPaV972YcBxtZzFXdyI5SKezBLvGUr1Mlo/5KU4dJaWG1NZ4oiSNoKU
kqP5MaQX4hr7WxyBIEpVE51wzSQY+lXTqe5XTo78R0Xrt7JCktG9orQwMN7KGgf6
LLL98dsewk+HGDmegOyeKy9WsjyZrABjNFWbD4kcG/83EB+o0iEJj2u1BlF9nS1D
er034ukcnu2qROsVjYwXyXyho3PCtaCrObgKFtf7AhuMo8RUjhowRWhD/lj7YMSc
ZipV8FI6Y+YF0ip9EJVFpFYdHyYttYEd8qSNOl5KlvaCdXUCllfP3UzJr2HZjy4r
XHNsp/v6fxRpBNGrS26ZSFzT735xCPX+Q4BHFgiYHf+EA/p5v+w8v2LSA9it6l+E
uuoJHPZ3v8AL2RK7xOJRoGFUjS/+nZaKdg9oORj1iZ14GyVASgj9ChxGjNON+4Xw
kQxdzkbRXuJk7PaEDVbsgTGDXmj75+5pUtb++iuci79bSmlJ6ubrxWKd0ldOjLET
uV8ALveN+lKABJY9grThUvuj3Iv4QIYKnXi2GO8fC8NVAnShC+33CymAD180KE/b
LTg+ZNShccsqO7vewO63+78IYfD+qRTonM6cKYwz5gMrpH63jlYlVkmXymR++AhD
b2vBY2ZhqhChpzT3aWjKtWzDM9bR6NyhMDwGlWX8e/O7wxSP7qhaiLXn1hR0C6VM
qh3W8f86nLEN2BLJebuUwHdHun2oyh1c1cxFQwAsen0w0aLbleUkGzSZZjzA/6Zk
QKa2Ej+yT8mbYs6RNRBzFZX158mSwHJNOwBuYVN7qIbd3IzLM5o3EBLL8dsR2PGs
IzQE+v0/9/qF1Go2ckmXe2UsCAd0vPm4QnW6qrPTC01hehw7Qeng2ZVeya/HSsVG
FM3NT0W590aRq3ZreaAsp0X6038IuTO8qkBIAKvGjRbDs5Acy7goHOFD4TyQFqb4
V9D6JWkBe+OVvmeQtTdmfdPpb0tH5urJpvFqszFHZdkISE/8emxC5vKRB5nDhfbf
Hn3Elt7u3kQBbYGE0g4mQLLj+tc7h+bipQ72i3jX/8M4jltgJPs8UOTxiD8Osn0U
IjkYxZup0lI+BYOgDnttozWwkFpklh+gVE/shShwAlhzZicHU19P89iyy3NgYvIM
lIDO5t90HhNGyxnXQpQTmp6bfMdqNAriAyleLrSKDvtEBtprnfTFsPbiSzEOZ1CX
15SW4wJeEhmeh04DGFLhowUSALXd71pJVVGs1hKrR7sYxf362Na0A9W6UxADP5+e
tyzsnBKmGOpFAye0B4ngE9uy6QUAMO034EbTowtKmZmkQm8OBp3CWBg96mn2nx30
2s1JLHzWZ71OqQxufMqzQsxPta5mbK7KhdhE6Y9aX20JxiEqNmt29EKUXWA4PktL
4Sj09LyihR7Q+Pt8lSl7nqKBOhZpkU3gAAMi0nBvmyzSM0fhFdSS2y1CrZfKzA0n
GdoY3YO89E0R/aG0kTl1TkL12fUoFyNFpEMG2v4IMyNqdlmH89wY11neXtJvj+J6
6psGqwuq1EDvvy5IzrPJDeuCYdTjRrWmFYgaRZ7Sy95suqS+X87LyW9jpLAoXfxM
Md3wFqykOe3igeIvmX5BAsH0TUHSZvbvAkzLQsRLxGEI48s/a98DSD+h8HgoaDUz
/lDnmEHsmQfJOEiY965rXBWhkRBpSquQbN1kzD/nANb368qUfve+nvmA0mu9V+BV
ZdViY+eahsLi90bTKOdQTSNEvKelIvMyyOweDrMQ3ktUi4aPmli9+Q9cozDngV9T
Lx3RPIlJryDzQtpqAciwjKef8GhgaAqXdhz0MaNYY+9ylKh0FoBiqJJMNISA+Von
vc7hKb0lUP7WpFLVlHNv4PNpGobq4K0u4h9sJYJlYrAtahQz1/PEXPbDMcMmWWs2
kGdxVkGWMQ8YNCoS5jDk2cjumGrKhdh+mSzEiuJHGSoDw2Ft6Qb/eAjqqjWpa9UI
Q7BQWlH3PMrh3UFIbIzFPMLs67bnHn5JP87etEcbZ77MchTsktC7303DVAttYsBM
k92j8FTtkdzwqNEcUFbHquUk1LMunwdANRyp9yNpS5L1XTtuYhGfSW1IxN/QHJUh
1xcCKzUBIHCDTnxUErZONvLqOdpBc8XTIqNcgYlLOYPZC23mrTGD+N0oibO2mhKi
NFsg/vGRcOEKcc5pVXMdJavMk9hcd1YO6Py3Jh1imuguXxGGjPMrPvL7lMjt4xt4
IdBrJl0ZjQ9BCJTpGRWHyb5caRQ0eO5QdxirP13PaoHITrdeatUIgOp8BG49YJNK
9MCG0LS5BCHbM82pAvJ1RWi3ThlRJvscStM5peMR9GrEUi79uBsL30NVirhX/Rhk
oKDE4ThCEMxZalFHrFfiM5dmHkQ25Ug/pEIXCY+O0BBjbG0pc5zM6JsDmb+BvOed
0Evd1ZiOo7dnA7GBZAWKVedlTYarzZunY7LavhbutQyG5wtWFMzfs6VdxW4pWakd
fQy/kS9kr+SX9U3783pPY88iRAp7Fvc+Xfnp88/nkRXEyvf9s3Jl7Vp4tpCwWVQk
i0XVTGDIFxKnWXslEiwuPFxrLXNttBGxw0TyBW+knCHBavEXs7MGWF25N1NpnVCK
fWXSJYt9ByIjIIOlbr2wDQ1p+uBQ/vfp77lEuimUuap5YzQ18fye6G3nGot6qjmP
Y+2G8k4OlZTWwwRJPAPrFJ4uY0tzc2kkkti89J80DFF7FT0ZeRq6RO13nyi7MIiD
JHQP1A77psFd0ur1qefxo3VPbBo7iB4A3tiQT33TjxEuAFQMHQ4OSkjTD2wbSa5z
dgfi5tolSDB+BGfuylKXez2ZF1KHKxvoRz0tcCqi3WHYlSrYHZeS+QHGMDodW/+3
lQavkxJgoEmlZ+wDiMX/ZCZoi8wdjEdwu+QBRCM5ljwPIsU3plwiqP/1aqEm4UzW
lb6GnuapV+Y8pNbD1D05YJojYVMdl+lUzZm91gvX++kHh1AYCbO03MbMN9dTxfGO
qE5cQGR0nncB4AV3let/feBSs7c3JKSLW056n4/veuTh63KoL8q2dka396nkfhFk
xSKg0prlG8I5PqJb7vDpb21AVdpKyPrO2fT21i2YgYcekgEGkkydNd5yC4TH5u6h
5mziEcQZGVxM05ojFTFXN27gxNetHeGzFOpWeuq7N+Uis7XlrpgTT6PuiGMa8+3I
7KIO29qQupyXrKSjAnJKxhL/lwV91BPE5zt8j6S7Ug8qguR6L/u1lPaGJPe7+tMD
l2/uH0KXN5WqMgxPFep7LLh3lF2SFspN1HRloUic8fUlRV2RA8BSqgo51QpMjXQk
J0VB0Fe/wd7UPTZEah65BD98rFc8GFI1zH/dq7jWd11Ch3a3VFOSnWpwddndtmOf
Vg8k4K4P5ti9RVF5yoUDfN0LdgmiwtwX6GaK+BUwR76IsWeoR0BoY9e6jLQeM2Ij
7GNkT7bDe5mhbLasUKpgSU41vVek6ZE1yE6kkKrWAYx5y7427/oVJo2/KD7NiE/t
hlre76Hwd6fOFMJwFjyLGwfhcbu4U4PplqEnVl+BItMG0eyROnh3y7WrUnZv1iiq
EznEkTSie4FG8tXGIhzOTI+rQKjdhKg9m1QxDfKx9FoO4ghGXpOOrHZMM2DpbSwV
L+UnPP18kGXCoHWwTS3TgYCP4T6g26iWigc5D9z3Csrij0herawRTPh2erdE6HF/
kDRbWdBHt6lyyKNRhXPZ0gs/ujWneIrctXhHpCpqKTHLj7rUs4YHzQMTjuPsorqQ
2w1B5x+1OEnSSY9BNtp95rXw4QlVFXikZy/8zJIl3sGjr9qD8QGNse8h0mC2yh7n
TzDqGwx4xQAz1O9sz0zslsmLAPds3arwBFkwZ+fazaOTC/vHqGUNpgJGGW8PxDYj
kzWPA7rA3hmBsgZwBSR4veVvRo1lhc9Wrr4hnOidAabuWnfMJDTltC9EPzOxC7dW
NHDckO1HfjrMdykhZrUJUImzmSJ5GgsvT3PI+kLBRJZJxa2ejYVrSMsROFE4deEh
j0Kk4hqqbzTeqyaP5yDdyWMkaq+YQV9pUp0CjTxU6ehtGB2TGB/SYEmLu5B6Crap
vT19gy/1jfUq7H+ynO3dxRXyVDMPVU71t3cgHhjEEB/JC5BBUPvYxzTyjN7D5Dh6
OWLtXQJifSAjncQf8P9BUdSlaVNhf80Go8jq1+fFz6FQNVaggo2uUrhL5AXt1c5G
1wDym7SsVym5a1GX0cJd99+hyOx2peIsrvCj5pktzUvI+ASbn6H7xrcnGYRH2s5f
Yb4g3BKLDSj11A9d7iCVpQelel8zV5PNWhcA4HtMKNjYQPURwoohaux5U4QJugIC
dgI3eAxxp4GFQqDFKt6YFSXWsDo7cmn2jc2LwyGl7NTeUZCEYaQanIfwFLPaNFdF
XRg1TNcJ//9hk39c6kzhTGeBEWRUYoVnPWa/N1rA5PHtNDwDNjzGm1SAt9ExvfJQ
9scTHvPXTyyvZT6A9zRtZYi3koO69OHbJnsfLAc8kB1S5h6EfeREbvjcIsKsEweX
bffic8KUomIlACSVIbm6GMrHMkLH9TtTKEhgPSAm2P+EHyvhw4uUkYfrMsiD0DvL
r+/yojDhFQp5//uFa9J9rws3XsysqQZ1DyysHwICF2QOcYBBDyeQnWLhI07AoSAN
8HrVdpz6pTc0YzL4LOGjcCMxUprevjG39V6Elf9MZZTuQ14/PC4JIoxW2Rp1mwJV
DvnqHvgUmoRkORhyXdORZaUdAKh5GgbIkvvmDQsb0/V85i4Jm0waHz0b/MRCCgrT
uNKWMV+c1x2Rc73sTlCUMNWxXab9vzXVskS5Gc81Dg8Wh+GuzRaFPXMD1CC0Ve94
nzrj3sK1mGQGxKDbAmQjFhV/cMnVr0WIl84GRksYjT/rUMpUM51TGD7U+iHcSSO4
EBy0XZm8Vu1EkjkhBuHCFmY3VKrpNuZOLpSOHvq9F+0z2G9zVKwPKrhwrNjTwZRN
fLRJDDUX3BUmDMs798dImCGuwG7Ny4vVtwyYzQUrJJ1rySZiryxpKq+dSeLnFhYP
5Xx3WZwEjV+UwXBOitFXlpj1l7HOdqAcI8fdDK/zcRZgej+KuLkeUov61PA9+lwW
wwYRIFA9w+TPQenYnrEfsbwjWrasBJRpJKstguuKcUY3srREJByE1zQ/eOVq05IY
I/T8BXG7E46Whu2rd0kX5o5cikJOXun0kbtcb13W8sXo1TervWSSI0aSmP1Riwk7
s3s1d0LaTvr3chRWLvHKQvjcCxQDfTMCX2i/vwV6k6JksTjooc23Z1MaKcLHwk4n
rg5uRHZcdxkxYW64PFYLYpNP/YfmDK6vPhF5StATybOxmanb/U1RAjfJbq2hbUMq
s5SMlk76vJxbwrap+0m5FSNSDk7JRgGGC7YTr3nnkYzpL2HUleTSUfAowQp9R7oZ
HrAQ1oAsnxAUUGKsOFyVx6bOwiQRIuyUF7HXpHqaZxnNVZdTLdRY7NSSOjeptWw4
rdfloCkxKJWY6Q+c0c6MeT0xDONIrXtvKs34Mr62zsO0e7meVqW1eaMUQcd56iKk
6OfLsxTHnrM3FolveQ+4ujI3Arq9+HsOYX6Ab1IfJ0uO2wuIONdzUjWeomvfN2FA
iHZXEZw0AzxmfUyinuapwF9dFGdxdhi8V3F8luCwG/qQNnasEoefOhr/E4+g83GQ
RRC/wpgzf26UwY3+e/naAizqtkUgeRAJP7VgG286am1ix6MJ7lSxEbi7coV9+WsS
DHLQO0qdh9Es1aqY+kncuElCYKBZN5tTxQEF3bogWKEaoDyIMqCMSBYELc05at/k
kSzYAOxUW393IP2AOBCnIJ9iH73CJ/LXBpYDEZtDpRZ/TWvYrfr9dFz0dt/A7oka
zsvmSTphHQpm+xAYRYmk0kXs0B4JZQgPX2xU17hj2o/jNG8ghvwFsSOzW0/r1QXH
JDjq0aOvWobWzIABdCtV671VNrD+qZQIkYjKivsb6Io9kaNLYNspqzOh8biMK047
oYYIEIXvggGN+rOdQBGflM5YjJBUyTjkmniykSXKbwSAtrTwbZsORj+25kcgnyO9
Ap3qfIWiik0UyxTH+iaz6YHOKJGEQxwpxbYXu+oZNavJxYfgxDK3jrqHMABOFbHI
mTxDbJB/c7Xxe+RQqzp7L1siuEzZmNGkSZr/+91xVcY1EgNNlMK++je8EvBipHhO
nZ0B/Z55YWReT1TP+hUyhbXW1n6dKlZjwDbid/U2dtrjQCdMnSwmmDkcPjDKPDXY
2ei4JNmkZSZqEkSVrHtJVDPLCs4bIg+FKKfjTj9jWMyP3tDMvePVxI1C3Zc3fsOK
O0C5vqozNI3VWEpS6WVJYWWJ6oRbvC+wXpS/Zk9NVjfURxnX4GXvHt1c0l85ZqsN
V9Cfjk4bemr1CAIDoCnmtl2ztrq9UQ1KNSUkMfmkCl+nx/cJljycMARr7K61Jhb0
Qx/qKvVW49ca/7dwUJXRgINvqZUKghJTYEov9787peZzqUKw0bgJbMCnDnOiqje3
bbIok2/fyXJuMiYuSYTPAKZTmKf0nlyENe27i2OLCO18XxOQMQecX47Syb/HDqUW
N/vyOQQExSYEzxrMl6FwmzUJtu+xBkfCQSi74u+9Saz9LCJ73V5lp2L9Dpm3VW+C
DmK+rnGy9HwMZLKf936V9XN+peEgSIwh22CMLM5XD35g/jaRcytkf4vJU+7M9XGS
AS7M0orw0c/aMZpn7ojfi1yFDOqKOMrHmN7tzUEX7BcXLn/X99D+O3N+3S+Y1gBW
fb//L/5b5IiTrHL0NECh7R/u2ay7Xw+gmvfEkLfSl8wdgyCNBNCAiYCtLj1JtO7h
1n/A30h53LOTllaqN6Gf+RRvczgidlo5gBKAEePPoaWxW/q0vaJRowPWw9YBZuaY
zxxh98LSRxooTo24TUBaMx7ZH8anr02PRwMk+spzgsVCs0wPpbaByC1tvC3WcSX6
8OkSshHEfMxWx8rsfob6sll/4FVT/yQXYJAvwwMnvC0jrzaBUWgC0pvVdD8bHkjH
H9GyrWPLHzSSWUUFwDabJvnYm/3Kr98t8iZOB1wu61NlWkq0Pxpjheyf4kv24A1y
lpuUNvVsHgQD+EPoYOUlu2f+FD16c+EE1fw2T5zfrrfWABtFD3po1CVREYR4BNko
R96cwtdAY1rzdG6cwTnUr8K04/uwRGhKILMkWKqMGbuuBB+ZIFgyEkh056YHsFNy
NMiH3ZEN2MjcwsQpZlsD1+LWKU/jDFRfRTkEwbcl7+JqdFrEIvFFe/DXnw/7784U
HKBEsMagGpudXxqAjMHlJqdXawdNRmDpvc/EaKpqonxWUSWDQ1ytKutfc+Pcj29H
t9wp3wbm1ucZ0HNRywlCGrTa47e+1yiKFamPNOmSMF4b8T4KtIUET0ztkYDpqxdW
pn7+IkMj40RtEesbtz6257FqkfySBDhJEC3QaFzCnL7MzHOyYTpIr6SSy4ICSrUo
IvsYqNxcDyahcELjXCKP87fF6raAWOh5xkggpvG+CyIp07YkFEDPHG/802MROlky
WyU4+BGYDk/tVnU/owvKfUHBNLVAxnHF1rm+FYcA/C3DklwkFq2/DXl19DPe6prv
TWG0IpHPwmXYIQQT40qy8Z0u3RuR+IJ8o39YxSzByJl2xazhgGqsbQ1a7sT5yAot
LSPuleHzfQRn8PhXXgNTiFc8bU45uZPpwpTJrwvBXPGuiL72WJUye4zTYJlXGVww
7pD5M5i4B3MAvhQuD3zFWztyiSPm3Im77eIdYmrRq3vD8evqyX8nAj75o81Qibhg
aSx8v3O5u8kQIYgos9a+nHZoNilRuBdMsaaFfbIyAs7QSdsuhdXKnP4zLobU4QAk
aerDbhc0fg11C8BGOCpMpTX/Xuu/mXBPjfUl0iQhBCqqmN5UVoT/FPO8IaEZJYTr
jb8O3gqSSwfIGWFFCmd6ras4No77JAvlmO3piCU9Gpg7yas6A1V86MCVcu3SR5UZ
ueAFAArSCzBQinZT3btj/WoWVY/43zvXdUwrC2W67Eu/Q5eMqHslhRkBPDAZ4rX4
40jbSGfkVIc/WjshXjX+9RLFIH41yCciLfXsu5rK6gNG7cioAQGNLi/N52iTYU3F
ZTCBHNMiore8mBfW/T90B8fAOMmQJkJ0VFMaMEFrozqRbm4VNX5/qQADnrVBKsXs
CcxUsZAkudng1k1wV+jjn5cUoME4kl8qJXwoQE5LCaulkcWAN+ItnSgtZaBCyFZJ
+RlkAYLMx0GtAQgFDGQJclPE5rgDWAutpwPTXdUe+hbMKSdd89EABos1COExhP+2
5RxtbtwQsAFI4YULHjdIWIC43lFQSlQjhdcgD3ttoB/2aSRELCbI1NcoYebfubTW
IPnti+l4E6lhf0bVQJpQQ9rZdC/FafKzqfEdLnpPhRuApyzqdl6ypRXd4mscg8H2
YFCrkg5ewr+lL+5yqFXTJQWa5d5Vp8mYo2MenbCgiGr+yU7IlI2mXv+qkvcooswE
C84rWgC9vGNutNvAXT0lpNHgf2JO2Pw9C8wcEXb2c5zYAqpAmPcdmPx7ksuonArh
fTnr02daJ/HJgK0/b+Z3ppufRA18wCs4IXf6vzQPySi58SY9qrOEEMEdqO3r/CIJ
5M8tcId5+0ypQHZfWVuWGQt6kiI7HhUQ1s4TIVijMo/OtJRXKfrOw4nKr2CeoO4c
jt8fRLEsBk+uVvq8YSQ505K6K80BUkNiLooLVoMHC5aG2VOmJt1eRJ8Q+VqvYo3x
etQdWVK5kYgcbAsjAqaow0VL/l8I7lmJx8wLgg7BHFNi26HNh5eKlKZjX5fTJeTZ
IZOKMFs5YL/szduqqFPXWSuqvpDpnUEGutNd23eoeEye2FhNaL/b3qgHgzvVYseU
GqBXqwFCI+XSoE9uzvzMHAc/Wx0ZaZb3F6K4DvcVmTjLfcrXuZ0SSqzX1vXyKQB4
PoFOyZw5UMkaOIf9jVFt6Zlbqh2b3GTdxKa7574prs1hfpwheulwKRk7HsaBEts2
2g17UW9h6+rghhmIGXoy0JQbRrZp099cj01MWX5glkJYj6qbtevppCiNKMMP7AcA
PFckrZhizcC5tcNXh6kD7EF8ZAFU3ExJ0sxE8VSVJ1nTvdMkRkIOzl+6VXvivx0Q
z3MOvjjw7J8qahMbULy/y6GPK1EdEqx8YZ2kwjYhlvikXJoCMDQbOQhKWJ8WOJwB
bsoiGdzwF8rg34nDW5Oigra71+Kl41YEDpwSeulzyCMx6z/entDT3Vmum9ZLG7Kp
kTRMfWXlJE44XMQ+8MgxUjCo5rS+uNHxflWaa27SsWs7XA2Rn3ZY8ShjQ1uAbWan
8+5CjQ24jgkojVIlz4Oj4U7PFTAlgBjMrZcIjPZGuEvHC0VgxTQwVMxEK7Tzlcth
4zXQHNIdv/sSAKWWyTT1fTcVvjLcWm6ZaB870LSPXhErLtCAvEmDSo6T7/SNpk40
GJQWNmCXr76kBNWorWYUxZ57GjwJ9prln7pzTuHAWOLDw6TC2MS0/VPPpnJjTmEZ
HsOA7riH6Nl3HneaxKzdQMVu48NR0V/urRYt3Naqa8xx7Q7LSlOrjoVGxLKdU1pF
6gBiHXc8QrRZ3+OHuUzMes3foOHHP7Dj17X87UOp7uK53AfcYhu6WtJWu5lCkBQe
T7sTcaLefup1N5NoDqObvaNWhFI97X4U2Xn/mohQ1LNKrfLeXyL18YDsnvtjaEQK
rfYm8Y2FfhW1Lbf9unacZIGqs0z0SiEHLe17XxG1dd0lR5J9yyk7IkG9GZmUyrT1
ZbOB9ZORWV6BMPArKF2eGIebfbJuP7MOLOgdiEFT6YzeeW0I82iUu8X5NZibGyoO
cS6y8ysee7ppieqUtQcCkCmDiQpVnV327Q2VDz/k7ZYAPAXfDwCPINO64PWdUE+6
PQ+RtXMcleQWfv408dGAyqRRCqRtGu7vFPsYls6k2QdlLkI/V51+5Y3guoB0F0qQ
UmvccBeCFvuRnDfgBF48tU4V+bRoSXaGALRrvlyz8tH68mRnMpMpyM5aFqGnLxi9
9QbSIENje/GYjDVhpJOegQVp/ednKXueRpAyp0cznO/fQfbM+ZsHz7mh7yh4zXiW
VsOzVQi5ic1zv0gOZKpNlX0y1TJcvxIC1zS3pHQqky2FvccW6H8S/EvKne/Qd0FA
cw1D8FYdoaVH9XO3WPgzztj3eVe0IUwpotAB+DV8BxGbI8XseokkiKH7ILXp0OYP
WbsTLM/Z1zozsxcwpr3MrrO0huvfxjHMjCnO1VhzkZdg77lsSMvo6DZccxidvnmd
S3JPA/VVpMMgdtJv0bXCg58zBl0A5SThWVRcWr4YNFMh3zeAPyjCwuriS3VEgchC
q3r+rCRKQpk3dj3b0S4hdHyzG1wkiuaBzQmxIl8KvaRG+ybkufw88kqophWSQPrJ
vWatHYRawtgErv5psf0VZCGyFIJI7RIaLZV4Z9tyVEvYHB8vYPDyNJP+cr19vWrq
Egvx3n0449H+xyWb8WtU+kg8b8ulQJm0XgP+v8LBxdsSLqGGwZASAB/3+mBIQDAj
IqwV3Kl6+tm6GNIBT2TwnWS3qopdIA5D91t1WXu0suclm9h7uA/9suA5/lBaeitI
riAZhCOE0PtFORIqy09ACaQbVc1VEk9lY7mZwvziwzveiXalPs8m+1C2/sGo+H7s
xRHOD8H5OgPpRFnye04iIeam/anyn3l7EwxIi8ZUGX4Aj3SGPUqdA9frjT8kcpwM
IuD9CVG7m0Xigts7ytvzYp4f7D7HIR5t2o6Trxt7wKmb966TQKlkYM+fai7ZHa5o
56wgmn4Nd5DLe9XHyZuYXJQ3SurUDLhUavFKoFQQ+wLcOGCRh76VSmuKNbpb3+3n
zbIwKjuwseckrKmMm0fWrnob5zo7ro+WXiFlALUh9wmGq4jrtR7JrzgV6tFVCzUg
WuonHPXgCwCqw1FugRIaeJDzg1q8/T5dLiAqt2fO9HQAo9pjBvZBMCo90ThYmeFO
U82pnHzMa4jtv0hIIASwCw2kxTh+5+PrqlgzLHjE0x16gL8YmQJAhD+hmSYRhJFg
6hrRqiInKj5CSa7z7Q6/CR0/iuAJeoK7l4RNyA6wRuIdYDdiGtQrWv4/bZI+1bLk
1YE9iTPFtxO4+aSLGr/tHQjN/jWjjMGTOFwg/OMVDISSWFaKlgCMTHBne1PA6zNs
Urbkl05NAdcIqmhJB9i31qTLN1Fdl6qlUk8C4XkSCYnaUIXDOzVjOcvHJ7jlCGKb
ZwkNpD5ZikeFjTwpylYa8P38dCIZNOPPU9PzOtMHlZGEoqYLNErSR56/4rdutRNp
dDKgOfuff3km9CFNJhMnr93QAoBZQ45pIccGm2j7i0/JqXUvpPC7VoMSRCiYNB3x
UxNiB8SrZ6Jkb/vpJXK19aNcpb5hv+k7v5f71gBlr96HE2v49T9+At9/42pIu/gI
+j6Bf7F/m9f7/2Plm1CKfP74dV/5mkSm+Jl7oxaGg+zE/sOxNbMjPRCWipu5SzNe
s3MD+iV0TQDH97gRVcrRrdnPwsY5xw7qF/VGl33JguPwEkbclNU01axFKbzLVjwF
uHmd+BU4YcmrXqWFGTw6EAPljUM9S+JYMgPAmqgFQJhbTOSXB/Uz9qBlxo9XkbgG
QWaCpliV1ukmxpxpOKf3tj5ibt1dpaPUVeqQCCOnaiRyMg0asWfiIUCjF4AdkndW
OAzDvs4PKhxgd0avxLvp847pg0ikd0EZbHYktb59Ds/Px8Qvt1fknYM1RiejEhXG
fmBGtTeXhj65NtQddVGM8vQY5bcCDDwI8fhw752hzvGuf805wP97egxv/QKW3DxF
tbmPSIPDwut0jckhUVQPi/mJN3wAkqyPE+MqYuxMTrki+ei/bSe+3OXEVg23ClOk
8k3M4135+AZLzS5NzM7m39/P4AQlXdkXDYbS2SfBJb86B3hyMR4nftQFSdPK+Uvo
ON593qvvaTxGf1X7YpF++wSYKnzQE822qTWHrgsKR6AkCoNtCp8/LqxU+NqQJ3FB
/FNLDIDvK+01BhX2cT496Rx/oJJsRU/8Nr3Vn281IeJHXXJIsIfH87BQfI6SClex
/6H7wn/SUFuQgTRRlcOCjgSHaITD/8RiUVtBUzvOKjoPcFD5F1K/mC2axE+ObVgo
J5RVyflmJdMpwAZrtYWxUM4a19EPgpmCqng3/mRTK/LUvY+iVtw7veBebcgZATd0
nbVUurUWh2yR2s8H475AYAM66bIU+AEllGaCBG+u8L2nE5vDOrxJraYPV2+5Kaeb
XqNayvdl3sn3dUXS6DoDvOMeQ+Z+oYTBV5qK+JTzAYjyCFUXd+kwmfu7ifYxFv/j
qJSl28Ok2BGpEg+VcG8dnpBUVGVE5547xnqxQ+flvJ7AavwOfngJZP+dADx7VaTd
06vWMng/urhrdhblBASrAMGeEXY+E86ErwAu7TI5344YirYsp6KuH21gAn/r2Ppe
sj9yMH/D7nIvWU1ML/vBx/dhf6EJ7WWy/j/TVzjSQq2W4nfdC7Vv0ycSm5n8Rx/2
T74u17eqwAfG3s3SY/iJPl3jXkwRSX8MrqlzgzP/lLqoO80JmxAgVVKkRtuuOECk
35adEymGyv91CDo5hM8ZwlyK7D9MFN4Wdkg0LefGnwslL6Ejh2a9K19oF3sxk30e
OgSMC6EcJYYaxEZ2MZETKAmrzvsnUQHFKiZCB45I7fXv2fNF2HbM2MGs6ij/bGQE
N9uzXJbQEgn1N1wwLLz+T/aiFQjC/wBRyLvck1AgxFq/dpsuA0yITrpV5kMsV5iG
EANQCBrOl+xDOvOfdPyuWP3jDE673K564x8zKpIh26JOwFJ78+6W0er85U7xZ0bj
THRxwC1WJ9Qk58mDZmhISffQXm+PR4yRGBgTinNHX19wKH/GlV2pYMGWGeGcVvK2
/kuffBgE4dGVHYs8pawbSGP3CxwKdAGJ/Rq/xSxYMraesX2uJw51QjdMd5TiLEQI
ew2PV6fRJOdf/7+zclq9CJbnmMtycYxLbQNZFNCXg34mBiNzxMZDVyo4PewMuSdu
4mkpKoNKsHlg4+l4w5V376dQ9cvdN3TVw++UOdPYykSCRoLnKRyCmzSdcowbQWEm
3cH5CCpYBF496OXWujtceZFtI/idaEjUnPoT2ZxYY8irQrJvCSj5+pJdMD03Ft32
AnXDRVbxtaopko3FRQh4xNpxCjbRYARSKgVwwJ1wBaVN6PxNv3Yx2r/d/1FirGez
/+mnfvaMpdvlrtGyA1Xo9q6cGwUbp1FO8Lw5X/nrYqz3LohkFmN9W4us7J/mtwOr
tD9Ak08dPWLFEeY2015H360l4M7sVdPXYcB4C8XXGC473J10swOACXUjzMeSbUQM
KDtAlYnU7TLppB/aHbSVe4HT15dwAaNHVObT+WAIo6aWg3zBLz2SR7L6iCXZD76O
HBTo7B2/YcfRK7QTaq7BiNvbUCDuwpwdlJfjgXAOoe50CeAjVCCFMHpFII3n2+C7
hy/aOEWfRMIxFpq/CwRRGg5wVawXiofHfL3U/yqkEB5HdA/tA1atetB4cistYcPr
R0tUSY6J8cYivPU5aQZ70xsZ1/k1kHAAGnsacG9MUm5/nxXkGfa1lc55tv2Zhb4I
KQVuhGi04B+mgm7DzWyijz2AM9eFFtO4Ts0pqd0S3EzMPiE4LF8MQYWjgpIWEAyc
SzZ3s9qnYD3o4WtuQOmbBBljNixWIAer3DnqiFxZBFndFIPQBGPDfQnq+Ew6Tjbg
tw5ZYNqTD13kxXH+dpOqqbodNqlsVPO+o/yk0MXoP4Y7TFifXr2KYZUOAy+N222s
ZPMKzjaAbOqB0ZekC7kq6cZcrn/tUcdartOaDRpg8gLCnJk6dQPmLaLLNBPFyuRW
bvuRqpPJ1GC0HBWiC+XrZ9+jpMDm3bT8L/tq1EdE5jduVbwPQ82we/8dw9s333Q2
TidAdOyUf6WGnccOnlQceFpl3YI9bd+91qR+ScouZEn+UqDa7ByP8jZlklyU6f9E
E6n6hDfVHdKN70oR6OAuDEuqiK9ALU1D25oeFXY9Cjl/sEhybnN6jayBJbh3DV88
KimePwDXmHAJxVh7Ol6TXRhKWJLOuNnM9w6JiI8cOcSt/Bw+2G/Eet0sLGq9lnQt
MghSeUW147HG7BqbT5gN5W1wWmM1ahsmolJlMXYIkgdLhVgfO7XJX8JyB7BVvWJ0
NCxwtb9qSfqg2nOkqNSex7Z72EXPTsJbP5Us3judd5oe/NArk47fkIC4zJl+0dao
xaz5G+EzoLFGtpUC+5lT4sU8oU8DRa+jTu5VJ4nDKz6jzzNb8cw939KBRIjZ+nWd
ORYHmn9xd5+OLD5N23ZUxSJTS7pKDxZIKYxHP0kDLF+TuxghrduXvcDtcTmXqEqX
8IfA4b6YUi6RH+Z0It71Law/sF3IkMGmdMvnNMKEqTfQuTxqixsmFgkGgEj1OyZ5
zUKFoKnQoWLlIisSvtiy3rVQKx1PeW6wG8N102VoXBPjHz4jwvZn7WHwybxD3zeW
x4tcaYrhvyz5gPKZoCSSjaXUS02YxheyUDjrkU3eWaKn/FJ/4Tv0b71zMSz+NYgt
odfMnSRUs/SpJV0vlTJL2N6lzVwMcu515JOJs7p+W2Iv6oX6C76OLNri8P9PvnGL
0w5CHsVf3wHOG8DVRfQ5JycNNUi+02GAye3Uvx7QuAQ9PGQADjBbfdmugMJ1bLzn
nvqkgkWcf2lwE9/K1iYxR0i5suU1dMGcoTv28PuIn4NJodZZvgy+cZWUlaY4oiRP
UWzI1fIv1QjL7/VIRIvhyVwWqGyecTXktcTZ+QNU6/C5djc8jcgG1jCIMJv73r2v
zGIUcjH49wqrvbBmeb8B4D4XFldSIDM36oiGxZXZ69xZtXChdz90jcAh2+gnQxbd
5YQbdhpbrpiGbpyW7ywtEvFQkqrnKMrCRxD5oUZfU1euxXV68g47oLp8NiWU/AuE
NLT36h6NwRSBulLSmmbtw7B4IxuPeOB2DtrT6VCgVd8tCICcIcdugZEPDp1F8kUd
Xb9htKVEUK0kVJZcBnpku0xNDoho1vij+Lnvq7b23hccvH5mnLCWfYuScXa7wL3/
auCGbi8SfnpXcjD4Ggh9V3tEIO6MDoxwk0ihtPtbHe6qi9fzjSDKQ32QyIWkN5M5
sAhpzZrg8mdqnQZGq+CuQ+V1XxHsoPoxwragCrzQ7I6Ql6NJsDIHqo6x4AQz5BVa
9T741R5G0RkM7MaBnS7c3Ie1jxvDh5PJMkta0VYTXsEmT96PPEco07rn/pPWG83c
WbITzlb8hDJvjB1zmV42R+neR0sJ35e1j0Hu535flQAi1+Bmf1pyUp8O8Cq2riNU
lP72sbge9kaCDzwdv4IbBfSjts7McKFBvKEWsbVEVdhiz/Hg1UtFydvZuf6mdtKU
cxX9WcBG4bC9LC/X+1JEpY7AgoLelhv2RkHf5b5vjED3qBqTKw/F55/WVzSgGxoo
v+xpYk0czeQPQUdrtvSqGuwRT5mUvBuo5q03l7zwIHxuBmnvMmKj6ULN3grWAHd6
qtACOd9iadq+EGZNqXwvuRmBhjKiaWrhI5//fDt3g/dfjb5KEdR+mvn/fkDWxwPZ
Cy+NyANNUGLpDT67Rgf4Sn37wYRO9ypBUclP7cxUBucylkZfz75VzpU9+YoMfq4X
tIVFhl8ljvjHq1b8Z8mOaeAxrzrNARUdn3Bgrr46Ei0Vl1qOa1yHyd3qfsVKApxB
3e/uhgCefFgEwL7EVqTY2kiu0jJIsuUvLFFGCOY6pWA7TeKT40JB5dmPdBuanF24
cZ+3UaSeRgakdvmf4x4jH+0G2edL15B+7YGyNABrBFQoBNu7n1BjndwDDEgEZqM4
gqQ1b/XAuYn+Efi3Wu8EXHWWA1OIjVnRbnaetcjZQk3nmAXTha8egkrEeYL6kfIw
rMOY77BmVmtpjUX3YAfupatxSYUu3m4TJ5JitvOLA2WrZ1Ng/ckPUhtUFt2NzJ+v
K74fJeSIHvABjwp/T1knQUF4HCnYJdLiB0EVVNMMzd4TE0Z/CvwX0AtLKl3X/NDt
rWG0NEZC4brCue23vSrAfd7+DEqvtwHNyF0AmZu/tX9ZmEBfhqbXzsCoOGDE4d6K
w6fckBY9gZMKdzbG6+HV2NdQBRXxnWa+JvZpimGEr5DG8iOF+tw1wBEUf9mKTlPi
fqp0OdnQZT2sq57v65TKgtKIlMaCmEDJCF+7p4QNjcGQT9cCATThA5S2Ppg1EfQw
c8LLrllGL8Hx15nIwlua3NIeQIiccBLTOv4UjEndJXZnXjirEKOYTZu62uiQo5iM
zV0dAUhfKP5gDGuwXpifIoDQ36kE9q5SRuH6U74aVRpnd1FT5BkJlPlvCyDi0YFW
Cu0rWD7oTw2aaWsoSsmCH8L/SMvdD/NmZvD+l88uXORMuocFPEJ0R3UCz+hzhasz
cAM4tGi937Ex5cR7coxmg81ibkmAS85cG1R6vvsSCFlRHFlnaN0UB3qPUFWJs2vR
03FhvlNyZNhFTJU69wtLF8D8o1xH1PPe68k88T3HtdUh04WtYN4fCbZ3gZjrN64Y
ljfT4pJTvvLN/jCWQoxgS/esCCrTvdaFgA53BwdCVMQ7qz4aW40+NCafqX+A3VS0
1RFCllUgf/6r9C5gZHJwE4JsMnNr+GkPRA72cUnNr5/7HlvI/OuEdtjBb3GsbVY4
McfCp0bBwW6JdW1H/MDK7QIdCl5sPvETNHLhSajlU6gIuTCr4CMjY2UmL4Dm8VVA
pjcUwwcIg9ETXHLnoPP5uY/oESCRRzof/+js1I0Xn2k7hYkr6mrgxheXCateZZ0P
7TEddoYLeSJprynmcp03oOazMaPw5whQ3UV+sEfIbacDnHEDf9ffp8Sr97ap/Nv+
WevgoeoDcDu5kw2GDZ0UgzQ4xRpdv0HK/ArlR0Cw6Ld9mjyDyXsPEze8zlmF4A3w
zu9rAh9PWyFeE+9sUloNHejQjnrCg3LD3h67+RI2TfxSC54ayAjm2zEykWyIRtYy
jGvAlAMshvPnGszqRRyNesy9LCfy+cXydo7OLipoQu+TPMHjBgUg9otwL9rgAzYn
o78bSS2hP9q/jyonMIXPGc+V66R1kXqKXP6WFQ09M2paQXmUDEdUCrYR5Z9qt1CA
1jXeS9FHfI0CmpgYHZvbKxobYv2NrSZTucPcI6hAdMUT/0pBq9j+S2fjO66eSlqs
UiEJAr5Dcixwqfhudj44CdLMzlqJ+hlBuwm8VQn3ee+aM1ew6GNdfyM4TdHxl5j7
KNKDZIaHF5ryzcAxCfXu2dL7qGal0d9onAXWeNhUVP3ZqY2jRQ5w9Q3qjqWkp49C
txcom2NiGxeZOCIJQk8mTZRTH/1A2VPNWAvd8ErME7GEFWchdVJaiZK7Xk36hepN
yJwY26KjH63G2PFLmAb90fsdKaQ6YJt2ssiza4pJapvXXTN9p1v+ePJEJV8PNHNm
cbUFdF0yXGIPUHOo0nRvAZxJ5TJ3Eoj3vRVs+MrTOr7F2jBn+awpiC+98vPT59iD
R9XgllriUfpckwgUtz4gIGp6aZvaidZHzqv5UaBF2U9TVp6eCf0K4nxnKISJHzrk
JWcBDNdQKOyQXwGMcLHFGV4TKLBCJCkxbX/wi6eOQTWPr0UNYZQXTvD/L50Irs8u
V6m7Ds15n47pzGvlgvmRGB6XiOEONos3RKrrsrT7fvU2cDvAcS6yc4YsaRclGfKB
wCsiRXjReHDlTfP3PER1GJWdocdHINjOd4+k+0EOCmf8fcwXq08petlnrSbP/wd+
VK4cWYSSMNcKN7mFCE88kbEyJeLF3n7CJRHVKltDoHhuR9wu82vilBmtDDBlIzaV
tTWAduo46lKUYIqZ1GpYofraoupTo5fWE+WPKQAuF9dmtFwgaBYMuXwUvCj/4ad7
+c+zl33KYNjxkUf16MKMSDnfiGmbp2pLN3afF44OOzAlwITbjQ1kSbeAI8uitng3
1q41L5JOF1eCq4ofTf2q60DdlchBWYJIBP/JWCgaAiBAD5WJJLnDspRi9VVBBFDq
xBToThK2m8QRrS4Xz311Z2V3kX0QM2b61FCJi/fKLrGnCeKuPSUAxZGKHR5/4aB7
/twZex4gKUvVsp3EVLXGj/DWdyCYALVdqmEe7eoRQUikCJZ7NFAMYOjxVTl7nfXz
s9XjHOAPBPqIek0JNxXxkwb+IjtlwmfFQWWkoVU40ln79qkjv6UYSy2Oa1dK7pKT
t6ZeLUZMXUuwqQeNSQrjIFBRQK16CseOGu6YN5fafRIQs9on87TSxh6YqZP31iwn
D/Xd3DWqZwfJYeOBRCE/g6hnRQVmEEhpM9MKBo7bnTihCou5rcGlFIhFA1AH2x79
gRpBYfrDSeOo/VuHhfkPRz0mjgfCLxmdnDIJ6qM5OOU6l/5SGlbOlH5ZwxFQhDu/
wGnoM/f6Y/v0K6mZgYWBPqmkHQNZdMAG0nF+WHql25A/2G0q68p5dRX6K1F1cUjY
wbMEhea9h+4AWpi4TuE3uw3rA1+8Yo+aoWKzYNjYcKfIK70UzVN1ip4XegHOvtm4
SDJ3rMn9C1bbSv/3XmhrWh7+quPnHQVCugCdCLkmBdObNxcEDJQosjdCFWcMviIw
lnlp40RC0KFi0Lq3aYjGgHK9H444AmvSVdWer2Bizo43vQTqBm4ZQav1UW0vov5W
iqEPtXAA2JGdOJm9vhq82N7hqtChHApIaXSFbjU3Pl8TZ3jRc13rtlpsp1XQcBXo
Taw/PgVrvKAgbXAEg6R37GCq7iFIGibd9OTPQoizaV5zsIs4eP+7GNoruL5Km+EV
iMao49J8lEzkw5lcbHGbLMX2AMjIKZrImCfz1sRUw1DD9cBO1GCpwRZOFVz/PeK1
LbfYI8bZX9iwVNl1JdwzIkTAx13y2dYow0tEYruZ6d3MYWUgZ256XASn4MWBNrOj
VKl0L01bBVGKO2BtZ2Kwgh/dZjs6xE+/SUXHTjbRk6LolXcrqrxwj1SdOhOEDPNO
YE8EKutG6t+6ksqRMcoziyTlPyxMRy038bz+yXi0g8RMxeCcDzh6mBP+BNvUvOBW
JkjnGktgQ/Snmuy64W1QVuoP7hflJ8egCKkTl4abkDa9/QAOrv/0lt2glzHEhAHZ
c9qH2MIkeMcqYsAccQ2CQIpPyLrvtB0jxDaM7I2g/mSqZpLiGxKMOY47tQkHYk4X
0PG3SiLPppoOdwml2yCX6vRDTOe1Qobmg/wifUBYBo9ikCCUWLSSYSBhukTyJZB/
eYDLOFjLQ7lCE+SE+jRuYMUkjyN2EDAA5Z5JtFflde0U+3rulPh+jUgmXOGjv2zc
6Y54ERLVwFVdKrCGE9d8F3MAC+u4asEoIJ8pn4a9qG+6J4/+AJ76/LPdgttnl2cR
keag4pObGWiUFHhXYTf1t8FXrfS7k/aH/G+5aBH3y3icxAuGtPuvfnZRgesbtUFu
Pan05QvSxb0KewrAQge57tLiwQQn96R/9xB26CEW5Rifs3GmuY67cRwQ2BpwV1Zb
F/aN5nyFK2G6ajL/yoGOfEgMg9LkUQbvBveMdS0SeuPbINWfTnhPVxDWFHLlxr/L
poFS7rwTkahWD8vH8lyVJ8FPbMlDqpXH5Z5d3pQoONH100Zil1PO26bCbybTg5mK
YPwvzSkYZLb0HY9lWtiZBlg7qqu7y6sILAISvJ0ItVKLHnijSMxKaH80tC1yKsYm
n8oQKi77VUx+M0t/ekXvpPLfd7aGnNW0yxLxVGJDhE7esZQiEi+18oSC9Y/q5W1+
MftpACLelhI6+VIPX715eMzJqB0YyXDPimRvaDLC9TgK+QPHHtT62YYdIGNkU3/k
Y3tyxvP8eqpWoOyx8F09ziOleddMsyG89kvPkqH7iqihvIJG2DkO1Vx8zcJ6yrmP
YmnT1RUIrp3NjSF/QTSLGz9fYj6N8seICLk5Jkb0+UPpO7ZJ5+wM0RCgcLnjhYfq
gisVr0b8g7+jvSLjlJRSCqUv0LIDu1pVTWA2Ae7dP2hdnlpxt+zaKpJRFKbh1368
Ua6siTKL/XFi91OCZOn4J2626XlDzhpo51qQzygGZVfGdUCZV58Qj60My/0mRgIq
Cm7dqBHMkWdb/azREUT5qLjI1+ZBR9nO0b1PD3lPknNM2k48/wa6ktUhP3eyWK8f
5Xhx8/zUuiqfUOMsiEB3ftKLfc4WWuzAjO8+DTxoT8Y3a4NUxBTyYDxriv8oZI48
6xPX6c0O/w0gzkTdezif7BhT/rGQXHiRVisnUZbze4tL7PoHOfupg8eZPelCMpXm
9BsZVAMEAGa+miW+lgs+yYdo/iemE6qUv1xisapdwhdjooifhYqu/P8dOr/FbGgi
iAlcZxvtASvSP1uI1ktoqZOchCYllpyvUetbSOHrSArRKacVP3aCH4fh9msSWLwL
D1QTn6OI4rS/qScEuhysfDFrU3yaRKElAtTI2a3aBkhImQpf3ouLLSvsB5gF6WMy
qgrWlQME3hjNGFLtgneF4llqtzf5rDqVYgjbvTkW6xaM5PEDn3IjtWelQyk3yek+
FQCLVvNC1CQeS9mbJ0Aot68WnSPU/ne5VrLM9/PfF6VGNApYCOuQ7Cb2Piz4zdWG
TR1JIv3zoymYfK7TIepSHOSYRgKoG29p70waAcepz+OhT/cVnSTbWCgx6fgwcH6B
vS0YN3+4EU421z5vUOlZKkdQog/2WsrtyFzvEyMX+viy3c4JQKzySFnGw5O0MuzR
9tEwVYgBA3IB996OCpxWHDi1eT2OvmP6yXDriJfHCqsKmhW+kq3JVndssFqmB2Sg
3xqLA9g+7avDuI8e0T8wbUNAsw6CqJf9u5famogXQkJH4lMeK4NVBlVr9JCiLKgs
NwJqJ7pkPUrui8eC8zKeZ0Ex08glRrOXGAOkqF6AL94/u7PGqUeHiLbbcUhg7rFr
mz0ZIDXNpwNG230VcfcQdV5L4Z+AKPWJzkehmMOC9TgT8DeU22vI2x1Fmh9MIU7c
wzXOfCtZjTHh/2G+JVQUDFJg1uULUI2+NEbmk0sjY42DM7r8421BQLNM1sVuMkzY
Hy8K6X4MWSxZb2jrZTwUXoYW1o7PCsFkf2ErtwyrOdrBFEqPonIz1zwx58PqsHEx
fvIkWvVnJZfDnAJ7nUnQN515XZXPFNTSJzLH89AvdDXv8aLa5ODyabHZuT9i/EVY
9cNsyohhs3PgUSBI482SiF3hucw2GSDUnn1hx7QM0rzHsMdWEQpCasChIZS6uyTW
rCxvt5mjpxriaw3CuwOqsHfwTANfNUSNinxC6J36553GvXQLP5KVwDj6w/oajt55
pzPjth/czXi1O/kCsMPZJUDgBp+d2Ka3d5Kuo/TkNnkNZw2wYBnbhe/q5kfd55J8
blPL7xmvp831rhOwtVs04tuwv3ToUes+qhF5zvqzHfa2zcQ65t1fjHVs1HEK5i8Y
BdiFNSFnqlePf2BQFjs+zWFzLTKMMNuf/+Wa5Dpe92vIbhYMQnVW8EAggWr4EeG+
0A/Emt2n+QDzHTMxt3L4ro/cBx4gzERn2eDfpCvZ6dP3iyXSij6W9/OIkVAthGHE
lMgDbNTxKIXp96ARj0UteoBvj8qWicfbRudqhIsr2AYEyRYuOP8r7lwmvoGYZeOW
HWZl7k0Hs7rwHbhgZzQBJFIJMiAR+GK/dNLJcwG7mmyBVU7bvAI0P9ru8XZYVumi
FKQbqwcMkP7/czzjOlQD88LMXqbtzqVyX64N2j3dQ5Jczuq9JmlaQKfx9FdHAf++
H4b42S+X3Gxnu/CL62Q8yEIOLXmw69Gno4z6BeYTOC/DyZfv7/qoZVp5B+vgcywD
XkA7RYACabwG943KUPdoIoU8FkVBzRi59hktSbi5B6r6oQ4exVLqqwCSLfwKzwBB
4H2dR5pYJj7YUjuyDsjC5onURuFW6SEMu4G1cHkVXTORSEbT0Th8NK8DN6MuRPZe
91SRYG8W5mmUKoxCy3tqvPY/cBhwoKINv2KJNosf2k6ZQk4RUyDcE9swM1D2bZfH
vGtxtl7tYc/usHigswHfVTpyVwFnAid5q6e5yXFQuKkX8XuaOZwLFM8J2o/7ZxYt
HWm/GQp0I7L6cOyAgyFiGpF7d3VieGljCB6veMDYlJNFFNDLSPDjQ0zTOBCk3GQA
+GJoygjSncEyEKYng7RDi794RfBgtHEiDDQXABuD8PMVFMvvDq86igrCKfhuDrUp
q2m7xhmQw8pakXzD2EQbUOMOJ/1ouiLpE6qpTCQC+TbW83kF/7y/vieEbsQOM411
NTsxl3wMzKUNDa+e/8GLEM1bu+ArT9btyXSSyFMzNuDvXz0PPjGTCZRpb3XCmtUz
9WqzHSk1E5MGfQM282kllhogQ09yqUGoyoOqtVjNI+sLMCG8k0GmSzUY4oow6NP8
H2xGLKa8EaoKg5YAacr8DnuhqBW7seKfgqbBCvNcCngaYJsreEruWbB3kQFVCkWX
IDIxhjjraVrAzqlOTyuvKG1tKySpUDJb1cNKR+Thq+IuBiSyslwjQcj9wBZVPyfp
HFk1VDclM9MgUgtQHIigQIVz5cFl3PAD6YqDifHD5BV9YHgoopxVdWpHGeINo8z1
aGGlzz8qNlgBiMwhlp8afch2dr5WmffLFVB2PO25BvQmCy3kXiIv0FidCBNwVxbz
tcSpb39AIroJJWvY4+KQeN8VPTX5ONfPAhCJNcoh/uMs+KKEXlSgKbpgu/iP60RW
VKdndsisQiVn0UL7WrUvpHEnN51uXQOHPdeK0Rz/d6lqYx5mchM3RU3xXp1a6PM9
DraIilqy+SgQ5mRrX2RpumTxL7X7az8/R128Ho9O3txamhaUbNOJXNv6KEcrXHlj
AHNoVZl1AtkYXnLDtQAbb4Iyme44rkRIZtOtVAFNevQXJXXt+tOLbwRttBneDwlC
qwiyvjUfwg0YXB20RRSJiFMSupwhG1ICCpD/hUgylUzUfqiULnPS3RV0xiuqHU7j
kAg4eL37pmyAIusT0JJm0255uL1LezSgYtLjezSaDpj1e0ARiT7iPCNHRCFRXKU8
rW2D5UthWyOwHFA3NWXFXqH+gPUFwvitGgXbdW6Ocakqjom0ghyPGh9MBHO0YyDz
AJgbrYcho898qQiHabWdbpfhhYq+AAsq0jeq8QpVocvIDTn+bqrnsQnblr/oVvaQ
rf44MnjK1EvORe/UXLM5cElvc9OZ/K/wE3nVd136gqI/8WybfyutMrdgxPdIg3LO
EWDlLoPteQ4ZoM86KFyXbRV3m0Q6io9H4ZqZtzXNo68LkhE6O8PG52uyY1sh+0dE
kz0KZwshgFymLGJmMkCFe8Gj26s96l1dr1/XmdkV8DjF/9+70QKxY49jaozK0NVh
03nx/JJxyzfyGMEVrc0IcElWHZsmAUrsThsu2p7Td5oqA3pN+TJW7DzgAgWXAi+P
TtN73uMrnC8Q/p1Gi5w++T9tznZBxJTGi7jG4s1opLb29LrhrRdjMqX7WeBjSgDl
erjSdHhhGnRX7cUp/4wJHCMIheON21zeGpxK0Jl783gcI2izpFvOh3OhTj3wK4cx
CZmiz4kEKxoHUndymgf4j2+zZEXINSlE3JHXZSmmr0OUUt23VQXPZeH78qEJEhce
mMtq8I/fG+Tyd+1J+FW6MpyCE0Qk2SNafZvRdeN42xR6aIrJvD5V4IpoDcI350rK
blBxClpsVbcNpO7mq4LFEjkVCfG/dwh8Ldw9I3QpktBjKHvvjhiM3PGK2TbzmEg8
j2Ki+gDq70QKlBvfF/gd11C9Tv+07H++tSU0rxWMa6vuXjR2/hBYAPyLO1D7fF3S
ymvIwA4hsDqiUDkzQ9xioUtLp4zD9XZG9KKEaM6UCu0trF6cRRXUDHh58TXVLVJ/
9egXQmbpsGZCU52wZ6A/bTy/rK1Ns0q2ABZSCwcBFuEAMiLdqTBzYZqTTO4F6ZFy
1ufpNW4l0jeI/Menqmv+QOm3Nly+yHH2+eUMhAbLnO9QSeibcqLNGa0Cfy4tx6uX
2XFk97qwsTxin4Kdkv/8W4e+qYHpkNMZIQkWMBBVHi5PtEV6XMPhTHkJuTn7wy4A
jYvSPq7chsXkRGrOKoEDNx+qgJAtMHAvuurt793bHNCDNLsaaoPQny9/CL7o5e6T
GDKtox04qLtvezmxnvznuHsyMdiNOLYGQ9VJdMC6FPJDvHHGD0FNIySZZMiMDjin
nX0py9wayXa46WZ03VBtvE3IHzTRtTFeMl/TY7EOrcJygtgZQxFWB46Q+EfeK4cO
dnzq+66BP5M6IIaW78a11JFovHDqtbV6Gkxy6Xn1jPSPC9pYEChsmoafiHPhmIDa
WyD8L1iQLVZRRJUQXWY5VLAGCWpA0c9VGPXtvZH9JS29o53mKz6LkwRzphnCHu+E
E0EQWrzTxp+HSrKk90NTHTt2FoN7ZV3JqvRee39KafhK4W/oRLjC7cgOIA7Rt0BL
tWv4KIaxmxjwWMfjV5JJxz5+hYht7VC5REg7q6VOWWlpVn+zwScZoWsrIp5hCMyx
EVMxqghFtSe7TiTs2QBpCDFPb/uywi7iDtLwBhf65rX5ybudSIlpQQ15WP9Ylg6P
FD/Grb5gKkxB9NxsAcd5HMwQvCgJknHx0NZf+uWcBov9Cu/v8yDufd+xhLt1p5xa
ANHea0SOf2JKk9dQn5E6+jCDmK9ZZAQGcAv3s0yLaNcRCRiF2pFm6iVV9ly1bH4L
dJXP+9nE4C4K59LriLWV/UpE4I7pYuXxf4DvlsCekaTeb1wToWYx3khql9/cS3i4
8qgfpWD5Olsrv7FqPTB+ovjzdg2Tc9MgMKNZEPQ7e96GGaowoCVI3IPZlQTn8/c2
9QdmzHr01OKElP+5kwL/eGUFUUU6cfG2zIcldtCM8MtdgDirnycDaD19zTAb21Nh
1JdpTVTtopYdfub7eXQLdk8SOShARisajjtZtY4gRjb7KBxPggLKRMpbNZiAFbmd
wgSDw8HDY8JsQZ3Y7cGXeDxflGEHWxoDIoiiax+SzhrWt1O4RYMscQL/sb4P6hFh
D6dL2aGR056S5rtnEfWaOa3fV4u7E30RXV1u9QQQhZR7CaP0umCYLx+8QPr96zLE
LAa9YDd+5ohipowZp2h6lt9nsFFUYqxS+PgEWsZJZZu1jZdXQ3NtM6jbC7VN0uHL
0jq3wK4aCjpQ69XedO18eDWx40XyOV/s8inx5UdhF4mNHz1JmVHPXxBggrrAOmqy
4PsY3L5ljW6q57L7lUTNnuuJR4bCe8CzcJCELbB8Ezw51WNH9N8iDi5BpL42Xcwm
XCxilbQL/r+jl/nN6f+7nIO47nxlzUVENWZ2TRqpn8hjFPlb0h/tKGPdpcqiQug5
h9rRRuNPqiLlM4mSal5xddaL/KMeT/2w0xUxV2eqWubjYF1R4phr160TPipSGtMi
CcP5Oez5yVKn6MxhA7B50jAuo6z62A9bX1gmxSemhiBXpddocolbfDTkYzkqtbnd
1NaoTn5zA1ofFeB87Hq4/b1UM9igN6bqAo6YP0GWOhjzBn0o5MmKfcOkNN/+P5FL
mmXQ17pMrGDTj2p7UN/yLWmkPg7uwpDeAlPW/OuXkSro7mn+daLE4Jvzwl4ePNgW
JpNyIhbzOMyIYMKLAGiFY2qjVY3oX4dJxcobNt0OBOpSK6iQLpavr4ywrPFx2Rsn
gCUM3uAhd6WtnLz/BOCNl6WJOy66m4Lj8HvRrBpSbYFnSzzzev0GSwksnhkUSIje
CSQjq5MVdo6GDDUc3KnA4NXNcZc88UZhPE9j6Nu3kKMHJKNQVtxrYfUWzIlsTwQA
UlptkvqUtEJrsfFK9B7k1StZ3wbNffiPfXbMEwgAgezZkICkn+em8eOoORbpLa7I
H5n6gngiJaIqTlVMGHHgSzdJtXn5ypnr6icgDU35srMelqMfUr0kZvqdtLRY2ope
HmJEQRpNebR1OAc6V4GaFLWDle0Ko5sNMNEuk6RpP+JIO77EfYcm0PPaPcMjnAao
irPVZZ/O9NOth+78e8MCsjfFg5Xp6iVEqDvznWJ6XJ5Jaq0uZPA4KrWKk8wqCGfr
3iPhijJndMdsfDaDWSMac5XbcS2sukDUNjuGjb1gBXhhzBmShQJxx0thpX+/EPRN
Z6cCGpE0GqTUQC5gt6waPZpyO8QHEpXQ8B/+C5pa4FBDxA7S8UEl93/DeUUy/Wg8
2itTxSjpienobOjl5S2gJcsFICzSREdDClVOZWgUXRcMAniI0iHdMFtIDfIkqiF9
H3e2BgV6wy+CDcQzdAUYC4+zK1jXbbvL5YG4B9LpM3O3qn7AlE/UzyB1AuNe4VcJ
YUJi8yxD7b3KP7YaMw4TlLzZ0sMbIjaB79ZDJMXtc4IHYKB+P2nuCHpiC2Homvgk
uuJueuEeA6b5ZzLkP7OyUSnDvCtBHlWfY25ML5T1FptSm7f0SG9OV6WJuH6qqf0s
W3xXxPQdj9Hd6hjLGS+HeRWxYw8xQGwqSn9shYb5uHQGYGvKhXof85ZFVoXLURhs
tv1k8BO9fjSMz1swcYpJUKLuVnQTh+7uHMQtwnVdBOg7QOdOD7+eStdh2HpEQSfw
BVNqTtFHcYSTZ4nmK5Ecc/skrv3J2Sh/pe2WWplpf9uhYJ49/qoZI+Lw78G2s9GV
auklXT/Yli+b4BuRQyD6qH71Dqt/ZqSDxQYyZ05ySPuCTJPHhGrI8V0Rt70GRqjt
vwHY/VW9dXaEZh5KUcXt4btbOULR2LJD7gSdzmQdF65Tm1lksf3sfFqWS/pWa0l4
PG/QgIsTicFZtKdHRIxih7qKLvj4FFZZbSidfwlsF0MIN/M8t0r4NoJgneKZjsT9
AkUSsQZGsVmh+Lklz3p6RSm9ue8Oc7Px4v61E2iiO88vzY5WsYrv0tT+arsc5Wzy
4OcU8T6cbfdMJXoM8lzjRALPdn3cqYBRVYFAerp+hGKSSYVo0PGDF2rde71OSiic
JVRgDETOnmV7FVWLZuE3PMZ/etGiV9kvuduQ4W5GPhwqrdW0chi2Na85U0/fNOYN
bWVwPxC4uRYJOazJlq10x30j7EfIdYnyErO01kMCtWtszkgmqAAo3wSGQR+fcTHC
emSarfnz6ga7CTxUh/7MT6HCusolBa92ztCc0oSihTKpUB3l0acoxwW1B5ZTcnbD
6oC/ACqIBiCOC1mYlBbXquo9xkIPC58g2A33dV0PTtxi5TCn6KejTbYh8fc6QJQ9
+XpslqcgsF8MZTjsum1/d0LvRFkhBBl1k3h9QWvXMNE9O4MbqG8th2R28Rz2KG/K
WAQ4eylNXtWULKUmUzNG8fN8hI6Hq1O/i14FW+ZsLVQTZoFSDdJlLHSe+tsulv8c
X7T+dM/i1XcOkPq+6+qijVfBphH6CKKX4g1hidmvujIGN3EInp6hn9miu/usbQ+e
y0fMMqZ7Lj4bw9jFk4r4H6LOhL/30owc7YpkEd9lI+lexhVGBqIvkz9nk01DXPnY
MX0OXzI4vl3dMW7o6jv6AP2iPLyRrD0wCV1bAu3NrQL7czpMiWwuX6iF8VL+CXWZ
ldVpj/9HIrS5jG8NemYIpdU5ec4SfYf0F3/l8FQJFtQNeQlQxhr/BmZqzKb8B47Q
4VL5purF1r/Rta27BL2GOFTq57d5zWa9RYlMEYNi/LuuwSK5bo3sC1S+LeXzHx6u
KrRizpd0t6I9Q9pP6VOmRI0WyqQohjteG3cwMgRparctgvBLrFoGBJjk0M/56loa
tRoOYRAG4uekj67VJHnoeDyjCnVBuUAK36muVaPvwFtCMn16V1YABwjzSod8MIxV
BQ2wLS5KxJL7ridFPKl4gwYuZq/BEdCNy8WDmGlGpEeFoG4QjGCJh53Cqu6rrKNA
r60x02hLJJnBJr7kGpYNHoA45OHtUFKd+jsTvCog64d0oxZsAg94LWyvo+1pgF7/
XJZAhMt2v5ne4eDooQ+XGHu4miU2aPB4loUoKFfc6j0J600Iogg4ViED+6XKzW2o
bXUHc7OR1iz2pQfUE0OISFwyLbAOaQzWsez3uMsqr3sObp6f7qL3hjNrFSXzGn8+
gEB1IrgaDW2y2TQC0sKgeX80f0IfCGrLKxgl1+OzwRoKO4IEEcYFCWc3sV5JUKcl
kdQAFBGO6JGOk0pa99F0Ee5c9On+kth8Tk8OECnATT0WJl4SpA4dJdss2A4lL3UG
vVXxj1Wpc7AL8bTs2A7sPWbhoiLhEpG1sj9w/NvL/ni3M3KGnr5EqrHE4PHkViyj
ICsRFevLuBtZFXPORq2nRMNBSVUfxMy8MKp/oe8Hsv7gIUQv07fX7SZiwW56nK+w
7VmEzX2xfZ60i9YKiRrbjA7uO0ahDxlF4Bt4gpteHLxjMUCTPNnUghDVommlEOOs
aDJEqp4NEJeOCjmeMQK3RFwLNiz4tbwpvhFAPLYb6k+5BdQOq19Pzh+1JfEg6wIA
pYoTFjo7TJ8ZiW517oEcEhBjKzxX++X2Ga7lle6BhXnA+yddH/zPMKMFEj10Zulh
dNDdjup+xb/7p1a/Gk3kInvhC/jj3nm6gjviRSaOP0v60rkq01I2NjiQhwif2Z2k
W10e/vr1URhgemA9ATKuWgl2hKkWkdFkH+3vJ+MdtbW0EWMH/AH5ZCjLI7MiHNqH
7viMxz4wdAlOilcn09If/0usU8Bi4kaQagT6nK1ZlhSBO0DF02zbWc8sly7hZ9WB
BVAdl6UHuod8D4uXnOltdgzQWn2WoDk0bw1vu1YDqp8PmEJ6CxzBg/fE0xuOkYZj
3sHpedB39y3bQYx01VbXPQIZdJ5VSOhbBHXbtLWiEZBgLoA3l+yT9y19QYz/2Ejz
SMn+LZ7ZXp5hKH7YSJnTw+4wbd23q+jiK4MwXNrf2HzW9BZuXbb0BICjKf1ARtls
cvFxOq2WOr1F7egfo4AdleDBWqrieaH+kyrG3zke0CCRiDf16OQHY0rQn/TKh5AC
LDdXWYx0mg/2jnrie2lWpgOg2fHvVSQd/NIqUDO9vwoUV2j5E2Gyu1BGZnP3d/AH
4iamNqWbXcW1ccfrRXRXmc5D2B10xfjzd9RRotgrxrK0+6Mz5LIMT/8KUqdjS3gD
87fwomsn/cVU5cuyWB5yVkeNc31muricxfopikmxfawwwCTwNvQ0Rf9QR9vNIJ/p
hAJ+gca7+Nb31HWA2rbtWSwSnOF1kUICe2T6HWaAf3z+do696YN4FVm8HCvXtuAG
0xpCSduzy82hWyUr8CuPaMhUb53yFRDPn2ezHUvUaojreEJEKGEi51i2ctfvHCjx
f/NorVD5DVAplr48dWOxbQv+PnYTHWXbQCxDP3uoast2fV/MwjBUp71QB6WUB+Cj
LmF0RyQRf9FlCdwrqoJo/5Dj3ws2GFNcRSVSLfuRlpP6+69yVX2LqNVDLb5ld31+
el61+ELYW8Y7kBIEcQGmfynRlUl26jPbDHztboKkSQdB1sM4uO3FSZHzgmz8sV/v
qsKzYfYJCsL3wDnD5SyeyApFlofEiT57E2m0dOzd7k/woL+p1LmVnSwpG+QNceZy
bSeYYlOftwW04IgJlpj80UJL1y3B3EtFV/BKXw2L0D0MH498HNZYXvnvEN8mmhXN
mHD5jaQWWB5ZASUFpKcuuCkg4yhdJIZzBPMfOKqOOZwUYFEmskEk/HN/s9Goz8r3
N10vgxcFUI5b3ORka7O7oYhl3gD7vMTxUT/SVsNO8JeE4zyZVoD0FVZ+54aZG8/2
fEFEMZldM0yRoXjkIXrIuYtwNtBB+GXKi5QEEmWaRAz+2LB+agWutHVeWbgI3Hme
QbJ2Zo71LXnzeZuXFqg69W/MiciWngVjzos/7cRB1idt8UNKrFW4e7RuB+bXwPKL
iMmpqcBX6BjVci6VgpYSlfJjbDv1+woujeyIrdqeMyxUjwU/YJDxxcAo26M0E4qT
/Ca3NExBi1cNCUFlW5zaHZcXty8CAFf/w2XwBAy0t1aEYvf8rdLDY0isI/fhZV6p
vuuD8UvSWFTKWscSunV6FX4j1/8Hb+QBHI+Pr3TE5Ie5h0KuNGOi9Yz+f9iN2Egf
hQcosKCHXwg9IKMv2Pd+uABauCGj/kRdnBwsX1wRJl1KcwmhlE9C4kN+4XoC1NsK
4ovhErPitzB6nZ3kxU6DbGOGCQDzJsXMVwYwb9beVOZI+5x9jb7+1JS+TPpXrE+Y
dDk5OJWg8I4Bf6ZG3VhV0Hj0sDJcNuC9aTdXDuUx/id5aCfmA4a297kFtljVmoH6
lSC1/BNPY0PUbM4FBrVMwlGyOmpCAvn/POhPkDabZB2p8hMKt0yNoEQgRAMMW4/5
85Kv+x1TJxltyQv158rlkVPATSWCFQKLTxMtBrRNMjhODCaR+m1+XCYDtMND/wjV
vaLJa/q/4BpeQOMHDezGGiHRkfOMQn3082eHNCFGSAyhKJ5ARkADHJgstMToHWle
01QsK32DZTRL0syKqaVpUVdKRvZpuh8SFpEYTHRkgLLMTDpW1XDUfxkq5q7Lj5r/
ACpPoVRudVid42OYwMKNzJVNG2yv2vbhT3R9V5ExrZlN3UhC5Q4pc8AL5OF14P2Q
6edSe9L1sJG7UcT5Il6cdbhpMEpzw6oV2BOXc/s7yOE2mMT6DpIiyjGk0FEEYbnp
oEnOOfBqEC7m9CCnq3+2s6ajqJri6PThtIUfUDBimdFe6tsUfGzX0BaFAvU8mir5
oM5Jicv3fLgGShgngLYHoEdua+DUcu8FZ5TqKjHU+H9fweGawFBW8QwRSqHXUHue
7hmW0emqP+2Xw95TPlrP3WPBoa+9EW/fmXNiTu82Od67LFxYQ2OQ9MwgDHfF8nok
gzn2AU3cHy0xL3+N9Qe6r3TofKu7NoJOMsVlNiKlmWzvhzR9CrYFcb/4LL/E7iJi
RwL6EfGRcfOqtUgaILZ256oax4N5cQhilIU+U5/Njk4CvAwPg8U90UmowhMGsbtV
byVpp5N7uGWDIQeyPJ7KCxpVED3nHso2pJs0j2AYI4p58TLTNQ0mdFrlAO6Xxhh/
WK8i2scUdRWhubUypqTfaWtadojnlWIf9gTeKo0NVf1TqPfq2QMf7ybZtrY9ePb6
6WWCcRP2sAUSCL77HZO03RLNXoh2qmElTn2995jBDAosE+ro7X/xNHvCo2OfcRYq
ibS3h8g2NyjMNdjTvFEjOgMqhZyUg37d8xoxvhtaQH2plLPj7s5w6/BdMlwOuTdr
cDXRNafQJ/U2hb3glRi1p6oQ9YSDoxOTIBQNJLLh2JDsuX9MOuhnDdy9eyULNfrb
9Bq+1kh7P/2zESU1AmdqfbfLJ35ixvPp9KmJrNdqe0ik1oAhm7HFHAL4PrII71O0
LNQnBU2urh2BApegjPn+U3hxawUZfbDU1KmKB9chzaIqmaqPk9/IptLMYMJ3drln
DeWnsX18dpsdI6fZlwQH3gnvRJxBXhlENxo3bynAizqSMxuZ7pUTE2eMFqmBjeGb
YfbTWA0ad4xvprFg9yS7xXvb3DesG6Qa8gx2wvy5cwl42+GTqKw72yI3ptSQhCPl
yFNlnEtkay/2UJm6ajlbWc1uyIjsSc+lT4reBn3X+SANk7yPPgz7HZKJoYb2PeqY
ySCtNkL2WTunKUXKxI363N5cSevRf9GBQJDXAiT3EimJX4hOJzerR9yucAvnqy22
ZLc4nwKQUg2Tvqv23mNU7d4poraKyCcRtI3hMe9GpBhovrCU6VKcuJ2bGca1wmrD
O2nBh7h/A+9QTdimliKrKMLNLM6xiVR+/NENms1x8Rdbz4QcE/ANNV0X81k1/sUL
xrU1Eujp2ZEnW6Nm8xwRK8I7uInjQdvOLHGGKWaTgEccpgskI1ZuIDqQAa7WMWFk
T+eQ3Yze0fgq4FfzxhNePgj/LyHFVgk7p/4GPdy4ssdzDXfN9745s93CT3+lou97
Kgm554yodBTX1aJcxJocUFmFTodra2c4GzNs4RWnB/ZqBYhCjnIAgSLTpxKOfJ9J
skS+aHOXeYLGDE1SM3hTk+AUsZbbHuNoxoquacFRi5OkU8ac8Zo9x6ePwoLyV6Bq
SCSSbDkbfVfeR+eNWoEYQ7hXoCu5OUoXFADAo9qITgoRsODcBaVbyEz09+4xB91C
G5iEfs25LahGBjDwsASk61h/mlKzZo/FCWRHE14kxSxDZXr3fJ/PUyC3HKK+Ve9c
A/njF6FIPAzG5pZjas7mIevPC76QJ+/DzZfIgbVc1Lb2IQ91+tc+bjCW3DtC4BYJ
vbbNdLyr50FyKffI3ufU4qu/0/x266+FSSefT4TkwmoAJ+AhadK2emfv4EuWgK8P
Y7rFTa/c1lV/NlEnjxlkVrnEDpwGs9zCcVLldvHYDXiwAnei9KX4y5CSx//2I2GC
zALI+agqGdDFOVa0cyPmnVkB3qif3U2F1fYwOrHIp9YDhFB35GuhCpbRZU4b6BWi
b6BTB09QUaTptf16WW5O6xfhhyssIe9YdY7Uyf2Thafxqk9xUqxdYJDfZx7audyy
WhLTuOdt4Qv26ss+u2Anq68tS8FSt9UYD3XERZ4rMJWkAycUkDbhdWPbhJu2G9jl
cnyKegz13HFf1HAGCo3k3lq68W7MZKCjx0oVsTsyfBQvaSW1oQLq7SIUv7UvhYM5
8qgUsXT68oN/eFxOnjCVKNs0WNTWRuh9hw5T2cZqfpHIpM0vBFKF03QjGV3wkrGs
n7xUrDfyVsOIZTPV7PPPv/WmeoB4IUIQ3pZ85QsP8wYebzYO7f3bWeMNACMM3DlZ
BRzff3ADIKp9UzvOf8kiXWkc7jEuX8d0+6vtFy8V24GjzbeyS4NgCEzLA6uQp/wc
ycp2PTW5LGvcRc8GrC0qxDMtdjy6C3yGsFLBeIbu5XzObd3quUABTvSbDrz/c8vL
yzXbJYGvGuxHTNAsrE1a40lo8dka5GK+bVMLvaE06gVSHmeBc3jYto+XO7ZD+qgD
wXYll8NV2smUDxBj97tHFXYIdTLOYj5JtBNxnk7qzJIq4xfHDF+HTixtc7mHvJdj
ngVoJ3JMCe+11aZlFCb2OD2h95mtAc/XePAdfEIY351Klta1jYQ12SN2o43QdHgg
FU1MuNjLUoPmJ168qg4ilxAALmWFs915SbCB5OiknkQUzM17nXApOf138A45MXWM
nVlQeaRctrnI5Dv+6Lw5rxDDEAcEFiVKVh8QY+cNkRc9Z2a79Qcyny2BeOdumRad
LQivBw2P6z7LD+fSFIQiRiHeEsLDaL5k1mlw8xmz6h858P7GrTHtjwhK99/AXzXn
et3rHXUlHfAHHyeN2zOgkRfLQ3PNhC9A+WCpUXdrVAIu9Um4isaSVnjJfIm9JR/F
Wcd5vJVl7EHf0miAdHI49f9Hw3x4QAZxv2W3kZpV+aY/+XhUIOf3vQpEdNIW4S4t
MM5TTyGeJ3zMT3KQXTCHl/20VC2jGdvwu7OTERTDE+Gz+W8S/PIqQYQbFSmF7Wcz
vrEkj54V28ufa5xwcnNVzxhEdN1OLXSjpfHjSJwyEkuVf2PIXAQEQmtQm/1FclQn
fMbn/y/zFusJkHVCZQdJSpRbBKIZliDBDAHIZT+I/9z5wb0iam0Vb8c74lpDOP47
D0akpXOkXH2B5cxstcl5iCgtKyli9P8IxspvyMaUpMFBBek+Aj+Gy0HLlO0keIah
1KEwPMD1Ikq1I0nbSUULXyr7kmpC0bX4YcnU4kCsC3e0+Eei207k4JtQumsbg56h
tf2k919sE2octQG0nz6XLSmLfMEuQi8obZHw+qg/7uxYttYw0yOdfZ+Td+i3uQeN
vRYu0/IoDwzCMUE6Evu/IBOvkufk1+bI43HOW3HyuwKlFJ9EoDE0jFG7Bi10thz9
pX9f5qGL5zXdqdQ+aniKnMNoFwTWPNzLjmCSIHelQc1BVU9SFDN3vemf8XI/krZX
23wYFgMW3PCsLrKtTe9FIBioqUY0ZfUHjIolQx80yTLvurXpo4BkkYIqmFOdY/mJ
lFlupn3H6xZYXS8cycNAwj2O85CsKQbLjz19uap7PPefnV5s7V2UTwn7xYFMnhJ1
quFbNzMv8OyPh6qj0/bVHhI2nmNHEciurcIb8ogW8TUw5o3J+mMSEqdlzna+d5w0
TZl04lKdpfAZt7uW7x/l8lHAilVNxIb6fNsGnj9DVRFhTqUqF7L5K/UxMCS86x6i
Zpgy8doHEhHI801Ge+txOQ2dQXt9tvfUTqiJsnCgPEjRrGb7DLsD5OqcRA1btAnj
yf3EZi8LWgtcrTxDOHHhy/sYf/ewLptwAqHVYe7+hHavfm199TS0pCTuIIdcbUQq
Nk0ho1oF9z0SqDC9ZbrQmDismjSt2Ze1hxe7fKr0q0MbxMSD3xjsqswDNqNt1QbX
jWm533PM75qJzaqYpxPnsLiyCXsifjmtjg1MSfs0giz26EUPtYH6QsEfrEbu78HY
801/bWxWDcGpYtzKBGeZ1jpzeOeo2MGj9YO8nFPXaLmis2/MWrrh+P63GI+j1Jrw
x09S3yfdHt1W7+VrEXXyS2bSHgzDeywPQTrJlTgqi2pJADt0kjIsA9IbQzD31wo+
4GrjODt5rEGj2ueV9+V1OM+QdjlTjFkXGpwk6pbF/TFHbzl40pZfKWYKwWThmMD3
pK0ddlFddin7wMnjxsXBC5AA2jpZI1bFLkVbOksdyy+gte2rnPHfXsG+PayLiYl+
moFYrMGZkZqM10Ma7x56WQS7L3T64k8WudP1YtvvxQ3Qmz8Lrq9+KOB8CAOwWQyY
HFuw+QPNe4xShd/EAUCk37OlM0kiSJ91DNgOw/cEkpQa9FHN49mQCQWTmBm7dFCX
C3xg95BHV4sc9HFJKCi8qpGfpwR7qWJK9jr9P/7NpZxWBEtF9owDtDmw6HsS5qCM
Gxf988czmC2mZa/SuaAHvbvEBeXcLd5gGO0Kb720Yf0Kl3w3k5QpNUYIXyLayPcm
IthuLJk/Ac9irYtu8bURMSiHwPMVI2t0hjRemLZKseQL/Bm0jmK/9O1qWYaWNoKV
x/aJisac+PAac1hFpjX7wPT5RfUdIBu9pYXE2v+Dd3MaDGGiHMOL+MtPeF3Qas+P
zPCXOuBp5GDGonhYMJXiHgbk9K5EJ0ywdEeQH65REG+MiPBR6djE1Vfdezj75DGw
tjx3+wqDi9/e0gdGq9hvD2KFnURD9sQj1bmRYL8CEF0cP2OG32ev1/g7exWDMYf5
T0C1fV8mSwERVQnkYQX15YXUi8L7Bl00Y7XztpbJqsIyf8ydAwZVYDICXtxTC03v
Tr9mVHieFzFFFKRIuB6NPIXHapwulcHhsrUtPGUvEDmcliAr306QabtYL5FF38Aq
G8I2sDlAc04olg1jygwY6/XYJ+l5Uqg66YffLASpCioyAzf+AkK+G8bJ9ORrvTDZ
uZuyjuOQCej+q58BNTU2yVFqbTa/49RaOmjFDg5MeqQw+p0m3xKvpQejclZI+xxq
wEqHElQLAgXsch2TbIi5ZdzryT4RUaDjcyFdjsleo7613H3mwcsnIAjdxWuKyY9C
sBl8k40oDv7ayie82QfaD27Wl4ZmXFDG0tuYFmAbrIWc4VxPyYiR5TCnKQ8nEMJz
yRkZy0QnCyHwmWEZuFs8jcFM/WEv9o2eNV5ZKsk3Qwae3TzD1U+fQWbvOpSJW36r
b+b9NNwoo/09WepCtCQb0begSMW7ywzZ7CmmQ835ebP7j/xaWncJPbUs+8SMVB1m
r2ksqSl/g/+lZhmhC9GRopBMflJTBPRS8teOtoqXxuj2k+UCysAa8Cj0PH9Ad0de
gxiuOvdTjLFzGOqzjg0fIxIRGGZ9hC8gmNbWqp3P22BawCpWGVGE2950nmbTsJ1E
HgHLn3uunGgQnkRfQWxrhLOfYwVYKFNbOdNokwWCjfyUNsG3sSNiHClbPsniR2PV
EwIn6y20uPg+zI0Utc0AKzVxaWZsnkC9P1tJWhNa6RPMgUSYm+M1Z+4jqZwvGEu9
DeNIQSdj9QeEdG7Vsly5agCX1FL94odYKPyXuazRkvcKErCKjHHdU4KKrecTN3Ob
y7TnxCr8qV7gv1szRfAkeAvBGQW1L+nHXdFVJiswfOwGycgmtNNiI+Mktegb/KXo
feadsuEu2JgZ+TaCI4vW6I3H2K2MIIgkk16nfQV+V8X99SmOK/DAbNwYhWRvrFD9
93GBwtEL4vbu/1Tlw3ijSHlpyi0rx8L3vdfiWn+8dKRbxF4xjQrH7QDmPifc8tkg
QiJ3fY8GKNL86QjdDb/P5ZqBpqOFdSIz4ucmfsA770YJ5D55rr/K/wK6mIEMChLi
OCvka+uHwf8gMIuQ4Ro534Hh5qYYr9fkNqbChtIvoUDSaGF0KGNv6EM8/EchbsWD
SpiHaA4dorSGEmWGMjgXKrXpwWulcIBpIHT3QMdkd1gAnGdc02BAL62ggUi4CiGv
m8S0XfkuXXtn1Y68CgT3eQG2OOxZ2WAPy18N3ZuJMu3vkNyG4EZ/R001Oue9ZZDL
IHYpxeGSoZ9EKR99rVqr8XozNUm8xxxKqMv286cu8M7cxyAHnIGDeHqRJHdASYJf
ymlW5VNz/PdRoOKpHr7hvC4svCm04C4gJk5MgWX1xDf95hlCXRHab9WJhcOPIrNm
AE+5SSIyKip5D02sAPReOg5LrlOGS9+BgFEvC5YLJHve53856umuUgNBmjG3h+iK
CAUZBAqlwrmcp33xNwVO3yWGOYv2qog+Io0+aV4nH0MO3hhDWeXDnxtvrt4zZiEq
3gNFNkuBbe0RNQE+FYvwk/bwf6Ai6aLqsE8KxWjj4d2XcHVnexQvbMoyWo3RZPZk
SJtEPHfv9uSXHyy5uWlCrvo6JLuKGK2zHTDBtsUtYvBVUu1NhWGmIgNbLR1fP5Zo
phkxXG7Bly51Jma4usYt9AT8D5EmOp4V7xEI+bD+wcnJL7FnAK7lpf4Ui6Mh41TL
Q3oVs4nI1uH/3FwGQ7YzGDKAMkbpW/TODpGt1X85IpVz/04s0dBANP1YUPn8gQDA
PH5IZ8XiCyPP3nA1Re+fqYU/kQTJYYQ8yaq/w6dhvXTovCPKMXXzrc4p3C5anC+m
U0ZsVGDFvBYzVXdtDAuLAHVCsU7xUa69h0pN9LRttirKUPEn0GJ7rqUiCEIivxRq
JdhpG8mcochOaloCixNaZeI02y8tih67AC6qHYK4NCS7nhlfqDeG5Z9yUCzXH5Nr
kpHjD5DQHsh0gnRn0y5424Yk6UyC0EN5BfP9S4eJfRvJR/mjo94VUqNr1HHs1WEU
szI0Jf7yOXgFT1DkdfbgVlU+nKWSfvhiYoTlD0xxsaLhVhkuOR+hNOmV0j8dWGz4
Zaz3w/V8y+xvvBWcITvZUDZjrxDIdPcO10uwOKqQ/mx29SZySpIZmC8MX6dZKFe2
EKXfohAbARNXSkZb/QqCTgnSEGWJPIGt8DLgl7av+QGjm6i8rRaPiVi7ILyLzZVO
G9MpkShJI68tB7dEhzbHhEUg2QwS7/zZR6Sn74/URBWolBbYHlO6VPLuaizUPiQI
gWBOlW8T+hIJmfsAGoMpzEqbxKAN1LtX1eT+gnHTYh+15vsHQZYAPkNWh+dfr9Oi
atZDSGVfZG9nZ91kr+usj0RKruDx0hnsg1jiaI7YW05zZJ4dUdeQA11haJPgW+Gg
n7ewgygIIMHp7Wq5J2lUPgrPrLS1mlCGDS7Ij1GSPq3E5FY+0jNlPzA+76r99y12
W5OSNy9FifbE87vnGNlKuyQbWZqev16TP5NBki0d0NGG7kGXDIjk8h5Tpb4cYaB/
Ntb9nTuERbyKFwZM/FHS4LmDm60lGUjAw7z3ki5j64pqrhkGxjeQP/G2PPQhIE5e
304nNA01anafJ/9hw9Ydp1RfLNhLTcV5ZxdGzSkCjMjiGmzuyVShWJ43nB9VQ4pX
h4MEDq4ma2JeakPpeZzmtiemqqN/H/q41V65u+JRQX7qPtLKmblyDVBFy3IUNfxg
V4P75W4Ihfx8GuMURj0RvoOEcIIp+kIwxoQXLrtdQzs0OtWBs0VEjQMOdQjTQzih
53qyiNfZAInEIHrSFTIyqFOWXqZaE06ztkM9ztAX1BDl8gghDQki303GXXucX0/b
827N/LBfBxdcYM8IgyKXamS7efHOAlUlc/lT9lJJXkYIzowWNNvDRciHG5jZf+uE
uPrEBdxCO0V4F+m3ZjTi0KlC4Herj7PwIfL58iK+3ihGq3Ak518mktRJC7JhvoIb
M5yP53/0gbFjWPwjuOTn8k3eNWXt7RVPOWqmLAW2b9h0X1nboJlvvUeDluNvyoAJ
gsXhbTx05j5TqBxHOo+WGeNKi85aRuxABujZbJK4PWjePPxQ36IaypR5vYGQdALq
vxfwwL1blwTbTMkc/iD0jDjaIYPsPJXGx08OH+WP/8ObkOJ07E2VvSW/S9vDOqcU
YJcczQApCBI0nCE0slkEBWOUAwwtLil8N7o+k3znP8J3C6YVnL+PXXF9csNufcVN
lDM+WPvmbsyiu4qXs9sCVdhKRcyci32q0wRtoqeRbj15P873ome7fyzyEd9xZET9
HDNotFD72Ve6wgfQ2jPhTtkyzQg0uJHBdJRZmk/8E+i44n0Q2e2J8eqfwwUAPcnv
gXK1gn80dvHaua3k+rzyIB1it6+4pgBz3quqcDuXYebLwcgmmJH8bqrhLBvZZSLv
CzT1suQ+YLJSzcPrIOboviVbAEztFzEQkj9d18+WELmAisoNdKkPbzeEwtX2NPIc
xNcUpzQaIGpQy1oNsmJNSjsg5/3nYRKsyvUYVwK4FMma4iJtlZ4mDvp6ifk9/j6Z
AkVL4J0CtRf9BctDT8e1wdbvFcOjcW79olj7LpJmQaY9WChbuglVYvpkv2ndC+39
r3E7QqEc4tYdAGR87kZGFJK+Ic0Gtxn+KEMNX7FTeGr1JzbhPC5JT6nFZ0KclPQ+
SbXnKUMQFk5r5o5zFiH7qZCR+bNnGbZ3PQU3EsrrKJGaxwfZXKO5DaYjkGVjJR0b
zrri9spEipVBQlMi9IdwQu6kJc3xi7G70UoVuq56t+7qW/jvIwE/9NzlSDvJXhuB
Wy3d6Udffc7mumNoOVLtoRz2QL4d1/ZufWSQdQRv3xhUbUOVxM2o1roBFqqxz9G9
r1I3THVjBIkOrQt1D2a/1PXD8XoMazEyFvg+p0hMsgwyK0W8aRC7PtHQI8BnIwcR
/JjMT98PHIMS/MxKcCn/d1EB37bnM8kmRfCFdUZmRUsHivw5/q8qWdU3AzMhNCRX
lQ8TLLxM5XOaTMGvz6uqar2cNgXJxM9iyFnDAgAzVukWIfnpJUnerZKXufQteBZJ
MX6FWivxjC5CzbjwNUHI2kmLQqU5y5J98w6Y1Mf4xvK0b/Tv58FxEWT+B6DIdWF0
6Lr6kdk4x+JcAk3cyshVJlqbxXizoPfbuig47whrRByCnK8sJOQ0LU+txxP4nMRs
MtPVPcGitdaq9hC1KUWHtDnBsI313tm2bXHxarApwhl7fAF+aBJVw1N3lAhJbhNX
K2JDoV4nAns0kFl+InHlq56tQSIynxQ5abTZ147yT0grWvS3c0EWom2L3Asd4bYe
XnlNqr3pN/BPMidpirrRii1oDlvx9/Fp4KkKJMJlKJrljVZuRxSXW0telQXTCpsk
72xpGrbQjbfHbFu8NWH2TDHLCFlaHakp5lBL10QEa+L2N//zdXRdmwF1lwwMYB8N
fVesPwbXpoYVQls73x0YoKsNF+5MocZHVMsirnQrqeTZVsLJfjVwpVErHeOE+1A5
9Pn1ozrcMHtqGwLI3HxN41Bbuu23Ty508s6Ozr6kvDqKa9kw7+uRHHKzd9CoAxDX
/RYEFzt+K8QmYncDrY0KIJ/lr3ET976ow7jFLnIlmt8B4+Fv90U1L9htKXLwUxIl
8IcgvuUbYHprk5+nY3tEHLcFtkd/vTMuIMzL4cru4C1ZFMi2vpB/hgwZ9GeNMvHo
X7793FSYgd+TJ8s4eda7TFI70uT+nEG5axQDhdt4fWF41LHsHR62vvu71G7gl5Y1
Fn9jujM8bG3FH7TzckW7kNMN6PAOwDcQOY0Roc2UIajqyOyozTcOXd/LGOwExAJ4
Xq3fvUBbT0cW3u4HIfJYUlgiO93rVTPZXtiL/9QkbyDveMOUixgdOG6mKpotoL6z
CDFZXSoAsrl0IUJgBJVu+BjIGPtWQuI4MVf4A03fTpADfT0yxwwrA2bGLDkEiMy4
MMAWaFTK5sUiItGLFxjQX8m/akMvyyEZkCoLHcgoTnwedpCKNmNAVvGYPQak9R2X
VXCEY6sZOXxnB07Y9nDb+Mmn960uNrkqYuJkQRwJZfC98j9nldPzbZ4K1K3HKBfQ
SIoXLmqLy4vBFSjcfTXkDYPNM43P/fORzTsHpfSeb/xw8IsnvBNEsAVKi8yWe3y8
S1sBqb3SMN0wxZTA1/2B1bwb/WUBaQtTYm0oXrkufU/WsAjxV47KBpvUo3wlqh2w
XUzYCT7gIwq+9MslbMgrWyV5zlHUyQ09ZEmneqEC0ixOelidZh8syrTidBAQzPXF
lK63ScKx3OHrzLd9udAHLrlIsqbqetOfj5n+DapqxuZ7A+r/pFf5g6fF9KUNmGBb
ZAL5a8Rz4jpISSYhuuWNTVrk6tDYqBZSSwlJVjFCbDuzXHysBG48X4mBwicVxkk+
IrFC3pgkB0o5YNOueNW0P4kxjQpyVVN3Kh8u+CNA61v4MpjxNtmRqhPX6Q/x8oDG
q6DIexbgc49e1PI8dTCbGt8vgOEIXgTKmLrDXMLX+YClvt8xGTCG7e0xvG5HAfVA
NWadxtBdUrjyCXuIdbII2HwDyjuLlUln3GAwd14LkA26cYrehAROQjQspOyEvL6f
FJiFxTQHFCzQIg98d7rKdaqwTrkziJcWlzaO2tDnuobMwLzHrGVRw/slR+L7gkbY
QxxePRqteet+enp5YNJbJ1GTDoLc48iSJCAIiAg4mziuc46IrPvECpYXy+62yMY5
ovTSVorT4qzKGXcvt0PWKSPiFxCvHx4tLCW/I3UwtU8vWEYzytDzlbTexLxJ8Od2
8GmHBLppLlKp9MD9ST77AnMmIpHR5RkEqQz0Wa5uou8liADAFC7jdfHNy44+icn3
DbaL+EjYqYeEJ6MvbaJk7FeHN6rX2Ys4Lhk10lfR21baWOTG4JylFZa1cxpjODMv
WYfhi6QbAF2TSZUTOfonKnHTRmms1EzBYHsXB571oB7NwzVCQsKKiLLo3JnB1Fsg
cPGq5pigJbzaeGHZIFOgwtgl3H6LBY5Jst/bQhl0RrV8jXGi5EZz4XP9Zjekh1G6
h2j56cRQE2mD9/p8CULNDjRQrz7xX8CitX63YHrSDDqMLVzGoOG9Kr6lgW5Hv7rh
JtEvJJJHFr6OynQxgnfaWU24oyJl8c+8lpcqjmG9gRV0hOOpWCqUQ8XPVaynxWCI
MHy4D+/cFzf+/LH35cBhs/QcYlJXcj8ZEno2P6mM61gAOlXawY6b7j7YeAql9o2P
Si7hdGL/5iAOlnj5/LpX+uWj3+1psmcUA+2KEIUNkpoYJNTzGteQJIYlpcCsa8pd
YQve8Shj+1WRI0PnE8QekGresVi7VH9TxIjz1mHKp5kQyxEIb8isQM7zL00s+NPt
7U5gX/E5yT/OmlrqykjK8VuB9/mbGcbfP9I8eSHEFJM7mHrhbfjBrwMhMAPJnXT8
VIxS3ikHEUmrxkuK1VBfzwxGfEE8ua9TXwB1VNV2FCGiuKj3TAsrJBnS41cWbGf7
k6jJhyP+x2wkQ0moGTG28G5Xe0IKrN3Ubf/Hy+dP2uDa3W7OGIs+KlWZrgPhpI2Z
jETUzWfSqM3dvVuTmhWbUx2C/cr5urzhllOjf406ErIrpV95LCrw+ui2z1xtBs0h
0uVj5L12lRFmcKNgljjrN4v1vo0Q/hDIeB+8zySBusOOZ/rV0rqzcj8cccltwsLr
wS6g8x7VjHiXDgJKnP4sTOwbxAKv5ax/yuv6kUFENJN33kCZLtKxhzglO/6UJkm4
BPBOdystuhJSIEHDZyu09idhFdXZELEdTD++xHDUBv30029Nfh0QBwgnJwaZUfuJ
cZD254PtH4EJcDF5AzrqXni4w6Kz7tpgFAOI+JPyZmNOxErHQo1SZs8ONl9pa2FL
3ObyThkSngOlmzGBPTJ7c/QVG3/JX+EDDy3aNoKe9kaDGzSm05BduXGCS6EEGHsf
L3H8BsVVhs9++zIauarnl3hETUE51YM0p4eLwe3P6+yJL3jCj5FqjsCP+DSfy42b
5hGBxKa2AU9yQtIb1QcM9HGlpPYENHsZFgdaT49vccF2m6uxxIMfS0BVWCuPnaM0
EAy911HS/DZou5FEUl1i9plGySxDwrl6dITtKABtxh4XpqCnJnanc8pXZ3Fyv+zA
EWTomCgxuJBIS0xDByyyspPEib/0Sd1TG8wQjm5p1kdwv94FHiD6VMnCKq2TNCF6
fO7OMCHgVi1/fHl2I+WYhSJWvJh6TBbAuYDSRc0FNAMopfr6VZ3FPZ+2A5xufSXo
mY3MQc4izoXMmC2yv4o2S9oNL3FvchqV6NaOeKE7IvlpAgmvmWV4VtvtG2xvfpiQ
FYA76ucNzEYQvU8PeKvyqgPraqrp6+RrNQue2yUH//13+4kC5spLlPfYtEGPqiga
LvspSZ019uK5Z4Tm69AbHbcgi5a1uZbpXVhDZw8vLPjLbqLCSnAQEOnT+OfIOm9G
KJcuZy2Xn3/Ae4qsCVcGiAMF9PVmhD2qYCHN+Uvn9jxYAx2L2vJjlICixMXBiWl2
Tri5owsxwAGLy0Lt0jhT53yJ/K1DFKOISU2QudT2i3oQTyUf+NJ4CSYnzF60Q/Cw
qc9bSimY5BquBO3NdJdBG4LA9drd7Uk8WgSqGbCjGKU61lvx8VBEudrzdgEtLsEz
4gl7TtjbfJ2bCRWPh8zpKDc22X+bmViDOAXpz++PD5wNHcBID83Zhs9htflByyZN
KForO4zW9sWDwP8jb/1Qgu5TjtWDq0OSjxF1uQYeyKh84eVzgzL8TGbQwHLrBudc
5e9sz0TCR+omYl+a3JbKUu9TxQg4OBM1bGpWFN9Ev+KButALrYzpesY26QlIRQiI
FSGNR6Yey3D7Xq1rvfK04b6dZaqGq5FOojy2ibVIOptprkQjW+1OcURnN7JzSXjQ
PwhHN30hhGJ/JkWQ2+3vrO8C3aNE0lb5n7ZYlEgr2+1SKR++rU9fYKn9+y3ObUKC
vGvo6bcua/0C4kq/uOzdTfZksbeKpBM62ZQaFkgueYRL7dfyHAIkQ9+VeXSwsdIb
jxqEdmgk2+oZjU/uboNJEORuuiGsOLZV1ya9SloUIMVy1Hl05oIu8lsH3ycy+Yea
QWc/BzUH92/r4k/yuDJfP85b7IEDFk41NPHOOaupmMbu9ZbtHhkRSvtoNJzcFT3W
/xNHvDTPanijP1oaxLBbgCIVz/gmzRbH467KwE1QG8aRG0cJWEC1qui3MfXQaD6c
qteg/uyQn/Q1T/MN6X5bkubCYItK6LdZNIhHnGJdnr1aiyk9/PyWDnahVbY0fhKq
OXmb+9MqmbGAKIfBBJU9fAkC6aCLBdqiWOf78gP1M8Y/ioDoJc7DJFpklyYLh5dp
R2enxk+7oCLqEXV5P5cuc/5kDq6/rP2IffRKYWzMgG7ya2ijCDECaFXTvKllDYPo
yGjmzSVq2i5isrSrIjZydj68urcb3fSQYt5Hh27YjMJXszd2sMDMXkcLIDZShvlP
/KSffcVvQGexm4302nbzBLFSr9VI/Fu8YObuyyzbafRFPMl/okoywZ8g2u/ToLYR
Nnp3bvQgpTd7ZDwZCRJM3jaZigrDdA9HxFMTaO39NHLxWjPR0o5UE4D5gaPGtLKv
FxgXL3FhWdfcajtCCVvNZXr+QUdya/hMCJ/sJTGiqjxZev7joWDpb84gYtYKOdih
Xvuf0mAGg6ItwLozEq67wixkrld7Vr2JXT7QTZ+kIPPcNqBo6MQxCqB17HnbQYnH
hRodLd5N8LRjBoA4moE2Qv9ru6IXl2B2JjvcRuv9CjkwSIUodAFhTyK2b+8fKbXK
JxfkgTATSfc71y1HAMQSIb1j/6jVA+7SmPcGPRVzmhEsS3k1C1sJNn5oWsC+iY57
R8kBu+FDwL+gZAjF9EMwRMkyzZobyEZzhHDMX/LZIwVbPGzz42Rhd3iNWsWVJAwe
oVeCz9wD2QwZaDGDv5+ovPLssZC8NvJDImw09qOHR/b8KZowjnt+xPiAcC/R3MYk
d87p7s3OVllbP9zDPIe5BDdhX5rpjaoGSFQ8xsswkso4z2IAkrPAqL5uT8ciJbi/
FMxJ2U0eFiJn2+Z+AOiLmQBD9/7MCbb0Qkv+40GXyIEhuTr5zhwPdmLkd/eHACgT
4aibNOHbzWj/KhWHbJKqpszvPKQDNKVhZIERA6hIWYExE/Qkci2fsvun+zcbyiKN
O5QpR9k6y3V/MbwOH3GRRqvgtEvkMGrnPz4+mEefHfCTu01Rcgz06zrL8shTq8Yc
v+pN6s+y2hSLSAz11g9sJoEjBDCv6I72zWhJpzrhEGvLrNCqYJM0JYkKoDxfxbrn
6+j62sJkJq3l9HvdEZvtSjy29HSzim6UyfC+ijPYln1cHrWzNRmkTj2hVKz1InQ4
7UTDEMymmFEtwTMysq6k7WzgoIxOpZTzq1j9cEpES1I3xkZ7qLFWHG1tXdRJH0ZP
LghV9QtHD1iuadvxOw6NQDfwzS06OpT9By4OGHJk8XC1/xVb+W3URV9GhOiIYgwL
4hhKkIbw2HypgU4VhHi/A38DGFbAbU1nYxGW5h72jQeHYnRfXfThr6KDpDKftsIl
hiYjAeb5/3kfR9XxB2HoGaWGCZAzc0hydMxtcNvqbln2WPmJHkZ+3fWkv87Xoc2D
tbryXdqlmNqZz07Xv15AnM/xJpvTruEDczwBfwQ2J75CYKfvncLIv4DHkRn0Kjw2
fqaVGy4BWzL5GARUB8oEDi1fsetxyXBZ1nMun0U3B3otPd13HnMeWqpCmbls/fOx
N3nWubCPD/gKKV4mJk6mQpVcPNvMbBoYdJWAoVTSRZhsT755eleayI6u9wleDptV
aQXB6E6NRx5PuWDKddOqQqefIzM1Wm6tmJWuXxrQb0DpD2XFLiS8MawBI9O6ruWZ
GE6yU8roI9uO0yAHx1dVtP0kjXzmv+63AD6S1qzl0rySIJxnamxSXMSZr/ORnJpw
TuC5r+LQjga5zeAdIdVo0E1N8qZ5fqUknLlej7I7QmHiLtnw0SJVshb0Or6faGlj
wLGL1ktQpHlTIGXM9Kkys6iYn7Y08n5NHBib8UcOVdngCcwNzdrqlg3btCSpr8sZ
7wgy1uMBj26h5zRCgHbBkLuQWVJnVPv7EjbOsrM07hy3dBcb4cMFUHX12A/32+tM
PLQjpH36/riCph8LyVkfme15RBfI3BhpFMaP7W3trkCqnF3b9QH7AUGNoK2fBUY2
Qx7Yjis1rJSzMH9Rw1KLG2bbAu9q10YxBINX8+Gmzo/qi8iqXKu9GctK2BoPeDvp
9hUYI/MKQQ8FgYj90ThkbDP6HJaxdtd00s/w9MXrHo0lI476KbMbdJFtqaHiWJn3
FqBDeTl3gLSll6A/J1rZ50TbWI5F9czAJxuQKtgKRQL9117p/GEGVDW5T2nkQ8WL
Xg82Q09SrqnCy1wwx/ZtDtyiASwyB9C/sCsxQdRdBmMshODaPbXsgXB/tqhaIGXP
sr2XJKZybd8iyLSWSFyLcXXZdFKniUFUjJ9gTIxj3MZiSL/RZhJBJbmYgZ3pGG6R
YSSmqxjA/JIibOUhDrMqjdgrCJ1Pwrck8smiMaBEKITBFtCudh/sLbkipLfApFOI
i2HSn0T+JKmmOVEzDTmIwO9/lbBYKeUCvZ6FASZHvT3ScAormU73pOicnskLCb4A
nSSgMp+K7/DgnkwSfLV08Z8OwNcNMkNIXMwbNkE5uqF0J0NzB/aR1OVMkCUKYn0i
cEmBm2a5+HnVEgsEWP9QRTfqgQu5NkitV2SGg41AnuhWrxq/JzNKhM7A7AI8n1VD
uggTtb75YGVW9nQA4zucJchUKO7PMR2kuNQYo9zO0HbGDzH6fdfzbeuYi+3z6cR8
Kw53ZSgpTqZlnJPeqr/eFsV1zFxNzUYt80nMb+GEvsWsrzb34P+C+9lsLlUTZnKb
d60iRydeqZgTiEqJsyHf5o7hwZS2iQpU4C5PhaUthjSTPeTU686Wbv48xqFbRWu3
WtY9Y/mqSGZE3iQEerM227huvYvFxWkRd/8A16qdSwUAR5ejAwk2JeyZe5jWx0E/
lKXUs64rB4NlAORkpiskBZm30lRmSy2ggzKZ/t7pim2KmSsE0vXT2rzksZDooMOl
WUWsQ/JNB6tdBrVl51rENRs1IJBtlIqc1jJ7ng0FYq6SOv5gXMfzfFksEjvIO/a+
VCrZ4GqOK323E++e7Bg5FD1BHJvqhzp7Nf2wWGQcvc8hiorzzPqEcUnzW2+j5LAG
p9Ll4+/KlSAudPTKriOI55wOUDz06z0iE970tK/UmMuuc0QCFsT0L19YF3O8RNBZ
Na3VAbl07Ayam72MbQT4XjqYNZzhRBj6KzCXnjG8y6cb4z2iLOTJfeuN5LTuxIKY
VC6yDhQdx5yiciyi+MQjiVFkepFDu3HoonDfHIBR99KReMEvkSyPIAPXb89l6Y0I
IXL5dxmGXUZ0dAGEUUFioLz4zWPG5BSB+a3jdJdxYAe9DhKTrDe2piqQe4PyqlWq
ALJn6EyD6EVFLOdsrceNH2lArwhsBWZ3okZI/PeylnlTjAvyHiP0MTOi/GxMrFoM
bIKMq25jLSMTnRlCCRFPyr2nCNnHTO3QjgpnDTOXqh0Ha7rj7CTn8lUgTpnmIEWw
LdHyF0YEjPi8E+dSV8woYTM/due9WisPs7pcfC4Q9il8t+TyGSqmWOaLXY9bC0l4
jFTeaEipuvAjzppPE8Re6Q1JR2r7sI6emzoYHT9BcN7OV00UU6N4Vz0InWSwMKhK
pLJIpAJrweYleR2NTXnZTaUKIUgfc+mGGHpSekvtkzIAmXIAodtp62e779jcDmB4
DR6ZZ2l5kZJt5jXJknQF5RS+3S/DhO3HGJjwfgw8okzHd0WWem2MH+IZBHLkLP4C
TPj/iLQsCUYN2BYZCLnVjYx4ZGvAnI0tQfYPxAdbvP99UFD60utYwEQ/TxWu9kCw
sSwvmTy9/JEX84tOK2eQdCrXSZBmRSsWaV5yyC97fKCtpoDYYZeOluVuYRECcWVz
gl/nW/50P5BcwsiqwxyZwWPUfn5m0SqMcNCAZMyjICeam+deP9XkW8/pqKP993b9
3Ub6jft3Bauh42MjW3wE3mUyP6IiatMXsdBczf+CLDYv7C7gK1BbohqW/ttEOrFw
QAvIp8Jo25K26rRvtd6TYFQobHBNjkNEPiqxlzbe4/adLM+0p4YOQG78l3hwpinp
RGQIFDRpWOc31TWpkJGySJDVVz0FbgBeEpeuzAvgqz0rPs9cH7OZQ3QU+IxuKOXQ
B7DVRNrDyDgUQcc29XCDVFPRthgR4UEM6k5Z9Z66ijr/85SpdtNVBVFPw6vNJZCu
6MDrEDUd9QVzG5t3eMQeS9iuqJFgFtNu+Gm3rfoSt2pqd7wuvkX2KXJW97sEHrsy
Npvzt0WmAgQrrZuSl/HCBHYB3mbx/jdkJPWngUAJnE+rZpqyFmqpq4yGPF8Sr/E6
YWxKbyTJu7flHQlokrq7xUeUvK/ABHPfIKhSDKCBJhwj9WiwEYgXL+nWtraU+McO
OIQQHxBQBK/Ms9K2DQ+NfdbC8zjQ8y9TdofRYY/z3kubpJTK9RCs/qlSEdSGh7b/
5+zEglN6be3traSnoMQAnwfAKyzmOF8Ys7MVxtGGPdn/0XJXuYV4Ww/d7ZABiKfD
H6yiGleyYHRNBLm/4N4r6Y/r+ex07Wwklu0kkqDDx2wpLGwKT+vajvy/t6hwToUa
Wr08pvK8U3QUZ0htkHfWry7ZZ/ZNeszgBonLD6D+NKELQfE4oU3a7Yl0Dk7E+i2M
gGhVEWAipO1/SBnNJZyXoXdhZDQi+w+Q48PyGl+6lkhrQn15/8rv89KJjZJWKXca
8e2PsJc63MUbeAJv9uKkQY4xl9jwm/5VYIvNRPUyZZqExJByErROtLxOaZkkkxxi
sm4WOX9upbgZBe+bUXn1oElLMjcJ7/4Mi4IWuA2pbrbA7bTNF7gUU0peI9g1h/Xt
AOWrJ75JjyKoVhioS6+tEMW8kzGz1bByoTAL8vc5y+5iO/cmHIdrG4Tqx67+eNDx
IJU6SukQDL1d2NL1yGzel6yH1qTvfnai8QXenQPZWxb1afYfwZYHLxQ+R1fg7fwn
i9XwCsG8clWrS1OYxYSekxyG0TAnYU1xXx9srNIFEroy1gbEN2hA7N9V7b21X1c1
slWWaGVXE9xuB8EstGdHEwje9F3OJSn8sYLvj0sTEMOneJ1Tn/0oQ8Rfo7Bm+jm3
kFfTXgTJGKoD+HMZhuA4naPbDgB9Qf9nxz3K2lOuY8sWeBwlgMjPua+mjf4PchTh
+yVps5yUwEd4kIARc9B7mi48I+0VsDWjwpNPEFXc0VTavXDmuC+s5HLZxrtBLd1/
tjRHLru3/bBexGM7PlepbieWXDp0UtB4B/6lbMeh4BWpDLHjVY7L8gnBx9p8q+uF
8VUHWNjSLWxlJgXh6dfhB5NpRoDnZS2RCnQwY1gPBXi1v71HQYbTTudzl5tGwUiY
xLJ+3YnqVnMubT8acnw/igszxzyfsEkxD+xWS1Jsv9pUQZpX3pHlp1IY8OtNv0g0
1ITKtKnKwUR8dWFBF1y07u2qO+2wAqQVJQ39RzKppCQ8Z0pDG6/9csuSj3klue2y
hib/rh7YKOWpNlITSnHz4SNH0fkWQcuGdaRxUGP+WgXkjrYmoLbX4gXlB9e+vpN1
evkKd1ISzu3MOvs8fxkUll57jEmh8FOShcRQyYbT2iWRoawAp1nqkxGLimkoUWMe
Y/9hAHn/otYb+20pEt1vEoq/d6UU/qxEMMK5bWzlcI1n5ygDwhKCsgCpuK5AsE2E
zf3Fpap+EPy9ufqM7EeeiDWkyDHlT1imJkmV9bEdLU1vQtHXsgfFkfY9NqE6IXZj
+MgefY3878yX4zLy8pSYOTG4Ss+VCorKVRdvw83qWDkDaBfIZLJLzWXvgxW0xYJm
vTYdOoTimWnnt7GlOe1bDzGmDI9sNtn0LStWdt+4WI3hN66Lln0eUor0S52kSDle
1cvulP3z3o7jEcYWz8eYUK89GxPWkYrxI8hkNquJZMyLAurvaFtW/h+RXy8PGdCB
fADbhgnmV5PeCSjifxEYpsSiQCGGsptWRsW6qaYvztmhr3CPZ6m0g+uU+SnQPuvJ
MxItX3Hn29ggt9BYMbuB5NHJzi5wln3QUymvkK8xC3TY5FSkzYant4YLm92ZN/hN
EH88SPbPKKK6iKuda8PROFCB7Hils1QEPx/uQkjUFLx8A3dtbEO2TCrr0pTjht4z
XzPVi15bHbRqadQNCAnuNooGY77Xas2zRS4fUbkbEJlwDTb3SdebB8PAPXr8vnEd
9T6wbZe6ATlxmkEkKP/B558tuAtIjwR05ZuZShoSlzHgmRApxM5+mgdKbRuLPu0N
xe/H0J3NNyFolDGddxf8zEKmHYFVLVL8YEWTDpG3O3zCIgOeUaEedfA2oJbjX98Q
wOy9wxcDcUkTDFISnZqdXzHOwbHcysm3TfJ1IXtT3CrflElRyA8nC9DeShFDGZ60
n2gWOSQWi4GZTtvDgiCoMO2pZGKfMrvzy7ChUOTUAKCJdRkIV3CSpkcDXw2jZ+g3
ewxWKUmU7QszgA84vGfdZ+8ivO4KV6NnXsPQzFjj9yswbYQX8EYme5k/MOZgIcfT
/NAuLivbJ6qHCj8wj03wonKUH5YfQrZfcQ8PFW6xN4IjJe/myJ/9NqpU63lqvmvW
KT2l8pUyhbzF+vi5jZb+BKGLMMPZiB3gbCBFXZT4D+oL3xQqSw+JCkVvErx6A1/+
ojjU1ysIWoDu4Vw3ZxRkNuhn0/BPBzCBHghtD7cNHYpMVJwXRdEpHbM1ghh82F41
zVdr+prgeCdWa0XamUlHLYHXWb7DIjivskfFASd+r+amP5T2vj8eY0aj7oHKwSCf
Ks2jGM2daFY3Hsj99D0SeC2ortgX82IUFpEizKGQYcVOe90pdJ3TvlLulkJEEfoU
rGwc3m5hzEVQkGx04UBWnhPvhk6PRrL1DgfTPXWrMFL95nbRn5HojXZjD0tK9C3J
zj4kcgA4Wfv+2XBrmKMkf871b7lSFQtU1HnNGOrmpYhN0/pp++2ciDp9LnX1u7Du
Kd5swksva9J5NVQhKCtgajqOnn4wNK3RNzHDRKPQGZmQimOOwywxqvz8a3xeCIFo
Qpuo/AD9flENRO233IVGVcnIDBjQNrX8Z8IKOEQ8MJEJmKq4lgApJw4SEx2avNOq
4rZteq1bwtaKASqUY61Q9c325BnJzEfQsI2rP1/slcbR6mhsrsLF2iaDCWiR4EAb
RweDlSQkyLi2BqXokZcPwCYxDc7E1srin9Bdg8dNdoQbj3hqY4GUEHxa3OfkvYXu
NY2QxBj6ZsaQzX1gzwqP/wZuir8MprNrqQIXASpnkJBd2Xe33ZxGHQmhBSOKNj99
VQWzmdCHAqSKcY94Qpo5/se5UXf5Ir+S+//cqpAgrWmy0NQNHWCE0FfgRIjMVEeV
b5oSvwxoJ+ctOYuSyweQViilymkTAFExZxfWi9AIddnrKtBaSQK2/UfbkKwCItLP
Ll8zeCbh+79n/HJFd1Fjcrm2BV83+ZHuem1EQvZpaMZnLzN9XC5XyGrRpUudccga
PW9eiviS0j1pHnjc0N9JE2+hR0lg9HHO+K/8938v1YsjD94KUzP6/U2CV0Rn1moc
4pyvelrzwZnqI3ApzgSJs/Y9uH2PsPk4lHrK2+hF5xWzn+toJL6rKGnlLpXbP0YA
wIMIsiC/2AbPuTOCL60oN+25GYJ4FZeaRN9mzERm290HAzhR5ea0yXaHB+7nQ8os
CZVJLhThOv4MRC7iGFkXbb7muZQQ14MbqbnFnbiHLeWu7SGn0akVekZIrl/ds7yv
SF6OZyqFSXp/b34Gi2k7fU+nB1N+gurrPqljrVLbblfdhTEjGHfcnk8a2JcI5TmA
5gmTtrj6JgOOLlIHswt4RsjH/tSyT52H5dC3BPWq6llzJsqsOx+KWZX/Q67PPanG
iMi4aXfLi7W8yLXWdB8dFprNgw9sAusLWUPC38CR0q5/EIf978ApL35Jb3xWaBcs
bCRCaIet3ywTnqPw0r2756jgIA1ypqjlCeOfazdwyoly1pyK/OrSmisBQ3DNDP9b
+Z+cZjiMiQye2/GgsHKKt+b4FYowbtoxMder3oHnsb3jBNTKuRLCYFYPIw5asoH+
L4wjkMHk6fRYWkGLSEIsF3PGeWgBcDte5GNrS0jt2gcMVRiHOFCQOC9dwHus7F/S
J0/nfWiaphJsb7p3Q2XejfskSU9i13Nq9dnY7rC2ux0cUQv3Nb3YZoxk+mTk/nFk
BEyvT5HS4NlgIZtaZPv2zhgM1J/z69Yb/UNwwrU/gas5wQRnfX/WaVBW+t6ZU8jR
vyglrJZufjuBE1ayWuY3aYpgFuWCXK8Bpd/csphafOJcbLpuRkicbDMJPb7vPOVX
ByNjdx5QN6RdEVqb77rDkh2jtzJxbKBoCs9FtWaTNmDK7O2jgeqtlxRB0vZY2Pof
fs+vyiaEwFgZ3GAqcj0SFxwTRCDVlKB0tnZfNJyT5j/fFFZ65KMU5VrJdOlO2Gp/
Y7Kb7lTf+u6AaFLOn8vsUrM0Ru6Q56r+TecyoZTtNCMg7ZzlV4NRqjgGXrHZ+xB4
hTDbuBnfaGIGm/pMf5HT+NgleLLIDRfMeYqWUAPcGeFwk3zlgULUfLHry9s2mPXl
eTx3o9R+jqeblhZT34g9KDtamNq9RZwv0WJVDYB+ecw4qR/dOCXebbuBDywvqjkt
1vva9CtIbhnPVk9LKoX7C7VW2nZVJxl0lXaOaF9RudoWVB7ZgVBFLBfTqql0XZ/T
gziGgsvu6d5BriMtZw7r045KiQOy4V5J/naI9xp/h/xzVPY+os45wubvOZLbq29q
X9u8njBgS1Ypmh7+kPY/oEdIozcZBANIFV6BEBoxOpXcNZd5rPNSPm/ZuMb6KyOI
zpdcqjR32xXgoRuCGrgLDdmlVsemDy67meoa4JFN5esF91e1XgNov5QuaHbiVMza
IFkDuzs7LUMN03YWbOQUvZ5MrJP0gVkts4xU8md7cOLDbDDIif/ersOzh4fwt8lP
FE3RCeOOC0DmMyJakkf7iZLR+c1zNKHaKHgbxTIVUE+VEV16rWIz7i6ObN6th2xF
0ygZi2YGHS2Q3r7+RJVrLCGkCdlsXsXt2cyClcsbKeUMT2UfisXU4vu5/cBut8Bc
oOqZJhktif+kFpFYeZRQKX9YSPMF9NVYHMfGkfT4+oO1bkgOp6txGLugjL+sDyvD
TC/pRYjkz27LI4UoeH+M9W80xAGGLwKKqGISZ6I/ri5QAAPHm3fmw7quwTirPPgQ
Uq0cGm5uskCEZXPSGcDA6hPcMibN8tXLtWVHib1cTK2FDjJ0zDTqEfhZOARfDF8q
TPqYAW44wz1l83jeH7lSHrp6zyedzyBerQ/ReZbNN4CQ4V20rcAj0u+RE/XN07/b
0wqoZnKwCXgKbZLi4eiVQMNp5jIs5locW7nla7rT2EVfrF3h0sim4QEZrNsLjEVi
MxcMZ62jvgAhBge96FYaYR5dqXbeZv4aewm3ud5n3jW3jEZjd76zGduLwCcyYbzh
GRHzoR1GAg0wyBPE8uF0b0aFD5SFkohNs9Qa2B/ZxvJM6uISG0cwwuIZ7YV7LBv9
SRDZs/qAUR4pJfGx241aDsC5jw3cVkJLVgjHOOJi+nbBZxtG+rr9N8ul8rXDNrEC
iIGiuFpdvNNlXNlr1VXwHyjIAwjnBrtx5On1TSJ7e7csCGNIBcmiE1e7P4D8y5fh
SC7mrIjlynZanEst5YX3ewh0Ik6POQAgN/mbWHMJ811aN+wlhHXUVow0Ex6ko7xD
o2bFIkrhpvBDvp0jz8gxq6TsI3LwAazcSfGpV3PZQTZEeou3EKwXmgVEiSBqT35D
l5MU3FPvz/EqylW4Yt+u5Cx2a2XHwb9dYjW0I5TVjPePl4mR3B9RouCipjUedWaT
RhtjS8HxZvWTEdvoC87S715hAe1LBe2C2osVvO6FudbB1FdrSTIzV5raPqu7tiDk
WZc660PgO4nIdcU1rdpvZoWCLyfqO21MpwjHnRFe8PnUDWfEwUPHY0jYfcyqz3QA
7WMerbwZgcbrFaYJk/zGHo9bGSM8kBethAfYHCXIoJiG6dJ+aGyLgDRcfAiS/Sbm
ZlC3ihW9Rv4CCk1k+FwlbZILeQgckzfc2ZxygiHzkwwylnY4eRuExT/V1ymyVdFu
ZTk/enwBoR7NEAKNMDMH4jVU0Ld1PMD6lkHzFtaLLoUbZcYtSAodjtKBjoEePzha
a+/33YMCf43UyZjAURL5ELSfCae/aiOIpFinQfZqXJZYQun22DYdfaDkEg/LFzvm
2qXCDsSztlo8gnTTttgAivrwEme4fwS8C97tNlCKqsX5iyraSHSUZlbyqORCEQpj
qKiUaAnOCT4b8G4bC4VFjwBIyJ9DaFHnoH6IainOxClJvrvQSjFY6JvLccX2mykr
GCm82X3m0aQR8KX89elLBT8EZ3dO0LIU/+ROSQt5QawBYudXhELBaaQQveEIFsjJ
64u8IFNRfFUaxg+nfyadT6ALMfIG/O+dlpJuLePLpkmFWt/4dDGUdLS4Lg1YRo4X
GGafv7krWkLe23/TSqNiwazu38k2nKLz60cA1+BbRKKzZ6TIVfhHQoAkVtVbHQJ3
SVs79f1Uth3E+ok4tuS8C236vIp87n8/r+d3fuCWoKVv45tqGo8JXCzjL2apkJjs
92ps4L9YeZZ1mS49Vn6J0yifQ+Zn/C3kXejM2MQrmyolESYbI52JhbfxjSHfklDK
gQpiYYoA75jDC7oS8WqpxxeO6wXPyz7OSDZPTpIUP9NCOokdkzb/7R+JI/1jz/AE
s3QPplIO4WlnlE5vuApEmaLjK6400bnbQfFaWZXFZP3TqYB4lRORxmV5C/YAfxtN
P5Rv7gAJz3AblDCftTZt/6bDt7z5ZfO5ENqSiro6gKoApwySliD0wvhuVEo033Kf
aKIJWfdM2SHKdMZYh22es6GH2GcLbo/DIDfNohyfby6IzyoDS84Tt6FABa1b+oJX
BRcVjIprNhPeBvsYKrfbPGSwfRbHJRTJi3gA6aOW5c9nRTHUDW0ifV46yhbpobSO
L2HlxvgA50VnGxgBYuhWeJExRh61T73t/JgpO1sMtIYU0OEkuABQqRU/Hh+7SC8j
rpGtO2+7KPcx5yN++NPnfy8I82XbHHlZvTfvXvOo379XupyiQpR6oc4atjkq1kuO
xML3hKsQNSKSnqa1SpWVJDl0SM2ACIizQJp7otbT0pwUx2X8RkiS/dU7JjdTPCix
lf5OpkcBN40G4e4u6cUhY5f5JMc+3llW1OMn/Y5U9t5BXHMMG+T8A48+s48rxmb4
FE3kNq5JDXOhjnBpTSS65pS2fTW+zYWZJDzWLBjyk0czAjwMrEGHVW0d8x/fCZU/
ulhBmgD4eE8lWaI9aSHVRXC/mLZrJH8EHHQ8c5BYMM49L8Dz3QpbIaERI6GFQ1r1
tYM23yKh5CM2zdnse9yzOR3lQqOFH3R5ksP9NZkp9iR4c6Or4TuBXA/lvTRlsfKC
/jR4a4RQLbzpHQlEWFg57klMelgxN4siD/Ue2yq26Zd4cwZhdUWGhHcnHuvYzKws
zgkga8zpcJZmE02DWBmloYvKQCXB300gllSxbOeawgAlQA727vSFZm2q58w7Q3kH
xNMYeIz5rEjxXKT5XSv2ONRkIy/9YMJmghaKhs1aYHHr6sWQECW16RbnCOmoGgUi
rIe17hko1i3ue4FiUIkU8j7f1VJ1NqS/WLqwSUBhbd+waIAmS+OhD5uloX4bRFN1
1mFcoeMOtAE4uwckgaRP8LfDwbGc+9+Cuq1qvWa3b/ww1pMnjkUMyiM4ZBlEJg9e
9OMN9eR2fI5Yx87CQI7/MhuRxJvtaaWAEf43/PTdGWElMB8fUg86TdD9CIa1Gdk8
381QwHFcqxOKPXDwUMw/BClKYNfxv4UNEUZs0PiCNe5tS70+cY5FjFMmY6N0PJ45
H09ot+ookKQfntbhJC05L7AG59atea/FD966lTjQB63TJAETR1uS4jlSVv94a1B6
Jftkvod4Lxogs/wnoll8h0cFAjmIFH6U3i8VHqCCoPhfqGJPs6P7y2IOyCx60tOU
+psssTfeoefyR6BiGWk0EKdamvdYXVMiLY9i4KbAxauWhdnySP4fKHlt6BNulRfB
D2ZUmNZbISalqY3OZR6uatChSBpKYq3G6VCmuOyjGvMGVVJmjnnNAwK+SY+pz1zs
e7/bI3PxJlKHmibaLvKyqrxlL9tu390rtvoJzBKlMV9SjG5klc+CzEivzEOJ01x4
Y2ujkOKRzm8I48xgwy5SBO/TDoXgLkw+rxxCseF1soFMyWwNqbPPG1bfYjGBeHgj
62PLZgFjo3YAgZNeVQVU4yG2mA1sdhauH+8Q8b8eHp5wSdOKqWTMV5QaxJYLMLQm
MFshSt6omxPbBX+IDoAtPfAE34/4yObx0JaaukGhHQyWESGssGGVG8Y2AeFCGyBV
u7seELP+o6Ar1nCHMS9eTFv7y/IntQ5toHURKoqTl8mcPJ6JGmwVxb1WnNOYzz8v
MubDB+5Cfy+DOF4etHfp1jLtr5yHDZNePwnRs8bVXybfxowhN6y1N3oGUrWZ+bg8
LLC7/rCbNyoconvDmO47JMXYLuYqjqs+tpCdM2dEJF22s1QVADEMjEt28cmYZTFS
3i/KMOQ+67Dzfc+d4d/pSCYASAgm4lnh4TOHBFBIcyCiLcgZGndDDanX/B62Y3Zm
ZplszA3lODwa5XUqoGdRN5aqvxs/i0CyaGCx/tz2v5rveX8PsgjVOaWcoD7HyN+v
zptbCWfX+u7KxTLrjhhpRd49JvdNYICnJmdYzAtCLOVsPPu0U/5WJ9pAf0mPMqxu
beeruAsvia5EjFMXTlFdP1HcMrGYxKMX1NIp8r+Wtf7JeAvJU/dRDqmbaeLBMplz
6h9GEXiSpg3ksRlsBPThrFsbQ4w1eG5BIRBP7SyL2nVBFHjKQVK4+9q8F0ZYkp/W
mDEP4m/GeqJcjhY2QRe7wVWAm/Re4I+bd/7tvq45N9o7cWrih/1gL74LSiGlHTgK
JfRa6AtPAXO750Mt6iK+KKef+lFpoQi4Pgcjln/p/40/BQB8q+NW/VDZoM4HmKRI
gCSMnmpXU+SuhXVCQdVrLXKxbWDWximL4jRghiF6z3PrYg5+u85TQy/XN5AV3L3J
iSdOEJy9W02jGP0mAJZ/jA8j7i0KzJAzpWUCH4k6pKa86bCdZLNR+70v/jIxIE+n
sK/GIcPXG5/iy1aJDWilC2ZHuvZv2LHiWLGXJ/pGpW4see+rMr/SeKLzQdnQ/GST
qONJ80A7PgUPxHMFK0Fv1eDrgpy7PWq67SWOg/r/c2jOquL3YzcKp1J8PT20V7SW
64CAvxfF4yaHi62BKfhytyHPccU0ZRzoABs9S3rwZeUMv+qeSRwLGI//oZD+fgd/
zz8UavpmI7L1EfMuQCJNP1wDQUm5MVBsaiQP2m94qp3r7aGqzuhrzh2XIWy7U/qQ
o9HjMqFDY4xqBWVOVt79/m0ukP6fw7d2dxy+wG+ptTmznaQcfH/9NIXVRKSHy8FT
IS+9utWrVPZl1Rfs5LnpZ0uNMqOEJfisn+Iqe7Juth9r/lpwIMRb7CDMTjWnVrwa
Zed4VuuPdRpInFHQtQTcOy7AclnSI7vZWyevwbnkgNEaYICPfsHZvSFqioR9EWw9
hYOYBai2chyQpfnemK2xxGIz+aprbrz3frEED/LyR5O2/riqy2+MjL01OsDZaj3s
PQjm0d8FUJ3sppu4Sc3pOlnWLuGUkOFLsipO6TgIys4QZjilGgKYicX8tUnmF2jA
osSy60EYtqLwROx/j51o2HM7s8QHIirBmluaTudCLF3910o5mgJlAXR+mPvKgCNA
NHCWWJMVqOftw10eQ5gzczWVdTm+SIv3C5T7u5ht1Dw0UzWt6NlYgSmEauxfkZmh
4c79YqoMQCkcJYuTye12K7O5WqaQ8FVnQFqo9a860r+bv6jV1JAe37zjjZFphhzs
WiuG9htYNCFsX9/ubae+Qi3yreHO8Onewli19gKOVgFfSYF1KJOmk1+DFZJYQA4L
Rdqd3T6STHLlN0y7F0wHSrc3ReELaSDMkxRZqmBZGSbDvlDaVSgAXi4XfMxmDNzV
KRrMc0Ptr8DISPq9TE41mZiBx6L6MQigKsnjSY+085VDisui2vvKb1N54x++J1/3
T5+69D8U/+MQEr2EC11i7NQEqVbad9so3rHI2HKIOaP1AdtFKoUZWacGeEiirpYi
TG7S4jNV24d1TAiRmh/EtursVSxfxYoOSh7EP7iiCjO25RskLUdFtATb7sw/sFRB
YcJTrfs6aeb4GqHEwtT2MjFQ2JdN2a1Lnyfcve5eCsemcD5Z83L+6yYcuAs5N5J0
z1jR2isdL3fzgdZc/FZM46nLET0y+8vvbzBq49+H94R8K9maT7S3msX+P2viHIq3
E51zFuntN1GjRTPaklTlyTkWv7wIKViLPYIxTZZ1pQs6K/KWwuS+whoavOUUALLP
ec/LBrECJ/3uUgwIGF40NzUP16UXNUzbiZxZkBZMML6bvmYepyhwu99FgG78oWkQ
UWskYrcm5yNgbuuML7pIkdCFpHRdnZFLK7FbvPDniT12t/5dTgIyY+2bUXeVNi/v
UQ+I6saqWP27TgNvK2gpQLGmAhuhYL8I6f2efBOntXqN3q3Pxbv+dcmxNmNbks8K
/xkryFfBe4GHpxEqATN4niKS6JPwvnqDqdKouFehNUCagXlXPXIlCJ3oyYECXphq
sW1RcHWg9eEqX8+3Hggu2EYFgrus9JYrCOu4t4ft67HnCQ2raAZgoJ173aEhsDA5
yYraSXxZKzhAdnfmVWcBVDh/ULSXfRoZqs9Wtw7ywRkqSB0/RAI9sTJL9DtSpZEV
AXOuXWScqoLHj2usNH0ipw6ID/xAOra6pbedePFXdPZRgAufRS5MY3SG77MmJzXe
SADtQKNmj7g/X4vGM8MUho2AgyxzAVGHziCqXlr9IkJ8/MXczDqx0PG70DFSEOXt
Ig8q8wGKDe2VCZlxscmY+vsXvSixDS+Lzj3JaSrszgdCqiGQn9f9LtpyiPcnlLLH
TI8o/7+AYMUzF/uWsyiRO8kq1oSgbYDBmmXltGZ8k0CR7yeMM+nNniWDZMVDM2Xp
34GNyGJ3rdCY3HmPwGGEdiY9d7l5LJWOZO5EleOLLZc4DQnRbm6zotUR7Yd9oGp3
mDxgSrjMwxY+0GEsYRURlF1XGEi4k0JA3yu5Jv0TCiyRWrgC3Rfeho6ucAJkVPRE
MgxNmgjNgvdlJPbXd/D3zKrf5dpIrTB3oRlWJ0nAL7UTXbj0VuHniRLghl0tztv5
dgaLAGa1+/V3amaBewRvweRwlDRfi8OOZ/TKPtz4IWRtJikav4/EALtguDUtXq/h
284fhrVUyQOondGt+qMX2hxRYwvPhakVtgwCGgP4cSM2a06eMxeh+4gUXIG5w5Yw
+UKY8WUSdp153yxpR3hPVB7KTdQPG/PuiH/D/r9c9AqlS1lWtyvmuuBgyORx07kG
Be0Ah2XlQ1wvnkRa9zQdDBwzx2Zh7AOldsKluxCude6QM39AiGMfySAaYlkO6YWa
7dvTyiMc7akhNUhEE2ozxCxUPNrLzDz7SrAHCoZiCAiHgZAurrLGbLTQZPqPxLi6
E3cedCjaIlg6UYkeGTGEYpgH9NwnvuKea5nX07/17gV8KA/Zopb1KDy4/IIrgaAI
oyup8hvwdE1MzUYEH5kirPw6NoDXyvBGzaNZQBcCRPnS2P5fY1lobjYFPaFwAxbK
R2oTkQr91UE6B6lxMBPlIPKAwIIMVUbhzrqoLitMnCsCtfBwYulDZmCDtmR22M2T
1DWAQrHxpXhPed674t5QySP5quT2Rt8xXEpDTPScUUY7U8IUDmao4BtaNxcDnTzn
vSiIiZ4bGYmRL6Wg8ZcWEdlCEvPmgwLsBV/lNSIRS1Oj7tpy67V+rybowqQmmeSO
9fnszMJDgAn19jNxDtNUN8m9aJrQWpvSNQEb4+0LPNkBh41RsIBBJ1Q333LdX4/O
i3gD7Usk5wWw9DhLmjS+LkFxZiBZDifzCDxpYlwIjy03qfypOosE2AxnQMk04dM2
VIW1nYjTLWFOZzM81i6yd6JXu8mcnahQSdThT8iUTJYjgu8DWf4zblxKYJySdWCY
NiuaIKvtO4pDqeYG4HqGTH46CNJ7W8h+F3P7sXM8mWP0amSCtScaRkBl1hi/v1Fs
4JlEc43xTE4zZ7me0y+Txo6EudZqyckIUEVNAO/TKpqtHKJadmHonqBlto+SADrs
NSQEr0Bk2hhdnWn6ma69DN2gD2b/MjnWlTKsKRPEHrgzTNUGwByjjXN8ROFAhh87
GZBT1E/qrM5BBKrbyFhmxqtdOveTP28Q8BC4j2MSB1DMr4Xfn1I4iW8HQFS2a8E+
sY3jXHKdE9E1IQ+VN+6mQxLD74hxrIhHThvN0JcgXt8IqkUUx6KEsrZ2nb9dmf5W
JsbCFeQfAbXPAixOqsmGzI1WAuKGLODlucnGZm/yOkycoNTCh7IH0Y6sDKzG3R7g
WSSlEA+JjM4TuTrUIF35C5yhN9CQumQm/Po7lNxQXlnG9060vlfHJRbVEPAHwzWO
HiA8o/qKt7ZwrrK2OHUjKjk59Tf/es4OFsiaAASH1twIY3LJgeLgVQm+TkHyGiUm
CYh8dX/2Re4HbUzIsbM7nAQCM3//DSZ8hwUNQ6QJQ3t0HvaYgU6RV9Ubm1jMIs0T
CGMRcxe0Vr6oLDNsPNSu3J4tu+MQnNPI10FCR4QCa75SPmVkwMFJQphWyxfSczvE
mkzEwTEBxCSxjqnctC3KuNX5jD+oJRHOmeDbTNnFvRTQUfoAS/k2WyWZKVLB6LX/
klMSi/5su+vJ9AVWPJ7rPSNCGVM1oQXT1ZLM/YFn1HkOyT3lV4IGdNZ20Sj+7mEC
xpBlDJEGP7/kgHQCyLDUJHmVPu6XK/jZKNcQ7S9dblVBgmLJEjJGlT+JkVJWsTAM
3g85UMOebqVB9jActrBBcEQQYLtFQGGCFjUM9B7Lc95tk0knytpa7ixt6lvjBdja
THvhv9GXZaULzGqHf9kVDdmY0Ic76yJS/dLa046grpSi2PPsdUUxS3nznN9nX/Jb
OB+rRtzFL3yMJOaDYHl4Z30n17PNVaotjm5s4Hsucdh8Gbsz5IiLAzEF24sSXHOt
k7ZiQG0CzG9Q+e/7ymjjedyH0l+Xf0/9SPS43LDc/3v5F248R3AMgUCqgaU2xYap
bYh6EFIimbJKW9UOvAJ6JnZh30L87sOT5VLpX3NaWt9A4ZCheIEQtrEHMqKW+fBW
80Z8Jq8bNbR/fYxOl1n24auN8lAbI21WHKdGi1yQX6KuE14SYuE3+Xz+2UdbUF+D
XkL4skSs/Y4t0jpOIh+iCjnUwJojCTk9TSMTs3AbvmNECYcOSX/wmGRAsykvXLsF
z0b40eA5gLTQM7wMCwUYmBcAmNGEKvLn7yCsb7tyxKjU9T4IGLhLfI8Lhx00M3Dr
EP6EFWuL5bcfvh41K7ltq0iKmDLL3k1//9/QT+IxFz4mOocNUEuCZMjqMYuChI1j
NQYmsMne+vdPnX+pOJ0A7ICoaRvMsZlEQSSJQtV/n6IeTbuJOD2Pl3P2gdjxrTXC
ke42rkJ1DEUiSOCFyTPyVlSpCcoNXRjFlZr2do6EXDoi2rIP+43W0L+KIhIoEpGD
y7coATKYsPPpYRZdh+XoucTjVoLtFVlwdpB69wtFxIoC5f6sA+POg3GwiPQYnWeM
lpQko9m5usVtpoNZHoHyUwnkXtPcqrD8k1Bi/CkSHBtdgISgicD09f8mXA8YnLyz
kCCZAUx11vb4CnC38zhkfreurYiNgAgPzOcdqSviAFCS0k35RxsCYK1kxnkgzOsU
mwOKc+0IbW9S2uJ3sSDM49tV7A8md65bE1yR3oiIayHkZLdMk8MOwqMntd02g3X3
Dl3PBxwWkPzye/DLWy+BOFBzqsLsrAqn1v6CEU6qHjhOjxDiuIjfRcf4YBR1VDgd
+s5dtUrTDqobkQu63RsK4QqTbFUYpkMdxojizevLTxaO9Wn1+CVEt3TiJRm2ImWz
8IqISifeUIfu3pNLgje+4hhcoaHb+wdhuLOrrJB70tHxyMlWUs/mZVj0fRJ4J2BC
LRsMX4RshuHw6ALmTddruT8KMtFUrWbvr9wrK8IrMZREGvnqXkcvgGyeyua+A7Wm
O9BR32XDfHEe53GDwWlqAjqJ6pLg/u75zVPU0WET8oLYhFSG/qBtkTogZnHhYiMO
njiKwcS+BneBEsvIfDjphpWIbT3hJRBy4tU+jHMCSXh2LBrhOPTfdrdqQkDs4yoq
JwlQ5IVEydW8xDfg5VEuvon/HBzu2rkTsibiPJkqRJl13/JVJ6zkg2G+5NHOB/NL
qYL7j50+ATNXwiODtQCIJUy6Lsevd/ejmyc9idJSRqxU3ps9ia+jkmVqgN5suVLl
bBAkwgtjsqZaO986/Aa80ZmhUhpiu6DecEoAjpxzvpm0WaxElCVoPynV2wyvuF82
d19mC2R54IRs4UTHi/sTyr2CQd2IdHG4CCg4rJGxexPj9vXlnBW0KtukdfSBd+58
TvQ1mD6LaMLKvkxpnnzhYEBETheoCVnrYv2nafSN8RipfSottharh9GfyXWb/Jst
gurFd818ENTYZ4eh1000Yu3Uj5kGWn/VNB5mHMPrMuUDM0mGPL1u51/vyha/vE4T
NPMJnqfUi4c99WYhMjV68xan6sKjIHxa2g3Z+9NBwTONIBVu/heWxSyyjaCZR/r0
Dgozl2uJ0/D1n+TieWlFHFnvv4LdyYnfEfJJPG57jA5/1upEz2IifO6ohzXwHqhK
BdDc4mOpVt5gCUtN+7h7KKsj+ZD/z8e+rOARVaj6I1/i+SGrv5p8BslFx9MInApZ
xHlsan+cVS86k1M2F0KjXnOUyrf0s9w9lXNacTrYc24L0Sdt6huRz4Ks9ovOLK6B
5YHhEj66wAVyg9/6q7M4NfBc6YkY7A0puLYXKvE0AyaCnSbZxPn0Q+5tsEDeGc4R
1HVBUNKJAUbCywPuK2lW829yuYqq/Ub2sfQ8kvu65IzPhQa6nMhjkE30mdazFBVu
k8gEAwIkrgCBKjkg94vi5x66u/39PqgPESHvBQvq5uTFoJwEYmV5BiNRzKP/Jz6n
AIFmu7E/nnzMqmJRON5qWwHRlrHgCGMgyiOD8qgiamKd2+iWZe2iOn7r8yIU5lJ2
BgYZtpMTqzZuNRw/Eff/F24O8IFBgRCJWJAsR2MPe6cu3DffSrnW3UWyI291I7bU
YpztRESGM6qNtxl47Ck2KdWc6Bjzu1gFdB915lXfRIaKN+ElniILhjA36utisxn9
6qQxCr4WYDEWKzgaNocPWCYdvvWO7XGyk1aSA5jNoEOvvLdKyrqAMbG8noo5EqXX
FutCmSnRcndqtSHM8YUOsRNISaYichkX2rbpgLj7rfu45XWt2b7F7arYIhCi30jS
6onwH18towt18S/690cWx6UFthWq54JEAu380mltH325QEXbZ45zgmOwadzPJPnc
eYVjUvSPmcaoOVU2ek8oGSNvpD/v/iJMn6YiBSTl6W+QO9fIlKiG+k4EUXL+eJHB
aTKN6gZP+KQtlQTyj77V+Bfr/0u1XqG1Nk8POVCk+J+VNji1Ps7tfISduBHHLs29
Dj3K5T5hRdmiB9UTq9U1ZykaQpXV3Ju9hTWRXVQmwhvADhLEkWOxWUNekrWvEohx
DjgxUCZRoY/7rpR/u1C7iKDusepcIi+jlRySzouN1JQ0tWuiwx9d54qO5hn5cuTZ
R/xptN5mCrBZCerr5/hV14irtklYY+pKLSAx6+J8ajguBF4n/iwQ4kT+X4Pd6uqs
5q4PvLIGTehDvBxwqz0rSaP5lex8P9598z0dBxRd6Vv3JvhkGrXjLa34FEw/qKv+
7NinP87vTRD1UbSmCva/8aU/fRAiI7GgZAhYAjGGYNeceMiASr3N1QXrDjpBq7BI
84Mx0xBKtIMDCpsiSn3fT+q0ooPRABL3tD8RdXdivEUegPBGpGCUGwJoiq7YXCFq
NunvxQo/YY8tHYtUbxEnnWjA6k+S9Dy5YqpZeSTq06jIyOMMyBwuxI+Cg2RS/KIX
/LqozWvopWic3sNnfpmFWi/IXBlf7wl84BkxBa563yPMgbcAfoWP3SzgFtJvfL/S
YZZBzfd3eljBjIHBU4UD5sehPIrSGfoZFHa5tA92u16R2QyBMZRf93+4f0g8paUp
CSxWjnBp+ZR/PQjx6/+kG8ER1LVlrMDxgKwf1X0J+hsiyW1asqdRSB+Qb0mjS5T/
sIoSepjsX/Ao2317VhqcXkAVnLVUDQ82Q47pqCCcxxn33yyUsoWUAq9xjyMH0+M7
h6OqjPnzqbuVHYFs7AdaysEJNGtAofIKf487UuYwvCRZ2wz8+l6McvPjcMdHpBtD
Wgw+gpOQNrlX2Jb8obj2SbVGhLNhdvc1bLpNCIfoMoHM1k4a0WRHMHXe7qcMAfSv
gurkxdlqHldq2C3o2ME6VNypPib7NIBaAXu1V3t0HjuzoEHXqb/W7WJUiSL3HgbF
X/YFo6MfNlVRb99LJgdfLBN357xdA2oNMlMZnVWO0H7cAR+CWc+OtXrvmr6kSf1c
RqxsuWY2UhWZddSRmuJAMHexxYxXn4+YYVpusMQtuLlsRVkDqexefOFO2KX9u7KB
bGMaFHMKtlqDB7xJWeDQ0LmQNA089HPgVrWqE2l1E0M0cyOenyOnDte3wsgy54z9
eWxydnMyzECIET/8Fg2ZVHEp6trnnHD0WD6GoHXrtt43tmuZqVA+VIai/j6pZmgF
C0Rln4gskLUDGbj8NM6+c+SwhKCx7+W7V+YwWi75jbYPC7tpsodHFGtg0x6a2jAX
60x1lTqho70Qn6S/un9WKGlfU+6BccifRGxvm7I0tO3nVTSekexos1hY8GMh59uw
+1Kd1MMzaf2mil7NSCcmBTdE3kH0Xcz3fHVAZ5e7e1KRsrVXzzGfaPrHOKfV0IA7
ndTjBr2Ps+I3IGMQarknjfaGIDLG/2sfEM2CO1/Cevu7x1Fxg93DuJk//u+ZcoOQ
YyKQCKDd7n4MIabTjPGuD/Vv596ni/WA6G2z9+WdZo7lVDLkhCqkH8eGv89DY1ha
yeiN2fCXNuDSae8z2iUy9AyfnaDCrhZLTXjxpHPdT4xVwhGaIPSxBvzLMzssHI1G
eMpyg4uIbn/EpOI2w5xaa0VaUv36rGipwcfjvj0VVnjAE6IbZoqqYe3xblO77fdj
nxw4gXIXqQseTcWwxeeA6ulNCOQCvQvllZpXpqj63nmOLvyYJHatjiYazYb2Dd6s
ngr8XJBjQtiWVnINVdKPz5d3QTxP6lwIUM0pGHSzGcdu5JSy/8IBOhy+LJJ8lQWL
ClSe+SFZGtMbXto+MB/LajXzegg01Om/Tcj5CdA1VI+ii3m+UHzkJsEHJlJthJGP
fZVaO1iceMzbiCwyRBUx9QNVh6xgRfP9j721hD07/rqD9/MGbMlOEM5S485UJqyy
8Vp4dn7V5WEv9UwMJYeOSaOnhUJd/+bxIgU9KHrV+SdzJICSANc4taFUrEeCAPb+
PQKLpDwXKYmm0sRUbDTkSyf4X0D9bJlas/olMTA/W9IUTdAVEjCcG1zOCiBh0v9O
rMVKw/IO/x/LDedw/zOogsKDONVqaz7LAYGW2dfA1cXRQbuHqtMcqi9Nbum0y3xN
48GmqXpb4oBOF9a/7HlX2fhpiSKwjBAIOj0Kym/GBhQCIzBtOuvaC7+Vd3oBys4I
SPjnSK7q25Mw/m16s428B9aWLEFxpuhMaeIeoKetJ23ouH+Hx0+ZOdAmueE8ndfI
LEXGTf3Vpi/z5cNdWm4Nr4ztdOV+OISORlzrp5WgdVZYANAYfzNULHRkHhTVMOZf
ggwV5dsmObIXRD1XXentWGNr8pnALEX2YgXcv2WlBQ8J7mp/RJPEkWhraHqxcq8N
ZPJRtJDTjRzwAK6RgODs7Nne40PQra9IGMINzOngilh8dcA6h7ZZ95ycLmpmmow9
66IpoM6I6Jh45YFCyThzFUgUzROnIP0onjvhV80RJRQZJLGH9U/xdZDqMo20y+gb
d/PNxFq5k+Zhp4tDWzFqYZSvMuNynRmyDC4b/GajckKDmhC32fgQzyJwTntHYN3U
QyOkyDGqtBS/E259t7V356C/ZU0d6SouC6kWaUT3waCudz9iMG0+iDH6PsgOp5Bu
mfKm6OfWlYRrku2xCIGmlqxaBUBM1W7rmGNIaa8Kh2HYXHdMmYpBwHmBqsm53XIj
k7tro8ngMhiiiGFvIuJFlsqcQKGBZu/LMpicoHT8sVMLhkO2GUtAT3uqgiJWalAj
Du1zSVQmOJub/Gv+daVFFSgJvd3vbr8mVw7SrAz/Q6XBSfUam+RMXRet/Mvn/K5E
x5sCYT7f1ofHnj4A7Iw5clta+dAFw3J0nfkEcmej2yxt3AXwStWKbhSvptmlsUAi
9FMXzin0mdZqW86CBksnh6ZJusiSMzGaCEqAzGkCxDAxW7RCsrJeM/4m34n7BNfK
nMwjeb4OioWRPNCyOR5qaUzhamjhg0KPm1GZPdE5R+ibZfaHHLV5ynR9yJNLjxvw
+iFRWY8Dp6AloszuXeIol4ipx3gYQgeyQr6G0JE/KRcvyki6Mp7HwWSE6PVIOks/
NotiS4wVy7MMFANasfwED4F7NiHVLgwllbvSAkMjgpHCFxh6SOWQRX0VbmVhzdm0
b1qfYvbTw+wzZm9zKWvxjaXeE7XxVTmqV1+uVEqsjWqOxKk34QX7tYsuwv6fTStj
ZwcR+3tTt8t+/x9O+R/GwfGPh7/001P01bvVTLKqmOZxkrTrMsvC1EytXqpYk+P5
YahBCDw6OkTsTGIsZXfMoE29T7sXXfMwo5hS/w6yR0Gx/eA66/PMYLpm1Tk1KDtl
FJC3uIHZkD3Wrw0aIUfWvPYaVDIMe+npPvIIQI0TKKCpEaOsm0Wi1MRMiddXefiH
XSA5vaR083WnwA1PNSIO94wUAcJLCtqlMhIbRh4oHcCj7rpTkQ7Mpo0p5i7YdDvu
5JV21gJvC4ZiwL08FhPfjEz2KPifMcsFmg5W5OtIPK75OUWackV7UXnzrosJyYhm
3u+SbFJIthw9i78DLMwY3Qtn5KaTzjSiaAij2oVKwYdfy3mm3F9vbH6Xi42CGk0j
7nTRvzf8p74j2viXX1ipLOxj9ctWtQi82K9vJsf7MmBOUlESPnWWMxQ8OaDmCEVv
DUo6qP8JzQWMeuoIhWSwN3xyPa+nkgnKhmTV/uW2QIEg2Mjg57jKLt8y6Lo68sLZ
fJkinX7s56Q1AsCtWk1EDH/POygjXt4ts/ghvC+p+DT6E/KNxVvIU9xkbCf2SKQ7
N1Aa2/kFqg5uj+wUnAZrFKKobPFV25MO7QHDSocxHY4+wQHuqoM7/P1WPPsDbA6v
YWmpVsujyESYYZfBj2ulqJZTZC/udXDo+d/Ol1niKL2OSPHy6UFWTqGfMWo2u7Ri
viC5BCZxbNpzuS/oprlX4g/9K8IuFBEygUrwgZaSNc96RxHu5FyV8uclqOaJ5PJu
cRCrApR/WminVtWreZ4GlGwSm4C4vLdbl+JCCrN3CR3Az5qqbkDVsDhtaoDsP3lu
QgLs5hZ6OiMp14N7dgDqSIdAiK1WXv+hWL1ZqzAOxfrBWyHm5VYSKSqkyFEJgIU4
MRLKJHeBvatmKwMVTdjlD8kCzhL3u0q7tJvCfJSyCENBnxZ1J6ljfiwDY9+pH8rn
0mBahNJx/sRqcuzp4Azy4ZG58SSig5TLCPkV+7BHyhZeyIutSmyKdxqiBC7ysxri
hgneSItou2DSQUFfCaR4UOZNBkuXmctApo1rPMXuxJLiCO5ftb/ax6ntlnSex/+3
I0cjd5XKHfRRZY5VQVmn3q7xylFBbaDdI/8CBXhcaOIK0VBG+mPzavBIY4Wjc3wU
yhThjpoAJ7SzjyZ0MsJ9nWfTojQqSU0VVqPA0/xglte/popeq3OfGwuH8tNoj/0S
w+qP4cvov56BB3RxBYKnTOJbHe4+kOcyXC0QsmNb+MBA6+H4PoIIFwznLA+tsArF
011uPqe72mLCoGTemgb12vh1JOpLRIsTgm2apk8JQu55nBYeZD1eYk9aH3fxFD6p
Cf+eSt0HOxFu22ybz+KQzxtl2O4ERp7BOyHe/u7eJIZnILqxDh2YTBvvAfVroR+O
g8ypccvEuzm/s4QMviEJba8+z5BeS7OffqLBRMD+swhAGZQpjlnvp0/MFkASn6Da
d/EFH8t3kcbqC5oA+dnfIXHA/gvp7eh2lyq8i5zoT6dQ52cszmvCg1kzWgOaccTE
Ens8OoEFsDcJRqgNTlBWx40SafzkgcA/Yqdv+sFgkluhg88FcpNJjGTb8cgNojTh
4LmmwZWTgaE4wvnG9/kjUbk4Hbve23pZvpswra7+OcgJEWDBl8+27RNhexGqK5r3
GKyiUezK46XSVP9bGEGpEjGlidDLrco7dIyEmOmwk4OlHvAqZNu/KhTlZpPTfl17
E0hhmzI4HqCTnoSdpZzXVx0znz8nxBr2PyYG+i1dtn7OQyLkksqeJ9EKmVQpaCZK
HYp9YjAOvaNWs7fAQbIalfOodrU5R3YSIUcEVnFhAvY1Tu5E/JTJuMAklbKbr3VN
pJaoyWQUVhGGxrV4I14+HdWE12DxJ/QBzWcV7rqd3/cXrfetrL9NGyBijxI7+8xY
/+XVom25JSAZtwwWDwu5z1mc4AnTsInfWzEG2AXdB5eHgcm3y/7sjdB+Y88I4LcV
Diw++MQj/4tyDmK4KFakXunmJBpV6/bAOI6l9hy7Mv4kcxX4WmZjmP8bDSTTjurA
ZuslgiXhIm4uCVfK6FaecZqFhaSrcG/XBH8Z9a838Y6aszE+dgqv7BIG+zBRoW/P
472SZGs0yikETSnYqYZYY08y0fDyzdqpLNppSQxfxoefXtTNZOhPfgaiGwNvPthE
PTR7OCi4aNR+OYDgTah2YV5/FO9+uyfkUU8rnstd5IPn3ZrULsSGNPOx8bi3ZzRC
8T3MsZeQucdcgEEKM3UjR3LyPSnv2cUXSfTnbU0rVnlQZ1ssY9Ilx7TmjgmM127K
SgN2SPWDHbva1o424dEzxwARUVhLYG/Qjy4QcG6BXex+Xy4as86ONYDdOlsLvJjC
fai02TXZsxw7ya1b7LQfXpsbKwEkocAzxDXwHMbixOZhiY3a8B9GKkGhrydSGT3o
F8sIMR8/1KfxsCbEmi4nEy/4HwBOBiSWyzce57EHjU1QCrFkTLRCh6bW8slcB+Wp
DyJpSf8Ee35qDODLZFfBa/y+qAYC8/WI5jTbcG1ldbiWrwa5dySAeVaB1/Tyo/pZ
dMJA5lb31tWWg1xuLktT5BHhghjVW8SdXkokmZw0A5BzgO6Yn53Q1wOo8tb7yGrL
jLXocBkMh0XCCLRYhOF0ZHF0w7lOteGXI4SM7YDXkclZarNMZbPfzEpnTsa8evi6
0aCxwcud2F/whO5CoI1VJGgAJmpXUAQrhzakJm/0X2tCtNeF+cShWPwvpaO7DYYB
yMSM9oZ7Kado6ulIvNsEW4SLBWX3CzIUNNIcOMGhIvMHe9LL5x2CK/8XWzeTCTnk
xVsascbM2ISj7EnjtZK7PsaNzlEbLjqdkxFC8j6YZtHhdmwT5vatTW83OkU/YHfz
y92wMX3YibVld9ajAg+njjiX1+y4B3pOFw/MCQDUdijigjkDOUgQOuHebC6RTJlK
7OCJkosQIXBG5iF4eAXJ3EY1OmgZXyt4JLFDT/OJrEzD/WoELdH5LQKqXX6JB1Uc
HZ+n5GTgBsdAhQ8rdpCPrpzobmH5ysgmfGdHyhibSMdkkGXHCdo5nu6L/t5MtJwC
6eas42kuJwWDGQ/AZXI0PMvSN3S9jb/RVFEtFXlA/ujQq5TtJXk/2bgzFdEp9Qj5
PxSbVVomtAafViHirl1EkpJ5S2V+HQFeUpXyrfa2wgutw2c7exVnzMNG+acubtQz
pNjqsfSHMWUabNEUInjg/Ek/UsZDyiSkIx0+2egQN+V1On5FaLGw0zCIrN5ucC4W
KnFoSNXiItKCsk5KmsDdcHpME3rqjjxFsAbU00B6/Mnya4FN9NqCeUaw08mb/cid
18fznkyUGohJCODeYQFwKtznfZuYgjwWlJDNCodDF+OBwHcT30ppewV3XN3HA3Cf
xlQCMgZdrXUdPxuTsbQeO+cO4tsHMhN2eylTD1VRyI3jcPf13cLWNwRzCDc615ug
gYrA+gCZvzoTncCDkefdDgBgfU0tNFrlgD9uGdQj42jfrfaMMday4geY5qtgJBEo
ioOelHmoh7ojdDy9Ijn4hYBuHnkCc6cYczD8v839USGlfyaIp4QPkc+mz36B17kn
UaLM7jPIlQ486enEQEdNtI8Ix81il3+sA9/RpA9i/ANkX9Uea8g7DVbfSM7kL+GI
jgmXR9sXhby9QUKh74MX/7fdc6UpQCOhZVZuJCzY/vkqJA6mUfK3O1w3wYcEXFQT
676QZ1hul6s8SIn1IMXiMQhnhUmoyW9NdWKeFF4ovK7CLhva/bn3xISFvTRuc0sv
P7QGksmVrpq4gt341ZXU7Bja5iq1lE8yK2x52ZTtPONPPGAnoaHs2PimJ8RwyFHx
/5+9NpBxnuXoax3zd+PjxyuT60mUZdYAMv6qJKDLGzTeuC29nA5NPcr5dsnqjK1J
Tr5ODohWGDbp6y8rh5qhTXhBg+8Qx+5j5Bp+awQ0Dn8AUXWysHm1AXWLZaWdLZeu
2BQXrPaqng6Za2g8Hq/C3KmzI6qBTQgTiA8yj5ZPk/E2WRPdejTU4koI5q+GYPHx
1JKz7LQhjM+4mLdxAJJpzqfaDBmBDzlORYrSIW/YzGL0Wv2o6f1Z2Eiuq/gtexJ3
uwC8dZgsJN1jsw01TmXhgAM6xGcLLXyrzBBofVIYZXPAJXPT8Gbjd/KeINWuc2zw
OmLXuJuTKL7/Ogkf9GuPD/Tlk84Koc8PZM4byKYR2rnC/Bks+Yf3L1QC1pYc+pae
P9oLsz6nwQPrgKC8XU/CwCyoVYIn6G8xHmOx0V2oSkR2fVFFQj+5Guoc8ROHRMBE
VHyYVYk+kbRTE9ZsWuRHWYe0NdbLPhnZxd4qDOxnVTWtVEuFpkh2LDfeeVpn3Dgc
67Hsk9zbQuLF9nEzuMQlKIiga5obnu6tk1idzvKsUnGk2VibjIZ/L+G8PudND87Z
N3diKt2A3hPcHu5s+lRThh82s8+b3+kkN33PNTBzM0YKQUCx27UjgDZPFHagcwW4
DhFo57d5b3/J8+xucpLWtLFEc2/C6cgbRYXcrQlUrg06piok4TRubwZTbrmk47Ys
gb01NdgIjgqElfdwEsg3x2tvDkCslsvFZzPJsx1RvxNKJ5AOKQrLHpiE2Gk+JvFQ
xcVMxvyrVHmE4mtIwaPsjzcebz41u871+brATwfyGt5AmCmXA2eau4Zlxi8c+FZB
EGLpviv6fpSZtwhfXpW0dTfxR9+qb2EaXCOUbbUdK2ZzRNc2nDUFbTRt+bfEZygo
MJ/FYFnvL7M8ZcAg25sM/4gZb7UQi8fPWcp42UQONutFO6yfSVXGeNNNBGbq+bxO
xkgAabU6qryDz28Bw2T6lF0kZXsFlGGE7Odn8axkJulJh+wt/fY9vw85WZHrxGHZ
W5poof3MmM9ygNUc3dkqHhVzpTzk7jEIgngk2xIHrBqmGQT189LkI/GfQljSp6WI
RNYQ0IWp7Tm/mpZqfFKApBEOx5skw7CNdG/W3olnQrCEWhggLu0YO7RD2VfVq60a
bbjST5CDHMQdeZfdgBHZvWLTSOtefT87x1A/Lb8CiaVTGrEGSA9qzbzwj3uVfr98
xoj4IM7u73h0GDt7gdjqABCaXxQ19EqX+OE6TfBTDLxNtEshBg2faVnm/RX2p9OP
FDuWioWqq96XXyWJ3E87dfUFHgcSsCGM0OCRsxIY7T5Sgkmwf7fKkgnWLpDSGr7N
nyW/jDOCtf/fwmQeXJ/bhyDIYyBicaIe5JSvD4iT906mO0Yk8w15DowIFRrUS9Qr
e5awujaGn5EqHegOMPqRvycvh4jY8BHDvViKYK8uBfBmsxEEX8HhL9nehl17gXg9
FeXOdLe/y1JXgr+NQtHVpSngic3nBWgMn8TyoiuDLOWOcJWglzuFPuyOpHP9H0fJ
xNvsuKgN8nmeCXm5EVFTRsJHfqCkhv/QCTnHsN/zg1MiMTCqt9W+0C9ZFBNvOY8l
RoVMBQRA0g7DfFN2C7TI9piK9FTCW3M2gbOXJUbNOZMxAqqo0qiLUGFFj3Eek5xd
XWCcVKNyxwTGhTxpRSZtKm9FWKqdwg0ujb/XJDyxFEyDBXJm9ZDq49+9FmSzxiPL
8uHIrKBVTyKZ6m8HJytNLRJVqtn8C1tqOQvOGGGBnl/X0JajuXy/hfZty5o1WtP4
oXyyfFVCdKCa3ij6PsoSds7ttCZr4ceh7anQifW8Zeu068hMnUYEjJuC6srnrVzr
LJBXa+21tpPiE7UbcWRg8y1f8666j9vNAi14GT2TWhnYFlH3hykls3YoG6aYjVKg
QPM1ET/4+4xLOGEYhTZ6O/dpD/N2w/GuRRS+H9iarjjRkiFivjZm0JWZ5GyldyTj
ZDfKLWB/ffcduOP4iIlhAL/OA28ZhBobTjXV29FMO/2+RIAbXBbpsJ20/g0MhEZ+
6x5/OpNO4zldCBaKgPKpmi0sRzqs0xrzh5kZhK+U0d9H9JDo/q5/ROpzg/iRAKxR
3Jt1GyJmkZ3SUDGfix29RpkE1ceuXR6olTOMMsNupWMkXe1fK17/79HKNGuIIrnp
mQ2ZaIUoAUEkGoP7skEsEZxBaXZ9O4trFuB+duOOYBfG8kEL9N3G/v/vOwqTaHrt
Uciem8PHtGutKeXYWsfNLg9aU5XO04BbTP5ps1XIyp9wM9e1ThcSB5L6dYCpHzHZ
OT5Bf/F/ev2AS1vWwnRHQs3QtQeRTGeFYkR7enf+xEKVkJDvAsh/7tf0ZK4WGfCr
FbOCRSwLHJ+tP8O+nwvyNcVcuJoYzXf/ritwDjrR/hoRNZ1SKn6qF7Dc3hRLxS12
QDCz9SCb+Jz2Mus2v2FxQrvP6vWTeKBvNcuIIEAud1dIAEmzcmz5ukDr0lk8s6wS
mpe5xQ7n5jUL1+l1m20eiI6c6nw+601IpTh9kp83ASM7PLG+JVHea1a6dTscUc4D
i41tqlivCianWGeIJLfPiCY7xFq0hYoBfYhuK4dOGVu2HL5dAqarhLHmFn88c85t
NlpadBzfpxYxM25q290rwuO3YuN4s8f0GQTJqEJEN2DovuNBYW4h5/Mw+LNYgG7z
41VnOfOVbNXetPjhqSygF52gg8XgE+Sk5z3rJE+ygmzqWc+Ad6RGInT1SNTODKR/
ckvLiTdoKw6aJpy1kzMs06F6z1z7lI7VW7OycNrJb1YYfccp+lIqhuOzaAyLAQBv
RWarqRB5oO5J0hspd+Q0XZzZPm5y6yC3KvVNCglG3CeSyT38yI/H1cwhGPIZeDfk
BkagOt5LM6ydsaxNZFq6pz4AQEvdxKjdfMwTbRKfAy0TjAXbhsyNHcXj7iT7K4wa
HsyFKIV9j3Hmh3nkd6g79n4AvkhuIEWfOYmLxj6EsSfhi4kaJbaljUpX27Qs2vnt
fQaf3CwPHTyMfQgyFCc4q8xK0ULKlwFbJ2gVH23W41ywKopEQcYfGvJLvRrLrV0X
R8mh1hY7YFINopVGWFPKCKXKfMHYVOpOjLXjvpI59WdvKVUHbV8K1dLneEei34T+
w9VbF27IveOPHvs8q/9FgXe/c+RztdAjKhbcw6ENro78lTbePTUw3AJ8+OCgesAq
IFET3hgZSEb+be8Lr4Kb3maY5pd+JKOTCdNRQkE+YI+UiBW8OK4c1bY4sK6R4q/O
eOgNf9j+ZfSZvmSG2WpV74MEOn7tZDNh3RsFjDm75KiXOTz8ACMpHinMW1NY/AHm
oCM2J0GNHLzXsSnLJnNwZpSK7T+49LF9c1C1HNgqyYrkNS/aZfH6QNoDlb6KNAuM
F1a+zEiMZ62n0B3JZ9Vxp5g3jA1D2LJrneWbFC+iUPK/jAEeIYt8AeFadHiYSHwH
S1AqG3jvtNmmUX7vsPbE0fHsDR9Visu6s91bq9cDPH9CGm63cBDiigzuKF+chQmn
8dbzi03A75lKxoOjgH4snHRWFmepO/n3o1wfJVN2+Zl3aEkacSMDUsEMX+UcjOm1
puex7iTak2t2tMK1f4MnxRh8Hsw2PRs4rvXU7jwsbwluMGnNmPSMVn8GlsF+Ajrf
/kGCu7FYiByFUmr7nZEvNftZcNQ1jLJMis2Sxwe0OOG7kCWjefZaRVsv9idpefx8
mXLu/HercKbCNDVGTLZtYdcngEd8TafRnCavDvSRIRaXSbtiGWrlu6r/kJ6MAzK5
Or3dYsFvplVddOLu3kS3xIxdy1nVVZ0qpokKVwBGRnL0JHCixy1qGgtC9FKKTT8W
3SYAz8ypyLxe7YjtsvfKM1iJDlmFobhfBs4LvvsRnjLm33os64GkQbwMV+JfUThO
WX2V+rkJUo2eopXLVdovlE5ZPiQwAwFd5YJ7SZ5uc+1d4WCtJVp3Ua4icNtqpNvI
dX+n+OTGT23gSprBXb7bSr0wDoHBfefnyO0k0NhRKuzks6m1p0P0h27Yk4QIkPQe
yGsqcB6HopflqyYIbrR6j/PIJCLjPqp+tfqvKfAllNItCVDW4A9103yOtIsoB6Uj
uttyTKVb1doi5PptWQa8lVewC0xjq5hvuSpoQK/1Y5ETyOGmHeni8iV+BaHY2CZA
rC/F9mxa5l9FMCie9TPZ23EwKLJY1u/ePneEPShNEzm74/xheBvNSei5ndmyI/xu
hq5Vhhrh/yGDMwf8gYDJc8EvDLDj2TUt2onWhCg8qomTTKYFUwfov28GNFzLZ4RM
eUT1oU+xjJ6fa88933nTed7XJ9TNdVYZe+JQsqwHCKCcwcautxwtfmD34KnDjPvw
8QUk+OYcwIgDkgrh9osnZuyNqJTCLQzcLqo69BqiIFl1SxWzJsKT52rL0UdEBlA/
2Dz9auV3bCdZGR5wJ40UoK9rfL5KdJZQYBgFIpcJGGX88uArNP8M0jHzXI2UqEh3
H3hg7qgqXLpUjBfHwQxk7FpOnFlHsbeqH2O1UPUuMiE2Rg3enKxy3XPZDdpYEi64
KqWS3xTJj1vDSg/1AlDZ6/+xfnOZsNMMNpIbLl0itvKAFxyGX/DmVxUStiZ5pqUP
N3C9uzYMO+6eCabEjnbyFLK1CB9revuBOyLA+CNlVtKhdbeVHKPoOh2rMREFAzWx
f/nuPzp/Nh8ZhuvKYj4QJsM0kOGgCyFlSV0QNyJoObgECJyU8O9piwSD3Byn3zGO
v/e2FcRv096kd5KtBUHybygpt6/eHpTjIjLMXwmHXKoTrvBYjt05vxwkCl8O0zfS
IGrczakhaG1h66I2bZzQ/RpcwilWIPV64eLJHPiV/wFrPDL9r0N/UsopAZR9Z9B7
SXJXfhNNGTaaIk9MJaurYmeBE+4nlzMffhHkyejjD5smGoGFAFsAjrQaI91UNm4J
0Tz6KCRAwUA+LObUkajTxlpKTMF5IGRDeuiFYpcOiunwTMjzCcorwVmeFLg6uyxR
b6BmTaiSVSI43P7+9OEabDoz+FNw8ZNajD49YUKXvBrO6+V12nFYFXDDz5DE8GV6
6VIRXk+b10p60tfn8Aig5Q9Jvjxa8SIla0yKqeocNfTq9kyJVA5G9142InqquVj/
5xYHyCCWOwSZgjyPwj4y6N01B+XtZspI7jtoymfyCQGlEii8ZE3FhDz9yEnzS7Fe
VXYqRJGF5hA92IbxgsBe2erZkx+PWOANpPzPRTEmaDJ2kNpapYlPu0w/q+BwnSew
xUZxeyK4/T7JJVkKRZp0CRwZbtB4WST8uyf3UOed6iTVieh0Pgh4pQPKPnuqYVuH
4ODFkv+NcyHMwUwHm+AFBkmx/CayruiC4TQ+3fFCsJLyvP25AM0mdb57LUHqOle1
KrQTeZh8K43I39Z2cXUIe4ohCWmyTvBpAaLaquJYQ54uR1L3HgTqkrO9gPoOKMWT
x81PUmgZ6jZVwHV8AduJpdEZiN88N4h9uj6MP9mAeYpbC75fRiK7bOec9isfaNF3
ulnEKhbC9r7XBShRvFHDkzRdZdMjNxGogkXZ6Skt1K4qDXIxv3cmcQxfvWGNbaKY
+Dowo8Zl/C7pWMoWJGDQo526MgfNj1A+UY2WpYJhsMu+cCoew4cUvS8gvnc0Wxta
D5WwR7DDE4oXkdphkvxTm66T8wO8Lt3j+LbKi5paLJUN/EsMkffcd2cQMd9EGDgr
gJlwOmwGVGs8Vx3uFLUFexoDdJt1rrEeNF81wWm9xwoeWRkTr6aDiCJZSoiaQMAc
IQD8PV9mMylRptpLcNJkKFjXdUldi8n74vC358BGC+M5NYzWU9W0tQh7zQpkUe3g
gmIz1SXmbbeloJ3jQOP2pyFsWDFt5vkLWzm6vklpIGut+VQxuJwijPJu+tUk2ypa
Sq8UgFX5tmU03rDER8stUuX2ytRdBiX7gtOctqipqEpgOM9IvIw4JTXu8PhijywT
lyVMMXobM6DvUOSFYrcZeIT9gjmReGgSo6IEfInoOoMvyNxAgTXJUqIth8Tcg4Kj
z+AsXdg9+etxJ1BP9vpujJvmRxLCFSaMLwtn3I4r+luig4uFOAYCLZMNfHKH9ctk
nSEASLwxmAAKzJwBYDYX1Zf36LRiX1cYWxdKB8noKO7qjAEOeGluagVxljQ05uCd
wN42gWbEJp234ugwPcZR78N/KnJN2dRPL8PzRMU7VBNS2rAWbANlpXzrkt+XQqG4
2H74j1dpMUIVGnW1oGchzYslljkT0roOPu7U2K2BJxNMA40j9cQvymEWDJMtBE71
PBQ46NdGcSx7g9GPX7wdmdnH/UVPGL+aeb2g/+MjdoZoX6yP/FKzhEvQfbcYvoUd
uA9cJoa7S4IiZK2cXCVFPo/GS24K6TThTebhjPB75ZVODLhLrw30y6uCOQf4dLDQ
rIsi5jiU8tMTZdvcn/iejidBjCEFK40vr0gFdZ3o0h8rAQHOrZ9Dzg9/wNK7xiZG
RjqBfjsQ/5vcjkd6WfGZscSOKIe3Sv6xoK3mYUfndYYxQIYAs7xxGLOzOzuGq5tF
i42YeQ6+s2De21EUCbtfQpG3Ecj4IGEQpRqXRzJnF4c+KvX/N1c/54e1tj41QoHu
0PVqm1N12www/Mr1bX7fddUF7V+fsy6A+rlhLWvNe8FYmLoBXx9lFV1uho5V7ysF
dP/ZwmJDTFJex0B4W2knYHVn2wswiWirGJahC1M/YtsJ5SgPsxxq63sz0K+q4Msb
nQ/jZM1z69lOVkXCpheqfCev/P4uKi6bTShr+Tj8zFR1xmla1UyVKxPSa7oVWYLt
EfWwzOhOuwITYwODaxROciHvT0NcbHXiQMb5sxRebzBNKV0+2LqaOnPZfGlY5B69
dU7Z8ajJGb/3s+S2uReZnRtoRzGdjmv0VDAw6A2m307QImFr2p7OUfRd8r/jUirg
RWLMxL9ibI4PSgE6ushA0gKUptYo0o/pZZXW1ehbYecZleftR1n0Bz7JgFN0lD59
w6+DxpCeUjn/LaGzcXdSnsVgVZzRH6gq85U9XGwvaDLR7oWaecNUA6N2oi6OL1n+
4/wI8lrmAsVnhD0/9/jLY11XmVT2vdyI4nI+kwNESsB+C9jEt4Wz44aTUWGwq4+L
IkYILhh5K+uU8JDVrzENlkwVmN9yLffutI9A2NTPxr+aO/1QhW5YM7sGV9646TC6
/E3JZY1x2jXLuqRC7RnVprb2IbG4Aw9oYcjpwOlYYWxFPwPBRS423Ji8J5LJ0T02
7giF/3emTr02z2DHOBrKvKNZnowWS8dxmCret0qkljsTzB7So9Dhd1iPQp7peLar
coIXMw6WjlcLEOmMoWuk0dsxTUVhMEpPTuJV5ifcfR3WXCk1jZPsaJhMpfVIERuq
ScATq6HceMR6nt08cGoXbXUuS4/mSjAFEqeUA2HmTmQ5p2m4Oz8vvcu1pgAkjX1a
OztCK/N0O3Aj4vE2PAkxZaUAXRRXk7fvncSXP3KT36Bmld4/bwMQMXgESEUK6Xwm
Q+Xhg6cWID0c5A5G++VFBBn6CARXVamP3YB5oKwIWlA3hVcrWosb1aCEqKq4R0ou
sBSLQhGRBSjkM5wSP81BDde/+33fUzUvWgQtVI7tUQ4BggaNt2kUwcFmhflmqps3
LmqKcIcGI3jDg6RaFx/Zr6cIicuP47+ITPljR+vUbqXpwC5CdMPdSJi+OkiEV1pF
mhjVYZWzkRhETFlGa62GHphEc+R23ZflTY/K5ye7qmp/FChpddkwULBxixl6zGdk
oglEWEXtd01EF4N48rMKf6Y1aOCWb82LvsAn3qKuKe2fDjaXaxrDUMm5HXhzTmoE
Q5mQl5Kb1BxX6K6XUc+gjadfr6ZdqY/tmXBFxIwAvjQGIP3pseivn4t1KDxEM2Sq
KFqA1GDsS1sJiq35+6r9DLipCAKaUSIivw+ktXK7At4LInikDJpToCJQBU96akji
uMOC0KoLGaJrNTJKyVdCE636xyWuq/Clx+uIr2xbipFsFQAYma5/Fhjp1VRQciVt
24DeTZTLH6LsrG308lbOtQA/0kR9SEXIACIOIs0NyfVP7jY2Vf7Lwm9r032CI8RK
Ceb0UBCAqUhaRpUyglXxq9to4vpqCvRH5w5uA4TAeOYVlAQg0cGcl5h+b1hgFCqf
V3BSXuH0YbRCDyaEuJF3lPMI+wPlnO08H18rpipO1qznVnm1khGHHTthJkkr3GOh
1VMdFlldogVcvEwYlBL9oGlkHPbd8RjNa4IjAM6iG+n2NytWS5V98qwEeq/MPG7t
DUYE73wVPWYarTHfDKt1qhwVZ1yB27hkJVRdv0JOTCmmjWeDOOIaaC3PVruu2CZo
CyuOPhLHdZZuzu4MInZSn6ZSdHtONLDggeSbVbkz/+WdtMZlAz3JnKBMTWNHxiW5
V1+uFTZHfTIqbsH+kiZTsuznvi+aYfky3MoqDDfmnms8HZTGevOTHoUhMosDwrXk
8chyx5vh9pN8W458yjkA9GMb/Qe9bU80uAN25ffR6eByedMRq1hFZoSqDT3saGuk
UCg2+dY+IV+iFQ7J0oZqbUL3Yo7o0LxWsUO0qKCnPE7+O3TX2DhbduH+U1Eov6Ai
33uxGe8RMUUhr93aOkLFiMHws5u2sTp094iLmgdeEIikIypk4L8AjqcSybe9hsDn
JPti9mu0Pkv0IBOa4vOGl0MvLfvVEWmzosc32GpiszqunA4Iy0D3iTdezAEzmYak
wKwM5zhOJb/ZJwqL4HkNqdZhyvv6XTlUgRGjVrx/J0NEiU7gTNLIVqNPXEA7eLev
ytyskJuYin7H/nCowB/Ah0PZwgb2f4+vUCILu7sZo9yw/htooZCsLQb+2xBy56Nf
A04p9nu8gFJgV+tvCN8QuZ/boG6T+9qv9nQdIgzRJmIcy4b7m1pYp/k3+pV3n86t
AJBQGkcV1MRRuZBU7qNjTQNRIBKU7gtumpvSxxWe5ggoTgQeweefrHrrtpF/0VdZ
rbge8eodJkwdvWrPyjWxLfIdsquQ0aVqAqpVYbjQXrzIkRKsk8jYYkJmeCzXbAMc
jYD/7BI0WXgeQRSZBBbsqjRkwECZaqZomyZ3JUcVPHaJmV0byB/Qij8p5gXnWigI
tEDbYUEeGoDrnfmSZOggzLvMjEyItQTUZcVj1MK0DmR2lPv+v5G6Kx58tKkOHXf7
Fy6CFYWhxixukMLAWO6Qff7TxQojNSuVacOXJQTP873Mhf5bTbUHnftIs0iyMkOX
ecYergm0xw2Gq4ExMbqXwPaZCD/1zMFaLu8BKRNrdLu7LOSP0Is2Y3vBszQGGU6Y
iy1+hi/YbyouYDWAViiKwV8yiHghA3ABZOX4H2G+3PAYxcYq26ntC6uoPYHAmOmK
MsYFtSgrXIJliivf7V//x7QdW+Jo0J0Fsqp/P/SxyS3ih5TgFqroV2hzXmWqPK1p
G7zEqc3ppw/ywuEtyUI9WZPYS6HXVYSbhCaBYUD+gfclqn5V5m0ocNSJ0hwtO5aD
a/iFaFlcCVWsR7etLLxLh3pxsqKJOClBjawIDFl9CgSwtVVErcYLHIADM+WfAcQj
GnBTBxMJj01minBU8KJ+MJHFulbvze8qac8H3JlKWbKMVbx5wDG+KmFhUeZSFEmg
t+XOXwZEl2zREsJd6eLABTgWFXlI6SJrgnK1YOFqAvFhAwcrnomLWV0TwvDeD6Zi
ZATkNueAf3IL686BguucaPJR03wk8b8MTDRWZlbXe66cmJw0LpySSz0pbTAUTrjD
5KTQdyVn1VL8xYix2Wa5fH9PfGplfyFlnNQctHfiB5QdOAQUxHiORBSmPOus21Y8
MmMp+bLtOgvO8BT0mgYntFudLGbTgKNtA0aXCAB9jENZkTLsEvppcKEW7dwhNsLs
M8eehIH9UcWZTeDFp/7L9If1DQLZ9Hi9ourePcfMp+0JiH87eDLrTxiUfTLlSmkP
ZqjzYtUMyD4EHthfl7C6dBo2era+zhKax5S37kAsm1crnhK5wf/5EJoh808Qs5zj
HBLtCQ+pTvz4+D1MbQqvHB4Ooli5VfXlKH1scRw8M2uaBqNII6kto9SOjKC/06Fz
TK02Gs+w8a/UFJIoFS6sfwFFIgGW6+Nds0H+AKUu2PZsxrWNT0n4iUeBvaT3dJeA
NH9cHci2WebEcj+/ljitYctLeIRrbmttUbz8H5N5JnUnWK8ksJuEotjnjHK5zIMh
N5oGjyrWRsflPM3TaZPDp3w1hknpc9OqpB6G74sAfUfD0oHoXzP7QAAPThtCPJCN
0ebsJZ+bVWW/gpPoXq43ZlJ7yO+CSpXSgcVwKpWDM+2x+GErWTDGwTpX0p49aeOe
o/flXo/s3Nb1K0pMuSbjwPV3Y+VYTQmvybscbEGn+ft9JpZmvWsesOXfiqcoyadt
+DZ70tQYwrFgRJ4c3Iv6fezzYSfa0x85X7zVRAwAjMe2ujoI4JsEdOfvU+WRZ26t
wiTUUhUSXBf19JSw5lq56C/Rb8GQojeh6mTXfaOU/+oksZkP+5Mt/bdPIgcvBcyo
J40wcmtoEpBGIqZtBPbkZFUs7jy///yXJyey4PLiOeKXA5utwuGcySDmlZtHJbHU
Uom+uAZ5JMA4e99Y8X23LlCi3ZKxMxPSNOuvIeHDO/LkhTc5xCy50h1Yn7wGyCRJ
uMFOdXMqQJvQ57eI+/6ztvLIyAeEbGYF0laXFRFnqeM96h12znDX22CY819N1MwH
9Aul43Mb9PzqbsEB1NJng71pAuK4Ait8lx9TsqPBR1mfOo1QvNJVidWFR+1JvgZb
0IRNuR1FpNRuB/I/3/teQbA8UQalMnTZrHp67BX1FfPGOlFJua662kL0BdfIOEXE
2J+G1IoyxUr8kVXMD5jCKwDgtZSuG2ePNdCBEUV2CTJmDO62bLUMvzdv74bwefE6
TQV4fwh54q/krQufwLeHq0lnAtl2GWpRs1bFj4xRROnz7CwCsQs0CA0KD0JhAnsG
kgWsfF+ffsjNCbdIfNd9xuMdMfex1ph/VHER7UJWkjxB9nnLz6IRODb7wjbXRKLF
6SrAWk0kXrgLZY5jz7CcHYlEudcCCn6k+9z7wN9ho0lnayn3doKFnR9u7S69L3qh
Z1zboBsLaLp4WfYVuteynOktqDbu8Ei2t1Y3XNrepBVpO+FK6g61NQ1G6L/7QDuN
AHqKWx0cwICIPMGBUZDoTdHcb4wZ7CevLuq32szj9AbWeCABV3J7thCQ3Krcovv6
0sl7ol2tiIUbkDSeNb7XczDNuqJEpvdDAT3h0/sL+eXS0VAbtKXQ0KMm832OcI1p
SeMgiYHAysnRvMrEDBtjFjxX7nnZaybCJ8fcmzOxtFzFfCP43Nj0AFjPuz1xYgv5
Q3P7HVtCiH9WVQSqMcQrj7r1cNC1Q0gIPdeA9Rtne2ceqHEo6maifo2eduKynEjT
QJcIf7UbV9uvUcZeDQD514qE+9FNETfW7MLCUR9A9Wcmj/cmH9x7DmDT5aZJ49zL
fwRNpb1o1qXPGhkekvWTGz/aG9sa7P8WRbOyy7BFh8Nm1vukfvkDtfHvpnPf3P6z
fAH/jcV8GX5m1dxwmHC4yWyyuA3m7/oiMa137VkW5E7wyDgMU0HU1Sqj8QooAHrz
1pbuLtIwf00pYxDComUUVzeBFk3Aeqjpwsh8S++nJEoLaYAVu6VXNnXltZTWJuGW
P/wpUF/KVos83OIeqQcowzwAw3mxVdMeiQS+JIwS2QEZaWLvMWOHSuqlQIcs0AaB
PSuQ0IEAjO8MrhSDjlqLn1a4j5CrWdoRqzKWEJ1vgr+pOrVAha51Var8J7sTOfOo
e/760xnmpReZ+iam/TeM26LEDlD8z0sv1afD9lXfI1xo3nijKuzn6ZaZAiq20BKV
rBls1QhnqvkrwpNZ/PG6UczHqVCn9VXjafnqlFjyPMAxc44UygKS+fq7U8FNzYd3
uJTuSKQqZKh74TuEudCmmQJmzcDCzcTXJDcyjLwERZjlWZ87FrI/o7fYQ09NqAWy
qIIVSdxTvuGfVoBBW+klGlncKnfYic4qUMcSWo5DxssLhVdfX+noBFNs4Z00ouJJ
iesU+or7FsVbVlNStAPSDzWrtZQULjfewhqYCbfd4mos8x0x1c9EpeYDwZqM3duc
omTNFs2+5zgo6dUp3SS1tH1yFyKPaf1XZSc3vmtBxi0DjrZDoqnItUMAdCBZGMT9
S/cmIkhS6nH+4Z4P5BNdidIk5iPorWAKvxQyxlmfrbxEAzbMnYcttFitKRDWxJ7f
iqUDgHgYKWNWl3+sKv49w0I7ZEkI3Q3RsGyOCd7aVHJLtrTf2z8wQtooyyPyQH/q
oBBlLCV+iCRG/wBOlfXO3CBglKa004tvR86Y2PhY9vRnwdMNCvQpJn/pl9j2jmkR
9mGrchMTpg0HN9rzwQKo1PB+WOuvMGkwTF+GjNFi02MagPiVZhpAqk0Ich2xtczF
WBLhrZZPrpzmyxxOaP6XE2XmtbQJjwL1a4222PoLJ/GSdG6V5qf7IaH8TX9QHqzJ
EcTZ17WjS4gOupr+HwJr5Lka0j4GfPgOhzOq0ZDU9osCAODVoJsvN2K6UrCeYXow
TbIyeRnx0TZnJF1q9atnhVV4DT4SMjsaUDy2FFBFsSUTmWqq4Gmtyfpu6iYv6g/3
Q0JmUrDcetdY5Xj0QgqFeniHssbgjZ8HCF1STW+cZ+cE4Gmr6dzlR7JpxinkB4NP
0HIM0ZWCl84qcPynG2KLTJ978TDBiXO15elOnnLKR+ynaPRLslG6eS5d1ncADWnT
en8aGyt+cDnPLbE0o1LZo9vLoRKailEQnpI3Oo8uuX318c8kJav7gdm1pkjh4/Pb
KkIexlLpCuZEFuHe6m9BBMjo/MG2Q1zfos/IdcZTnMVryjnyGeWaPUrYHsurUaQx
NGq/yHzLyzgCP5k6ofcq/ay56Gq1aVN41RpJ4jmWSb5iIQWUsNSZEa9kfIdo4g+f
1ndsC5U5pQPc1oYefaOEdTWwKQ7SgcNc4P3S9BHtiA/nuGB+Fe5lIes1+YoXN9dK
H842DCWj9GFHk4iyOCyI/7KbTZQUMOIqrXKYKPnLvMhEK9LghxXtqDdEK5aOhqwk
MUKANEjS+d+1+oRzs8e8LR2/trKTI2/GNJBHgXFDnu9hXGzR5bOef2rPvD+PS46O
ogoAQl/868ya4piC3VDyrx2y49yOUkXoRjfpv9EcvBUh0/md95inkNUxX7nNBhnH
EpqF3NITlZTd1xtf5NTvOxefRzn7XK5zGoTWpB/D/3FdrHEAwXMoaFpBj8QIvEcO
ZqvARgN1pigv8wMxTcdqsn27ggJ/iulPzEjdE5Ma+WEDbBXP/7/AwiI9MOWaz2Zk
jq8cLgYFNuPzRIHxDz1Sa5MKRlt3bcfgRaXBdXbwZjzt8/ZClPm3qZsLgeIxlDDi
girEk8ve6R4Dc20xwJFs4YzCaqlEo3GGfvkezdu6Gy8S52ChHi6uU5hwqLC6g/nA
F60YJFCqVAX7fYv769CBDSCYDM0yw0JEf+fnC5rylUuWjhI+f/XoY6SXMEe77TvI
fnfU1iCwcFjm/LDTKCd35XZTwldbcqiQegXGB6QuU3BysrLT5S7vRHfmRX7bJl5u
NAoIrg2F0zJlLcwOQUIyAn9fxxyCnny8WvyChyCPK541tNKOLuIiou933pUnB9a2
NN9Rz/XIOS8xZPez3q03nb91aIbpXmrc4R3xbQ57ieF6aLEANA2ql1U4MiK1o7s0
K/tmdi/G2B/KP3dfQL3oolzN0g7DOhaHJznzA2bZeBgrXugBqavyj3Mk2C4fd6lO
1H1SgI9viSBjFBq0bqQaW4K93xWhk+fjqwuriGr+538m897vR+AIzGcRr0IIRL5W
3pCFANp9wP7iD5Jyhc5vgvHl/pYmvDE5Ttvx1pSM7ObNC6ALIVXvOFlU+MKY52xK
IK2zGk+AOPUq8xRBTDHQYlmDHWUT38OwZSbG+muI/MGJoev5ap4tpFiCZ7e2sQ8F
+LxrT/AwYDFjN9hxUPh0/bOZ6aP/lsFDkMFMRfFtQVw24tZ0EJzkfgcyMJGeXCMt
QfkJcZDmdgBaXgH/KA3UMDSB4NG+9xZrTlAyRwVE9UDJtScfoYwID3PCVGpq0iCI
W/pcBzo23PRKDso3Hc0zKPeek5avwkXE5D3NGT5jev+aUKBY+kKnSUx7wapj9meT
vZrkE2qC5a3rsCHDqsZ1CAEbNO96+mcKe1DEM9G/wTb6Z6yYcmCKd7hIS9oaZHvs
tegIr5tz+UVR5nW4uTkp8BWFiL3bwTKwH1okuEvROexnKHKW0z9Z1GmrsEdZ1l+f
WH/TP2Pd0sc3eJdlzW9mUhz1xqR5zvQGj5Pdbptbyb3cNzGme7m4MOKg4JiRmVLX
lCs97+ksAQdKfnoOf05wGD8FjueLN70P2PwQEEijPyVnsYnDVfd0RkTguTnqUBB+
NGYePGgMuhpWMAXBQD5JFk9TeR3se5FdONivjeNIEX2oUVdd7+QsMTfrVJdrheNk
vz9DYvtv3mvTjiqZDSql5C3gIYo/4BGyr2CCc9ye/zPmibM5NMrf1KQfoJPaUzs4
B9BVF5fRXdHasRIQtFj7sYtcfcGnpmxxFFRT2IuvD9FwyPVKz59kZlxkF612+zoN
To1dJrpRX0+qKp4PAhibtP74rk7FlNYz+yYW8nqwQs2HKZWvaeW8bG7lyrOUDVV9
41kbyduzpEU2vviLEJEp1W5E4w3y/YogDHt2KHPbvhsVOl3cqMFLdFDdJMLEhnx8
iY79kzFFckeOLzGZI7z+1vEbZ8mh3CaXiQfCA6VCugaF//TvzPA8Lu4tpdk02S9i
W17+DPL6MBTpLlCM4T4L3OIH/AZJ/KQW6q5M6z1rTRL3YN0DHipuEkJpty+y8Yjl
t+o0zhjRHCSBmosL/is+rXc34txl1zCQCBF9DAg0Edl+iBXZzlgKhx0ZTQ15RMWc
dETRCUhwnbJnwzIsU2kBvFI+UkTbPKl24idmStFA/2dZSlglfWU8NB1mBHu5U+64
+Fdcq1/OxRN1i/sRxUcUK2MGsn5YQ0YI5ltyZtRda8CfxtVRODEkyTO/et81UFq7
pb4y3ocEfm+QGlD/NuGr7xz4qNCZaVvB+fCYDJAAH5xGaxmn798zblw47Njty5id
YOmmB5zGZ2lRHx3Na2kwzifnG1b5C61e8gipMGsnZ6A40D0PjuNlpe8f+pbB+P57
zu0VvsGFVBwBxFg/+OkBYcm8WmeY63eLqw22NsjnmHJMcloBVvUsKhGt4sawCfaI
RIqpgpvwozcf/yp9nxHauMW8UOBTqA2JhvmCyV1MyTY0+aHf985n9+MhseStBLFt
dll0/+22fANwR2VZHyoikAPxPhK/0Upos1/N2jY2LTA9DLg0HdKfqyT1PRlEEseP
H2TW1+cK6jk9GYPcQjeSLXMCxqrGauCJmGtG3bNyPbKd+fc8q4/TmWe2y1wLpd+P
ohLgd54Ot27oR/nAnsFlILmwZ/JPYw3o616ozN+ipRXPTMjh9VpdgPGbQJnHcAex
by5xOnXFN9vSkY8e79ewDe3WU/ddWtKCknbEtV3dz3Am4sKUBGkdsuOBKTgryFZV
jehDwWOhTsTIDloUbKCgUMochLC9s2jSZPzxgnKA3LTsXFIT2COrMQUhK/4ivr6t
5yeYHJLIv8JdL9suJGnssgjlsARDjYLr2fC4Qkzf+eXW13Tp0u5PUzgYRlUfugAz
gC5D69iFOHGUlfegTaHCWUarCFxKAg3o6z9yKOBuf91Q+XeGqKHg4v5N/Z++XMDB
0O/NUkfE6HUzo4aaAM3vhDDCc//B64f+4JCEpvNNBO4tWGsyGQBnlMqe6OcSFuFN
RVfRVKtOhGzdqLV5C6w6+I9FxJpAyQfVE0rrTlAFAE/YM3KagbqdZ+TB+B4LFAUe
sFF2/SkTpPx4Q5wOPh/uZkr0vjP9o+pPnTU5uWy9uR7xAxXpTwrIsaK3JNpykTT8
4jYwzT2WpcFXx+T7xTgkU42KprwbdFBk4jdPjrZj/WWbxnSZd0lhC3+F14zJeiSR
QrFtWoHXejusYRTPJs1oCRDsWY0hAOnH0fbiy4PdeKAkzA2AIzKZnVCG9khEzYTt
CsKOzUl+2F6vwxFHN+be0Qi1rp4eTCEOHda/V8BTKfvbYgD3RZzT7skKUkU9GCfG
82NC7xm4eUGv6MY5O3zlYhVI86hrov7vpdYYLLrD1a+dOnqqq4N/q4qgDxui151w
W1dKn/DiYfR3Ks4X2joW02p8gSAjfVs+j9YAGmOTohUCPesnDwgF0EbqxstjCt3c
doY8x/13mf52J2eNoHN3FHfMx16haBYFC2Cqfd7Stvm711W8WMT8/a0MGqVz4KAT
JFaBmbO+aF9YmmT9pl8JQYvMwSqT7cmqwu5moitHuaUDo6D448vrEYpDBc4J48JR
OADoxm14N4rbcDNc2gNPr7t7k784Fy/iabss7+u8zZKekERmf3nnBu6jFsKQLVsY
QKpHrMaqIT3gXxlMSPaCJIIKeMmg9hAuGu8MxRwj7kdq2kbesBcmWbHz0xKcjpIU
HOpBNx9rVYDqVGa5COFrNSh6hXmRTc8xe51A4m4NJuyaBkiMnbCAt1meq83KS7pA
vgwTCsvdQgwxj0oV2INrzWRzqcIIM59ERS74HPnKf94dejqkxEEeaf5i9HW/huUU
+GmCO3YuJgIfvWtifrxQqeQFPTP9HliGrIExBMBt5mfWdph9csu2gnf+iCLRhp9j
kLsWQogeRXyt2FL7zYk7E3FEfkHM+wdS6/sw53LFcN0JJqFdgcWt6PV7YOBDS0wA
uGtn+koJvfkQUlMu8yZnvFyr1gaAUqgjrWtvhiKzCDF+X3lbWISbAhNy+1iMxOlE
zkzzboIfBv528/twifAIgYFkQCSnF/BW6KVR42hdH2JWxF116QL2/M1UgkmP3ApZ
59i6YzNz9wMbG0sxFrFAPxZl8EO9G3rF0km0ArTkpTPH6Tjatj7ylWzw5f4PzW0P
hDr9NN6K6+mGp481HlON7dYAhakz8+qujgPhmnGZss/a1u/HjZVfHz5ET4GU86TE
amz3rdtaHW3lMI6EDha0E4y6wixBLYTNB6+X89zYTRSInnJMb3iCXwHTkIR8Qr60
BHh5cmi0OQc7+vh5E6IkqvKF69zkqu9aAlaRwxFOViVNZwy/PqOZybXbq5cJEdFG
Qpcy3l6OQDoeQtVng9Jvwh8vXtCJf/EpXq2K19jRHtvq/UAoijSOh+T/P88VR5wB
dbGZOF/42kIt9xUyRFsbj2VEUJOh1C2bIwpTIXDvju4Ah5kyM22U5aHL1Zm8sAWO
55lKIFo6uvyGq2J6tPSdL+m9CKG3dXCoUBV0HJ079ojyzJ5sraDm/2ic2k9OVTl0
mnBRM+vXgM5/m+1xBFDDSqNrsenosFRFhdrxxtEuDrUFa+krZjXXKXjq0CQhMSMj
L35j7ZGnAOi8BB9YS5AaTcyiPDQdARdcKhCEN5sn9jGyg2iO47WR6p7HLWXJ1vgI
gCKiXI0ELHRtte9nHcDoyVJTN2E7cT0wN+R6++9Ey+ZpVBYlAarvJrZnm+OVmT9c
nLUjazLL3JdPy2pABHtFffhGnRVML8IeOw6dYgADVatGMcBLZnx+25Kl/FhHoisO
EUj9bH3ZXg9RbiJQ/xu8Ld0gdrTSHwuGkceeLLi9sjHM0jgyTBJ9Zthj8576cqIv
eK58sPDmvP2Di1pcMSWHckv6yx5d3GPIsoGhrW67jWxaX9I35BxXz7P9ujI9kbXP
ps71y6zWBxbzaam+MKiEaVSMXTpsX9I0xz4X/jyQXo1DoqSHA0xjN13l+Kxl8o+/
4Ul9+ijQCnSsigMcNSj5UXWdK2himvVGLTBZOjVesiZpolTe+Nlt3BiaQWR5Ev2s
bcmfiNZK37WBzmfDxnxO0qgCRQh+2fBNv2YkXD6FsoU4RSU/ArwbWs06B3uxKvm+
OsDTIsst6tcttgEatM6jspE+oMqhmKefYR4M17NgUBIz1FhJOE5tm9kXm0vY85t+
DFwDBOLlzYktQLOQzcdVCGZZM6XW6XzTENzQ/+wibyScA2z9unAhIvVfMSXNO4VW
/pvnLeVpjbSdUs4Gpshn8G2B2oTgf8OP35Dt2JyID4haftlD0MDotYbs99VeiLCN
Ba5SezTFTIMDmTM6Z1JZe8aaXgY8xXitJtbNP/DtLB8qjUkNuoWdu31bFWdp4n0R
LemFp9jX78ZRYOcHGWNnlto6R81S8WzhCyxxd+QWIhYAi+HbzlMdSGIByjQj30eE
FXn8q9ufs8fMDoIcpr4mpgOz+H+bFG3oo9EFkTB+TwVHVNphzoC70Nsnm3/MM1RD
bROcHcX++Vz028r0rC1q6NbfND/5EXKnw0SCjyLn+x1WzMfRsmBbQzHtfxw/aa4M
R7msydSB2AFMNjlh9vhGvfyR8qV7N0Q5zxFTZjwWzJ5S+4pJ57f88kuY8eKSOdRS
F5BMLNDhPIxuP2k9SnHeu3Rp1Ljlc2BY/iYfVFU/eE7uKSDptlhrKCVl8uphY7m1
bJ6hT2q/ajn1PtoQbYIJSUCYMNSxgtbCvOjdeOPLC5QfPTEufV8HD9akfvPHMcmD
oEjq4l/4f3PxyhWFCqWlo0KW4vPUnKQLpIXgiCfUeKm2ictOVCLmOonbxQiRb1Kr
OsY2IB4pp3CNqmZmAeGrwq7Gzf8IdqLvYeGY5fYjn2jcSYWSfKsE9o4Qcja7CvH2
a08f0podWgXhvAV6DoIuiFt3hzhyMR/4fz9t9WP8tK4nSrV5FRsbbVILG6vJmGrn
IbHI/uWTaQQMlZoVdWMR+jhN0FuSGuu4p2teuJW8uAKF9w5lZppnNpQdbeVtYuAa
g4g3R+VH0owVJcfqbE9FF0Z0ZHa9QlYpAxUV3oSSyE2dtbGIblUK62G2wcdh5TBo
aT+VudTyCTDcd/xi7M43BMQv2BCrdKfUe+eEQBajMw2KW2HKwP35uCs6GWmUDgHt
a1vxLdiqvXVBUfpQBDq5VqUJUqwhTgHFV5Qr6EeCVtE3dcy1XgrPzhRUi/5vG7n4
Qd4vxRdiIOOWKsinJ7QtpFl7tijOnkmxiVBJvqvBSMsZkGwBuSOg5Vhz/63iXVuJ
bG4ImHoQq2V735jBbPvsu4mRKE9RoIpdX/A398cF9xy2O1XeiX2xxcfeMKvrF2/R
HxdkH0FO8I9oJagHnH3r3sQoFaBZgRBHNbNqA7oLPO36wtTRUC4vuZ78jaD/b26e
xfFuxW6rnFlRQl5tQDf9YKw4P54Babk6wOFw4bncNuyG1FfymDvDbt+t6kpBAXjf
GQMwa42PF7Kd4S2IJA330/ijX/jUPJ99zlAaHg1AAgkdqNEjtXN5vTRQ3lNnUlyP
H/e7sBAd9hiJ69y0EGye1b50/l1B+RHlWtjfi9CQpudxU6ccwFtHgzYxFgrbatDA
BNBnQeGD9nOb/D5V9WddXGtbRttY4S7JBMYQRjRJMsSmcaQaYpcg/CKz3sInKpnx
YFWgu1Pb8EkzyRTQ8rcxSi5KSX9AIAlArowlXqsWNdQOMnA7p41Tgb0TXdiJVZmW
QqMp35VmLkY6/YQe+4/uEaeY01nAK5FXd3w1u70dw2df3fW+KNgBYDV/YnkDKI7G
huFr9WhBiyiiDZbooDwEro5Zxlm3TX/gHEj1g7fA9YkiCKYwO1nM+qx2/Hb/rCR2
J61s0CnyAs7P63m8qGUSM2SUjBUsOk477b1dPiWTz3iIW5X/a6/fIVFXjFGoF8L0
8JymwWj4bIEtnL45hghKA1vbTNcZxSOxs2rdp74wVsWvpltEsaMXgmTT7u+JzGlr
WdsBMrMtA+s6c7pMS3bC30TrH/tUR8XaZv6l9KnGZi3nyMugURlYahT3myrB5ddp
wnmnniSuAaslpPXNAq63ruPGdpKosQlZZ1BHZh0VtxlF+qZgn4lpi6jp/6peARLm
UBu0z6UX2WJL+ZM/lIIucyTufWCqw73ZmQa8JJwwPFaJSkslXuoHCIHiYCRJ7cN+
O/Z9WonYvA8u39j5paXJujlK/gUsDfS8sivZJsK7ChBavAEOx2yMwfEqGjdIgfNh
wEns32Q6ah9tpMNIzoT4aCikjmqEoyPHL1gpin2gd4FMrPZn93fqTYMuW3+ZuxBp
B6hDg7BEqDEgDvfl1lZtBNDeMiqTBpdaz5iErRNnnuHyey8uz6/1ELkFAAuVpVka
3iXBAs0ALkn2UrlxjMY+9MzNO28lYYBEIyGuwWGCYW4kedtRekcj/9kQPnHTo/HT
CdvTyF/cxh9fITSA5skAsUxeEWjoI9Vvuzk1shEwQ+oiiwTXxwxl29UyDslAzsLu
u1B4/oVT7jQjEh8i6A1UcR5RmKqwwZEOhaSPpQ7nYLWJfcZ1psZpsajM5INPwuAg
wl3G96GWVVdVQ65Qhd3EWF9B9H7/pDvCWbZwmK1sgEe80VShlr/mwOajx6X2Fp6A
DeFfy1bvXsYxyDlnQ2mLUTsRtub6DF/2+5J2OlH2oKAcDhnVBua7PPJ+y4UPMj1I
A1nrxDdIi+AC0SRLZvJAamPcTNMcazXKvvNo0cAY6Wu21asSEiOeY3qwffL9Ewhu
x0z4V7RD+oOPditb6Gf6A4ugJt6BXxJXWprGiGDo1drlIlEhoTK6YOMScUAZ5id1
wbiNJnyBVQ79AUQIpC8d/2H9BrRN8u6OXAY5z+O095ntM4Hu+n7RsWCHsAkXmTQV
MxznLsLGxOB0f8zmKuryU3HTFpBWTptZdAl43Qfda1GbdFMEWfFYqcDwRLHu6c/q
UqQiMwFMTWrKjoETg6dRsqQVwz6sJosc70SorxN3L1EQ2a5pVXDt3jXwOSh+29jZ
LvqcH3El51aeLv2/lTNF8liCnWR43cUf9qp1ULxygWdUaLyT5GgduuL+abD5VeGE
f7rHlxC9ZTBoQE76fiWqWcy0j6rqHwUpbGLK52AQ80vQ0O4wbGoo2qU1ENnoX9RY
TSAF65xj9VHJw2i+ShbRLLXtfoRTTmPWWvR9mvG6m+GJjwPA9GzklLJYuSN65FwC
E/bOZW/bvdzDnPCmyTVhBl+6KCnYs8aFwPd9HlT/NNqrQzuH87pooaj+2hRfuqUy
Lb0aYlkUkOHXwGUGLUF6ccCEb6Lts2yzcJr7xTwqaoxTKs1gAW705Rq+ou2tfcAr
F1t11pBrZWx3ap5mUs80+GUN3Xx+heRlgDrughoT/R2WAVQ0qOs1UyHCzQHFHquV
ism3xL3ZgbTdYpzqLKck09Hjh87jU7iLh9wpLCWpP0NRaMHGIv4Zm/of2yFMBq6a
M4e0cRXuhpuSsk2FU5cPvZdztzCl04fwWxWMKBkE87+jfaEE/d9RxohCA3Re2T9h
1Fiug0ZL7tTuDPhac3mFG32WTsgASrmcmPrsa9giIDFjfx3XSy5OMEXK3/q1frRr
o4FYxRk7cc2f6jaOiN5sjBej8doJyojq1WBhhrVc5KqrLG1lCMxzzoPOT3G/WYbl
GrahFbVZD97aAGvg2zMmdqo+I+nwH+hpiMZGN6VI/Ot+OhAaFl/iLNC7kMd4S/cr
T4e7l8T9BN0KF3zusSZrjklUIKNAGHKQWS3KXKFOHlBE5J53tJ2TB79pzHh+xX7A
QRGa95oC7WMhzAfcK3yB3JtrQsLiOQFQZVA6aTwqVkJH+GV/sE9OLjf2qj1RTrzj
u3SJuTLmt0FE4wlSlqDbtl90idaZbNhGBuFibuwWjonV2gO3ElEVFpX0SLnk9azp
UJ0KsFBlkFd79HlaJ1tl6Mo9eBu6luyQwa4Tio9+UBmnqjxiQ6AQ63VmTDqzycGT
PbIqhWVfgUT3pY4rKjXjgjizhiJEPqBqCGELUH6XPPunaCme4ErthQQx6jqrYSl+
euHlBEgAn7QnRIFT4AsyOO+oY8fymocpksE4NfPUvM3Hib38V8R3YotSRg/Opbwa
cMv6aUUn85eHYa87JpeB7l+9uZR/yYviheZAhOSbS464xGXBdpPItnDxyETgHWxW
wK6DYjVWhWjcqyxDg2gakk4fJvXQjpSIlzrp5IX28PAkOk4oZOnQYf0yvlzIFjEX
iozX+rN1W3175DZtKv/blKK+SwFxsXNhKKWth9NWBGOih8NynSf3QqhZcMBt5FGD
QjJvhitCuTTW8StC/bZ6iR0e/Q5htNApoSN5Cls+dTIzCRK/Ap2QwiPFKz9rmh29
yjWoznH745MLiXI1zqZJ8jW1EF0eC4RVNvzkYjmS3AViL97VlGgescLqiCnBQrrH
41l+eY1PG20VlblxrqUGeCJFKGujDHYXufgh8D4rLt7hBPB64J0m+FvpJ9qGPhFQ
okT51V/lQ9O4cwVlGLrLeTl4k4Jdh54ix0IHFTpiB4g3/1VAuC9YGjftpmuXk4Zb
sCA05AwuP9tLDn31pB9otVtEL4KSxJ7C527r18J9ACSnDjM4ogx0vdMU7M8TWlup
FKYYcomioB0kLDbfQAKXKeiJNfXXoo70QNbkdMfeH6THDjy7QzOC9TtB38ayrZ+T
FpVkq9hqIW4dzS0XiaoxN/QSN1I7vgDHxqm6F24wsY24dzLaXcJgceuLwecw3AlW
CUfO2ehA+LTrb396ihYR7CmB/6iAvdjIzJYCs3ZCKwAWadkezduMPvpV618TlPyo
QZ3NNLcUYdNejLcXwzhcvLNQjQjO288GUS1oZtBVkvl02vAdTSWem11W5+Hgnd60
lKi+R5a4z4CbI9o5gibp0AAViRoe5HL/fdmB+6dlBOO3QfH944Ns+dzECdzFbUG8
13eKDAZp/LKtkJrFw093jJLSt/J9YMLKOdmeS/Thom6uPI0pj4C0MFUJ841Kq8hC
SFZ5nQf/m3/Gz5JQTpf78KDA05m7wmvKaFHF9W8XHFh7ldc8HiVJxuXrdO7181ZL
uOYFiB7hmaDi4/NeSLI5CkIBdZ5+sTbJLCexHICkA24HD80HFEXvUNcrF64qQEg0
B8ptKLph1o4YJuXKTejYEC125k2KBOUCMGdYwpFoMSAzGV94Qyg8ki5bmA3QYBPe
0jgJqO7V7rBvI3T8wzOt6OZVTfeF2Q6CiTmyXFWouZMviTcaArq/lI3nCg5JCHI5
LRkFlsTZBA5Yx9VOPxAS4GJYskCrxclsu0R0IJD/P8EUjjPO7I5uQ3kavUIE03E+
e/oOS0KjAwq9iAI/Lp66+qhBVeHnn7nTovO6hMDsEwqLhfmkBAEcnwLY9yWshpnP
3w3WlFkErrrK/gCTfXrVaUR01cmHKqRO9811S76uCw30uEBSFxynJLp5yVuVhaVx
Zyl2kpycNbxhJHjhFqLWM6wA4PwYYm0uXrIuFyERdB8t7jN6rdEiO5TNqGXiHjc5
h16t6HZTMyBqCCIctd7i3soqcdAhPlC2EguHwJhYThEPkhJPmB/tvcvfWqd1OYJa
aKsCKMgWzyfKaNbB+y2/3sfl7hAW3eZrZpRElLjSMv2JEFXBKDljcbAJjwYSI+AX
9fLen4PVk1uDHrA5eKs3m1Pgn0q/dmh6eWaOaAFsi6Jh1Xo6ltpJQ67SMV1S6Pk5
MvtszzLUD9gAVTJ6HHE2G/cxfl0la3g7y7fIDD/5nFFVBI4OBBJcUPIf9HJnpBe+
o//yoLUJYHPCQY3T+39+FYLVOMYF/p2KE/7KXbHQa9RsTfOMoVj1dfqcv0fYiIOK
3W95s82ESmc+Zkn7mTBAHDCbwrjPsApb1LymZcUY7kXUQiJgWesncB3BG90rSyAL
AV3GlkkihsbA3KPbEZJ/ncNB707IQY5SZSzICHpa2l0O8d2tsXjnP8VwySdIE++W
zBlHc4YrY9tjH8HfjndbmrmAS2XajxEZzJq6oTVodMfReC7hxajzFNTJWXyVJq6+
Mhy/Kp6UnAjiBDONkXA4h/JUNT6CCGDRpOvgmgea8X9NijGzJU5+kW8CncUpSyjU
7dLCkTieaVXjQ2sP6RKK94TXFMfVxtfZ68AFh/8rI9lVdf5cnqF1DE2oV/OeDtTg
8h73A9HEam3mu7blksZcOWG6nFYjP8hBpFHNqFMGunnUOYzcReVdJMGrwKFa2mZ2
wssFc+32Z5FF63RbcUXGhQZqbKDD8ifSxRpf4u/3xEgfRIFYaI+OkOkcbu5yfyuM
IqaKdzQM79snFlFnUSuVNUsIoU9ZxhfqbW8GvNTYOCgR9/uQTTs0XjQgxZxIvwJh
ZXldO+Yt20/gzj//K3+bVBuR+tYXLh1YeMR9ysJ1WU0/D4U0tLk4W4SEYMl4In2g
SosM1SxAxmT7h7C/KPtCSXMh2gemifHg2oci1M5klmoLHvB+rhH55xQwK0XciQuX
81oCBn71mwKEx7y0hxiQOcCMp6RMRBG712Wq3v5i11dA7kuIFS72QcfSzgwQiZPY
b+HDmIoO5kubakk4GJLx1JnPsfCHa+2P7mLbI9v7PjisG9AamyFPF2otf4HHreNy
2RPQQHveuBD7XEVyvwgL3CzhgZwqBZdH3vXNz4c5FV3Z+XoWT3CNv2rdBGQgH/0h
hkoFb6+1ngxD1uGRwcA+Ul6HqgW227mFhO9AN3sN4nDGve7f9ghryqnvkPkx8jzD
4WQifzrwOPiximQUfTrpTFChUxnBVO0+sE8n9YYZi452c0TuczcoNBN99OnQbTPk
JSDe7eLUp6yKiQPN9NGUxQCb9aafBXZIN1k3oOu54zkuaGL9XjiGZEi4eFTUK8dI
bfnO6JYdC3PgkJTmGn9Lj1UgzofroBiCdbq/+9ztDk3LyM3mLk8vqstYpM2uFfYa
0mgXv9sTCmkmvXUK+CNeAUMK2VXgxV1lR0zTJTjD1mQbyUXnuZ+i5rjqVmuFn3bb
QuBd3xy6ClNm3mV/RztQ8iyGP1kvBEi9TKkAOHaxL+WakwVTpRW5YGgK36yb0J43
xNGBGWxyR63dr1k4twCc7S3/bMGHZK7dXwkCF0javZB5MEzCclbEGPxLT5Ys84wN
6Jzvuu1Nl79lY09ZfvlNWKuZhpyQ4PX9eNtfuCjP4AL87m/m8FVp+wWsxTifMfze
pjhHr6ieuFSzvXzp/fJo8xS6iXsR+VeIP7PxuaRFTiCvmnmJxILW/MSCfQXCJ+uA
mMsW/cO8sDY8zn9vV6NhboEP4/fRowtbnK8x9+4H4b+xfEHaiBn/YGGutBGNsL8x
k809Xiey+BXLnRWmqIPK6DmcZo8zgSSCSNPZRBWUIkCkKV9GSpLXpiY7anr33mxM
9fkgotjk/GubftN1jT/1xxbW5T60B7auR1m7GpykHsD55NdUKFuRDwusYfj2vEBp
8fG6uNxUHW6FjzSBPAPKI4KL1zYHRJrGaTvnM5TuXWzMPQ0CZBxOS7Szxr+2i7ln
Z4G3JgmSgHDJkhNTdMYZtyraT7NMFQQxHgw/ljzyYbGNsqHqOuKg9S26AqgxMSlr
aSUOX06+34IYBiF+jRfn7vXEDTZg3crKJLlJ+8JD46rdgRShusZ9YuYCWdApVaVE
NHG4vXOnddxHdEmz8y5n1fpqBIXjO4jxBQXzr3zysZpGyMBKOtcl+jRPRRlQ6gzJ
YF/5pf04LjjjaPiorEwqbDKBYDaTiun+RFZSZlDxsMjqAPDkZUdekZjZ93aE7UxV
ETDI6xpDcaHD936NGv1BYb1kDfbBtC7smEDYWJrGAvQ7K++1K+mcMnX1xpSnpD7T
3rbhE3KjAJdeNLlHEJtuteJsgJctw+/CFLBNlAfr1xxtG5bB6dDE0WWad40KaOdU
vzgLBHdtW222X1kXhzeus+0EARc+wufR9bZk3x0dI6eSg39pzFcsZAI7Rh/AKcSU
ttKI7DxYDH/7Z8SMnIXEQHpxNOCU5z3muz8C1Ks9vZxQhhi1J1cgTIvFZ5ftEC8J
7wvDXsxxsNUbn2WM/+ynPeVrMsGGoHCMl8Z6xMri5E01nAKciC4dlIkU7YsYgsy5
qpkfOoYmeju14LbxeMlEfaaBTcMVfZmbdTJX8PlPYMBYyiJaOZ9kk8EcdThUfqYq
y3KStPsAymnFjGtFevkYUSIIoir59baPh6sAY8w4upabM2KtTP9PLnJlve20nZDW
cpUARSVVHG9z1qgQxQ2zQ4lMbje5SrMn43+fWjOC9EB6TfJv/7UEUmc4UGiKGyGH
sqZHp2gEebEpmP4zBWpNU4Oh1S9W6sQTqjPnrrySUzJzw0sCg3BeNkqseEKkTe2V
Tq88IOSxlPU8CEgQFQZhLkSnuSFdcit/lL27/fWtpV+2UbMUkFiZUkW0O7JjY7iQ
wIKFSHaOYBKpxI8+P3BVLRUYHRtCzSDlrcibcnlpoqzZHmEBtAFoV7lepYwuX5A1
/YBWabm6milizryO8CWRczPVIT3m40gM741k9U/3ndD3AXX8hfWApUMhZMnR0aRp
QFVL4A5aXWXqrdhjlJ+hOBZEBQohT8bDNFi51arsQJ/8bidX/hGBm4gW2CaVOP72
2SgkbzqmraFFGJDf6SRqTzN7NzAWsgqyRIGL2o39TXoZLOwBJNjnHnV8hNj7Fso9
HP5AQEmrJlUIwezZCjGHii7Cd538/tOGWZSYBQFCOrSSk+0IUuO85F2hiGxPk/Wk
IWqpjOUyLTayrExcEnFjnwLNaqbksngSNfzgecEKWvYeqf/ssfUTAxxCd5hjGjK9
RiUU9st3vG/yjBzu35I51hUi51sWAp+rQHwZE+Ag+Vgh+G7KGoDA8c17nezXX/IN
H+O07VfPh8XDYLlODmg7T0hqY+7rwC5goAJtmmhfWifD+U6IL2bapLw64VMgOV2Z
VbC/LHL4gI8N8bqU7vnNKtCKbU3U0hKV59d9zu0azHLuYKRdaTVgWHcovNQVXE5U
YV1uMTIK14qDF001nFYnwaOJOMPZzG8VrfNipCqzTnX4ZIWohfgj10lkb5yGlfSh
vfZziV7y84lWuyVXC65HeOryTH06kUwBtEZfJrbCB7BCMxSJ+idVfS0lJ1Dgs4f0
b8lVbTuM/9QahzYQhJ9T2iUz+Ql21Fust8WMJzFc0b4Cytc/DTL47AM51zovuElR
04rzTX2GZ0JZOo8vGlWCHyF+m6GacD0CB7IL5xamLxUnVAmX7XB65oMr9/t578Vo
OwbUULrpnq2bVbDsOVJ1omRq+UnHlEjWpt1M/O1NfOD/081nzFsicgXipdyFZlbK
6nH+IyfnDCUWHpUcNUbKKgYB3bLLerVkNcnYn9WZ2VsqyuYsslk9WUngvWxP+OKF
BBrlOD//lVfzBTf/EvBvVG8EmD4sd+yPJ0W2flX+79eIoBSwOJ5wCpDOHtbqulLw
d6Zngna0vyXixlRbrpWQpHfdzsP9hwwpNpUGSwD/Z0xP/5ppi2j3Mcby0RGO3soc
zUCdo9Cy18W+ftU9PrGviwzAJQ3kzJKK99ADcuGLqS7WxwlsqvtV4d8S1iSnoS1w
ShzjdUCkdPtQuUgXsCmLrGr2ioi9DoVGP/RB5r+nezxyHAl3sIKhXR2bmIvchRuJ
H/vA+tOKlYR+U8XjRzSWmsedkbeG5jKnIlKxtuSFkv9VIoJ8ivnnK267Jw6RAp1e
j8MfKSlkEHp2zSK3cGUXMcGSjWu5gomSnBvfBbvGvfX627pjchNtRVD19EQvoanu
Wc4lz8SUpJBhbbUQKO0kkReArqkbRMJMBBuJLX0+gPc/eKRkmuvp5mczTfHklPH3
S773Bohrdk1NCJJbEdby+VcJ9jWT7MSvO+jpXF3tHdJzJdvUuSDY18Loc70tZeX5
L+Ib+G4tw7SsjjLiMav8RcYXHNBAnpKk6uDHYAcoeGKXSTh4qU/14EOv0XJ/K/eU
GlzR8g+drx0a9gnMj6wq1gOmOhAajPz+RL/SvWC5M078zVsm4f4jY7Tj5kYmzEJY
bHciGe+dPNr7RFRoH5YGBnvUVqHswhkpbrVzc1ByrP3smSVn+CDFq1f8Rc//kbWR
QvYr4FCjohb7r+AQEEbQWyDuCSTBHXEeyh6XIV6klUYn83N9cFg4Php2fWkaV4Yy
0XvRCmbTK6l1C4URkme5M9fDKvZWiA9Ex7u/cjo2oV52OBSItwLORrdWjt55I5Hp
uEb0zE9xyIO2uubV9riasxdNBdAX8eACNcCAOfdojwIsJLlRIDHU//Y+lzuYKJFp
7RgfyBfy8Wdr7/Ws1b0bLyrwLqY3kD/Z+szSDeeoYd5Fmg9blg/VmrG08QVyoWMJ
zOWFlRv+N3vauKv3oAC9mvkf/oS5XKnNC0nR7OKG4s2Hq+jtF/RwyFU0Gm1mTi9R
inEf0XL9MU63E6bBYLGst/05ui2po2QWdzs89yhjvHHbz9QcWciFKWK4ppNkXao9
vRW4Efv849DOQUTOKBLEvPNBZgGMScbs1v6smBvQdKXxaKwouFCbAklN3DS3bSR3
UXpJqGIGGeOy9Mhe74e3FvpmI7DOtam6eQsRVcbNM+dl/XfU1gvJS8LoxSxqjZGp
GsNNi/GpIe3S9OBuerOo/9sR1ql3HD0CeD3SlBuTifv2eDaWKOKTA2+XMKmN1qAV
opF2TmGLULLE8+024Q68B/OWQB/AN6u32L8MXwGZVX2vytWwjrk2XBTbgXAEZOXr
tCTvsR0RfrprD14s/Jd7Q09JhwlNtoOwzMB4MZgt4Rj7b2vOUc1r53IDDWQE+6an
/3skGLL600AwhvMEmmveJrX0RUAi30PH5gZRpSjBu8F71vw0aPE+bzd9atpJw9vc
Ly+cWMh+CW1m3C5XiYPsv0LvxSj1/1+EkWV3/TxsiLTP+j7Y9rbH6aXTgzwUP3wQ
p181eiwdk09Dt/JhGHyw07XVOsAXmZsOS9oiur2WULLY3BWbhHMmuhRrJDJ1T7Cv
s6lha1jFpNPDGwjl0yQ+r2wkVezVZkLHwLm38qzTJO2R8NViinJHqfXosk7NPFA8
EiMRNQLoP7ucmkeSvN87n/Nlz/0lSt5LvqjT+UTD8quJzmUKV2GXfGhyoCBSQzUq
Vw62RIr63iEYNA6bcudAW7Me1k1yyWL8Vwb2Y/K80LTeEsBFt0F8HtCsFQSlxI/8
bDV3JH6zj0z4KdfQ3Dr9CMEt9pKu0s80KVwqjVIzt3DLE7QDrjRVulw+yTaCR7QA
T3hdneu3ha5onuiaLDhZy4WZpf7ft7m+d0q/jkJBZAw2TSXWdfxNib60AUEjoXpu
WD12vue5pwNfPX0ZIHvVnSzVVDOtBi4vmV/o5fnnQHUWzgb4/r0NAZpt6lJr2vgh
L9Z6Nc/ZHcafwQ2miBCq0bdLRFL4Yutf4XhoDLcPKxohyTuKLmHKhyp8bH+ciHng
hsVUldO6OzhhRIhmhlWI6EINeDtF5EbGX8Glttd8+Jz4rI493orbWac7IJVt9sz6
CobARReSTVt5QweKkEWTId37QBKG88cbQD4x8jnxVPONAsgwMDCvav96XpZU+D4Y
mb7k3roRfHwpSsOfG/4QeDq2Cxx5ZmWb/07BdZ87iq8tmufxZmTbSZcGb/czRM8i
x48hpbmM+PxKxltTYswJCxZocr0x49P5c/G1F9d3VakQMDzYyYlRnwJYMM3yUN/C
emQRuxMF6s+NAjtprcG0+nqTPmUaqwKg2sVo3eQT01F3C416Gi9tt3Dt8yIj5sR5
/Rza1DbC+Z4fZPTWjjSS0wtuv1jX9msNcjNrMXREH5EXVBihUk7d/kjCQywPBrg/
O+MTzlI4TNfG9RFpn+C/c0ZzCc/bVOPAJqyANBD2Djp1nrx2bHjyLMY4fw8KK76R
kxZYmBt4yzJY/J+OGJjKbi//dcDCTfmfIMiozMhRQVPqpUrkwtYaqG8nfxqXPSwj
ZMG3e6ZCG4nmgr/8iSBemZgdsgc3iM+Qm1FSwMPngtYy0r4saQHFgonfHJXg8Sxl
ttQZAF+ArAwO+Poopo/yx1Nl8ZnKcxyJl9SuIodBN4dXvuYADhtte2WqxQYD+xEK
MOQF+xfFG25QacUOrpFwyW6DknkA6tkst56qGyuI+ip+e9AXuJVzhFyzE/wJmSIu
IgNBG35T1vIonN8+imdZO667pFnlqsuMpWB5xvb5U3DI731tKlygeKleCL7PFa8p
X2xAS7UUL3C0HzqPNjPEHJS840r075XZiGPMtZC9J6H0InzTOnQtaD/kJNtorl4E
ZZs9mdC1Xi2kUxLXot4SJtgzojKtWZEGhrdhaYJNBhDMGOtH+ss9BJLDfuMLhtV0
OWOR/YbFUKEKUxRmq7PeIGVY/AGv9gDwFVj6RPbl2D9aig693vlPKoMseX0yWrFp
0b0cqG/CiFVcLegOcRo+no3NVn9qrYHdJQxPR8k/p75TNQ8J5OJowCmBDQm4eQwr
BvGY7H1k0nYXBJbXsZBascRxqJSAEGy8JDVxPb+/aql4CnWgTOplm6cUiMCG3vM2
41nPi/vnGJ/Vu7F6QjnMXUxALBE7sVft+6rP2Q5oyDQMa/GLpNRZuII+dVqN15TU
vzkd7Sd7bCo5l7r2uFoKIIDc6gMxdB7Vw0Ma1U82Q/F8bE05lYRkLwF8bLbl/kVf
7SKMtHAm5MvOQgo0nRaOondzPhKKPchDG89/TQ9Ya4KLuQE/beBTTsspI7g/RY5A
fHjfXZPCK5HPQAzyU1xA/qhHqRnq6QyLF0YX4nLYNNdBFdj8KadJSR0HhTOCtmjm
N7pIjqCM671VqbMtCV+SouaFhAJZX1YquczDE2xByDLRGZ4IXbY5cuh6094eyL1E
/mQ2nVZjdQtw6EkyLPz6egVBNe2kpoq9JHjrKvD0cikxTD0Gswr2X7BaVPvWJiRH
6JTQQnpui/2N4w11j5PAUhdDFG9o5/4lg9BTa+UMRXiXrOcg7I5+P/mxiXBGS1Jw
/c13QDZfDXp5o0fEnhtvd2axaNx5McqTSZ0/rTYrBXigHwXMj0Pb/DLf0nUxsq7g
oDAlU+GXAv/N5fUfCp4q90SwlJSchqeS7GECI3j2dH9pABe24w5aOWnjMWQsvMDS
uHiClYnI+NoOLrak6/1e+3HroXuhyFootjJlXWZY6Cvph4R4BlkRKp7wnN4zWgXk
dYYYC8ZoKezZ8q5XPpbrf3oLUYjO4K9GTZHk/gz0zh3sTFcQhTBsSNkBd2wZzaGK
Ud7RzF7pUzYkvcK1+ppllU6wnYFb4ViUBlh7k9v/rKphp4soemphEZsAjBz3bp8F
aUe5lBwuEtRLvkHmISBOmtDp7+FaOL6stwKkiXv/E0UIfsGOOtcf+jNMfiXa3Opa
ZF5XtRbq9CH1jQLp96oAPXaMQ3HxuyUH35rpNb7fwhQDlxqbeSvqRwaVFNNUyNFj
RoLsJV7KFQtk8BPl1YI53UqeByhLxzC303WZzsNh2ATlkEEMCGizZx09jZo6n5fl
r4uiwYNcC+LY94bRzsGa7b4i+V1WrLtq+Ac7rUKgVofys01rIzC2LeN1Ynl/OLVT
KckYYcuEj7HpJ3oy95QYKDxfURMXkpDHk7itXVnj2XO8DKMpPGkQsXT0lb8i+KWn
yiEJiviPLbDnXD1pehDdtC+NA7VEAty2H7mvM3m48XMk1XKT6p7V2d2EwMz+0ZK3
ddt4D3QaxLSotf7z+bKmxDKSqyYSfwPc3pYuglIj9LQQmLjYmQS8B2/rb/wT8gIq
JCx8+KabFSw4ayg15tz7Bup7wah8jNeo8pNqlBW6T10s2BOIBPNoZcjAeMf0ZonS
7HN8S7jcOmwSH92r/zLzABtLWH+44Ix1fVV2SFFD2zV8FdV5Sw1W94YMWiS0mFpQ
bfKKtdP67xl9Tv6OqZwldY7IGyPuQEk3sX8QC0VvFg9uqe25EMcyTijj9BDPZQRT
vUYgB4iAeQu48rfeSfLnGttxTNDmUAmWXtlVQGCg4Pl/4dEgPtN2volVt/rAm6f0
Q/11QxS5t02ddpqkelPT/HyIA1VfywXDYWVxdXCr+WSBo7Mf25jbeEazqOw7EVPB
9mgp0s5Lr2iWeqXJoOazc6WpSEwX+hOLfITKjyIz+4t8qN/qgne1bZ8fbditCXjl
7MebxSnQJYEpuh1pt2S2uXhf2pa31lcN+Tk8L8kXXP+a6lpSOo9jqfzC2k6mSZ0o
KOX7U3GsoQyxCjNSudvz7n5OVLvum8/AX0zTJHIW6SOrEw3CmhyMrZAmR2HdwO6m
GfDXvemoridBV8ibkMWGvphkolkkEoKR7X/Sr6FTOQop/cpveZ2rnd0io1NkLEFr
aUTFR22A6y5zSEH/JdnilV33xvoE0e1pcJGRbPY1dD9v0yiwJ9FUh586ljH4jJzv
E0gE/es0E7u2z5PxAUnKD/LVhuTPLKIigwQ4B6weB2fYtqyWZ1H3jS/CzpzU6ubZ
r5u5NWn3MAAO2LEs8uR+BuvG2AKyYFeykgA/q//I4pG5F7n5uBE+7TGmfLjhX/TW
zltRkjCqgg/i3rnJxREj/RtPf8v31oIudn7CUq+sr6ZBwUl47KTbzJ34TyHzrxMp
MM+HwnCren7CZV6eohPq5VgvBQ/x4tAUGnBnLNQncN+SDpczNB0apYZl3S+H7VeN
GsWpmJLAHEhiYillcar0gZFEbLSjSLPqy6BtWaobAGt1k+5+iwdn9xNDakTDe0mR
ef7SjZit98QbxeH/940qMrRTOWC+nMYrrZUlfKp6rRWZ2MRQhwnGL4ewk30jxgtn
PWX04mfZ30BfsrZlsfYTas+ZAgfegCky39DUrBHF7fks0fciYmNTvE8Q1GhwUJ8i
menDKL+N2/miPMb1foVhHeZN3j0tQKTjlq/thh0inrz2ArQ9kryD5YWHF8LEeAsg
surXAv5OGe3SK7V+8RLV5daT94QdUNSPoaoFxlCBZTKZqEJa4kA9OvHlgaHbqS23
TLRltgKFadBkcRBhSCPRDn31kHqJQd6GR+rS4ozUOQxZF7pO2Y3ulkucnSO723dr
AmF1mSMYZ0/BOUrGUXaAvvCN+zTDKN7SU3+68MIVvTS6QCaZCmq8tzFjfhZLVSgg
FllX7pxJFRhNQVceosypB6NE7LzCUOAvUcLjxJ4FRqZzZyP+UvZ7DAALrur7Zfh7
FmAO3aAuqOWAKew8T+QdiKLJBefOmqepqz66zX+ShOCyPnR3F4VIHQkka2A5Vrv9
0HKiJGeSkIkDUligIevGZCA7qOQn1mMydmXnBsKcrVvCtrXR/orN7Z5ZujTgZLXO
aKIsYfnRI3Xw3h5iVu39/eWQMGPq4REV+nf2IPiZyrVzl1H4TK0glY9XppmgQYNi
mN59OR2ZC2k90e6K3C9sZO1M4prvqCNs4VKEPtGzVO43AbH3AGzo687Wnxm2q2za
R/xWuMw8peeDRSfgIYXSZezbNs2CIFZMCogDDYag6Ic/2uJyJ53kmMmIgghCqXkI
IR5eRiYaidwBPdV0uKGkpVjuQU/8KPmobeswHq5rBYHGB0xfuy6G5+/E/fDQk1MS
rh8CKWLlpVx9T+ufsrdxZaxejDp6G7YcdAtOsLH+LlUef8No7nsnw8+iPkVMU/2d
8yU88sUvAlKK+dM4qkGqYvnObJuCnkz9PSobSbxakiFBJAdEvqJ3QDsL3Vtat4NM
ay/LDcASlbVcXU3EbPWChjdcHMlmbqc2qwu3DplmLagzfEnNtMD8dLjgrBdZqMQM
+mExDB7NNQoYPn7KPL/t69pBZJQu57Z4kZB9I8vblrrK0wwJTqPGA1794EhYq9/R
oLYiSdUVw4DetEkfWTxUAtrD/1IbFvmRqmC7Ch1pmZ7TcXPsvqtvbtVpSbUmER2s
41oLWTdLAFGLWcmuUPc1vhOS9xWg8gx/gv/wabXbPfQFYRORLqdkKu0EC6eRXRg/
eMiVpR26ORC2hzb9DHxzGuxg4DUQlW8IeCw9FPcr1WvLQ4F1VypaB60gMGVumTuc
IUl+lwCfAleSoAHE7aA0FRVQEIxtx+XsBQWjHG1UYUTa2/5yKeNN+p8owuVDgbHi
mdXQkpdk71bIwAPNDW9Tk+/dyDCNmjtmSzzp7cn5nW7HB9DJGt+dBLsoICqIqcjF
VADZOgIF0TKsmGmQxgCDSUI7zE34aSCSSBEyzN3yQXP7EKa6pSYSUCPyBF+qsrwa
DinJZEOyj45asR85ubKTEIG0DH5duU6wb3TCj9fatd+P+McN7J2hvPgk89XQ9wCX
0hnv5Vn9y+5NYklbplmUNCjTzny5X0PBZbQIWZEqHD1zopPBVieIf9jaITmOLTq7
0Z0/F8uafgR7YL/3PgtLWljnfWEtVtmP4YsjsaUotMDVJv7MNzojpOfXFg0K8ijE
3ULNyFTlNmnwBuwBe2yqlgIyLorMqL2a0crv05Cr9P3XALhF+vdzwcDZ6Ps/tU+B
exf1KvKi9+CmfhxfqbpHeK3/f+bdaVj9EP8YKL/X5HDKZFErvAOe7qcLs3zSS7U/
mMLkdd9jXSAW5/SK0tsOG6S/pBJjtSL40BU5JnyzLNlU4K4OLtX8JLjsl7kmHgYi
P45i9uYv23VYWZTlgtO5ILH/EzPeGXl6aLaDUKmMva2W1Gg1n7PYzWc1grylPbpj
W4OVocO+HGrQYWlScphD8jW6mbUzD2qKOEebRC+lXHunPNw9OVKEJXbBrmrUdLZw
5OCTbpgWoaSLwaGb8AwSq3pOdBEwLAtTHBwSoHvj+t+oX8hsgrzl/SFsjXMo8A5Q
5GrT7IDIzs80LfVLk23IQ26mOLi0Vk1LEzNZhwePRxFGUrQRu7vJFMnFdVs7Uh9p
moifO9eEyXVvHRrV8ZpCnDjubpwopTBCFFgBfQEcLBf1+t7XEOHgw7jGkW4qTBi9
Jt3T52vPnSGnSK5DOnMwWHM7SCQJ3yiq3IEtDCIpjKCM+4T9BaiEbcqs8nJPalxW
jgM3+HPt8Yy734JZjOLfkL3GY3uSh2vG2tdm6WLByYr2N7TVpJFKtG8oRM7RetwJ
DK+NFAkzfyfWQeXee+geEjOqR56N9V2RoGQyQsJ0urWnOP5DbI3gVAwnGmT0dE3/
okECrijtBn3GSWmuAMv0bEBH2G1WKWzdAJuECX0lx+1ugFSXY35lScxjBUfj5+Ms
6V4WO0IidWO/p9BZII4G3vTgEn3I6Blch3FJ/YoPDNlveVagFh9PEQdp8ZNb2XEq
IZ1lNjtBp8baxKEvSJ7pcyIFpK1qzVhJEzCfRcl+HgRrJ23PEXH4AB8puXr0aWcN
Ap2GLap6oXfsMFwAo9fLx+10L0oTD+znYtZ47kuajBf2smgWJHdC/r6ZBJhN6kb5
9MGVXKVvIESofKB9nJniTtTRnumtmX8CfootoBGw2XEEpG+ZZyTZVrsVUGcbxnZn
Pi6GDyHHMeanscbfCeY8WKRoAKmCdmkmktlFTYvRS5r9tzeR8isXRzUR4QiXz4AQ
kl6UM5XES2ubyRaVTLkBQ1w++v/G7IcvZeyrHwxDJEYvNI/BW7JyQFgyo2m+wH7F
uEKd5/z0D8QqtZe3GLP4JZbHZANXn5jiTp7zTbZr/12/Kz3F5Ywo1eI/K3oWTrQX
Jr3nh4AshxbHoUEqd1qf1GbCNeBGnlS/z+jLGpM4jWHj07g6iNXCbZYEipy2+CGv
SxpwR9WmXBA8OJvY1QXhNwKZRhxAm32wwEOABY8x3Jr+xgEXwR55Jzbnf3jyWTUf
B8weCPjhida7o+6iWuDeDYcaWdbXMoaJxohYQ1kDGPYt0IiYTAyghQx7Ktp+nBmE
ece6T5ZYlZLPO5GU6XAN6ocaMqu1biqHblG0v3WZFv0ZVCE/l/xd04bGxZQyBD5K
JaZFSl2pXQPyuethxbV1CxdCgP89+LUNNXO8Bqb9SUNrbaHwj6eGRS1kQxFJZedM
bWcVfjgtxkbROv2avd/+g7D+2ESDhD6MVvljpewSYvSAD4CNwLV6V0JEZySc5taG
1ZQutpUf/TsFy33fCwNttmfR+Xc7SSqh24U04YfLkoKHKGsSNp41eheIpcBn5xYX
ob3ctcK1JYbEgnN0KG6ImOh2jjny3mX7bZowUhN8LRZFATcUcOZ55HYGl+lblbRu
yYQudGeKPSk4kabGnwjM9oNnnXTP7q+RJ2HFi5j3mVB4sPfcOSjYpeFkLaqWQQEH
V8qD33NpJPZEB9yqMcjP7ehwARF9vfmktt5joMAy9kilTGVyyTaE3ezsmFlWPEmu
DslHm8Lqkw8N7rnoHmXAvjXhUlGrbRnqEMrK4x5h/dPCrXZ62694XfgX9KLsjf/o
6tYzx11Mtejf8m0OZ1EpkIQIKxEpI6p6c6bHhqTfqotVEOyTvmdKGq4Uc3B4pjjl
BtV0hx6lsg+k9T6RZLzL/+ESHs5UiYIqhDIHx8bj2k32xLmOIDfE2+twXXt9iR7F
N5b53kCpm7QqH1QNxrvPgNrR/RKkkbrIuZsXF//SBq+m2DWuVsg0hJWBYy8Na2DN
+9EK60v6PgjsJ7LCr7JKyRYUQeKbVYoGX/Iwl9MH4D4MAibebY/BFZrsNY5Pcz5j
2rrOt7+B7bR2FLKOg7GeY4j42qFdScVR6fHBUjYA43Uhg0NzprAlYthrLvLK5BoI
rgbmn+wqHfShzsDHhcj9/JQW+t8yP2OuyDWhAUwiYJ5CQb4nkdpkWtQPPnlUcy35
NCtKorP5kBgfcMDnj7Ls8+WqRH+oKI6eqkfaRYILua99R6f/FYmcWuLK+qceIbPG
hMcVMvq+gZfmvUogmvQZT7ZN9KbzsU0N0JA18tHkys+omQQkeEj9nEUmyJEnb7ud
M4XIrYJf2UXrHMHqAffUHAe8/sDCIMn5ZG3fULHjIO+y3SIdE+qATAh50P6fPfm7
aM2qEiLPr37jNobnmJyKprOVc9BWiAwnqWDBMdTgPlp3C+7qMgSGN2DgowR1BL91
fcTZ1E4Wt9vEY4kNIdZMy/7zTUEKEtOGm7HRYRuzSS/yvWRQe3yytzMYdj/63tCy
R3RBG7wVUScrYBPnM6JK/p90uPxMNs5/+tbRhs6XMgjKJRSSI/LrofvusGR0ULG4
p4Xq3EyhQH2cRMBzLVQhykw4XTwNUmxtkkwV/wdajvrxleTGg62BS4e0Qto/24g0
xJgd81bZzkG1o8d6Mazk7id1b2p+DCosxJz4tt1QDYyMkadu+GE3KayZ/WedLQr8
7A2yWmqWXsR+MAdzNl7Sb6ra63cPGFrVhNr/8gA9bbNpKP1s73FW30KN8RoZHmkP
8icPLSGk8ZPgn6oz0nrgc60h7ootQN0BMDbuYvDal4thxhGmFZCu+r0QNysnEC7e
68mEaTfvyeQ1QgouiKV/74p/HSuEggt+vG2PhSJAs3YpXBLdfa0laxE4ARllK3gv
34xdnV/Q4fTwSReXnkZIxZ8SKEigrm8sA5YW/l5uoyUtOpeGz/Zt1GJh0hYlasm3
TZAYo/ByP5p0f34SpexO8+DuPhMk/oavuR4UyG6hcRKco0qxcGQd2N67sPIzPa3t
3ycwJAeC8N2bkBuVMluuzlKCK3wGENwQ4pnB01v4g4wRvKQq8xYmlwSwlFoXdhZC
ZHRjkrEORB2E79Bj4S3czD6i3moihe7Zh/Mn57GZJPV965n013SaH3h1QfAjrMbE
gnCk28+H1+sKsTLX0eKCOg8nBz98kL7dSdYL+WIhAEPP8RgO1zbabxaUW17itprP
W0t2ugt7ho3U5t5aokHx+/qfoJx8m+OwRqSgjRcXubDC9Ukzuz0hGpfkLWHK6pYu
8Cz2pcCzG8rFLBUBpkQcxxxsY96+O2IlcqbeJNWDjfrNBwLowBHz7AvPpsvpAyCN
Pds8vzO2z2DE6WZE367mITOnVZz452VbU8YvntN2ImAUC2YNSzxRPfahX0PCMw9d
ZlbZp3LArKGH0ffzq77koPABjUY0R7HA5vgBkp68Fwiu4He+gTwco6mja0ANj+bN
zHajmn+KVmEvcec+bLJtIvo6Fe1a/g1fn3InNu50ypdY5cmSVyD36abGFrQvduXJ
YAJpvMHNc7SRldGwsT8wBJ8QIAoYeSy+S38HykavNXnmf0+wnJh/q+Uc/dmU1Qf6
VHarWBJf0yckVv9oU7c1hwq9RsShDZq2yTKEBb/LnADpqyn8YXDFqODcAgw4ApTq
1/dNwlBsIDH01Tbo5GBJS4Onoy5sUwp5cwyznpjes947NgEdBSAXCHTfAr2QLuQm
ZDQNSX2AlisX0ZMyetf7le1MZhrCWWbrnuiBUkkfsCRpRc/Wbg0m8MvdhYNAm+5f
/hQ6WJcaeleQCn7G/rG9tZP72Z5TRCZ0JzRZOV423DII0IehWvKQk8W3u1izAoxy
5yEYpyBcT2Zs7sUAc9x8dOtMQt0yXcwf63vrocszDOmXqORzdced8N4k7FBHeQzt
CPyQCCUkQViV+/BDubyDbQJ73uF/+fGkbbS6RbYX4WpP6OKggsFAKsdjjqQ+NfGM
1enazoS5pXEsDdiUneW2d0QrXG87ee9BvOrt2ot8Y6RE7UmSqXWgK90rXQPxvOJm
GCxr/wcNu6S7JmadQtJleWqz/6HhQ5uiI3hb5PkqI2MJ2w+YlooNvar/c0WDCD3k
TK11LZFvdUL2NgUulBzneM6nKJ3OezoJErIU4XdJeAdMjE+/K+4BqsGvvbhv742t
2UUM/ntLI00oRSwdPKvVbHJWzQ34bs2p8t4Q5UXzKH4gW5O2bwnF8MoHUIPiKiKj
/Z7hro7s0/DJFBfmtPtmRM3auk2tQf6+hK6lawQK1bSgjT4YUQ06KOqekRBZEf3U
YJgezM+YOdhdvSwTKtYVR7gd70Z0crk/KYeKkKRtjsM3Vsc8Jy63N2YtX5vOuqt9
G8EKuACIOogCPfwiHmMa4lHZ9RZPBrxvIckqujTR9lKDrbWVpg0ne69ERxJ4Btgn
WJDUAEyfc+2J0djOKxo7Gl6jVZSUAmRXS9pYqmjMrrwTO/OgBJg5t9KC59mXxySC
JOz6iRMdk5sPA8qY+VKbOXgl07t3BDOo2FsLNGmiZuBC81XFY3HVndq9BsxGrteN
htIhdkNNXIZ7Ub2yypbQWuFjkMU7Etf0fVNzOIg/3qn3VJHhHXmmf7Yy/ddluI9S
pfLIeKN2eR21ZP8InjjuTFhyBuVtcLJgppFKjTyyX7pYrpPT0ohUoa2kERuEf8er
sJZXPfJf9WkSX93HQAf6wnMCJcjTTRzD7hxVLRbJ2zmdg5xHkbVg06m1M5AvyqqK
bgMr8WM0Y683JAKQbi2AaHb5VPVhlIPD0c6ZinQ0RajjQMky9C2TwUFqpjT1f3mX
/YGyCPX500FUtwJww1EyiyvHSi2z75s3/bM/4c4y+S1BInD+jwST7ouDbUXsByVw
p7VosxsWnqCGEOJP2Jo3wAvIWsJvEBpvHS6HPZKkPP6fEyoo+ZxYltIfdZXLnouu
oGIR2FfHNTQss9a/pIlaG0V+6AU/YjZTXUOoSPvZcgfdrc8uuMA2a1hsNo9ikeB4
ntaFxFRIrlkyXvBGPy2Sv8XRewfvSyHGLEJXZ1MkE7Q3jE0e+QESMOh3LpTrmecA
/NsHEUJH2l+jlquwnu6613SW/WVfAnAn6lNYMO16jrIsWcKeFUvLyOgq4WIjPPws
jP0AKfUarhDZFxKaKIKR9PYVztOtVkq9UqDxmXVXmNW0Z412I5/K6pQ3Cx/c+gXh
hajbUO4AOrNnJZUEWnMfhPqiZwj4n8LuUyNiNs4hpK+gy1PAz+SDtAzWJNxFi36g
mOx2M2deKdMH9kQUue106uDHEF9O1pNDqxt9p9VJjG5+8EYY7jIOnmm5tuDL+4yI
ZsT0UV+gWVfd3fMjhGFbivQXAWBApGbsFw59TS52Ulb/AShl6qmajsj5r1Mi2N/H
o9SQAi2mfvYxONdSe2pJ33XkMwJTlwwAuD4P2Bla4Kd4mJFu55oWlEqDugYL64vv
EB2C1qTEcoVckJ+dnwCpd6gRslmTLNA0fuMPdbQ1NbUN8LFsBUaMqrD2t+t3RDDI
WjWttrDSkDCfBNDKfhrXLV6r+muq8MBACiZf8khHpOkpMPdEOHnuX9Nn9r2uGabN
8gX17f9HfsAMgo1h4uCTgCGgDcIWlooH7x/SRuh44IYUjGFEERsFce+04J6g+xGs
IplqIn14WLOgjdReNUXFtOHIIWoMS9ac4m4udJxkufE/lroiCUHHjtnybVHKoaL4
K6a+cU9I02DIhswXq8LJYkn+GkBcM7FtCfLmc1sEKDPXehYeuHtsioekI3VTOL3w
eGETdonAScyEBQhUp/ZP8opfXO2TIJMTQv9gB1cagResOGVUJlV6kfqbNkccRSUF
A+As9x6e5Q+TzWaq1nMJHCSU5cdLW+H58U7JWeK38w8+McDkzD/Jj/sFK8bFfqcZ
dqDUA0XE9Q3uG+uOwYP1fwn4zmmXPy+Uvo0UfqysnYtifk4fyQ88vwkE8UUCpOq8
5HKh/LEp0ILIqGS5O50wAgPVpIeKAkEgmypB3PPSaxnaP48w66JE4GjWItGubAnH
TNa2ytCvCqQwfId6cbfdX/jQMzXy09iNxO63uOvZy/7wYVbotNRtBgaU2ygP7jrD
M1b5UtTMn8eex64jOZIHhR8JTNUNd0X/MXGe6kRrBqR6JofD4kuEWGJlETm2g1Zu
QuhgGLwxLc7hPssgzBFt2k5z1ld6Ae6UvXFj9Wfz2s8Y4HodIdBcYFLkNyFH1Tsn
d37AK5ZKDnIRS7Bu5jlYPUuitll2vEhhDtfbhU2cyMYGDwoop7ypAz+laAdMtxB4
SlP7ThaItyRwzNJdWRgBaD+ipep+cry/RHmL+bLG6cztYOI8qj24FcF3hi3IpPtu
qnzPAx4uqIX+MS/TyEulFzw4TDbTvmn/z2X3xRfIxPmNjBEz6zSoI7odENUNAuVl
0C7EM0N72lM0nOV8n5CXGrG7Jr3Jxw2NTSPR+mlfG5ZlVic2e72tPVNU/Q4To/SV
1fkcI6xlIXONgi8XCZyYvpNbASJVocp12b1t7KiwdPGaPnvKB7Z+Xs5o97/3BPYT
xJkmCyxsxYwvoS7ahnNulne4r26tgAX8lPpSjGWVSMVROZc+a4GAKkKYrLfNB1eL
u8XQSUtkclHNAgUXrQ2Dqn/Ycpg20v6Vkf/zI1XamgLo/Wwd/g2qBPI3dQBwU0BE
sexrRp6DCwZzV+IQkeadE+trfPmew2m0vIKnGtd7h+nuPMvaZZGh3Qvx7cWH4izA
H2vIYAK6lYiAR9M3PKFxqiUfR65MsoFkKu5FGnvh2th0rIonhbeez3vcg5vE0BMS
HF2VsZy0xQg1BNhv4kdFTz0X8Xam5JRRS9sV41VTFsS5dP2sUkveMjEzStiGnfPL
w4aUGRqUx+pFK4apJ63xBO9/t5TxO52jQ3ozShB8stNR39xWbBT20Rjg8jFseQMp
Gqp4d0wl8B9PTNfL1yJrw2x4QH08RRSkR04Pqfb7+5dB1188gqhM2Dh/DSdaGare
TrPl9SsIwQK5MJ49cO8pjC0VhTnWFc9CX9LXa+GEL7sDRf1hXpi0VAer287bZ2Pe
7EhlZO5dPdLybavivWQXXWP26ESkI3eG5qIuqccxyo30tl3A2kFrOvldGJYLqivu
e6q7OyOlRD1pjIf+KWZoiOULYfPqubwJedjcHaYgWGeLLrd5OP6U6eaLrfZ5sxtH
Nh6/eV6QAGzJaCBWfglUd7dj46x5MWZvzq4hdD9apVYdLwQ4H9uo3bTDVrqVR7NL
KnC6+wntEAllMI1q/L0cqRYOc+QeQlsMIDtsFq3pIscF/yYqaVgVmjqG7tYu112c
s0azEoiYokVVU85blinvtRKmTtywK9mssy1lG7zuaXJ0JlpRIdkPXbFKGxOmpACV
WCxkpxLTtoBn578Vp3YA9+eIxLHCAlWrk5BdMXwqVRwWUvUTM+hn6irb4zaM8M3l
r20p40Y492FYpvPhH6vFRoB/hdmXIBxRhbaorFhD0wJ4xPfNoxQK5cZfkh0XkNjo
lbB/LMFTegM14Wt99/fpNJthoNBbl9kSQvTApEJmE1ixGw8+7PpxHsdus7JaFkf2
RIjzNUND5Y5x3Z+jHyOt0Mwgm3W1yWzvDv3DMwpfrayVxFbX8i1fxIlmkq7oAK1D
JlEfcHjxbw4BbcWeUsQUbIQ+Q4qaM3HUNdpT8vBL15P5QU7ESHzm9LU08aHm+GhY
x74y1Ks0YUQiqTba7uLVoTxZjo4OyjJ8MP4Mn0uq81X01fXAU3VacS/oNKCxRA0n
tjPU38FNxXjCFk1SQlWU6+9HKAqgTRvVM+OJoUIi+X2gIJ4Xo/s5P7uE9OpEV+Kd
TC+LFHWiio63JAwqxX6ocG6pNO0dijFQc55spRCdmsOoYbePkcdQSqVGf69jll6Q
52SOMJ9TI14I5V0seFKhSv1/VuUaBHj824WDtv2K2hjrhW3bYAT6XjoxBpDXoBrj
64D19hDNr4motVeBYEKppGE7VEbY8svz5wnUHHJNAAaStcmrHVxbuN0l+UkrGmPJ
3vrjlGNhBQ3S60xeEXHGTvnHzb2RxrC+svgDNzJW18Z0sWcg3LBAAJIC3Ub9qEtb
Hf+LLXx/A3bx1QltlLrXx0qIsQUbbzG3A1ch4rvYeWANRoxbSO2wYaLqojEfiAL4
cI1fb8tnUeYUY/P7PkPEEg3dRG5IsHKnyCIbe0azjjsxNHFzQDymfqEHPraYtva2
KTVk6YlfbtKEq4QFikLar8l6gXjcnh3DcgRYgvoOAGkLRV63qjKhmFWCr07P88s9
n3FFEGQdI4JTPUGE1dONOYG268AoUfLh3vmBfwnqAyCZ9IqImrCcKI0a4i6/Z7PX
yGgHt66u8g4hCY/6s53PR1WC6asrSwKH5LBfCrO5FXh2L9Z7Y8d8ngV3vRl89UAo
Rz3XNk7ORtJ5W0yaJ4l/1dARnOnuX/CqkyjVVEBcgVXgNHVDccxZHjbuay06vp4t
SDhz7MeZt5O5gEKyfKbzhxEUqHB9TiP4IsLOy3pSPy2RHmVOEUH191GPkAyYMCEr
w85WoXJJCz1AsxDRI23qZV2+sH9Mid2y9+hdNxi1N/GwxKM7BgveQ6GxRJSIPTaQ
7qoJoSAx/wSpdH07+y1phkyJKdmVNjeoxcQH0UJIcba1d0W1+NJfLQ3MsPpEK+0+
oYI+VNNS1IJQKks3hdMHcFVsziy4f+9ceibhs1nPKuoYhtLeCt3PUoUK5nP70XAq
PxENojgLfI3yrSEb2HmWRI7XGxUBvggGlEqackwKQtsck4k2hp67Mbfyh/d/yMJn
4jpxtUfgzOa5BLxYXzBjHrUjo/xL0LlWvhVK/jEnWLUr++/s9zU0eGIAOzEUC0ZJ
ofWlbOPmNfzqIwnhNO6pDgRNJ5niWqQo8XgiKw7uBg31fwad2x9Or3g8c4EYLeEB
BrUDg3Guzus4J1XGu4HLkZmrAHD6iyKXOuxtqfJS+iYV+0VwGjPwPMeGWnS9hmfV
Yonq0Qvyp8bDhAS7yltm1URNoDuQs/1MEjnIzDQTkIj2Gya7kf4SKth/xx4DS8W8
mbywaU2qfVpy91Yba19Rs0U2+Ssg1xTBUkGzg6YEOTr+sv/CvaB0rYKeS1Wqti4f
4C0YK0BydRZT38+hQeSM34Bg8dJkkGjMXzcW6j4NzzFD8gvu8agTS8PsvmjAekts
JDvN3qIiB23Gn5h7jBypQPmJ4nI44H12+AKLWPPx1RjyJZcjklfWCPp0t/j8SlCW
czkYGFX+q+pUfVzFpFZNmXk+0XgrITVZZXZyiphu4SivUh0qFaKMs3dMAr9AiAkk
65y7gDISdZemMZYsgy/J+h2zKsmrv+8o92FDiPyi/ojHHRoUC4DWVr1ts/ZymKhS
SPbGjF8jgqip20arJUlfkzE2Pb7ijHF2aH4vsASC0hvTgVHMJAi/rgFunIU5Qh02
eDM4YAA04R0Ssn18RZBzWgOwH5S+UVlX8qi1jIBNw9bWkjAflBjD0fwtGQIeV1k7
vIKAmTWV3dnaoij/Yrr3FPS6SztRuafrA+4f/e1YLp8JClNR8Ltbi+ZvC4t4MgNy
q04d0GYMAgAM0HnCuYQOp4+/n1JUFsvaCLVqQ5DJGf7ZLLnN8EPRa7WDQ2YfePyF
yhF68E2J89QcMNo9ntjVeDJ5KtDb4fyzEGEdDNv7tfiPS6pzk5nLQHGhSsepElGv
z+lZF3o0Z+AMqLXIn4wiU7aBYjYWTHQER/7UKawXeWJ8p/OJyskMoYqdzbvO5Swb
fDtj2BH2F/vXc6MMl+BAJbnA6XZJfPWV6xVULLO2XDDxlTN32PRf2yaCE7qc8h/V
8ue9sLwqmsKs/BjuMqxYBlNMIyUWkCvApZwfsiuubrilgghGCEDpvx0zXz3DIA8n
Zzd01NGJX7gZIFnY7gSsNfAEPfeQCeXG6BczKbRT+fsUL/93IEecVYNTlveXPog4
BMu1Wv2Ct4hU/BbLKHuIlcf2+TKPc+xeWeNKa9b4BaOuTSf3H94d7u3JHvtmfLRW
tLzcJSwWoYUTn4agHxtn18dl2wcLmZMCfnYCLEd9bAbrKmESAthtFvKnU8F5BOj/
VjsZhhVFb/rF9fj02C9x8VHPMoYDoLRLXhi/2YdtzKLzIFA/BTAgZG8x9zcqnjS6
V2XvSmnOBUPXu4UD70DZRSOTEuD38HqeP6QGjerqJdZ2UPtv8CF0fe7l+Ls3fjXc
XLe9Q03HJBxBZ7A9/gV7ajjErVOmI0/JUdVzcP+jaEYePH8hmbvzW0Mpozo4IR8v
gxNaSELYprQvRze+0+mprEqUnIBzSkmJ+NaLvR2HkeogKSR+RWnvFQxm4Y8FhtZ1
rTdnzwlnXpRHaXD4Kloplw39QD0qEEznCTgeoENZJo89HdN28y8A0VspT+WwoWWz
BkQkuGfuViwRPIEXyIZTZZJOCtLEskScucn0Gk7UoO6U09945+4xdLmHqEO/9ecv
aqCIdbA8pfxgQ2NVi4J49OgBwMylqXg4V8cN1uFv4r5IWDKNvApQxY//CjKcWLES
AhU3bFa1i9EG80GhSjrWSOXic5Pfe+phA/bgCwKF37OmSvf2s8NEcCeTUMytmkZh
6w51U2BafZblA2PpvnrmnFqG6BhZqpw0ngNnznFE0DrhnZSIcHO+eSOSahB6EZim
ZOSttiVbP8evYPfGtXkNhmhqNRV7bLO+dKUnmlI0MqCuJaDVeK2J/ak/EzarThkh
iVHF+2d/vUV1fps1Uc+mjNY7MG7jKwtmyocHxIZ27S+jkAo1DX7kkQ8W+YSCa9op
EwhirM4nno5hgwnyzdkPkOW9TtLgjctce/d28s3oS/XJGbD9CkUAApXX6r/Apg3F
d8m0PKQdkYMxwSPHUmmAVFfTPIxdaR5I9pVd5auQZrD+jsYhA2gSpWOR2AA3MMUk
+zHjLM1AOMOjEGOX/woNrnALsBl4IEqgU8RRMuDHKJNfF4lkd7bLYufBA5myNaRr
LKxL5a8dyxK8YCi+jiQRfurW71145y/6L6jaAM5dko351Ct8KUAYGtcMZf9NLe6X
HSphRWh3czzgLvvODet2RqimA+xa3DBJAtLcLN7XmVWxT5UNYOlA5qnpX+9ofVVK
YG5EdtsIrPzRwT6MNy16SnAf+DIvGKOCvoNXdRCoIjpd5sTeEdz2skqYwPXs994p
2gbw5RlN++3sEfuFstsiU+ZgES+/LO532bYqeQjs/f+e4+u9o0toEftG3zW9jDgp
/N+jvXqYjbBunjVjIFMgjO8TaQ50nlP9UUTFgqbMRaT0/s6nCPxoJkaiP3+UshOJ
KeUN0lJZvtuvxahRPVa2boTCSU98A2HiMM+PMOfMATkUuUdqJqpzU74RJa93BHdj
z4fADghSCg1CRmeWhHsECksPaE0P8xxMyJVqQaRSQ5NAx1GwAeM9qGKDaxzVoUDB
kiGUO72FAAo40n4605R5XLeREDGBCuD63ewRIhwhINkrTHDd9tsLjgmLEFKkZI2o
3RaLyKpgl8oLISkGYmat19XG0WWcCZl8qUDmW+mQ8Kgz33sBixyxaHT1MN0wGcsn
z3jANlDNJ2Gj9RqkHR1wpjWhm3R908znJEsbSzC8aOkAGcEmzrv+cPmSrbYKFZmx
z5D1wb88QH4UXV/7WOftINClazXckVrHZSQJo0NQRRP9AJVw3E8u8R+jx70VFOKh
CywUp45JqvUbh4r1999M2714x4oYsgbaZ2JjswqgOYimHyE2KJ+EaYplKscZTouc
llP+ZbjmS/XenAeYWvAV6Y7z71mET45Ir7pCHep60jeRX2It0xAPpMjoH7EOc418
Q1LtAghxZ4Gi2Ph3V5+jUJ5zjzWTmzQ43ilCgJS7qVWjbI9g96leETJzmaeNZglh
eKp3H98Ff27DmWoQlICtacri3vFLkU95nNQfGWugIdZt44vG+0L+RU8yYiCn96g9
u1L5R2zBjLOIkb8LZigLtq94ZBt2W9xxWlcLSABEcXSgkh4AsLz+N6kjtOR4TeWT
xhyHSMDdmq59VbMfgl3LNyiiHxu0Q1M74Nhab/n53h1+ehIlyB1X/OhVoXfiofcO
dmwJNWiOs/Hht/KoV+Mzk9jAwYiWaOwLEzZpw5n1bzfBkBu0Ycuqdqs1aAUeFAOW
FtKV5jv4WNunsWomW9do7WNiSTEqA70Ojj6176mnLRIOO6024bLsxLhz/vs1YzeS
vgDrlJMy90fXxI9qNnp36uYv6p9HFkovGmOHYfzpC71uJ9kMBjl0s8HBcY5e3In9
2IPcxNXgxTExuJkFSi5lPcei4RAUaQkb2qaimJ9dlToDl8WHpmqhhsoeeBl662tX
h0llnJRpZFXDkK+zoGFWuz5Pm/fc0PEwADjyDOL7g8Mq2nQ06QY4jPbAu80GW4Ea
Pil8jeD/JjZ2pE35TYhsB88wKG4JZEiYn1+v/vA3/deiU4ZKUFY2sc7PpmFbT+Tb
cTWP5wTdr4YP028yfdA4dbnBq9Y451GbWdb7u161AsW5FPYcQFK4Tak5Si0v79K2
U1rtq8kN2ID/T8wPwXaqcLScHQx1BQ9nEstwko9GUyxtr345PPf/wPFtRU/6wrRP
c5rd4aaFoJKxyiUI0t8Kc1uD6bDDC1WjahblB0/JsFhSL8Gso4o8XTDE8Ii/JSi2
4zQ8kJnYQOAPDawlzCafcPpqQ2tXazspZwZ7Jd5vZSA0u1Nu7AANqTqT48j3W3mz
uwpzIe5LRGHK39p25gJkrAiJ8I9Fjw9K6MKxxlQP2tZaUxkR9J3tlLxh7s6YUynw
96Oq49kCNl/L7+BZpgehEhQhGHDe7b/sjP4tBBcdv6PenO8Ec6AueeyN5b1pjzbU
R8NVQv6LzGAtJ4JHl39pBYEL5o1lxd4cVGT4PODULwBn2E2Mht+iSCfC6E+Mtr4c
rVNo+Vz4iJQ9vafPUvB//4AplEGKjz3rKnGAwXa2xNADmWubEJY3I4WtkzSXH50q
0SoHo4gi2sRxGIHDWtsVmiyrb8RxE2b3n7AROEs7rIOgjbPmmgfNy+jUrErFxhZv
+0CRkkXHiXseBSLZMRldqCQZWOiW4HbuTpbK54rR0naVzzezPzd9k0PTq0GThS42
DiMSQJGQr3qpwLbfrNgqu9pkiPDT5av3QeG6tmASyrJLgpJcvcrSiscUFz2mOt8V
KF4vDMu/HWNp/U6KAMeeYpzXV+hNY7h/hcn1lqW0uMa9xNQiQ6ugu4SZKhDAIvLP
rRO1mGQ+TisBiJGNDDljjdWQd7hdsQiBmmDMmzRqjBDKT8ZtzVKpZBTLeSkyK6Dk
iT3N92+F+u6xCCspQXcNAG/qxBLWUVPqWy4PwP6dMiiWVtGGdhprftyXwFeYquIw
DNcgPSy8rV+HaN/YnpLjSWLb3eXTARkLeftA11n8ixFvIyv/gMhxS6shOIn8HrlM
cZSQy1HQWxyR8KnNg10VB7Kz2TNmwgyUQ6ATzDTz+8ox5NizFMdkmZHiS0hQ4jg/
/A2r7c31UurFowWBQ2iPhnQhmEIVvYMxUh6oE9Q5459PEWGEXbYV3DKlzlCGrm2F
Z13g4kA6G8YYlcXCTtLnJTuWHgPMaQEb2NVLO5DCpKpTo1JlDgkk21xXeq2j8RAX
b8JnNMWVZjtcnYlwMtA1yKunvSd7nnx/by/vt9hC4FitgRRNLJDzktQblRusOjTS
ZylUVj9xECz4iz/QSvey5HxcfkuCV6ZW/bQQ5a/VTqAmrRVYwJ2jX1MLQTPB/iCK
fhbIRY/HJ1MXdQp629qDBhFFMztgRRx9U9yvc0CaN6T0mPIq8iidTxYaHo31G9Qz
UkNv47yytmZOpPlCvik8TB7yeKDnmbOKMJM6/ZNBtR588tqUSdPAwY3v/kUlID2W
jAPw696KT9L3acEMAzUj3tbG2jyzYkP3iYjPLTPYFRufWPij9prpvK0YyZ18imZk
+ofDXIrFJoOIwLiBEqKQHdYj/JLQ/HpzeTLV0N9J/3mWaNKKHaM71/HLltXorhDR
Ft7FK9UIs0YCWdKyjHWIffufnTuk/lnTItOgYZAI6EA0kACq/wLGh3Iloc4GieR4
p2kGc/Si6MG+T1gO3HVUEdqa/H1LmZ014YGEN4X4d2D5GJh685ASV9o4RB2y09Rs
uy8f3RLgxRctiIczgeYDWT1xF/f7Wy8dJCOU6kjwk8z6geJhLSaodh6enpNjuLqq
5uJAeeSQbTjpwJpG3cVHssCTCn5roB7dIbTpZMHWBg+dOxyJsjtS9tdmedlbWsLp
6iBqJLjFpVIdCsy79byWHnMxQ48uUYbcmTChNZghM+G5iovpdiCZbeNE4MoOS5Pb
3xF26/+8nzxuBnGj5lmF/1fpZ9+W7XiumcyBOzqWOoD0hk+b3uQ/svX/HbxU6YZA
HeX8FhtP18jBev0fRXj34cDYmyrhUjqxfOKxGCDkHAzQONi04uCqNxI05hHI8gSm
Xrruyx9kqFI0/cbWvtOYHXjYZk8z2zsh4+eVYRwWAU02DOB2ynE2rxrbMVFYqw8Q
uO/YVkssMTJhFWjOgvyiWauzi0lDkVoYxiN5on6BKgLh9zxEongr8gA4dQ6xn9X9
zd+8BPEfvcSAxsSyJ1GjCcaqqGke/H7J96Az3mY3wgUYMSUQ2g5LrftLsZbyqHVP
MwXHSrzzmpwnEzko9Bf5V3JSQghRiBE0u3bT2AoO1kjqs9q+cxwAxzWyJjJ/8Cyw
I5cGC95BlPCy+gDHs7P1SzLuEdcv/i44gttDO3nlvgsrtyAVXEj79hrrWYGrbaao
Qmc9g0UczY/MfpAvgiS2pr1gjg5+4Bl7iL0k0N3sNbB511TKgBuzLOWoNSp2Zzw+
Eng0f4PnETBetcGVQzJhLvN9I9ZunSPOU2NPQ5MICglRunjYrkhjuaTve599XfFX
NVxONURsuXGYDyVV2BVn0jMrFlaal5UeBJKqTdDxuVU+myVyMcRUR6eYSO9qJmhN
xBzM1BRnvSYlp9tcVIDPr2yj6Z6vm80biis93d6abSoCSpqVws330pDP44iJj/K5
/tPrd+479kNROIumyhN2pFmF1EBVi34Oe2httwLZbpFKnOOZimlw85kfnqxF6w25
81yGY8XSG2Xns0uX9XUW9acg2ljFCvUm2bAD5mSlD3EXzSEknyE5qGofsqEUVfGK
sA5fyMpWtUsGxScVIIM1zz2whgQ8AMubcX1oJvtoQOsl529rgPEAafc5kRTREoL8
Y0MsW8oBABtPgcVj1N3i58KuD2mjJd3A/D7Td+D2f5aP4DCFWhuGKnkOTwGh5/nk
spKZYyNOasGwgSgm0Rm8QBDq1E9tQUznj0zbtJ/CJHbtARW0Nwo8V2fEjRNE/FmC
bXac230qQwO6vj02dHyGOHgoIoUWd5shkd95StuZ7A7BXeycQexgtMjS/wP8IfB1
916jzu7kPIiwJ/YX5dM3TtiW88U6lnG6oCWO76hUNEjTEtZV+l+SNS6WtIpNfGdd
l/04tmpUkRvbB3MtrXUkI5WHS/cUC4Qp3G5O3EgzD/6MdYuE+bOW2vf0HtGPVUSL
Mc7fSYf0NR00JvcHRlWckZPlpgQxnPCgqYQF2SJzAMZA4vqRbz0538b1bzP4rZmm
QGVLrwOflCZ6fmgeA8bSFbzMQBKTsnWwVS9PPLvRqk1woU6DWLObJiaYFG/HEW1q
0JEc5RI9FRXD5kZjVP1HKqemHzM5RJxfc4/FU67HwQgSbI2kOFDUptKQOTFvM+qk
NNGtxY4j8/6DIIwZUyvjyka6deDrLCaXkM+inGH1LKWE2i3Xd5WLYIhW3bc5O1Sg
paaD6zl+5uIpbnYptoacf3lC3DabWU/1iX3XJgeX9KwVRrjYLcQQHgwGRE3CzaC0
efQhq/ZXUHe8q3Ck80wclky70Z8P9RwZhebP10zAczT2CqAimKVxFyzGqStd6Qob
ROWBd8jYhJzfrEJxgccbZMz2hxUke7h6NFXVUrpfDwRW/DBWxN/f+dEEApTpFhMX
/LdVtwhQMmxc8Nka0mCw5Ef6GdwOPSPemn5y+DDDFWPTQI6cE76M8SqzNkGrwnsM
a4sfUMKq1obMdk7VKhoKy0MGa4q+sDQe+G0UDGG6GLYptMsW7P8sGRQTWOp2ObsC
MsP82k4MKjWLjfp0ApwW2QaqpLFyJrqCEIeVl8z2JnX6vSu/DvpWyIElqps+E16Y
0vOsQhiWTsQk6uFx0YG9UDNr7wb1Y3FEXvedfitYDvEy1BMYcr/eY+X8QKNiQvLc
fBPjbhx8SLdCQ7vxwzV5lwfdMMaSc+34nKtYR89hbcrjAmVDC8mZReiAXPTSLCYB
/RJ5Pelbl18jOkydGRQH8IgUZMT3z3EDNWnR2Cs+Ow0vgRazE7Edx9TjJ2mB1di/
U1JQEMnFMYhbgHg/DBSemOJgfi6kw9NWN3Ng3I5HcHGHkxP+LAJhVe096YGpyHSV
GbJ/mAgR9eW+PT0LbzkDMVwCCm3IrdmMKH9T2+mgRhuySoi+YQXpU8GRqwVCukjI
NdAKE9kyj32dNcdRhuh4f5pYmncOLgcnAvdQ3Gcq7E2TV4jBTeMZp2cOluVKgt7r
cizHD0qLIm9soE3AAqmTqkERaSDNoQdyIv7w+wOnmfVPCsenA8Ea9AxJ8/1+6cMl
QQw+dadQgy8sqohz0+KFUOQVbLIwLUtwP7T+n5cW2+oi08SqS7HXbbFf+kLP1iRM
SAsRaBp98COz4A18FRBckOK2hZO1oMTIz0Bv6NK2IzoEkEl2Tu9kefGsBLjv6Utk
O6bArU1RuHiKra96Vp47CXdTLcMHmWmRP2jg1vBt/ExABFPfzjW+uh4GiMZISPSa
L/u3G8bDCorpiec45vnxiJAQ12uhBIBA5PWOC7BuxiCU35b4wdaRHAVTUHcwJAXs
2u0HmtC+O6rbXs5eJqmFUm6XF/a917jBTeEhclIukzheLozuZAHUl77t4RH6uhvT
Xm6jewQh2/Ywy/tZxeIpxMs5AhL4dg9kYN9cE6seCamLMcYGRO5zpRXCc91/PT7U
qAQK2R+oTg6RD4fOoQr5iMunXo/55gbBUPooNziQPEJh/D/p7wbhgHYm1wEVbEJD
OsxvT4c4Myz7vVdx85vn4KeGpnkYoQVl3Nsl/tEZGtIMVEVGJW4CwcjYp+RQ5X/j
ALQTs6HFElesJas80iaiyHNbFMsJSKB8bOe2yHetUWrEli9p5Y5+s6oxFXADkjk1
zlKsVnt71TGHho4XT76LDmT6MzUpfu4RPwbY0Uf4zP4aFzcp20k5hTji0JKC8dVe
7z8AVq8oPeM4w3eX/Shbh51mBlUC4WG2MuqHC83XdSqoxjuwR7yfL7IiVG4o5Mzx
KzDCjbijrxvUL/PLo7JjfWS39mpOnnULyS7Sp1A0TcYU3kMdkPJ44+7Ig7QbBf+n
nAzbDU/X0n3m0Aqc96NOY0GZA5tvVo2OVxZLJFO4vNsIPRq81M0UjDlpbH045flf
z7mCOdyggzA8COYSydIRj4boFd9LpJ8jAP+m5hph4I3L11o73NSfFvNEXLoLSbJN
EcfnaaQqJQGM4pOJcFcmhk6APq0PtXQYxlwWe9WQScdvD3r5ZVkf07sf8h3S/1NC
g3CO67oHOno6EQT5TrgSPLmMSc0x2/MMK79bZ6lXBUbzJUjLXAx87dvosmDPMz/b
hwxdq2XWQ+yE3xFlvxVno6XOEpzaprzBadbtXHA/sL2gEkZ1ptok45VbDaFKcTTR
L7kJ7TD2DTsEXRMVS3DCLnqTlDqyRHbjk0XF2O+gzaXkQ3HPNmA1y1WOpeVxLPpJ
FnUke8wjrVfGwpMoZDGGDbLRwdAzgJVU7p21sgYqbwczTwzngkqLQQrVt1D2uAk2
gAxL1Y5jBn57qmHvtaevG2HgT5qKx5GvrTr+CkMfCsNPl4Ek0KbQYvRdqX2RmEsK
AaSGKxSLCGThWkRO58UlSdWcNApdWJA7m0+EprtCImJCohoQtp4xvG84tyMSm5bn
rXFxE/6zS87wQhFl5y3RGVJ/RVZkKUZt4oDA35EFR/Zr0fC4NQcpUMEtQ4VySoPN
3VPmNIFFsm06o9haNnNiDNhdRd1tbfHZy9lRHw7surjSsLBFcO7CKecF2HTXzCnN
8wSs/rRdhS298jBbRI3ZB3hWr8ICWbkmkBOTtFZxkoAhJgwETLiGEuUbOoBX+aWn
A24rcpbMqHqmsCjW0ZKt67R5yxRV6uOx3A80XxZEt04TwlnXcaMXbNfGWjTLesM4
2/fJB3y0IlDtz8kRsaIifKloAbbojnLnELzNlGz5M6qOutD+iPqUDZB/TlcpXRho
Yfzo9k8xsv9jOZgl/ncxK4/wilCjLWAgHwa4RFZdhAKGmuW6uBfXjkVa2Ybnggie
3A0uoxOT2dfnUjsMtuXgXXRUeCUMaWYbsbkUfiu6564St6tZvUIkn0alAyymMk/X
rPty53s3ywzHbXEeBC2qr4gAFqRFlbqCELZk/15xFXb1uW7dNhppoB5262nFKxB4
tIts0SSqI/oGqJEy1bIfBJq0PPShvwKqtUg1alhP2YkhoGt3G3qX96JV8qOvXeOu
5eMVDFC37Ty/VHsitmg79AA6yMINpJ8b7ap46n+vzes8dBgxp6y3Jgx66L8fr1Ps
8spT765wsmRCxBfgrxCQZii6YPxby9tyjJY1i4sr6SP3tcqAFbhZb203YLXtrM62
SuuBGjRnJ+4vY8wFrO1l7oGduysLmtj/bMyEuShTcRbQ0zO33UlSkNyFGD1UCRnX
5SI4tAPiZnygST8y1fYiYvuDu9YDBbHZuOq6EWNxeUA7SyNbRTDrTu82s7rsmPAN
ELtbeEs/uP32Dpivnx6InEtGxuJvPfDLhFKxQdJFeGXDrLgpZ66ASbQoLFhyCIOL
JPQE7ku1gcThflcwyD9sKJ3VD1FsAeDwintXJoyw9tBu4wPhSxolfHQMTLbMle4a
fjrKk4DyDpZ7h3z6B9Yubb/YTRQn5MQkCTUhzBC1/q47b15LI8eGhXWGOVPX88EZ
wF82WRXH/VuWCEEoe0k/mO6g1AnlnMbMuVn9toxQr5LVtYk0RSYqKLlcoTZ6l0j6
6mdcGJGcQ3Vvxy6xspFtlxLQuBP9nZtHOzbR0Duokxp1/I6Ty61cQTGGhebzcVuO
xQHyXDuMKPJhATtksa2A9uwIgooD3vkLc4C0zNOKk8f47SjEz2dzrEMv+SfCKaP+
LkyUb+jb2WQWOG0kfttmWt7W60TZqBuH65hwtSj8zBHFaN/SkN9vkK5fZV6r5nvp
9MSaHdI2ByVrJ3e+3jpn34qWonRUwtrsT01L/TfS5AnsE0faimUNrc7gKLCsrLkh
KXAPw0DOofGp8HZ+UeAjTeWpd8s7ti+mAyPp6B99v/OtMbCH6lMIwjmGf4M2IJP3
jcUt32lgxI2oJ3sYd5tGHvjJ/Y6XUWi3Ojbq4X2kHRuOzDZD/YHgxA1GSo8kXz8a
XLg+TIJSNn/0NWwiv79/8VlyFAlnP6HKuJbZffNn+huJnKTSocgB4fJhhqELA1Eu
znyw14c9o+uPOxzaSVOXCkgLg/f3EaF3oSjb/J1DQijXcAvppGOVcEzyYBdid6TR
nz6dZ4sH58+hHfbA9zFQMxeFkA7X8OeY+xagkbYbwGMZNxLtZiiIaSHAgUovAuhs
9O60FW+gFLl86+YrSeUZyAJPKl3YKrlzQIxwIKjF7Y2keYjmDdrswTAoqBtTqeLL
uvDqC/jO2YxS6w2Z92zbDGTptYKvAWpyZuAas5mn9AmV1WibzzMIlfJZsH6ZXnlf
oL3mzR1Sh9+6EalAIiSEuQFRS/MySNGUfxexooAH5ZWpT5HtjNfcxX8r7lOIRxrw
H//QuhcAsoXDICUNaD7jXsP2IKNy7QMOuLuWM1Q/SsPpnweENlSPRU+FX3I8uVyb
/2Akgtgexln4Bya8hJAZDfHgecgEVE6152b9yn0AeZnjR5SvBX+KOCrrBbvWuZ+P
LDhA8QrG8bXKhABnMKmQAwE6P4fjn0NhEx4Vd6PpsVGk8kw7c3rZXC2W/et8MZ9C
RjgpuhpYVypigrXpLCP52Bp2kEbkq43JczbOMTybeG3unyTwt23hTY3txMn5htW7
mkDkvhc85SVHFtU0r2fyflT4O2hxWUU2Jad/NUtC2ryyWYDF57vQSXXzkR3H6wY0
AKJRG7XLYizRYqo0HQd33DtKe4HPnifPLO2kX5QXXLP6NGLkVf4Qjbd3YOTpxi7n
HGUXK1WkB+9YSiuq4u8fT96Xo0A2YpoQUQiXI20zdLIgeRhUnz01gI5jaEfSX4SQ
D3DOGgWke+yWfKBeixpGsIoYGlpWi7v+/yK9NKFyscRkzcOMqYPCX1G+0XdJUm/1
0SWKIH3eweiIrqUk3P1GfRDbQij/ablxmK52ewBb4KmqC416w5ar4ijQarHaPSFc
FfRyT2KtLVaP0S8uZ7/hDu/RBolL5fOueYHtElMrBZ8Np7BPRy4ht3kIxOU+QK65
7AqrLeHov9CPeaqvqvO7+8FnKCvIwRRT4mHPyLimQLvCE4GDK/ZiSLvMXs06RgBg
ohGWLWrD3xgFwHNPG0VcET/biERq8kbJ1ieZxtYN71Lr1RPFZDIFuPhfrshlvKKB
g6AaOckxIuQT8z4GHe+ifJ5UR35VNrlvB7nJWhE2wL7FDM4msQysiFyMFIYkSrSo
QaqYPdEEQEYWRF4nT7SW5lhDpEcLs9XTiE/defIrtsDuw6s+mItnKAx49K4n+jFf
Jfi9V0SmzsxrttFDai6eAeRRn2/V9KUZVGoGSE3Lexxj/G+iOOYWevrfVsDyB1PG
o+6JxTn9xgkXINiFitLFQ0v/pDR/NLoJx90aGCnhA5+m6qd09Kk9kbwQSosU4atw
/J7Cz4ek7wdO71MO+XjNzxrJb3u1OQWTTMWXPR/3sWk7FvyriSPMkR1huI0hiear
y4hD/P4MkDmD/CPKjIzheJjtE/Jjp3I+0sK8aR2+Ee8Ekb/pQq2HJmrbn71e6J4l
pe2zorDEEW6Uq26UseKXb8H5UjZjo5g3SIpEaNpcx6ah32P/WzXbbWC6MeVACFvO
LuZMDhRpyLVYEDd7917sCtcU9E2/FuJMhwN/WASLBXljLySdUweMbLlolRf3jXqS
u2Z9EkpXbOo4e+MLjJ2hN+zb2kOHriHLbt7Elbp5Qkqdpe86d6GMCspYEErVx//M
Vh4c6ukLQPrt1BmnQUSrwx84Yxyl3jG0Y0ekf1L0NC9w8azqXbjk5m7VW6/msBQL
RpBQn9ySiusjB5/pmURwpPQd6HNVlwsYKOVfy3SMFmX7EzRQ3pAKpcNTMif5is8Q
Ftf+V6b0RzbCw8uoX1TkPzsO8dND3IEp7T8IS211pdGpN0HSjpPcdD18onW9+0t9
DjgvutCiiro9lPLos/o8pQhwUomehK1guXPH9VVwsu98raTdUKbFoHHQMq8UEHqi
eCluhQR3UzxzPWSC2TMQxQw+9KUGchJPI/8BCjHG/1bgzG/pqP2+BUUPscCxBsBA
VkiyErkeeT8Bn5BzL1+0vZ219Tpj6rKUf1x1Ub0Sk9LuCGho4JCp1DK1OY1yVFtv
xg5MJgSBfFR7D/OfDegV3QhLfqE+WpkQyE4xLWaVgREiGuyhmS5dYqpqQY9u5rBg
t1g7bsglMD4N0aSdIg1ilP3nxyPVdcKnuHiRVz1rGRdjVj+uAK2WpQ7Y0Rf6Hese
f/TaEEwUCGluMxfg19GiIS1IOr9FVJlnkbWtAs4zC/asoG9K5nZ3rkmv5NTJAeD5
nMbuoG8Jhmh9YU61T6kAoEijMYOFaI3TVhE/ehRxbTzd7B0QMYtk7Gc+2T3ncsak
tBv7Dw/81HiOgT5m4thpnolIGbBsq/V4jEJAyei/SBM4V1Jo6MUWZvp8ns8yc0C2
THMsVC2+IL+LPcdT01B1O1p6vliVpEcEVrcH6JyMh3+Fpqgo+9sLEhDROh0iGxf5
w514Xk8am3lDt6jxdeT5F6xTHbRi+ANVjBLxKmQCNrvncvfpV1vo5rPqxubZXFRf
W+UYrUjgmt+myDIJIujgdOV4DLHiFRPAhmZXcm4pt0qoRqfzMqvjK9OoMBnT7y+4
v+GNOCj//6dSmVttw1+0n6ok5Rkt1zheFNRpSO72QlSsrh1h4/APZoFBBBZY+twz
3JFChjAFHGaB+fXuwmJ0SqCRrRYtXdyKkG09tdZSy3wl+OL+X6W5YQvLJWDJhH0R
AIN1qx7gvLmU5Q9N5qQ6Pa3lVuH4697Sf129Mm7p7dCPA3iV/PKtYHEclN2GyRXG
pDgBsy13fAINiV72CBWM522ILEAJN0dj6N4ZvxVSvWaS6g7RHCCXmfDEKwx71pP1
vvry638w7fRCVC8cv4m8Jzs/hePLtLiw+pMF3z2VmiTrkv2G49nlsE+mpWwppD5C
xd4pYUkPIdTyg/VwAPwJ8Zta6jnwTkSBt1lxH18mB+Hx26xw+Czu9XpR0YgRAcce
EppSq2NkybVh+e3p2U+wp/4SsND7WVEyLj4FqzSHx64RKspZiaQE7syJbsOIhcZc
ZaCNwLZxD6K8VT29r98F4sSPsKyiPIS74+vJ6nG8BNTPK5AGWYN/tCX3tty1yrsc
WnT8jDtTHhmMHszZSpqcEePkPzyblxZUbmRbZSOXsBajGFN0jhCo2y7unQJeviAW
v41PUtmpbiOQ49HTVrwa3SJ2kpPLa7SIbVOTDWt7wkoy3jE5CpycLCX/ghtrIJfg
fYZcTYZdWUdcJ4JTOign3g+fdzXNpYpINmOu5qjCvlNYoJ9+YdGhhZmdxlYlsqQB
OIs7Ela9eythiw5R3E+DneDsA1y5pP5ei9YdKtH6rfR9iupCLerYBNGlLwJ0p+e2
GEGcfVxukDCSeoOy9zeGqwqLMMhYGZhbOqh5jho61rFvq4not22JGGLYolTQsuXo
rQu/aGm3JeWXhmr9vYXDEBX9UBb644OwGDU9ZH1J/eVoAMUYsHW+Sh/LhnEiuNnK
NhVOSU/syKN0LnguGmu01W45swtSkUN1+6KTZhO3xj5Ir3iCxnCKiFRuwv92bXEn
kQs9uq07N2ZBGFP51ZtbzB/Tt1Iie+WAVFKOOahTKGTnAqrWMVdhQPiPA8xgkw06
Q29cu4RnqjSeRc2rHIZtnmImhv39yBjWambzZI56L03s81koG29hDzCF7lqXTZmm
YJMybDthLjisqRjzKGIjzXrEFRXPXtL/ghnuqZLQwPbCdWGFdYAE5S1/S0Wylf+r
62a2aFK1jJ9tClicbJdYOlh3lEw89lyABs+mIP3guTdj6akTys1h1X9pQebl2dDV
MQ8L7Nt/9lYctVDS9SPH+YAx8lx2ZF4OpV/pX9/36xI51cxqdY4niHHMH3TNqr4z
32XRkChGAoWulFXINIPT8wAq0kQEkSn/Ukj01G1/YS2pTNZmxGdl8Qe8nskApULw
ismZPm78rp7znV2IJDju5T5OUylhFG9hFSyTWS7aYNaGc7IT0tC5mh9wbPZpt62X
PcFZ1+Hez9NffvI22tTKTYCulsE77oq+8w5uY7scVzivwrnxtparyLl7V+eo/O6N
kY6llSTanv0NtecVia/Et9Xj/FaO3kjL5GQD9YgEEYhZjwPzpsPo84RP02P1Pp0x
Bewf1syOI2ppB/N3heDCDsA6M62uxmwboCtLkE9oT4N02/CoUXyGlRUAD16g+AoH
CawwaflQ5Wg7g4Sg6BJwJ7+BwEZWYsQRlWjIz7Qsc6y44fUxNYAGliTOMzTgnLG5
pjOOCj0tLKzXwrVaslaZCP9oH0bTFlFA2a8RggyFMpyg/IcTF23qp8W5N56sXqAb
Gr5aiUAToV2kggkwy1FOwCzmcBv8zbGgKXv0yd4GLgQaH+YqlZ4eDDUZKNq1gJ1j
l6di+zn8V829dhPIaZTyVh74lkW+mYy6iz8XACNTvdpBwa3Gg046pyQql9aiA9bx
xC5Dd3MFjApP4SUWUSt9TvtH21HwGaWJOY8Va/ZYUZgatHhgdZMBSO/ESjJa/FZk
y4SAn+KwZeezBzVb5S73Qvx0/1Dw3/ZRUqtqf7RDsVEs8l/NpdS7qJQGhawuC7fp
XwDKvyrbm/KdKHSCdHPovbwwIFq6+leAXII+nyQxycwkMdGXNiCEvYEENPT7klUa
l47dB92QCNb3VIFM0imUhUjB0ArPxZdDrJukwugTkQjfdhPCHIbfRtYPjOD4EYwb
P0wgMYuHcT8ftaqVQouY9dYqBRkuQZaBg1hYUp/4fMZVWDXty0YQmsxYduwajFum
8RXaXieL/gSVE3zJ2vtMBVmZ4Gd9zOVTnGT+cG/vR1lk3iJLxpMQg50EK5ZYQzt1
DOKt4zdYnkfFxAlyl4GyKrvF7zADnMNvxvi6vsIZV4SjuOP4kob6NeHvy8J3FMBD
7iXb/ck9slrbSLvLbXgo2wQx7G0Hl/bm7BtP73W1lhhFxkB+vHLOGbKZ+pGcrYEv
Z0+jjOhwzSjyK8P5rjQWrnrcm9+l6NmtW/gmqc5TsOMbLcBNn+Tl8D2frMd4zEUS
oPdNQ2wecRn2C4GJVjTRm8vWEFf0lBCUayRZcpW7LrneEx/6ONLn7zOeFPO9CZv9
xlaS0uikzx6gWcEirkCfNTOLUgLh+lY7xrpnZqpxd78KJa/sk7CpKnEySVCyeqGt
OpsotEpsGjrBiyWkU/I1RSBLMS7gw++jT4oaNraFQgXdwfwtqcuHfeRGimnUJ1Le
GrxuCA2eheCkWM3Hlhqg5DCAwHNiTe9/hKfwzmgJ45qMgqLDkLslHr9YcYsJ5OhJ
0iDZeui/pAa785MH9QYjTzo+2wZTk0kfzDBkl3go6gav99p7UKleD1Fhjulwkw7u
6bGHBRAmMQGSxAXE+J+OA8aTRBTo2rhrjsddNz8EAPiEGqs5XPUCyhvDHyjT/BDF
rMdjpfUWJ2/wuMbIYWr94RJLOPMq3+BI7S7KY0AfG3VZmybW/45EU5+FHTh4hTi/
lbrzNb24SplmcB97aB6iBLU+dfzgORfBYAPNt9yY4agrHb9a4FrGWsSPXLasvGN5
0BO0Q76ceLLtxChDB8RC/EuO8w2LhU2BGG0gG9O4XaIzE7+oRZ91vqeQtxJcpz3z
2XEw/DGJKE2cP280EzyRxZf5FmzGiqjZE3pqdtZ60Qh+GiQfD56k8MNKHDT0+2GD
dzds1Gh20fnzN9rdBpLHV7y7d3IB97wZSqhv70Xbef+LRkghF1LlM7e7s/TzvGck
Q1NZTTogbaeB2I5hb4sBh9mVeKC6S01/kqQWoolv8FQJlksh8beVDXHvHcFCzHpR
nkALn5oRgtNW60RT2AoN2RFGW++kN2+6qZRnzfKk2j98ZiesDSWF1RF1iSw5V6rI
T3BVJFaLPHnLwZWn//kogGYfQ/Rv0aCM2PdMNYVVaAAcjXqzIU4wB46R2wLzDVST
1BsGL3E6NmTY6g2bXsoQP26s+5j5wGGYTcbY69TZibggU4JsPlS7vZnebBYA+roJ
zNkZvl/7zV7qTuqCWdN7oZEvSxkhoulCzbqD4dbLS+gyY4M4t9ia2tsSSrTCjs7c
zrW0MoLTbMU3WinHzuXGMv8j5uMwWU8ummvvD9e7rBbF57bHJ8SXDsGM+ytlo5Bj
mmJ/z8Jo0cCvKri0KpYDUKvoHNstVFt63ebZw+fxe4FSiTIPgLUpIBZjnQTgYx+4
2eNMeBTBtdC2N16VqqgCgAxeHEP1kNtlb1rR9S1dOKUyS9NDv0di71TFjgJDZ3V0
8UAXZ1FWIuvklMjThYF51Xhg36TXZKQ2dgkb8AoOYc33YtwnbLDEwYRC+Noc0/SZ
l4Kl+e1kL1tBykWDTXsxpvA+4xhWqXuvL28k3irTXybyFrXcPV7di07wRA38evWQ
/b99Gt5u0YEfm06hWbMcXgGnyvPcLZ9koIOav4EhyQJRvkE684uLY9yJxVL0zSJD
r54ZAYmDhVFu4TCxeiGhLa7AOSQL3YfljH8rCvOgxqP8HnutTGfVKoQLQGdlxheg
3nUtQpDWzt/I6+6ocuGquuz3NEXHpkDpzAttWrdImDVBNQ3fsVQRL/SX3/R/1KKi
HPJJ+OeZhHJEvlS41qrV4DNeBPBzv26GrX6gveuckq7aezjdGimTv3Wn68QzvDgB
5FJzPqHIEsTZldLB7pXCNLnE20hvgQz3jck67l8sPEqK3u5yz92Hdru/Di5cH+dm
gyXsgq5vYEcQC9SxR1/DtM7dwpFybCRmraGagWf2RG46idFcx1gt1+BfflOz5cQ4
q+2idqAazqagFjtu01JMo2Sj0EwBrHgpzYgqNEr5E3W2vJQ/mo1lb1zGSUl9p9hx
Ys4sgfb6pAZlHGBZAB404d8oucBiMtqprm4unMFm4VB8xnAws2Ise7ZGkUzuTUv1
QnHyW0HGJjtKZORT0DNgOdhzBunnsuFga2wiK+DtP2oN6LHCTovhHgxHVwvkKMSJ
GdXsDBS5b8i41ESrzkOj9jTJtC2aRt7GN9MWmI3Y7KsZ5y1DQS1Hf2Wati9uV/+C
2yLTHQfQlbuULVngoI57xSazeLa6DefYzy6ALFaSLWf2ZiMKY5mlB1ITdqf4B2X/
tb8rN43bc4kRfiMKSXjGgRKclYTSVlnH8/EU2YhI89PlhZlE2dzvEjpgmlHsq5jm
zQzNkC37yHAaQonwVxdimeAR9BTw2dsZpxS5F+8GA93qkx5q+jRW7Ycrky38CgLJ
RlQ0KR5mBdMAlXPB98V0sGTv3xosPiqYFRDt6aeZl5gJmjB6eIYM6REwX3WNTkOM
eugOqy+wERD+qwSGSvjW5qjObVOcd9iN8TPcSLd3bnhszVJFdFbnwFriqasvaGR+
p2/miVvNiowfxkuHkmkeybNRc+LO3bUwiKutiF/+cKzF+D3t3RwXiIpaXMQRJkpG
3SpmcxhvAOCP4E76XKo+WHnZDgT2a1g9rhSoTrKDObbxPv9lpaizhWSZBWm4ukah
JONIMXv9wxeikogqpYkyto3zZF6bwWU/w4dZiVqixUmDxBo875GM1Lr3VZJkmdZt
QxrIT7eJr6yjINfneomfHNRWiVis5GquqIT78p61j/Oczq+AvZqdYBEjUuTlfk1s
uALHY+bHzCAwiDXCJa+lhJ28+l6W8XHs9aEb2f8HG/V20V4eXtA8sp3cQz6g/ydx
ZDd6hS5FJh0iW8CFrb2GPWCfzBTvvMyQ4ESIrcuyOHJIAkhvO9bNubdj9SlVmb6E
xVYDlYj4BVt0DIY2BSEVai0oX2Tv0DRYoPaf1DMvsaS8OdoT31DlKcPsKWP9WGoO
Ifo6nDSV/70NcftJCPPY35v57fGj6ynD3Ni/YDQr9nYitIdAN5WU4d5kfwKiW9tI
S1SYBGXhKG7dXEoQKXLOBeEZhize5CjGf/5YFjQWarNhDHMFo81jr40N+bNZdTrH
QE5obDjQp3fACcMAWptfj+uO3OJlqxDX2XZ6WiJrp2d7KzcAAbqKjhVXOse7Nnkd
Kif+6QkU/1skIOaAttqVNsmDId5UBuwgs+RYYk2P65K2ZeweBYOAqAASmKbPA8qF
TWKFjUE8yLcctgd7toNeGTHzkjbQRAuqTc2UdeZnmYPiQIL7qZKYwLCvIlVRmWYQ
cE+IdebTy56IrQMmVOpKGe3yhr8gDnBa/W+ojrQMiC3BxDy5L4Tqqvmqa/e5T4KY
B554zqhNoSDmoM5AlhAPSxjR3ApWlAhgv+2UEqRd+h8Npk76l+jcw8guqXx+2LwH
fEdazEJhM2EHiRMxX0Sg7DZNrXf3U+hT2yfLhytnnuZu4uBvhfBMjQ2Bt7jn1nro
EVI52rNOHobEhZj3p5xdDO4rVYwyNGmPIRFQhDYJmIw0vkOKp0IB5oyQW1O8mDmw
tpUbkBpWOvPxOwkIPJL6T3jg27cyRFzWV4fHf6sUJk3CDjT0oPEAyU5jQhGS9h+V
y55U7avg/Alf2v5X031V88DQ0sNfehY7NZrDued+kmUQBUoI2RjsqTSV/1got65x
BagnC6UKQzeiOFB8V9Msj7cAvBdKk9N7078X8U32XFD9iJv1watWRU8sNsDlMKfA
d3LCu7LlImiZQBt0cJoYP70ToWxS4cLCgvugUUyi3UQRNniXSkGZ8lqRKTyTqSLO
717Wa5Uz1jf8rI2OrVRBl9ISyqwrZkJUcVfXsttbFPkeUhm1THv3wJfUOsuePdRx
i6Gft3AWzCm5hfi1uGkptBhK77ucid5QNt4ymttWTvhsQFjiYKZyz9CiTbwOFlq9
z9TkSxnBWYAYhY2UXHBaPcYUVPCnEeQOAa/ObZ9Zt71Lbeyg1RLJbOMszlQ3Midd
PV5FENEXZrmgtD+7U9zFp6jWzlxfYHRVZplZ0BhvU7+Q85Fg5jNfGfL1kFdxggoH
xxlL3ZxSbi3nZ1GDG+sDbUsBvXyT4bJurhUqC7dnD/eSww/C08SHRe00iSlcItft
jqpJ2wXGYYEQiW1OzifM6g65TFsMDc2k3nWNZ1zFW20knD7KE+nrXWh1BJrcIw2Z
l3stH6n8yDKF1LTLDzPJoYAVInK3TLJBV5gCR2gdOUXt/aFtdXgqL66qvZjD2uz+
Lew4LGIGoY37T9KfCxCNPHjFMY+FoYDVQMCGtxLgmOzAzyDI8WMbwJbuvN+bHiYU
o1NIQ55VOqOMish2q+1P0mjz1B+AqyEPmJblNZrIVZ4hHzT8KEqnYltnVAIQ2ybM
AG0xpjGjm8wdxEe476YIylEnuztpcRfQlvbylcAIGlzLplhPpsBuvsuyJw6RvkrI
Tu4CtkyhznfxiN4tVVhhm5bXhkPsstaPL3ACNKE5Frx/J0/7COjBvl5ng2t4Vcl2
CXMHRe+w3wRTC9vb0OGrP0OShVitoFso+vTVfmqVFhtM0Rqa98S/hcu8ylCOeYBS
Vz+bMNTpR6AORH+vnQkDJ5iTymSGGPvE5xwzyOXoXuWVkW9NVADxWxHVAV7mXdCI
TuktpLc/a72rsBIuhSYZ/5Q/042KasK3NzQEbKsotL8hW3l2LXmJO5HW3F5jjOI4
k+CVgT8OGRs/nylw0Y3UZTiClavn6vN2wgVEFCZQ+8jtWSaPTqndcwWs9GKbiNP0
q2OIC+0YDtD07DFXmewax8XfpC5xW817OSmVlwtvbHEBDvDCU2kAAc/dE5gQZJmz
kiR+YCvA7LKTq6FTEMHgDl0l/vfsntS7WO0cPdh4wfuJXxZvlVycvfF5oyPin7+a
tCJwPGuZsxXzJ9t56d2fIuG4DVqT97eqOOu/eGDVXPSGu/YtrNXsB43IswExtdEE
fMeAm8CbHucpnG2AfaXUYwVStI9f+TmRbZZ5HJtd1yOuMjggseRT3JduXJUblQ+t
tDpcdPYtrL4C/Zm/RbQLV7+F9UC+ke4r+4dGogOXxCshUogjyz4x3v+TOEsRkKMI
/XSUO5PsHqUhXhISFpOb5jvnGLA5bm3fJJVfRWDscAy300LBUXoJX86nfcwDOnAf
YtYlmGuITJSys7b7bJwRM4sbc/vygskqRjfWVqVJQWVt4XhHaofnYMkbwrGqSUb4
HRc7qa3scU6L1exMgqwMTuZHrT5xbzufIwZPQ3f6Zpvbgsu51AZHarjYa7Cign34
epkPhv7BUpWV3aWD6Iae3okfKuPslkI4DpbaE+/q9sAYL33kxuQuCFN5dJXUkM3h
LD5XCspolTUkXoyZM55ohhc16mQW/6k08o2g8H3ViRB2DqrdolIrzXqYJwYU/bC6
gQFzTRrpd00JGi7LrpSkFj9QDFQXWpy5aAQsq/Zgu8/8IW8hP6cB9lXKdMDBxm+F
tg2wrTiAqYaoUOdEtCQd2avdyUfCTD2U+geIHDKkLTmGXeKxHSpY6Zp/dQISU+kh
Sm9+K78/niJWX/6VR7L6Xoak2nmUhmwZr/9WFRhGha0UnIB7z5W5xYkDwZDgZcCx
stXOJaU/rdasJe6hKy5OPdJa8vhtgp598FSrH+ToECCw2UeEg41fK0rFgJqg84Rp
ZRdGbGADADPmTuE3kMe2Bm/N+lU94z17mVIGOb+ckOXIPwQAsyO9ASJyloCYSgCP
iV8AWkuVCi+6/PL1ed48heaj4e0M3QKN3DdSWi49fjAm13A9eUgqaxh2dyVtn9yM
S98C+X0wKHZO6zoj2y4EjZPuQCZVq+s4q/ZoSYtUsqbvXG3oFxRYTHLI0U7Sz9zd
3P1au65FPxi5ItiWbOfTSHMtTX9Z+r2k0JeGBazsOmWS8e/Dz94U2GN9iN8pCKPc
W/vyeq0UzbNurBXPJ26NsO3BbG/Fe//mTA5YHyixNXcNNy2G/nd3EK/JsA3K7Oq8
0npCOE9e/oALvq9WqEfB4nZKnxQ6L0nmStsAMzVjPSNxHoX5imMs7Dn1OUx4ao1/
VXTWDmnORplGhyDWKLyG1O7wkzRadDNNSHDiaB0Iy5+nEbvfqWHQYL9kHX0ZKHU9
bKTFK/QP1ow25usc16vulGA176aGlZ/l12rDXayiWCxz2ZB/0HXuYzj9jO/nH0rx
eNB41Cbax9vnAKllKU865tjCdtVLJ5SXMV1vunX2eUqd/hqNehuHP/5o/0r7ZaBL
GrLwyLvnq37QNVRTfxZVMc0aPTLutJ91AcmVSOD/PHp6cdg97E2i27pu9jeOL5nW
ljSnLzzBtduD1UvZ5a+hQoL1LJeTYzfgK2R0akq1hLR2MvE+vmBTC8zjPuizPfk+
VWP1Em6rknaipz4is1YgCkB9rmuzN8IUxZIPw2Ys0izEk1k6iGloAnXKoH24xfI7
p8O7du1qFnTXf1bKKNyz6pWu14EDZ1Midn/1YOdfhS66JAS7LUqS6YeTQbdnc45J
co6ggv/Ilm9R1lCusT+XqE5wxHBuTlNZXN8PeyQo9vdcron5WrqdT+r7ykhsC5/X
kjDPFRnFTQ1lJlAp/1m+ge3NPGOtQLRUTomUBzfSUEWOuU81KfICD7f1dW01pBVd
BYBwRJ8SlSpXojXh7RaaOB3X5vWL23MrXAwpYN3HoE523mi6OYHJemeUAsUj4V1M
rIjNgOdJbHGPCt8HKzXMvFSNLBK/Xa2Cy2Pj/JFnwEYvVlkx+7iYhxN+ouiUJKlS
Oj2jbHFqdH1piyUbm/qeFfvIyE8m2qCMp8hncztoN8B9I1r/GkYI3JJJYEHuDy74
hyK2AEmDeBPUfCp6+AyzhloY4HvivJWysCYamUFfIAT5XX5WjGwT01QtIMwvcIis
Z+7pJSbvhA4gt2DBOVEearyMHsuLgSWoXnBOQva7beNG3VMKMMa0UDdeLSs52DuA
2x6EVEQVvxBRMzQoszhFeoIfpaHEyXgYBtG/Xba82Oxqstghb25XZQCjwZTU0jfD
K5Y53R3OcjoM31Uk35OWlxJ8jXmWKgNB3uKe2P32vqHky64jLl2hOnYcBkX20HWp
C9NFZl4IBRmex+02FU61cazWmw0O+fZHvwaeOxdV7hsNveGIjRP/aVpyO3dmUYZ9
uJpgDRUPVuBAJkAfqdcOe1PNcfIRKHb+bvClp+kINBOSCzeoSXCTyP8XX4r2M3OX
RVjR4OJublv9ONyFYimqUo5BEh8pw17CwCe1LoIgNHlmmc4yKzmgavMzjwGirv+6
EMtAir35T018uul6bCxHVMM+h+WwAPj22cb1HcjzglKL+wMi1DgChcBrWEqFvCrK
49GRtwtyYYxpNGh+Z1uAqSA49pY1WSXyHmyMaWnBlcMWNF+pKtkdlXoDDZMbgLNE
YWP49nCw5pXnAXI4RLZOqb0q/UZwbUlf0o4Kx7+9wMPJsqP30UrEMmGocv5qYmId
YFYwLlgGV3pJIwGtu1QbtlyCZpLV4DFabEaIKE33ByoPatqTJKcfbezPOwEDRuH/
EfsFLrswIdKDXGhMzc/YZAJLZHnyeuhJq1QQ5by7JnWvIaJvb+8HIh0vpLIod66j
UUOitVEvHuBCIPZ6GdAkHSfpDgl4jYO2mEiEQdcQQmvwLmUaZqvsjo4M77Q9IsqE
KVKOYJE1ftqQZlOKVan7cBrkL5s04K1HouyRdGJznVqPzj10Yr+J3Obv5cqzwE1c
acpbp8fSgN+pGpsfRN2b26QqDF6IRgaZ7QChemBdJ2Bw6j69Qz60EjgU/mFnpvvG
VRgeXYD3R8NSfz1QIirH8d/y7VCDM+ZcB4BNcjgO5mXcSm/y2YrE3rrZL6A+OUfC
f/Flsi4WfEEh9nHf4ssHryK3zThcStLaohLBKya+EnQxRHk26jRXfUscMIT0Z2mq
juWM9b48n8k/m9oTsfVlF/jPb+Xa7a569toHpJyEmLmXactBWLbMBPUFMHMIcXBM
gNpXMRYyM2Kxdjp/sVC6aOau9MXWKB4pIGRZaVnRiAxuI7WyLlFmvnX+bMiJ8Wt9
LK6y/HPi6Pzk57y5gQKMJev7SHRx04ChT22fabwlbUeAW2iB9+gT50BomIZc+V5K
W+Z6D+yltT/0yc9bCJ5/MdqyrHbNkRPJ8MFSk4GNwYvOU7L2gMK3urouSuSVOySX
ZQ0J5u4zllLQ2AnyqrIXRmoKXQ9hZjYKHlsqihaXWuyAk28F9OJJaIzNvdRVTQ1c
ybPddNfik8LOZATwtcjZZPwdRlnG6T7L0cbFQm0ptIAI3pRcGTlHMV5TQHZFLloC
M2CHvkgFmnc/OpIhg5KNEUmTWzOMVL8dUKtL6n6LcrvSBPFPVndXf4xmoNYWXwQL
9yHCe51EnRmcyEiAIz88iI02NleA3Yz6EDdYIGfWHd3RCoVw3dFa8bT9+fn5jm87
2BZEjlGTacqSZ+0M/GPjOTQ2q8oRHk8hRSpj2Gy4633YyAkbAtKV63/U8fJfdFPh
4VoInOZ+JtwrErKUu0MCqBWUWY6oEQ3PiELw8ippOt7I5Qq2wVlwjmRmYIowPLAH
18HTr38mjstNzHF8wnGeSqPl/c/NXDx4afDkk0WqcPHWYGVeZ8hKgqNYtSozi7oi
M+rUdtNHHM3FFVcjSx56pR9I66I3iCSX/E2e+2BOk4NGDAsUc9FE8M/fPe8HWz/S
8IMl2NjWkvSQmyXRueBoQdVzmXvdCafxw4lobMA9WXi+6wCRr42AbZ+lj4r9U0YP
vidPdnzwI+odqehY8VcSX3vT1H82Ulq7hCjVGZEw6WJ6Mvhb+FmISPKhLtUwh3Gf
jArCIiKMD5cFWQALyDLrUZFCjNqugnBkC8T4YhMPzpO5ms6p/Mke8XL1xKi+09ZM
DwIP9L4VVhH1y0hj54mmJmixbi/t7mPFKsZRgJ4INdK+xE9zWXVjg/W3+B1/gFKw
TUTbWMHKr0UpNiP2doQSq/h19yV1az84TD5EA1xRgWDrf/6s7FWJfPHj6SmW1Cg7
jD1oiL+CzcBGKcDzTzRpRrVEn0bCs3ODTg6ifZ7aqRdtRS5CPoEMpCcv69Hrx34b
jfLN2CxdlkwtpYhxwU7LKQWhEcrH5t2zFD0Xw2ARt0pZE85swL/LcsDq+TOgbwZ5
AB3YWajnG0mWdfN9pZJ2UnjJ3ckCDpLXPqbyw9sGJ0f8JR1InnpXG6xWtKMb7L02
pjHQ8NP0A59e40N3opGQabFrr9+oBMg1cPfVDIlqb5a+2PRSMpF9FBeeZeBQWPlI
5FpM7Q2ZYsLeBhUc1VKgrhJdb7f6PUCPSoU2U+bpus3Qy6XnSlCgbRc6sZpmX8Ny
agf/Zg9fKK+h+LBi279kFVvc7Znnijc2GoO2TE82Al1mY2nMgrOv+ksxVtFevc4F
1DO5uGVGILLr/Zja8sJtTcTcGOjSeoqfB8DPFy0zeOWoXpWxFCX7wmoajAu/x0Ti
cb1BOGseeI95yyx6nNg/OsSuaI6FZDZWkI5PtgDM0nAgIpGk3v9pwNf4pgJUmzoY
K02kMWsdMhE3arvM+gUgKNZaSCX4NcwA734JYPJQMpiCWBm2EZNVzBB5Jus7PjAQ
E2mnOEuOkNEPJvuDgyFq6m2CPalrCZifEzScAIwQrgIPyiDWDL0nlZnk9A9RUYhv
k57ZF2ld5qV8o+HhRDbHcCA9tkps99MpmKSEuL7/Uw3feIZVYTvLTQuH6MQrhNop
+EJESVhk7XyVcHkuKWbxyqzvw8ApoU0N4HS5FABLemMh5hUDp3aB1xHodrF/Bl7X
jNnXu9B+Z+GHl/T/JxhHkRnrI4PmweivPHRxAKZzXlKSmjgET/bYPzl1jZF5I3uW
rOjJ9NbvfRI+VJhexnw7+3KCD/9g5JR5f1b8pSOlC6+WaQOcRe4AkpGtjLwsU+Ai
VWeS/xZTcuKV5WlT/KacRXRClNcQm9BwdvVpH21TBqq/Cx4h+fJ9WcA+RgMQI7kN
zD7DonaAetsJ9FFiDLEiNsk79R9Mmb7vEmacmDHt+vVUxGBHeXe2vOU5To/s5KrC
Eg1jdJjZGU8iIjvy9sYiDkJAIMraMOTGXcbHyV9NODU4NgqrzGRYqfJ1AyOBK1X4
zoV26HLjxNCsj2em9Zy8G4/rDRaT6niAOgHZ57CJEc16mmUBG39JvtKGDXWghE+O
qTSUBORpZ7tUzvH4a+P2tq0PzQr2/EoBqbhOUczU0Y86afL7PCEbOxqQU0TiwmKx
ii9QXft2EojYSe20BnhEUtE+ZNc34Pe9uaooL8OxZzN3TL4p/jwfbVmlDMVSbiZA
jcDZFIhgQUgX4ixLRz50ECOYMKzd/tfgNF67eIkH2gBVc46JHE2IKNOpqg97PT2N
sghwS4JKJ3GpRhl3ChH121Envv6Dmp7AUucqz6dmp3NlxLWuIWolPugXC4eQTqE8
ow9nLphO2WTBLner+uAiAA3XJn0dSZGpYVUu4Yk8kOkXvEjlf62zbexxKHxQxTx2
Wj+wTNhoEz6rH4Tpz8cKeUh/9Y+xH0wpRkLi/ZzqSmI4QF89aUiRgSTsLNYX6qIz
pNei9F9mTtqFWHf3vadR5KDOXw5M5Rk9zJypqiw0v4bAw1TqAdRha6YH0OquxyE9
ul8g6aoYk84XuNYBpf0yMqQEkY1F/x78WcGq697QsEOkql558gBlHfAWW2Kf1joU
ewxzJm9lXUpl07OIQRC0SKo9PERFw5cQ/O7fVG2ABWN9Kcad76fKkpm31j1bxr8M
jNUWQZSTs12oVUJ5l+/jxkCqntuDaZ4AcP1+ppgw4ZasD9Rk1NnMA8Omwi51ao47
CuVHVuznwqyHZmtquCYclCpODDB8r5VijzOsTUCVDEX4fKgINBMh23qniOldQS30
VBTIYZ38lswMBtxEbfJ49gAFIvFaciPnn8uVkJolc6PwF7Zhkj5+ye7+hi4lWKFn
+oLk0bOrGwy0ntsFtpTAJ91lX7jVhVEzgYbtosRMbzqn/zVPEmxS2KrpWUDdzFM7
rzFITqlGTnfO4obel18Fm2sj4k0ZTCAOJbvNlHifSiLPCBvtiqVsOQgRJSB8MEH3
OwaN9QxEBSwvWBJE/pJ6teCLACcWiCIEzc+HzghEXrRvhK3lNVk0+SLM+uQsX8UJ
Ev4phP5bLBLGR7k9zkasaMV4oqytJBUw/IfLuFeOiNmtKZ2IYMyWI0kqPf9b/vpw
JOxikNqXsTGe4tQDPMgVC1/wovjw1yZ/cI0nk/YxyNmXDSOzgI7wpSitNx7yCWfV
qW6OrzyUrB8bvMLxOX3QUAKgVr/RmBTrpv/76Au7vhAORklnOeG3GmG4QD9PgTx1
PFz7UzbmJfBdbPC2jkbx8wPSK0SGuR67vjHOjDDSNqCrktbY18P3HPYzaF47LxRu
At3U4hHgoMk57/ehme9SL2q/0C6cmNZYjmKiPYbMpn5RBiuJ2g759JYg4T8RR0F2
kFzeAkQj81Yq1DUjfZxNuYUM7CyLdnZyvThpzlBp8fnIpj0/27TPpF+L+SM3NmOd
YU0gRVUwHVgmXKeVFDgBPLAi1+M9Xkp6qPxlqF03JKKL5eCxibmHjDlhOOcUU8+1
J4PqJGCYThq1QXbvIl2MZKbUria9xM3vEpTZ1fWyC2CfmEI1TSpZANnMZik4+dfA
6uZqLUhSjUJMwEXchlI72pCvuF+A9SA3xMhDiEQWhvSfhoOMg2hyQq1K2BlkhGIw
XSLQZuuvpy/xDB2UIBqm3oI/c4i9qms3A1IU7YuHYENsy+XV3IM5b5y+7TrM4ADA
a7OZlKrfLfB8pN4aoZz5MyrxfXBIx6hoceNRRuHb/iLyH3A9Y8NBs7o9fQq1t6uk
oMDoTvVYe7Tcs/I0CxKDM4gMj8mwz1PMOs0G4fzuOnya9qF8HbVqlL6TQYn1jzwy
FyfjqsAuLUiAGIq22yhUq8bXtwuMor+tXjX76CAjJoudZVZB+k6iuqRFZo1uc5/6
pF0xpR+KngXl6xrrBPK9kwKxyLLuf5Ya/bndFPYdOHE1eLbxNOkn7vwSVrD3stm+
p6flDvnmeamCD32wTTFh3ahctIj0JiHpqOw66bduS2cvdgnsBNLGcGgq05nd6xFP
AYvoCR4kHebtz1Pkp1B/LUSE6MHID5s3g9t++bFgQ2+SBgfMYdBXNO65P94EyJKQ
TBtM7cyxE208oxKXcLoyqt6SFYY93CXkBWwehisiFRxTFZf7F84F0zy3LPwyTxM7
m9aStBPvzMy3YotaNKh6Nl4DJSPE+feDrueqWI0jDcs4asp311UzidJ9VyqJ/EeP
PdqAeI0JKpcZBSP3gRrmeWPhqp6G1Urz43hLyerqOg+n3J6myAA7dlFYuqC4byG3
uoWUZHv4mbDjm6KUHF098wXuL9f2gaX+MLmoYDwBLghV3zEIivYqufGtpOEZB/Kl
BMb6wXwr8Bd+F7LI+qNcKUHbyXxtCitLp+5PNAgibrEjr9HLokF5TefenIgQEQ6K
2DYidtiP3g4FAfwR/91JgcQ3WXVpY1kb/mSwbiCpKLSTotSuK/EEXiCBDanwVX9m
tBWHJGD6kRcYXdVg36PX4U5lv1FttUBFGRjToXC4bSah2jDB3RexYDl3OHEbaJsx
ULfTI+6XvWAz5gDMZNLl3jP+B1XDtFub/fK16AvRACcxcB4+vcuFcxx9dtWU81iT
O0mQzrci9wyrQp1HmeOXUVTdov4g/PC7kfbFKTKHMcYlON3f4+tG6LlwKOHzl7Z0
agLpnzBlmtcKOqElw8H4x34ueanZjIrobbd0+i5qXwEVOmXEqiSv1tqYRWtfTBK5
TAxyXfk2tDVd7gZ9wo3auJuIP/O0UoTgNSXuw6CsZOz5i7B2Ce4ecWE9BR9YqBPq
4D8XbgzJ7OijfvTJEx+Hgjh/oP6o+A6a6psD7KzjbyKjnC/m0SvAiMlCqMGJA4l3
uv4Ly48hjq/XGPT9q7873vUDWmEivbf3kJTzy3OE9fDsQn7OF0yVUX3FCdQeBCwY
nPARRNm/lwOgArp+Y2t8P1cwysW0v87E85alPHPVrs1Kub3gzP2lXtQ9OFU8Y9JQ
cYBqcTF1oUR0iBPhg1lNiuzTrKozs/bDdNHkJkCc+YQ/5J+1Eu5Dh2l8k2ig8IO4
4fYMmEDKTU4bEqHb/DyWRTwBkS00RVKlIRmS9MiV2gARq6GJPPMR06sQ+AHCmD5N
4nQgr32SAchJg8KA4wAuUyivvhXXmJCTnCNlEkEK0Hef0o+FCWHYQb/GTRX+k8GV
gVFdP9FYIbUpnPC40HOsuqBMjHpmGywR7XSNxWaG85/NF2zhZAkpRyKBIUkYesBj
8BaFBLMj7FElJ1fdcE4twGr+USO+dZ9toyXC50cRS8C3Bc9dxYOAP//ziO1y2Y5/
wgsr0DnHWqp5Pmc/KeLm470aSnGFp2P4IGdIhzJs185k+PJp1iA+1swzf0O5wjH7
KU/OBcyU87ppccA5f2aItwHAi5Iqg6H5qEjcbJSK8jP2Pn8FEem9A0zRd8jgsPN1
xySUHuT7erGtF8JGLrRM5EcJuzILskrVH/bqOxm+rnhPcepDYcIP51MH6h7Igl6X
BGAZvhi01bpAJ5a1lhn8lMXr7D+wk3D3W/qiEKDcXhKOJ6FGb0eroS5EFsGlbGXE
kMT787A3jJlmsD+rw654bN+v+bpDtulr61VGikbfKKVnHBw0lgXBx5BEhwwf48Lx
TIZqk3BVSADOEzW6CT72lrYl++ow0+IuGDTE/vr7Egq67DmDgVuvvcF9p4mALPu2
omH+JG7VRBDAwFl0dJTxE5mMCkWOdJcQxS49ZwI0hg2EhcGnkrPmNEvmkNdBc7c0
pR1ba3Wo/djbkS1ylNFZnxa24I30L9gNC1StlU92zEvP4pt+jF266A+w1WX2YkT8
beKhgnWRjFzadrRAGzmryaeAdHZBVF/5e2bFsk+hjqv1tmiL4vD8gqy9zrJZhVj7
gGQXZZzGAhNW34H1d3RHw/7b68Ky3E41iyceuG5JCmz3++WNJhGt2Z05Z6u2EydP
+13el2A32cbB3DmRts4FShzlLKQCpMkLdLGlxsX+5TzEFYKmba4IVSuWcnV62fe1
kwxsCl88G9eYO+w+BoXCjIMWnNADJ1Y76GTX6Wg9ZjMQdclHiX8YAIdwq0PoraPQ
tH1yF2IIWEvFKhps5370BA8OS5tx3UpHY+wxDfMWcAyc27eng/zALJdtHkZslpKN
Dy2W+HFvwVe6+2m59mZHfYAgsa44rzDFSMNqvbkNaUfPknn3Hc/MDSlz43fA0C4T
5r6WLqe+tUJ0QWs8XpuA5EYgATOxFEEjovmzwkKqfcNb0lcpZMBwR8dLFoOTV0f9
SfeI6L9kwAEUURAMXIue9Pu62qfVJKd1s9IQndcoj9+B96L35T9/GZVzbV1BTJgV
Xv6PcN5sJHoh2SfpaqYFSPLpinWdQ5yaYH6QRSjNe/W50qnVXyUTjVCLr4uVqXMc
G1DxxWr37gRvNZeOCa9mpPRc6vdYPA238GJEnhyVwE+3GbBM2sNEliDmM7Fxnedi
XOyw86wR6+kXN+wjgmWR2MPSDHBEnmJp2Mv08L+IDSZaYMvzdAZM3PvYT6Fg9tBF
1Xxzure4vXEgE3Lrc9uN3WnQrNAm6RVqkCxT5FA0thJFnUAB2jp1Xr84UsBL8sos
T+K0RrHV5D8DK2jIbXSSQX30LulP8Yb01ghz9T0bPLjHPTnsFeJlPtd7HNJV7ES8
uLZdrV7fUC6tybuTfOo12pmQAu0AjSg76QtYxIrodWmlNx6vZZo75EsRNyGV4QtI
5S+fy5hKw1BGqJG2mHy2zswc4krywPDnQGLeEAiFD5JqdV6qXSHax5EI6SU9jY9u
JHxaw5wcCUZ9ZHgVDMgi7Rqep4/j57xohdTvFTJ7BxkR50/ZQLNQvpJN0hoV/bhK
2QWje/0x8j8QIrnAK6cVMoNda+SdiLwthhQPU+wkru5Kh6Em5TDSOa3QoE3Ws3Lw
eEydzh7FDruIVmbdZyemkTCIw/Fowx9hGfwZn1MAeE+SELGyiu4nWvRML/8fI0xn
ZNIzTpRG5Ovsr5W/YSnKKpWVWJq8yGIQGDdhdk21ksNr3HZIWI47i4qNmTDMKFol
U+KLFgktS+tOaHQh7NAHNtapz0+ESHxCUyTAlWJ11DEeFtIqRVofPZ2cEzCEGg75
OILlAddIjdKyDRJox1sbPMKpxNXWFml+AX+hDctWjUXU5BJyj/prDfmWE0fEk9MQ
q7bLnZ3rVN9wMxrreefa21Nh5JyC1lV0t2rj6N8GU+ZWE/4WU8xSGxMdnXkAAGbA
OnzpgvtWpLGzuS7w1Ml4f3eBwwF4UDfexGR9tpNB9UB/X3s8/7tN8L5AkxKXnQYV
OMt18auyfj/1Zlros8ls7/+yEuKGxfX5R7klrqQ0IsM9A/0ZzRqvLVNQ/0AZOvFW
4497IZljURBIM6CWOAzBk4Sve/345cyqoqoMKXqipc9HgyYhE+84jdC9/gnqQQFG
0qwQj7lZUDg60zp74Oi63JU9m7XKToc0zL4aH6R+vXzbsfUQP/44DDeKz6Jbw/Vi
gg0H29VmL3SwucP05vPhOEEy0VjHq7habFhqdF3zGjKpSCPw5hSrF4Riotx5bfQd
7tJASfF1SYxjnPAc6++7jMniyyNLS7f6+OAtPivqTVxTOrOL0X3NYPhyX3wpDdfM
+kP9/WxfPrtdCKUBWDAm5sS747zPikhDY+fN02TkRw8oIV2JIwON6yyRceKgDyhD
DRu8h84BAHj++ujCmVKmy3zRc87BcBDSHZS1fozL8vd77AM7YBcMJYI29mvBJw+2
X2vBDzwI8T7SLWAovgXcICd3f/Ex5k9p4sWG4cPfOJ21AEUh54lh9NP6v28rkviO
hD+45jdxMfVVd9+9xREcFUof3tgKqof3syU4TUUc4PoNELOLdElY/yFFVbdUQJFD
He4mSy3/Al9rP18fEAEHKu3YNAkFuJlQW+su7WFXB4Ztj9Bduhb9FaBTUVYs7vQl
91PO0lO7qqXrhxgQ/1SjHkJcalAoq4WYzKKJDHy6Qqu7n+tPlQy8BPIsAeI1614D
t2ukd+OM4sxLrT0YtjCjn+63fOInB6vOSlLIhd+RXA32zUubYwEViU8RJvc2fg6v
ZvZawOsj00rpLzQBQqfy4f8y5Yp9pQYJr6y2SiAvbKYFr/81128il2OKIji0qlQi
E8wjpoPqcBBaFyRkbnC7dhxmHtkU1Oommoai2ePZRYWMoCZAt6pmGZm4V+lBZECm
oTW9esqGmkPtbgAK56SjB15KJjW8qAFJm34ZRjiZ2ID07/GdHbdHUqVkNx1lyHxa
gJ5gv+OFrNOetDgS0GJasAXALiuhchQlcnjlotrKo3FW8Tk5I3vXInoQFq2SpX3X
OI7NyNA5IKov8ivYz/4qZyntjKNusgiArZyJNuhZnJ0yCa9NPdFxeqqqCt+t/D1d
romkNAXdF8xPlue6tr8WeDfJZ5QFSArlUX4U4FRo05KHuJEVLDScFOvxOZXXzSZW
n7SC7KQHO0/ahFzQOgmeMk9k+wpOrGt7Q6GcdUJqOcYh0+JQNXB2cnE5ExovPUDr
xZC42mwY7FSy9mCztredzEqH6MvmLyZiXcR+29wgtIvhz8FB2lJWdmGvNKEC9mbn
piJgIBcXC/9dUEHqaVN/SjD71my49A9VuerpRziN8JUyCLaRE9yXI9b+B/gWk1Rm
Qp5O15MV6zEJZuhZt2fSlb3EUDKzxq2L9U1cIcUyTzXIlBJ1xxKF5Ol+2hpk6sQq
xx4zqgRWak4bp9C4ac3MbaFYdLRm82gSAhf3DJOTnRVDI8mVQSOX6UziABlxffVk
nqvrD+Ssy8hPf5PKscXKEjw6Yre0tiiM+cv9FzdzKDK9WMDzp2tdYxMuF8MLEvhf
m+sbYXnpndYWlM/9x7XAui2u1VhsLg9crMCtQeraId9f3rYBu61j6JLEkyMfpkd4
a9Bbgtflqggu6B6f9AaySNUrgAA+K7z2l03QZWch+2rlpxD7nlnFTxeWmP6zii4K
y4y5fmv+q7ozpGgcYe1pR2MXTYNNTP1BTBD9+Yu4aUrqv7tDghsxZYGf8Kehkq13
d4cMgP+x/GJo3aHA3oQtg9no29yNqFL+gNF+0wiiYejx2Jba8hAT9OfaQjilwUPb
yR8IMiSsE2jf24KN67ZTyW/FcpUvp+1vjPg1y6LgcLmEfqPBFVGA65b38aA/0eeE
9RHT6YHD1u68DR8lcvpIVkGi9H3rdIPEqeq4OaVRhkiJtKuGFihoKqbbyGujN9l8
VtjioVsqxMGG4OCPekvB2mbInqljtOY5kCQYhNCBnahyoLZ2s2PCI3EMzJu4dovC
OrIm4BiQI0Z2hz17otlfKjxNfAUVUa7yUsoa86K7ud3ExzbjRkv4iZRBgRfGS5yY
H5p1qh8ceRQhrjwAvLlIC/tUE2hfC/Jk44l8JxgPY0ZrJETr9wNeu6oHWrTXBIEt
l7YZ9iaJwUfiJdomghQ0LDuZWbwqQ9HUvlp5QaTltWNLlOWAt4pWp68w9srGYv1R
hWDH5qeNVcNT0gQzNJuML52AkwUtxG+diCS5vTlDnOaQE14DlJKBIK/Q+WCNWBvU
ZhzAwg2MiMYugUriywAftDwheLiO3yXHsMy3tyAY3V+BKzwmBgPeoUwI4cg1IGd1
IVEB7GfOgU0hMIYBWuDhObrFg9KvMF8HjB8bqL1W5KBGVYMifHHmrhTzodBYINtS
DGMx2IXpjS0EX+753Wq9QXCl/GhGYL7ukg6LkBQLW8PSIKstfX2VkDQbWKvXPb5O
wkgAINJl6k2Vur4mDPUrGAUKBpAfvLH3L4+9mO5lcMYHRuFQvtbAyA+nkXma907l
ozhYpa0eWSediNCHOGKR1Yfgj9gAzM6MoFAyJV5CCBjwhj+wwkS3jMjy50Q2eMQY
f3M7otXfzBBTYmGb3rZ5OfoyZZW5jt503UHZlauZ73qNhXJcWrOFoicI2HbFcg62
x4+zISmVKT2J8B65EVcT4pG6R6xA423IC4nb/wEhf9jzPOGPyrAMZPXBWpPQKfxt
GeULSbHEmkUMPZQAb2VGirBKUSRrgRqcXf8Zyqvunj2Uk/oFiMKE+WFkOwpqOCEP
W1Md9a4O1M0AX+yLCWQa+YdOg2m9nUVVwbyrNcTbRelbGPHXTjIBzf/JB2kAb60Z
WXI/0UWt3zeDJNaJj+c3GMTqzyadQwAFG/Z6F+cNcgmkedDBUOj2PfYvRbwBNfRO
AnPpZLbv5un0+4GzFb2VzhaSiJQIESuzA0Vf34oqyrptmaq3BIYwby0NKuzavcgp
hqEIL3+mR6oTZTXMzRNoI89UqFlurdUYlBgmLmqkJC2YpinDPbx3pVQJbLHZMWxV
ueYkafNuj7dx/fI3lBVpqgZAd0hUDVtErvcNdfiViue72ay+swxrx/ZnAuOZsqpH
POEzfO59B00nn8R6abTq/fxr6VZ1zzerx5u6qlFVQQGztnV0uf9GXKigyETUzNFo
u6XaWcsFT00IrNIdmUbirplntSiPGcINVDmSnOS1GRArJSF2eMkJhYXEGfmBNtt2
IA2DJh2n4WezAYzENIASZQLYw1QnqrfYjh395O5GFv04B3b9Y/zYB4Zwob1vhk/h
CbyISTixvSDXJnYwbNwsObNTQa4/Q+D2YawySeSvKmbOZrfoW6IEQ6I54qfW0f69
36e1CF0LCDgS69iRs+HLIP4QZkH/af082Ajm2GxF29r3Trh8EKbmS5ustqpGQlVR
n84dYxS2i1hLnYi+EypbhgF6tpE869jb9M5JWaWrid1d+jJQTSOq1MLOSvzwFMMD
3Dv1QA4M6GLN65oYChouiSbfbBjnIUkV+9mbfOPVRAzO6wm1YTgLTMdwW4+hVUoO
+5X3XeSyaCy5Ds9mblv62j4Wav5aaQGQE+8G5JWa2nWv6aBZf7SXV8+SfuutSCDU
+X+Uf4T5r2jEsv+trWFNdlO5xD2OPTo9dAPSJ/hFUxa4RnXuOl50I/UtfwtOCq7H
0KrVd2YBXRqYlGIInvl3Nbgehh4J519/Lov+xqu6ixdYhVJJ+8e11avIRs6x74vu
f/o46RWr+o5WI2Xb4D6mN9cT9jZyB5Q4czbsCkedhcVlXVglOwwZj7iloa9Ei6KU
hqABlKoJS3uR/nAnLLXvHIjv+pN4vPzQLu1l4hb5CIsk8mDa6ohlL/5bHDjYZtry
D/mHNW5pGITPUysTEt0iLZZP6QGI/jDtXUUpc2UpsyI0J2EGPXNi3NqMlRUO/0UL
u3aQYBlFwaBp4uc9A9alUcdHU8NaZMNaiz/uOuXO8eQL/iFg1Dn57avPy9KVStjw
t0gnZwh8ISDD/LrrllziglSBmrK7KyZqrPGJwptEkYQcJOq1EC7e7oA67tFdKfT8
C3dwsKV3GPQ/x75mxicxGrhmAdfyEJNXABwzLgrHVwID397QQxvG8cMIF2blITZz
ASeIy4GsOCjX9f9IsLO1aayRPcbRbXbnsRTTSZOVq/InoioML6NUuM0oQGvrOxBb
3bXM4PTNK7/Uj4WCN1sjqiNbTsGT3KtjQGNONwQO6dmb5aGPbm4MRy0cP7UMGjd1
2HUYNlKdzsPa9w1m2FxLGmHRog7eLTHV2sQ54q18hzjzygmco3FOz810xSKc4GXe
lnx2zI8sVlYYl9a24JvE8ci9zF/dgi8XC4NaS5oVcGxqfWTrkxuWUrbkjK0QBEV5
ZrD44vMNFQcpejx+rBK6OQQWsnXoBkjuUioBE2gRhENFpugv2YBH73mco5vEHEHO
UpHrknB961I4I6zZEKF0gsNb8ozEtt5kKBSUJ6jP/5IrMuYDQSTQiiZDq0uJnnjc
sVys6SF1A5dT9rYwbTaLEcP2lfM4tB7Fpx4rBP/B1fPjEV5Y8+ePlrl5djD5ADZV
uFtRaQUAmD28dgL68rmiIvj+HsLfbobBOJdEeCjrQyo9pnoy32Z5N1yGsCpJ0+Ys
NFOxa+gBkvVSQJGqQsmzQgXG1oI9o1CmbDqInA+7TcxkxNvFEhACbbls814PEUjv
ostHfp+d2RWFOngPQ7Ab15Xj2YZ9VTWFruUC0GCQdcdjzhT0kgURVLbtGX7ILiYd
0pPRrG8AP1SWek/SQCBFh87n+/DQho4GlHpTbO2fVw12ACeiovvkvpE539hGla3R
17McPmM0QQKwIOWn6Fz/TgIdF/Sfps1YwO5OkuoigdK49IouG0ipFYrPVqXH1xhQ
R4Z/fS9TXR7aZngbJ5YL7SJhMv3fIyiMScK5lKdRvxqiq19IHETRA2x72Xobvs2K
UDwMW9kM6reCp7ZYmKReekA0ApaS78GI8VEVfEPop8IBglMHoKKg9XCo5ThWh+dO
w0eBN/UHCniPzjTlVDIyfuGKSo07Yoo8jB4RMZXn8+7IhG02lUmkAEJxcHnHylCm
KeCZD6SkheHEKwkK650B4IkyoexK5e4XWXvKgcRHM1MiuufNx9WjGcI9oHfhRxms
wXNkeyM/AnKUOCQg7ihhq7LeWf/bpTeRq7O+4eeRSX5ZdXz7frHcNdW93zanjQNC
wNIMU1Kczl9IUIbIqBgQ0CvOgKUqkZtZoCn4KXEAHhlXQ/PsWtwFDqclRE4zw2et
dJfxYhmnxuNc8+IEgydOFmBBY1/mldl8al1+iHOTJck6lkp8J3/MiWnqF+D5xYBQ
7sIdASmWG3hP4TvQeDflu7NLe5x7KfnqaqjHq/FXXOiaozMc6hH7srW1MbCKlN8C
UYA2ZlRV/AxJjUKBHKyq/asSLRDEtvicwltEg9bra5jKK+3Qui8H3czpmB3hXyLI
zHimTclWH80qgkaK64wsD4wnHl82iY8l4H/p657kSNNRWREnKVrsbYnX7KEpyCqe
tEWMS9nB3zo1kIzPb08mSEbzDg5HIR91E1YqcThtr+lY5GDeENzCcBFWt2s4Fc1O
PKDRw/RKhxQVzSaRAaXjK6dR/Cp4Co4EtrWXdarqO7yM3JFNxpAZXu2nTOceCI8H
Z5cvpvbch0j/1QDtBy7eLmewbQIjNN++fn+J3ggaBzn05DU774fFXaQHFnC41v7d
DRnIwCDRRb22NexKQXlkBsq5TTH4FttVxb0r7DZ9dk2d2N6OorBw6F3lUf8XtjUA
I2IH427otnQPXIDfT+2Hb6T8wFZyzupSWjcpCI5/b6q/sP1/eMcRNfMJT+1+Xb7F
uV/zAPOc3ymaIrmzjpTKvmYNLbfXhM4DZWCH03M2PWo62NZfKTErfjJ9nJhFlJKR
MuBy4rvub1FL4RpJaalcbZ5A6WeMTelJJu03N+IQJoClRVKxnkwNjY/Iv657ISep
uMz0ZfsFAlHcVd5RKDt7WXSIU8BKfU8TNGli10WjBB1WiZQ/Addgq8xKVz2Lg4wC
2pusfD3oRd9AxeBouTvEMITTcQY0NF1gj7WmQ/L2za2o2CalNksQx9ROcWfaSTcb
bGGzPsZtTAh50kIDJ8EMDLFnjJqjMfNpj8cmf0O9KnBS+SQ1owMk18io32ekS93A
Nry81lJPhWkDLH17X6E9bd/+U91ZQA9g6C+GR+Ijk7Hfxuf4yvC6i407k4Mr8/X8
/dJWUDQIqumc2zgSx6m7PagYJI0P4ppWEAsls1EU8p9OaVu0ryeDL1NtJ1s82hQU
/XtfwWlopXnKwFZjBmbngVlyP1NDGI9m2m0+/YB6655tyCgHy34RFGDnkw0vN9/H
3ploKiQ3FnEPqZGJ9MNgQpoBRVRU2hg1zBQ79um/nlAXzXwTuMziVy5UYyuEtzJa
CaWdedfo34q/svNDydCWLY/vz55YSHll3w/b/euJcpKiNPi6WfOrkF888u8Xmpdw
soE4NeixHO+Hd0Drbtuzd6ZO2qFfRIEPYxe9MpwZ37/qfIbTBoTCDXzLvjT1jSay
Ml7I4h0SmHuuMl7MZwOOKT6VcCzx4YPSiYdRMMhdWc9USt2F8FhPB9E50BuO2vng
59b9QrEKZ9RJUyheAz9S2AdVZHF8zc2/PrtQBQdQ4HKE08dyNLjAmOZXtglBXgYS
tZHaAmJJTHJBU1TnEjNr3UZOY6q+pz2iHmhus3885ucLXf50ZvwbfTK+e4SHCS4x
WBOtOJoXIwlFONxMipg70opO46xuRptC/2YXVOfK3wti9kpPoUsMzTPExHAtF0no
m/0TjWWHayN7TUSP3QZ+xVQPWURngZQX2WeNpwnIKEtO0GpeauiTxzEQGphhWXvq
0Ux9Q+hPIY1mnbLDc7ReHrydg0uS5aaENMeAdLXWtU6g9itSuIgBOzfz9Peb3zif
idf66F4IqTkbTUP0w68inJYUQKXnVT8ydtjkpnKcOo35jVYCXVdlSLspMx5Q8J1M
zZc1SxkQ3/bVO7IwiC0cbUya7bbO/9zBdW+iFCbLa/ubANqvCsq8SXyyXOXUGqko
SJ2E0IJVf7nWlbpmzxH5xWHQnX/qeWor/zjVMy0zp1j4Uws0Y33GcGLYIG/G32y0
KEeARp3E7KUGSbbJy2/2MmzWlo8huyqIyJRUMCMLvP60Xm2Ohayv5TSWhYV6onGK
NIdSO3OPwAOfHwcjR7qAsHWbEft1ZG7zAZhHTeqRsqVi/LO4Kn8N1fZPRCngIUV/
Y8YsPH6XcS46ReQV/cuFC/FkXTnjQqF/5hJyAb6lbjxIw2rd6BozV2lrWKfqi+T7
JIuftNfg9q57myfDCgjpbmp1mlbh53i7XYt4Mm1OZYvGcHtPnkuUVfB+sUnYK6YT
7f3uvQqIz8Wu9m9BgPOvSWcL0gx0EqtAaa2AZgahqTfbCqBbYOqj2gQ1vLOkxX+F
6u0eCYgwx9e3VCrTTU3JOLHa//ospOAoLBBR4JIqOjKp5ZFImERkKfTZE0ayshaK
UqZx/LSBU10KiA6RDSZ5BHERzNzYDKHHcCyUvy97l6e3HTIwDaK4gEWGbN9epoA8
hXcQ2Wg80O4huarBFluwC8zDUKE2YINtngGBjzjovrezzK1p+LHLKbzJKNlLCGIY
MkPgrKBOU1NPSNCJMaheCGK1FrET3O3R5JE0aIovLb331vdaHHFe6Ay4dDfNHm8o
2x9VQsjhtDPB2Ink/65y3ZT9FQ/fpQKyPo79DvTPMqi6AP2+WAJt/nCxidDJLD2F
xdsk1eR2IYjNvknioJNGBNF/RUSf2pIiDYh1lXXxuNA5falW1ERIGAQ/JkZKyA2o
ti2JvUHgXGkM+v4HtdW56hgt68fiA+PjRCE/HpR5UZ+feVvyZwLFA0YTrvWlFxyk
03ikwrrj63lOrpAeY7dpedWfH1zrfeSuEG4ybTHXDOZa/V/KyNI3Yv2RB2t8DrmH
C6mCaDX9Fh05umXCQDBRSE4K9zgeTl20nS5eteZP+lhqdiSlXtqChkw+B6ujRvqV
+MjbEI/unzAfWv/LpoBMCUgySvPfiaDDvz6J2+Q4koRQ4vxl5Kgufa2n3Wj2pjU9
uQ8z4YL3LKcf09ZkB+dUi+Y/sunEVrpgPhgpkmF9iKOX53vn2Z5IM/Wzy3uJTSic
KkwSq71FBVH3Vl7tfbwtz8XPkJQc/8U0IRLQAMxcIovDQu2D9y1ZmAl/gj+JRoq6
ol2zzIHkPVXnmd646Y8IRVFL0OSQrsGGnis0JndUYwIsGOWT6/t2Bchj32P/WRCt
bOPQE/s/FuIHZM4qx57bBd7qg2z/usFrUUKobGViYYAwS/gfLcjcJ2NRg9m42EvI
jiU8bQdPAhCURq/ppBVXHSTB4kkbe7svdOZLaYp1NQg772zTWOIMoGOgH+994HHj
5N7zMs0mGYJwNTHzxy61jpv84R2r4UD13n5jKtrVzpQ+0jXDjZTx5GStT9KFRZ0T
FGy/r5UIj2Q5iXs916sEXinOZzNIwBp6hCB4qSw9ZSusFN6lZ9iCwx4gfnHUuGT+
X5OjHvD/MUeN4CyzRR8qYGZ+6Fih/TRsGx1PM/cgKjVB5bWFdyoBuT0UkLotn9h+
AZhdglPVKqkysLhWN1vIwMjBWMieU8C3pEVCrDecmlKzAz3sIS9tEJNOt587zjjs
6SBGVbO501yJvJ52DwK7tlye+ncurSxrSEpqaDiA/1DPR7YB3LM+H0d8PHq3gZ0W
FoVVMoyhmww5fcVf3XXOqRabvHnPXKwFJLc79B5wPJg3fCQ5xp/y5QGb4+KlCi0l
Xwr53LC0i17rrxHeEw6cW+qcq5vB8XTxuaTy3bDjd4Obb4bjcawekH0s4sQblBzl
f6GK4RRhUfyg+rvIn0dQ6sBa1LclPgeJxdZ3Ou7chHRnmPXhU8ZBJtpGT+f+u7I7
Ss1O3Rz5k3VtXdDPVfcZu+BRDR5WxiKFltjaxtMhZotx69Rpjg7fxn0TnU6d8rMF
3X5l/MHe6K1GtUkGaJnGhSTY3jfYVE2kj7TY3/Q4FFGj9672xuXwk8j8ZvVbd/ON
TjvX5k+391DZg1kgp6RflSQzzYmXh5Okgqx+4vyYY+4DCIBaHvtkki5iwDuDa7Wt
ZfjvwkLhHPbjuKXW8qRAzo/ryOwykPtmdqIoaBDkqFdNzZ668rPS88gH0+dbLgPN
bSei1dcToJxog6597BLGVErko7w4kDt4d0yEM6EtuibLDytfFO8D/0v2LJp1ofR1
xA6QQOOAQ0eGhlEhSGfx3EWqIa0M47q/lv4oiq4SIE8KIf3HAN9j0ZNNkeWBZtd5
Mk0LYRKIXs7TFzryE1oKrymDRjEW/4hdY8bcK0RaAa3BTvjhvF8+JJITZAKYQV0j
68kt5krUtlvfRe7KKc3exWjNxSKzMInoh9OMOw0DcfeKZ3r96AUUVFxNoatckx5J
5EGid+e3wOE63GBYML/wxk98CBChK7ILMgUtqhzosRsAwpzVncGu/+7q1vY6+KjB
fHecMbNhc+kaVL6Br5xz4vbn0vekuooxca/anO0kkAj1TmE6NdlGMhZ3jTO6DkHt
HuVGJcjvHsi46HDUe173dnZKKxvsW1jp81fRrNdpzz9DgYOI30PtF8OOyYkFyBT4
4etX3UpVmrbuj7q4YSmtW0C8hCZ4n6Tf4ID4WWpBMNsPKWdPTnsDMhaS9mVEH+6A
mHGrZBQyt/baiip1toe3G4CTc4+oR3dlWWXnHpGRM/1/XXbVjBsp7HYm30C1Yj4I
EN2HEWeIvxQjCs2Sl+F4Bcoidg+2BkPHondW9TuUHclccc8AERTNF4pUDktQHUoL
FYJQ5a1B/UD9f0zWQMOVY/JzcOCTcB5S395iQvisdumsbS8kI57oP+sDf5Sh8Ohy
lqKETdNkZsmRJ9qb4gzbO/l8eYqrgL9GCwaLeQhedVUkuVWUoTBaAyyvCY+wfwhJ
3w2vt02bXIxL4xn5pk9FOPJXGZ2e2RwdEMq8gZ4MSeVJzxiuovuap/6JZPyHmDts
pE1W29SwOQog6Oj5vZ4+JUELL51ceBnDGHdDTez7cjmn7D3lFIjmWH3o+fmqjedi
hD96jjoBARJidEcA/vN2u+DlrmQqCt5bg8TILCUy2YbiLukkAY8kBh3I7SPQKcqE
mpxxreVDwL6332O91JVTFu8rlwngQ1XfjOURHF0XrPs821DOl9IqhFeNIbR3/WvC
bgztfOoyoXyTBH0yvtVh++V490/LITSroXrk7/7CYi806wlxdOWe86KYsqzFlF41
eADVPITHUQzxb5pQUEw+6SMKPyBoiAJFiceZ/G2gFRTnrIsOR6zUBoj3OMVmG8TO
q1icuj34vBpTbxM3ZFZWuIxd9fK2+ZEN8thV2YsXOm3Rw4vNdRMD17As/FARGOEq
beJZmV4qPeCkq7pRTpQzHR/O84DBjIViyaucsg5I4wAjFYt8si+PWGf0lya7QsxE
rBHmnw5ykfbt6oy/CLFm/+z0g3PhX1vXFsV7epIRtBqGatyI4aS743qhQd/YUDSG
XzjmTMmildT8b8v3yWoMJZTGW3UxABLghMnGJZvtr3BuSHl3jed60lpWfAMOiLd5
vO2eVpvCg18DRh0GWr7mPXe3DJhsxB6gXu5xdp7kFk77dkd5vAnuJLi7UVlhuvcV
IuNxoimWe06v4whTTFn+mtb8xjnAlXzWTXeMHbaCN/r3yNWuITZMsugnuYL4Uu/N
vMG+Uf0WPPXJySVSTv4CkKGYfkRVG5Q8NezRg1T5jZOH82MK1FXKQjLkMVwI1VEj
SsPZe//FNtLGoE4M5p3c36mZEQCnL1MdXyMAtPbHSjy3SGvkIXeppapvsGYwuCSB
sB0EbHMf6iJ6Xhtg4Gf9mSayNf//wr2tWWayhBjeRnu1wClyw0w/N+7rzGJj9PeL
P/BmrjYL8BZb6WE+Mryro4Ft3Vda3EnxwTFXOEAoYA4bIg1exBwhLCPc6YFGuLjS
9SFSfuT0vq7JfivBrDmB09hMf8CbXxsZeC2tdwLIPJnLeY+oLryBM+85qbKO4YVO
Wj4P6iuJlmr5Mje1AtTsKSiI3Os7aTQZrrFdbXr//lbZ1WhqQNIb8gDGPfP8vChs
NflxXyN02fCgw+CCle/2H3Fp0uHYR0qKOydxIPGVP05I12Q1znj8Ph00iZrBfaj1
zmSR7RnOxmhdmbSc9SvBG9H85LPIRZXw2IKAGy3yIisJ+nl1A20QqteeDoTduMSv
D1cVh1G9r2Z1GFFY8Y8diR7+OhHUMiQGhHjbZLQPSPoMnf5p4pcoDlSenNUWSoyA
AI8TkMXitLvR2CNNng8eah1DbGUp2SGAYT3rcXo6O833xp+a0hdr6xTnwnB5sbxl
vspXIsf0PlFT9a8e4ZkJHSUvEac9hrOngEtT/OHc31WVUE08WOe1p5Spgm+gQJtu
QqV4QwRHqpMXkbHI4bQa9GR/KEBb0lB56SlNhGI6H0jpKNS1TGqXshPwWWUnU1wh
TX09NX6kynI9PsNG3F9LX2NloJU6jIJp1kDyBUZZXZEn0E8z4Y/jRzYWXncMqyZ7
Z4zi9cnfU8xH2pku7NEaKQ/kihooMfFz6t4hgmT8rzwpt3w9yo6Jxc1VgyqaTwTY
HBxAq6Xo2bW0Ehr+H+H+KPUsU1X6KxpwkvRMxP2tXtxJuyxJJAMgizaJx+OmgMZK
YJfht90QcegaoyXL9+YD01yBS9Rxr6C64CF/NKiDG2EJpgw1uTxA6PC5VwdvYgxB
WZlwwvfONitd8CGGe/w5Y/+4LgKE2vDalQ+Kus0cPgm1SaWrHaESjV/pe8Gc8SYY
QBOCyYovIeLTPYjhAiFLzkXhmcdlfBlXuMye5vA0lVLCgTNtjsyKtliAfnl63AGn
8ECbECCTAh1m35H7iZ50NYVq7WlUqmAfYQYKLeI2VXXKGRX5gFWGsG0q+5pAwWji
J31QZWbPseYp2D21XF+yObg4uulJrOqnUGiWlbHAju+20N6qYCwgl0uxx30/y3Q3
I07iAc2rrqBcszVipCBjNY3G6fHFxduVYSEPKJbdezyj1/2qLyx5j2twTmF0SQq2
F1aBP4VbHjUVn5tBOjQq/j/XdXLskE7BKE9Y42IxJHcmoJOlZSnuCy0HA3iC/7Pp
6Nayk7MyT6yP8O5f4VqPJ80bg3GTSMSHY8USSHFS2qLQonAgcUKv45o8/LyGAV4+
4DAxs+oUcnctvkCFKkGdAQFJCGqoVEipz9KRYnf3F7UQBOX+clAF2RTcjNIGDZDS
PDZEKr+T9ji6s3/Qpiqqd/b/OsfiHn7agvXuFVtMmi36nmrlKpUpwVpP6brh/LUs
UNarZscw3W2HCH6OWTdo0vGmneajXm2MyRuFIBxOYxxUBp9Yat1ii/PDaxOinlcA
WihW1ee2hNGZaGKdzb21UU5TkJML3TQcWzxCiasSPTwT8RK0/9uYOkW321PpQKVK
457PrihY5xGhkqdLB3hNg5X0UpNmkgfhJrgoEugyyaQz/FiXgSYhkNAlIeh7cXDI
w5mokGojyOwNazvbuMOk648TOr8VEo4qyjyt4PVPQyv/UDdQWcidledFuH5HUw1/
BSgGTMTjiAJJod0LkslybHB5k8fPAH/IYyEBJQCTKV/v2Vz1Mj8yepClZFz5KUHp
9Pi1kgQFv59pLuCYnfNkTA3qbuLYAQ1FtiYWhcQh+rlNFM3UChCcOvZ1dFRSxEoy
UPpBEnDtaq7FFTJ3dfs0TbyZbFruaj6qvfBnS5ieg9DolXGCSOf9vnSF5amRgcJc
VuJBQNYNXHhThhNud5zQghyVEb0SAb7/N3UONYAcMvnivCqv6foBkI05xthm09Hh
q21pbn9S4B7YR4dpSzdMW62Im9rRCStQfPflK8JjKzbC2CP6/62VqEP9xg/m+eAj
jwHDk4okCEhK9bU0X5A76JkWa+ulSDrBqiKGKOaujkJ47xv8KP8QfFTDkf/t3YRO
ZGmZpaVMeUExhHv15+Z//zn0sTicH5TM7BX/ldE++W0gVr0l1/nRZojSTBwi8tU2
zrus1ogfeVlA7Crfgyi2aTpFEZfU/6kfO8I369P0m7+/dUmyok6SqcpQhEeg7eJ3
U8aHDU//p9w3Vmqbl2DH4IFwrR4CuqM4WLfaPfHxfLORoBCy9isZccOBT8AqQRBw
WI+DafppotYU+lA6FcVbY0r3zMa7As6/R7IPciKD2zsIJIN1rHSEI7/FyI/KEHCe
AFvMotj+tgwFj2kuPHvw6a1qhH8aEkys+iYpNQkGF1Av746Y5GJabHuB9SNoS63r
uMSURPPCehMcgPl6a+vwxowNisxYeUigeDqWkWbQedoMCzJ5bNxdPaeL2nuHpd6n
15JsKu/3E+bmiEmIqs6UDTUHFuCzEfQGcCLm/e5RoAiR08X5983BalfJTm4lAtSS
desIP3tp1FVqLFxUgb0kE4CqIpzmBz9bzo+aDcRH/4nYA7L9nFEGIIpJs5b0W0DS
wHeERVCC0mTMFdLSIkiGg44mk9Nd2J9JX5/CT9//TzxRVDo49DLA2I3EC42txMfb
q/X1VH/8d9h0OzGkgnDMneFufg05yG7UBVyMgQYIH4xXDSR+omk1XNCj+mdxhc4r
dczdXEhGc06eAtYmO93lUcNFUW/z8Kx1Cw1B0DHI1NfE286Y7o/v1shoY8uOAOQe
9cr8NlbQic5aX7xgDcPG2wcwq+jli6BgZwgJolzRq9wVsr5d8+mqfoSgxnkY+WCa
611PKt4g/qQHV6WBrgAQgfgWBT22zXRNbM6JLkLbp6vVwVDvlNxEj6vYTEpoM+xE
bSk9QFC0y+DZ1iKubADh5LXDNoPtWuuNpZMcanF2TuGYTtTPF/spCDNV4JuhMDd2
Jx+MqCRB1FIsBCU9vifyBF+BtsHm/wMKVgki0tnytHUiLlO9hjh1/qi3x10n2F17
hMuMwTFCro5f90axr6NB9gV/ljeB6W/ZkIYuE6rc8tM0duBWZVEM3noLsrQMb70O
9v9EV4MLIR+Lw75BYMB300Z9hZp6OGkgaRgAjKk0lEw1soHOOhf5FZOZ6gYLc/+c
bdnBOD54KIsyz+t2wn7J00DUWcqksYtMdri0pjx8zhyKMrxj6UfW4GXdHy5wIO1W
a32gaXhApKZPirVrUrTEh5YZ3Cm5imJvXwMfcE6syfhzH8XhyzK+LDWyihdmGHD+
ALOapBkJd9GD3Xwg5O6zUmfqY5y1oDHqGHgMNyheITcw3Q3F75o+tiY9g9y8L5JE
ie4f2skpjuTLLLLaCpokGjkHhFzhB8QR4BfWyMNdnwNONz8XfSLOQft9Ih2Th9P+
WNyAfdKb+zZ4FhYo0lBvVxV0GW9CkSVF5ur7DKR4iCyDHeJJ0B5K7noW9eePTo8S
ejNEWaLe8s59jC5CBQo5fq2N1QUxMXdCGiIWEK3xgz89CPki9q1kuE0+l2MDT8qT
VG+vBsI1GrTq4fWzi/dsNSDlEx3cnCvExJpI2dBeu8zGm9jVpbXipMc7kas/a+C/
t8ZRlhuQ6sId6hkRrhBRVoLTCBR/aLXK9u9FNq5Ryx02ia3tLxVWM8DWOa8452Xk
fPPonTv6bhdLmFW30vYmjJGLSoBDmYURTdKpxwKSh5g/83wos8I24B5FiucDL6tk
LVIZf/yz3/d21TVJwyycnf98tlc1bQgb3cGlxMcyGGEmzebDzK7spZcVyEixIDXY
R9lm42aw16DzEC3pvUR8r8kvyuPYR9pi6NRpx5eWcCjSzPGy8KrBS/p2wyE+pFXz
FbzVuXmmMS1t/QdTFw9MGOBEAm4DZGz1DKQRnuthDJvie3P5C6JyvCiQeL4bgipI
yYv5P2x7RRPnUdLX086ifY4tygRsBNrJEMUSe+VSVc0VX4QXx/j3VhTIp/Y9Xg0L
tqdecOKG7+C5k61gogSo89ub/OUexoYGny3lYrEPqUYJ2lDtXK97cR39H42p0pi9
COlV0GS2Za56XQG9OKpUfv13QncNgmCbd8NLQlF8gY1Ht49SjUJjEOyykDU/bqBm
tw+VAXVPPUKoOVaT/Ox7H18SwnSgfppoDNwtpjajKWbHSA1x7O2eC+mLgQw1gZMq
MurM+iCPs3NyRcxMoTEPdXMBvZ1b/WW154Fuyw/L/ssW1LjZEfWG/T6BL13ed6Id
pLy6ZVqTzIXjjd541SKSbySgS9ozEInvGuJ3418eaYr10uAu0+FHj6pDQ9ApW2K4
JcvvpmOjRzwg4AxtCIYBiU/hiK1nmQOD8Q5wnpLaEw2rySSw01fd3fDLu0B81sqR
XBll7U3p+9OnydiTzp90R18q51qmNyrvW2waMeZ5Us3xfE4rNlOI36cbFVuQxNFQ
Z0exil2HjMb7Wj3ptlNiPNbU0BxXTiGyw75KMcng5iMlkCQYAmNUQ7DcPNP9lWKX
8u16Y601dbSn5GMkBS06bYuiTksE1+42gX+gMUBXZZJtDFBeSWI1QWhIEee921N/
/XWgANp3Kne/H3Ud1B6gg0rEqQoDx5V9XVemZNAZ3Ci/RZGME2p4xB7IqLa439wN
f2WIbzk0MiRL7piDbFWUBKVECILzs69RKP7AlaLN34qm94M7V4M+J24m3pQhMx1D
zcwqaFeEF6i3h09O664pKJshq5OHX/01UPi9YczZR1sEEaXNJlSYB+CcsmDWCrJd
550wN4oQJEaggSpQ4qWIgYMNuR0SxOq8YzsoqrXrYx5q2rsySP1MjLOm8BvBigls
f/CD0vAxJDbEuSHYZovHhZT7PzZW9xjMmr4Kzrd2CEn4BvRVfw522Nc3N7iA/JyG
ef2uYdzVWdQSNJWdWHwEoWqWxcnOFNRBk3gDYLQzWlhUkg3GZrTYnX4WG+VRjFey
UFrbG/l/b9PMjkMIjqDU+x3WcPnBZjOrDG/yo5cLv6f2kfcvxFDdUJj42IxxJMzd
iR3a6U8oaSGOLvRUZc1Filnh1cj53t9tt/6QZeVPMqBpn4abO10tHZmLBHNs59Ju
rexu7wZ6ygMbExrXHsEwbGg1F++bSubfIgeJgm6uUiL22KdiyKIFDgjtFmHw6NgX
OIM3eqt3x6car/6VhTKU7gQBLS9HTPF0llSvExAqEGtpC9Od0WRZ30mjUvHwrplf
0tEI7SMemPnzWNNrkP2H0N/YjkyGKETQAtWAZ12JJAa2xReXILEuI7lp+96DewZO
/T7Q4220ldZf/LOykNIGEFj8hb4XYWT0veoWq/QM+iHGpJJjQP8Vi0z9jfZuNkKm
LuRwZNGoTrF2dEfYCQL/vLZanM6zQoUj8fb/HlJdoOI1a1bKtG0YFy+ECtZM9aQE
RWRRK0R5dfzmTyRsVNGcM9LZRJrh9TlLLolca494/6L5x3+dkfKJ6H+5UIke+Fh8
8AibaBb/Oa7Q1OYpQhQk+FgACeQJYpdlz12uVSq7YjPMaOwMyvgZeLOuA3NyXJdb
ddibVJPI4o+gMQi/Hs8juawH8dComwJM4FOAxSVuJgOs+HUYfMaw61X9IRgdQeEZ
6edS+MNnpD1W00wZVvb1/fq82v2TJawczoEPd05jbV5goA6Yyq9GOibXpNF6d9mh
OZDF3bhSHVxJH++nQhCHHE4WQJyuCovvWQdIADdAH/UU2LnneFHucvEpr8PIBO8T
D/kUvp+OrTewBXEcHome/1v/pLeWNfo4sKHNwgYG+eIi047BUUVnzxjOjU8cTM+A
9vjdO9yIJ2RhsjJhiSTomAT0dOsZOSNPtdxmPEIheLU5Kku0o/BOf0tFn2lNLeuT
sxJCXPNHfEA/WQvJmdJV0vHHmxcjNT+Gk4WrbafTl9lreXcGRYV4k+MYtzfF9BIt
dM/uCfZlSy1AoWQKSuFVMp6CASth1hjIoWY+HzwsgpYQVWhC0IWd+/ORVXZiTCam
tsRPQvaSABNJbDkLutkUMosyXT7iTTrC6LvoG4y2+OiXXXJ6hSSd+8AJLJt06JK/
7owH9Rwn0u41orDlHgPUXrSljfY0z1q3bozns9seph/fbAaHJdm8WE++toyknJtH
Mty/qD0etGooRpsCHLmp4a1wG1NtFA8jM5VWzXZXLxb96SLiD9KVDWEFnisQ1tq5
X9JfzcFNb8/rmcwBH0FM1S1CaHcfBZEXzl3KiziSNEhKEaaEs9cqot/UMCq6Ahp4
u00WvJgCBd3lNCk17McbyQZO2KxFx8EvuqW3G1OEJFqp0G4xKt8YOSjAocGxbPFZ
tCIm3zOpFP75ikS3hS/P3fhcvKOmVUHJIBm0/Ex0YUsV9CMWczeDh0ax4iNtJl2N
RiBhvfhLD4mdZSTrGk+vTwnwo6GNXaiBMtPOVcynnWhkN3v6nSGEwmCq83s5aK2D
8WrkwTEqcwMUdJANm72YFzsIWS7Dp9mLX2pWU4RP2j9jIYN85Gxf64yckSTApH9O
Ql0+TC79XOnPVSwcVmXdVOWxTFdkZXnkZhQE8CSrm4OBWlIXcxSQ6/cpk5wqBKx+
J41Wtyzn8O2tCx4f6ugcQDIU+G332AbGV6j4MmZtS9/VaoVIA427CBrvpR9Tr5uX
YN7gnWd+fmCf60+hOXYza+q7CdRiYvfeNBWS8/nXhMOtVnBNVuEC0kw7HNDx7H3e
aHQGq/ag+9KTblHyBjM8fynrzOdjepFpIz8MzGeG6sQQyHSogtiJr1VhVIOC8uqs
kk8/vTFoKMX9D5o9q0NQS4AmunWOY8Ha1nLEWDysgpZyg/mC+ykdbM74zaXFE4xU
UpZ0A1u+2Pp2iyMIZFqFWrQzAklCExJJXoPHPd2qyGJHTFlvdwUtfA6tjYUihTdG
5CzUHPRGfV7u4CA7Of5Ww6Zw18jidaUkM4uGGLBxT3iqMI8aqhgFmCj/rIrxHKji
GUyKwPv8AkftmaZSdRK5osRPUnzSxYaWDRWwTHXZ/yt9qvZ/wRqot/O31lkYed1/
D6SdHMf7cSXobgkyWosaftrsqLUeM1NbAeTEzw1msZaaOGtlhWfolgo0IZb8+mph
qMqomq1Dg9ie/V28A68Hyaz64pWHzjaSF3cMsnVOapuqtd28gp2Q/pXYUrPeCAAU
IBUtgjjxou2akFznDAA+Pjm3iUlyRV4erRy+ByXaNDEApKz5LYS0VecLalF/lwVB
gg3mgO6l1L8issoeYtA5fvCP1lJXHZJzsUEvRCeyKNTr4GwBAwobOlee3rUPQYb3
nptvQn26JqIwBnCawishNkBhm2WybeQAugaZ4mTDLvuy48PUCHW3eZBiMVb77sgE
CufeB0chQamY7qAxUmBhdFvsy5mHigJioLNSCSkSzwYJjGwDuLKJzDlWyFrqvj+l
vfUXHqq0nTKT6MXG+Zp2hoMq2KoSJKkdam6b/LnFk9oeLo/O3dyUlmL3S7FIybQK
alcAM6qe+qTwR/9LH8BHZ14H3vXVs8MwD37SSsKZ8AIk7mQB4mwbz31vX9rqQeah
jCJ6vK6g1XrMriYjmtKDY9F42PPehMI8P3nRPJ27V0nWTiJlM2L5IH5X7BKPd7K/
Jg0v3rUwz4lvl1vEuRxp+LQD7Yn1hcEW1ynhYKckvaTvUQZ2UTpGdboGeuMSnFCa
e451z1Dg4GrVJSGeRE8r8N3gNLGDGD10dWry+0RKih5GkvIVbhvCzG4mF1eVzV2k
Hi5wEQU36/kDi21fy/LYGatBGOBxQ5KOxNAmCLwjJMDWl8F2TAXN1YaY3LQgOYc+
484hpmoYtJSdPw27/CdnfhjNlw9qJSISX3u2UyPC+czBbthL4WmnAdpyHcq3I2hb
mAM7SVv+jt6QqwvaW0X7MHVkTjXZOUosrkNtXZq10G+p7bGF3GG29VC5NI7Oac0D
8HuTcvwYpTt2N7GFd6Irl2N79AB2dIyjcnX0nMbMyL+zxF+1pXThn/9auG/wKbTB
yGyyL3nVnRbm1LBblcVxtBSvj1mswtbiWCdBHKOfnSelme1QHC3WQW/1IJYqlXZb
axQpjn9CKEzScDCPw/cPIZHa3fOGArDEHf2K7poHn5+zq703R6nTZfuVlmmzCt66
rLHXSQAuvFvo1gs7BajBgqYSJOLENp6vym+AclZTWHQgYC9c6G3tu5zC1U97U0g2
rQ08v0KHeNFayVAHZ98047m3dFEXWLt+HvmWhYg8ZGHLb3EtSSfyv5jvx1f9zp5k
/wOGNZysecQ5UdhhpsdRDsUKQfs1oMgH1Vs4Fwm3Ty1mdU7+spJTyy33QL0J2Ytk
ygji0gTj7ytAMV4WKtyXHlGfTPhnOf82cVsR845y7jcu4VNXv1a/85W9qia8B2jE
SdTkzUuLqW2SnKOleTnX6MKfbqrfvpF4cW4qth5+iqGZJCs5HUogVkPF26g2BU/x
h3Bk952VhFb6jju1H6JKrVeQ1v2vzJpMByzW/FSgOf5p8D4RDjtpS7gQ6OwX9k3j
mEB2qyDbT8Bx7VTlE0kr1+aZRzDRBJmM/a3VGNM0qtIpYJBfqENk7xlHPVEeJ89Y
zankTsXw6johqz+K9b4zEg/6nwL8Ph+kayvxwyw4h9IP8sFhfvLTB8VMDacwo+p2
dPZ/0/MN431zfBst9NwIJpFF44Ahpe56x/FxL521Ob0TxsPhi1OPYdxXKQzVmfjm
uJbZXl63pLT15l//+rMvNLMOaK2PfBi78M28gfoyaGRhjkKtUtVHqzZCT+bInhhY
GTsjY8Ras5MK9izwsUHKFXqUJ39T0sbxKM3E5jphsn+lwTeInwtQewJNbeJR/HDl
B2xT8If2zyOvQ4jro/ekBojoI082Nt9TO/t7iiR6Alw+pfruPfiYi+0dleBsJkJ2
bzhyU4IgcPYFl/AfbY2nb5+svaa1qquvn+iNk8/skIszqoLY98blQYlXtU0YSgxg
iQYrhYHVGrC8NWQhDMrx5T8ycc6CF/W943zAv/8Wi3qykjXoIJ0pJ50QHfZu1gog
r3rsopCoNSNwThrhIMfl0oAu3f49dSkhlnT14MGw6X3Cq3xMEm2pCvYREynM1gRQ
Ow3qhamgnuQ6A96HWyEoHVMi8w2jVc92GMjXGd+Me7MhpdAQZu2D88ttwbugDiCj
KFjofwJIZ7F2MAcpsIZL2s0D8K11I8PyARHQwoCDpqjgZYAy4znLD6g6a7xUIEGi
km0Qc0yLCz/GFtQZ7XJYLrWCm1JN7MXFNBHIRtyzKYfuyLziWtxQJRXbtQCSqAyG
kXOAp8uKogA3Y+7k1uxZvGiAI/HrsEU5hD4yQZHrc6QIalANuJwCZeS2y5tG4P1X
BadrPPakLKfsr5IybafqUnApukK1GPUelH2GLYVNrHjVx75f1hj28ce6GPqDOqE8
5ipxZGByx9AZily90Sb3hciVCyjetWYBAU0cs914cqxzKZSjUN0/nL5uCaQRyqMC
6Mpf6HFrSInZZ9XXfogheS3pzc9vBvPRsdmS6+1fb9TzqMpqzwsLWPixwfEAJQcm
wRPwTRtqfbRi8RnjO0fkJfeJ2Rqg2T+Hz96l8qmgQPG1N1/q+9bQgQMP+QxGN+pt
Qw+9mmDNorJADPNq+sVx40OGn+sVPx2kJIpYo69YUVDTWy3ZyzvkaPW5nBbZosoB
2n/LMPsKxdMlP+/HKnFwgaEDjVZXa58vsRg08Y6ZB22Qk3annuBMWGrsvLrXNfEG
harYNBWGCsq9JYdcZqLBKXujC9JMAGys0cgNFMLZvD4GZFeZxfNH/wcmOSA2hwz9
ALBA8b7Ev1djUbaIjDwM8gjKfuZ58gbQce2Z+nDrXP27SiuSEM7LWswsD/RaepWR
dj2Ru+LqiWHA/M/IXU/ZlJh82R2CVxazL/wmWzSJthZEBFVsQJLbcSaMRVNtzddO
NGKzMz60jmGVDJvIcd/52n4v0dCUCix3b+xVwG8pY02EYLGSWZqySq82Scp2JRKN
jGxKpIudR9UO7d++uNbfZ3+1RSdaso25h5O7IZ97TUwU8vF/3ZQKfVOFMdIaOaZN
C9/U6S/HnAvPRT8LgNPHnNchhDCkAOEFI0ZQCNCdoI2pYXBfgAwiQraZtISahGLr
W+Yy2xUfERCemishmBEp1UcDwzGX+zVuCWOSkbEAohrKkxSyz+2PEX73l3+nY+Ne
PHaCS6pZhDFLdohJ4UGuhfqIGdsSUFaFKtF+j9V2X7a6F6V0Rj2D4Velrugi1rXb
Zk0GRqMasrBQ8hRNUV+XzMus+oAzMYX/+wFaokdY47z47iNvQ8d5uNtfM6xOMJRI
YKPt9TQa8Ss1LZT6MopsDrqcMs2VPcgrwEXc/8WN2e42FOiOBgIdA16Z4AbiSU4y
3D1N9L8aYd24JjWesW3zOL2FxvWwXZjWI/LN3rl6P/AOBoIiKuRts807YE0WL95R
1BOo2siDzSCDolRVmtYcEWyJfcIxkMbbm9JIc0qhIRh8PrB3nm1sIH3MF5LZ5HqZ
kQoinOHBZmvHnTVtei26Eo2aoSPrHyzn+9VyQu7pDEzO23DFBvGzhHpczrbbI3S8
HxGacKnQ4I8NTMmT3XP5apng7+VA/qGlVoXPO5NlRRjCyyTIOaYVKdB1uTkPKV72
J/A5O0Qk3G9MYDDwdsWssqKyR9hK9LyAimPvqJtP07sjrW23564x5Ufl8UMWN9WK
ipWiazPS2PAOvGgXS/opQmVg3c9Ee0X9Sn0ziRyeb0sy/FRnKoBEHEcEgkHOawca
CVSuJclG09tiKDo9GnzmJ1Ycz3C0tPZNJKg0435m4pW7B65zEatO2bC2oh4bxfqo
LDr0MTB0J074JBmB3VEZ55cj+JcfkxKN/GlcRflKU0vlXgkKn2lmCI6VxixC9THb
yBic4VvrJS1qr2YwpiIQHa23TTx9YkRq6ZUZf7hWK9kUk2yR/Joo0L+5fJrCO6CL
1JeIBS46tEUSqQLZowv81to2WBjrl6lPVor7FjQiEpcJE8fj+cGcfhhSuNHAPbcI
5R2eooXbPxdCGNK/nfLiefMWuSjpw0TlH8V9xEYKtyjZjYqwNRDS+UlcWVavbh3t
tFEDKYekYZGt2c1qO5WJslXf2Cmn+Jt82YAElBCa5fjm8Iep7oDnQyx49DW1Opsv
l0yMs5ev4PhfZwGayMH54Qa0BK1GbN47QxL7z9uUK2Oke11uHD1gpuO2H9YpRlbu
lpffxm1fEr7Z17vLWwa2qaH0nhgJHa19X8V24uWtB5snpi8q9KGjj2FBwi9NfiVt
WihT+g67QxYuhustmsMQTEqEgZcfciMad3MrOWFF5rx4NnksUqw8773XXXNRisbz
LgEyZu9NkC/JNNo7B+tLBAX0GtSq75TnrdNb0bfnypPJKTYV38+UqmaCWKfVlftx
cdI4li0XyCMLe5VeKG6KGB7zGa8Ap9M7BAoG3//B0wG3T3olbZNYEYcp3iQemJzA
LqylJLP/9+ZlANzrZFqD7+Vl105KRaPDcnV0cOYFf9ZqNVskSqpBU5yuBwK4jEha
Q5fQeza3Hro32hekgflmM1l0Ig713tZMX5UthnbSpvRvh4Zn+7cHUP18x1Td4DCL
Wj3oR/D5f2rl2T9DVBkTYwvf/bymPQkClJ6k7qgc02aA5hv/efYfLJruOhkO+vkz
GCGsxSSIA5ItY/BXxso3NMGFJUkM0Tv84yHOQvzTeZDb9kS9vuIIRzTZH8X63C4G
gdN5zDzgyHCjQKHn0vISqh1jQWHHpnqDNRCBgttpnIVUDV2rpiFpKkmQ0Iyjhgz3
XxTxeQtWCosnPNFe7ytKrvxDhBzXaNWW4b21BZlaG9UoUKD/V3z4jEYphedNW61L
jbYGqy/uR6lRcPdSeRaXsS/wbQPpUO8fflZj7xnitdsilbvKKGW1eN4l9L068pV2
XTlgp8QY7EdJH5J9WGkChEuxvSodgadtoq+BbQOChuyGd9DnEBUCcNOdJ/3MR/o7
+SIgGT8GdnptwTCSGh+Jcq6iMBiVAz6EeHglnW95Ki+5VgM9N8zewObItvNHGXP5
VL0USbqKT/mucUdZShyM7y1t2XfqL0Hwjwp03e2/2dW5p3lExEJKUori8rkvWLIl
bS/l8d4aeRrNh1zMjjb7vVa5kvWnPG3YkRq0F2PqkvZuCeJpozePHU4txKblxS2X
OAohMBa4UlN5SKVqJcQLfnE7C0nhM70tCm/lS82vH5Jv17X5hYvcD+/ZadRwDFCX
skOxzkzL3oVWGpHrpHdv71tCX1e+TA+G9b2Tf/Z8QS2TU8jCinx6KQiVNWDZBQFz
OGSLbwpbNyIirvfApP6uy8LiHdKll7a0cR/5QkIJz5wPww+AmP+sAD9FK+ftuANm
0j0kfEZFxlCg5drQlF1E6dmF/W6FBYsTyXw37wIVed6UcoIYI10D+gZL7iDnLDbo
oMEPqTv09bpu+hyqW7cymmDMSKUyuMnM31PYVtcsx92fRDc1FYrthHxEmSbMim60
9ztmoLzQoGeXODNNxM+a40Qdx4JT1JIgNLYV6BeOoBxTwiNa7iJgFxfBi7jZcUnY
pPdrHgjlgx24xi2AYZo4uAGEAEX9EKfeE9PpVG7XFKyY8QQmO5bxNIWYX2PCytfl
FSr6H55kpgU4rmZuBGJAc6d5S7tQwVZrKuclNhEq4mRcT1wAPmqT6JfkdBZu858D
l+7y8fm+xfH2VJH8Jp/J0UQFGQRL8S+qpTsU898kOD8Sm1p5juKzlZCj1Pw9nh6d
d4qjahyfLVc2s9/IsATtSPzOqzMZCqU1YuPTz37v+dJvcoJYE9vPCe6oqIcioOHt
ih1S/gEkn049+SVW/SfywmvsvjPPai7Y+gIcmKkT+0l2hRUVy6f2Zaj+OmJJ6rYL
ewFxcdV+vw7oVjHoO8162SPRGO1fbWeDjEy6HrcKHTVgEk5XOi85sMCwIGbBUmn8
HQnjx8g5MrpoLiTNomKnpngvrLDOKKLVqFhXWsWutcxnkA9T8ApaJdAU2Pm6gU61
4b6PsskPlj9TFVxg0do3xZGspOmILJWxNDCApNPedbwLVj2UmyKe6mR1wIujOYYH
5IFbWb1TGyLMaMYLUiwHUg+Wat1mgan8YJg1yrQtO5rgJ0pBvVNFgr9JHA4os7Yi
E1xa9kWvfPzSc4rGuq8E4riOFZNlBDtXbL8OtOj6oSyIlvdFRa0VzillfjkXWtLA
mjSLM+jlne2vonfhpkw0qaZ0CmGmp+o+z2zyag3ICt7FSEFXL2lwbdBNxgrbQRDb
/QGTzjatoIZgdLvfiSTu+g0n0r5EZ362FKGRx6LAIeYAxm+Efs6pVEXaw18gjyyk
GAC7MtHXLQX+z1xlrkykdzJsLtT/NmwjFJMx/bw8LAZAwhJxGOcdgwjKJBtcdCvn
6r8O15QnrsJlNLamxKuGqohiE+Z4QPyJ+ZLG54XaIWMYvfvBLi4ys+x/mW9C2Xad
kHFUbtL/gv3XFbT94p6UZNZ3anrrHGrZR6CE5yXkwIL1opNBN+q0FIPK2AXV3cG+
XHvzvrXtAXJGN3ZIu2D0u554pFa3GiccQM67nbIqm46XgW5dVRuM85fG7yW/j3Rd
BJt7Hokuw8SceXuUvAkY31XaQq3FEu2tEM1j92cnRQn9PW1CsWnTVe5j2rouKxxm
YiJnKBBtx7pAGWQS7XoZiqtlnytf3mIO+zxKMAQK22lt9UGeecwGfDX37hIlg9DY
5dlOrRCETfJycF2ODrVfNHwvqUkumGwzg6xWIAIb0+fOIXgRLlwRhBTg7RzXZ302
5MnZvFKImaeywmXylbeHa41aDeDJPDUKBArZD+VsqUNw+rykCeIWzWHYPAvMejMX
FhuwQ7sl99r17214peWyfTnYxNzKhP2AWJqPUI5q/l0CvkijNrZSk3WHaR+bdKEj
MXO7R9asLP/wIMxW9nPxZ8zRseTSnGa9nuZNuGG8X7BzJkxsiNvs/dArKQDtjVjP
N13BH2YERSgpQqvt/zFajE4RA5xaJKkVCLvuV4tzBfvsKvaFWg+hIDlKADTlujcr
mXjaM+XjPcD2fUO8Oy9i42Tjr4LELjmgB+KoKAkzT7k+WXm2xw9CO4UOnHsaI2p4
HCqtRH5FUzK5a7AxNg52lPTplNSX9nI5mFFe8ZnI++u/2SXlp1Z9WEGaQgeQAycD
XnyETKtd8Jt9m4LqxQ44pHUv5HsQU9uZxdL+1RW6GDOm52aiGXa2UVDWJrc7zsCY
sJYhK/C6xhRgDARMF6zLAFzWq3gti5aJaUkx13QPW2yWKMsscm/Adw8UQa/kGFAa
b2HcpFMS1BO1etNAoI5U2fYjwLDp+AgSYI/D8I2UEPlNj/dCmKg8Cx/z82dSgT4c
XRliPikEB2O6HdWoZJPpisJQUReg6ErCXBHSTWkwibf7hfEYO5j7PdYYAZTi19rT
+GUvXk04wJrijm0jfrlZsZqyTqAL9h8HCeWPYwHRnwY60OBPF846bRTsaKeWo1rr
Oq8ehRWgzS0CR+qNepPuTEmRsMTDuBYlYJvOchSnytDB7ibdrWO+1rgGMHmBWvGO
eJ2Og6AZ0RK9VJMVb0vDbPoWS9IiMIcNFhvK34qF6qTXw22729FCY2MbKh6ypebp
dg+ViRDyowWy2vQKRtCq4DnOOCgEUGKHHeb8mQvos/C0cqkyvQe2A/HaO2og7D81
PLd8z5n28QBsDG0PqjeXz2qutMPY2x++VKiMO1yINR2eUcMX4/OKrGq756lMpmYC
rznLvM99iJAvikQyki0XvOlNgmC4PZFfFaz5L6ggN0ckojc0zlhX/npLCCMyIab/
oCk3k+9kBzL5F5GXwK2DZ3sk5HxRK7CB6VjixmxWRlLMlKoEMVNBtWgnJOppNY8Z
66J3uGTXktQUvndSW84qiMnbkwzmn/9HIaHTElLyrO05+1tp+uQQ9x/l7cX6w/D5
H61JhxWG1AIAsPYSsvgHkqUS8++TYk8l4MlVpPAbvxXBpL6Jg/E5uXG5BWvzZQIg
I6BK6FdqXqQO6qop5/3sErFLM6WxeLROv8574PPhrHmMFuHsqZSeLIjwkZoN6bM7
UBdDsg2LHE8hst4l1B3xjG12g8KATPaWfEsPO5FXwJLR65R1bx9buXFTALaUuZoE
/TXd7hpaKMQQUmbHbZuRCZj2u6TXhVPxhLiuclr2rjnYyvfwL1mmCUPqL+5IIz01
GByNpTyVGjX8LBmLXr8tNZ9r4Q0JZY/avXHJ4EoaAgaOjGq4ZprbOod3FXUMmt/9
4IivyIhUeroRTCpPWHOPp6M1R/lZxmhar7vQ7a62AmMG8q3azic6CZI0mqcy70nx
mDETkoVcjFaBqkFflHbFjXCTE//B7NlVZTOQ+Nuhh8IFBhut12Etr2L28oIrVxoO
T/EpvOLV1Sbz9SYiihJPxlOUcUB76uKbOt9MYgmXNBaUwacrtpAId+4cZbZARU1n
/rZxzgw+F7soy3YRF8O8NJYYdg7KhnG5FW4gIPgq4zxzelMQggMMasxfpmY+LuD7
MS0OUgbO8pEv3J9LXk4aWyXdJH8kVtBi291yxwSSJepA6k9dzTgIYwUOan62CcLD
O9YyssFjwHs4aiJzocQPFG4qKXERBfqL63iYrhOLRS8fyVFWSwxFz3ia/7reF6vH
pCs1nX2d7PPi2x5qzpteSpP34N1eoa7OgqhQA/PM5PK10WKG0QZ7Yxb3a6DtQaeR
FgLqmCa+G8dPHUiSF5P6CG+aGXMPwy/3KlQpph7Bh3ItgUGYcrZVREsGfMp1rdJj
XuCVi/TgttY8i/Rjl6MWIZtBxqyUTrFQ2I0PRpYQVJf9WAKafu8PclflNFq9zxSc
SJIs3ngweLurOnZEL5D14dWEoLxQB5RdkqMlmW5aPKGc+dDd2c+p1TyrnURZyH6V
4iU8dCv0wv+D8mg9L9RzWkBmD9m2NzrL1Ez/Cm8CQffO53Qe/E2cJWDgRkUqSdo9
MbL17FwLZxMxXzBUU0BIPrNiOt0o81pi2uu5PLCuhIvSbeVl0pgSnvs54YaJIA+b
O64wI6p91e6zdZc4sgfGdVZZIv7VtnZsYydttoCVsUw/yqfuGzl225HxdAuQnjBl
/hNn8m6++Wm975DwgFZLApWqMd9kKXEpQcx3MvRupdT1ZWxcv7ReU4NzBU8cQjzw
fgFcVk9qkC3g4aiiAFSw5xId0NUCuajinjoTzSlAuveuYDr53gehRVkkaR8i2ENm
Z7V7eQ129xIjrq2mMm/CPD7XTVDuDW2OSz+dlOJr5cx+E1l3ouZU8DInq2lvrdVD
PA3DUeFH0iEg3qo1OV7d6VEGTAHZgrn5cy9JtSB01T4fCVc3qqw4uLIXix67+Yri
qc8+uDrMzVTvF1UxFiD6mvH2riXOL9y3iVF0Dp0yKEgdzmhoj5SuUzghxK5BwiwV
ZIoEXl+2Tp4ewsGNv6YQH1nXVeBoNBHQmKuDQ55qFf3Yl9cDBNMvgcfGj6mf2tCj
pat4AGiFhvWEa2IyLE5eYEMaE8EnlbXVc7sn3mi+8j+xo+vZLHkmQ1Cj0z6UkX6y
qNZw6Ti75ma/AFMVIGBXHcq9HmLfljCzq/xM8M7k9ANCWwWS26+mT3kn/TdOENAG
TonlFwUUYHA247jWDMg52Hig1/2CNNDOIFxbLrgrdmIdnMo9gQbFr5A0ZX5h7b+f
CXgbJgaSSVAKJ0moQ2qtFs52x8vzQuX+QUqS4Hpdgv0or6m/QQdmHRN0Ka1feMce
+HHEpYMZTcQT00khb5/CR3yxpkkQYTWiwlZPWkS4kRPazviKALc/JKDoSAQajhSk
v3FQCPfqmx4+PUsCAFJ98GyRJfYsrOxXt48M2nGmDqNlR4eQVzbTERJG0W3CY54z
d5j/mlG8NKpLbzJqDqQDmCAMM0zRlJlW6aQ2fpu27nWVifhLYHXF0xB2fABH2UMF
E8Kq6YVpVbvQ6KGlNxYtTp984S2mgIYUynZSoNaw4H9qrIVCDNg/c1inMqXEVoWE
/pm8FRNG77oVenvCHHlOv1v5yRtRVHLGT6EQzIaSfQKK9qWzw6QEKXR/vbKrAUF6
f63WHlRfFoaiCrXpBS8QIN8hKXnblONUE0O0ZudOMExOQSjn2YBroRqavYF/xKie
nirva5DfrMJRLBnT4NsKGpHbkcydbLlwrVl+PeGnLnypPKzTMUP6GCwtX/ogkzoW
3Zija/8MbFpaBY77kOQTOOEpDrfABrie5xDU1PSFNmnR4k0htVIKUoTiYkgIpuux
+FfGQRxY0bPF+QZqCwyNerNR7ZflUimb+O41X3S4+j75V9SxtTxZyHRHkwydgT/T
rZAxFfFqrNfNKBHjuQYao0OXUuXGjK3TLdixtLF+vn+UPw1w9yAXwoN5dvCcTB7y
385tf5qNbx0micc0Gw/C2o5cydT/OFq3GS0md4z5dulwAF2nU6YoIzw9bCmQExqB
sbVMOzYn60aO4N2ivQiUWj/PDAoo7YIpTvchUxJ/GNi1vc+dmrpdH3TDUxhcqWm5
pyzD2cSFUdIj2DHW+U/QJOPvKeUvXETjmIvePiu8u/9Pz0WpMXG4ikDm74EUdp3f
2gepYZFDsUHFiBkW8KKmKYnVyTF+VvI/DmqKSTF9iEOxWG7MbIwOUkuUhgsmaTQa
KND7g6DnwsvCIq0EWSPjdvwI9eH+zWY1r0aseXpwM2e+GVH1vtMfcXKwHQ1ok7im
l8EnkRyK8X242nKOQpwu1VEaE/F2YaFGJP1hMDAdIB+IXZocSkYX9u9UzeMD76CD
/rIY0jbih0YQC2RGWL3D+c6XywBs5/J78P4l3pnAcUnV0ChmYjLyGQ6ABiWJDTzg
Oh1+7lM3+VOV4RUarmbPDud+jFXDt+6RDLTzKb5o1tKeKi39i8T3Phd3b27PNbz4
D3XJGcZQNTSV1xkoJp+lZdgI0xKrlrxQthI9kkw6/uei65ofNDWbCaZsfgJsYkGy
y0tSY0Jr/38mwtYExy8JzpiVLgN8LI5eUi+AXBtjkUW1iX4vLAT/L5lvFwm7atIc
fouVr0U69QbkzTA/jzVLufDrvTWJPWJjsSahaxsp1gJGNMfaodQa7ACxxOyaMoxk
R+IvO+fw2NE9Il1FgzLn0oPJTSLzyNFsb89GwnqOxWZmkGOCqPt4uo+aVoKZJAYq
0+ugvk8kI2dcCwOWKw7Su5S/qvjHgd2wAzjWPRncno0kzDYoIWmaYTRBYaWCnrmr
Jmppqgo2Adia3F4AuF/soMoMnnrLO/uA9xxfcQkqAnMYKRX+AB+Q6Gl4jMDuTaqH
KJVzck5HD3JPK39+RIoXcadYh9uAoVou87I3d18XUJnLyjPUjGZ+ztFx1IPz7M55
muyoIn7jke1GNco6lJGlOZ+3wIokIYx3pHtb5cnZY+hDwXEllBvsc31gF4K1/IWR
m4KRzxdq1G+4Ep6PdeR7MKEZckOeVLVvklKWJVH6mDeW37/38HqwtzS4rkHuvKaH
6hE9hZqrcr5avoUD3WjTnCME0i6jIQ6GhOVzpZLwlj/w7Gj9kdocxjV+bQ4u9jqR
Wm1/z+nGwhvLU00GK0RrdmLgWIb0KiKNYQa1/HoxbtjeGHAzG5cJC6F4lUCdwDCx
v2+fGkEUbX4OGfrePZp4/+rxmipk5BbMeYx4HXx7uPNo/J9PpZ1K7VK0zyAqy1z+
yPoQTpHoDhAnsJQn8HwdtkH8KvkCCckz3un6fhtzk00/7a7+4xM/1xZlgvcrnSug
pHVsvOf7LlW7ErldebB6P7BLs4HwiKy0nExmO9HCkFALafWkRmbhnoKFbuKgXVx/
TfiT0b8H+81e4zvp6VA+2FvFNGmlFi9Nvqa+nkid2JNf/Md/jpEXQBPArNjB3uod
82eGjk5p7KMTO1/Q2x1aTPpzh68SSev2SFvXWT1Y/qZmXXpgh6bvg4YDRk0RWF9j
7cZuaGZnIwYOlSjal99N6qbyKfrrSOgZADJ7OzzyUo+f/tj84mVbu9Zi9yCPtVy7
0gyv5/JZozUFpoPBjbqiQyvbBFe6A2sOfyaUkqKDPULkCMlreudV8egOUGdBti6c
RA07WtHJixxHWqSihj81vdB6ZafkVdaYmrH0EU+kF9Iw7uUyZSJKSEv75A0rwO+n
Jf/IMP4j0Uxle40oetmrYiG2CjdN4dEpRZkiiBz8gZ7O4xYAPOkrexpzEn/OaBTe
agrFbfCKaYkxV8XAygLxrwn4v8EcMxhh3NUfPRElLR3rF66PwRs3yycQF1q0sCpf
QejbtliyQHHVWvedmdL3jJDDN/41pGRuXjW4m3p/NbYKKh5bsOYtYOwkEXhop00Q
q8yqeg3JCBoMhuTfTye+J6MS4HDWjR7GNZKYNSfbk7acC6lCT8WTX0z+iW0+Wt2z
z//1+mMIbXTgGHAgavcjJQB7hcVMVR3Aca0PvfkiI+6spDygKsweDbnwokWzmFYr
wDRM84bXWfxtkECRFoeOM8rIn8LnzWqxSRcONWxHqZSzYD8lA0OBsYUDqqkliOTq
FTCOpWvM31C8mtYGj1L6n18mo0Ju+iMcSWNaPgda78O34GNObX/+yn9M+oyHaXiB
6EeWniqlf6liy+sqHz2Q6KJikn84MxYsFh8cl3Furd960c+SsgqxvKqZEvbBPXTc
xv6GQyChYox1WsLm0Lk66SY3MhnIFYa8qxBbPGGRMvenALHbtZ9clhLTGObdqfr/
3trSZ7KDlzh2YJLfaJJtn3QW2dIUyeRqGFnnOImmN7JtwTJodCWKj5z1jtPNtAtq
YxykNwRfRwcFLrBp0vjW6jjiDC8ct0mSuXIu+MRV1A+UChPdxHbjDeNKHmHm6VLz
YeDylXBTmROSG7vcHLrCmhfURG4FxN9whw4NvlnGGvjcf+umi8ryYak1XjjMuUlW
LffJ+0mJiPdFJPkKvYDTEcPAsSPdk2H4prluzXPVP9iSUm4P/ac/dS5eDMNt+JSk
H0/zIcY79dUczi73DMSg1DONkDOW/4khPlxqX0OKJQvtJrOiMkfojCCREHAPpeJc
He0P2EQwMt9hw/egQnTT/Kjo5962HyJujPjjnvXdxptql/JotVtlg126Vo/qj+dG
1OVT4bZJE61c4pZLui9VfRhMmKPnVEC9G2fXR0sOtbvMdhdRdtdZ+FWPkThmpb7j
0mtw0hIPuLlfQHIo8OaeEbSvhQtDclc/Te/Tz0XwrYABzKh4iQah7RsJyfL3xfdb
XTL2UEqC5Kpx23Y0gGjOOEjQ9Ta8hflaiAeUAkG/tvefUq8jDwQKskcJGKiTrJj+
YWvYdoKeFlw91vd7cknKRbcnXBkEFmecv2gr+CmED3IlwJZnpjTMDKJ/+QVd8ECQ
mMbc2wCTPUDi2e0dIsmBxYF4sNFoVjtGqKQG2h6sGfUkMcM2k0TjC9XQT5a1aJkZ
MFjcXDpJjJAK7xNHbye+CMWIstXQB1R/x5C5PZ6HwXI6glndzh5xlzR4+Jue2pcV
V18+lS6c+xtI9irCHdoILIixDXsaYA9//GkdJ9pUBfMvpVo7E7ikCaK+/mgH9/3n
XVXak0Rp2RrrLTZh/sz6/aZMTOdfjdYSlvk5CZ0wUQWbtUmBs/UG4taE5tNAE9KU
Xhimz2o5ouuMoL5RNNAmTwC7Vl4tQvu9I7BdsiXjRkje6VsJZXXIN7MHoFEPE/Zf
9DiwXmnVwXrpEpcBMjbOs8m75x5cJLdOanlX9fmiI3v1X4Qy74cHOSD8QP3Lgh6m
pwuGuBywc1XlF8Y565AB4cw4/Ntkj7MEnuPat5gkPviRwM/qO6EQ/WLx/pVVQ4lT
I92oDB7DgJzEwV1oTe42jxZN+m2PZszYQFX8VVFvcr/9XIBm5z5KTRFJfpDCPPnB
lQ5sHr0rklLT+p2+mMurRtL/zFXEJw1JVfHlpB3X0/Gok8STPdRX3lgA7rEYekFA
bPVwHWyJq+76AgSdmoxiWYjVoIKD4vUtZoYaYtTgYRbMX4uXZh8TrHfdeEdsK8HA
PMWLtZjF2zvYvfK/3jYwKUM60MFO0h2R8eN5eZEpo/orwZptRjMAxCuL5Z3EAsvl
uVtOm9IkbghPDcZjmC/D9JdtgUv3m5CNz3YEMy2DHjTna9g2HSRCtmia30YV2CK2
F++68MdCaGxgkMstG7VxI84oGwj/LFrtuG/fQrqJegphxsL9IUC7n8HHJX3OPfFz
USrLr4mrIRfhFsyHWoI2ezLxj7KCNDUPyhFQLWzFEqsw8s0FBBoDEWlaUVfjBvEE
5fahTwe5ajZZ8SxAAwvd1uXnzpRxBXSfbW6tWkHTFZxFyz9q4b2NXt9H5xbO6jWz
19XMVLKDKnyrGvxusotc1aJPb4v8/4QNj9NUw2LRQlWd1h9SFAlfSc0FYi8iGsJL
IOYdOqbVyrKG0zawN/WLIeAlaPgfzKNuGd1VXBEwIYVmNAA/aP8cV8fn1o2Si5/I
5l5CMlyKBZq7DcdX4ahE2QJh3YeVyXi+gjQXCmGYiqBwTBDj+5AXLl4XHJ87vra7
o1tciJ9+8bZcFT76H9qk41UwNf32EbseJCL0gQhMiir4FXgfAESg8+ahqeOvHftQ
mFvooA/Qo/88liRGDtGZTVvAcq3fwvAi3nRFbbOEJWsqxVr/8M74KBr2Y0bvP9yR
LUAAK/mDzNkQ5lrZ60tD6x8urExGndA2xizqqHZlfBvkwNLidNQS6tqaoGWTqJSV
nVSoydHhWZWd3hekMn6tcz459RhusTGV4f3c9KTyJRNFLguGc2C4JShHEKsHBScU
IlP71FrD33ojhIaJ9r1RxYI6j7wi1DvVY9zdILaOFmBAO5g7/KMb/GVsmeff/akS
vs1bGcd1PKM+c9Zb3VJPk3rc+AuywAf+9mEiJBjZ2Bm88+K+U1L7CeAeQEfJdo4w
FDiUamz6P+yDmbkGqa/LJBU91QLDMcf+ISF7cPU4DZPbP1OfWmpLqCBPk55L7LYG
LX8giB2cYiB9OoiaPVTw08q3LwmrNqpndU0cZxZKDjhMHHcXq6AJle4pWSl5u3xb
p4yaMHGATpx/NRgGcbBiwoBkgJiXwtbXWXdycCHBeG6taNzZ2XdPfZdzH/shgGR1
PtwfYpf5VE0V3ONDRuloZJAaN4gRF/K+gocMY525cAjYognID3srWFNvexaWmnKE
VsTul4CNVHNkK+zDxXDwrkL900DAAlm6C/uyj+c6UA8fr9k1sBHFwXDSrpcSuTxu
J2KLaBnXis7uG9plNt6xdaPd33hGrcS9XjgG+3RGVT/UF/T9KB28WjwmGbgzAsWe
LLvuUV3vvee71qUaAMMw207+gq3k8WvIL5ao7+RJ0Ow795dT2iPiaMuhb8ZgyL9X
PZdr4hwhnfAWvxmQPIqR91OR3LTBhRcpAgE9UbaPOSpRJe9fyDwEbQdwWuzGWF4h
KO/wujWiAkfGkiOCUaC/NZDQT1+06ZO63FQV9FcpmPAWWnSz2kP8oHDF+2pTqhZS
ur5si7mZ24jhC+3MTsH28p051O1kDlOIwUh+v8PKaaEvYrmJhNbwgn54JRP7QnWa
iwrAZvLCRn0++sYtbKmS4krfeKUHqqLxzi3FsauAtkGRkoXRM7tcguXJCiPEwInD
Gw33Z7T2AHbZkMi2qmYQvUL6ty5cBiP+1N+RTiURCT02W83jLpImgJPA9IqVLuYA
fc0Ax7KxpSBGssI7cjxrQR8PLQfSbKcBLbOz0/KURHZVZa/+OMi5Sie2yf0zQCAO
SOqFNQp6aO+ddS3ssnx6HYb6fhNAYSy3r6yv3grQ5E3BWqq4I/3BqcPWSLg85/bz
kb4fXvr2uhvWMoevdaZJxLmfTW1/qBVU1V55W5gDtV/OleodZrN6SPojFcV9t+0F
LbyL62dWtqp+lEI0ZvCkXC4ry9NRHcXUFdmVEA4MovHX3zTOcSCyY5l/3S8GnKnf
HFriJd1RIwomYDg6zoka8JvUlbTa9KVPyx3q869vZ0dCYtneYP2hPs4UKSWcSuUp
GUx8YpeQFHepTgYXQvxYmF/N+SduLwj2NrZxIKFKnTdnLdD3b7uZCzpsG9BYwQlS
J9F/GXfxo8iXNoL+3eRrMUIPt3/mHlHOe7hFG9uloRzi5mlCroccIaSA0nJr3rxa
rSoP5A0PItSp9+Tn/UpxRzRv5+8MIf6FVEAgJS6d8J0uSh17yVBp2aU842kqhzk6
nKHlF2SjjncO5XAvm79t5iDAmoFAQQW5SPIp3ve8rqjZ/tZ9QegR7mDzX6kZfPcT
lSUycN12W8t8XrQ/Qk8ffnfJuMC9neqw4WyYraqtBhPqPBbpLG9g63wGezWhPegq
Cp/uibwHzauWOL3ZSMkwGEgSiv0UwgEIp/gaD27SgzGZaGzMKMMWiybEtkGXU0gv
JJ5aSjS2X0Bw00/r/WODmruop4B7RpnIC5nedYLAN3U8zyurVlVVoap2CwP7/mxO
3crTuSxqkxYkWWQQ/Ifpy+HvhN/xj/32nh+cd+kioyaQV5+kznGchZhBrZkZa8hU
bMZDR+blFYGMO+oQzoTWqrA0zfKjbxfvMKXkONhVyX4207o8cT6XBuko9p7r7uTK
v3XK6jecsO9yIctDvbPAVeXxr9HcmML8CkLXlPCRpy91ThnIOeWPxYgO8414r0hd
shE5L84R1ZtLEayssAxBL+9xwhVBRgA4O0E6VROZeISC38ZgDF2gzutiJZlWfM7f
sGXLk4oOViJkAe0Ho0cVjjuJ2XE9y3AlOY8ing9KLU1ZHigB6cDgfBfGXVfHbH6D
MF98TO8YAweM7jwTaAR71ESw0Tutlp746hjA7CHhLEecK1Px9AffOWesZTkAAVOv
FMSkJHLlDXDJXumZZ9FA6BnesndwQ7n5oFBER336dzNRSsi9+5lvXZnpyR5vgtSy
UaMtcrv9X5P2A5OYq0LEPH4PcdquPjUWjegPBtrQqi0lWq1fPZ3t31DNkXD1wYwk
BG9D9g5MPFk3rTilB6EzJM50XrXsfMEsaKRc0kztCtODO/fB9ey9dzxM5GSQQnd+
L9HkMDx5DXbRJXFLAqwQwcJkkJZpFyYI75vRhP+jqBf+bUA5kUyhqyi4VA/TlEYn
BnA4LKfI97Hg/cl+Was7SxYKKsnTCSc/KmhhbyR34NkxT3RoliFZUx7YcnSavb4b
UUi0qBZQq7OEOny5uDrdj98RJ8P5p952Z1tS5v7QYHqOp+Sm3nUoVk2+N4B1b2O7
T4JyldexsqXgVVgmnbXboZCTkUW9EwSTgMVVwSq5cw9u6C5YFtPuii6q/QAWdFDA
9hOH9DXCwnp65NEHOW1aBiXnLnDLeV47YcW16SZ+jn8SSJ4u9jPMGQe+LQavdm/V
jHXZr1hHzn/FFbdDTzm+Rv54xaLNcEsVZHWgenjyygQUdap2ApzhWCrvvXr8HGMC
1D0KdhmaUevBHRfdkwtPFAdB35gHmcB5Rek1f6Nwo9kYVPJHzHmx+2ig5OvHm3xd
zRFjxkRO92rt+Ee+ASdKyPL73ugYXjdfA2CS1hbNY/jR1ouIYbYHXZwQ7b/h3mJs
zsKDWmN6LkCw7P64CR4gMWRZC5X1chiXZ7nck5wBsxx2dcsM0o0LmnWWERw0oJdK
0hAeoW8SqBPPT25AfFlkqMoxo+LkU9FCUdFViHGoDfAsmgczmqS03KmM4265UvG0
+fnfxLAs/hiMMGSdCRizeWyrz23Xgninp0vG/9M2DN0rUmPwlHT8vbxn8lGBOhp/
z4TYAwTakE+OFQFIQcsbf5sSnY8NudnXVYmKyGFmpEcyl35Y+icPApcP/COSVzKO
i++UXIXwm/DRDtnTdogjLy/w9HLSzywCAOK48gAFphbWoli0/9KqYXEaq0+UzHy9
WQ1T5ifNs+TCDB2NiNllZ2kfxn4f9VSF6qqQTJEFmtXxoxBP9f+x56InLwqin0IW
nmTJ1Njk4d8+mT/xpTqk/0bhVr0Xics7hVm0xxhsYZU51F4ge9/sezaqSG54Pl8d
lX4kOChYqpLLjz787n27fgECo4EvlTQGEcdfyt4lanI7kWIfcIVrQhsvEgsFwOju
Vq/2AgHxsbxuOR+QUluhLWawIWeae6h51XEg1LtsadgbhVieeSnHXBU/fblrVwcw
0Om7z76DF0l9eClIw6e74EfHp/KXjMJfIQvNqx0LFiTYNkUUgK+jfRrVYl3qCfJ9
FLTSg2OIcPOBq/f16kgLPl92jSRdQNcdcITp8vd4l44SGkfw8etYXaNA5eNMBalH
PljwvnlUjrKv/uEwNdNdx9xPwjnBCUtGUgDOvDcLlXk/XYnL6xhON5dpYmtJxku0
p+n0WdRQu0dJP7Qv4ELdw68SEEiD2tMJStUYwuFC9l7T6vTSmkayWvW3ZJpn+4TR
pSsO5GUONVaNJ3p9FAZWZEIBGJiTrdOoh2aZTvXAULlWllHEVZJs3Eq7NFqNVy26
lwG+KDzXq2i/SPopA3EZCfWuQsyVDHj9PX6LAXP/sZL2o2dhpX1ANxlOe8ZYMYPt
sD/ejXA8rP6VuCQ4PBK/WwNXWLZUgS2vlnTLlXuGDsydx0J5bVqSzk3VzgcjdITk
kG7vJ6JTSfLWg4dzQcjWKZjJ2qYtaldZyeiaq4LOrXVmbeq3U3xv+ONO5qGE2Utq
5U1J1MeFgwQv/z6834Lle1jfJj39IfIJJCtpXBVfg6tHNVnqn+sRnWwpIMBJohRx
M8qvodsM2FN0eIY7vL9Nher82pAtcb5SVW1H8NlC7ffkkKl2FuayrYQqSzdhiZOY
9Shd0oMEYGGjwooJm0f8sR6lKNw2FM3b0vRcu531Q0sD4LcTRX5G8wYpTjHHpGp0
4hIyJQMJvJThFCFibensu4n0l0/WjsA0ydAnQRMPpafFw41qQD1rA9c0eCm6EZy7
GJzBhivm7RpNtUAGSjF6Vs7I8MHccstH+UJvpsbFYxMq8zCaFsnQw+322H9luNJ4
I3XBVHZ2lL4zMky/c1GccaUgJqIaI5yg/7o1HQB/jAD8kp0IpZTsHzYOMuCm7BOh
rE5py17XfgcfxJnUGO2MpvX84O6ikDjDwRQg54IrfKU7lvT1uKuOHTUgHhiXgtyO
yq7bGURHCEAA63Gu7Mp2jtbU91X2wk5rIbesrW+0+57reSB3Lt2XjlkLO1I+/eX5
BZY5rLNmsEVTvrH4f+IwSQgMRg+kyjd9En4vkw+e5q3Kdpy9Z+q1/kKX2ksveSbD
i7SZ1wYFXQ6orpoXc9QiRw1Xjzn3C0RpoHo03aaHABqtHVIrlPtCm+ezAwSIBjpP
XcqjtYmHB7b3sowMrI4UXWMFms1fFRX5D55lmwRJHCsVYEc691HalBo/RKzcBBqy
ggnAUZVXH7PyP6z6mwxZiXbI3k3m9to7lQ4fXTNMKjkcgwFp4uBwY2XWc/2xmA4L
XT48wie3fPWS2Hvx7IaPeFyVj50jBW7Z9Ku/z7SaGQDaYDNmF0+BPYYy2bFKv7SW
L9hz47rXUf14PKjLOnxC9AyhoT1H3a0TejQbB1/IpzWsdwybimbN4ct2Xvg+8VoG
/3K0iDmx2LNjtvwUzkIQEIx51jGREvoQploFagDT2vnK2NCW6jtyZetPLXQf5WNc
F+d3gUPzKXeqCsxj+uYOQbzYCXskhK8cLgNqWGnWn5Acn29O4rU4Wyy4S//0fuzr
AviUUuBfgS38lRhJDljimMFspazJEhMwBvGGJxpk4zu2rGi8/k41Zhm01I9sv9ta
CcvRmxbhwgK1QQ8P43EXLa9NClmp87mWNPJFN2vp1TbQZQhRtLdoWFJoBiocV4Ce
yfd7gTSSfH/xlMWeSeRtIlUVpHLc8imtJ1GRa343eJvQC8O+btwaV7amyCAs0iCx
gn6l4MwTQRRf8Tgz0cegMSQCngm5Mo1XLK3doEekXUGXI6zr61Ldo/6O/4FbJlqw
UYd95aWZPV0+SY1QG1Vw2WR1w7RbRUx/6sasBWPc6SLLHg9eofvw/YHFdsbsKJko
RdZdPzMNzrVv+ueOxV27LxIYCGsuh0ff0p/1AxJqEqP2swQYmQxgXCPF9IfrJo30
cvyxALw+BxINCp+BkQvZ4A/O9rzxNSKVu9pPbn6UQZeCn/6G9WGSUomVJ6cWm6Ba
eWhgiAqwmVhW6zZN1Hmpo7l70MipBvmie9rawmP8n2DLBTcUwXo2vrgiZc1QHvnd
BH4aLGZZdwjJIWdOZ0l/41yTADUgGecv0nzpB7FosHGfvw3XQ3ph1kbKzMed29aP
NrsXw6oZdlt/tYRLJ8LPuApwEo4ax+OECN26ZN3TpjV1v6MFpMqX8Whpnm8lJGBC
fvG78wdwUsz7H9nAmrUfUQEyOmo74bVgBpPBnavBYuS49O19/BRTXehBJamwo7Ql
EVP1NC5GdBuZycL2ux4XD1+KUkEGJVxiT/JkcZrYcUcxTcwKD/PJqO4ttTVZV1cj
L2nNaVlUwaTPeH7/UsYu/EHzcfxptNB7IdASMDUiEFGVa1EFtQqSkLIGBNPnoiQN
aOfTvvRx/PnkEN6iKV/oOefIgv8PkCMeaVad+gkxGACyhQ1sZNS0Iftax5xCMpKx
GWPOK4YgCxHOr20X8wbO+lapPri+fmgF4CvDbvRKgCx/vY6WmvGi7TfLNrS7Ool3
O6D6m1tgj1BM9maFxJUogbZ5dT2AlmkY2Q+bbYe90My8FpvONa97iUfQr6YGlBsh
D6CrRiOBneeLyBx+kAcaC+C4+uwhiMDL+MXWJSHZkxFrADQVZ8/wuBZSGgHWz7jb
7hFHlDH3igq8cnUd5kTBt/v7AlX3QqNr56irIBYkUytqj9PRSXW3jAvFy7YmoBDl
DbW95wL3XzW5ptP2CMFs2SPNTdEpawAOMV2RIBEgMBibMUVLnxSAvpBPhFFDNpIo
Xsj33yoIBAO/vIKBrNieAHEH7iADpzhvM1qKiBkaLEsUiUSKGfh+pOxCP6r00cOV
7mNy2bRCFGqZYw1DKNV6xCixWz7zavw1ZbRYl8Tn1L1TxsQKQgF2fUB9EQOmro7I
PysKGK8Td4XM5/U25c5EzIuhNXxnkN9jhUmtT+ytJXT49ikaCEC9BnF61V9GHHOG
y05IiMXxRSC9QRiTVC/JNBZq/AjVbs0M7xxjfxpEAFzeBD+Et0gId91ErXH+aN5R
K1m6mcXtxBdbJPy0a5VrYUm2obIMm2AcEBmor09aPCvZLGS1yY4tYI7YrOHrMpi0
yw3+NVa5JbEbZM4BhAqlAYBjTqS8uKMe4ehN+l+YhJ3EhwJKZBIEdVGEdVnA6pmM
oK4N5kddrMOf3nnpmQy5n4ENWqmGrItNWcmTYffFrQtdNAzMhBMdSJ6Illyx1OBr
BtuIwBPrHEO3GJp4povGopBDar86x3gKIWrVQU4FUOT/DvJUJxHH31rw0XjIQ9Si
n5n0uGqYEGNhj0lwoktNPSsxB3onltFuLxBvq7knEETCwVM7hEXFFE9jdrt8LsG1
9xFkE5FQDX0kkF1o5Er5S+dtijJ1mgTTo0b2tWh480gB+ol6XH0+fma34E0clgK7
9fTiFoDDlF/J1t/0VaJDGDr/YS5ax9bLAP+PK3Ewn7FPWeVe/GWiG0wPLf73igim
U8dPTyH0hH8Xn6FeFlWFd99cuPPekxPdjk2hnERZt2y+3aE1oF0dVQUMMwbgqIJ0
XEFaK8gbVEPAJ7uMQhWps1Fai5UVDg3DsZNATgEE72Z+5gBlltgr+mc3qOiDijqp
lPlYWMet8bqqPy+tKfQ+Mz/u+smV9CZxnQ55oE4v2PfCMCri2kiiV0etE1kLpmt3
3QlDKbb42mA4svX5sp0dOR771brxe8s067befN4W222dA3tDtSYeQdw/Lr926EIn
+S4OCgofJVe+M+uQBZoANrRQkviuipHo26H85MilCapYOp+SGUcHfsnorZS+XUWo
/xq7I3sX9B1inMpnZaYaoZjKc9Yi8bDwbLHv9PzNBu+nSF9AuQtnKbGngfyrjooo
emaNYdvE6suA8qLOQDP5XpYuNs8MtxF1UWpVC/kaThOZmoydld0LpG41eckxZWi1
gJNaWaVQhvJoNHxtHGajs6tl8Lbrv6xGql1RWFphAmZARb3Eqdwc/NVRatlEauX1
nzn5Nd22pbPn5EdxOZbbKAHtwjgqhd2mPHwoyfoPOpJ8Hu9c6h89uc5OIoDEuftK
M6fHD03VTwyYft7mtfo/Gn8u1NFdY3h9/uuWoe6LJtiEJStGHDCP31n8HxYqSmej
cK8pYQGamVRfQrH6ZnNhgXZ/uG6DD8+EIWnXixfRB3pRj32RUJ8f86VPzGALmWTc
uByiDZV2fC2FZFg2eVkbaoxZ3FSIT8IvwQvtAd32Ws95qcx03wJW5JagQUUifkci
/4nXhU0G5HhiUqL1DQlepD/MzVJgGDgRDdn+j9vvVsaPKHAoYkDoGfrWrJc6ow3c
y3xkP5htQc7bs6YLZCLOjF8n2bjxPHRlEdsHYYq7cxg9ocBqyDmYYBrYL0G1qusZ
czrWr/boLFuOtrgtaT/Pk/PybzUSzCh6ys9d9V4YOGL4k9b8JCRsuB8RT0rJsSU2
nh9aUe28akr23MO/lTI94AkYgKRYl8TSWvcUTftBD+D9D0KvBXMvSoNC3JLNgNmA
THDoBwGnxSmWO30DMX9UumbRH03rJQ21LQjwACOouQq7sA3rQ/VF+YlLBTinmZ7C
rLrZk5bOUmEna7W/u8beN8KCquJj7adZf6Qw66VGhUtr0pqEm4F1qe4MRzzbzbk5
HHm63Y0juYBcBkDd1JaNVrHWlRL4kJLhb2QmUNBm/nw3VcP/sbJEq226bHZwJQF2
CklAHxVRKWodIPOEb5j5uZfFhqxex8CgGVjc/jXdqWa4uKPmbcnKplheOOVDbFOf
UeaxyRvAKZH4GPj1HBBDbmOycuFojMuuelVD9FaPS+dAPzTvNMUk/Dvxq+gsnse1
CrR+evxfXL3TDeq+x2m4ODxyP6hUW/s2oW7bUYCNKB43b8ej619CIcRk/TPnjvMt
9ELB5dkTmGmwFNIJa/LpkTeOgls2Xckfxh5H5MlB93Xc30yfHzQiyFjX3L/tWpT8
o/8aW4KB8xNxJ31rTg2vbQBHRurxOXyF+5aOqTPb6yQ/1xtf985jN+h/lJWMYhCH
sFhdghIKv8B0pd0F2VPrOeajfwu0KpUoAs6lwV4dZOxy/bh4/B+ArAw/DI/zQ2qk
e0Y/w9HjbNpyJB88c34fMQL5K19Uc1+aj4gdZwfwzqRbCfFqK7Pa+bU35rpQmrGb
M98M4SIqi0TCFuiE2l0Z4IjIv5mKPkKgEgRKUEGniPAKu3wbAzjDrnLe95chngTk
mJT+EDPNY240L4viWhgrQqceXgwE55JkrREw2uvbq7pt1BPfxvwPwZal7EA13gOt
vvIzarnq/kL1ECl4Zrj6mcImWDSTpuybt0EQ6vy/2LHM8EncyOhN3vB5uJmkhWqS
OQciGA9mlbf6EPVD9s4WEwOzVnEXDm/LzGvq9vvQVlDvnspH5/iVhG3Ln6sRkrh8
1nk0ngFoPoVP6x7LwIbppTNrReH3wLQ8tm1Ts3PRRdx6kNhc0BY0gzRiMUR9Y4s7
E86B2rOUNifXSaOE5S63OsYJJAvsMm7Rz/WsKNiEN1up/CpUiCXm/GDkmylK1c2e
kVBSFsBhkRQQrKUd/8Ccmnh1Gqduyf46KjldQiFtLdBxETt3v/n6qSS9Wdqj5dwo
52qySBXh0eodsz81CV3lvjdgybeY/19VtcCQbyg0spOebuiAVMkXb2sPe7YMTfWa
vgqSLnsBPy608KVlGhtrnzpsx7Rgs7u64qgHLF5vguJ7EVsM7akU03XJ3zEqZ68v
StC51H2FeMc3yQgYXh8dUh76/WNUO9EriWDrREK9bv7QDwhLNC2wip3jOJIdJb2z
h2tZsmh8qW16F12TEb7E6qAmadyb6Pg5cg9EWMxcMWiA4A5T8AvOOZbE9OD41JFY
I6gThfl/0Y09O2no7fqNhB+qfDCtCgnqY/59AV3X98e4D7gVR9jKEmqAgJlLkGDM
dM7SBxFj56m9tRtAjpeb8Nk6g9BF8+wuTb+LKLoVDvtdaHpaE9pYRDXgFr4rVK/Y
mkk45Y5Z/e0k5lURtMXgLVlamysImDF6jo15EewfdPs7vk/G6jJMfYYTN2y1CP7e
i1H0VAYuGC6s2hDgum9HyhSmsFE4I1oTzssS14WhTKv3zXNlW2m6fmhA8QDX8hXh
8zVOkBMTSQiNVKyhjwHHosgqjYQ7IEouXzgWNVOhwAj+aqlnptaHbPq+HuqItmqf
IVtb6d0NUhuZGnjwagaip1tUCAeO6KTdHpV1fApgI8lhbNEU7LH3UsPwgFJRTSVu
bDVPffixi7oiyGmBtTIcID7N+jUHoVATV3FJna8jswZd78zr41/oD8D2HCze+/Ww
tA1teNXAtPGajeV/cUleqyqgvQ/AMusO/CP6EixFWCZJt+HeIjjZ5U08B08d8+pM
8VPSCjztw/3ItgcijovkeuIh5lmiODVImZvQaSAwtUi6dQInCEoh5wnOD3vc+2JR
QwJ680RFPFo7N5xVa8ayqasZrLzYvQ/DFyNwRgihasUToDEGZ7uN8yV12p+ei1xY
aFEu98TqGmfTe4rQewxBW5AVyr1F2inKix3UvnjMiJQd7Lu3qeE/cx+RsaI6DxnU
z8Be2mJzEZ2BcmsUGFrGQgssNKXEqduSPgoTN2x+qji2gWmrwYblHoGWHPsr7nt3
/fGvuvQVHmALi5/Kw7YmTfq//U2T4YIpCTZdTze/ocLYcV+H4wJPzBUR2D9oKi6Q
1aW0bN8ugWwhRQi8SgJTEe3kPbCUekVK/x+vcZ4XbDcFCvfjBqr/YCsAB22yJB/A
KWP46COz44QGORv7TFcMCSrvQTkAlGAdHHVGVeSk1NtOIKwDdToWXkEsNnNWI3Fl
Lx9t0SzJwYlLph7BNYzA14/bZIp9b5cL6tuIyryr7K6jJrk79K1cRkoCT2KG7Jha
rnlx1v07vwZLJNnQsUFr2diSrI+rqG6QNVFToH3icS2baqd1TqzL7d4FGkHVRnFu
Dm6sIxS9Dwft+2ym+JExVFVxlc8Sn8vkrqXufMvGyhD1ygZZBJLtGPbHNUBWTkWy
WMqmWEIJYWGHhTQRKHQntqOSLlgxTxgy4R6+6dFyyCLHA2A5M6PYFofs0vRfZrKB
fUXXnOWAanoCl0AzHmoJCCvwjlMPM/GjVjs/a2Lej/1WjkyyDDwG4nY4hPv04E0p
VkQkERX1RA2sAhWkZgGha3wX5PFFVV6fnqNiTMLvVwSQSCdPiGeBU0Ul1olOY0ap
v94G0VJXm+GPyXOoxHKbYkHmznCzQxy2jrYVjjJpOeJvF10Y2cJrbYDo1CQTwZtm
HOuXbC5GxWdDM83MDa83RgLFt/Z7rqgLoYMSG5Y6qIzFOCETOIv5THa0dmLAxO7U
ayrERdYfoAtrDjGs0f70gdFO27QHJREo+i0Dxr1wZiD/YBWaDt46C7snwYUw2vBU
pqpikPooZzcGnTkFSIk6XNkZf9Vek/3enIt0f3GjdLmr3CA0mKeGGYhbLkwxtwJK
L7D00PfjfRX+9rdgi1VlxnO/5fzVSMO80iEPN+DTUgtKKqo1jJQaEGqUOdFVfmJE
Z+mUAVdhiPVb77M6ZVRzB6FtA7Ye5Bm3ei0Azcrj/ABJGLa7NbIrZHC+4xja16rl
k8lzOasNN4MJmzpwW1qbY3jXT20MyemEVF+gzbSbpn9/PsUpUkWY6fD/S903tfEe
EmJdjMukvDC8Od9poUOIcFAgTg5ACz//ulu4X9eAQACNZyVqTqFdlV/nV54kqcOW
tg7bzAQnrV4JydQ97Xk3Yfl/ZnwBXAFdQVpg+cy4ZMKb9VvgN/cIck4xn3r690LD
Gx4c6W6QUslWzKJztmXYrAQk9wxk7cHcnrgaHtyAms4z+rWEgVOGm5uLrtQBBHUY
Qh16IEabUGI4NPLbIiEuCDhQ+pjYgPGOlZxNOZmeYAuyQPFK/EZxYzgi4EYfuVcU
iYU/dIyispVVfNmPIC5NwxwIAUCY20hSZJLvOZ//4oc+TNzmVVSWDJkIb/ANBFUX
HyBKHFcpvxYFhP6oy2pQmMepngr1QCxmndBF9CbbuIk2VwbVrfgOoJKX85Py6PYM
9+EuEmWMoqjaC7f+WurtdZ0To/nhpjCX9e58TCU1+qfMa3jjsxXyIkk0MYmPejo/
O7C0kkVCOdY+pvhqFsj9hfGMGIYNsD7r9D9vRkN8DQ5HYZScxRlnzMgvTmp92TZE
kynss8eMo1sTYhRYrZEqih8QJY3hY3ZPsrdqAcwfvudEJPpnov+c02gW1KfYmAAd
S09Wqq4QqDwE0cYNqrswcgQo5/8KcQipm7K4K9mhjqKd7EJ7HCUk6tFBK6RC+jNn
KO1ZwsobFTIVg6BotYRwxb0Tlxmt1X+D580yM1wAxi/nWf0nH9b3Nq6kry6gH1dC
C97kWLF2SREoo62OcY+CXGPrp8QIjAiOfh/RU2YG2xYNeCfe2zeDKZxxHCpPH58b
dMBfyZFSaLWHvIkJ8G64EXB/XKBXUGAvyZ7IUl0YINyHiNfUEoYUu+FlXUh3yk3b
LyXebETQMkIfVLXU8KtSGNRgDfZMrIE9+11jbdf9EklVWRI2q/0C7FOu1ZuR6pLH
8oCqGNcUdXMfXjinwiMCZjN4C+0oRq7wWiehSa+4Vn91khEaboKB2g7REa1fGYTy
Bm8m/GYotfytFZZcMpP7/oY5ZbGOoSRrOMsq5TBJYeTQTyvMXid/iFK1RFabxjkd
2Y04UwRInyK9OoJZG0Ra/m2SXYISzuh+MQDTruUt4wqGlPqiY0SKuqPsnLKxDOGS
vGAVCufDJm3qMp591Pjw2q3s7q/Ib2sQ3sNb8Y/z9EpRzwVyxIJ7hWZNzIlkI1Tz
GiiUW/lzb0iSA4UvaIVWO229cdj7+roZTdWm04h5EuJHStGZutfrT39FM2Zw5Eme
L2FtJrKv05NcFJMgVPRdSS50u/qGZcJL3L6F+G3gUNV4QXVvNsd/PoBUvcta7ee/
+9HL62y0q7gjXbUjzWrIosTXCo+LMea/PMaHrrFwFs8D2hZd8WkHEh7UGUg/XkJt
n1eQrjlVdMOsO/x4MrAHKA06o6LV0ngF2HVRAd5p4Td2yhckTheQAcl43rcPPVnk
LZgB3dDrxR/Pyz9RxQCW3MDmvGSi7Xvp7y3pSKU5EFktg+tFf1v3RoyASsoFNtZZ
GIE9Y/yQzZCOdT5AgxrXGriXy2CyMYJjot/2rFqJmryAnMQ+/gGwlQQs5jflk/UL
NSDnrabxumduAiCePIY1+b20GwXR5QSg2TubSLMMJ7tmm3Cui3GtElaJlBclmWWU
78h8ofqS19ob23cRdvFTIY15MJoxEuVHL+W8pdrlcwB4Xp6xyo/iIb4giUvqb/wz
e6zmSlGg02M5rpQxvOWp15mdaHLC3tX96N9AWJ4E9JcP9sHdqgXf68m3MW2gxuig
P5AK/uUyToBPGl94vq9s305qYLz+wZQe72uJmehjHlfii/SV6DxUbdSwyPBJuzRg
/FhISTOjeiwAqEJVaVU4nsaFNgt/N0xX7K7XXj0moy2W8eOPQli3GyzNdExKYu0b
ZZvIYx7Vy9e6DshT+Zh9HoY3akLY+bgOuakYqrePH9mcnCTbrLii3DL/BRW8KyBY
Tukqc6FJ/+7dHpqhfuo3iPOLMnRKHHkmdohkgQlAAzDpm3Z8Z+3o2KYclcsaNo7G
0LNTxepyttAYu/bsNu4PtWtCP6XBU4uCqR6IuI7rDGxX6AIvAJgzLjJUwihCv0Eu
WzJ54SRgnFW8Eq4C/ItEOnjdd0IDCX0OBZ49gibxA1HPM53JVqE3PL3MyQmIpVdv
3jFru94F63EI3WlEr/b/ZDU/qWyBDR0QZKPar9uqg+L7TkSyI44q/xPWB7xNOTBL
xXjkhcRfzVpMbJUMdfr7dB7WdPQvTG4nbiXVFPBc5CVFxfRFxrUB2S9WlDvfq6WA
kGZbC7J0L4MH9M4DCohSO6jU9pH1VxglEBpyx2vylEqfGzzkjcoEyyuVLUCkQv3V
5ilIqY/GVN/bVECoeZJugbStQAFePLXz7WOnO4uR9PEiOj1mwl778C7JgNBVbdfS
ah7OcZtjUNWCl3NxmHNTt3C+w3/Ovrmt7qndC3r53oPT51H3o6jC/xbPp76EWD5C
Z/Lrfiy1NgdS8aLIsSOEye42lzRi5UBE4HIH6b9crwQl6/4SwX7Ve5pegCP9/KuJ
r5cc5PyRsExEuZL40Q1jH5EyRjiTe2OMfLwGugMzVhKRu9schXW+xunTvLP2w+Al
4LNPHNPOddwcxZIMACDsAqXK3DEG00uT/FeZx7ZAVYzQ1uqRCMvw/lfbHRPMHWZD
3CvevhC6tvXFu7Ur3XiSPM3CgEsoaKDSacffTtD+b5XzX35vqhoJ9IYtO6Yg79Y7
rTucYnwzEzxc0bye2qo2KRErVM5GAhhdRsmpivh+KoznpyjSvRcxLSSV20EUvBW8
SXd6ldCwZ0mXSIccs1CTpAllmG0yricT2A3hcUmvIic82k7KyE6rnozTtzAEGD9Y
YiZy+8dhz7lW61juNVAaSnfxZu5qikMu40pRBfZjAsPUkeoLaqHyRATvD5gMEjcY
IwSWNu4pLZwlo+fmNsHA6bMaCPC+NwrGUgaNljdxZetr1VzG82GbZL13A/IpYAid
K6eoPP/6RzqGsjOkxLZW6KDqL84KKbhOJ7XzQB4KGinsK7VIRIZLyyXlw/FpJLp7
G8R5gLSaIw+Hdv8qb54LIMeqn8JRyZu4DwxzdOSPWSNrV0019rk6QyVxynO1qZ5c
CXL7NeE/QBohwY+DUjVmPUeocuLiA875yQwXAI2DGHNJDWV07UHBEKQ/0709ikn+
TZxU+QkzbZ7vSHb1k/XFnJUBp7ThdekYYmM+uhm0bK0/yL3y7s3oriDM0ZmqYiP8
MVpfIzuKoASO0ax5S2S1eqtA7FCNwUtJgkav7Li52JrnDvOeJ1mqZWKXF91A43im
RfbjKVTiK0Im/KPldw9MDChwvxvhUZrMnswkh3pbPCjLZVU5WDAeXg8K/0ZwuHK5
lCA8fjeQstxi3M1zIillHw72LdCJz1jAuRJKexgN7RvpymnWwt5rpcJ56DCZohjz
mUOn01NPred1CE3VWrJg2MJEm1og4PEMsSo4VINhBPnftpKX2memy9JMtovZ2UIM
2USkPp3E2s7XzxBIPTKP4s1jS5AH97KyqBcnnq8Qh0+0SLxox9VS+FS3qOAlcvOm
H1GXqzqyTtM5w78FwZofFP9Q8qsxZ2B3DIgVkWH6VgH5naRKj0Unc23hwA22XuVq
TkWjZeIg6YCZVCiMd++6zhfS7SihdJ6k0Gzh1wpasLzOezRg6zhgxT0vWp5qLl49
G9YeYtvyE37iUsx+ZgxjPTOTaOAk1Lkjzyy4iuwZrz0GTklFnUacq/rtc2gBrYjW
JivDNPcL4kevb3d+GafDTX1a58FbTD6TrPdi0YgDQ/3+UXZ8Ed0JPOPCRe+s/czE
9ZZ0jPcwAe9FwlnZt+tSAGexR7+x93kiwj4dHNxaF+9yNJM/dSQkiKIx6TV5E6ID
E42GYhkey61goTmb8VBwSgem9+TFRU1TlJkz3bBpkyBxhjdV2nTINqTTkX4EVj2d
Jd1Vw7/mAWbxAkZkYSOhOMpbJnk2+K5V9SmRrBjsuQ3ENT0nW2plyW5MLcGRpUYd
vk3ZZqzDFyP8XRfgqMh4rttusAEwYhEDIOGNaD+pXRbqLcqJQHIdvrb+nlqhJ8xT
eydVcVldGZ5p3rBn9XxntlPMfuMBLfcqUclIxmCIffwVnq823wo1RNlq3EHKMufD
15HQ7DcUsdDxtCU9LilUe1/igtSFcBd0DmbCXoUKDrTMHyPg4Ay+HIpwVw/ASrjf
o5Lq5kDBU+gV6BpABF97k8Ibf1s0p05UvUfYSUij/UGw2EvyRZWGHEOkcHv1bXSU
ivXzzri9xQM4pt3QJ9Vn8W+X6unmHEo0u27NgNMOV2WSKa36z1pr1rVWI0kQNwH6
77r3vmGViDnbnbvNZotBsOTrz/hFEn4d4WPYUDlW1nY3eOUCiqul4C/U3DSOIQN0
BDsMbD326BNK7OrS1B4EgOy1dG1MyXlCAaxI09Y6/auG/fMDXINQ+WPBxFJZpk+D
dCx2lfRrk3CYD74jhrWo7jGzlDmfQzmwEkWiknWcBcM44bb0uo4MWXZcAG7dUUlo
KUAMfSQy/k3zC0oP2+xqc6RVaNxEwuuvcubIzL8IkzHGuMvxQRwJ6Y8n7x+RWtIL
xmzxn0SkCQdXhKn38LcecsQoPxpEo99dear8vsUZ1RRQjS8ibanNXe9RQcOXox8D
hs5El5BIfo8egOoYYI42LcqqTwAAcqGWb/yRoNfnZ6lDHhWH3Csew0ab3HMFtsE3
67cE+mUeWZVrEfZ+NonJOix6l9zQSPWNgkRLiEsHXa3qsGPtnKkXSykTkC7NxSD3
EkQgUD/cMItUq59wD2vVqn6br9St5OBRknrrI52zvLnXjlDfoqdbWdsbc+u4Zk7J
bpr6jfwO7/RqlcMKZ2Z10yksnBR3IbzHyRY0srC6BIIM1/D+FBs0NS9TCXrq0sUE
3aZ+3A90coUJpv3RxxgZwREnsqUEnrBdAxx7cFb6tkKtZ23iNGpO9lOJrrvy/DI1
z1M0A4q+u+ylBRbhF6HxkdtqFDXbqrAtYBnaGEXjbhgbc9+rybq81HbrO+g2jo/m
ORfd/LlKXeXdLsKfrs3TozOF8Jljt3m5E4Jc4tKmPZaOV1DNI4PYyhsCR/R3wDfr
AfiU5TISBGdSp/WaqZh+AqzKukJ9N4iDlpehtmm6uXixxvrXOviT2/RzGjqO0gKe
gCK/+PurmWBUOkKRFPchZvVsgKLdFPJWCZpLDuKfNNWC/cUAdHlzuuXEDuiZVASS
Wb61afEQcUXA3I34viM1iWMrRMJOjj/HC94MKemkDEMRk6DPV/lmuTdgtpUkZsoy
r7zzcBAu4P8VU0fSDxU+j8D+5G6P2u30SUGjHvvm0njDOoSEifSPYY52sayowYmk
wjov0P6npYeUw+2VAzJ4U2AGbBM+mKyCv68AR30caPl5Eppp48Hk5bTJWDX3/+m4
52cp3mFiu9CIABM+qLFDltYSBNlQebsV0VRWQlwtqzv0LnA9pmEbnnFl9/tOvgTo
sVAtzxBhVKQdyxbqSdGwMG24vnXHTykJTta5RkndjGGqTGx72RwdvcMZ+4LZApVM
NZRh+GHUflIz5XUSe+BUfMI4usP+gP5/zNFlgYD9h3HQ8/j93rCHRKeyPbG3is0C
8fwMtrJGxvwOE9m904wdxrNeVdbLlc8P/R9kc8RFMQzu/KjYeuwAIWLh9SWqiRxL
b8jcgcEA7b5Wpz8rw1XhJxg/grB0580VPssVEf9SC5iFql2aFIsO+Cez81LOgvLv
JlMguXBmihqyDA63hy89yAqI8/asUZ1T29Jsk0un4bJQh08b8U1ax3OLRBuPT++W
ydl+yk6ZhMm3BcHbfVgyZhyPr4l/N+TrVxNwksWdmD2pVo7CCff17xm7760ENgzX
c/21gRCzCM3J3L4bRr50fdEZs7lCF4IvrLDH1bnc0KRMd+Q292NFiuS5h9GO5t1L
JF+kZID90AoVwphCj1lPSjtm32AROlak0+CL+4q3qyY8gQMq+VZ7roismkR6+pYl
Slsvgf5pF7OWyKu38k8VNOcjhA3yfxmeuzKtcpIzGSpEwN8W85HE0rpG/yGDZl7F
nwa/RVAyliLDRBpScUOsXi6Ok+jr9uPzcBZZY4fgK/OMyi3OpCdHnRZjOFx3NyDy
37KvfZGBheiN+XoTN4pe/ziUzLKUMR6sM/W7Hit/g9+u6fJo4RUHU8tBv9ZguIOM
3GDR5KJbPQG9HwwSCeOS69mL0FdWer6S8j77Xhiq/7MGo3l0Dc3RyCK0GtqpJYpr
MOPivNiOmopMgMPfpzPHpi7sfo+HX0VYZfggBlICnyD7Kz9QHJdATBlks88etqVo
PNpDdNcKQJvAPn4Q7kwNGWacTl7znTW00L0zbypz6rYuKcm7go6vp+wuUjVhvWN5
pcfuY5YrX+G25HwUiuDyWmGOKSpePx0SEWUWaasNKRsXLxAkAigQecZl4ieoPQOq
3F09QGFZ2RqBtw2Daf/eqemjQ1ScWFLXEP83Ygzu0b0mgW/x7d1Vt8jskMsr+8AQ
W1hGd03P6xUcXSUoo/hLsMeXmSk1y1DJfmoNuEQIU44HRGZPYgJjzZd20BWTAnzT
a/fuF/T7QyDOo11tKklLWTYoMJc5LKqkM6ov4w0+kPqChM44mr7IpcN1j54ifjWi
nrUUwkg8YTKxygfMLCKo6AmjLXu2PujRcrOG5lWIObdeDFSGxfG0zId9Q70fyObE
29f2pBdxlQekZR4+41uS060IiMAenKpf6Jms/gYXwvPMsvs9rl65W1M6xOFZOoIm
beZr4ucyNqXv9wrIQ6vrBN6saFPRju+xxqG1zoc5XwMI1Rja+pac2XZOW1N1Ggjm
uDG0FVJEWDmoM0N7NBDNkKei5WqZFgRtn1cCDbF1874qZknY8pY4YeJvMrLK0WO3
p5PQTw7TTnahLpy4QpXHxPfyhkmTnNmQS7lrcz6uY5D71pwqalTidKlNQaCG6EA7
ePA5pwxmmwQ1sidnkrt1NPIYOvQ38wD5cNpRx5B3aRg7iglkPrZ7VvUcP7VolbgI
iXKcdq0WPyGk8plHf7HPan7/QvVvoZc8LQrnON41Si2+hBakqt2X78Dh5Clat2rS
rRCuayGOldZqMTo3BRdoZSqeXBYNv1HAUd9bSYCwhKjLWSwc0d1mtjCqyz2vyjGv
C7by0w2gFhJhAVE7qy19G5pDm55iXPsA/7zATZ/kpMO5HKgSA7OWjvB99lvFzzPU
f0egVwsx+OfpnYFObIhrNiq2T00ggv0G0D4zOa7fuotmmQYFElIXAqlL6ba+0Vrx
fZl6SY3rjDAbAjjwmL16neT347D9PlPyNe/C3l0qtBa46fHKW6V9KB1SddjVZ/Fz
aF6mZcn8UcgYJKyLhi17rAL2nwlOz1/9EQ7R1OGX3CwUDU07xL9tl8IKUwfey4J/
zxm8FBfZQzHirDDn4d8ePSxSgHZgH+rAbgE5+KdY6/fNg/Omj+RHIEbO7DGn0NOk
2krvEVFxxVvjK7WjUZ80p7tD2ccthc2QoKPZg5oMKs0QgL6M/mfsKMLKN0As3Mh9
qNNmr/pycCn93KC2AxIHRWFjpZVyYkzSmJR/2zXnaylfBGJsZ+tq8V8Qmh9cU2tz
j6dWpoum9NgKgzl+5nHwKN/pTcq8QZJDAZ7+dMWS6VVkTsq6fgsTaYnQNWiyaM9N
6PFIa/IyMhuFURvpPwP30eyOrlY7qSI3n84lhSjS+mEkjV24L8K/Bsum8wbyeSTq
vef5K9YTKMnoNSltbwIEn8YtNcQ1r412fkl/FQS3IpIW2q5yIEXhAA9Tvzr8mnfm
evX/KeNMUB/qM9mH6w91yz3Zw6vGskP9UC3h/CQ/dE+Sze3/rmpEBel9rhQmqpIU
dPzGo8TkGAqmgasQesbcRwootIDbJHtXsDWNRNmKPBoT94lhOVUarpI4RPq6e6YH
XBTAeljas2jkuq35pEKbfbmnhvSGxL7WuriUAak8s1sypj7SBZeFIZQVkhwpSa1k
78Zo3tJvRmbRFngKCmLjEK4T3e5o6Gjn5yZveElczYDBP+YJLV6bhpn8xxxqT/i1
GHWCgJ8L6MQx2Wy6BFWWzEEstMs59FNBfVl+B6jEh34RDThI4Y4apwI8DrlFgkpE
wp3cp+oxxUsW8dmT9nBdLequRyLMvxSD5JUxjAA35D+T6HgnThYFWmXmtY3zWDTc
Mi1FUYyFRqUBXS4B5GkJFqPDAyNT4u8v2bAZuW9yx2T5/3dj/kQdXbGdK8usVKgO
8TsTPAFxsrHBs0VMgyu+mtqm/9egKQU+aI/uKIY9rvUMpyQRXbQ1nHaLeQZ+SJ9o
u6KVv6JfEKaYLuYJYWlQR5GGAp0X9vdzVUEA+w5Fxnbjd8QP3saBaNICYqHmcMrH
uYkso5aPgHD2GA/bDiqm4VcWE4V7WV+Bda+2VLLPZ0kgDxhLLXZG+zIeKpNosY1q
5sTiIm3O9kxqNTy4zHT5MywntMcckLYXSx3GpQIyQN7nIUPlu/7lnJYIASCsfXEe
LcdCYGPrwJdx7VT5EgXXctvZ7FGRU8uJDy6F1Qkz8NyV5eA/ccA71ERUV/R20vjx
H65SdlkuCUCqNG6Zc6w+oNdF30Gk2169DfNQeZqHBcBAIhQb0teUQEz49KpwGftt
w6DsuMWr+cFx0FQLMq0qns9jap4FBINOIYvKzzYgKqpm8kp+HL+wJ0aGHdmORIj8
c+yZ+sZtSM0oVu3CWuaxwBFP+lly1t2wpkVsSMorbctQolIX6TBovDE7r423C5mO
Zwwh9a0jpOW8nr1TEc56QtHN4gJBpy+aG0fGJBPOQ8JhhOiyMNHfnXDTjoS0Qzx/
7T4xPHDRvNxVoVkEjlTCn3PPuv7z+TjKAYCp/3RgdvVYZZaGNiOEHpTSMOP84jdf
bOMBzuZC2XKrFRPKeuBsX/b289hTlmx1hcVFLhXgJincY6QWedKbh2yPTnP81PDt
DNzBvX51R7ol+3lAv/80IauuDAVlH+NAKsqxVCuHt65JXLnM+mSpeeAWotUvKrhU
9NtfH/DHEHWeoq5ORCdMLqPldKZ8r4P7KDCGgTlxz71EAf137HIVWzQmKYTYHESm
5vWK0bVSlykp1leOoql35+wZU26UIWB+kFDHV4b4LOGcCbpPe8I2ICzR7vXLg9tV
w7pXXHd2Pon5berHyeSokWCUW+SdtVz3W9fmmQEHx5L5brNUAR2zZEczxEHv4yHR
R/SCuEXeTGI6WoJbjaW3uvHZnRvJpdoyk517MPJ8Mmjh8Z3uI9oaKFCrS9WugE27
1e9EKaDeyIvzbaxE4Ihmpq7PMdkvA8ovePXlnyp6vyn/2rGI2eCwnz2h490myc8M
OxYBMUkEUuO+qTuUVrroq6K0LHYD+JGqo/0GqMLVb5D04cIm3z3n8eGwQ9KK5o7a
uV67pKWRZnN1LNDb+CTfOnmJSX51dDpOFnGqN2HSGkxgtrysXpW9hsFc2BxUHLon
+xHbIvieYm+edf2UmtcivbzWjB+UDE0y10l/xk8CANxDePiUwvUzw96riea43ZN6
AnzXW+7e3Y3lwFMA10+sDMucfNo93PrvvaVUb5gnoAxMQ+/ilzWwxo4FTQkHzGMT
VFGN+2dj1vIjDnB1uMoA9oc91SpU65VPLI0c8Ha2TwR7Fx0gDaC4hD1wBbD8XtSx
oMb/JjoIEhCY4qtMyOSLihNckOEX2hci2aMBahGd+u8PqqGOe0wQfA14ajqSqIIa
SatbcNk3D9Ldk9ehOA6Hd7gHXttZlqgNJk4OWFkvfC5ey8W3YKhd8J+68klEHL2K
0AcW90alwee6t6agA44TmVAWlboHs4B1inqxphcetsmMvqw6oNzZEQX/bXPk6Mr8
tsHC39yuKJlpT7iFRw6KYw+anOwT6uCnZJdYKOBDWgNv8S9IjXLGe45Xx7VjShdD
tOTrRkz42tC2Ef8qVupeYXhE57gx/1m+qAMv+X0g4TtyIoqMKJ1v4RcBWaz6oz1H
hlXoD3+sY9mFo32mD441lGkkCswjurTj+dCQmkWiokOr/oQLNb0UQ4bXjxZ4OszZ
Go67+qN4gc8gMGPwLJ69Tg4S5CqlW06PjuRczW7fqjmii2OQdziDJ8glnWc+kqeP
9Ehp43rIK8f49YHb9+AWUhUpfhHyG5ztEpngfO1NetlpOsRvw//2E1VtlMD4f4zG
hdEoXmGqSl5p9xK7yA+l2TaQmeN+/X51cH+ggu8pTKGM73j748114FkPf6C071tq
BTs/TLkrRSqT2HFTa241eAp5Cv8B1FE4oXfbDmw5ppoOFcl9WNOVKO/bClIN8+Vr
5Vg2QB88Q9ZzjbCzhHI/dZwnaGwkOHYpyuzA812ZewMuLxCWGYDOXYjBQhf2vd5I
gSsqL9PQus0ZvrH1Ub1fGpzo1/AW2gVDmScHn9Jk+STZfPWbCIJ6wSFoTsTYONc+
zNHIpJIvVVu+mPr11xLAgwjIONx/yYbazw0MvlnTydaPRhSxke05y24bcLYtLVNd
J458bECo0NQAqeV4uh+u0Ow9e65TUXTVUpvuLaXKz6N6mjE6iuPSHb7ilROaAzHP
IQJOlqKHiZSPeMchSiy02nKfb6xuueDyWC2uLgIqU0GhUcItUCPcK73DHQ4BCkjv
UekXsZ9NcFRRTx6T90THmrJYjQLC/akfLWQsAiruMd5dMGg2T+LVqx4+hpoJ/aSG
Ig9sw6+xGl3aOPYlao0s3YtwIMB8PQE6SQdRvbezAkxBB1fRJZTX0U0Oi5l/1+Js
5xkEnyOjhZq9iBtNp912kaA+8uQ4fuZpK6xTgPnCREhTy1spq6969beXIDFwxm30
EIYE5agWAIPWZpeAdvzaD9BvOi2G0wI157WJ0mHh/mSdjuy4hHg8gTgKEWjtvhhS
6ZasbfBcab2brdD+vgbd8bQp2OuoS9SnFpZ2ZbiWq/NEW0UrYhFMEw8Qe8ZJAs4P
3luJCTeTWyCWOojr7JFb5AlvMAvcfV8asK5o4fZRN4fgXa7CbhA+zF0zCzjgOgIS
wfA5GA08HZegGttcBVY2/MbCMFTa1AWwLGsOB9JGa7MT0vv4WQEcM7GUeo4Am207
zhWgH+uk2WkYxnbPwCMx8rZzz8GFeMGLDrEiz4F9qSJ08F5VOW9pDKAwl/T2V/MR
h99P1cMiPtX0GGh1NzD+LBhyPqUgEY/jTxCwl2joXGgSFmJnZau2bsjRJcjmXWqz
GOSyj9c5hmde/qk9IxfdVSbYpU2s5uVs+eCWa/NTOb6ddyGGiWrsjdr1LqaDXEBQ
uuJIi7oczZwsCZ3TbzeAMdHSV+qneQav9X9UqhQB+VvmwlfWA4NQGAvFTNK7iiA5
p0BdnzbjNtCiTqtA9Sf3K9LFnrLT2LycPZIKecmonUJ6HuI+JozfNdXboXMhpm07
JdFFAiAKwQ2sR++LaWpZvRfZCm8Fb6+vc2ZFxsGJpsCBLBosC3zelxkEOkZOT+E1
sh5bZK97+z0X12hp6NeM2QHya9zJTB9svfdZ4MdNTV4/DkVDj13LV1CKXZvw0BkR
/eLRhbGF4ESslyJ7xlUDYMOwc3mOBtS6jCHOSxZJ5UHVieo0nFshVXSJDiNv4gt/
vZiKmNt5V9QSv/cVhBm8Ky5YmTHChxBzhPka1P3HrnIdR+nWXAxwis6yOYPi7bUB
dD3DpvD0OX+XUK0rCiSa3ECkpUMxyFQJEIS5KpB47ePkEpKF75NKkxJcBulsXuEO
Q1V6f8/dyJZ4DZ7RWekKwBKe57STxF7tP4IGoCrxoRB8tcrqLNn1C35NMFtLhW99
xvgLseKpVR/lqlL7eeV77L0JmXnfKb2ULGFu2GKv3/O9T6mjeTuVOk5gU3ZTmlOv
oGX09t2npJv4dPeu6gq8eD28PKVB9006Wi1O+BN5abWyHoedB9QLRzHpn2O60xzt
T0KISNt/CeV3e0Bk/jB0lWxsgtSt+/x44yvC2bLNWQ8/NenzaFx7eRbA6IZ4et58
aA9j6OpznnpfdCf6WmJRGTZztACWCi5x+jEkv1kLqPZ+RIhKHALwrsqI8+xC52m3
zADTdH4ZqVGrD5wdP+5Q++FemucYJPqShvlEItdzgKOteLJjhACVqMsQ6A96kjTf
cbXcyuw31MieFZf0thq4ppdm1W7sqx4ODiWat/mDe/1YAIcPjKqFc6eTywMy3dhX
EvHwHzqpVYcPVBc0Ml8jLtmxD08fAGJiSMWWSyqC+oZH427/SRKZOz5/bag9Kx1Q
G5NZycUji9YNUYqGukkd3qpUwHxruKd2G/Ms8TOC1otC0FiuI/aj3CvhoOk4syXU
67ZijBje8xRAsdo0oDzQoA4lihkooyMQq8NcZqghiNzW3HsKWMFjU8cSDzn9QYoQ
dDWfSf28er1kXelhuf+0QUS2V7ejVm6NVIzBCAcoj7B8g9cm9t6p5uzydwrN5W+B
ToHAvM9th6xLm94KmG91JjmBif9p2yMw+1yG3rk1M4aTnuB13BdGKp54tr7nvKEQ
h79Z4nfns9UCcts7Vk7li6pgT8RSZgL7NCMqBKO1uRxoZaQ4B4iYdJMZfwwj1t/y
PQbWUc6FdkwpN/Ry8AXzwWahohZ+CraYFKDYRBj5y1JzTyAmTDQ7NMKfBRL2ljgg
kE9+RwXYwUNH11MxZegtwIuLc5yxjuIE2O25J3wqEwRNzIB6U1kJ4PV/flxLJeXA
pJH+B0jGfxbZ9RScueIljYnPO9yrzQdDLORc3uUflQ85NE1wbQDa0GjKOUwraUo6
TW36E7sbQ/3Iqj389oU4U+d9fk5Rdqeptglf4sJyFhhKaoP9hJwakvW4q4q2ZF0f
ojhL6juplxo96HUGtn6llrdAR4X5WrwOCXwjENJeQEQ/Vfr2PpH+ao31vouUri8+
QY7JsZ1lwMIgq1ImpMur4LA6jqUFW6dv7oS9PfKBGq9SC8rnv23ELtWX/CEfdCCf
JnsXn4dgErXzMoDqscg6BoMnhLw8goQ4H1lE92I4oS+1p+gs/MYDvEpp7d9WgJAa
getSPg1/A+XXKWjg3zUIApMPgwHdH8kfPVsTdOJm2WSURlG0KcTN6v2L1JDBis47
SgwEU1l0z4MfaFN+fDuuz6l365VcssxohBZzaDbXZuUVefpSaYAmTlX7rdd69vj9
yKkBcnVrh7+KOwnszFovLpJq9ZxI+y5kh3EvqF6w/7BBuWju6q4n8Y1UhM+hDMJe
iGXIOhj+E5Iu0erHGWqVmVzyEOzuE2AMVX3WIlhyy+HQPj35BfRcxc6HwJzyO3vD
K64WQvK9FnVm5YbvSY6ZDIC8YlM4JbONK2IkEE8vuonbbi65dN79IgxtvhkVJYQe
kqSuNMeR6y7lX6VqKV7ic0+/4YHZeFMGq2ziF36V5Lg54LK00MQdFS+1WpS75gfl
+Creqmelc25zSHfwVsCZ8dZxBX2tsjdSrWKSqao1p1lh4fZrgaAIIzF7QNRUVRME
PXMYQeL5Z9sdGE7dGIz0qJxasudDj9vA1w9jxe3Y3+rPUmRZdVrwgjqheRyhULng
ZCH3T/74mPKOCtg3u5DW9pCc/0IelF8wDaOCLtPpLRnWxyEG1F2/kIw5cPIvRycL
l7mfMuWfr36CbQq96IGOYJ84SVBdOWojMPPEWcBhHFnUwWuHS/wjbTKr6NcPzk6J
E2AYDICtBuOdhDdXntWNB+LTV/mRuggxEulg9H7PkAyhLGJRuF4/++neTOe01u7m
mhYSNiGlW7jlGAGflafkYYjgi1D92WjHHMR1lZtmlVZzBVRNLojll6lZC94KnO4/
215JhK3kIGALWIUbXUJtsOmFk70DXfd3Cuxx2Gpj49v8KHFVtKlgTlBUQLfZB0hM
08SWXwuAqmEf/4pYbFIaYvmgVnfIP+0eMdoYUeX0xnnMXBg31PPMd/HMChJ5ySr4
mNczoaJdrfSvrvgMZNiFP01gtDejpNmQGYlv4l3NyKl32fHxXC+DCeThFlKYy1Nh
Fjrnp7wmQ40JkObg7AYzRwc04JrZi/+nTBxu15/nqpkJ1hbVQi+7d6aVfYFTyx4Q
iY3iIYZTqCl5q6oCfy3T/yHXPZ1NGSKkQqHXyvb9zu6jZjkIyIz0wiPPA6DaSUeY
k+3m6EyFHwKuNyNapNdr0Pcp1bUOwJZu3gTnloFGLvwPRDMPXq+u5saa7Fq0iIXg
gttlNxxDCxdpkpnIz1i4hZE1mRn7UtHRq1n/RPIGTEUZutys3248x/RUuZ+wl9kc
3ll0iIYpkQG38mz51jqLHvbVGPzBVBCxgFG7xgIN7NqW4YmAycNUSa7l9esEWdN6
OoRKhYTRJ6gZU9ZHnOgIjOZSpck8qDMPACajdlvGlPyp73hY+/nsmOdbCURUF841
EuuBx7NNZ3LRdrbAv2OoOxefvAxStAtcEx4nPzi8Mc0ArmkDFn/C4ov/n2SpC9HF
k+dsTvkcXY3LmyH2uBnfLCdNExtY+YzhwBCE5n2YRwPJJmOUm+JtmwLpr+Q44cqD
AAm86r2Sjss5Adbc5zOGWErMxh9enZ4ARo+JSaTF8BOn8slputxB2DZzlpFmkqhW
xiN7Hdt5RCxMjoYzQz+HxqS7dKtXHn+Bvc8yRVEP2VxYiEZ1LTxLNxWoyvfAfsXh
4YwQ5pL31jsjOdRV6P6XuYmlIga1rr4O4Bf5fxLCbqfp7UPnsgOTMVkPy8kJXP7E
M8y8VgR7S+XgWFsg+poR7CTdhy+u4mgqa5wJYKOryJRXOH2u63Ey3ZuihEX8CaI5
2AyGcoeQ2LR7jl8uK6b62b4lIrhPHFY86fMrDZLGH+A/wEn8gOseR1iIVFGA/Zox
sIEp5rHGBkxk4rmHXFV02enTQIxOnepAQJYX7wazszehE4Kzjs6IQKV4JbZDNYK0
7zAXCdk/g9IVPHo3zqSq0cdG97Jn1w2A0RcIxgYtqwf3uclcpu1Gu/yg64dfLubL
7S4dQCQPLdbVyjjh2/FbF0EzK/bcozgOdiHxfI/1Z5LlSxIKvaCpfHXxjfZG2Auq
83E9CKU3LQZs5c+KrRQk6JBVKetiTzQ01wpK09WtvF0oPo9tV6hyb8G/M9VyF8u6
CPJSHw7FMY2aWzlAp8KOBAbT6+5JO15FvrDLKLqleKHEDPzsfJPSttsmo9SFfh/W
PBeGJSyTm1Q8nxF0bNJd0/kWmKVPMqzj3eiaVigwEs/ZvCaTIWxqtSU+nhdLf24Q
aSRPfyiZOqAIj2lpmAeeAUE2BUKSaJBV+JgPKkNMOpKIyJZPrK7jJ6M1gNWH1xLW
VaEFIba7a9xMM3ngxm3pqWZ29U5tKZBy8x/YXUPg9jF4R5omP1RiqdXMXAVuPqaS
079WR1J6k1tMhlVuSJ4ryoVi2WM5kySuY/6A8Lwd44RkpRgigWtCh9CqxudVzBjL
r/Ck3Ty8y0gEIqAdlD/n88vcDTM0QVGZQAS3Ms/wsQS/Gbu8YPc07GpQ1DFbskqU
0+znAKh1vZxcHmb7wzkaFRCBpvNZwCSY83P5rnWDOCgPypEqTgwJePNvHqd2hPxU
YMa/7Bh6LccSkdCX/lTZO4cAltV4svvOMYfD877oxhmbQ2GyyYc8RAKcux5rLwvJ
XQnCefgFGYucddUmDIth+ZmOlxyI3RL0S8rg+5lcQmpmNSuFUvGyfC7GLmfzuLPn
O0kgioSxOk4guCXy7csjwmHhLy9sAlkWXJSZMXBoVapl+aH1pHQOVL7025b2jBnu
oHcog5IpJdunsvvNRfaht85wx9/AwlWvDoBuKVNK3GiukQ2fJ66BH3XJEcUnK5gb
wrB6EWLCYGANiVRiOWWYo2jBWVQ2m8SFNC4jAldtBbQvmlnli3jIBIJCqNo7dXuo
cXWY7ImnzBquvsarvHq6WHehWwbm4TZGz903x73LPCTreZzlQ6PQ1urO8ZQBk4pq
oGndwLxPkg7cw4bzp4wc5z4X19cRjVJUjE4Mftp9eP6jjWSg6zOJaJ70/Zi00L6g
Rq6FwC1lYzmJkGU2h2YfgZQ5X4wGBPc9gU37SQAIgsYwViOnZYa0ghiPfVAcyRBs
HxyxlxZn8XPbLFiSUKrs7bLo9eBM9ryQkCeyWbbtUMK3W0YU6gkB2OclKKyCKobt
h+6G8u2u6c5eLU+ukNC5oLryi2QOGTtRV/kfP/7/og/lGoTMeSq0htwLDwW3K7Bp
8/V4BJNGFQvxAhe9gZ6W5UmeGKrpKGgK/urlgC/37cmfa9HLA7eEtNEAVvrt+UjP
WhMzMew5R3ASQV2c7KtqFMiMqzIpOpSLvpGty1n2TS/3hHg4Tn7g9V1u09uJlG0V
NyrU1qtF7bdRag1kNsXLxk3D7yzPnRG0XmILw6rZ9Umeb8q31+AmtHcUVSOd2Ruy
1SwS3UENODco+wuNKCn3ihwGy6Mq7CNzR39VXCiGtv7B1di7PZO6hUN0MJmUHTMP
mm/YVx1BEEVPbPGxpKZEqXLLc7fUNlXz2FU4OpFawi+czu500IU/EyrR9EubG8K8
H7HyLf86KJyCs5YV6/ignsfgpaOKvIqNLWimROCERj2eDx37xEP7g2oici/Z5ZlX
ZyKbW8aEKwDV6GvPlkEcd3gsIlxxHgni8vgeUYM4J+xHxBaeo7YDJ4NPe6xc+0v1
H/uV3skoBrmwl6MyciCURwnJ84VuPsY/9XbYW8dC4TtaZu0JQ+BD+93arJ7fg1HK
EO9uKebX2/EmZOGYEPUe5FKiUUVI+2jqd1jaPvpf/ZLBnsaYuB6H/dxOE2rtRLJJ
n0UdDx6WMFO++hEHm/98TpYDVaavsul5aEqD8YJsm0tnDLlFIU6BSgSRUAVw0r41
E4X6OAu+le4SxTQg99I++8qk1DHIu78FCYuwsPpZq6aO84FxbxV0QBrUvX/3Uic4
e1LvAl/eFRk///St9wjRKitJLG1nFjNVgSddyJytWMwF7bxrGLeU5UpDav6VFuX1
hSlzyQRRnGiAdwQRDsgSGI1wVQGuGzmPzk7vwm7yuk7PBD5h/MGKSuV3A6vKRZam
dPUiYT/YnX8hDwUzk+mPm6CHv8Jk+oHVf+NP0KBCPx61nwvnBtDvxgFswz7CliGE
k36ahLW3C11UyFqhjVOVFXm2UDPkoHv7Ze5mD63zFjA9kAGFEk15/MxVCKyNkZP+
YItnwxwL+asbUY40v1TT98Kx9ezCOBhYHBCeVVScjDpNOXqr/Bbr8O3PRJhzlILD
ojXF4LW+Zmk38al8jLpUoufVhXAC+uKuz3NIlefTAAxrlhsKyKuQcFBMBZ7vLmfs
ckzk920GB7iBfHjqG4wzahYlqk1hQeLyCJAGtQV7XnqI/A4MWIYoWX1X8r00D/xW
PbR1O/EDUEZUYZ8bugrARh46cBJLpD95z2pd9gZPUGN8UNlkySrQBRiZGROeoo2V
i/MpnVJFFsaJKnOs3zVRhv33DfVsgKYlB15BFnQcVCQ5n39qV8JnmkbRsfT12X18
8epKqk4dRLs9IGlJdkurQrykjPJjwx6j2hgOVRLnQUYjxCYHwJrTWbHQ4FEtLWhl
/MjzGLatWZndBMpXbLOUCjZf7KmOFPCgGizKdNgjhPpqfVFIWhtr10oFlLHcNU/p
NswDJdRX9Gq1M0/pwmZwUSaUgJ1Y0bvuJ1DZFJjBuTp0/hSnOOridzuF+fAYTwUr
/J8OrLiDcDOYTiD1ScxHl1LWYqTEdyQ8c0ZUxGb0lvtbPG2X64PF5VRtRYrYsZ4U
eguTorlMNGDfzn1gSdlLl+87gXeqgdb2da2pZMJoBNAMPD+DRljx3m/L+hu6Nusy
i1Tk0c8qXWwWzAywveVJ18/WJOaaTiETZXIyh8jSXgkiwUDZ5q5fdOZZFlwlUw/A
z0Gh6ASG/zCJTjNLzlnBLKRTuRtoVBs29Ja6aBbobZC2m54fW7PLT0NDumKiAOwZ
UNvswXmQjPRFAbqfH+vnU4GYWjuaV2CpGRiDY2z+stCRYRh2WnBFPSFjDqSj7Akg
2EJyuoslXYXdJJcNGPqlCoVHT5+pAglbjcNyuKQFx+aDmnGRqBg0gXpP/YP/jKmv
dYMYMioddnfqXtxJTXP/Lkfu7Ikdim+YGO+G6mD0lOTgdn58Y5TG9EqBFiuxOt4c
FKYhSZ6+TseATcHXlhTQbCt5kjLOCuTj4/pYsMKWWY8pVuzHVQ8BY03poNJMG4RK
UfsWz6Ex1wZoVR9r5BkRkXLM1EwbLI4HkLFOZCpaCawhEu57TZgUrqT9EgpTTQTb
Lm1lTxpXH7ucLt4+PkC2c6+9wwHNjKBzjmYgAhbcUQnpjdRAWm8vlZajLW8GjgZS
jsZUjD00lhjJB0P03juA3VbiZPs1l2QQ4XHUyl2dm4IS2rs7LAVB/hBPjYxi+5Xn
MieHyLXLFjoJiFtxPVrmIaYrVw6fHCzgvsTyvmMmMdhe457mjGEB+ocEztJZGy/E
20DOWad/34aLyCmIGXYxhnMlDxMAXF3G73HCSKZ0mapzC6JDaVwRQJZnGlw2WTw/
3JNoKox8pMBuufEfwRGSnc9jvHd9dGaXRHYWPHAN7GBx+L0YTaf1rRUUfLHLPFiD
wWr260mcNS0ZclhqdNtkydlbI5yyek+xv+XVvKeVjVxemyRQ4kUC5VjrwlVF7DaI
8jsibZNnlHHr18tCV5Ah8r0Bxq4kfUqmdq9uy+F4yN/net9xMGxBkN0BqhT263yV
XyD3BXszWeFHLSQKyzlGvm3D9gOVj4ljK/Eni0BE2SXGWjYliOuKmPGEdZrEgbZq
zUIHTQA/UdHnNtv0g1YsXZxXFpbdcxCOWaQeoA/G327cRvYEpnON+U8lyh0aNrDT
aQaMg56fVaaCggeXmpaHoGc4ObZJo4jBv93MonNAYtNBJIjSiOn+biKshQRMxroU
Zvx6ylAjUOixYXxVAKzEXAnkAeFvEhi1okliLg92x1d4dtAmoqqdL4sUpgFOOEoC
Pl/UD7zKsL/zJ5dR8pOyQu7D7Uhvc9LDHZLvQWPOOaQO4Y6KZ/4UPQUJE1/Md8JG
M0AX2AD8J7JuNWoJMbjr9eiEd8x3R+h0gJMLfG/cHNAsGFkUOcpP5VoSqUFEylrB
zJ5panyeJCtzjYwAtm4ZK09PEA/1tLYlM/kt6AozJcF4o5lMH8Aes1h0pFi8MIZN
ERdNtG/MK728EV8PyYaygwz5FfxDW0SLjM6IZZ6qUQXNS2UWCv99lSmIbX6Aj4p8
MqFMEFUnPxFyh9rNLqlQIg/VAe8RZdL2V5FrK1AlqIRFQxa0kC79Lb4Tv4WhUkIT
S+5IgvKqFRpggSgYjwLO4v9ZTS7VtSL1z9mDHQFWvrRPbG7shbCoIfKmeUtJ8YrB
TyZ8wWGBzdTUU5KmB58bZKuNc4XsdGN7NTFgkQCl9utgYVVPiIiT69q3ksIvMe0s
zOmZgxoZtVyTr6f4UJQjY81bI8Cvt1Lqzr9IuO+kS2c/5Iz/cb8Wv9brUewrz4O9
UQR0mmoDpxhAcxhW2julymtEktMMThuCI8GMP3zYMiNhtxw4GPDGaHqgL56eMqHd
VnNgqu+lajiYE1xNRmBpOKnibJKORLMvU/fUAFidtWz62jvV2b0ZickM8rAbb3cn
ka8iTrAQpm0afRx3YWZ1zGSB+bX0s+FBEUgZbJZ6kII6hXmZPIcgjzQeIP6JeCRd
fi8I0XpMNs/5UB8zNa1rcIZz64q6xyNI7YqjfSth/R0mQ64Lzkr8UYLcLJkwdQN6
MtCQUypBxntvWGQf/EWlF2rh4VXZtz6bTW2Br526n8E7nNrJJCptgWoMm5Yy1BYU
vCMRcOqPgzmyqWrsO/0nxYWRfo+XztfWou3gR76s33H9lFeFLRsY94sEaqyoVZEt
Opqh6Qpx5rxO6Z1f1wQjKWMuya95/gxijDWFCtkO+8t549m5POezQ5G7N/43VwwJ
KixagQ/QIlaiw4kmBB6Mbo5WelnCC3ms1WFbV6qNYpeVZ34r5KsNgF2n6HX8QNVP
M3LqYcjDeY6x0RcS+Ak9MmMUO+iaLX1ldiDmw2xEMweVuslSO3YR37jlTWtJx8uq
FhT28TW8SfhgT/PJ4uZQscWnY62g4ZaRt7gr8ahBvX8sAnxXUPzM4/nehyPTYAb7
JrpAEmkEex2bsv4cMeUZiHC6o6w8eEmp3lhLTwmJQAAr1fjH0B5GJh8QBXh//Xg5
k5fyq0gXQkRYpYBcMhNepGIRENw/Dun9WODpp0S824r/wDI+Vmi92qh6Y2ZtOcMZ
S6iuxK/jxxip8WcO1PE4E13PVOCayjkCaRZ95BjegJMrlfFsA1uTtzsqYdRTn7m9
qItAo0aXhW3y8PNcwU31ANPF10zuDlvz9EWtaHfKWtaDlXp5sI01BG8i2vpasWd5
mrAPgSWNCioWXYWQs1g7jOobXoP3A6yhz+d/n+z1pl8+/y69lsHqvdzBwvtxOO8M
vgcB+Z8r/r7Gvo1WDHrS0xs5C29xUcN78aWGsjDT92W9NfbegJyDCsz1d/hKCFP7
WCrMuponL2zNONPMhLkH5eTZOTBoYG94XLBxKPYUjRH5QfcXDpD42/G+VfCdubOI
WMj732irBQsxlO9bDdao4y5WHcPQ0uvDCqPoZDaUNsrvIHLUhOcPmL0+DEy/Y6my
+82IDGrq4An0mq9Qvq9YodoWwtx+mNKqn4BIwtIiZ809qGDI2m6FvyC2gEFUd2hi
JYqxddYT1Wd0ov3RMUZcWfy9b2KIy0bH94cJdueBefVTIcGpjqzOvH2vSiFW1/DW
pbZ883boe92u2bhcrtg7kvwCzh/9XQKxEV1TLpzW/2CfBLUvOvAkIDp4v3QdCY6B
Sk7mH5w1KFC0zTiIJ3Nr9NPbON91UTjoSx+SFk8CW0swBqIh54Cq662Zz7Adac75
2yvb4attQccziBMbuq+PAcle8pewtbCP5iV0BujG+zCSIr8CihQSAD2OGzOtuLTH
m/+m+hZctBrkHoql+qLPr3DqLTl2iM8N/srKVCcUkKHdWDSm5/GPy1AYhMPJXKfM
FMEzVS1227UT4yoxg37sk81Sqht3F8g5/AgJXM8LMzRa4X6zAhHGAQgTrNjkZzGZ
0Ta4lpCdaGyWjyIKEZWAt74l4hp9ir9oOn4ZDGnbR0VFqfoFlrS1MUTNdNvIBvg4
p5FsRw+70hSRX5ZZbFf9zcfTl1ojea3eDj6/fkXKXuzbWkE0wVsIswoEgNLtCLKa
/Zwc1H74iE9aB+gy5rMRjvTN0nMIg1mDpvK9Xn9cAEieBnvqFwknlJrJ3tK1I0CU
eWCTZBd1jXRJCuzonie9kjfzUloxi3ptT1ctrPyUQxrezEPDghXkXM/+wrywUG6g
fYwXzwYhxNORygmjjNTXUsQ5iNXwL7K/qw8r0keUpPCiVvQT5KleglSLZVQGHMLU
GnyaFWBlttHdR0RFRN5NAXPCwQzWZsR+PcGDhOY+4eHNppVXFS4LEhYRiH0RooWm
HZlYea2rV4EkO+5hxp1f8ISpbua8v9eFTsTAeRAG9DTcl1eUNL4ry2kaa5eZmPwN
1vwEqQhbbapJfz/OZXWd3vQP2LJjofOl0GcmnpdlXwRzvXJVeeRH2tbnqnVkUJKK
AALHr0ub2xJFjMDxS9iXXEdFvJjSvRBBMjvo/GYUSWNbc4CDFaSniIvJK5JcMcbH
g8QJ4Hg3nwDjQHrCt0bVo+uHV1ICPRuolD1Ol5KCe1BfMrfYRSxgLkGsrWNwxyKq
12/Vr/AW7agADo72HphMudl9dWkt57aL9Ssy5YI6OAT5MLwu/qNsSkdU6AGg9BPL
QEn+eaqPKbhfaa+XPKqWGWDBR5y0nWYEOBHr644G6Ezegur44eL6uKpZu6Re8UOU
oJ/VtNG6H0VXB4286ZKzJXThXLRcskRnlSk8sQu4T6Z24S3wCQ7IJIrsRIZjoIm/
573TY/7tK2kOyxAPKHfWu2JUhzZhO2OJru5g/e6ZoRUZ+w7u876Y7cRUDmt07XR9
LRjP3ncDnUDs3NMOkRFn5T74DfXrJaUoOUsNBj4bLGL+Vq08ar0OWHARd/i0a7Ii
CoBG9ZlM9QvKSNTPOPh0+9k5E04AGHMYXQzujZlUHZSjoU041rTgrFfVpf3GwSPd
nvuYSqUW0a9FBpHMBxnOh7aHTGk9NpOZYTToGkeJJVa0h15RYGwhJB+QNmlH12yy
tarhEGgmqelgp2Yl5x+nAo4sQ4i+1dadITTSJFnBExYjBC3jYCi3rzUmiaBDiZ/y
cFhVMOQK8U8XT4sfUCaPaL4GYZzwDd9pqS5rg+CRBkVB/gM6xcHi4cg6jjt6kpyQ
AJndfPSWjIbL+Vrp0eIaPLiXnCbQF1VbRE2eSP1Hl5tfGKm9RZZ7KykWDtJ4rmGy
Mm8mF5LwwVe0UZz2/092VrXXe8YBOMmvjLFdA3gSOZntZSpi0pl5LoJG7WfRWuRy
59Z4fn7/VmUCcm4KSGFUO0oOpsabud96tuVWDzUtYATy+bEqoFYiQmxWN5XzjXq7
vVGfYNvqBWmk9v8g68qNM5zx29BjOeuxgXswAczj9djhTRByUzmrHGuFHZJ7fsgd
mL+f/3sRMpMDYFtdKvUT0bjmfm+rrel0i7kh1BRG/zIJEOzu/KGg4HhkGlo3D25J
uW4QSi3uzLBSw0eHTRNlBViHa8ZAGYloilou79ySUiTpIPfHIxVWVVDdZYf1xBe2
QIrJbU2dHmQwylQtCYyWg6uWRuE/BjftTg21mh6huj9QrO3vEi4YpK3c1nMpAzaI
xex6wZ7noRSE0FDaMdWd1mX6Ndb4sPJ/ato6arklxMjhsO2kU3psDm+92da5thRN
j9cw3tYV7Iyp4rwf7QqQChpxtbstzwUJ2UtRv2uekzdF6QgllB/wWKhpNZKLFY34
i9L1c+fOMG/qdv14Nq276qGHnEQGzhvHzD5NHjZw5Bildcmowb4gh0FlKth4DaKt
8iFSr+AmmqAKgjdHvGIb6U3y3DfCzYrSgfEkk4swFNBzXNCPOqPfs9wIrGAIXDIl
OtMZDjQf3NaZ/DGVmkOMySrQYROwQDEqiP3aSyps5w5w6sq3R+DWu/GIwU77yqSl
g6EiQ9MUR0P2DEpC8GSPapUv+EE6PbvtlkjA+MpAL/AzIH/SLz0E0nPry42r+UUH
vwgIxCBn0/03xsXquSbahl3U5jHibkn5V5mLCoXsl/L/yii/Z15/2YyVTbvsgrt0
eOEnlkvZgvLibIBVa1fokyIoZh0O+c50h+licsgAi34KFnQfO+TCc7Y/mUgtQoF1
1VI+zFDSZg+Q8MWJJEf/IYZ/+hwoYo0gNotqX2c0buDDt86g/sHVD6tf2ZAdYfJj
J4u685BlxtqPte7mdnslXsYAzkG9nLMWN2ThkzOPS/cqgl92O/P3rAoOvAyMaXTm
emZ0eRBShB+hsX2pIwF7JLUxfkHBpm4JWPBKAmCF1/iRDxJKtdB7VPRMUueoRXsk
a6ovfoXM2O/qy+rssX/01k+D4ehJ3V+R5/9+r/WHWD18eeFtrSNuPbbpTBjMdTLM
2lNXG/pIlzCBPibH4ofEAjKNsWTMYwgd2E+DoH7uiPVodidUBdYYjyvNH7IX5jdD
FEKS2u+473PnwLScsBPsZxeCU8q/NL3w5ucH0ZYHGZXiC425EoHQhzanBmE+NaNU
x58y8LY1VgmeybpuZlriM8UwOZjtPQ2iC4k1HK5U6cwEkuzU1/JFxPBuYoPHsv7W
2qo8XQyAq0k2zEyMTnYgmOIDbpNvq6ykoPK+9EE+BpCBXPn/huQHFCT7r72qrSw9
hXFdfRKMexn5j6IYvhBGIR9cROEZ5uQ4JRl7/hMBE56AVpazw0K+sDLKDnGLnLbk
do+Qt/4kYBeUKGUqrmDSxMaBHts1UKqO1uQs7tV5I4+6vvknQLYUee5y6BmQ2sIi
rElHfvpk91jS42WQ0a0XbrsSE6h/ZDP+tGXO2DG59QnX8V1WfOI+0GICIedRyvan
gw+udjUkxih0tP+UvP/QBGOD5Zl/j6N1I5Q8QKoxIrarLtOB2jpPoHxZEFv/M468
MGQp5xnKtP1CL93eqWYYuaw3fYaLPFJiczieqKGYaCI2TrvZbF+uzsZ/gBXDe4yI
b+dkZCCufmekIankTvQP9jk2R7lABOrKOFXzC28VidQW609wTLtKCBllOUivdxfE
xf9v17CCkkMx64786U/Ugr2Jr2ho9eX5iY7Cc/CepCDqDhD0SH6UHZhBv1R6nrzR
gvcxhy5k6ixJt0UukBHZFxdyUcWjjlf8LSc6P+XN0NdTOnyWmMJtzXIMFtooAZm0
nqBfcTYAVW6FDRYk8anSIgR5t06Zny1fAL8swQcFAmnbXEDBjDRSs6yE2aNqonNV
8i+bnZn7BLXtv6eYMooqOTFqWWogEAl3SbXXjMhJw2IrNTQz5nCHTX3Srw+Rezuj
EtjQzNJsYba0z6IDZUqo5Zy0N3AFQwk5WRWiJjnPX3rjtKAKHXnFKCDE1E2Dm7Uj
uOEqMWiA8NhnR+nLTLhYzNM3ekfFxkHQkpthZw6egM9CJrpLjhiZRSYkzXIPR2uj
gEYuW3AUH46/GVwBbxOXXD8jEqE5HR+BhM4rvuViFlAnK6CVUaVVc4GTq8NSEqQL
VLmTGXTeEctFfZhdnu+xiecWyis7NLKjIDobxlOGMKBqoxWYTanZf6OeLK0CdJM6
n4V2QsXvaCuUc781WKv0C25X000t0sMJiTpUAOIrmjqE0+ACUS78KV4GMBR9UKbZ
g3TQ2BOoiitDjOt03qBFhrjJdLmGL+8D9bGCbsEjyOG9MtUV48YWgVvyUmqLBfAj
RSefJ8sHqrMEdHjgET83h8JwZQHUynwzJbniD83rJguelgy073CrXX7mdkMPHUwv
0uEgV18mSwtmrMNdCzvjVGbiW7I0t7fYJothV+7xXN84ktmMXVNH47vL46v1qU9T
9ufaRQXDG+RoqWJ7BCS17vPAh9ppfQISi+QzFDDxnd3dLFo9Fg2BS1CX2McSW2RZ
q3/PpV7RBNfgIgKzL4Ru7b0z+gBxYdlPbxV5DjRoJJDx7/+NpHW+Vq0rYEeSbtKd
ZLWk21hEyWqlRCBv6SUQNXBTAHI+blmCQS9ghakDC8aEIDG2wEPcybpeL7laePVr
5jLeZWDkDVRoN4cYwKruM0zWc64TUgIcE8NIY1vcaCuZHtl5C2bmjf+nXLIkUlHc
+CgnqCN1Ap90IfKksr73VGM+Hj85826l1FyhkPiyTthDuwW7l6y1L+i4cq3Hav7W
o83AU9fRxbaj2J0kVW5Bcv7BHizdtBhZu3cnaDjMlaQ16dGy54F40+h3MuqlVK0O
lL/VwBnRS9JSXVXsvAT3RPIoE9XGkJDtpYlHPCgZJ0WbKZvOEujgiSAgvyjo7nzL
f+K545vF9K4BJfXSYaL9LjeXbHE0oMk9eW3Ybr7T0+hZ59ge98uJ4Bm+wmFHGKjQ
QIQGCNQpwXt9SD9eEWF/KBLhIhq2fmQo8EMs4fR6ene9HUD1W0DULwE4tXqkk1+u
YR00epsr1hMrPwn1++vAHi09+MeNqdcQ1/6FOBxLz0FKQDkKQ3xmPp2UOEEw6CYk
8MJOK+0f0iwRONUjpUdsZsXGz0VprG6pu80xbec3HxVHdB1ncX5Wd6GCkqvEMB8I
a5QK26IXw8jue8bIhlq/vLiTmtA+j4ELFlPIL5J+UFojKJSxGZCr+KQjlwIaqdex
FUvxTEYl0MQANuPpsYbXuHIYw7dODUbD5d1HJwyfisAZZJdhH097Aqq60o7/ev1r
ViYXoy+paXq2U9STbY0ZjXsI4hUx94l6Ax5OSfcPOCGRleEHRS+FPEdEmOWoRvwX
1+9wVoBAZs1jUELfRXfvPOWGZakRz/JQ039gsN+EuX8V1yGPrJTMGGyREzqGoQjq
z1q916U7fN09hrvlOy+SWmMjnW4Biw/6IHJcNwi6sTDNc6rrXSJ97H5FaYeNOAr1
e7whUlskiJvAPWUWsQcnPcy/u89vSylo/6dWL5nneC0hfO7P2YzYdzD2VpdybFAn
4cNbU2Cn6LRv9aqpAxKL0sG+i0iEFvTgHI+KjBawi/ayTbRR8v79qlgaU9Nyv4fG
7Ullb5NBVDM3kX9TjfcrVfBFZtOPFCh/BWQN6G1m1RvTsVn74dDy7WwrWco/Omji
KDp+MjSH2NSs1opQ3PuWL2ezucfwQwzyWAxP0ZJ0suiSxYGopFl09W8oVMPskZle
5F27PE9Uiq6mTwwHZbipSwiPxkXxjd6kF86n1COj7R7MHvGym5TUpSLkqTg1N6J2
bowtXtfEN3nghmEHpEgVqgjeOehniIZh/dYmYAsLgqmpRmburVdbWJgaXl1DiK70
d7vnqE/eOQzdmkUkDVerDC2YTE/8bY1Rgf8jmc1tQRj1itbhwzD9idFaZ2YNpMRf
dJHLz0s0Q5zDAsmxHxOw75/D4hD0PSn2N3eRCAlKcWmQ5FvrtUFYXJqCcEq8YVxD
cHh93YTdstNjEBO7o+pQZ5AvGlFovtHJHW8EUKPe9TOAVhz4XhbIBTho7enQz0dV
Wdc3PFqe651BD30Jp51QGHBI0Flc2i2MnNARzXHkvKlMMAQx8qt4BCJuxA1GEqcV
Y7XUAaLfv3V1lwdzcsOWihlnXazF5kyhyIQHjioWBTdiif4YMY+5shp8OhBecJc4
C8dFM0NGMftrbdyA3fV9Fm7aDJTvNzBllt7RF8ez/N+yGETN6O0r9dmIGojKWvnA
6o7MdbRBt89iCYd0nrHqmmQa9I96ipv8Hr3vTlBqkGzMyqSXJrwRXycDje773iGH
3kPpLtdUSvvMqvvReccaLapF5eTHydYbNNM5nILQOkt2qJqIrNPGv0ImaN7VHsYp
CQK18nt++/UijIBygSdXfgBIjPsljkKDYn/lgdC2WrrznY/Le1ANFxuILqqsi26n
01s1rS6mkF9JZZ2e/h9AYVNwzWm7P4/+EWszgTCja0uotpVrt+9DQbjwZoPQuiin
yJq1RGaxtVc+kBfawyrOUNtrMU+0hAO9WV0FythO5UA8VjRz73Gw9wrrpnmb/tXO
iL5hm5mKyXSYNIc+Si5fyQpo3wF86hc5YVzLdh/g2B0dXDgFhToMj/6DU6l9Rker
EFij2qD8L+mMJ3sr3KPQZSjtwg+2eyHGfAJeqpNU5gQWA/qyMcb60N3w+wiCs6rI
oxSGXqc3cGcHup0B+2JCxZ74OIbjya//fzIMpdj3U32OzOVulR/E8J1CV/eEwqM/
iFdo2pXSi0oJJ/hRQRqrQ52SqhV57GSU5H855DHsE/1+8iS/T6UJIGWfb1crmj3W
44NSRLkFrK4sVq6i9807dVbCv7OrdO+VNBVC47725BuY+EYsBe8kvUMotWuqzGJS
/slKS39NIVbK+yD6+gn/Z7pdj2cGVj+3uGEWL/InGFLBv2ha0H0caVj15FTKGgT2
kJMiJfmddUMnhT6U0uatawtfXy5L8/gTpPLQSJaAyDpw06F/5IVq4AzBvFxpQbT4
D4lmzrOSnmelYoHvASJrOLJ7hcKjBjh5YYwjP8QCgvDARnwr7cjGHBk0ZAR76dcm
Ni4WY+OsDAm8+IXvfHCvAqBsGf8a1ss0kajCzIMt0fTqI7wUyNYTFyKNqSjgIIUJ
8+LTAZAzpROremGCC8JtYfKEycJA+1JPCtgPWc8oC+Vr3yfngazA6cb1p4HP4zoB
4JqVQNAE1DWzMVy2Ktno1lefcWbQVrLvOl1D0PsHhWbSfgdOFWFSyi0baY0MhYNf
ZaA1FnTZnq0VGybJNWGL2BzaQcoHpGWOu46ry8jqDq8XwHfKhXG6EfD9rGCMLBVG
yADMZMgziXU1LckpCgJ92uDp4O472sbdwY94SDzn2QEbba1Fo1NgdgGXo3Ffk0la
TfVS/G4rEScox1iWMZW53aLdGUHlJ/pBRYWoeyO0Q1YZHX7C2xkT3bV0bJZ6XXw5
6MYFAL6vIuxKWe5PO4eB7FkRV5kGuw6DFsTjeroanli83/dtJefhZyXFv/lwRQju
LEVWFfBGSwUGY9fVC6zQ1BdfpgYDLExJQZgVPjXbwjP7B+h9gCWwcOriJIA6qk2W
bN0gMujy58gamURKLxKYGMKN95Dy9LJktuxouw32AjDg55Aq7YmO11w8Xfzx/HMs
LNc0ErL9o8WMNmPwLnWCmwn0DxH8QnhCw7q/lqmsUtM7Wsz9Wl9YJkNxugA8MTkP
q41vqZ8ssJevL/KDNSt92quKXOO9wR1Lyk85++HuwxK7vSnlGu3VK5LZAndQvTPi
7nP7MLxn4SfEY/wJABJlsek1S/IJkb4x+QjIyyW8MWz9F9SU6ohNfF/bTaW/RvsS
/QJhDhkaKYrt7exvhCfEACZPqHZdzMuf/2w0nHIRmWouTh2hWpjLiOAFy0H5JFqN
27uV4DmEE/3bIrfm1UM7xZkh+BXPr543ggImKI89uZ5qGT//UfGgkln1wILKD92d
kdtVRgbzSLtT0hAk3DC+P9Ep0tM2lWYYeD3cgLak5rAWBSjrieOLksLvXPVu7xTx
Zw1Gk9MfGysztAAAdng8DtCsLowo3QvTRqoOPCmJgnK1V1RxN55+whqGcmX2xfFB
zBiihzmBRhopPCsPV2Qi6OcFe0kO4JhUo84uiikvsINevINvVMJY9awXFa8Oj9O3
+WPaHo4jXYZQe01Uvp7tMr5w+vJaqFk9X1l3p4xqlvA/JC2DJzKyo/b1eyIppDTf
LxDjltjgEEgClIjJGhyt77Oh+FKlT/6QwDyUwhkq81THwIEsZjoFXvp/Gfbi2xld
My5gqxd7WHg88b6m2AQ0+MmPjOTmF2Tc1kYyu3c9yGdVjbCTjztFft1QICqcB7de
gHkityfv9o7MwsVPJJgt2gTmzUcslMMST+iy/a7X41bu6EqfBMK74A1LN2jXsF4P
HP689uvpt/YuLacux8rcw/iTA3iOFB1Bb3zTD0FMKBKcofLa0PXTYnMoK1pI8Uy6
dskXodTuHGJAVIm1WPuz3ansNWTyxzpJhO3+WfLaEwwkk296T/hU75W92SiHwQS4
9//MsUCIqBlTrUZ419yAmhhTN/XCPg0cGoOeK62/AHZd5OmddMHmQu48FGptKM4i
RUrU0in9eHEPOuzokLwMJtBFO11dPV5ZEa9123LFKtfAi6UuEhoUk9yrDxz0XVpY
oS+2TpCdXrgFKt3O+szRZ2rgAsX6yUe3dInZd8gRUmjHNT9m7x44NYyq2NomQ45D
7kZiEaoGu5Qbuk1OZ7/lGUrlVrGx68WN1cX7ulTY6GrFSYFcvkigexyG4RJZGUkA
ATKh6hY4oxaUkn5NWnldLHl/UoiMSvkJmhAz+Mw4sJWAdat04h2a2KUgC1VOWn9P
/qkAiDmgBOy+XXZHInc10C8GJ0X/kqkgx+LZ/Ab96f96ug8q2ues5i+HZIx4cbMA
P7PMtsM+mvpkaBgug17tUo9fY/0y80gFbBIjDpPIEQKJDtdkeOKgsMcKaPYOatcu
u2+xHejBRTJohF/k50A0Ltvf5/VEWu7hGx8qKl4lAQ1mX6Mv/pnrifkf+MOCIu52
lpLamLueP9BSp1r/T2zRGZWY5BSZw/jnkVJ7mkO6R7zU9IFvv+tzhAzBzWxK9v5n
IrgQ+1i+eOjeq6qriJBRc4W8oBPiKfkYloERxMPCHVCC060Iwvzd8ttA3Mza1f0a
b0lA9TW39zQV0dTNl0iIohwqewGcDI5jVWXHzGWPwDRyrNkal6/lNg0PPAViQDcz
0p3Qr31b9uV+NII+9DvI2HfxJYm+mcMvx0+FLkmjqpJJ4Ir4qtRspp110O77pVSm
h09ow6pl8UiP7HPlg6ls+DIN3hWFI51Uqo1eieyJw00kXjbAQMIBqHhnvrIloTkT
qDp9ZiYQjCn25PhF7OeA8OLo9RLxS38eEhRx3VhUhAkgUSdnQ+WC0kltRTtm7Yn5
Gw7lLT5CGcJ8+KUnCgIuY+7e2IksEC1c/1EMkAXdUKvLCfUQUSk8oWz5W4V0qMQ/
2qSGS6XhTOKBdPttN/RvT7frSWW2hRx25sEbjJY3D1mX62nNBoHOVZj/lofS0rfz
51v5CRNO2AGrB2Rv79RUIMViFsQ7q6q/HNes53OYL8U82/uoJwd3j5O7hto3uoWl
X91Kwe37VWfrlX6uY0s0UwclnUG8GpqwdRZkV41nOQCnyvtFrAE75V0Buu46fxDf
4rChm29wzhf68kU8kiy+aS0KKpRXzr0A2AMdIZSyjOmh7a58bExy0SKHvIxM04Em
rsb61OzmwGlVoGrDYoBc08QWxShaFFv0pDCI9hegyaG9fvXGkeSa043zSmLNa6qJ
HC5qmZv8IDXNJ6/FBCObeeTZzqQyfJK40Cv306ql7ZG4KZTKrpyTo1ueHBlMIYmd
e6nfL1dwm88s1odt840LN4TAmTU39jLQqWH20OvsXFlHLbK7yy8vXPOTpQO6PFHw
I0FIVIm7UvPyPAFPWJBn01EDuCn/2Azcj41jZ2t45avMtgQZlfjsR0bNHx+18Z1M
X4lEd0u/or3mpD2qdX6z5gkrWutx3oqOIjAYQHBJFkpVAKEqMn/4pZVaVKkZH1YQ
06X29u4vDxOAhBLOYCerUircQgAWkl7JTVSCKaZzGXvknDDB8/x4UluUHoL/QPsP
UN1khpAy+l96nKAHC+eSE/BPPRnI16JNlZR7wUDImaTvm89CIS8KO2RbUEJvBpdw
//HiPqVBdgFOPb/rEz+ozNxyfch9/CqbRAaOLqSNDB+Ixs1Rjf3Slup+yNTb6jRG
PSv93sM/mxqrwVhoZKonWxIB2BsN4+p+gbXVynyQPX2rr9mhRD3puKljl8JnDoHK
ms6iuLmCv+lfvBiHOqiKmm4P3io3T0MHODnI/l3m66x/42BULiT/uXz1ewSQt31g
iMwVE02M0N9n+Lbl0JsdW9H0Uh37rs9TKLh4TGVmRI5/LMOnSFLymF8txMGQ1e2Z
H0Ee2SbOwbup0GEoiDMxPtpl65y2JVY2iJDN6UX50LM8gFc79VkBFuqp0BRlNLR7
CRQ2zbEDpnPlAT98y5BIxpn7AYAvemvDnagOW4zFcRXhY/CXf0t3XyNLUka3tONn
BkfKrlranYfmxy0dFdUjglZUkGTu24il0ioZu79zhSv0FGjCoWiw2mDbrjA/JrmF
foP1mAOGZ/Si4tXxeTBAYxMzltbb3NjzPEYddyFoamRs5NLlzEoF5Xs0C8gi/LrD
tYKtOZW7u3aYIjr8D01wJQnmxqAEigmD0Trk7EA0QwdA6UJDNF6xftERPAC6rkNG
dNT+DcqnfsoFTgbB+QsYB4URtbzEOE5LDtVaLtvCGCfJ3Lmm7itWyOOslonfRv76
pMFHFdtVQthtahwpKTnVSC7UC5X8W/Aa5RMMp2+u5+uqeqMHOheEjbdYiMgcCPLW
FoQuyBRQfnQ937jZAHo5k4irmNHUBQHyxfraN/B7LzwABYTQqLnmI3sPlmps7cqj
GtL3c0BKLBI6cBtxWQuwJJHvZotIrTkc7zAiiFoheIRp6Babul3vjap2lC4ARhkd
NnVOur3QGRulZCR0D9y4MqWUgVO2Bs81APL8gXk/dbuv4qp5qezkHONVtm7gZFlb
C+F12o6jZwFMBula47oEkXXG3Khr9A4LJ94LnM7llHFtar79MVqOx6i5mX3npeR2
I5Bqh4S6loc8VA80v1UBZoIZ4hjXgTS424ByE8fWf3ZVBHsUJGjDh9KL8MEUQ1hS
YkK9nTmmT9ty0a3TD8MIE/wI1QqZtQc0fLRN6B56r5MMi5TzMJb9TTu6twznbQxj
fAdP5gmU7W5sL5wkAt3K3UiRkrpqviI3+VP+pBUdNHbLd4nlb4H6TX+/WLYqNOzg
xP6N3j4KGvRjz+LB72VeF+M3yvspZLDYf6fszPjewQDMhXvoSoY5pbD6rJ0FxKfo
J5qDo1y4fXml50ZV+64EWu0TpNYwADH4VQ8lt6FoiCtuQjCHtGOiCaQ0dD2RzvtU
p9Zt9I6MgEONy7Bq7tgYTA1xoxmdG4GfRW2QlG/k7G1pahbxJaMmteMf/iWNGUDq
1rSUL8lRgKWY0Bkt/4r8shBxRqlfvTrod0BD5rtFaQR1Zr1EQd0peH8JFbOzqVoI
gCXzrYscKGpAzay88Yg4CpomYDg+DlbCTTGH6sDyoiDAsYy+RuRsV+EaInQ0XjjD
ZalX5EQyON+A2QvDd53C96W9gSE+vtq3D8RbuzXxRZ2yBakAi/QbwmL/IxBQcoD2
PMVn5HPkEQXIqJAxd8IWw6pJGDqqv80HUN1fwAIQqwDNQE0/df+iWEBoEZhobiyt
PIUeqJZSrizkolvlZP2Eb8IiWg07qOAdct+yqpbdKGOBaM3ffHCYF+5RjFlXV7s6
YqFmBJQljTLuYtHQLXf/PfulpFxRwkuxxUNP6+K5MnyCIBKJCcEgJrWlnF/7M4Mr
w34yU4jA5757MG/Bkh/TrFMz80UIp1l5ZZ16glVgUEuPlZmjeSo4HE67aXW+AX6s
RWB2B5ZXZwpqUW5u6XpVS0+EIE8SCQRet9GQiEUt+WwEzASMhHvqE0VKJoo+UAOC
p9mW4LSG3KrbqF4Zt0lqLTjTds1+e1peCC9LWgSpgdllMB6nRELva7jh4diOl3pN
F/4/KQWuuXD1518ctUG9TUAUZAk/iNuO4V40giRXUCGQgplcDH4csmf/GYiSHfLL
B0PwuKo8gT7IyxHX9U0V9eG0/wjPZEUujvzXkc7QncdNluNF7gUUBqsW67oa5cHl
5NrRENPCee2xfQwmXF8CRa/l4JvJ+dz1laveuOlmQcWy3c324F1TUHaHEFcof/sg
kDq/XlYmvKB55INOTK/fEIe0jQio4HvKFWils95X4O5nW03u9qm3v26RwXVearor
RW9DzRLZIGa/T5K53aDpDmZTpUxZFmvC4msKqRmcghvEJC+s/rrcjyYmCTFrJ1UD
8kwSOJNdh7q7wcKSVt50+Vo4CRlPWS0O4/XujEbfjMP+Ipaxwrqdo8k21cEH0yUv
8cs3uw0i1sASjlO1Sde84AtV1yFpkSge4VJSq6JhNynFx6c6Vhg2t+VmUEQOHS1D
41FmDS1r+CZTD9HqSspWUuTKVQpbm0/1+7k2lh1hbvMbS+CjKlaRCmkoWV/3qyk6
MmPb+E5QvCrLhqU2O/Wlkdcvw7ljNXGISfKLKcw8dz1kGvLicIJeURmGR793OG9M
T3bwtUE3qcfOZsRdRG/h9ItHfAU7/Y+bBplvKUly8vIJikXH4s2t7QgKvxJwjT/5
WGhtjrpEmAC2HK/3xmCOGYI7lgeV4ELm+AM20qq373JTkMkrAzOqFtxo7YnszBaz
fKRDXVzYwBtsMkpQMjQjPVNux42ezC4xbJogGp5ixY09L5V6V+LY5txZHW6uXIN+
EvIAssuQ0AESucIFBERor9onnwEdD3y/elK6OYyOjEEFdiVHF1zEppMLjmsDqS4B
Cfj+6SbdPHC35jimEyzFy/RhkpcZAjMHHgrQa6g1R2gedB0bZjJ6oCPqryAfFD6j
rv1c8C3DOViM4tgmIGdTc1jbjKTbiJm4dk6WXNIMHqDUjFa6mY4a2MQzdFctqC8w
qM9icqSeyowwAms1kaVKeDSOPL/7+9QVFnhG+gKFKmwbFb2uFagH3ZA9Tn5ea6Dl
pmISt4Ii7YU6ZppU6a2or8/Kcqo943kR+SIGQnUKLpl21tqhXznUl3KnxTWEWl2B
fJUStM2mtXl8BPmx5mdkB2MG/uNnlUa1xDyMjcycLWHi07L2OZIIyApptoY0bsba
4lpAGsaT1CtaR2ybQF2Lqs8MRbKd2DL43EIuzJ2UDDJqOoGxTq9LwdUND6y9vE7+
ekpml/peAA40oJHfTQtMQ58F3hHgLBkgPGLb5gfo1/Mu47UhOFGCMCVKw5PWXETa
I6Gr7cgNPjIku/kF21Evz3tA79xOQhJqKBKhXkVUkrEwFG0MmGyMkMUrEo0foiSP
qeNY8UNFxjEmQ+sZISMVJsvXtB1CoG3mcDGKPLUq0ucBxwGzx/qMwN2jShjv6PNt
QmXOrBD63NMX2bJw5bqndIf1/EScpIQTBrl5anJT6cJ18qD0QkQW1kNZhJrjbCiU
Cc9Cut629AOPkoPTRDsmR1xwt88H9fhNusRniKtTa+B1+dXYPJbZ0APiUtCehoGb
gVHx60N9HWDO2drRSMPE0VNMeMSKSCN3mxE7OovXD8MhhGIGhkB32DeJfWhY+a9a
nHJ2nfztrAf+eKEympa5apvbunJ4JkOBrlvQj+MJjOBwNy7kSlC1YnS82CQgVzAK
cKn9py2VJmb/1HJtXMDefesHmFDli/lUK9oiiZJjoRPcd1On81JK1d46dn1pJdo4
NSzhip2tFLF3EuqqIOReCNA+ezMEEfhnKdefJ2D76B/FW36HAttNTv/bthGr8trw
tRgpUrRMTgt6fT4ktUjqO4rWs6MfEeAD1fIq52zGRI1I+R2r4zkvOqB+T9ys13kR
BmX9giJRfjBe1eYqU0wX/kXL0joQdaqQcmqj2w9syW1EEfSMHscjqHfNbanhYcoi
mSgtXzB1QUr0ejSfVKDkez5hy5ygntiCXd1y7JRit4MIIyaFsHNujXMVvJGuS17w
0X7eQLsKgk9DQ1zBzbTAze/DLuCcX2z7rRUscTJfwiUqINwluDWMPmq6s52SOVhp
0XyaysD8+JCCRvrKVO48ZfdmfooFq+7zRyHJhWuPRx1GoY08QEe5RDiXtoyjrMvX
u8NNyKa/FKn5jLKnJgiLokxfSXSPGPa29dvX3t1nlgDyzhXiTVKECmfsZvOktBA2
hLJuzDEaKGnUQkxGMF1u16UwC3gcczFls8TP5Hr0+JYWg5ZEU6/d1zBnl+Rrs3xT
KYOCEtUmkgfjz2e+uMQeYlyJbKHDcyq+WswsZiDV6XO5y43vfjoLppM7W5psxzGP
cBklg0kMXKDqTiinSqm2AdP0jFDmuxdmhvDTtknW4pgeojlgQYKGa494G5GX6QNh
H7B9/hTCT9dZA74z2pJyqwHq01J5I5o+tooB686ZvhVeIFz7rSwweA/9HVwSO8o7
DXaLCE8cg3MKIKzaHBHQ96ZrNKkjhuFR/9TCX24sf7BuVe7q2UrwcsAoqNRmPJW2
yr2J97NeCRwPokla/kox/bMs9pIuWoirelY874+dtOfxdttPhB+tj/MH3zk/MwPD
o70ZzwToExE3yu+Dcjx1SMeJyKyqDmI+6DfvdITmlyGpWD2Xf93eC97067EpjG0b
wKTm8FYoIlrYFCj4fUTp9/pq0ZErWNxYOg9ziCe30tMCeXcQ3aSmlEKFFwLn793h
A4v5SWft7UKl7+bvtlxYAbYXh03phKAn+w5rgMl5mvCiz33WjrliQlOCtTP5vWOj
/NqaN1Eg6AxksNtfvViNU21HWaTlMrsuCWQF8jZc9tZviuwT/A+xFo5WrsItYUEL
hGK8JvgJFGCaOlkMxAw/TR4J9j2GGqC+OiyVPb5nZwPiwyetdb0j3CDiODTJnCCW
DweNVDdzVQYPZNRhBSVmfzown5Mn+H1kNJDBa8CC33DzkDRSXBAi3GlILQGx4ss3
pGlCefwoZFCJFYjyqqC/9reWy2XEJpH9GY0C0+vU2mmXXGDRGWM32WpmFlRFUVYk
bXE00ke/nb5FmTMCs34d6kyjMMoWXeiCrpQEWuf9AabwrNz8v254mANjJMMWWuFb
u4DO/iayYrNmSjMhYBWn1i/SBl8zXTsf0tpJqvEIZyh7QMggDVCZkwulHrmSa0RM
NasgxAxRnqbGf3SN5FtMCm0hZPkduAIqes0NNawYdnWiEDJpZ9LGguwq5C+tcURo
uj2tc/dIvi0wwQVX7Jr+fJCd8inVG+T9Fwtygt7GX+KGjey3Mt606CrUSdWWkZpd
IGMO9GCC120y65lMtyCF5dC6OB+XY4sI1JuyfP1X12RyrUR+ja4GgLK9Z6msjBxK
f5N8nFe9nwnLrX+CyDdKT2REcBlcZ2bQMiZpMln7LY/Fo1d35SyHEUAdYG9RenBV
j/63vhFIDHJpUtK4fb9ypQ2wdcQnFrO7iKCHhbfXQ3Ab7NEcZ6X7DIrrsUfIcaig
fQtTV0JXmvW3sPttt93qMhZ+kwPynkuzb8vaE7C9+aydCSitjbfXk9Cs7D2Zz3uK
FM0tp8YorCGnekp0Rew6HPDn3fjqDOA8yCZmvaTQQjtriCihtQjpB6ybb075VJzm
AIwjIZQt8pfAI79PYMrt3lDQayudy/R3VY1fZCaezWkObpv2rMGxehBU+U2kqnZ1
2VCabd0bMJaAuASd18c0MfZ5q6suNhlL0UoQipfUQJwzTvt8qT8UW2ijnju38vTb
TCJhgM1fuNxFZqj+2xrSG9hpV9zQa8aS+E/rYvKmPZK1uUKuB912r5K36zViNgxl
UIWHlfvHsjvErZ9ZOoxMmXzBPLXHWmMR4/Axvzti8y2F8ne84HfAy7VSCKKZxMeK
8+bMbxqI2Q8q52nXIKdTwLSsm9oVDo8UqJUkTv7OOri1XS8FEO7Er5IsDB7oaXU9
x9z9eSWd2twKGxEGmkfx6jPdBfG8gaVCjrUx+W3dHOu0M0TsTJb7tqtkKQuma1hA
39Udht++FGODSG13mDxmfRBQluvqJ/UgO9GH7hUAhwwU20S1WzbRC+r3b965HKQ2
NAHvWRzvQM8dra6dapzQTHprZVNWKF7vdQdeAP5cvEHoU7hlowN7Y9t+21cP/NhQ
/0U9l7z/1t30j/UunhE+ux44XptOytZKVXLHodyva+Uz5fhvHjKXs+EzkaOllVBj
2bn3YV0skGfYQO5Vkh/6Bo8CF8O/hdpGIEIFTX5rdl5Uu58uOsHQzKBxQWsVB2B3
PqZ335H2tYJfLsF8tI937zVHg/Y1iRYI6cU4JV162lu9NNPX8BEs0OzJ6bf+0WWx
UXuvwmIo0kD8EYcNRD+m/mUU5Cjc+/oowSJGHO5yrWYQti43Aukf08SRdnxJc55r
Y68sljzmUag1EzG3cjvzpa87WQ8dJJ+bV+0bZd4RFR91AWaGYj4xOAnMrGt4CwNa
7n4YEwSQcIBfJQ11C9Mr4FlZTcIE5SdFapfUK0/OjMZMG9OxedjrwbeyBvFhgW6/
QwIGaSTAAdZT8TJyeXfUeDmZ3N3Jk06/ibXGA/2iJ6kFxVsbykk5tKAhh8x2B2au
qRkxyrV07TaWtfobPGRV3tlHX/GgKpP3GB6BVAKNNbxJf7qVPhp7ipa5e9B56hfj
ppfkbB73YfqcZ4/Gff7NslMOM6PJRFny6ilZSctMWV8JS/7RAVf7ti6ABLkDDQZn
Gj+vqxtH+cvrtZrTHAovUAssTITYzoJ0HBlos5Yu1h/ti3C5kBHdLkj1uSn03X45
fscIJo7Cwu88+ESe0zkIT5RyycpDceKob9t58UKRIuZjEvWd42neGVoDkPrnJa5z
oZ9CQmv19myUSi1q8QgIxhFyCO5UgOUlJxiiwvoiC9SvzVM9NR4GOhghQf3ovMJQ
Dfgv4QMkCpm+KpiqAPzc87nZLliyb4IWnq7aNY4LSk4GKXCB6T1xUwFu99164Nbk
2R49hRS7Wc7TQBm3091TH4ywd9vGUsBf5g86zwaVRPdKaWzSbDL4pQvFHAjNZb9W
LxOG8f8bH4ES3h53REfNk4uSYOJHdJ/TuiJT+AvSZc70Wftl6c3EQYSUKDEwGM+i
ApKq6ey5eb/IHO0nz32eYoFuqDcHPn7uMbTK+30EdCsjO68qjxxVfWtapgPzmWs7
z3hokMWmQGMnDZUfkHMJJuG1nlXCC7V3IrJkj0C4houEbCqfuf3cys0sg/rNw4B1
svHzBQo6yFprjR9GpOl/QvulWlQEuo7kSc2NJIiowoJrliLGstnxLLRU5e1JDOGN
uNFjMn696Zo8N+0V9gyGM5mkyW2RkRc3Wakpvy26QLuRWmHOhoFbWeFv2brZOBZs
TsToXxaCX66vpAT9mss+yKoLv+zqPNnEdEEpzH6UU0kiGr0ampnH9LIP0Dt+Fl2a
dnQEvNyMSxRjSIbhXGM7IY0nixIXdTcp/Lt2Sz4h9QPEV6KXikbQUu8syXxCe4KG
sI0Awd5W1RWFZEG2O/agGv7o5oME4BbdCJuFYEAqBtaUshTcAdcCm0nt82ZDiUuP
FH9iLkX8RL53fHQrFomeoIjMuo5HdULyJtzDyfE3g3LPfROvgg6lCDvkxMr3LfSU
wKvBsqiLQ68+J9TIPpNBZjpszSeOJJSOWoAOy6BkRco/pjlSwQIXHuIbp/wm5lj9
nUDty2NYiMX+fslnGM6gsatnklfCiAquGXwKvbC+ACE45IbVnaSbe7+b+luD842+
p+LNJp6YvmBGZ204FMISpRe9YoN7Hlysv1aJyMX94M5KvN+AFM4Jb39qezvDyZdX
T5vZkK67WO+OgvywzpBcMfx+ivS23TWRzJH9BugEKqPN55KmyKbLZBoEyfKOGiUu
fpOSz4o/IhkPyL5hikmqjAGrq09Aj1CPAVDY1YUte4ZI/UJSNgT7bSaiVDG6MFYi
xR9V5PxJGqlwo9z3TdnH6JukAj9ezYXgilEiqx/ZVYk42nSu350EVmyHlRq1xPOs
ojeXurM913givlgBMjHpHtbmvUN2B3x86c/6KYexc6f7NslPWlU4izPBQIw3C/lE
74H4I+daekDHSzwUASTmXl8Xs0aeR6Iw/GGm+tC3VSM1/qbWxBGerv4Hcqjoe+MN
YWbZhkBtc4n0lMRVTgWF8ZtFlwTUvTSOPdKq92L9teeCV39lENnz6suShk5g9LkO
zaalIRILjdNwSwObs+NDq9DeDZJMM0sZR+1VjBqGpmxlAWcPuC9RqzpOXhXBDV0m
RqNUJ/DCtJG6fftfUbk9pdUAnjnY3KujKC0Vv3xlPbZ3iSy/S6JmyjZ2vTRnI2VX
R/xr1GwfhoggWvNyXjSlWEdA7bKb22YQow8uyN1l5iuh67mj+AQibbXCSG0OqmYo
rqohhgZrVGD97/juKppnGrd92t1e5BFtX/DQp9w+uHlJHSK8tR2ZWTFO1KSE+4fR
iA42gr1hNwthIu9WqVHGYmX+IZfQkvdG4U1gBhTKWtflGUaUvBlJp422HDAWE8Ew
APXueYwbdrZ9S99iSWczfB3z932nlKc6Uw4NLLrVWrN93EpzJN3OCroP/loBeluT
rOjMDTvy59nqFpbY5FHxir3yBbi27FMUnVtIs/TDmDVGO4WqGGNCXntf2Yp4+vgd
n85tEAxMatj2JV8PHxVIKE172lWxQA5DHJfmp2p6v1UGnPxcmqFoGi3l/D1hqDWX
Y27kuYG2d/ev63dI5wJ+duiMXCwJq/894tlY0hjLQfqbVzAeCyv/MoNZnynVpCSH
C5ukvfoYqGDZhonE0Pxyb550l5Ay6Ihn9JmUbfESljMVnEMLBFFO+e5wHFYNxxEw
tUSiFv4lnpB9SnWDtVArgGGdDnBv5kvyzJK35b7lMZPtMy8GgUKKvJtuCUDJKTuz
OO5Hfk3uaZkSBlSJ6oDzZWAEmBcyEYu2AxGGqPDPW6PQ3pnQBQM/8j7hEV1zpqBp
ZWdWBEguNVypl0BzefuOrA4G9InUhcx0g9hXYpFZk/qMMUNbHZixwTd1wy0d59iE
EDhbgGdCZKpVWWxwY9axxRn75tJuNZU4tccn4nGFVyd0/2K0R5RwoVd4OfKo/JlR
qpRNzgYU7u74VIjbgl1Hzq/MAoV5ehfy1rmanT7U8GL+iCyN08gnfDaBBKPLhZMV
UlNBcDro/A9LnlwtJbN8AiDBlrH0DjLqD2NhLS+GOXsZJoewQ9N4bBTApFRQn4CR
N6pOWeAh1+DTvCnbCsR+unxHDEs4a6uBhwZzDiKL4VHyJus6lGmBJmUcEp2LPp1i
QdV2gm2W5xgC64a1Q8v4lVpcVSCBiFnBtjmhSyMFh4zuaeYsjBeAYb+A1trOqApw
XVYDYtBii/LNCNb1+bw1/n+jUQ8EUoZ6i19vgTuwfeAE7t8GZ0GwrOFNt5tWwq9e
sao96e6nJ79D5v8v/T/7C/anuG4XZjJdRWMS/ameKiCQEeF3bkjZGIyRA98rDFna
/d56VY4KztqSyXkzzzStCq9VH4UGSSuZs4IDj1x1byDBIpuTIgF25Xcs04xjO32K
7+bm0vGQ8LBz7ezx3svbZ0LfpC1Onuf6ydw+HJy1Sy0qurRg6I0eUimgPo4b+O/l
I6tkARIuIjoqnayOyR6PnheygiuOseBDjkvubK7IEmcN3vKe/BCkyh7Tg6PNJDxq
qA163AqOlXrZiA0P420MgrerecC88/u8rGPlUw6KM3vMKKtn922211BZmI/Zf9ul
rvkoRwvn5IIL8WlGMBplgnXtOKkv4IWdX58oNWMcDeVw1XutnpsJhsCSe3+1+r99
kqf1uplNUG30YxsDN2qGZdzKeHVsypr+xHOz3wpcd50sPYE2OA7xO8nN9v/Lh4nZ
QmimgN37jtP9eeIsrYLXdi6fF3mWLjKdtIvFTfRHC0rlLd5D+y4dU8eMfrgTdekM
0DqM+6Wui8p7QeFWN+EZputOZcDsn3PYAEudfYOgNLdUQdISHMRBpuTRbL+E4kz5
FVNwXx6mpL2QnMfL9Sm3XAVIBG4RNny4HPS5M7uDVyXuh5p6zVBCHUsx/GBXHsE0
4gFkZKN6NcOw8eaOrhOfn8FYBxrjc7R0QmjefDFLUtgldFhuOOYSz62fyKo0YF2R
kfUPPcYdWmNUhY/VMVOgnmJHdTMHxxQ5GTaPAlmM20rhtX0a9x9l8U79WOxc5ZWz
mqG3irsm+c/lFZVdHaUP1MWMTBKsQBjljk5II7fAais9yO1ZUf4CncivuQ7q19+j
c71CwsbcRHjgSLUl0Ov6GwYqS1DzGOM2etAxC0YiT3fI3OK/tkMlCqsewnFoSIlT
wxv8jy6p/YO/ISNhg4Izm4twTqvkrbos+s1TlEVGynMGhvSElT14b0RMtpDeaatU
as/FcmdjmPK8LIC/fXvH25YrPlrnXBTWZEjBc2UAXb1xEc9sPfXzh8b+dRuOszmo
Ks2ACoAI9MFnBit+myRcKGhXVzVDV6TW78DZjioFUVian4kezI1kF9NELtG5AEYQ
8hMXcOJmxtWKH9wb75DDVTWpAe5AwU1NOW3gtuVwnnca98ODquaFGL1DCZpYeXj+
mrYgi3P98dkIsog17x0FACWszAxbMLa7dLzmSsRuUUgXvRY+o8gLeyJEAiEYjo0J
8T9XUuexJmKes5WLiXU1aNX3W4iUoyMEDGAy+sfoMz/ygZEWhGrc8QWknApwgcw5
YRQ23JvoknBmueOyh+F5RK966v6YuI5lFeY1UoE4o4mK7uWOPBV2GGDnlDH0QD/k
L9GWNLM9MArQuoP+N2m1yis1M4hEKSmviUkQDlB8XfQCRDQ2qCA2WevQZekMVtkE
Ypu7pJa5YFI8cOKvR+T1eY9P/5Bn0c6tqPU3gXAmIB/H0HGbBd07ocKqNm2CrP8Q
0e93QA14K46Pg8pd17YMuz0F+fHD8J2W+sWA2JJojWsjuqHBgigY6VXgHnk8UZVb
aXAzsaY5o+CuNTYIhJYrkDfXuVHglOXbJ5pVVyCOl7mKi4iMu7bQTHMWg9FUHK1p
ky/J+V8gyVxSKa8n+/PjWRa53TiG12XPSDFRQIdz3Ee3hvhRcsAzFqxnjI+QwgwU
+L8oJU8/pbqqVDXluK7hjrRPUnLLxS9MsR32SfU4ZKJZP26jRV7yO3I7VTNnwNwI
ohmwiXIIzfWa/X3QkTIBxqXKqZlmiZyQn9fvuXW6sc6sA6m4Lhz796/NxitDVo8m
I0EMV5N+NR72t+mzf8GZjJGWwhDmkyjDbFlu7Gz48Tg3UvuYvnmx7IGErlcqXOIz
16qWV+TJh2Vn4WSc1/ENz+YU2IXT8fB+5vJRW40WS7VT8v8fyAQ5q0IIhxxBXLrk
gG82tKaPh+SmfVXzHIfCnqGdViIjfYfDxTNHzwlmYb2ISyvSN2Q6phCkovlcYKbp
5sxXW8tPcQs2C6vvDuVA2/STOb7HALPyXeaBS0aadzv9xIUnDO6xHZMcvuFc/sBC
aHuK+lCBWdJHNyR4etWF/RE/XxSZlZ5PmoyWlfmTuv1mBiXrr6pj+zhFRVF26t49
jtgqQTDqCsTAM25tfpot79zL5bmoETmfPoMiGqYGKL/m5Um0z9B0qveNM+1uokvd
8b63e62yovoX2h4GNQyngAQwKwmNVf9Vbni7DClff2K7PEThkNYMI8+Rk4X0jCWZ
dHQl9IaN/bSmOjeZnB9SXJjkg3zpgm0goe/7FoM5CDwzeGFJUC5zR1Jd041r6S+X
UWHaPk/JxruX2f9UgAitDTqTt0xvoi/TyvFjEebLsKqspposbrzscZnB/cjdZdOf
PsLeMKl+aWbs5El3Ewsn44BzSScKO0et0YB4Pqu4p0KIG6JkFNCQTF/y2tbwyHv2
tVyjIvENNn1aEP6JZAsY0Jm5ZLWBJQBid4x2r1PCDIvlOq9Uu1omrPzYKpZ94O7f
n71BZu98/D1GLeBQ+l+4FEtWUNxQ2McFzF4XJ3bL54hnDKSofOBkRDb9bypzKeZU
TNG4Y+OhGkjYYuXnmCfDYMxPMDDqVuxvnoTaSOhkbQOOfcr1MhIeTmyuPb2vcRZz
vbT+RdFco5GOSDsMpUEgp7fJwzwBeOy0/W48FdWj0vQtwcBBYBhCQiaSApr7afsa
72ApeNK0I7l0atuBODfan+KLfaxGwptjabLrIr/mo4Z76oyGLkSV2g2qJ/g/myN/
k69WTxgcY7YhAmhXiOuKzqH81MgEZQPw1eriyDhL+ipRZQ6Sxby7iRfAmZcIPTd+
/FVjA2OyBVgORIDXiwMtsCBWRimA+bfwETZvmXJy7+Hf/n8dBrdHywwfTTmovZyq
SLc9RfIZ/SmhcF3hcc3cVJ5Qc5+9ogmO2DczhNSKZc/J3gDYBDyHDEfDZYKMT7/w
JgAudbi3ZqK6nMWkQaNoHIjTko/ATn/AKHqrduBvpKhfMV0YrJ+9uTDHStwC8XQQ
BVJfkWrQgY1Pi1gyEWPFmRB/tvqC/6mYTgOcpK5BrdvFIftL1tQemgFhIS++zKNh
sUrHE781ijiMXV8zsBQTrPCBEX+7yEO17cWEjUkV6mvzZBUE6XiU8Zo6ynjloe4b
t50F865pgT/KUTmhe6l2t8bmu+WXFHdJCeIldB9RqlNGPqArLrpZV7Nmwj58doUe
P4T66lar2fUNGCuN4alw4cCEuIxDgbc8Bi3dTufzRAoC/qyUKgFTZqAL6nT+xSRf
pLh6iUoZoai2aSsVZb/wwJ/z8keIpuPyTHn5+JQIdC3oeb2E2YU9gYD1mdTMyaEL
AE5Ihq5jQ1Do+9WHl7mrgnrOAV0pdMWtkr7GWlOZGLgN2d3CGPxdosa+PS7yB5T3
HO/UbBP++c9L6QB8bkLmc8SV8v11KQgfqBi5Grhex/fApdHMGTEMbPbBD70XHi2z
AtvHsDQrMrisjCnnotoHIx3UG+h4ISRWTSvxRF9pE/3eX3tKQgn9dsYEvmYl1McG
jShyLThVU8HV98DEd6jNhWyd/6GP5maEV6DmMQ7mdbO0XjJsu//EYdMU0Zr2YMDI
NOXtMm6Bxwg3g4HWOWaeHXTP9RPfyiZIzEFMx5OfO83Jhj+jyVweS+k7R46OnmRp
bXWTrvGHCmIm9sjE79TsDQrySCZWt2HTYISPS9OdaXz09hUg+5RbHU3racp0RGAM
1ALhDRwOwmsPuxzeamD9ynA0N2TcuhSdsaE8B6tsx5KKkLDpbOgAoObt6ez5E9J3
2Wd9zAqnrvveFr9tr7ldsRAWlN+zQ8cekk5WWsvVulIBZdX+ibuvUjPRASmsyeWs
fYpG0oGpniec4mONAW+erNI3n4b/dyevgfmDpK3Rpc1+/ieUyyJyCGSlUSZEqtD0
9PCMVN1P1HAR4nXStMdx+1ssICaYe2k942++DEI+PIf68bixgqZEvpJm3RCh9wB7
+x11NOqt2k4ELld1d7DjFwaTGbIrUqQ8cXj9Ertuax5B6TBb+imdA43Hd3pr3GuN
VdMqeuVIO2u524qJV4yeIWcn9O29rae1hHjwpvbwr2J5pcLU7cjliGPyrwJhO0mY
78sTHbrEvVfEXBhiHpUFeNI6p+xBx6N5HrUcfJsbUzUBfNmCjK428F+xCZG0/cQw
Gu3OrNFy4ydCklGpxJJI/Al3bqUdVsabhwtagqpy6N3S1x3iKC7mdTHAnpTT76Em
F205WYg2dHjKSwZy/Us2I+rybYtgqHrZBLRv/syE5lDsWmVXkikgXpV3B0yfvh+d
9YwE+jTlylNuhJ2GTmAqzG0l/FK0CusffjHlFqMacjGdfwaiiy+UaE9rOYGbxQ88
VpghWmHPs+oOWJmXjadyNFG4tS0H8eRdfWXiOiSGlqpl7eMAtFwJq0EGzt1aalya
SvI9jLUzPkboLvuJHxqSjy/fvdjFun2MoIvBjF60EZesB5sd7DvPLx6FCCJmxyoD
u7Q1u4ktMHzC7MFDbdB/xdkk7fxjMOX2O9u0hXH9UPn+fGUVJYdIr9roU3tTeOas
3MWf0IkkNI8Hyl2kV4K6Lmi8SXPpkAbtEfEwDDofD8nGfOwdtfN/HpYd1UUqr6ch
xB63D84Y4z3Fpl7sdVJzrIbbCJ6NZjVUX/OvRWhP1JrY98y/aUjl9S09gs49YuRb
sxjDm9u8Q8RhSK9bMOrHesFJQRk598+dUJI7WC+8jBpzM1I2bSsHFnkr2+j9aN/Q
fmde969uexX6V1KujGHhJIvLPbBS+Ti7s8u+6SRpwJJwF7Gq4ge0pxuitouNHIG0
Rn3ce/uFN/T1Q7Sp1eOD/rpUwTlKU/U+pFoPP/143gngK/erBFMq+ral4P5y6RCA
rabjQMkSIIeaAL9yggpLlxxnDHPZhTkyZJUNb3qquG6qJe2a1yLRTTHd0UaFssag
030M+88h26lkBIMxBwxUcMPBzOd5PeBMZAfhLXVU77tm3Dc9RNOeXeXZ/APl5eNX
KpTYyRSHctiUr/Ca7ZFIT/UNJX3RwIIb7yiM3Up7TcANiOB++7Zk25dpbUhQPIOD
aUWJwRDetq86Cja45oFfifYhJsPXhIknJlnkEqdTmGekaziuvbhyPL7bHbZJCN9Q
ZKT6P9D2mKjz6/NfG5wg/6UFt66Ul0JY3ye5t28exxLjWqIxZ3DQtspvXQYf/kgd
nQ2ja8hHGZ+8dzI5dZbMvk92a21k6aXchcNyoIYd3q/WIm7vRLWVeJySQrFlw7dB
4nn1gbNt3O6l3TkIH7zl0IgMu2FRQa7IEihCheISxkK+Esz2EvZMO4MUrfNF9TXk
pRcX8U9IY/GT2RW9uAUjFZqDRK5IIWpnShyc+/zKIM0Mm534p7XmufBEyj3YQYiZ
ZnIi9O0poOTdBb8jbQnbF/bKzxZtLwW/dnL/nOzkLg78lrpZruhyCb1E+ueY3PLe
BOxmuJLfAsyovBZeCtuXqxlaxivGNAr8I9SsTHxl+ZEDQr3QBv7iZenYWwXVRsiZ
q3G6lKSThCSfgdocUVKrpQnj0lefQ8wvCTgqTQ9NBukuKDwMDVsKEasXoAAgOySr
pFyGvv8nJ+cpb7jUk9hJLWxM9/xOKtuqNomdRDHFHIomU6kqwjHrkSkTxHhX55dh
g67TUTRDPSAPCdohrEzxe4NeBn1dRHOVD8i77ICanQFamSZXwnRjdJkcbl/knDjM
OnZHnyQaqDt/sdzcyZUQgPXEyCbFqXMMp8CtDLfCsSV+t0KqBMgihQnUW/Teic0x
+nrg62V1RcYe7O9lyfwtPu9ACQGOeBF5H61cfHTZTzrrs366W+YlVv4hoiqvBAL8
3xZkTzoWSpa8H0XNJZipB9oKmKTCPDiUNRtRjquzu+IXI2oRSatbsInf4Nr/cIJi
6LAn6j/bo7xG2pQgQBe5f8CUa8FqV6pXPEk5oRM5peXne+Wmw/YJ2fASnMUK6/8+
/f/Y1JOOWlFKAg+FT6CpWIY+qPqgZTC+sGvz7Q9ANXkrOp7OkNG9EB5m3cJG0Dc0
dSznqnb1yijKVkE3a9HL9fHKzkV5y/6xC4BAmxzQM6x2PXV7tJldBdXniFJSAcIi
rwEods+o67t7k1xDEgj6kadCgRna4hbY9IX+wpxDkbHEfnD9XnKlCAZlOA6dYku3
gFwPiQoTKlCGjnt4752Md0DZTOs460CH8D04MuiArc7JnKOcyQAyDCRkW6NMZPP4
5I3usQQVtqHU8j4B3z2iFa4k5Ka8m3Ms/B4mPbVgCofdbE0uiCVDHHzFNM93/7Hd
iRB59Y80DelUfyqt+mn4FHAo/X0Q+XM/EfI/1thmbGmHUIpxeYPvPfYXpsM3cj6+
tBmw7LRudlJc4zsmPA659FAQ5GZ0m27BWqFy4cbEeBPnNx453EMp1aqd7J83YpNL
Hsa9MxzwtRW0NUMTzM64kcsvmItkKuqjpuzZwr8XejgABfSa57CgWu2qgG6Z23w9
2Az4yTf61ZewTRdeM64Ne5hBoOf59o90mgjpPezMnFtLs/PbWe8SRGhtAJbvoNFl
EoacWWRnDkwjUB4C7LEnnROfoyC9VyZxlSHEAvFI92KFZj0ElE7WxUcJ3Wxi6pbg
tl6wgODfU9DFywSv9oQIKV1snBCawmWKwp5pQKq9QFAfYmZ1qdy2uZeedYNoDpNl
Fnr2F59MQOkhckc3sV2XlDoYtQRdyF3lI72pgUec9xrCzstn8HcMO0VkFeL1AUCt
yQ5GxKdfalEiLrQF53R94rfky7Su7XYGfRev1lZhWaivhjDRgUM+kAqKBjUWwrGF
geLcBb65Qc/+NFueJoh8TT/Gm0pN4jiAWRVZoPWh5B48Uhn0cgn5gIMA9YOku0rl
eZRuqkPMUT17JSy8CFb/d01kcFaWnIPsmHIttuDiO474eFyKY3dTkSV6X2tsPXp4
WbbvjhJ8DUx+cROh3oWIa9b1+C0hZJ9dh8/oItf0+U4vJN/Oa3cWgYSE97w9PvOt
b4D8tjwfS+Pit6WuVYS3PZT5s5gNOm1FuyKHEmQJMRlolQTBoyUm9vwNhA/ZDQlc
WwCbsbmKix5WKp4xGoboImOA+4qWRtUr4jfLuu400bfOmlp/4V46Ahh6pSdfmNU6
6F2XC3WN2fg6jWbaE6kPzlrQSYsSYOHeSOc/y2IjYVOltoUlHAFoLFVPvL2np0uV
M2enRz9AjQUO6TJ9V9ZI4sZ9kvOC5eT6yT2dVrRI+bntldgU02qewRLZJLXR8LNG
RzpK919FEXY61H6DzQuJWH/SI2pQUoOD2t6JuAg6Se03vRFiW2AItPTOduLIEsaM
t97rPJpW9bUuL5h0p02tGa5SVAMe5sU74rvKfLxemlfx3rk9CEXed1JyE2zN+RhZ
YNliMx+dCOlfVYXITmWnZyq/GEDGjlHv57PE+3KjdPBSK6eUyjJPDZOUzfWOkolo
UfZbUy/Omsp+CS7mCHH54ARyBlhIgv+UFXj+ofmmOBQstTkkOEkOEwJM+HYR/JtG
okH2MrArf+Ceo+byWwwP0kJN0OZneqewFxi34KU5f21nF9ChHOZRpS+lxekRjAql
ZHYDaIu9yNOI77EJdrzhMH6BDPCe1zOsy/LzMEKdmSCBECzILvivcMwszVf2B+Ar
yMktlMpQ02O2ARlW1Ik438UwnhXqBoEktDWpIJg8SmQ3CILUCTYRIa895B+T4BI5
4gqISvln7o9IL4thb8AKn0/RJ9CJBI1QIRgXAG4g/Ys5YvxbKdvdwqTRIi3gu5+N
FsbT4B12QD0cgRC/iquQdiBeocl6E7rSsv+qICjmAdI1vDwoq4iP9KoCDhrCyIPr
XFyovN/6DlChQM2SCRO6XtGMb5AcgvTX5eY+jQ9UM9fTKfckYTrWaklh6SelL94r
kShTGE6cYop4JZPc0H6q+5NDP/6PSyrUxYDVJo3GKhK2nlk800hAsaViMrejS43d
SDVz/kuPAN3+iiMrECt46QSHFA0sIaH6qVo6yKLTcEd9laaBOVHkbMM2qrIrPMys
ff0wJJ1tDuUp/bs9KMi+RI3j80ZDmWmnZuDcN7q1XxU+s4lqLyOZmqPnvkVxePTr
C3MG6MplgnKNehN2idL/GZkFpTPnkwVBoOxwq88rabD4V2byqDtOftngT5SYbsIl
Borjduws/pYUfi/hVoS8nrnLtxML3QPdzTfW1nU+uzK8gpQZ7ckCWw4Zh5XRYe+B
SEAkpV/a4mDoE1WPucLGhoM49FjmUPzB+e7inwByaqo8cuT9zHPPuu3r9nhJWakP
l6q/28W4td7zkZ7EP6OgsXRfETP1YN8q3ehyKO3XiLKjjh+COJMsodbOvwqyrdrr
9BgQJIf0VL01YAaaIxay94sA4rsUPRjNJcnyU0YBg/RaOn2UYTglg295Q/C3H2k0
HfuhMgVecSEgwmbhHOjAwpAHPqag7m8oEKh8XoUzC+6gQ3QH4lnCjkgIbXTHleQ0
KgLjs2jJojLYFTClRfIcgadNuToECZpCHM7ZFXCI+wirctu2JP9facTmZb/2KHiJ
TnJ4wAb8wtFTqMy2HVv64wBljITDvuRqRB8f1KjhXN7pZP1xSSNWFP/kcEWeq3Qq
UtL+NxkiQ6FHbaksXfGICmzXXBl97xRMRsxNRIbu5uoGneAJyY5M0jNi4x8qgkQa
BuACjs+3bzp2+ydQFv4Zkw7+CYvGDrP23eYf+fwbZigPzWpDGA1Rmdh1EAaDdbVU
0orNjpog3HAibxRmPyKG2KdNh4otfjxvVUIXAMrV02ttfQAgTbQh6QnmctBQuGn/
0nHQhCSIpAQ93xKPJgDRzk1i5IawJsPYgmUQOQZe4PixlRRft8If+TVaEPCM2UQR
LJpx7zZE+FZpUERZA/x4wxgNx9zI1s1gTKW/W8LtC3bhxW75SKrN1+V/VxKmKOIm
KY3PZ8cjdGqHgNOKQxZe4bryFf6nanbEDEi6lPVmAkTkMUhq+kQgIZ5TMy1nT4Gt
zpixf3WUN95CVbw0Feu6YBE4HAJgVE2yaAXArBuUVn/XZv2Im/8Oe2mP2B9EJ3Vt
9d/ghtPBy/3PPq7si6dRPyS0fkbvk0wVmQHKJNWjWspiL209Df68cgCktKUiuJHD
B7CfkR0vzcVg6nsNDs00YSN+Mr4UFdDzy1TkBU+o811Sd/dRASOCbK6kZZ5fHM9N
WL1/hAnhxCudEd0FyySZKuOlBsT7HriZzzeeQsUfDsqSjan36WCIeFq/zrkrCmIP
wpm/jvpznsjlIURVJcCHUD/T9ye+2dYdP8EwLtltpAnbjnIMepZzNurXtGrQhPpo
6HLi7Zx4C79eN15EHG9YQ5SMI71OtXLdlWuxFWf/YxqyCoCRNUgvrypmp8Aa6PRS
15zc4NcEpca3HcXs6dACNklPlMzRZYKvmwgMHp5TQJn6F/y58icqFERnniENpxyx
CwYdwLZHHJSkZBgeAu6IRpwYtgN8s63/u1zjjZTY1ew//ha+G7wIJ1yakmdwHzyA
jf13cNCi/mUgxUP9eQTGmPkOoKJfPPJK4eTWX00bNnoLi9/cO4mniDITvQ8j/jjE
Qt3uPPrk5Urk4ogcQq64MqpDcijQD0HAW7gP7s9co49FuGevY0UYFOnti0ClvFpK
ntFv8tgZuh0AhsCKOgqIqxb1F45o0yWGB7WkQh5g8L20VV9MvgwWfCwk5yPxOgQ5
rTMxnO55e8VWyjFdT3d5Zhxcv0rTQVyxKO3sJjs7+XMCULsdQsf7dY0fG6KTaayW
jBo/cfgDiOnuLWAcEk3TgXbCv9zUtAKt83p7rqvxaKsdXxmM6ltPqzpY39UTJ+Zt
9oFIuxOnx/TH43Ulrnzb+B645sIyXXg1S90pLV2T3ggcsXXwYvakft7KghsZ7Ifn
68Bh6hMa6fnsB2ztMYonT0+YunnEQiLHdFq8a0u/mse02leqVwNvqvecGQEtHIv/
7bW1W5NtVJ1i3SU1honQ+wnwfgLREsgOsYX8m9jPe4FUcxcS2bAlyEtKzi631CEC
0EOdYnzktHaMMIMmlsk9R2fRH7bk6O5qGk5OT33u7pBWQYa+qnRs3WitPTJIn611
kf9hMnh9/r+cejZW9pbFm2sQRek7V3uhzmjGc+HZPT9CwOlSSzJJC9UxPU65h1hP
R0pO4j9kJrdE5Npgf9KwVRJGYZgRDXqJxVbIcWK2gs8di2uV1uyEe3EwaCPeyt0w
6eJqINe511UIu5e/oL3hQIq/6J24RmIX2muLmzweaUHYjQ/NT8UstFENiQNGIHZ/
3+EIEQI/a9FAoyvSGN64Vay69eeOWUnwiMFP5tc5cTtwHGM+40NQEdLnPuICa+SP
wlWSvG3FUW3BYUcCk3PpvBi8K7MA/1CZu1wB2F4ibe1pmWqDWnigXkqdSkOM5+ui
71PtbTXO5mln9gN7zC1l24hIpLXVWqez/4X8n7sNzAglWJp3FnQSfHogRTHToHfy
8Xq4Pcvb11rJCcijPwtQfsiRTqYnLVpIcxA00dnfrY2TagpTsriLrz3f5cfaOI0y
7rz2kk9ispX0L2myY+G6BmVxMDAQZFvvie2WafkVzm1R3Y98UMts71w0VWoY1LCi
fUSRsn1RJ8zoKnnlEvxOF2XUNvI+SxdIFtiOOxs0k+d0HhmtE/DEQ3n/UKMIkywX
C/ZtgiHayfb2Rn48gX58qB/y7dw1iwgtOvWT1doRlUCIxLdkUvtaLDj72qouuUCE
KW51ZvJOHxL3xYihhk8Trb3crk6SAywTErVKvbK0c/XJQ7B923jK9mfymmV6gFoE
EvssYyGd7jioyqQhvJZH+yPM2NAeNQoqfP9gHPRrKxTeYEN266Xvha0QAdwGrpoq
8ZwTaMhMFsyt7CxHkAXGVsAnEylKPVSqUBICoeyC6NbRZkNP7dtZ/RubBJE8MdS1
8V3znF64+rmF2Kj9r6XFaawLgh5VkzJ5OWVRIzZ683f00ZNFHjQBo3p9o1KGqum8
eNoh2SiatFSt6Y/+bHXeupBglDePlw0QkoW8QaOdi6UKQK/Lxq2Nxok8z9pfX8a/
pWsxrKYgQYJwtlZ9cS0863mmsBfyf9m2PZcnhiH0sjJ0e9Olhec3bqEpQHSB5gCk
x8jl+TpubIoqg7vcrVpzYtRtnlm2mHcj0VupG4IpM0puyFJnEbSvGpOE0fZJS4Uk
TamKQ63vRo8dE1Y25cnlO/5b42SKwdcdIBiYjVQTiZT3jvvSTlRzQUONnDIutaaQ
VEl/9GkBHOFiCuS/8FuYXUnJ9oYqLiXctNzcUhCOWFfuTV7+PtfVv2EMBEpFh7VH
SOZdZl3nAtMGTTYUcQeraAqfw1nzOxwn27R3bbLzvlbtnJhgQUeMrxg6+SojAraP
4m2GOFoSv+MqoQPlh4SiuH1lQa+n80WrI4CsuOndKDR4rD9jtIzMkGWRFLgInBlc
Rs0FmsXf1gg2upBN0mU+ytMkDzY4kRpEjUydGnlc6K5qw+C+mTL/vauTcGsSXLRp
GwqsqoUc/YkFlvcDUwjJf7DpvpQrsKtY7kEGmavAq96yYA3vNw+9NzDCTQdyHFDP
5YLUsoMaP2PlXcEtmJ0rV6HVK0sPmVXzsQfKEDocTGfbMp9nclZW7MybxEQ85w21
uZz713crO+J0iBwPOHUSVIf6CX/JGyV3Suati1nmID86gweMw9gQlyjJuO+pOrhP
wM9teq7dR0ntesRTOOQzuPOKEKFRZ5s3KVsN1YryoY6TmEQhCkZxOWaBoWBRT4GK
4AxE/onySa+A7WHeAo23iZ8e19OhCAnw8rvrXi7RwlJFX/HZwjR2AiSS+5fH/zI3
agqYg/cjnCV1tutDxw2nB/ZBHLfRsE21ZmNfGV9Xep8KGxSmerrPob4MZHOl/R7i
Gq757ck9MhNgZyeWUtm865NlxDprnjakH2InCqRFKY6FmPqJCuyPHVw15Bg+Rw1L
eQMgZGfoz3EvkgZIkb/69fQtRdbimjUY+kggqRDO7o+5JudwW8bUDiyeqLPOTxvq
Yap67Ts2FKkmd8fC8WwihoFkR/EO8LFQSnTDvNfuk3NfKLchrXpnr4YUWsal2GZP
S7UDtedPkCjhxK93amRY8ymawLSGgcQi3Owh23llw99SsKhnv7EUdPUZXQmxHO/y
sCzNYtLWCF37pRt48QWUUhhH+SSG73MD4QeVaXyaWOzYxGHCkf1Lk0CCQ2zEBABN
bLB9q7Iqsa4hAxDooZFPDg1ESf64YIASNbnLQ8ZtrjMBPUG9L84Nk2aO1zoN6lpI
AdHgZbsqkfv5EB/WPUsR9F+m0C1xFqgmzPfEpEeu+35W/5HToGoSoJuVheBlza+w
vyeTxGcaJYLuPpA3yk0IDIWlj6ARLhU4qdqZDbouNw+BI0YeiXodzmkCyMCDg0Hc
LUK+kcbGjSD2XzPFqU04SV7oEwQzsKGteQRi1TPpPBexcezDkZ1kRWWpnlru2bFp
GaaxpUpGcmpLIRiSLWEtGJCqRVTN12NM6nETQRcSNJHOqADjKEGbJj3VJj0oPNSn
TSP+Gzzi2aIxFEw0OiHFkvLxCFFW+qeeKMbBGHcOhHd3Bz/81Fq3Ypj5iwC4MKd8
yWsDFekDdS5t8GreSyn4gdDUVbXQBnxPHZ6fjq2uDI1A/Uz+2yWw5DThK9jPBVbW
GQWV4xH7jWBPGGe5ErpruMb0cxQd2xvVGLj0Z46lSHv8uNohT/PTah98WN3jHGpm
W6/j5DPTy+IgHBHs8A3YdQXtTA7CAp2xr/FoXdT+vL9vHS6yEpJC/Hgw6Rb0apBW
5XnRLZxvc60Gv3Ld7KPD8R90r1wQJrNXdk8zlHFqf6xyfcM/dOgRDP044Gjp842T
ieAx+UavaeH0Fx0R6tXc43Zhya/0b1rgPFL4YdQxmbN1dDRkaFtYm5LLzkyKkyZy
cjrlIr7CiauCdP0ckOlEulT7qHfZLkWC0Ow/kkmAEVzPcu88e2P0wbvqadbRC7r0
MML3xYaX1JRB8s2M/h0BXofyiRZMjfNmAoFbasWDhlW2XfqH2YY8zOgF5WBtlkcx
LKssc26Y4K/7zxiRJxZTrTuq50pwbtjOG0Ui/rvyj5pliLDVkbFL+QtO6t3e2tAw
8cQY6dNcU3+qX55KMkdMz6NWtlCASueYtrv98G8wgxYZ5rwgOYfElxRhyU6e+FRl
nxrxZrVutwZWLVRJZpXepmN6hnU66J1n56N4ZKp8BbTF9nvZfdVeKRlDZdtkieTB
Y3YldEX5nSabmnTvcahPap/EEmaPvqrALijllLF5WTFOiOEi/qx4LZjrA65Htx5d
vKFFmdYiDK8k8AG13w4MR+HuQmpoqpErql8wh1fp91Izwa799D5ZY8DJ/Qb3rgmk
0PaIZRMTfzZkmiXSR036Lj6aDAwHER5ZlwfzZglABK1xIPYGx5Q/BzySr1u0XVoQ
hFUlc1V/lh3yerlLHFeyH45vQP3gFkdB7N7sfqmQDMow1RI/F1eXFYZDg2UbSRRq
mK8gZbc5iHh0SZJVNdDM4/PqDGU1HbYX1b8cuPVNEXl6ZxWDVD5ZH+7gtb7zSy7r
6rk78YsBbiWv5Zi2TsrRiXk9A5z3DLqVfNy7tRek84GyerpnBJGp+mYVbmviKMdj
PVDBQEi8U3DNaI53mygKWekesXFm+k1gN57jlbxScs8sChgpHRyHKuL8K6JNA+fu
Syl0pOZ9bXG1z3yYSwDKFwFhBYTJHs4cu/FzvNbcKYW8lGiQAyd5ff9CurTDsnOj
Z+ZGh5WliTumK7vyxIdzVPc7UeKECFc8Q4ykb6DQdFceacWuUPS2cdw5sGO7s5TY
T1m13f7dSQGPLXk3hlp5fwQWlLEI592Q2WLDZhX+WcD2xfDYUBhdMz6ATwuootxN
JUwlCkCJTgsSiy7n5Iu9204tewVYCk2eFChfADikRzRqlvwJKm07VuZxOXiaF6mm
S8TAWLE8oCdA26QgupA1yaN71YXu1jGOVmCbYuTqqJkiWj1SA6d9BjNobobUY9xr
67Qynf8OYWiCkwcGJU+xIKoyOGh8O0/5cWaz7OcPzVQ0YyHTntxFROcGNKJ7vYPp
5im939AA1KeWyaQHd9uKezKEHuIPjqWnlD9r/fYUbVzLapxPCJRQ642CBsoeHehw
yUn5FHEBp4JoWrNn91KH4H0Szor4VR0/Z10U4Yi4RWP9Eq2de0c8g3/kbdsLxMlH
Y6awDQJWmLONYEqcUXmTevzzi7TAd+YQfFi1injrD5aj5r2OLfVsOaycf4zb/JoC
KYwwggiq89Idzf4qREAgv5+437kvhsPWbDRQv6McLYwkxD6n0gEZ6uGA+OOWk+ur
68ojy96CPKShrIe0UMMM2+kJHifVuhv2gONADVrKvtyoQM+6vJBo0AMQ8KQNoPO8
5tIWp0+9LV031WicE40xmAm4OQzmBKWtU2FwKS3ObTYaJvZNSPj9ocue2dBlO8lv
QGmMdrMZrA79sAaP/SMeJ6bcfoCf2QUY06O2XGMZ5EtVy9Uqwiui7L4bkLn7lwgn
vFbzj1n+uCdgKQHC7SmKiwzf7g8oYonzbDTT0jzlk4M5J92/8PTJ6zpDZr9An69p
i2cs3AKrwJZ/W7lTn5bNvdes1b5BoMoIVlOZYEEgde6vavdSP/qPyGbr3IiDtUnX
WLpjPc413JbQrITy+tCqcxoj19FSqRAVb/QKd81teDIkZ1XNOWHYxAdCYCwGu2ND
MAEz1hwlKxdlJrIgIHnjS+BPO2PI/5JqdcofEkhzHriw4QvTYIrDrY+GtvtwSPlC
Z8EFl3fV8nujkykObXASbdn9EExFzPUMxGHHKqRHdBqHoN3wZW4AvakIJzMFRJwp
ZUlQU3JT4qGJ/LTLSGMFXVe86+6MP3za0oQfHvqOlGu1+si1QrwCMaKtHYkr9/HV
riHIO9rz+h2yJEc3WcS7yrUenBWrDU8V8eN3ikzys+m45027aeT5HIHdZx9WZ701
lt/LMhLrbNDny4ao0jiX4zz0nbQiWqiHLQxOh03bW/af8ioirOkCrxEyRNA87DCV
9JEglyZFplZ16Zydf1prupix44seTHvy1ulp9uFV44FqoizZQSK14ReuCL6khzyB
1q0KJLG4cxGgy2HZEriZN0aS2s8jABd36d7tVt/fd4pI7p+PS37TWptC8ypGX8LY
dC7lZbkSdLDi603xxq4rOvXPORgYOxxUweERl5GsQG5ZyH9fw65u3jySI/+86lHA
aeoBDth8i6EuTiHU3+952bXGxInHOpxUPUxWqXi9f502PxikBNmzWEbkRoutt7fA
Cbnnqay72ouiKQaCd/e/d/AZA/OXvpsXPBTGbESRHFfrGP9p8C0fayBLHUL5tCih
sqqHSaGZ3+zrj3GWo4HRS/FM0g26deVdzw/O9KsUrMYZQiLv7/lWm+EZleDSu96/
qXGyP3K0nA6Fb2EeuKJ3z0KvVt4U+8unwi++ar1oIEvXUx1jg8+Yqt8n7il2/N5z
9icEtYDx/QMg810+SFq8cXebA/cyhvPVqsEDzNbNn8YBoBchuUqEWa2X0/KLA5I4
uEMrvnAv/2ldk2c+AL3mOYvK7a+xCCUltN64CFDmmGl/ijODlQSSKnbmaBvoxedy
XtQbtFUdno2YLSlNaAOzkQQoswQoM1ZIBqwpJPhA33Gn9bMo9zkd+LKGIYnUoYTI
YKuMffxPSktgV9z0MprtNnKur25yLBv5oJrjmryxL0ifxaD/mRyquhWOMLUaKBEY
I0PoDEAW7iXH216TJFGwriY0xF0pb9XwbAPVpkHXNH7bez+wLsGZ+TUHBns7dF2T
mOyaOIs5eS2ladnj7ODSulycgHSCmVLjgiNwe/tYmScxYDH+kMgmh/ixy3CYmin4
rTwmsLTiQ3PvhcpAPdy7GRJ+mhVeIiXGL/5Lpi1Ih6vzqpsGot5Uhl6tzt1k79WU
Z8fwe6xjkWR7YFo+bfJX5R9sQZltAVNw3n8iWSg27lyHosGDR4PEh453m2j2hxSI
zyAPOO+jYXilAS/bzyy7oeiNHlwjBXTs0VJ3f6j8MrBuTDRRTq00uk3z/BN9rtC2
y7du8fpjCpjkWy9mqFyOmmnUYSeZfWJaktY8ApaheGP6NGvheWCy2VsvmG0aaOY3
lX6QcbydSMqYA4DtbXnHEckClcnajDvFUjYkY03LdfP/YBKjdzDssKd1jSO6lzL6
t6y4FtAqWXwfY9hrP+gqLP6pBNtxoGompBBLvyCF0J4JrPygpvu9DKt/269jiVzO
AjwrvC7tGQiQBESWt5j1zclaUx7oR63I4Bo4broryYe07EZYlVfE7iC6lY3TDvy3
Gbf651IZJmmYBjAmeF31LraO+qZ6ngxx5OxbYaCtPRVJmu5x6jbLH8yyKntPqE8J
eChsKsGQ+r8n11jtYdG5oTURrmTMaQ9j2TNL98ucahfI4C/xTpGHBNMTw5ifS/ir
AzGx8gvciH3Er0QFSlPjpbbg0scM1b/49HkzdbxmrXjmppg0q9SzgQaXN5z7GMua
1FZiRIGVS3eE1hXi+iAfO1AoVPWgTpW0POwzwGBjaZv2MYSpIGC9XX3RXQ68AIKH
iCiU0PFO4NDvEkrDxDCGO2YFBeT4w7smZ8D1LmUOyvGPId/Qi/4GdhJ6ZNzRVRkp
ludFRjyM6mKmxNp+LnhrLdTHycw8qmwqBS5j/mEJPHbO8V7hOV3eB50CKl3qQS4F
AKgXRamj3PMK2Ewp/40hBpAEEocjzYaLlwj+47ZGKzYgj2wr7Y/656g2A+yhQVOx
31pNQPU1g1MDAOJH+2L9ArcSJnoLnMXibnaXzx40FTr9tGkCBOO17obcf8raVOVF
AWkduLit0NY+O8k8OKq0XpWdAFwcKN8oCdOJ0XYDiIsQXegKbHzFCXDRtiRxIwfH
2rImvZWZJlPbyjCkp6zEq1JhWuel0hYjYC5ue+3wsQ+u5sejcDYc8sDboYM9tWu+
42G4blatG8dBD45/SjZW8egJSjPYQ/PRTItPvb2x7XzmEOQTGFYurw6RatfYMuHQ
fdxvQser27y7cS4pAgMy/9NGyzRdNMlcEg3HuZJXMbRoQPGHBWQFTBCDuSbL137M
pzxay492hdClIMrG9iwCvYPC3DC63DDjFlzxRgwh5s6ckqLMEGAUeO8Jepy0r5UD
Urp5C46KwjmM8p7M+mqI3fUPQjM2NF65OdbILnZputxEzmNkGb2XMWRYhTEnYhj9
tH3bbX+vtJ8H/erQrDDRe6TDx49C/uIaDT6oaDYyO4jSqbTbV3XU0SescoN4RR7P
Qm53/un5OTg7DJMRybCgLBDSKRxoQ+yNlQrDge+Sm661/DcXoIfI0kPXraY0Xyrj
0eY7d7mOOQZhp39sxhfl8R/VT3HwxgD4cxf5i7yei3vPRULAmfdqThor/AqyD8JJ
uCa0bN6rJAMGkzLfbvdiNeUDDWi9O9tBS5G4bHYS/cMwZA+s4csC+ULVb5yeHSLl
ixKXRRpkZw9471wrLmDgz6CK7gRfMbRKbNntvoSgtaAcUxmoz4QUGY7g/BtPXJqo
yDLg6RZY7O6ww3DH+wxIt82pPCbPiNuBSgwb6J7nAgd3fPixunLLwfoKImldbaAx
CwMdPZ0slE2trX0fcSmgABwT8TG92YaShj2nChXCkCa2n2T2R9uhO4DIG/zWHFBM
lmzv2h+bfLg1ICuP9ez/SUT2VlcQ8FhwIa1NIQrchP4lLD5WnqQkFcrVPyFhalFd
TZtpPXqtgXnEaWlwbJwPhEjJdADN9xZgywXuWlaNPVj7RgU7Fxs51NFNNRS/cti8
p88PGxZTArIKaLi/r829TdZl2fTfNpvsYJXbieIAE/knGLpDSuQ1st5sFhRkq6r7
VVU38dWb9B7f2q0sQ/4nHuUzQUPB3KWvgxCIUlc25QnI5Sdm95PdNaYFLeaZ/QVk
zn7SaUArImS4jD3MJvTU9lh6/OMJ2AmTwYYsnj/UgiAnpfmMDmgssUMm+N32IvKM
lexS0B1zL7tPrb4UmjBKO35HWRWOlXrKIqDjyTMy6H7bKB2e205DLDqgnkMlEojC
5uDtqWjMBzbPN/h7W8MY4+FISCfH8akK/n2DLKXFt+EjjqJCt4KtqBXvDsp9wsVD
1Hot7gWQZOoMwjU/9xt+rad7Id0woD4C5beq54kKxS/lfoIByn3D+4JPUqwiVbNf
0C/Sgilw/FBVv+KccCNzkfHFz1Ux9tTYnQhdzqEZ+PWB5xKfme9Kq38zSP/iw6Rl
IIV0MDETv29Dyu1ZUJtOpbsfV0hEaqcTs4RrCmAJAMLHskjTFcZSIsNhSvEITHu6
aYKM5PMRaG1+fbbhLXH+jEBpjFAVuZn/OExJD26x6wBH2zRWQRmxfCg3+p1pGuHy
AUrN4wn5yY+uAuipcewlXTEV0kFpNOlpO2cqo+NOFAXg8I7WM6+uYCiMr3jdP4Ek
RrO+22wgl3iLGmZY/U3Z4CvbFq0wWgzIPPnhKcVO+6X9zkcQGoQWA5NA85WmdcJc
zvv0vAzEkW+9QB4De/WXXwJPCabXB7SAhq2lp1+pQS3Gr2ov7naI7ai9HA3djsks
BY8H4nWJVzoYi6o3q+NySrp0ygTzVf5LOLepQOnOXOsch/aOg+dAiNBnntuDTDls
oXymxTJKC7FjVJs+/UvoVgskwA/PIFF413htIhUENgCuVADGM09GAcDsDTBiDXaq
lDVjgXNULONurRvJaM7IEtd+ghBCEkSgrbbBcaqeNNKFJjDpT12uLLvAiyjbTXDW
2057b67MD7GrcXLgwJUNQ54MWcZgEh2/v+Qsf8aT7KpSMOqKVN6ufrgOCOG2cgV7
jvncIoHb5oHVa0rNwZ4zUdgpzaFTliTCfMAgUn6wVyfeVwEhZFdrsHZTwhQs5whM
Ph7PhWmGmmM18dA5Ok4yzuZ1M+cUh8mvVpr0ucmbUABQgqAKp9mXz3akEz8YuXHV
OS1UIatcaTJxAkV+FFv31CtvdQwSFdItKoHDU1H44xAQTw/C+nnkdLxpWA315zE3
aCgyKOm9Hs5nIVGAbTYNO/5QGzK98E4Nt4GH6oVqXRkNmt5SKedFXLbBvv3Z4yNO
F1a4IElUT41V37jxHFiT4zs4eDjJ3iYFyNFGeJ3dl1MzPpRqZaVZly4hhOINZ9a2
oldDhtSVuIKZpmajzGngVhg5IdAOtoxYd5esW8DJft+aiaNDEixrv8dWDf1TyMdd
PTmuaCSIR+FrkvffXDHEHywoSa51okAwKatrkl/xuCzZ0nM7P5scUWgo/tqjAo/G
QzThS/gSPSsElUIeiotX8TAuEG8c6amSBqKyZK45ai3fMigEV2kOLoht7/edG58I
QoUIe0DpgQnaFRa06vhwxsW5xqm7vNg6tiQlJf9YAGE1znoA6iHXnU7EY6YvVV8e
dW/x5Dydo5PTUovEWYiUYfbnbA3shiyAq/91sFrhvQ1TNXNRq39WXno4ruXktmdw
hcoVJVZYLXbjxqZEjX/a8xxTYty/phOHDJF7OrbBsQoR8U3ma6oRgfGNeBdJsgGP
YBpeKWo0vklRVlMBzzbDH2P8QAZcWBfaoe46x2YrqtPrThZ78rL6OmdVLamoB9aV
NqH2Z88qK390aSPsOL1WOR3ioROftEuF6dliikd/tvrHJcHffbAoSK9MFJlPHY44
q5a9TQR3/IjQgJY1hPMvg0YdLQgg8gGY7e9Dheh45wVYo3EaIwzs1zhBxtymMpz/
hCIZxUU5lonP8OVeVYtGQm0M/P1TLqXnTbEhZ0Pk5MQjpLqxKY1UeJl3UtupRtpL
lZoFSquVeQsNbMbHNxFeD0/1Mt8uPGUUohu8ViJoFrsNz2U4gaMRY1LqLS4s9J+J
4hoqhOn7ZoLDotWOd0RRI4PK19IEhZ9pwK4N6sAstG3Fa7I6vNpIzSYcqjLIpjdC
iMN84XdIB75GSWcwDfjvmmZLhsW7cK7ltwfTyL5a2DIseSlsYI/h0mt36Dn2UBLJ
4lcs+3zmVHwcrNFHTRYeUBQg2NytNkcJmd2n6+B/jxcVtUCz0L15o2+JnL0N1fFD
QKFoNqwKNSW6A4NK1K4j5BxNQpt7jvAQMiusMEzqa8lk0KlKF8eEbsM3hHp9WNCJ
2vb2c6ToB1vjE4v+5QciOjme1QOFLrXMUwdMnTqAROwKBlE5eieMlG9BoYDjFprs
fvdMjmx6Jvx3Kd6F3HIBjqH8hCKRHy+2dtsFJtiATVK3wDEjp405Mi6+xVL1gLc+
ovaCvzUKu8wEXUtGswlxWNZNftiNvpv2p0cVIAi30OhzjT1oZfDmMawCYEZO32ud
f+659ZflFXK1kzRzhUeLhlMXPQVJxR8NPK9yTTXBzZjH+B7AcE0T4u1KT2TE0E8R
sfh4CAT9B5eF6SZI1fbU4G8YOLKPHN8ivFn6GxqUGL6TVZMOSMb2E2XORsf+pT92
WsWx1tV5N1tmwANcQ4ebboVcf+A2IU3uw06tDvSV55+DBPHxicmz/YREdhYUjPMG
BMYJp7epkiXxum0RpJhAIgze+lCEIXpbOmSqMsDTm8hc1A09m5OhBs99hKO9BM6B
Nf/QCbhmDPsxHLDoiKimKR4Ypk2EwiN/UQTx2TREfQcbatQ3eVPhJygELPcEBOhr
ZPSsAEzdnL2dGf8wa2sCIxDBftTyqwZAMGXtpSEyhbMmq+Q2l1XZB7W9qsiGYu+X
6RBP4XNo1XA/3jaNOT3C3YqWa3jJIKZ+j1lZFuCYNosyky4Tb0j7qffLJPdfToi9
ZOHHJITbB9oD2fRhCP9sgJffYdqmV8UKOxoejBkIXPSoJt9pQWx4WSoTcxvXk0fn
nHjfDVsoiyY74gEreVaYvJHkxkNGX2s7VEuYbGDAU+FoCm4NgtukRuya1iJDHAqM
iDoUf8VoUQnqiwXs3qDhQNc2HfAOJNM/OKaIkODasgUteiE2sTvDm5kkNbk+qqqA
BHVI5+yhm5RCENTSIlU+oygKF5TeZAxi/5v4RabShjhqJYEybFGqXbEr/Cv1sCDd
dkgsJ7b4BMSt2pRD9OL2IwqTFMNjMWUKPfNFMal4YpjdgxJfwPDhIxgI0nLRWspD
EWUbtg9ulPbte/NWmmBJ34507TT5jcC7gmMdpLcHINVnhN84hjHiVVCabCGnnIJF
kVEHML8n0BCLmmHomfN39ghO/iQ6Zr641afjvoYQg9j0axdp22/CAPQCKYAtiVw1
kkuR2PRvRZLutJRkMOmdqoq9tvqmruGzrTrS4TPYfNQ6GKOBfovH/9fMvVIuMSMG
6MUjTUoYvKY5ispuiwQhyujLe7RN8H4vmEMs5kUTEdnejbbLDMjviKNOMrUQIelP
aG/extE0kvassMIN19Ou2vlo6r9rUX+O3tEuyiMYn2KWWsr6Gl06ZGzWKH7YU+1T
VJpmvB9OpkAO4brCx5lFLYr7jjZsRcjCa55/ZMbiqudlxLF0S+KEPY9AXQf+lv8d
3lrHshW3Wc+4HebCtPAKhXc7SiB0rbL/b+NNM6+WYhPKNYygmU/Di74zIRBi0clS
8MiQ7m3lgo0wCaGSkoOb/jK1UnBPBKthbgp9UPdyQYBNhRChTTCQ/FuUJXISSU3H
MueWZh/YzuMWLD6dQCGrXdur4Xkddh7JhKDXa8MGdzhLxxnGSx00ODl6SimxIR0h
nNMSL+D6Co0IBpdgR7PXfwledcFFFSp6kFGqnOTqzplYq8CvcsOWaYO4VXY0pPhI
q/XNYv6ct6JCVRWeorfh4+T5p24tg/CiFulGOtNMGiaDon04oQPg3/a2Plldbn1x
KsQHSwdUY8yTr+sIRu+tmp13fu10BuceDIWhUVU98kPsNda0wsPCWdMT/zFuDPfV
bxI4KpOPmrsav4u2TbC81TKC6NidIPY/Zn5s/5zQCzuGJaPIvihA32IZZapsWGOr
DFBH5vUy+mADQP2E0oNawFZ9J+XSv009c2L70EZIHksXQqkBaJSUME9JsAUzftOv
Taon8yU5gl8RWq5oi9NB4bCuIpPjVMkdIfumgg/A9GzxQKQE8c7YFZYi8v0AXCyZ
YQmkxadYZOLYaQoIt1tQX+qkFG59TKq59rR7638cGiOdT/YZYT1E1jbDNqVqpdH7
u1vPaiELJBqLl1euEWxt3l+WsDKoucEfLvv5MK2RCfIRu7pR7WN/M9oKKTcO4ad3
t/MwC5Wwz8VwrwxkylF3jwXTMoIwof/niRH1iqe8qUnntT11AMhILEFTVoRCIRR+
Lg6eHBOCALw8oFN3iVajVDIhUVs2uOx0BQxC4HhYATjhhgUAB224iOGwRz+smOC+
KfgcKHfi98joB537dzrCm6+ZG0kQsLAmp55jsdcL2yKE9C0rC6dbQtU8dfdHx8cd
XXl7GrJFq0YqfFZKcoWkEfblzHCmUtS4ClRU9pbecRLc30HDNui1dtXS5SSsy9TN
lJV4ZR1Q0tx4tEvCXr296aCucCbeFu7VlLYHDAc8g8iEAtFsY81iqjQAR1Vzm0H/
dA0PTpX2U7W/+7OP3dtV7m9ZjA1bl5PCqhrqmPADLH4LkCgITEYCBhptwHvvKJru
5FlIfdn8nthEHIr59dCSC0cwN8RrF7IBnL3WNzKemXVcFDT3h1L5tWkAbY5PL4/c
vzl6LmdMxJsLGFajE4WX5yfCcXvb2AlIsGnZbs1VIKnejoo9BBkXaJ++tugEXjr9
9itiZ7BwMA62uAmUq2SjT9bzzFy2DANABG3pZb1Agdh0WCM/TMZQ8Of29+/Ok23X
4eR2y4vGjxAYyDw+Imk3nwr1R+CxQwU1v+LHEowJZzte65kFL0H+7o8gdIiAz7l0
VAn2Cv1sGNWi7AG1LQ6GfrxhuEbAy7epVtItFRBIp8nF/4fdjWFm2EW2peyfSeqJ
Fm+AMSW6t/e8E3DA3WGT91bZ3O2RAUWMRXhqSsd6YrWcl3QPXHQq0cTZNP8sUHzm
5Qh+DloylIwbw1kTJ1PFxb1mpnCQ4OaVbIzGSVtbSxMyrOlSEb8PLnRLxpJCu/PB
Rrk59tyWPlF7AFlY4jNsl2On+5qDfEay9FPN2l+t3Rep3g05g6s5OOUxM9HoWwmS
g4ynIxDcU/sTs0xUp57Hs16DD2egrJdY6MuIfbpYoyRMm4YUHQd0G2Hskt7Wljge
eLw3GfsY6OMWdp2nf9IqruXUg914fu6DJmkaelHAvBLnjr9ymH2XAocuKe1nol2b
icdq2uzaeivHV2G08et3RS0EN6INEa1Yyhl4zU3ndBYcVdc+dqMba2mLIf/iEVCs
iimKMZqK/MupDZBZwq0/6GvMkxDVF20y3YVmcDFR/+62qDTYH8dkao57fHXx67U+
K9cWrWE5TT6wKXwBE35Pz3JO6flq75SOORwlmGt3vmKNTdMBvJUMD5jEwWvCIUPG
Cm3KubmjDgqygnMxaVd+mmpw1OxJIAKG3oI2xlX/W4YCms5TdL7HSgbxq3W0rsvm
izbYz02pbQNPp8Czuhu8YjzAScRdHOOhVmW58ZZ8XNHvYmybOtWe6QiUOFwi2HGq
MRc7O3xtmSuH66YThtdfI1EWZVrJ7jJ9fIdYDY7VooTtRmMtAfZixjS0g+wSs7O1
2CGw+sCkvByUptVF3CaGyH/n/lPWo5VtOj5wUu7EpSF69HNxce3Ui6xeb8zhHB7q
wWEXC4FZtXqDHLYjpWG54qHWmCd5wnC/4p+8TnwyO40RI+dbaQFonDYhGydFlL9T
RlFFHUnfcbz8lEl2kfvJDhbir1kD18a/co3RMkp0p+LZPKk7bDylav8onSJe3Vx/
NE1p/uz61Q/MCkB1YyyX88tACBEZi99jlglw95RLNUtGIvJc/0lBN8L0jd36GS/p
DSVeFl/wJAIwkJvtZCoTyetRe9fqr99aIEVg5JnYU2rsT85yix/pZEMap4h+qQHT
C8BbIqiCsH/Dmgw7AW40rHCqPCR4wv8UPjGr0e02K2SYl+wvBALD9Jx8b1Frcxbn
luaTjR/8i1AIBHlYqMgEuxU5mhvwzs4a9uE8e+q96k9Mc6BI9hWl68g90xGmZo3t
+L0YSbVuFhDOQY1ZGPHrhrsVYELynH0IwxXD/LoLYtKWhHxv1UVbHV748o6icS+r
yQDjw8arOoGOtkYXjXzpKl7hslodfnoXycpIpg32tY/vTgiOMEkccoFFWJG7XdYE
79HvssLRht0QWwM/SushAuYADHvJrHbKr7CatP3fBfviakFMJYspMnU6iLwf3ABD
wqhIM6IqEDdCeY2Ra9/WdpTLNxU5pZgKAP/hZC0bS/asquext20/KPN2BZC57Oyt
m1xKffk7/XETZkTvwr8HVnR1bweg11Y7C9iInuMMl+YYyODCQ14XXRGs+425Z/RC
WELDUXODj8iPOYAstUjTmcdtommTGXKdRSNaMJuWPwacDeMyVnvxmSIsVtegtDgI
0Qe2Rwvw2/YuyfrFXRaJOZofdML0fRmx4RNwLYfXZRHUSItCCtof1Pw16GQin859
YiflPnf9SM/1nLFZEDzDNxotaks3PUNhayp4ogLpNx4ReVgBEjn3xakooo3kKzJn
cGxza1f43D48aLN4v0raGT+RWlx1MbIi7smPyfocFdPdeU6Dm0GDgFuhgK3qjuRK
Y1xU1qP1c0GlF8eDV8N0tGvDE9ukMHkIbLv0j7mXJlsX3IES8jsec47wdAhyf7KM
WstI7D03+glb5mmu3Kf05veMd+7YgBLZPDd5c2ZZeqAfHLRYiX+PQJluM9Yp+WUu
+VoNBHYrz/Z3olrmXInzc4swFIXBHm1EhFvOF0QTa9EDhQkvbwu9Tkcyl4TAl7R6
/cxk947HoPyshETycrnw8Ic6+5++twWJBF696k1vYF2U4hXN0678VNkhgz89rNYI
MlkqVZPShx0pp8p0eZ75dOG/8xuy5K2oyu3zOdBsq70+v58pgmvkI/wlL1v0CC51
rh9vX8/IUDZ3d7uuKBaatpLohQasg6iXb0NqmkB2lmimoAdES8LeuzQ81gZlqexh
B0qm0LzES2c15PWHLVxt/h1P/B9ru37gDxGYH80GmtJ2ZT1RmUt3RPYFvqi9YMW9
V1YsCtZ4YH5XU64NH5K8MAL9ji3s92jAJnn4kAQUjJmtnCD4kwQXGkPGu2acVs38
H/j1YhWKXnuE0nxY1cTDXOsA1cXKrd+SKWnT3Cinoro5zW2goROItZGAfTQ4inmX
KJKkXsl7MTJ0B+iFTLVGdwLgUCibiIBG6m4aNtRjCjK6TjQiehwQuB7WktxP8OVM
rY7ccqIWW5URKZR1P9BKCuq+UgFSZJzICHjF1FEyabqc1U91qCVEmdJV4ZHJroh7
S+QJ4bev282bhnYGMzvOitisUhJbp+MWqOj5MbzJ/zSK2GH37oAE5p28Uo0qdpv8
Z11artbbUjItlvuFm0DEgLDGGPMSv1OiWlf2hc63XF9SHg7SVZFeZLjqz8mxo5nY
2f//U+DLB4vcJ4eAPCZ8wBZrNpMlVRosO2nl3kKA6IlKC5v/rHbSrbnT8lpeqGQI
dxzwsYKJcdmWzRmzCyqKVhY+GJbjLQ7JuGNcmoDlKdqu8bXBB6TLO7Tvg/M5FWPZ
MKRDZLJ2lf/S6GZ+5LEZzkOZGJs1ZVG4BPsOKOO1dovCQ7vzIwZZOUz+p7VMDaIg
j32ea2rYaULLY5dmUybcfuP/qXmceCoKhOeK1hwzMzuwzPcQcxF+Q6Goid2fs4Rn
FdxHO79OLes+WenfQz4+hpA+SpENITfEcTeeRjmHrwX0BNm0Rr5bM9iIqVlzSJ49
Zxdf2OJya967sbAfPV4U9SCHbWgSKt2xtGIkURifWF+WRakhGJoizQQN6rlfAY7p
INt28teo/9ZFwOjQ8MIcq/5J+9e2ZOH8yN6Y96/8vLVOcIvj/LRBrRvg2QfLi2uV
OaMYWFCl0e+xs3zfzlBStZ7l8nMuJceSzY1jPMbHi9bjlT/z2mvCIm6vaOz3qDQr
5EXbRaO3jQNbDPfh8eWAKOY1nUrjDLT2vmfasqvH+nicArqjBZ97pHyFGN3jva5P
DQdwaAQnY5orsn6OLiELAJVy12ppnsuHd8gYZXVH3mqBU4qyDInvlQuiRTmpVLYe
pxJiK8XF4GMl8VKppSSMJmAO7CLWFczODMNT7EHGUvW3/0cf3HBX837+3VHM+UIf
11txqoH9Aeohxe2XH9OGmFXHwHLMNWBgqX5rTLsspHO8e/bu/tbm7c4JxQcMuwvf
GRckErxzvVO1m9PS4UW68UJBDjpFDF9c2qN1ehJJA4OITrRkp4OMZuZqcAmCeup+
9/vbBX/ZVqf3mXk/5H9LN6u5icBNDu9v1llCx23fny+hCpNncA/nPhci98sxhTYi
jbKotlMW3vqI6POCjGZlhS5lJyTbNxEZH4b1aSHym9BoSd2I2rqDUZMct71QHLqB
QLcq43WUkpJ65Xi3VHWOd9AEwWqeeprMX6x8+BnezIoAJAh1nnUXAhqaNrbv0CeQ
NMFQafFTGiBZCZJWBvs8km2lQQlx7mQH7MBVNewUS8tdq1mcrEIXqpoWulb8/LP/
A3kqtt4ohtmMEWeju90rBO+71aEh4vyqwJNEHUvzyZkEv/tDR4FwLLHs0b3TMG1e
tj/6VZeT6aPnGI3lzqAWGXEiWfbooAjQhu/BYHNyka4vPCMGY8nQWaSAQlAOyOHn
Sn/ddv8xokSDwk/3bqCnTiIePc/oqZkZG8Ho7fayd8gxvaeu15t/OOWFN2sMy1I6
O0oQoTLMBrUi7CMVJTkVIm/h7l22r36sEd37buZlpbEKkrxidlmxasJgw7p9XIKl
e0FYW5K189gDDo1+YoODpTeSs+63bIR75IF0yzsHpAMflu08zMrHXwtdtzLpNQAc
XtDZK57fj3oCFMVJCDmyqrBFFvLW5FnSmjSrXDubRicvKWnvBAZJ+neBs0VePMWK
G09oN3jG+xdsHIfsngoNqxt3p2pDoXb8NqIyk0UBxaEkvi8npc8EF73Oo3X1/9/Q
SCeDA3U2eniY44uKSDdz0QjiNFoMJ1Vd+TBrQFUARRe3EL4JDvkNz1jkbYa3TSwj
sy5I/Cy7p3TKamKdeA3vkQCMoS3C5pSrF/ajZyXWa0+FKZLGNRGTF9XIwprt2WqN
vPX7GNsrCzSO2buUZC/yYKfleQ3aElA0QlUMSq38RSQpX4HmMOD7wA7YC4O9pTDx
51OdrwRO5vdfcDChjLhEXbEFLGzvnGbEslgaCMMKKfono21a63+ZsRoX4hKw50dI
OI4cMYKZTpeFwkYIRvO5GJWGtS361k0jg2VBizUTolLbQSDNWALBrhcdLsRql0nW
ZdXlMYWwWshkhAXXUztnPXfc2ef5ITvHaw7dTCTWvOUMp9WAdvHZ9XQGQnhcBGMn
sDdhLQO1RVYX6sbmnHYR9wAuFW0+uSSWyojwG2NAni6MjNAhkGz/PjcEK5kOJAJW
mKVx6P0RkNRRFAzzN74c3+lc9sVdAHI4xKRsrlP6f7VLhb8BSFtMISnwErd1scjp
UiaBGY01Q/mkiJli/PnFJ9qnnfrSw4j8sUwWH/qektQzH1eI1r4GivPu6Z5TNkHj
XM+65akRS9n4DhE20ux1uyYaarxiWormFT9ukyyApFjn3jOhfzx+3We8+4jukQBm
QxToeaalnT/YzUvQLaV5zvVBuvsuOuvymQzYtfPtTiZltsfubOt4cSY152PesrER
BC47qAp3VnaIz3v3XogFrvAAxJt1ztgtLYLvF0OAOYA0DC11tBK3ZNPZsELD4e1L
lXP4bi65ILanaAsiY8umQ2z9JfPKVhNEKSjoWz6TFqzWzjV6Uu94pO7RAZLUQ9uC
UyOEI6RlBtNZc0f9tDaVx7c98fiCnH2rLZBwvRIIfMKtPxl5yIj6KzfzxQCNCmRO
E2E7obmYY5aPK6yGiU9PIKDv++z3lCDUdmN0FkOh4soDXnz0a1Eg4sGZrlCPnSsn
BmlckOziStiHtUOEl6tDfXW1+lXJm6PNroApqcZsznRRdevRcLWqFKm4LlLsFjjU
hy9GF28FsbHyGkD44IAM9xCCrNaxifJNbPDY5YthpF6SXEx0edrygjczAAmaeyub
XZ3vv3hSE+q1GWO86j5b4nXTK44fbKVAtsYFmftlGp6bAwvuib4XURsPgoBAjg0E
EzlLpXkIALTs5sTdVsioxPtidKanQGcMG1bRWMGmc8Z5df4Vw8CzkvE6aj1J40fP
MVQmQda2owL//CEXii3RfxbcmhAf/6cptsZFBbF00/FcCdOYIdKbUq5JBPz1HT4j
cYRRF9gLHV60jWe4wxSTZPRG3yH32ulOgznVfkEZ3FEKL8xHN9+PzU/oOZ9NjQX/
68fKUXy99vmn9BaLujhotTS8E0QJhv3Y78UqkfDrCY1hesXr9oA++7IewWzbMmio
CEshw5t4PtGjGiNgFiD8pC8oyVKEJo4pIJR3VG6GOdGlWfx1XHs3EQA0MLVUYo2A
+IISzcowS3ko3hl3VcAFZpGXlCGoaNHWe2kka5wxLZq7iL9GsfmupbZ+e+WQuDgM
L5XozWuRktIpznkQvuwT5Eurzlzbaiz8AZk5NrWn73GDv8LoMFEZVFcTM+vt3T+i
tnxbQInH5A5FcOzL8VgbrICzz1jlaKccS4Ke47iRAXqfFmanxLhrsDhebSk3eXYZ
I52rzTI4dpaJw0Q44HoTVdAlPhyOZKuwenMnZgNWwu/QMTTqgiXc5oSw10DFc74l
yuL6WHAd1muEDBV/PQovNa/GwNUu7tuUmFXXPBwjuMtVRjDrnehuY3AXh/d2lyla
sLLYLvHrVb/40nHPC+SmJqcVQTj7HX8EhYrwvCsHgC4Ovt8N6lDLl2hOuURI8qpK
TTeravzACUTs6hZNzkaKyX3PuTJyVHzVQ0jdZ1h+RdL5+h+7opGm6HsmDaw0RL19
pM7k8tQ5BEei0sYesYeqGF9tMkBtsWLmgSKUaHNy0qFAoDn4mv0ymhiAlb7us+jZ
ZpikQwkUbU8qw0YbZMXXWPRoekbTBiYYFZIYmRxEAaFhwGRa5QodjQTwD3Gt6u8f
sHDWqXni8h27f0/62L3WLARM1+0ve974TygBaG5Wev3CvUIFfJpD7Tbj+28qC8nS
biab8igUHKAqnjHIw915rtwAZb7a1hYXTYa/bXWzRnykzXUbjPedXgCELVriw9Ba
XHgmJi6ALQ99RMTtnJDfdjDdo03P+9QsXNNljcj4jJeG6in29xqNWtTpo/me/M2g
zhmUnLyH5mhEhM+lqsKO/SsiEs0h53WClAZ5I6aFNsK5O8OOAmquRMeniv/BuyqF
KebnSdO+SfM1Ul1U8oY5N4th3RX7ZOEVHAdubhVDfe6rSWy3nCfuh0jBZZf2cyAm
3MQfeXGxgEdVFLtSFvxADjX1ReMb/Z9m6l/EjxhJiAwzSeadSW/rCZXwC9qml7x7
1xtYo1HkNl7Qpxn4KNXd7uGcsrD9FvePm8rsx27woQ81doFeVPJTqOL5G1zZCvm2
TfKbxNMLYxvq19B5K/j5oncNYYzat5/3oQEukCwnCk6Osbs1/1Q8mVNU7ey8+pba
OqizHGrtvyCYcOX5Ky929PSkBUc0/ol2fUNJos/u37/nLnmXfWW111gue98czy6Y
82kQDjX59XWiU8xhsgwd+489cRU+o93mzmD4H8H6u5Y8/v7qeaAPElWlL6hKl30G
dNDnWq3mR1V7unrbqMmwQJCu17W2wkjXpfxkJ5Pmscv6eh5EPLe4gIUVXxXX0EXz
oM8CMKMrHc73cMu8jOeBl8cYoKPvaJgR0fEtCbiWFqxrjju4y6H4jMjCzmAN6FMY
kKeb5gcGwkB24sMj3I8WhzKYCb/t6WDxVLKUnWKGk5yC7ZzBzdFyjHWBm+luR216
/soZAU9aUs8Vi9yGvBUtrWUc9YO+LxhuArJELj07OKTsWOCMc/3cGv8RukaGuchS
CRXJJTpcJdfzXmrq4h68LCNm69FJe2ymLi/KakVDDKBbMjxUu/bqMOQZ4qfW9oFn
E+tPJnDfFVXHk6Wbuyf8NGG38D/JmcMVFXF9Mi0nYCOd1zLD9+vLztnP0OlR0hdf
OthPtVSjOek4dPtcIRxpIUGXCcvj1Q0BI3dQKDpfMvBo2l/eHnqwjDHMXgCzDyrD
a2z3+4OCt4pdj2Gv8kqCNwB+qCtE0QFnPRnllARo4jGytpkJKpDHHb8ejwCvqq9J
4/2dsjhvWI71GWh/Xt+6LgLpDeSiDP/MtdHdmOYKlL12rI37FKzGoYYOfMuwKgRJ
JmGQazTvMv5jqqTbsDZlTaiZJP7tr4SMbH9KTunzxZTxm/YL51ezhvYKUedMk3rU
LRnmGkO2jwBNnO7nIf2OhkyAG7T0Ju51Pm8N60V3gwHLNpGRAar64m5xUDkZKrL9
2qo2FPxP6mGXAYkhouP03qa9StMjuKfTs77vFYY9SHscgq9Kd1pBoXgWzIazXYgg
TNg9eAY46N12XruaGvdXQchkUMBMYYwVWb0xcZegyY9iThfNZjgso2l3u/8bSofg
XivbaMo2PUJ8e8FaT9BKkrQ4vlYT1olAf9ct6F7/UO8XlXOAWUQCaa4UoFAT+ICu
2j/gW3WONowsOFOO1rA63f82biRLKOvMj5Ee6QZENLeaPDdtlvPIHCznFBZK/l0g
JD1GQWObN72EUgzJgKknp7i0L4hzyQfFIRYwV+uPQ585LthbesncrOtsRQ6XbRuY
pqpVAznHPvxoIQl8sefNLF9tRbAjBJfSz031Qw/nOBvApO/yQG4gRPU79pSwgbj8
gUPneW/reDLTt/6nFb1PyYDkzNPU00LOo8gd/CayC80TK7jUEuUFqMTgMceNlHLI
Y/Z5d/LARcnphhsINOmERf8tNOT76sFAM1dSRM3lviIhlTfagHni4YoX/Ki48bme
l2vjS0K5BFXWRf7ABedAbuK9yJUk5cYw4xR+mySAKIwWInR1OIo/C8bOzXajCG0P
HUEzPETFFOWxtFFc7W+Y2qjip26wChCP0sh0aFVKZbSS8vQfNbi0RG99jIlMbXrA
OswIsSkGorOqLuj0QcvBIh933JMIFAC/v7m1g5wv+nq601uZX+HGoJMlOKvqSsq/
iFMTVcExN9nn1MlQWZMIqIOXPDxODnrfm4vPWg5NKAh5olAieFHSNPZMSscOuAro
E1mwM0LEnH23q9j+P3foRqpGwEOKfGGAfhtucanI4WHj5EPrqSI3OtSruLBAYuOc
k8IEz51Y8gVPN3vR+uyDZFzO2RkxyQ/vrQvcwXYoVM8z8IOt5BshPMBv/BLdjEmA
PnBhkwC9g8TpsV21h4efC4NKvyp5usU9mF4L3CiYPVZBg5wqZdfdgdTi7Ja2imUl
fU80JRBcUabIENy+niCWkjFZRVQltHGRbsf62DzXVtfCxW2MlFFOYwCoig2r1Fhz
T9mRQTYpuIMMM2ODiKsJH5VC4araTxtxARjLQk050McUwo6uj2GmNq8OaPNUbF0m
rR+C9ZqOs2psmYKoU4L7HV8QuQvWA4NmpFzhGBNQ708gtEG9krB5iAVgLIDhERrJ
IHW4mFqkJ4f/BN0O4Qf3te1k3SbJSW1mUJLSOKsuAok+MZLZHnYAJEtJXTCz+z83
ScBhXE3s1vXZYuWFIdJeQxjNkaUezDjXHh9p8DiicrLIGU7JKAeqxA7DfwVccYA0
nWi0ErK+hPeWo8W/NLbc9m+vT9gHWAuryDd6MU2jJkPmxGCw9CkFKHHP18MrIVv6
F9c6SqajMCsWHGpov7vytt05xQ4Iiki+HrI5DikIivaGTwc0zGmWqDLHnL/LDicM
4AWmlZNiYoytfevLL5V0Rfdv5jMk6jZ2p/WZ5uXR9QrPG35u/pqvJrHfAlP8Go6j
3HrEWIETHMZcOgUfBY93GstmXItbDfPqPIGJhcaPGIJbF6I7hsl00vSSs2/KDJKG
NOYbDqW4sb8miNZeHoLCkaHO0yhbL3gJ0pJ4RvADZGwH0zNJYHYXDuXVt8bJQ5eL
BciFeXAKN0TGQtAuO4ZHknv2XL3V4SEYRMlzOajYzM+r93+XCbQ3MS8GsYVl+sS5
jP+LzH/RYRYgJl5mNkD2Swd7TmZDjJajt8oiJMhPfROMYjSe5tdWAQ8H+6wJleOw
Jiy07+FvpBdlZvjKgjHP+yN1p2oe9A4GZQtRU+ZysyHM6p5b5Ee/NkqYomusa5D6
kgHl63f9W6zZcI40OdSKdkiWgX/LY0QES+VtPsyX0HKSaqNy/bmFM8uQ+lsEpm84
jINmEKmZ5vVt5ThNDYFxyU5c3NyLT7lWXEnkljXCfbE8lZtaT0FnW7juX4v1CUde
TNcyULAkOLk6cURJcodR7kGeYJyAa6WrNHBQn8F2XkmDH9F+a3jg8o7eH5rn8AUB
6BLdV6ZTOBIJl9C6BLsif7jFghK+6xHiCOugS2rCLAamvF8RDqnTk23rnrG2OgfY
jNGrEtE2moQMyY732/OHiQx1ged/JCNJv53peRGZiFWjirYOZLbD5gaPzbAVX5Mf
QybiaCoXPsSfpOy/m8/55HsG2rAFa3ULwBQ0F0/B45xv7QkXV4kzZZUBJN5rchAx
xVdNzzXpjaRChI/kZtW7/3oVP4aqjXJfyn4POjaNSo1k3BJUC/RIAB6GHLTq0izC
b2H+YqMpf2GQ7Vwik3P1ilmYUSm7+4tjdDEQKz7gtGFy1JMyYiA06n/EOj6xEPm1
NV8gx3e30GjHhs0C2np2YARcQK/d5gXejssiD47rfNPXNlDN2T+xMyTy13l/lWqs
lrKnsiZTNzSm5iAG/Op1zOyw75V5oiCmvU1Q/Wya/Rj7yorCGNRoqKYZI8lRq9Oc
xco3gkBQEoyEcolmF+MgPUBBCcEBmIGNmcfI8ESSlbCINz3hkBlQA1H5dIm7Ih4/
4ElAJns73nnv4536ZTK2NARHQEk+DFThqOaXaPSm4gfnwzvE2LS1GT7m1EaBSgR+
9wr9O/gglh8zR1iEM+dvPlE6PB5ULcC9AZ+Kyu2QWFt4jfI0htmku/+CGikLskZl
AOjQNle893lPfmuyiTlvu36Gznc7tknwjquiimv04kfHjjhMvkn4o3o8KInPuEWS
JUbCYOfk24ZPclhJzXfOJ6fhyjYNMYabKTgMUOXtohrZZoVzz/ghI3uEijnEPHc+
JLer8nW+sBlw3Ph8c7btoLLr4WCZ8WDSYHtfv4qJ2bIh8EgZS+gxkaXiIb7Sdw7l
2qcgQOyHlclr3bU42G0koHpturjeHbJRr1eMxnDNF7vv9VGORajf2+jAFOPmb5Cx
X5B7UcwHTCWQcqHvw18xiJBdxf5JRsL0wVDgL2xVMCHcDZklLgvBeUtjU67Vp8fq
karvXWBdbWyO+UzULXAxINSNM5qAudH9H11/nkvXRbuOe+mNxbMIwhlVM44HWsOa
BG4XDsBTd6pgtO6/UPJ85aVEL3z+oMHciqyw5UJfmkAF4XY8t/QuuAXIIbQHes7O
N6uUdFKIc7mLv5INjxEm/NIVoGeU4I3H9jf3R+vyvB7AWN1ZxqgVZqog3zVxTSAS
KILScRYYA/n5GIvT49JsgAI8mP7RqHQ/8vXPtLgmb19PiHeB676gpjZLr9rM2aIe
P1GveRZMcSiIn0xfgifMJSFXFpeS3Hwd27lh4fByBZ0sEf53qbzJRO1EDFe8lPKv
DnD6g4rMlpzD/Av6RW2CC42VnPpEPC2f0OUSSePM7fCHiXw42mG2SFBucn2PwWW7
vjBB5jH3W++Amk3JVhPyje8r5uzNiK+ZhJOpKc27Nuxz58SWnBu8UNxM6ZcLv0Qi
FjQyV6y/jcmguLP9Eq5rF10apODyrKGHM0HtPQlI9dHKLcfe2rq7h6I+MGw/xXPO
aGSAQ7UIEk4oBV0SG26/Hzna+CghxFuXpXHWnD6vymE97GdGibf8FYB9yB9VC5nI
kJEz1J8gO7psgVl9OiHOPfKRf+fyEntXeKMabWahSnamcTrrNmRkN/HFDyll6Xvt
sw7+wQgMO/o79cljsfNw8bfb/fpKs7aQ179fm7CpLZUl8XjdzkeyDgR0Rzjvs63V
172Hz6OSQSnGVq2N7lLhPbo2BYoNqROuxcr1z6OHBm0t7Sw8u+0KeAkx16N5dHcm
heQZNeKUvpyydas1vN3kVSHX7dVRcThTOXts8gYLLY2nelqSJ8czFl57ibvbblbK
OZ/aFrL1OlA9CY0rmOXw3hdgDLjz7cbkH2Yi0v6f79IFdNQVPrWeyZuuAj2m+nRt
jF7RC0p3nHJstSPT+n9Ci84AFYHqjdVrxs37cYCEoYIpeMRX/Um/vFPznP5At4pf
gmEIrL/mKycggW4m5AYRsxhB2a0C96k/dLX7nfpWNw6nMpruL42LZiSCOYd3WcgA
y6bxzUnnBqHjQjibD4Y/HUVRCu1hXltyFtYoKxm+QR5GOhAaupgQ9x5SyIS9K492
PMU+pSWg8gOczeK1zbEEiVF1LFGQHO38BExdWaol1zoxe3hvb6rtz/Qy/lTH+Tpd
8Eg/WcQr5haewdznUZsPpnfidS7JOFEgJixeLpZRRS6Db32fVBCDo3GGyyKBXGIh
qvVN8G2An98cBrXFVm9zLx02NDU2HqzP1Lh1hcpJCkeqn0U9T0wn4o36mfpnvQBe
saBtK7lkNzNrNFocr9kN3TIGIFpQOEA4XEarFgiQjsA0X0tRiOkWpqI5frOJDBEw
ef4SjdYoQOdl0lw2vHY0ltO+N39L9gM5CIbY/FYI1Ufn7DkEx2rDwQlBvk3nVE19
5wUCFAxtMTRd4VuoA4btE4gWK29pzzwsDxhHnrvTufk/HaSoRfuBQ7D7ZTn77Arg
31az8Tmr7wP3v9UwBAIAFrCu5CF7xmZLD375/uFH9NR+Ep8M07mrxw/BQPu7BPx9
4e5+KqF2Ri1ds0foy1oZJHTsakVmeokJ8clacqPprAlUrNTM7ew5fvyi1e0jr4tD
tqlpA+abopV6wh/XVLsU6bw2eeLbn3NGQuKg5/ZwyLX/VmJmfw3D2clVDXjnjTC9
pZxhrfijBF70wP0BSXQEBwZVHYrUUyKIjioU+I/BORj63pOBP5oUBzoOgU3QgQ8K
RMntv+Z7USkF/nBt26W9yXqVexwWfGHgTDtzkvuVtpVO0/IAMOFlUekBtwOCMSwU
USdLO+aeoIVHbDYEzOxRkeqss9rxUSxDhY3LXU8e+4PHpX9UVezcb//1f6zUr92U
GaLBG5prvTmOA1aMJpdDdDXY/a9SqMoNrhhUJoKfjFfwgeGWqz2YvxyjBbkrHWJM
NcSHNoiDvuk4pdC8/VT8R/H0T87f/uU8ptXCp4tBem0C1RkdtT0ZVGNMRdVA/ZSp
Ywr/Bp81JXZVVzBFeXg5/ffkwEi93uzcjh1NHP/poo7FREGTuSrAwfHib3/CoVyE
bLm13N3hr0isfsh+liquY3cxhFNb39hufIEVcOsNdwXcSsC3RwzDf9qqvGIx0fdJ
J9eLmVOjX3V4z7Gj3kerfGs5WvuTk3wF/mjnLubfOcD+ecgzGTN+Q+ZpQ6XhIZ6/
ct+R8iAAFM05U0HpSY50Dbfn0D+RhlDfUE3yQ/Ir5ydTLLSf44TT7QsQuhaVjGGn
f0aRs/FZQW5kKnzEfKwWyV6+nWBRgPxulvh3mPBdm9Hokm2o7pO+YLPou57UjzM/
mx3D4CY1OlVvJ2a9qSQMUlXLQDIRTsAKQvSqwdTPUBiyeLFu1hQLwlqmLj7aph08
Fl+1Xff45WFOgww80HzAiJjd+X4yW43ZC2AibYFubMjdeGgGG/g6/PwW2qOkYaES
KUV7OrXcnNCYVIMT8xOyCYTDyKWKS94P5QMtj56pScHh/ZnkUSEC8eWZKohcw4t1
DZQV4o/S83FCHnh0cmR/TDCdbHm1S8fWBDiJE42DvMrP/cITQjx5qhte3VXIIonP
OJL6eq9ryXgd0+d63gF0t/0vp5fjJ5sLUr9HNxhsrv7qOy0B3CMy+xGe9M4Y4vYj
EclsuB04b7fynm6BjftL00i44pW6Ryd5+4GMGaw93QXhm+r65MU3ywgqpB3wEN85
fhM579x5HEMCfXEpk2hfgfrN6xoESJ5yoksi+MQim4SAoeItWWI0eyKh78dv/JpI
PAsgKPUzWYSUF6uSmZX0Kjqwhivg8BEXd2755WNI2eXxux4S1khVo4afh9lj5AZg
x/qTZ5S2zqdKwdDpySq7iaQKlKXPXeO0NUe8lNZzkOY/KArOKXGZIvYFIGsZ1LEh
VjnUAJtCXEHzMDZg0Pt+viqz1tYOGv5k4ep7frXEwHcuERauKgwg5oW3LH63P6ZT
6xRh/+ZUm3TQDQy+IWtdBdy6q0wRLqz1Z4jyfjMpgB0kgqXWsaVMYpA0Mi/9bojm
sWahuyUNYDV88R3SNXkhCWLIvHjSEDQTlrMzysfUXN2uYrgBH0YD2e+zJt1bjH7w
7R5nsuK0o9zYKKVIaGVBhKZ5EHdho+etPySirVqrVJZgRqILn/pK+rDiluPpTgxe
yCSB+0O6EMB4p7yaXX/QYX7vmYhiLgBzgRjSCBQMdYv9meyFQ4b1t1VKFoza3PWw
5OKkmFLH/3ZkM8t6XfdBvf/j8nbqeI61V5UoQsIW1K6w7SYjY/jxQLZ6r2kKIDc7
NecFENkLT9J9F72ErABwkQidZcfJgcwRqUyTBVSA0NarZ4OcQoDnmcTXkwUElezM
mxKrnZPNZD7g73p+NIM+EfUZtv6fSF3v3FX92u0uxAvMG5EXnjHdZvsYYmm7nKfI
dHQilBSMRP304EezhrcgothVFGOzclz4mIRDZbbUTD4wlQERj5pe92k933AJnXHV
OZAFXUc/XTIpKWrpj8krLROJ4tm8U8BF+2O8wdm9hsKas3dkxwteLiMbnK+gqqrO
C53oq/kKbI+0LRB26N42GeMWOiMpjE5w0Fl7U7BmTZ1S06KoASI3Hran2uet4X+U
ommzEjDeHizCYBeOE/vbcCnRFgD/Bn2gOnh86bY8UI8Y6PUTheVmtgdG3orb9SJJ
oFtqSRkrmFcNhZmwvX7Dgsd2Um3e+Z72pHUelL+GD1jLhc6b5bt5PQvbgNNEkRP9
Vvkx/mOUWJHhGWFYwRRZgqisoLMzL1MMVtB9Fi8hQMqnyNH5xgF8oHuAxB3Xp0bm
RxrR0VRz7vsVVXMSo6Jy7Lpt0YG/QoMmxGzrlYgv/awtgxOPePakM2YOfQ17r0vV
FGZT4EVPfNl+tnWB2hpob5lqRNA34kIV/ymvqQWMubPrdGvRnFAaKPJ0SlTQVao+
e0NF8qjszTsEpl3SleXho4rOiaas7CzbCN2wKKIMGQGJjPu8JpElwToG1v7qtUm4
gXeZuHZVspmlB0CxpnYF0Y90VSUAF7quq3VVRQeqoV9ka5E+gWTAcEZwVZfq99GA
JrZYFxpywxX/M6c1zuwuco7GIJGvtkGsNy5D7xM4Hzoab0+Eci/kEDK3qiBkUgFt
2U+4Ea+W5VBo8puoQU6hFQA+PZbQb0HIbUtvU2zSkE5uZwe0X1ONvuzv7Nt+Ug9J
ZwgJghqLO0X6mSwrx5fyZ89gQ7nCukDhd2DWkfDvOLJFx/X/3fUlI3quo6OhpAyE
ZFNdVn9RhEK+GD0soP9i7LDsS94mKCbpJZ00QsESKjPnB1ERrkLPQVRbSVhe64ni
92GnkeP5WbWJ4oHFKmxpWjpoF4UoguvTe+GTHQh7Usgrw8WwlW+vlkM0wN/UwZQl
SkVtoILQOwEM0GUzs0E1vS0hEUsy3n84/VMW7h6/kL7/MSryFZ9Rn+qU0UsyWpBi
uDD1qtxtJEoQnU3c0wVA8/SMYj2W+0fNUuPcZzAy6J7BioZzYvhRUIVoJ76pHQ1+
dpm54bog1TA8qjivAXF+F0qFjrbvTIcZf1R2t+9lVvcQSpv2qfGYbLVtr7qr7J7b
4qK7IH1mUwU0InsCjgXJZGaVFkqmP1xWBNdgIlGHmSCcZrIQ9xl5TC7gI/CSPBeW
k2bPNv3juHIZacTJtAM3G/1Y3iFkxL1TUhNEZ3rJpqGQ7WxwQ4p3psxGJR9+H5dE
Dor6MwMUO9qkgiK83dFIh3ZdSw0tF4p8ibGkS6NjQ38bxRSKHj6qve1i0OfEnqmO
yqTaa38lKAFlapjYmQNfYdidw0V8MdvDDlOWE6ze00nKxH9Se34hKcJts2+bLZjm
noYqsFozY/Jnd/WfbrktzABT8t8a6ESsGOS8LVpuhZGUECO4y70hWRIFoAUs56gV
aJux7O/i376SD/NudUXxP1OQcc0MdpyzltyzI3Hmf20BFEZvvPPesprqYLzFXXmX
hWLqeO1pB5k44xu1hYnWrPru8uBChlQs/Ov/bcPmlV4xa5FuP7bTRGOFts/po2Ei
B5WQNCiwTprcW28r+17bdA6cYCJYAt8oH3Td/iuAbHYKaa2OJ6jqbmKfoYUqFe0L
BVPOU7nz/6SKEUSzo4NO0+3vdHtphi3avK5SmhGerJd5s7pbiwmXyDgX9bm+BbAO
Ze0QnFdk+DTxHeI7TytJ8dwfLQPF7vEx1Tw6wTAIkCqCmylKvlktKJ1YrOd8kAiq
AdMRujvOfxpBzWAxU/G/XfRt/FG9lWMsStapBL7sx3K4ERTIXb/HyYFfNaYaR5fx
j4RuZdap6sacwYbuLDZdm554uAdZD5stLtVUJzQ3EmgZzUQFKX8eYWigvHx+qH2J
X4CGthzI7Y7zce3S4UcgI7LCve1+0EkaGo2UPmtiE9Q21iW+WDEzQwHRp20OrPfT
PNzv6tHIeiUut261R8pjs9Bn0qHIarzYD5dwqA9oH2ufMyA9HzD//M18baOGqEEY
IhwvHouPWN+NQOjoTiUU0igZ+iYpEFkomyh9xsE0t61Fv0igPcmEn+Up6VZpsS4h
VMTXOV+z/OgOKTiopuO2L63n1rdgSjlqIpZmslM5bAm7zxJoOLuZKLkn1P3OZD0y
83KSBEeGEHlA27XZhF33wBf6RA5/iFdvapvD1cruyG/kboNJOiLJ/He/sX+Xu8lT
Rbve1iM2g+WRnRboscsGC8m688LuMD+nDWYZYFryek5xTtGWn15aTRmOUS7dK6wY
kw4P4VdZFAsPgHCSuCMO/slVOV/MpI/ThnMWoes1affHjddZY8/dx1gxdle6dR8+
CozyxsbMyX0I6/xMmyQOnZqkZF2ipNLQbUCSYGRmgGpKDakJpimbZeZjZ+Fe3zv9
xnDt/zd7VFfUURpRpwnFZVEy+9cxPjLQdxhHItHUMFosgVX/uGmZ1i+3aBDzf4KT
/3IlXRD0ykAw9bWFrJ/CzWi3HuJB2WE5KmRKQ9DpTiF9IYFiNQemps9U6wMHjgLx
WFmIPeDJ47TZUHaN6PUvIydJ2WoIlPPdhpBEIsJPG9U3egNemiYDQjN8z4E1pT5Y
tdJoYPZtZkv0MqvYN9NuIriGM5AHe3rNhLSdhoslFXl62vQBQl/hnt0xBWdYdehe
kb5sKS+6WRikdWXQWJkpdp/s2p7qcTKwR0/vXtY742gxhq2vZ2Ir2HrwjSquaAJi
IOW/yjw9PC168jb+tztZXoIMw7tuLbtS0xeb5iLoEErGO973IsBlCbP//yoxm69V
ApIxdP1dCcp1CcaIn23XBHmUjzMcsqgv3I4IXiekckIZvyCSiVKxTDau6eQjU/QZ
D3nD2sn0X9OK5+673Is+z4pQn4ijSa4P9KsNJ6eUTCnNRHV8mIs9K+y+jv6dzTXW
GcCbCrqQBEZ7o/PKSVpNP+jQhiMtOuSMZBV/1tCazsc9i1zdpuKgYrwvmQ5iUnNL
51sV1VPdq8WgQHf30NUBjOqKweQVJtkr3QvsrBR1yMnaNSvjO5hYIZYGno2Xn5RH
/nu4a+r0LfrlsjLuvwMQiL8tEyW04z6BBUPQl/Fs3DJs0D7ls8hu8HkNQeccx/I+
mfIQkLSKgrzdxpOW+PGMqh0I1e56ySLR4as4pqu2wTngSvJwYvxORubOnHOpZhdT
7B29d9h6BW62cqvbQBd/Ml72iqorsFuTMitxW+KnSV1Hqm0d17C6P0elkOF021mm
8tPCkox/sZof13K1TXCKTrb5I22UCyuvuXQiDK35qcLzBvK3uxeBMj6KE5Ayd3an
hE6IAXl8eOjGIuHAFBi3+BSMCLik+xbHq/2tn3rN1gjhf/3qclCw7Cq1u4U+TGpi
EBU94V8h9l7OvempfRqNPnBmDrkx8E7LNqLv2W3ObxFrDp6CEWEstGio3C2Teup3
V/ncGTLLPr9Lwsbhq0BR9V2fZhiwEDpZ1K/JtfyRviGsfyy1p7PNI7fKPgOl6ox9
TXBMlWd2pFup/m4TNYFcqAnvnW2ZIP/Dh++fZ60QuQyN3mwGmWRry66FeEw6JwpB
G926CeAlI62sBnTmug0kBvEuRAB8zSflysIcazfqveajyPX2v4kSg4Qa3T2cKmXq
CUJch24DGj9RMv2Bf1Enr/LJWyXDg/Nh6T8GLr0J3m7WXvbzBECLmUlNB5Fm2abQ
DUlGLh/8+yqHtP8Op6/J6kG2Tf9wVa/YNDrIgl8YNJRtTKvIk/Z3MIzrPD0q/4KO
3zBfb4lHXW2TObU2KQJAvC1dGhEvNMZCsYuejWc4+IYVDA74v5MA69hsgT/aVC2X
+pR4KkAt2tciO64UEgvzg/LfRgB9Jfw0wHt9WLeobUKdDM6gJEGBLt7p00IuacLl
AszaYJ7+gy4YWx8+xSUfAijdR4pMJd6v6PSiy+pIF99VRtWx17UjMPSjNnM7JIVD
kV2pEsgApCLDQcwO9a7aICpxlSM7vfgTeHutn7FVsYOKVmaWs1+TC5q0bKOzV85o
BcjxNSh/YQ5hO6Vbz1uzhX1QtxIB1qUYOH/JLek7pULv0Oc/SbjPzXmEpJgUcT6v
OMfgr3d8j7MN6zkN0QZ9Q0BreKZh2dyAXS3oV+iZ+TFu+bn/UC1woF4JyoesWU0H
KtHk/Z3PJdnnA6DdgXSru/x3KWnwmleuyBxCzOyissLNOkwxMX8mtyxglWRwvxxB
dt6OiGfCdNKizTqwyOQnOXoRht731R7ZyTmcXXHD0f8cdVK1/M0E4BEnY3aePWF0
rwPwx8J8Q6Xkjg1LHxUh1TnAC1Aia3xFBP5OwzC06QvEO+xmuP5QxHPdjfNiCE4z
+NoRNDtThLp3QQ/P4iAfwD4AMzXh+LxM4tV/Vn/4arMnmmYdbgHWS4Cn7iBmjSKc
f6Ici8tthWSIzdYwIfaVpqTcuj0Vi638SBSPmkhp0FSyuEjFpDIpZJHD0MFBnnD8
McaOCTV5ho/ZssppFsl7R3F19DPRCECfz+/25SjpcbYBZdi3gEcjSumHFCdNVAdK
/NFP7/tygI5nBoC87cIHyoNQqEh8JvQY1/dT2xEQeUE4gWdfvn370KbDNXoDdTf1
/NVNvZtcLVEtqmf3vA7D6jz680Y649mVZZQXZELHrkS499pZdUCmPST0OAIaHYE9
UycA5e8YbryB6tiTAuUUbT9h6pimQKcQs/yCPooMtPKMy6edBPVemA8ctiKoyKlJ
71tVNyUTRofWOpIGdRsbrtjGdd/n9MxB3luntMTbvevnGdsraF9+0XzRkGQ/qNeq
vgbYHYsdSvKJM4Y2SzLihVzAI1oO6+vJ88JW9QH0VtJxcBr9wsz3dSAyjM7LZ65y
FB7CNDi5N/dzRG0XAUGdAoyC8bOE3LpfLVwucHTxagVZU5I5ijueA3/wRN83jnMY
db29yUoH4XJkYl+PK/wRAhZONNp+hmYmEvGMtulfeIrB78SDqRZe5ujro03Bnxwz
UHmAlRiuHX7DVsoJ4QGnaL2FkrumGhABUqDtCytyF18X1RSoqDyfx/vbLbL8ozhi
uXaU4H1KFO6TAJe6QsTJOHbu6JV3mN1g+vIlrXywVX9tsnm/e7l2Oah8SR616XOm
TlrDsYrMYA5Qd1aVm1LaAPdTMrRmLHU84gq4YJkspQ2nfVZRKXAbfKz5zLmHkItC
7W+7g21qKPkrKtB813hAS9g9nNZTCqxS7+i4zILt0D2yNtDmbHGHBu342u9mPaNq
sX0diOS1jB7meNZYRMg6LXWXd7fHNZJSONcdkJiC0PdotwQB+aj2i2fg7uuwW0sZ
DNgzNyRveIzW1I4mSlyO490LerHS14UkTCDoicyy0BVedBOIbRGsuTLZK1Mpjam4
z7Xz61769x+MgELJZ+HNEmRjdNSOFnOolbwyVwx611ahpY2MbsQ71SMxjsGEphex
j9dfpWI5K4fFdSXvkL7/FF7xOjc8WNaPSjPFm9U9GNOScfz4vqmoB49Cvu12rOPp
hddvD/HWU2kQuHW4w+JXLHLqh96eKDpET0shKCVT7BpEnQeWTgCHKHDCv9w6oHjB
bVD9O7sjeQPVVc4Cht2NuFNY8QxX3IJTAa2FsMqD/D/53H6qTpwkPSggpvjvUCAq
alfcrqch3VN0Jd8fFdRULzwGT+4p4zyMaQAQBNQLhIYF9tzgwPrVFOfpWSbDgh7v
Rf1AOh2zAAHOU0yDOEULT4LWk8KozopDTS6Xqlk43sbTW4oAn61l54tNgMxT5E2l
OSUStpX59ddmi52p6tAdHHG6Z2+QF1QvnhnJNRrLwdA+KUdLx1cGPU2tIOeHv8F1
WxYGli+f1Zlp1/8/q/LX6Dt1J1EqkDmeLNWy02psE5h4/38AQp+ZGk5oZH1Bv1fb
7uoHIAVVm3Mp06peCxmuTT2p7m1ARACq+fC1t8aROnyWCP3hmCGyD5ADyPhU1OhI
CVrLkjpph1KeMOcrCXCrxYjvn1auHYR3751Pk6EeuEV/wq0MJDG/rIAGSyov1Lvo
nd/vm8PnqBQq7oVErwtZgAn1KQkEe51BYTri/0qeJbZhnpv21tjOfB/tQlP3cBIO
8wqUTQBrf3nVciOV11ND81p3DLm7qEs2HBOTJwsS++44eLUcB9PW/wCmyxzknpeN
uFcdohIm/f8gDL1lMAcmUl59zVS6pB3FpieD31XofarLEysF/po3L43WZEs/BBAB
QaolIplX+mUnGppBubn8oxni4uJrcCW7ZkFjTLtDU+Ub3u/qvfB15bGVrHD5vNie
6CMiGsJdr20Mp/RqFKx+HVW+xDjOX6OikXa6P9ccktAK6M8hbnD2eu5HJ76aiAzr
CISSdJcgDqRE0Ghqeyxy2AlEeIitMS7qvtQplal8EhMr0D7okz6GvDQZbeXPVApf
tHKA4N2Ci0PkefzzzFYnqVH+rKszMc4nph3v7k/kSrwnM73i4v2HsQpVsufmoKAy
psZ28PB3LZ7lR80Wus7O2t0US3joXKZvl3xu3tdHzCKTM7dn2msfmtS67GEyJKyt
bm1ocQJR+9pmp0ptRur/bOgIpYSq9GqqFyc0j0/WScg2vBAwu1s8HR5C2qX0Jqk6
787M81jsZvntkRJT7sZVFwjyNkOTFBpCfLh1UO+0mHSppZfkaIPytiTbX7X8mG2A
9J1vcAcJ0zGAB6lvavn2rvW0HJbMgwuCDWSe+tuWRaC1PIHD9h66JliZ9hAVn1Q5
RlnWD09fI+cZPdlHz0BSxF6P+/a8HiRWwk3BqmLZL8qGNmL/rPCKyewjQv3FKiw6
xslioUtKe/9C9zCPTEHpLcu66qjg3Fy0eCubAZ96JqkynAjl4hTHOyRrxAGrhGcg
1pF0kMgBBe7QmFNrNdTTSUaD+CjbropubnXfPbb3P5wF976zux+0knwrVN1kqN+g
Ph148W/RhbON804cD0yg7HlDE1OWcnCezNl8TWUXk5jQEYqC7QSr0lJnCGQbaiJM
bG5unn+sL5XTGLpkSpY/bBeAP3zby2qsS4iCyhjw4gbaj4+H5VjJXPy/bmtz/Qm1
tzrL9+1lmGRBpOVakWAOoyLSH/0U+CR3wo9i0NXYpixvPZDH39yYceQY28vrg3qd
6SvywlskU/DrsaZD5sAaRdEWrHiKg+t4FHRLfAd5ksbhecung+EunB7AMMjXFNEe
KHa4youqqX+tx6hxeRX5//3NUyw37QR6+6BvhgXChkdiqsSdPodYuvpRWNDfZvZJ
tb8tf7qoGWjHB1y0tV4njp2TNnEV4R3cwttQXTkVZMFEUTsW9nZ8VW0M0f6G4SGv
XoPo7XeaeiyO0Z/RmnwJ3UPU91Bt5wqXy8g0Keee5DHyv3iWiwWOkfdLsjw+iTUO
jKRpCeioiStr5pDEVqhGXnrw7/EDG/TQJu2/dZcnyYv3zrlLDnkkfvSCjzOllrTC
mCuEFiFTWwvOIfPj47Z8knycDEiqh07DWghCVl/KATQejRv/JCe4BCVwcEH9LIEB
FVfeW61/ZrO/Qesy2duDkbv/g294xw374dEFvamHzqyNpVuPBUrXLkrweHIiidH5
A7IdvE+GGSZ5faoKDDJZcKMRV/tor1+AswkOzZ/8FlU7bbsJ5QiqHvxLA/ql6iy1
amAFEIX6WGi5YdhzH67GpKLTJLsnkopqANJa8dX8FYlNJJNN+5xNfQ9mVwMtqMiO
rtEO5hOdoCuXiRF7V3K5boejMzWeTgyKfu7RPbQHMw4NcmuD6o6gkPlp8zRs1gtf
+9+3MeimZSwIy9ZQqGiBPVdVucHuI/Xpk0Xj9FyYgWTrcQHM9hLGYWsJE0v3a+u9
LUxYwOgU1KAcBQ2u8jahHWd7xDXX/id9TCkdJNJTWBRyvDuYhPi+4VrxL79NxTUJ
Smst2fD4SZcryF17P0uV020CCNC5F0n88ym2vJ2NSq4tXtB0+in/r5gTYeSCFLq3
fjG13wVTBjQQvdqnLg9tLQyNB0yXH5b8wBc5VLqHzTE/r0bsLVjzMHLvbCkh4kaQ
D28swQCcX3fK3sGLj7QAe8EJSGrGZeidc40k5AKh/Bi+kOSH362sWJ3YPvU+wqWi
dqI5XqHyQKigN5pUhk98Vd9lxAgOsu45NOZ5G5F9BRBKxPi33/BhCnvBDxQvXgEQ
P/vBh1NoZepSJ7xAkF4tQ9lJ1119KaYuvWq7izU18ETrAYZERoBmzzt5eVVI1/9W
gAJpJ9d+PcR6IC2xwx3jjK9CV4KLt8qgH1lv5UTmzbQLNWCFu6n+WqTYWfihh3kH
gY62CZH1XXcbSeHnJAfq9TeOsP4wp72v4KIQGmX4hVUg7QXYO/KZLSfOrmpRu23x
DkAUmVB1HepCZ288whoMeWIwzSKk+JUpNYnlV/pZ1RAJEsRQcj1fyU4l0ZHrCKI7
YOPDfXY/yP4ehHxDP6i8ayV0RrgSomHJY0nJ56swXqPlIA+6l7jSazRSnGI1wkzI
GGmFb4l4tab4PxBdmfcDDaX7g3hoT46gMEG4Luiocjp1ic/hsx5UMYv7NlVIsEbK
D29UxusUj4nrOKATkGmj8lQB3rI4xmiqdXq5noM0Q46Q9Zz5tTKvnuBg5frcIoeX
QYWHJ08vOKkg1ZCmq4KIp6qNjAF84ilP0tWv36UQOBCqGP7DTnGvQPkTjprmidCS
7cazC6MMx1YkUBYaVE5uXjxzCEj16NHS0s6CghLgUTlXwMcis4o5oje9OJXENg2M
OLLnSTjbODu3RoOafHMe+ELhhO0shTccctLoHh9dODf6DcwWLYcvqS/7tPsKQxir
Mm8q57b5oEB1KOBzJTsEBVBMNFBjicM4bDXenswXWT9N7DySgMfjxGHLETrJgjyK
dNnyXlLqm3dVkNbhGGNR94FSFfoO1qARv8AXR2UFmgYV0ldPeNGJDR9tMTQbYZiX
1sEEDTo/8Y/ubJblm4xNRk0j/Ue4l5t6qI7HniyWXF3SLUPc/Z5etHKomOJCaGPP
8M3ZguoGI5kJS/jPo9SeIv0vsVz412w9o28RSvTeHFy5xdrcaNBn1nOU3DUFKZUL
X7CWoLXHs/CRbFUSvb1I/nZXFg5hUfXoediNZWPGR7rzGgVWLwR5ErGICEDpLM8p
vBjpkvpSZJuhm5+4mCEvj3o22SfJpHhaWOnnu5DZOuLnVDOKib5YR86kZFNGjbeY
bSDCzBQQDwyq5J13TSJz1j7LqBctmiS5EXqYCNlXRyk0DZXZ87Biz80VDkqeakbY
q2eVE0Xl5slmbOSsGTKL1RYh/g42PgN7rL/8LNXIcRRkYyszmh3TUj+8PUh/3EwC
lIW2Nc/tpWOoHE8Frz4ULttj82ccdkTrCitApSWShwkrifKScCiN+t51M4Jf/EW3
L5sjivRnEKwxrdh3GBIpVrfmtGEz9Xg0NLeOExl1Q8YDr2FRVdxhVvs4VMg2CaK9
bKnlHoXF+tXB9f+I/N1Odi2UE32qew9n1vShgs6ZTMEOPp9o1LBrjgeZnghVOMH5
CeANoz1fDp+u4JJN6WGK3jgPY0kPz7JpdeEstgnvNlDMsFf2DqkejQDd9bDKVnqJ
JnSZ3Qtg1fuXhanCvZ1IbBO7Lv9IppEnXPv8tDW26Im55mbzL9pZcyohxyS1hw4T
ZqE/HrdBoiZMbpMXdeYPsvm6hQW6eQCEFr/1rth7SfyFva3x3VYiQprXFNPDscvZ
pw36CzvUf4WRNFepNH/+ir+W6ZMoT46T7fIqUvZ0EFEzQ5B1VhWjLdI0oF5Xdu09
MJs2qCkvqihpB+OTaBwaTXGnwjvXekJV8NxtnawHZk9rJW7aqSQrXEvO6fK+8Cbb
Se9tRfbM//ksFTI+KBkZmKGbWPsmrM6VVgsMDEVbsyjvHSFF938ol6aQEi53hRQe
x0Quf2YKk/IvJsBiDrXeVwoOEB9Bocr8xY+/0d2qq8Tg0EJJwqSMju/ulBbDucMx
+Hvvt4D7xwQdPPMvsFIUuBqnRIxHZp9rsMCIvY2daLNOHJJlpWWn9DtDHnaZ5YTi
gUCPVTKR3KGfPm7Fy0kUnjM4LRLQpuVePeKProDiy9xCozeMHUMUkkBrSHftCxzi
cYeAJAoIb9XJsYtgiB/vWZSXVqMWShR4lnKZR7zF0oWsGmMvHtV86WVeO1iD/qDU
upDGO0/tbTMZx8NbwCVyPGnjPhbwqtf3h5pOeh6rzXzv9QALZI6BwOBILDW2t3pl
wL7JK2a72m/gmghw3Y0rVbvgVITct3EjcOvBJi/VagtHql/6yxU3xDM4Gb5CWCBL
gAV/E6Vm41+W4c6tyffINFJ+CfvYXaKHiiyyHIeSDvLQb9J71+hK0MsVaYTOEDWo
CB6hyjSsIxU0ydL8QI9UbinDIOK7R9yl0tMvVf4qNsawGK8LNFnPlPWcmcqbK+g/
LUKSvSl61t0GkdmxZobTkJ9bwBvYL5vEUGC/4heBjFzF6G214vydUqczG8yPluOp
7TysExQoNK1Fl0AS7pujQmn3/yJs7mvSpz1BvmVkd7kv43Bh4omfIRhTZ8oyUAof
ELVGc1YLJhTkTpm7I5uJTU/TberD1N2rJ0jpbd628lHFvzjnnGK3gtYYN+3R0r75
gy18x+TnbCe2geDdwYefgd6h3T2j00mUXl8YzQ5RXHfpyUbXlox+pKTWEJV43FSh
IWK7lo9BGmtl3EqDdW3zuYDHIPT5BFdrYWjJ/kUWLryIDOrLxGpR6Khobpox77N0
CjlhAJ/6rwljAuftVAcI69KN7u1i0vXfPGHvVgoMTMg/DPsc8u/G5D/bT2TQHhey
kmW6jqHZUV9XZ45GTmozo6Ct+3Hrpr2mXLb90uKiz3XVCIFSCmQ65RVbDzmIVWMd
AR/704yfrlTCS+xlX98H3UZzy7biDgTukRsvhwzhSxRHSTsjUlGcmiqYfhoiuJVn
b/GPJndThOt5GKWEQ46yPeazHPar7+arLkITzsRZRsZnKa8RlJLUr7STFHQEPn4j
vnZn3zOFg3jlGlKAmPaXWBKxJxloFsOxB3JTNFBdGD8Ugu3q6OQG3L+nZDmGAo0m
T4C6OFholDMRLI1EHX2/Y6+YcIyBBHf1KgBh/o2R+9H49gKvBwFTLP0OWtfSj2rk
dghL5U9sdR/eEhsK1emU4ws5TbtGpv1LXCepSI8bX1wk1404HkE5IcBvwXRWOQ2X
jd0dYOcHAJrTsAJ0zL8UgUUyZ1hZpLLc2UqzvrZp2tJnCGD1Yfka5heSeK9PY9sk
GiouDYIxPfOwFRsEPSA34jfVZBI1r0WSHfMb9NBn9SckygodhVMhV2T2Q1VeIQfy
GYNk8iDAQSEV9joStnF6aXEGUZMgcbdSM/wYinhQ+tOlqB/xBU0w/grxVTtQdU/Q
d5NK8IMGAuDTz/iwhRZ2iXKCM9WxX6gf6i7YbVv9JVRcjz7qDwsMR6bjzRXloXEv
Kr8GlX/F+U28kXj+Fjd9VL8+AgcdIMKVyGXLC7R0HqPgLPRLpK/ko6JrO9YIUX95
IWrMwbWvrGDQaTnqstwwPdt7lFx3eBzMUyzI3jjjRW0vsj+sr09UqYcW3g4uIIgt
RwN7PR8IBj/VEmYFZV8YC3RfeQh15h0eoLF43L+6Z7sjV/DHk/Pb2tGQ0jTjmpYG
ETGGxqSxpPEagHnvBiMuOj1C2msQq7sG3eJY6CX79F+aedYVB/o7zSOve/5R51NW
VRrODK580PVBawqZ68u1TFzfnCeLnt7vtT5Apvrixmh5gE0cKTV17UzmMXeOqyiI
sWA95v0z3aChrZA3BGiCYKVkEoJ4DOYBGvuuOEJPnmeuGCS5XRXj2btbAptBirr8
tR7K/Lmqfiq1NDEq2CyIKPNK0LRFEpGeGr+pd3j5ivB0z2Bf53JK+UCJTlRmss2a
H7SmbDd6ZHgb6ge3FI8eDSUVz6zR5cKJjSCmCwM87u9jGfSjpQ89+zcjwOJhYXvo
LrE4tnrfAuyl86BwyALd9/nRDyxoBEvZWqf/7nbCUGfCupLbAF/EoiqqZ6sxf6qW
GdSXYunDw6e36XWMGO1ZOS7W/X4CzKj2H3zs+YOUdAIKRXJuX12rYPxVJhkttYOL
pFJAaJQKpuL1s1JMA12xXls7HnkRvwLBsh9AdqPAyROR11hXSYGEMgLsuCEaYuYh
YVlwUu31odcjeyJgwNdPKwxH3nMMijbbJUYkSlnWnA4WgQ370fVbm8T8Z4awUCnl
1JucbkqCzMaM+yGXMkUNVGRAmr3X6XrL+u8U2rMBss0cFmCGh7lBUrUmpJFq6wK8
ORq21MEOndit2XLhEEKDW/h38rjNQxjA8VsV0UFamKO0x0aXKziKSe/z0TmRn4Gq
+v8b3RcH2oum6U4BgNU8la93IcPRT0XKlD+KZV2n834jeiUs4H3A9rm3xZuQFbga
kgHyo2Ei3CveH2LvPaJEX5Ohu/3NVQE5urEUDYZAxDgcOShf+Y6QfbEdNteG+lsb
hrPOFf0YTY49Y4iLcCrrNNXYsfHgzALyuW8m8+AXobQJw98foBeDdKbyW/0VfQq1
ThHnTYbaBOfFlXeH5ZyRvAniaufMEwbpdz71ei5ukyHAloQRV09WpXP427RLZl+5
KcWzIGQKlyodfFquSOy5pzGzJ1iuORFzplV8+rYOxEfMscvPLV5O9YSNQDIRJok4
me9InKWLOs2gE88Z+aZmIzJsYh8oqA3bmXhdYv1E2aXAB9VnJ3vBdhkBW5FPlfZL
zjhvDk+e3K0EJCm6Xin25ktdJgAqQhrQEVEhOGPPRsn+iMQonpd8gukuRqg3uVCP
zOreH3ntHEey8q0TuV5xATK8HrIFMR4cJKWx0hAAVxlNCwNnStRdQLndbAcZGR1e
gKMwbyO4HYI/9hJB2nADj0SDzCjnacyGzBaTRvZIX5IHOEm/we1fZJTMnrcmN4FQ
/R1j9mt7fE0L/UATb8Z6uIX3Dv0H4otzgb9YaXXX+MEfuedLofTFneVysVFfAPfI
2gzKd+/v34dba+ZDb2xCWSl2zSIkvBLKN0RD5FgEoNnARzC0y54+p8v04EfR7GS2
Ikum3Qpw638M5N4Dd7yJrRTxTSK64Ohy2tE3tyDR4HmWXS8iPnUdWfBx9JUG/V8F
SWzuONASq36/FuGEv+p+/KP6pZkLQjxtxmyrJV+QuGgMA1kSFUjT992TvRywAK0i
M1OHkKw9YNO2yqQJmBDrm/DGVgE/oaVTQzIupD4k2Su7nhhMxOp42W+tGv5qIB9c
gLHPH4fDyZq+paDwa3l4A1B2q2z5zC6yFJvp1drIsNthRvLtotpEHL60DU/Vdv51
zhdACT/J7ew/37WRU4dmOsyRb+oH/ZAXZWQh6eMcDb+lhpJ5O5jEHrj3gbLCkZIo
LVfWccNwkJ/TJeV2k4RnPJomGIrJY+sEFaQERableQIi8AIvOkhHASvqCqIJeQQP
ihj4P7aWBmP0zWx0HOcfTdHMA97xeM/ysC+KZ4MNEZ3epO+GyEEaGRpc2htH2Qwz
oz4JihJS7989gCztS5nqWPo5OrHUaaZy9oqAWKpEh5qKmR/xonW6uCwgqy3oFoIL
sohzkuaZm9op3GfzO5/beVBpVEg5nB7FBMcPNXHUfrd+w1XxLWsDQOS4o7WOAzvG
TE3oZGlitzYIpwtzbr9nyYjPA8UnCXHkCTkaKnasTUJrC+7JejU4RxZq+Z/7oigr
wfOszLHTA15QTzAqJuACRypUoxpESKsuk34VaaN7eRxcQzIjdN0tYy5gyjMz7HXe
TgdbfnSWFRZ1wk8aQSwdBJG765giaQQHK0cpgNC4eGC9qHcG5HrxIRgjsjfJwoIb
cG3N50GBWb7HA3RGom6Lp1FF9KaWnS9TLObHCIc3IIdoWoJi794S0b7eYbCz8K50
5VzKJLT5pjo15PJPTybDZwt2g3tnq+JLAhbNzCar1+Gsj7qCzugft2Db9yP7u4XS
AgnJW48medor92FsBCyOXqu8engrFHXO+DLKlavUhniGASRz2D9U3orTl/qGr4fI
1mLMsZ/MI7+GRk0edLA98j/5N1/C2uiYQ/0qLSXQiuv1QJgb0KBY46vAv4Y50h5Z
dRjgwg0EMxORiYtTVd4s97ieVx8iERlQhGCReKx+nPQcYHhopI2/O2gG1REYRZBT
gFTi+x9rsJlB9QMxc9JtOc4Os0lLcPaS1vdypYFdhLloZYCPyxwuR9OGeb3AQH9b
hPF+cadhWURv5d0CwuiG7h2+KcdeDhMCj7mqpG2eIYR59we8pS32GUTmH5kDknbz
c9k7OdAPLIQyLYuCsan+rxwEjcc0lDTD0qe8SiNK5Z38GQSs+NkR9S5/dSvoyc2T
1ofcxIoTTHJxIe3z0nRNFPBpx9Wm9iYo63s2Zx1kaJbM1Ss4g7KoEs7Gnbvc7USY
JpYyAF7+JXbZt1nBguIHsTqHUYHQEEHIjcwnGN4TBs9kbzrv/kGUMjh0vt3kkTEN
UbQtNvSRugYoqY8EOuZ1U7j+G+kSs6jbXGgh7xNgrDLd8jfq4wuUsAI2o96AOkxM
ajtEwhWHofONiSqIdcEPglHbhb5YsBYHn7xFVUmnHSz7pb3ZceSx86ys+AFmDpIP
d23I6wd1FeYrbpj84inQBSbNTMfe1/Yn9Ec8pDcDXfNv4wCK6LvLPVNKPABmfOBy
OsjjJ0qGLfZbxcDuxHZdK9vDf5ao4Sng3gZDXT/YFV5xMbNjeIWuR/vaBxSlFQBI
mO51PF1GbFexrzvfk/PID4mFy4py8G/3IqNRulmSLxYQwWWCsMfo7slccLrNjgfU
qPXJ529UsyAQHUTgATKXNa0WRhgR02OF8k6uN3BeWb4iwxGV8Fw96NUSyh0+WTKx
T6b8X6ULVS2y6jgeCxzeYt0eaExyLqHX8mvH5trBg446mMM1q+cY2WnTTMH34sC3
faa5pj8Q5vfFRbecpAxHkj13CC7mb52JSuzKTM7qTG4v/e3Rrb/2OKinVPCkidNu
b4klWEwOTtSAls4V1cCgUEHcik5IzPyWXcA67SDb9dp0vkdOnThMO7Bj3cIJWba0
Y7cSDRjYud2vXd9py3LjBwW16xU+Omd+A1lySR5gujhDhs0J6mxNMPFjjJ4XqCC4
z6wcWBnrRQH7AckR/Kutg+bZb6QkwTmu1+fGujwhbk0HDUeU2Bm7LuBNZWtgjWKe
Yqz/2b9ymJ99PSS48eSeJiIUM9YnXLFQUUJ+F0c1igdc21LDBHi23kM7kaxQCcXd
AQJQRgPGlFQ3qdUISmgR6+HkUIq5GoI2miVXlAG4jwICNrSrCZYFglA07ZK0bCLH
072FWkj7hM1OjBYhJbTI/WPDa7Q8a4UHU2Zs3w1emQcwvY+uAtciKg0kSmQNtUqG
bXvSHisA+2mpY6krzQX1G8s0PL8uluMSuPuAE378KGVplRGem1uqkWGkc+5OQ/5f
h8k8oxnRx00v7kzyM794ubIMESyoO9o7vHsCLBP2JXjijk/A2c9FlCh6JJuKKfln
aFlpQG/c4Jkzpxrd6fj4gjbl1QKo0eLnhH27KD7CkMENLV/ibOfL6Hj/av5ZlJEd
88G3RYHJFbkoCOxJouUp4H1jf7K0Y9hblQx5YTgP8rPp1GGoljRM3eXY7G83h6yf
bVsgd8ER70Kx/fBwKqho08SD+hACTmxI6TULsm9bw2iuS9A9ezUWLfZ+KXU8htmV
SMNXC+SSSL17bcQJ3tSqkMZtoe19SdQo36FTDaG/vo7mRX6OhIt9eOX4NqZ6D2Tn
j/h0IAhbh1p+RquItwrC+7q5T9jnAJknnD6FRjmc+ClHwLRpmWu6RXV1VhzulRJn
lmSGIqvuiRUI4VhhLIw+WBRsedaWZ/ainIRHXvLFihPxKkPw5RWPhXi1/cgd+GzZ
IrASxBZCYtm6vSjhGNYn62lYnySmKE99BcgXNvgeoI3lJr9txt3tv0nRYN80y/Zq
p4YW6FtnXceux5r1wiyfeUFjqtOuWAYJ+3yRs0WcitIgeDp83TU7v9KnEMsVIvt7
v3ExRgegPwwwTHWZ7mWYEHLtyltVrSdvgyS7fqoFrjGbc9+ekqg3suRECRzwSeTL
jl7UCQ+ZAJc8W3fg/aHIcn30UwRdWdZ/s2f+PofOVIDkTHzYFSDcHRwA6/mSVBaD
LNByuy9HmkbEUH8JgNToau20/Rait8ejGxPoXkYm78Rp/5lNNS43xND9rYiI9uaI
8Lr5j4dIzJpxpMMc3u7ah5+FuqSe+9Q89FJ/Uoz5HWGlRoAXFAzCskvi3uHkvXf8
XM7dhZqLzEYMXsFg8AtmnOoGORzfC9o7kruJ/4vXqAMmfoFx3odzkkR3PGBC7PxI
Cx26k24wRuQFGH6P3opSoHOv9tpUuzccIeragYoFn8j51FwU8ouXcs2+2VQJp2Nr
USyU/aa44GVjMAd11YPRbwXrcz4D7paY2dqLzha5RYbzznjYHzwsZij9rXO4uogY
M+Bs9767GDpNcqXsSGDKMwTspPdQmK6NWreaRU0t2kxwnbwRebLIgy6dXswIvcAB
5fGT5i8Yao6EI0KmrS69Pu/uq4/SDpXYzTE17XS7Eqjop/THSqfTxuCbwfWnG3t5
4YwPyLrUVI1hVQHr+7mWufefSem1/UUKwZyinabxQs5+xEKSNESTQH/7lam95fTS
NvU/xJxo8PfPMQ6EyFouse/sBr3Q0XKFgZuEmlqZS5scXLRQABPbGUEAIdQYHlzL
qNa1br48Ba4iaATydjNc35fZEzNDBWyYnEM7bh8p5DfW8m2y4fAok+WUNbuhbPI4
745uqqoAGWyH1QuAhPnb0pS5/QmG2SaIYC6VmfIxxzK2Am4kLwPEcU3QAiZ7WTUY
bTtK2GosPl02XZ419stH8YoUQwSlVXBlnWudDUC8PjubWVhaUh9535SrNlkLgyV0
2NcQ/2LFVVEWMkhkK/9aG0+rWXP3qmBAwpv6kM6jwoPrGhauHDoZ3mznxIamLZY9
YIdt6K0/98a3g0U8O0rQOvvxw1toAR05/7N4L6vBBhKPzCjyGYBD2FYUqlU4IoUq
5oT9OHAkn0awV6dKswQXTqPyifSQyijtINYz75SDnzPdPEHbEFz1lPBLxQ7LGZpj
4WuL4T/cQmwqbAj0Tu7B2I/7QUtrhE9JLyNNiDwF2HowIDoMNgkXtaUkF1HW7VMe
K+cHjFgyiotujCc/7nT/Dh6bStdCusBt+dr/XjZKKTpoprwfiWZ08InwlqQxU95I
zzWmz1ZzZldLGn/OFe9BE9ZHDvadL/JeCDSLHc9cLaXRDunvXL91Z4JSeANPF66r
/6AQBitXMLmovZMB9VotlpEqhaylH23jvgVJF/CZmhcEMaTMzDH2wf/92bef1ZFU
k5OEAxc822aG+YEO1xFE5gZyBR+SXUK1hUiXEAKtFuudZRMk89QKrF6yH/pA8UpH
1PAnhW7TvRLrBX9ChG3wKEDbHeuO+LK1RnKweYnlyvYKIBpsOnRAIpSOEPxx/pbN
1ptOLVu8qRwvXxjUhKbE43/XpijVZDTHhHm0FFEabxRXnMY+WUmN43MWerxhgu6R
d28Q3BG5VB9R8SprK0g7ATQOoNHbV7bD9LwNcfHX5DBWzKmhqooSDKXxCricKcWv
BV1H8Sg7676t75NdeOjV71p/J6onX7KjZ7cXHIFpFOUQ92ahr5/QqVRuCy21BRCI
Rt18EDkNIaAmglg7CEfuOCbrWAMYoCTyDCzPy39vN6PLt37kX9c3a+zGdSyAhc5k
No9Z7DtsuGb+H9z+fGz3tSm1r1//cPAw9fPokgKBIbz7FuxoRNUh2hxOzpE8LxiL
a4jg3UYdJVSht9IlkMo2aABByZKthSWMsd/HB1vDR6d4BE4YkrJobnEVwDiLnq78
qHyjG3wp9sUHLlk0E4QoUjcVf3ZUx/AHD8vnVhu+wubmNWhR6GO2pp6eRshWPeIM
Jof6NFMQlSuZTd5ddw1pK8g9sWdkt4+Nqsy+uyuAKXtqwr+5WjoDliRV2XYTh8SD
DggsvsL1lGuTjepODCz6nT+viHHbdiaTBdkTNoxQvPmlvpQCAZu15GQARHfgeoLn
x65KxlL5EbraRh1se1EGs7U2bJqnL6qunX85cb08RLwythfiXSbPmHVIgV8MeE8i
1iCpVgDqgdDmC7PK4pq14ChIt6Ndx6Uc/dILWh1q5ONf5n7ARlzsJHRk05xCSvIp
N1iwcjmHjQdyVEUED61DGk1h+0l2DTVoTt3Bd1nuwbCofJrw+6Qae1FGVVKLNAUj
Vugt7T5zY11veFON+tNvIS+RnWL0U5RmWhVBjTkE1kzA2cf6nlUJVQ1qJdHJb6JP
pNeaLxtvjLjSKpOXmi8v1tBAekMZZKcQJQcKKVpR29T9OyhXGU4ajs55VvClNEEx
LYsnH/Q+vTRhNb89I5DOsU3QZXrtlpYbzn/beKHV+XUoBZgOTOkpZqdPuCuQw+Xq
bb/DIPyusjzPQEKr1W1oP2SXfG/kN323KuPCven8kRYMyurVqS7WcDIULnAy3Z7f
Cor5gCujMCbjaFnWUxsvspq8sVs2YRj7yUb//4LB57b1ho4jjDo/U6Ggsa7Z8101
5MSVl657VHE60quS+CTOYouW0sw4oam9j9/WVb5/eqOko4oqM6dBoZjSe6PtGdUj
hQMTUfuMOMgbGf44G7eWmzQEv+zLB64KNs33/q1ElSMgpYW9YF9G0fHKtEsnmNbb
3uG1FFFXox2W84K8gRmyBuU4k48xC2Djb/Im0StmXM3yx5EkD6g8kCpB/N6h3MIQ
ivJFPQz2DG3wdsgkIKnM+MKlh2X99bmAfnhNRMTbdQ16O72af5IYP7NQy8QO2X0L
pX7l9VE6sjN14pEeydUEWMa4qUJaDI9VsixQmIxm4v5H3gMwEIlVx3Z4aG29vfs6
t8zUNtW8xMRXx/t0MO3SiwUojIIVR+ypdJQtesFyPi0/t8dQbAOiC24rTDCDeeEN
P4eyuPJbzWXt71oEYYEyHKrqvMAPnJFK92q4mt91KCMK7PkhTG2+M5dEueabOVzi
qVkWvEqvkhnb6/Ld7SB4AFVscGJUmEaKbrZBefuJKKA+mf0GyNDWw0Ai01HEfabG
y120sDqYCGfDBop4bgVcWPbC2OurUgomBPgIsDRe9qeGbjDJ0VDsgw+WMbz5c9N6
Fuo8uaZNDYtJm1aO/Bb1UwFsXvZlwQ+QQUnax7OiwEDIR8kNoHjAYC9qiCjYc7Pl
7WGkFxOC0W8drlbibMFLwm8snqRh5jmdWEEIlNnM7YPebNlDjcpaK1C9KWQOtA/Y
sIyHZDXUWy96pQUUu3EqYd+EwhEGcwm4yfir3LtAqGkkx/hEPAMi0J82f3LDgeay
z71l/HaxO6Yf8xAuC3w2n8f4w1rTaTK0UQR4WaBRl3E1FWjexl0KWnnBRJ04V0VW
524dr++6BOIcD4t79D/9hUxWel12d1cksO/ziy7+NzQaDm4kSYbvpZRQWfO2R7n/
BGKxHlMeFRFVaJWZrzkh/2LMKoUROY/Jw0tfqCoHxsRvwKkr7KfBC7xAlsnbx8dd
M0BoANKUYgI0uXM86FdkKBUzvx1WfzUS0lPoo2s40sBlVb0Qz194CjyXQVebhdHK
YE2DBgQrs7a2hWDetOP7seuJtljdeK844/U8BCKhhqkBfCJY2sJdxz84Mns3y34P
lFFB2w/+0+21DNGZY0ZEU6xVdmPGthaBbBDbrc02xO+ZUVndp7pZl2psCs7PS2MZ
UfAsJ7XT8ew4XoT2wGvoLg/CZoNZxXlP8JMBxFppOkZiilRMgCjU7Sh1PwhTbXvI
hqrcKOgzuCso0ap71W004+Ou7XpWwd9QfTCyJj1jikPRKg+bKPzDGfZBdCijuBiM
eIHKlvNeySdQnn8o+zIdInH1iytR3cfo5F3tFnSzYh0CYLmoGTplYAdiTXgpj0pk
E5lgjcq8TpujllKynHIZpy0aJzyR9Opd+c0NSquGU3w17KmXXEX7GaQtCYPjRPHl
ZksJODOT67tn3EYOY2wYPiLSVvVF5ISQ6KD+/R2fEVNOwmrJlzNmvXol/Mk88dRi
l7iaah2Q0UpUo671Q6klxKr9jF4hyC9Onus+EUIVYszhEHAi0TmbRQlyNhK+jbDD
wdmAqC5DjqOxLMz+deiyX/oCieS5sddmta72TKab7ii2a43dIwkzocgqsxWRA5jo
ehCPqZYmWJ9LECfohq3tsBHP6+rpYLJJYHJu+rZSJJnhkuH+r9UpE9r/982l1RS9
M2f1ICMpdNhSzDUUdNmp8Uxpagv3H9cCSnoyw6Ye8+a2yX2JUrbFVl1kRSLxdHD6
DUGMXlGRulJvoceKkpYCni10qiGmyXzqx978mEsZc/DZg+KG/jh7DsmYwgSeqixB
J9ukRp47A3FN+er2uaVUBg5sB8lZmxrCMiwiahU1rnbI/JXxw6BMh6tRFMyPMhcH
CG8ny+LDPwaQ14pCRd9IC5XB0x6Ary2lRPytHrS0Q73FJTT/EMpXtoDn9ItyF6pE
ZT28fQSAcxG53s1YiKS6lyOoUZdcScc+K8jkFat1QNZ1zs/1U8zBSMJHJVahpC/I
rla9VC9vmARlSCz45z6S3cpZIAZxHaUx+EyRHLqBhwlzsZFRYsAEngFpPsIsxp5b
843tgzgpehUORJUxPZ/r1QxP/q4jaS64gcwaxlbKbDhwTp2Aj6Or09FESbWsXfZO
qpLVgOMEVO8I0FOtNb3dhEIlQ2Y1CbSSexezGtoXUvpF7rlN71gk/c70f8C2WbvP
jZ0qqixl+XutsnQMqALogW/94TMlv5mdKq5nXWkFC77tbj9gSQgrnVk28PsK4Npb
N6LCZ47QijRAEZPFiQsA26o8mkL5yov2MaxtwqVu7QFAbjmHTT8t2e/8WrhEXVtL
strLaIOzQvlX3U6+vxUKY44fNu1A3aovSPjWNrngsv6QdOaDf7fCid21Fg46bwcS
MtJ8uUCAKr9o85zVcX65erOLiXSBS5IxIumnq7Jc9uJtIn4/Dn1UllrkBCZSw5Zb
jedvpwiqPt7EP1b7/uUTBGN2GVDcKNvkPq0bKXe+U4XmI3xLbdffCvgGc2/+iX5N
Fas4xS/jVfyuyaxCaVVP42X5XaItfCG7DSRxn4ikcytdhriAI+XHz4VKd6K7/kJn
uZfAX8rhJkY3zHjNobz4J5So3fBj9elT0hZG0dguGzJpwYROxS0A3EF9NfP/zNcX
Z4DseCHwergs33F5R6V5CcLMVpheIdoIlQqpPqWFyym0vuJWVB4GMyS/jXXulO1m
8GlhaKa/zuAUCRs8wRkhk1ZBaH/eZfqi5keapKzWOhvMR6emeeu2FUNO9KMYsX7u
9nD/dqUWGmubPhW6r+rCZBoFcL314rp+8lA0pVjr+cCsJ2r8pSAEUIDaLYIevaRY
GP5OACcIc7lGTwQm0OSbtDQGMENziHmms/igeRv5AsOmkIsTvlxcZ6KhP3rBua0P
A4jAcCiyXpbmuGLOCT1YscXmgXkgdpUykQeio9BU6VFkyiqUuGmXEIZGdZSL7Ea0
2ZXdXbPrNgIFAwR7Jujb22txCgLk0t0OHC9DukM7038fiWxDiI9EF3fBDvOot3WH
55P9vE0zSzGgOswrN5eViJrBUv2Px6puiDXRejjHpIer8YwFhkm+LzqyeVKEnsF7
pfRX/XQYdmkGf46A6xtAoyAyh6LLssRfage0WQ47XT/UalPkyULBic8rA4A9ZW7W
GvEnT4v23ecAUvKrADQ51ENiGSBP8A0Dtl8GbDhB/YPe2jBXCV/9VZv2fUQ7eRe/
xb9tX5Gt4xJUrtb0N6yAICrpYWvb2youa5jFp9pjkfYCRYYGWuTnIitrIpBA9PUg
pttrrkJ/LEU/agjHcr+z3+twsiBNlF/+9A5b+eKsOXkYhIdhBjTBUF0GrZSeHQ9q
5qxc+ijCQyePcPDtqmOfHl75d5MGOdrXWryivv2Zcy1S7pdgfFcJ0ziuclSZxu5U
5iqJG13Pj26aWDZiLCtKfh7rr3yQiO1d9dG5zCPWPW185MCp4/YNAeHBMpKp7n8l
nWJyxPcpSiysLA4Q+RClulGjS53FfBTXaCKo4vlUgLrRhTK8opo2g2U/AwC34RoW
1/L6jMGKSU3g4yKFq1CAjVL2QuF3uCYgBNUOe7t/kwZ5+bZA0cYpQ/AOMBnWhcOY
8M68HUfN93k/hZSbZlm2KA2rozKhgeSR3q5tKLYHdG+ktoPbiHWlBEceuF+pVXzy
l2/tGWX+W4rnhuZNSPELWvvihqfZVebYJhNgxJUmY1Gru2JiDtZRcvbl+lT3ey2f
QkA1ZVdKS3K7YopKNuTNXPKO7oJ3vW5geHkV+TDv38c0NyufnyVdiYlfHCzTg1YQ
3cP2ToYfy2tbqllGjMZZUPVgefAJbgcrh1OPilW4BHpOvLGH/wJCmwjqfpFb8WKk
ZawdIr1699u6Fde0Scw5HDNEKWyTFNAWO3SGQNVOBQzvOElbRDXb8oSS0jJGC/iw
MhJmjDBts5RVb0/whnngQIS4mVqtwo5uQgLtQk/PCBuKFgBJGLuhUx11h0toUZ6H
hED9k4SSpuAFrmhlQFE5bRbBTAC1LDOJoVVC3GmCTyTITLNKzySAWUkKvflqiWCQ
9zhgFoIj7LXnDnmL4/UhGxy0u6odJGbpC386EQQYFXNar1DIMVjRIBzSllxois82
sfiolB0BKP3s+qmi3gd3Rbw40KLLOOyA5qx6kROQnpP4mMT1z+Js+deReMVLPTsh
f5DNdfVZn7/Ee+d7pHWp3EC/jQVrweT1NM2YbtOWrmsjMME+MJaFluEuCfsUm7Qw
rvDskVfeQS4CIUjspspoPPJQhFBuZMk5EBVJQBgdXQu1W9VoJwAF9L7I5WuQg1yx
w/rrEAoL+kyidl/YM0ND6FOf4L0Ia64jXFxhrYz0dXsoKSsGGVy00J86Gv31A1g4
DrJDnx2155fvZyKOi3Pq4z7DGBxDwNC+E18uougxOkWkqU2PhfrZIkNhvZ5YYV3/
iVX5Twq8LZ6ilBnzYnOmIwECimTGezz7A7kFKiIm82cw7xgOF0i9A6y9t5TjjiYd
Ut80SBDOoPaWqLCGErHWmvW8m0VUGs+SMojeju/Xy0YLmpERkk27CIpGHHAPnucI
Y8GelxX2DZFcsRWnb5H1aYEULw8zLAt1JqPNmEuCo9Oi804cnrOq11JSFxcm4/md
40CgP84U3kZJqoryQPyAWu5yE1jml4tFxNyJeMghQbNCpC9ngE2NO6oL6+SPpa4+
QIZrjgfOlOrdXpk7twz4FUkXffgp1VfOiko9btzueHXzb3e1GYU2s4s87K+fC5ip
1wJ9I9jLKVpoFQcXmFHO7afr8KzlMNRZwC2O7Gpknj6wA+MUXWXRS29miQJMcpcD
t+22s2Er5aLKdeO5ZD89ZQsV5xSnPypTsuZKDSnAfLVVKNZn1uDfg8Zhyv8bBpPx
u3h94gMKn7VMcLqaJ5SbqKBmHIJ+9EtOX8qaLuU9EJGug8SgN+MNjglp3MKBN8Vm
FQGs5I2TDjkSjFZmqXfpTZCZD1/YsoCbSm7ysFowXk+p8bwjU2FaUEKqqnYH/Gls
LNYmIQB+KkaLwvRsHTL8X4okT+R7sAzCa1UBaYU+d5XBra8YYVOphA3IhIESKn1O
FjIjdsurZBmGVYmNJis2G9cs8Pcv1gZFXTTH/wMc7GwmJDm0kYDRVu1gR5DVSF57
hKC2Xp2OeAg6gm4ALtdELYVrNHt5JZ2oIEUz9JZ+kVxm3Fzqf5LeE40EFZu2Vr6V
d7VOzG0+oMCqXlLztUPGOK/zRi51ECbAXhpxB4KCqZcPLERS68RpE8YFW8bMrrvg
xIQvbKAJUsjSbySbeU32SmuulxIIfi25+KolljyQ9mkeFM+n1ljJkwkC6y0qGrZP
O0Ytue42wOMuOHs/f/pxoHhHX4nMa86eQFcnrfYq/KaDWX4XZsfMbXEQxybKux8S
Wlpa8WAFMMiOXPLmYpPT7b7GNPoygqxh+IUzJAZj0TRiZny1q3XcQClNsytAKR73
fFYdFmfcx0ttLSazmuch4rSF0Tt5dutSG5Mf8Al77kesYDWtQXWJjyuVnq/b59Ow
ne8/K0SkHOItk2+475InKX45lbHFDLM0hUinLiXRAxZtyMY8vRFwK+IRk7mxk9e/
ttGAz77dmy/WG/9rL2thOLd/ZFHXX7SQPL/LDxGMHVS53QRr3kydS7H5li/Hxnnc
cYijOhNnWHkOu+Jox3Xd2yvI+5jk2xm/N/CS8mggfXYe6XEUNlYcAFMvZAIbdZ9n
GrNouhm535erVA04NHHialypVdWSZo9lJVxnUjj7aXSbl1jDhzvXTlBRc253EXqk
+R37c6VZ8jGePm/YhuIIOhCncv0ny5PQIt37See3ST/ANro+1aJNAD1BMghByKwy
FJdAAIh6orgWu7cTWHB5MwNt2wsgQU5gXogJvM0zBGfdHx+qfJ1iTdzcwnT1M2SI
USXxIlgp69jLb0MzkggcwK3ABgOtfye4icF2frRhmtdiBq/5+UohJvTCiP6nr/DD
+Ngqa7hF/PE+cVR2O0xMn4Fk+kASgBpNTvsz9Kq8wEENHoSLITn6QtgGVAQVY5uc
EflbVtpPlWUsIJEUrl/HUJQMSyeU9yIj6w6AHCSIr0ZFomv2PhftuW4WnT0sEGvh
JsNiYOxwdADHakIrduwdtomz/FXsPUOoxzo1UH1b2pK52eRJ+zu4+QL2U1Lht7EH
AYwLFOrLaVXkrHUXQoMUERKO27JPDLAcRYv61Y1SHSKmm7AU86EkX2E8IRuRvRR6
v74Ulj5tRph6uhqDlRbAhM/iAl9nbdE7u2bmB7CndxcsIwcvWYCnE6XQbzipoLvB
DLbBMC4MUIvK4ZKXWZxF42x6bY9NQ7sZd2UHlaBa7v5/wsj+f2wIEmAGpZ1xmjQx
6wBiKX88l2R8+z0+vuoq/rwHQVjuhpycdh3wAEZ7TIB6TJ3km/fAdFGSiVr9h+Is
Zj4XbeWb/obCxTowzbZUt74OEzyPoPP/4BZd89MyWtN3gPuMclgWX8OXol5MEFMx
bPS1y0W0hcaoY9Z7iJpJCJIFB/WNTqQOseLdbHvtw0HLw+b4h4gw0tVjCyFYWbW7
xz8Nq206DaV5kHax8WZbOaBNWiTxqoylnmbwlZ+hW14OwT05D5IdMTZpD7BaNj78
ORYNYyycfQ/tIdfuJDJWwE0X7uaXWb/VnTEHjPtvtkEPfCP9MOYiJf+SEVm11cyg
8lg2ujczbVaAyDDtBq+wAZ653uOML0sGlPrYe/sk6Z15XrLRlpcIp6LWykHg22CU
Tsxq5Js5FWf7mwzEGciYbc6QNSKjAPuCy58CjuNllRc3PK7LgIM1Sobucnsdu5aG
ebgUE0u886oqWqUC14tnHtSGGgLS36z0hstw1R9LGejFZ3TcNwX4FdqaS12CD+yr
hBPVH2DvB7ZsMnnf8pAG1PWpwvF3KOPW21sFyyMB1cho43+LDrGcnpGAV/V62Djr
8IdjC2xkt9es4Mo+udtO7pgM2b7Jw1RrI9G+B5PqNxsbfO1mtOCG9Mf0A5gRgF/x
e3Ily2ZKqvI2nCxQ1rTJF2I+cMshcgBjgrpXGwqXJiQwaDgd89SoZ7ZG5Zyogywi
TLHj9Cj6Rg7X2t9SzL3d6Md5APDNtEocwFe6ry/AmYePY2eVbyEbImvxgdGrFF5Q
Xr/wfPEfX/+JSGDA7ztFw8JvS1yje6J/Uj7UHSlDBNdKjdVMHWumDxDP/yfGUaLs
osHn2/SGdVX09KJeCpHuhCcHHtOqj3gsUsr3ArF5ZMjzV0I2ms87cESGzn48rYqg
vZCoYg0kDQokDjMKUgVOdpaY7VqhnblNtGucIZr+rrsHbH1fCwoPSyq+3LXalwjX
1H8xTkXakcvjmdtANjfmjA03AyqISiphi3M9+rzyKvdqpIBv/9DguJoBm/ceWGu5
/RPcNzUnKJHZaZXMHb0gHtwOOMSV/lFOE7yzWlUUv9t+/g2sXVy1202WYuFAFxbZ
+655GpMgfimKJAjGrM2K/tFkMNAXz2rJA0TYbR1Tqy7stVlpz3XTaDvKb7QBAXgq
Dhanp9UVQ6QKwobTdn8eG+aN8g3h10kI6tQS+SUi5B7wt8lbToXuAEcYLc+O0LhK
XkWapCAxOhxyKKrIQpTiphVKPX3DYJVPyIFlVbgUfPgirQGsyoMpkqa8O1ARTtNC
PW2yitB3I5yqX6KL+XQW7v212/YfuXwUgQ5C5+1Srz8znkivBOEkXJF+tFpX9b23
4EVFpi8Dy9xYqMErdr/oRqQVU5JnNYJ46nFTmAo9B1OlO4hE8BvFHnCaJ+VSw92T
eTn3Z9M6bxy9IR7w8jUGcC2tb/rvHAbHkMYz3Os+5Z/bld6g7/QzA5cxAx94NegN
MCpO2HtRVWxCGHB8+JQMPGhMbNuhVrmuAIyz2DjQVF1WCI/229CZMFasaPYn0JDt
4d3kuZdz6FEUaBetvs/CJlf7WpqFMcPZSP/4ZGAFPLB6y8m9RUo5d92idhgQ0PBe
ug/DMdjxVzYhYE91ExYvAVzu0McShXzafCBxvoK/VBjlyWeUEbTL6mwmmcfsBfVL
6DkLmSaxOfQy29zyQ2JjFQS79IfmAZu1iBWv+DuyVN5aoUw/PR4cEcWnYu5eG+7H
5vXswOvI1IgqahLPJvEFWUlDaAhYxYSk2YOas1dTcoSJ8P3irKOi05mpyaeKIoT2
zPLIe9fIBQwuufusi7z04qfTgkh+ehcbJ1LvJAaST9A2N+TJnZPg3zL86iji9jq7
sckAQsc0a/HM1MBKhj6FcBVuERnIRJZl2bmAYHdkMfX0qIEvKfK+5RfDZZccMR4s
y0gV6cSJpVNRhuAYsgOcs7Rn3u1Ust9FWexb3VWRNFJGNO7fSBz4t/YiPUxBYNjK
G0Y36UGIRzFJIrKHVd1CdtJGJKta7eXBOJLw8ehUxMAB3ks2PeOi8NsVHG0UhHSF
zTw1MIY59BW8u29qVibsTNapdNTITx215jpPukgKFnMASjUzifT+Yavv/lYF8Pft
/wHmm8fj2RaUSDBTfXDic0ri5daaH4HF3lzbpbOcOee3uVRaTLcsRwdREYCYlXy4
z9FTkWlh/88fzFuWgO8T13AV2bJSSDuVwfQW98A1gwll5/WQSTrgNiNq+sE3NHEj
B/fgl/hES3EJqC6LFZqNRN+fjNjIND2Wd8L6jZj8TJsl8BVvjW6qKpU9bJxi2bj8
4xUXlSdwYiGiKZNhfxHy3Uyi9krCgmqvb4J2vEyhcgOpNy1DZr/ESoDT2eojkXJi
qz/TF2drRGhsauUCdB0bbs7ExdJhHExH0e3+16SZ7rhHDuGuuUE08UNuK/xTyEtj
Dg6FJq7IV/ctugMfxPkZxQKREZXTXwmPSUgXtcqgJ/UVuR4RCcDIWaR4wnyhxiaI
oNYEkRtp+LZ9H6q2BOYxoMlcdcEh7LygAQHDFyhoZDC5q2UdBUZQuL16/sbDfVFX
7tQ9q/HnmxUw4qWIosgNDKospIEJY7dknhksS1poqE6dGTTEd/G6szLRENSbWll6
D10njaSLCR4wyXx3LH3xuf/toEZ8hRO1ZDxypCgn3wP/jd5cyrZRMZguM/2xjGg+
oaoPndv9eK9cXP0VexFHtcjTHkWJdqFHhEkfjSQi6P0gOaMigqxjachpchGl0Okd
hDdvEu2fvNIrlFkXdktubNOTA775CHXd4QDZhjhNllH2xB8zv5k9tHfwmS7OspNr
jC4sCz+ZbADvKgDSAz8EzpdYCGzQTmc6JfMuABwI3ecz3KViodd1wmSe6cpxHD+m
Boj2fuo379FojImjU+9AMoW8pk8UZUkY4gsNvBDNIjAuDut/5j+h5WzefX2/GT5u
3eZpQDYP2K2BBoQTnh1/ckm0kHo1eJ9R2XROvdMCOkIm1Wt5tbyMAtN9ZCxA6Gvr
9lacQu2nT0erKAFG0vtyokW3DZdTt2SGUYn0znlSSc4Qlo/9KxIAkFIFNQqWyZRa
JH9rkDkNBZsQ/pQUetHgMTeUhtoHQei7RKNVuKkNQsOcnegcglcSdq9bh/AoJ9ed
ki1ZETwavW3xJFCVZr1lqWKUSfFDzfnK3oLIRya9ddX6y7C4SBDTS0126fl4+eaX
CuiKJPHsGVzhrGXI8nBO53C7SMctvYPzAbXh4bFuZo2zcHDSZ9YX5q65WMqVd9DK
PbJ9iW5g+58zMqRYnkBwu10PB5xqk2MRBI5fr6CdjNLAFOywAg7R5c6SVRAXv5CD
P2MVQ/+9HbaZUIu+ASvYEwH5APZ4XbjEZ6I/V8xm0NCMcqVFiFNSSPSNTTBe0cuQ
7/t3EmtBiVFBWQNS37uLa+7ZOY8dxb/5aBPqzKcvjbNJ6VSavQFmpQJMgQiILEkW
MGU2pamPwbDIDkZkgO8F2FaQ72y/dGG3suBD4sOiynmdW3uoug9lLbR4sEm2tdwr
uasIQ5ebavqgDi6baovmERfqSNdoJWItVHluM+aA5maDN3APhU0fSTJLVNVg3EcT
V5K8V2l7ZGU2mNIN+bVivdhCl9/K2pE2pYcwoTPKhGL8rNK9GxONfSPqhBFF2PeB
LJrunxpsAHgtfd1bs52Yp+19rXlfR1VwJEHVZhQRWtGDwHIzU88XaRXWq096Zae2
xuvkO7nTjJ6Je3qs/3rITNuGnU5W1RahLNvbVx8PBXRZgXGjt+o/mF8gIp2LPA2u
oVkmg3JpN2H//mJVEz8qscQOHQVo6E7O66vLK1xd3y1K6PqgJoEdwQCevABSNR7M
ZqCYWtUS3gHIMV44Uwi7cwVziYg4ntYApH4Dvij2EtH9RkbHnTmHbsK7rk3PKOIW
fXvSvCT/CicAWCX3JpdKYwX+MMpKcGx/RAAod+wmJd0sOA7PmXQ0XnSOlz14p1i/
DbrtxJ9VP5fqqti71do3YUq39d81YoaMLDwA99sFk4TRsdh6qBpTMSG6HLJYNRZr
rUbRZ0b4nzsin5f//ZJRjjFn/cOIIaPIthBFwzxfbk+/0NCNKl4CT2zOQxgYDJrt
YadQ4nvo7J8bqjx8rNIoqmqbg7C4kjbIaxDqNnyIc5RHUNmOj9qyWW2JqV9rgjSY
Ej7PcFfSAzdjecPqeA+Q62+ekzpYmhRPnFYzMxGuw5KC8qetI0gl5s0ELmpjojzJ
yMNmLYw5s/Db826+DYgnkuFNNLNly2pwsXlXKnp7NsAYR5vab4OGeAXAgXoDwAtI
3Fodhjm4W6Ix02i5fPKGRehhWld0+6bqvjYhhPb1+8o+wuZ0/pHfwposqeRZgRqs
cG9t4f82xhLpkZCfO6JZwCIO+Wm4ro6hUXJ8AlA/ERLSUB7Xm/g1Mx7xSZK4aDlc
2rasUvkfPpX+q8Jti0ngtmM483dcHiEiKnJXPKMSUOzYLnR7DBddbR4n0YamiPd1
ebpmsXdCBqIFLt1AxPOFTXwFHZzk3ZFOY956C1TSr1DFmbk047ptNGjvQqIpwZ2y
WPOFy7JHt0WAviZEN90mkHFC7hapzlSk0Fp+d1t5d47SSkQcU5RWu5mlY3eSyvyH
Y51Cye1hMeLAa68G7QfOruXyH1C7kNkc46ZJkXkcmKB3V4jWS4Gipt6xrYvqhYmH
pTFglTSPPHgWA0QXtCmb8KsNmbifCwUL+U1sKdl9y1qCSHV9GZ9dVdz7BywUppmq
swsciPXzecGthKqR1fptdBuKP0O/O26O5ditMrqc9OCZRahrH+5FOR34Neu3sK1N
Sczp3+6lYqWxqi8pQV/QCNakytl3SgBe8TE/FBbnsdhne8MQ3hcRZyGXZcwBG/to
LcN7c9Iej97a99LNlbygXa/URkPRl7KX4ZzLa0kQmzAYgKspxDsn+Vl2ebOvuU2X
7X8W/5LbMIpgdICTtMpCuh9gTrZpn8Y1ChCQPGlUgVqim2sdMxzDL11pRH2dMUBK
fnl3Y0UkMchRAoAG1UtrpRxtZK5JJYnARGjxkSjQk9dH0MlzFQERVXodxaDX2GwG
7+igsbB4utkEHWEES1gK3ti5vNRwHtPZIA0ftMU1GjwUyd2RcCSuenaoT2niIDhH
9i6jpBOyHvDfszya82M9KPJgrVQrXyL6cd7I5qzSqtGgysEa5uqKE0DXa97gsu1z
4JQ7PzcR1tndfqLGUCz7i076kOPJSfAl38kRPH5upoc/4Z8gye+2RTvzyFhDMU+g
+RFeo4tBYq4EMQdjOKdKyz7Fm6sqFpu3AB/oCaVGMZMpTJXg66aNaikQW1eKmeJL
1dcDdYvOEgTv2RnLc9ryR2vpdvszZ7+D+Q35uzDlU8+K+E4T7KNr9D7G5176XOwU
VsKHhtXrA5pQkqj0EuzHid/R6hrvGpYDC9w909KOkbI9uYTi6a8HtDY6+kwW/zm1
UrE5bvHaoWe8j8qVZ4Smuagc+SyYR6Af5w+45OyTb0GaFYYiBlPAJGsQXtnlZLI7
QFdeK7MKaVFpnEgU6dFy39YOBll2H+hSnx0D9oRefwt/9yjIze2/x+pV56weuw1+
9lrE1aOYRUvPlv1X4jZ0snnOcy4C46j4grB9DpVNlrkEyUdh4/urhbDd1+DMsig2
RYA9/uOldaClh2EXXeHLIBp1sIi7bjssmhGgg3X97V1QH3KoL0LuuVxrwaH1cCs0
4dfgnqWihzacIVf8jkZ1Q4aHJltFD3NLhF2DnI5XP19oYWxAnyGv3rEKf5ziPgou
AZQl/Q737pey4zeX9IAlOde2HnZDQshsu7G13qb0dr9nTSCW5V5ojjnUFBnRGUKY
lUte5FUrctX834BEk/2XOYnNDpK2vbBnqIGMk81EbSCd58UHxf4waIIL1XyiWK7/
erHmajuMigavbCnuHwkk6DL2FULMwG0II/OZXwfEAaTh3lbVW+oegVXso0JxBn+S
vFsuyDEF2FTpEfIaPHDYhrxr+baQy3gOgaJPLXx4JoQDT8Aqg6pgNF1OKnye5ceD
UZy4cIml5rIe7F9wlAStfAPOUNkcZISEwLxEjLXl1n3UhqBlrDjfo3bqNPQQCrtC
6rx2PZOa0MPFWmoa/OudG7A6KT8pxwr55KlxrQheGG1H4Z7uvqUAh+aBNSCLjwAf
cLEO0Mo5oAmFwZWla2PeYwOIYwZ+2Zog6Qj884LXftqiQMhjnt6hj4hQ/0irNPSN
50kla1mTw64kaY0wI2vKcz18XbH9ZFiJsF7+SydBna4NqAEorzcctf7absL8AH8L
75Bs8gUbYHAogPOYqQBZCsAV90cVGHcfbKKj2j2CBH1caV2kPTUel93rohTOk75e
mawLJhfMbfBjjs4Ql1i6W+yDSuyj3/DIYccHSad4oSrVTP8p9jtGwVkocuWtkl5h
a7OaC3d8Yp+qOV2d6t1UNtqs/RxAtfAZR735id69ZZlEQAmmQY4PXNWEditRWFP9
Nacf6qmj1WJqHPkBWN/Y3397ABVg8kVQB0FmoH5JDGIGPxIoN6FibDOVCDLabYYe
5VNN2BOS6Ksyn0XDkA1qhp1R11akoxeIuPmEYM0GlVPOPA8G9xCHWeYmrUC7vdgC
wuBukTjFGuzEluS3pm+pHVMSE9TGLTTGE7zItITZGL7DAfzrjJej4RvAej7/C7QY
Hfju9bvYyZLEg84sEicgv5IAxfRBwekFwXvL3ly0x78tFS46fWuNwgittzKeab3e
U0/KY2KHhhvRuaEJ48mG1Jr5JHufMTS6zpwPb0FbC+zlXc1OVdzC0xhBjK5OH0dO
mRZMFoP1L+x8E0j5oREGk9pACpLGcWluG8WQoPCx/8fStwRmOXS9WgwYEM98GP7z
hD5shQaZ8aDMRy6IKzQH4KnbaC/KAjJ0ddBrWFGjp/CdjzguJoNYMCqB5cITy04S
r69YaL9oyyJUxUr1kUmKNXtytU93ky95wgLRtGWgdIt0+DKyV0v2hqqHC7rqsDv6
rreXc8RVB6z/rSJUc6gPbQISxpW66sLJEbfeOlW45cneGdMMvIVF2QbvzOs9lQiZ
F3qVhAhO4e6knQR3oEMK1LB1QvEjGeiKrNudS64JH/xBXTlp15YQKg6hy7kWByAi
JKyjGR+XwPIKbfghGAv+RiNeVNJCPGYUcI8ZaxwllifElsKWJ1VbYh6eRlHxaml5
WtlSUI/yl3CWC7llHktoP2t1tqzO+0/0RxZT3IK4gisoDxzdCjEscEMhn5o9AUaA
E3EBOxLncUFidtpmq94+ZaNzDGOTSJlOXkCjGZbnyrBVnGQEIpA2rbQK77HljYSO
5AGV5zoj9Tgz2OYlAHucLnwCeIUDn9qZh/n2oa/I2ZCSzCiDYoQCNigg1VyCyyi3
W3Q/G+K6lJCcWvbPb7h0pL2HUWpbwEgrHt2y5+46Ai0n4anWit1SfZYLtycmGhiX
5JLfrGHAYmCRBHVVhmztyBj/DzK6XeWr8NmL26nPhQoh+r0hDd5menxU7WR/z6I8
pVSlSkcXvLa7DLQMnXW5Z7xrd1yyWdDztm+tjiojZl5v9XCWbDjvRzvYjKW1NR8E
0+4bonG5euwX02tUX/JN3rAIoh+pMhePbBupXOrpcpqj+7nzlxyNJL82ikPcaomm
efbc9UfYK0bBou4Hy6RlieHb7C18TIl9cllAXxLUh228HPkJkkLDdHRzuOlk0FSO
4/WfF0yDKulu5e2CrbT8aYBwG5s+y38A5n164IomWkCcaanXqY+5dj2NRWlVZnd4
e80dvmCReQsrDJTR57MAkKMlYWGhOQo4Pu6fxhlfMGtq1tTpZuzeHUgSlBvDA2Ym
6w9meeCqTDkvzfebSZdqAXDxEx9moeApbRDIz1b87TaNe7KeMy6S1QXZ64Jwv9q2
yFzDn9xWlkUt2+p8Yq9yz5Wk5aoZ1QVVBlIjsdqcrD4dgXB+gV8UEJGX0l43MUbN
xDJkA3XzZhKI6PNS2aZTYwgJ30N7QWXT615XOG63kyH547EzLsWuQ2Bl8t1MUlhb
7NyFU5FKco5DzawQnBObeekLJFC4q9Uo8wQeWVIK6LzyGK52PAWZ4AuAp2oyVUVa
DwHrNhUPE5pbBLAGssIyneekogYPskWHkZwjA58POv8/IXz/QZM8SA/vygfO/fKK
j0d8NhkUFG/PY3pTt3H7An0y394UXEwRDSDETkQ0eDVi5OYBLtCTnkIc/PrsVXUl
2bs2f15WSFfOrc0tq1pRPeMAUjucoGvbvxZ63PV40DnQN/p/+CFsH5/28eBwM6dh
GPg0pmpYPPSJcLFFkj27YwHp+0v3tSu1tjNSmLIIhJk6q8J5IyZKJ/i3/1qZ/xS+
7gN9FMemVOdeTgw0AdH9tXw82jpyLlld0oaPV+Ti2/bQiZZFlUpRo251w6ESKfjm
lQxvepDuMIy7m5SrlA2Fm4CYivBQrvupZ5nrrynY/2n0Ny6kbtcEstghmlqq5sZS
5O6j56NfMKPSRU7RqZA+KpZn61GrJ8tpNcjgPuFnIXuZUnfgB1DQxEPOzwlIn+CA
WtiIt0eAIg19Tz7NQGytcQsZvfQ9gby5zFfym1oqqIx4AiQQqZqU69CgH51VOM9w
oDTEK7NWxmcfQseTALCqRVvaMLjRWQzkBsDzvoFpOEB/dcnwQGYI4zaqFmO625ar
bRHqnxpvE9eJU6P1vPAWWCc/nH6knIwzm/j9c5KZzRK1THo4Md1RbepWanWrTS4A
IzMNtoANQjauWvnmDeWBbwx/L3nq8WYF2FR42Xzu48TQVN1Yi56AADzJFO2255+Y
QgrJcI2Vw4MRBiZyCodrKUtQCENIKgP54Sjz3wEo7ZNbTn3TBrg9mMepfoe09kjK
/bvf8gtKWHJKfpyEIVkAXFDyxB3XWaSmqK29PgtVl4DCxAYGMJf+RB70pB14buAg
6C0DWTe60crrAhK7QxuHotdqpYgaoIEvuuSNNXpDDef7tyKfT20UEOlJN004zeFI
TBnu0huJRGLFcKNPDBhiZmBvj7EJPOvoj9gKWd5J+ngrh0o4YwUNZzW0W9PRDgMj
1kc3+5ADV+NM4ZQKvCTgw1Zib+1D8O4M5Kv0Y5VT4gOYOQSL+3jX99QXCvdVNaJA
iC2M/Pf8aL1Vmv0nTkItwaLwY4cmTDRRAi/ewNJfz42cCfHIPUN4uSlG2AfFfMKM
Rk3Np4R0dboG6OqIdWp5XZZuIxa7B6xFYoLpSrv4mKg4+TXRHyCkKe4TA6o7GfcC
MLtagZ6mkl/KEB4aoLt32Z3mbqzu1Y7ocAgQrPaskQyHXwfNlrpM0iw6hFDVRHCF
Iy2XYvb5lzjqM3G0pE7jJYDC3+bHMj8sc8UcRaw0AtPLljQsdMJ/LVtmIOMfwIlG
3+1fQc5HW0NQP9CT7gOOiq0xk/TNJFvfnUreLZ6XWRBiPRlLGtkXvIMxwK8/2Su1
JFSest74ZhKBwji5ZLkrDCVqD0Ts76mOKfUI9ASAHJI7DG9s12n7D44EKzFx9eK+
VX3jC6D5KVaUSAStLSS+IV05sa4cdla3uZXXdsX772DFhLzCMZgpXnL1UsGaUt+3
k+QZFV2madT2qrtbK0C2MhNtrd1kGd5mWuTfk7Y9xtL1fpxtTakqkse2XBresCzj
s30+/gNlwA1rix0Gv025NP2fdnOuj69ZyjzjBQFUGY3Rva1O9HOI0QhBU+6jtN4K
a2b64MnpijqQ/Yb6OuHiHRXT9wwCFgoDhl6YsktZBPh2+3tGAGQyX1IyqhWz8/hX
fjTKDeVsRyQyh/m8mzu6WxF9rnfUzVKXjPDbg9sENJJbRVMYgsmdZnlbnjehLr6n
CPSwAOOo0NNf/gSCa+cR1bGxLQbQQnbcpndiF+2EJkGVRc3FUbJv5pphxnbRQjk1
jagvBy5hdx6lIsH/vcww7wDEBAIH6qIjvcxu+uRKQU3sFcKS6ygGgBfPj9B+iVQr
U/j5lHfn4NWa8hfnNjxND6qI6vYeJb98yO93Ih7nH9SgGxQHcgJyCT/+DUTqlS8D
AbfK63Tgd93F1aI3Y/pkmQS4YzWyFttV4KQVgBF888jMuZo2H64XKzIRGo8bDOh1
1EdXXzjBQJzk+Xznv9feeV4RFwaqLUkZDLZqs2thLMnq+hDlktxROHJ53KA3Qiqv
Hp23TtKKnLKKb2BCuMWoV9ZSiVGTGUwo1Mc5+QIMvfwFdxlP52oaV8alG71E6sFs
hjLtVDWqeg7se46LiOh+mSlVJVFB5iO6cof91iaX6yhMTCEv795bMge6o+lBQEDx
ZtXTkXpsy99HTbTLCJdp1bWZlcT84d8L5QwpuJ4QnGSm7/J/WyJfYyETp058uaEm
16Xa7KaLLFvkq0ZdodRYkBSfZsnwd72AXm7q9tpqN74D8DmqlvEd6mVco92yk0Vn
luZGsjPKX0PWGTRBpWIhjlzuqZDo82eTYJu4N04eXTZgYKOjCN0Il7uYazFUs4MP
9azCCx61fUH1ShygK8i4W9p9j1pNsnxfXOd8B4CmAd0Zpkp+c1EtgZJME7bKoQF6
ueoJXRCgL4h8/mLVkFCimOhzrGhrYjOOAXazYtpMKIsiEGYtAzfPjN9bGSuZDt69
h/aCWjZeO81ADrI86N7xA11zN3tADQ38hvNLWwVcwHJTtmL+nlgAQbiz+7R/EtDf
SlVyaLMcHALkwSshSUzTcxmKrzsH74ao+kFhDgYxQ5zK5etHkW2c5chH5JcUv5aU
JpZCpyqe5OPm94go4wrMAC0ZdY/T0Jw2QW404dvLebh/xAKnJo8Df3jz1OrwWAKK
0NXgtZzsGZyf7IJOmEhtgvoUN2Y07pjlGslh3L4JGhIWyw5GeQT632o53mX+fe/t
Sw52VRAUt2hjfghZ29q/DARHTuA96eZSWJsS4xZOYyAGtbLbLm32p8wbSmBcjrmt
9G4+nO/d9vgvOzJ/UU7+qE/tnGks/QJUU1cUDOzmGnyNA8QtijKhYHjuMZxe5UID
aviE4SWeQCy8GOlCZrv2hlnKrDT5gDCXIrGs07oezyzZ2ntkChObbAgU1322tCbA
dssrMpoUZ/v1XRK/P7aKyhZBKsSP4YZeDzLVFdZor+zaO9EB6expttxqJ3POTmGr
w4WumwNRqNYY5TYinDyaaP/4C7w7WoQpOflyM2N4eVrGpP1+mdypZPbCufksetzM
DyCjPbYBggUPhoga+luQMnjAjmCYHYWCVN1OMk5SK46uGjL6J3VsN8bu1BfP5npt
CdO9UNLvBMNEyZQ88CSbjm4GgYhvM2je8v1f2+RX13eorTf0R4yvnn+ceg49dW6W
OuTc+3LBCwL0gcm8YvsWXS+q5qhYBtWiyP++0c58tKeFBJaPsjgZnb+KetRgtYok
r4NkHBxlyNkbwwdHXGTB+g0lOnXnoPu37AZgH3U3/RM9rSQ/5WQlw9veHahxOUYX
VvQ/3OqHnIIK4OJsMm6lplg6wIEQsxN+K7X65VMkfClwis3WhltufJ7zSp1TUI/8
+Sbb5K43xVLaWkZvxcWyKfHRtFvC3tQ96XHRLNUfL8jQwUti34QwwxVviKLvE3Vc
hShJAqGeMyW1rTdwCLAwxg1n02SmbA46zickEr1Z+tuioS/8HQeMdemJU9ywPWWO
rqMPZirAEa5zMeVXLaWzwiymUIMtUSxlkceM9KEj4M3VWCH1O/SwMGSDYrQuWh6p
ENFWqfhGjU09kwsvJkh9bOqU8FQDFBgvI5Qv0Cws0NGyIxC1wc/prrtFiFwCgGFl
AgFcFX9DCfxLIM3cNlZahbSeAwmo7vYJap9kq+TFfFKvdGZYTqhXeg0CYKnTlwyq
EOgXVBzDBXcRDfEMYvXYz/wjRgs4F6tCfAj3oVGE+ZBhJakvdVUjCjqxEB9XbDpt
6xARdxeF9c6W27bYUnkY0S7BXDJdVyk3gNnoeB0P2gB2WFBXyb7+1yKjQUgq7NLy
5JerKSKT6DA0VSj0TlWuKY/g4QB7aoAVF40xBPySRCSV5yIfVM0ThKyb4J2F1+5y
Qc+B3snBRjVQTwE1fM3mSpSCl3hy9YIOc6FO/mXWGH4UYQ5/O1b4J1DAuqEhh+4w
+TOqZBLWAN6DynT8B23uiezY1JHY+9RdR1054YKtufsJX7x+Hdd0UuTHBABbJRW5
KlCD2jvjSwFQ1oSc+L27Gm7OC7AzCC0CheRoWdFY6Cl29DnSFcWEotZBazAmr7td
lko3MRCWo7obA1g5RMrkMe390Tw8p0rUSnrsQmy9ntY/+X6xGhXfr6fZGj4O2Fmw
uMuaj+oRE5ii40xQ5VAPuiGqMKWiyRsFGdFp3xR30JyzWg77NieZz4rUi9pEBQGi
Rah0kQVsz4m3MG8DIjXgCCL6HZcZxz7tv9yZklrEPu9O46u1wm9lldLMkwE5/uAM
eKr+vQldh77C3zpGB4mX3iMiPoOgJc6571NswpBpFHXdfofbxbUXhsCl4b8TnAJt
9S8Vs05EVjxRxhtT6qeWqnbDIWzgjWWdPKvsTi2iwKQFOjhk9AjXfTzvKhx7eX0A
MRQSwpibjNm/Tniu40WGjjvvUI9SbfG78KY8P3zarAz3YWvl4LvAFKeGA/KxmOHa
rRnKwnlwhWWOLf4ZIF1MkJgTggHwfXC64Ag+W/nGDHz1YsqsQu0odNKBABjx9mt6
o3bxM27Cx8ksEtJXBrtUIGqGJflhhsJqmmJRTxzSwLMdgTO7MtM1og7rhs6LrbPu
5cQvwQk1+CAZKYuxuCrmad3aCbaEb9VnHawpacWRbjOcTkwUoLQ9MbkrRAIX7GpD
KEflxTfq8/SlvjY0s0BdrURY+Bz3YuaI3/4JV3R2U7QmqY645X6/N8RZo/fhcoJv
fZ08JowcpLjBkcJQ8cTeaYfWISP5yCoJ782e7HhY3m/WXqpSUcfGPKwYPZSrbnEr
ugl8f2AuuWYutJlBEXpRwgyBvn4zrhedIpKfMnr5MHG+yN01+sbPGOsWJMa8KGAB
reJvvGuKGqyLHrU8bjqjci+0jky847kYXtMDj5PZ4ISLgkot5UPP68mnYGcKvR+a
NYGgiL9d7G5aoafvFKLtQTm2IUYlrOnWhpJiJ7GHBUpgdXmQ+7kkEra1gzTxRkYw
2hGJvfkzw0kQ8mAdPwIIakbSeoBqu6Nb8S92Bd5iUFpNE25OtQbmmFltAHxX1u7d
CtcAW7zA+wtxUigPWEzQObWGpn1Os5tNl7KIv7ej0VN0ifQ1mV9i2IkJKdzJlZIY
ntdpqySvzsOF1VpwBw3c6ryLjLuaSHBLBEiko8ZjEtSMeCSPiUn/y5966YDI9Rn2
+AS4xnkW7RPobwC1gRmCr5rlZBX0p0DHNMnrsUVPsJ++DBzvZA5PC/2uBG7k/RN0
+wyiH7KUKKbp2oMAlcJ8ji5iG137+wkno250VXIKN9ZXHd5DllwlSEK1CDaWPdXs
wFlY5oQyNB/X7wFlVRI1KXx2GN7HcOOP+63Z+6KpI49ewMKjgG+De+kKy+AN66Lv
BBdFsnGKrgP2oO7pUEb95eCNEsjbCwJKN+JL5QaWmvF7Lfj20DgKqYOEFkbEb+P7
On2qmLcbJye2BC221WLY1CuZNy/xjpwdY73QXNIsiiHKUzQNgSIWhE1ntRv5Vclf
eyWcVl6FnIrDm+V+90bskHyAYBCquqxRux2kjsEOiN/j1HVRMcVo2RnNapQy1/ia
duZbxjsQ6uJWq515fz8+F49VHKKiinpkF2MNlXl1cDH31WV3t8vIZprJVVlP2IqW
IhJo5KftRLZwmX4ze1ABjy5l4fHsYO9BAdOrME4F13DeaBh+xW6RYG7brgMdIeQ9
CbFmxk3qF4fhAwFpYp1MMOMDrSdNA5tJNZaNz+awC4Iy+xrr89qIcbari8Dpk7zJ
IPrVzQh/woyDQBVVbY92q0Jlo2ZVT4Sp3DwGdaQDHUZwC65VLgiYs8NDhIMuiJjZ
+Lg5akwP3olU/mqLcwZU8ZmqiqKWIk8xAD+b8B5o2SAbOl8yIkWW5oaru2ZHDqc0
CxpGv4gR+Y+cwPSRkZ+jxi9fisgxnIXr03zeFpyaTA73SRi2h7yBko5Sa04OoiJT
W+98CIISn+Z6/dPx+VQ4/Iog6MialQkLOdPs3fZ1YvWUUxJEN2LIsstm1crDpfx0
srvA8tofkS8Ernog8Ip6L+F4SABzX/xINgi6mFVznogv2oF1jGrfFRSC10Z9URJ6
i1R38y56rEt+GphrrshEE5D8IAN+uOxLDJo5f3BnUhyD+g6bwixLh++PLbPp8MdB
IM3LfX7E5lVlGkn09i+bLyzKQz4tG5MokiBk5jKMvTKPHs8nfUWTlglJv7CTNXtK
GhYQgbxsoPqlU7oqCZSdn4xXG/snwX5ekkP7o20MXIrc3dXvT3WWVttmphFfY4/7
OAjDvTCMNgl90kXvbPNTw8wyeiP38z3MqNcJRcJTYN8/M0a4kR1THRQLsUcLNwAz
eeBNeeY9j73gd7yHLnhFBCLtv5zk6lmuDtex0exs8aDu4u2VEI8HdZxkjt4zjTPW
SAJwG9ouScYddOz5srYrTwp8V0CwmtwncZMe+LPVpu1mCySh7quVExIHTMxu0uro
LjsvStm/tV/X8xSSVIR3i07MaTfih+QBraJnAqqprSc7FVxhkcjfP7TXkXHGlyHi
PMrdeIsj/xoEGypL9h3J8g5if/mcjg7R4N7fPzxAyAnc0s5Y04vT+dn4171u7iFe
/ZRbF8DnaVl442Mrlm53M//NHYULHQVZEdaRDPh0WQmxQX4mn+k7v0gOeMA8L2ge
v+ZDHJfWNKJw2KQQYFhdWMhtR/6q+/ZgN4Dbw6hnGlQ2afG8BWYQpWz7pHaR8W09
I+nmHLW8gbua/B1da1VgsdKOrR9jQka3VlxjZy7QCLv5jHnnYC5x4+8v3nuY3htn
xnb0nIeGjcRD747CDjmNvh68C5BCOkSBJfEd+BxUCXqiiQi09V0NjwsAhaXQAN25
yatIyh92pOv42dJyx4SUkYQWIIWVhhtfBHAkn/BkcKccXS+b+Ud+g620IdDuUAkU
TmlpzKAOOLNol57Ctmyc6uIDiTk7IKPsLbgnoN+B8A8QWWd3rwRyzWjbuu7nhMGQ
gHAnFGJCZ21wTHrxlXh3d6Cz1zQVATVOGeR3ke7RCNW9PEAAag+8LWAIuL1Wajj6
3k9sdFNWFltC7Eo/E18nds7ni6JLm/+0ZAdV8SJyQCKCs/HorQYnqhrd3LGG1Dv8
SKC8LDE+cZYxzCh57s5vEhTbeCGxjMFOWJ3WJR5IR0mU4y1vIxwnLd6lRf11xt8N
qN/Nu5YDb0h+k8qBHSpuVMnkjqBtZOaNy3KpD9wmtTyaXDSSa67wGZy8SRr0DML3
2ynQKgufe9XbtLDSCjfmW53XMiZ83foSRomBCpBvdrZpqFGYVbj+DDhuNUAHtE2X
1ioGPKj1keCcFMGyMeweYUDiEdttgwJwz8rgZkvnViWlYHzz2SPId+lnvgFA9nws
lz1Wa5gjGockRagvpVUFtcCclW+FB7KTeIYL4g0kzP2gXFHFgszpi0e9k66CqoHc
QsI1Rp4hCzwzGozpXcVOFw/se8bf7WYaH40d8C4Jmk9E2dTX5JvnyRFuD0Ai9p9e
QLiPDV+b2Pg8nOmXgwhOhGbrnJckDzTTdGeNBXhQr8wuLfKHbYGruwTSSHpTK3J5
5NiD9rRhN9zxgS0wUFJGdauKAmHCb4SeNm7eS6Y2Q/pzliCqODF+2LB7Ce9iHRGL
8apu3jfAe5K6++kVtfUmJvYPeqjg9mSaxaw08MtbFNU8JE6exhwLYziIOMGYJpmQ
Ttw/YpeE+7mfeSlZ0hUpcThGOf515ge7abhxOLccdR6MJ8nzWcj/GSJS9VASk2Jk
4iAGee+x2Kh0mtAFfSRN6LtEtzBe01l5VFWJGQikvMHUC5WzSXMzdWUFMcZHuJAG
F/s/yCui7k9R6TbsFTgOkk+Qxmuq2eAUpuejPM48DNt7n0vATgBGXLjx5+JLGr6A
fqEiHJ1wg2Tiwd7UiC6AtuoaQQ/Lrue0fvTv+4bogNqmUCHNwtvJrjxf0wBZ5z4b
sp5D0rZlpOKBh7Lm4xHkKtcmjbJropRfO1VI0uzudnQ+XuMiH/4ho8fzpEKWiqgO
HbrxPtLBZNmX2fi/ZEc6+SZ/6D81R3O2WXdBu724JIXmyhyRS3kNYk3Cq589dH+B
i4+yh+u58jHU0zCJI0UIpn4qpgW/Td4XN4/WXTFO2CnEYfZCC00g6O5UhW2LD5Hg
JRZFZwviTzSH8o8zsyELjPJTQeDBhA9Bo53eiIIZO2Aql2rGTrr3diPGgacqYSA4
UNwtKHsKRm3Ii1Fr5+DiMSPZBd6TzeJKFKw9lpr3r/Kx13Nxmm5oBfzdOkF1nFvk
95G3grLtNCnHMMiexyiFCkcUgob7Ikm83NPYula/IHOiMZ8oHr+b/r3zTDazEGaB
j2d96begufpYOb9DVNgAHUFEtTh8sDDXGn+a86AL3Zq2PUCqv/MFEkh+bVgWYzKH
AgQOQ1C7+CUCQ1E620HYKNKsyFrhlWjQ7vMXx4rP5WWF9CTUh+QFX8ze60ayxAEm
aC2qOWPZr5pkYUZxOcBZSfCgWCCJ85UH6PqDfo/XqnA/LehQV4RV8efbG37rdS/F
lOt24gcQVEGu6oxAAP+LVCjhISMpGCHkM+CIQbY0gdxbF5n6hESTxydRebqA6UjN
fzuKSGU6YBPXCdnN9MAZzBNVGMBSKVFmQvRUbk9cms067rKUeZXAaP0d0DQ+u8e+
2mG2udlfD8TVh8LFitgtgIK6uDnIDI0+T0a2ttmccshgJvw+vcYLGDE4XJe7BjsH
lHv1lH3pK1CWp9Ch+5bMq76G8N9jrq4OxjZdRguDpjbBOPO+XyquB+VF9epwwwg8
kI6Qs1s9wbfd65CpbgzCn//N33FyaGNM1wREmsY/cSIWLrZre+hMOZPtaWqSdoLw
hcX6wPV6MsnLpaQrmcf96pNwkM8Ai8Vn+N36qCmCGQumJGC6ZcxczFSMHlsY/+Uq
7eJELTkG51G5nu3kqdQvFj5MaikEnaCDlLCB7EDN1mOhD45c9hQbwyRJ33YlamYa
jgk+haVxM8e29ul/ep8IlyMGkIGruX6Z9syEcvdMJy6O6bJHstP4q1TqnQ4Zz8/C
gD4DAx+fKeXKhL/BPOtqoNXontb+oSJtsIxlPGHOKA8OpzMbztYAM5VFLS66o7uD
nk33iNUmHwSIBzYJxJ/haZN3SYSnT9dE4VAmEXbvYCXAXg2yLx6vr7lRdRcmNYH7
HUJFBFHVb06NBosrc9GL5bM809F3ZLBgqGc8zp56bz+uYgnhLmGxbD5xlACQytv+
FEp/g8YURi/hAgJ3IWLjPR1DGwxUS8YT14EhRKGWCy347DnihJKxsIDkOlUhVxCt
dh8kOSOvLdmxKHC5Ui/r7DU9MYldOu95P9NlHkjQyrTpzoemJYUipSKAtldVvBKi
5oreKqVXWC4J349IX0jbaKqvSqNzWRHJXsIBI0aAyoq9rH/R2GzCQqqY46tsoBAB
dG795EutM10wX27xdZ5MU0z4HZ16ZCIHWpA/taohvZPPN0JFINJ14c17UEluKLSY
Kp7Vvg748z9cSh2eucedGx6dC1x7nptt5SrN8NXouY/xwts60Pxo2hmBTQWQRWQU
CeitTPuKloHccZxGry1IB7zm38nUjULkRFmIW3i4qKpkT8i3JAh8c8+/td2QVVaK
m3B43ZgQIeEj9m4HGwAOwe1AHc7yHH0x+ycZN6vDhIJ3/o6kM7kz+czsAHlUoaBN
s4zIzqOR54xfaAE5clpeC05EiGbLZg6HlolumdO40aWIrZ/T2i/ob8Jt9fNneRU2
pkBpJyVB33vSMIJPDKN2ojMtTh07NBwT0A50q5AtjTHDrqzzY8w6YRpbKXcLDTSw
rDRJrSsjv06Pcv2/GFvutuSgZzQTAY4FtTAliJO+28xTEfN1tDvaE10cFnDmsZ+z
BWlpPSu4vNuJc1HwWAym0BarwmxcI/gP1tqmSNjhjRUvy9BgVS7mvSzGlPhEEcmA
/wHY8aEOa1Mn84DGKESNK6yUxAXIDAyzf8Gobuz7KXEW5TB0YRBN2/jDkUn62And
yYnL2NpQT7MyzUYzb5hrqthp5JqSp9IeDOLEeHyFHO0vopl2+M/ntjTQ5mR2iVIJ
SB2rneMRuFKpIFIQq/JHNHsPhDG7UeiRA15OuBIQIfA2+RHqh6T4bkurVli3rYg6
ptTcBPKy3mBd+jq3IomqWFS0Ir0hSt9XueoEFnKdifQPkpWfcHDymd0y0JQcrXi+
lGbQTbkO8l5RAFFuN4vQJjo+DYgktnqR9RpaRe+8C8aDwC5UiNDli92BXaNTu/7R
m+tSM7zbaAT+GsHpcQ4gAVUSq54mD2AAwJlyX6WchwYCaS3wPiawjf1xpqMWEsJh
M8/yI5vuFv8xiS9sr90ygVv/pm5KF1wBUzz459sJKUd6rrx0kV8F9oz5djVpMBSx
oy7KJn4+sPdSPxJmmj5he7izKzwT8C06uy6QYrsw6uk+GYT29ZUrYTloUGQUOnF7
p2M6046tTi4L4qvmKSJnIggKQnY0jCsoeOQZSFviFpG2TckkxMGpK2Swdj/5q3uy
d9EN8PbQytNImXYI1qAIsdLg65+rGJKkoi6nBxQbLu66SMyy0kaB5OyqlhfvMuWo
r7NnJv9qr74AwwJvVAMroURpku6wK5LSfP1O1Kk1UbR6sH4XYIC0pYX2cnq/T+jX
IyAo0ci1fKpCAgOeeFQ3SzRQe0w//RQMeGFAFejY/W9eJL3dMsgrUzqyBAyzIC+1
6gM0HuS9yGTgrwwpzdSz05ZH2dn5we0gOB73jbAc2+NTOwSKiarmQl25nJzPEoD1
g/cWX9sEWqSadBzQJupqRLS2tGJAU6tJiykinSMtk9qvz+0gDn6KyiYYcCPP6/3e
gKrtk06R92DQzbAUrXNjKsYZtfHpMait4RcmEOwmJm3WElDfm+iJos/1MBABeavu
00b1psZVPP5O2/i5RkrMU9XicSu7rN1+x0vE+Bx1GhfKq8f63aYryn3m7AHPZNm3
6+w7BciVuNU8NctvL31bordDBBKYcZc0WRoiayR8vuanp0A8qK3JCdXemqk5KwGd
YJ1pYBqdPFwlHRKSyNwJa21ZcLIqWlz5N4spiS5a4drSicnD+EjbMcc4oDKUTBBr
SRyaV3Zx6hq3UHSzdkn/8sKknp8/6xcf/M3Ejncfr4cKdYJ3HNGxwj4sNM0oe1Ey
trjCaBqmaXbfW8OEHi4Nd80bkvnGdeJ9crVqSh+OujKAncqn/EZM4rLk7om2PYT6
WCMGdWAEPJ6mOqMlotYj5HNwscxY/VIYzh08ZBOuUphxarthP0nsL/1TccyyHsKS
r+A5FlEa4UnuI/9o1GZ2ANkEHmTjW5EEhFscB3yxEjrHDZrTuhAcdi4AoQEWOwKh
Iz/NByB0aZNv+kcfe7DsV1WVsCjxWK+aGnC60dtvOagNyr2AICYmi6H3DmYxA2GV
XyqCUpjZCBNDzAk9tihSqRf4nv1yCFIpvNWxxf28Kaf7VtGRHfwipdZTsOdQDJkp
ZZS3hW6OKOI+MbILW91DNPUqy8G8qajTUnohEaH2EqoHNPKnqdvwa4gGpMSIN7xX
/MvvNwyjRcLlpApQWN3aAB4P/USPqpLqSni5VNwRkaw7NKSXDlXr7Xd93eM3tGvt
ZLKdBM8TA73HY2iMm78DswxzHV78DMywPtz27/2rE5h8BynzFdMpbjG+1knPZJ6T
r732zjPDwjqhI6oPzx3qWK8BqQHU8pbsi9Ut2VuvASG+zBeb+p9jei65ishjjs9k
24Eq46WmiuGqDvCof0IQEJDjAJplF7Ds3Wc6ad8yAfrUZzKoQclc4WC8MZ+EctC/
A8w5HVFTtt/bweKDJoRoxurz4m5GM6I642NINJ6RPvMNmnABv83Y51sW649Avt7Z
oqYLe2GvkTPyUohXP+kHhAJs2kh+k9QG84/mZtH0d0/0mR4rvyxlJ9hHthTcmZv4
0jLYJXXM/ao3Osbh26DU++Wu0hvr4kLzwNTRz2WchsuqJgLEcoMuQQV6XqX0E1Jp
bTaceNTPzPJEgH0X6SqjoDBh3cYp0VQWJwGn4+cuFb4suz0sCfC8tK4o+2xhB6tA
ZFysnrEfIsUsFNifd/azucduwcFXoVqJnLbrK3LF/P44cz74/WFImF8x9PyuzAvv
EjiQ58rRfYerSwiFDLS2EoTAkipAIy95wgzG5XZQ/LtAj38TQEACo3Hh61Jw1uL9
wTp6MDn/CyeyUWiB4FCH78WNyO+coljY5lY8nMnDaqgbc6dWEIlscqL2T0Nh1VST
Wg0DfmR9ceTmzzaMdGy6i64LwyhNwkMbjdE5bI0x0raVs8itmo9tJ6y/Da7xUByE
TtorPgqw6YGCgcV9urbOQmCZZAN/4566adFFkwDxsFWlHr4fmGnsNqa6UUL0JMio
0waLOvxA5C55Qasw/XhMeg3A3as1QYRB412UqK30IydsOfj78zSf9kgtrvgOjU0u
+8SQqdTP+hfX93YrEV/ESbqRW7y20XhkCMtt8P2nARXzfp3Wu9ejRVLQfkw0aBn9
ycWHaCs47nOW7yQDc2zxFb4SWqMJB/fU1ZrQmz5eaCsnOP1H6k7lhYXcuUWevkUj
fZ3LkKJ92MdbTu3Gvdz5YqIXE0v4HUy+aYebpQ9qdqIzlGWe1+mQjF3du9KoAZi+
fG3wPR3UbZCuPU6uyWL5JkZ4DTA2g1t2VCEbHptl5wmAj726XwmQGnNneO/fQIap
qnBSWTCOLc+6aPcZZAc2KdqlslMO6PNhF4Vi2WjmNkPFb1H8vSWfRxjlEWNM9Bb7
qBYVdBKUdRP+7FIfJGGI4Mz1XKTC0gYwIEu14+SBQePLfg2BaWoaS730HrU9WDQz
XpSb057+pw+HTYDr84Yku4qL3noOukchoBUH3iZR/9lHICDEZ0S++qpQVOjz9ZLP
GOGMRimDBcmD+FNDdnUKT4tIMiloazs+gZFXI6KCuZr7/BbKKtLBKidxFJwiPhZl
CrV8AQLET601CPYGjQEFEn03dBJ+3P61b7N+eMkJaoJmnh8DDdxysyUrqXlws9Ip
8mP7Jr8k0MZFqxLErwbH0H+ZEOfisVBy0SX6UpQxnrjCG2JkbwHmOltK8oeZuWwC
hoGXIkbDxD5ZagF7Tea0qpavVkdDaoagWxKA2Mf9S3K5toWCe5DT4+fKeTNXZiqq
QnxvwTXbZRPDuA1Le7D2ym3TIxYuadmwp353ZWoVZQHf+b2s5c2uS/HCpSMPxuLT
YnnqZ18jnwDjWGCmbqaINuC/Ruj9pKvjMXWCBzB5u/sLK4tA8UzfRDSGhCd53xTM
eqaZRk7+l4BVpzrxneZFX5b6etWr6/Taivn8vvFIHFp7W5t8rmS5cMb2mVeLHy6d
+WYGV+SYC5bsJScAs0ahE37Pdp2YAQuRLi+hKEcsf1rS4eaMex328bRvCUH5d0je
tPS/swvKNrvcVwmiuCzGsVkFXpOy0aX1cKYF1avnXh6wlwIC7ZE5RLlnYFxSK91X
4qOMKe8KHraJW41+3sM1oMsbvtuEf91vM50+lG2gg1KfvT7LPuHyKsjnSY4Bl2gB
LJeI2/uH7v5guBULYDm1dAMkdtZUpb4Hyf9qTsbiM+DeI/ZkLxcycVzYP9IAMYQb
c92aaIqBBLUWGdSmqX3H6ziUoxofb8+uhvi1/TcXxICZNE218Mb22WkXTzA2iqNV
LeK+IkMP7F0kK1KEWA6cF0S4mHLwvX/+oN8VXF/whOxkKqNAKrkIji97XBPs+ONc
ULZwsjEGWFSBBAWViXGnuwu7q7YN8o4qblfTzRo7uPIZ/z1u1vvBTaYiE3lWbraS
hXsI5jUktISS0zp5H8hDuw+YCT3PD8gJ6QVihxsiBHrkmziObgb3yWtLPqje0H69
IlIa1aiCPFvXUIwbWKWoJOzgWbN2jk2Ti4jP4RLT0mqICuGDcn51bJ1UNPVABm8z
RUV+RtT4w4VVG3UNeEPd+q+igTwVUHgNJY2X2p930hXhDkcnF5X1MZg+2fUEMsPV
bD5WejMvD7gALoVRaTjRBfQfr4Jzj4Oy+Fm9gg3knwNmSopZHaRwFhNZMaFl/l9i
HWbZk56nkDHTk9kga7ZiCoCiSSXA973z52swgWt9MHjqem3SHn96QsvnwPYe55XA
kMgOGP9qnnSeh2+8VeVgiQo9PnDQPSqBf1biL1AyWEuM1dp9Mc6Y/HzMxqAQyhEX
M/BUbMY6HvOFnFiBKCZtsyNxTn4+NDUYn2VTD7zF0RDRy0VrlIUtzedJOIatefx2
E4gIqc2xqRYDEg4WIuA815+eF6wJye28WOHbb4pk/PPNAh7n89DWNkzPT/Eec5hq
gGlZ1se13ILELfZv673MhbiOVnuO1tJXoHPx7tLyew/5qO/U15CTRxVzNu5Z5qxU
M8qk4oiZyF9Ruqeqwut5SM1ACnZyuLW+bp/KNyXH46BSZx6UxYNK3NYy9rp0kQk0
NYYIGeLFjpdjRIla8hwCtvqurLkFzZhdP1LNzh69HD/oohe3/eUpcVMygcQEePIG
GV1273GMNNQ3xksSKJn0YZ9rkq+0todneOx4g8+2Vb9/Uk0LasZDvGzYE9C0xncQ
d5t9QiLEIQjRC7QqW4L7xPlTLvXZxS/Mypq+CmsxyGlLKg1l/tPJ+i7ahRh1yt9G
OCXgMArTDcT4w7ad17+wEeUcQrQrZ/A7h6rlEc0x1ONEHYE2IK2+rfiAThU9uPDZ
TjTmIN4niB5AmSmxehjlE9kmp/FZNfLsoQalW7xIfigWoKDerGehfBv9ng6UEBNY
Bw3YXOz5Lzbcp24fr0NuSs0bs/U7qfTPK527dJiEp80SgBMscop8LHSIW4gT9QD/
gv8n4x7vfV96oRjlhBWdYPXu+hRqYI2BKms8juzPUP30LebiFSW3lbwVIM+VbQ84
5Q5F+5oUSlVfw5GL0ON1iT1E8L4nZfHexjXmv+bVazsKcSUJtPYoDhYUOso9FEIr
FYDzLjTo96d4zYKaNWtYeCcYRlgfGMPs5hXLlrAUby7d40CgepSavqe8SSehsX3b
tZOauLQt5IMeg7TAWS9RYcZUtZt+xHRGW649jxblNFrp/6HslNjx0OFgFBimnr5K
9M7hjvf77XCzkDbuF2+gWAPaKPb8QHXhBXxauypxgMdiPLT7vTxDatLaUP4bqUor
3MiS7mMptEqRGRd4tGcl0CrvwxL0AmrSIrhjmAUlkPiBX/U0/K3IYWfUFk7nnGHA
7nM3tUqUZ4XUH4Xnh9gPXXwl5EAwpsaR7J/FLVVQ4izXz+VcD2aRUzKATeBIVavL
gsZg0c5spQu8Yjzn/Vju54O7thzsz97PMOx2fLgsTBHFzE4zssv6mTfQ04rNPq2V
EM/xGws8g7PgH1glrnWyzISi69qPTjPA0WeKnsids/xXUpWoZ+ETKDOWVqN4DnUx
yxbmnbk4Zp2rkyIhbIXVIA/DMT8PTq+D8RB3WzAWbOAHel9UqtxXA2AlhBC0XCQ+
caMAjL0hc5nid7PV1TMCTEug0scsy1aMvHlDUkD8bJDQpRqz8vrbxIAGnabmWT4F
jTtMKZuz1cfpylZMzR0IbXT5gi7XDWM/esqIlAlPuaPI8LQkUb+yNhJ3PrYewfhx
a8MaVLvzqavRu31/Fd0DnceffiiK5/7vCJTB4Ygcrs5Qca1jAnBUym/kp2+1pcG+
eUlUAm94Vcs7vS0b4YKSPjfC6iFH/IEdScCdA+ZaQGmtN5juAeLXvKy0yjivQ8UU
aSUUG71ZXIYN/XezVNKG45nU3u4wJZi9SSuHEqNeXsdYF4td7/93wBLkaFFC5IuD
W0ozXFH2yTMGjtgV71linqJUV4GEyT/kvkGT+JCbdlEz/dEj6iw3YaJwLwlWW5A6
AMqdMEFoKmTLkN1lDiFD0GYEuamyZGfswSr0G2sBpjSqbVCZ8fbVfwObE7zsmUJu
5wQpq+eIQxlZiIVzxPiRlFOG4VcApMnIV3y7c3N4ROvUeBF93eCAVGIXK5GPfQti
hruCsIMrgJS/bU4x8l8d4gMVdQbCknXZ9LBBJprQaCv/d35xm6GJeE1BNtu36SvJ
2wD2TGB13AxyJr/DJn/Hg+/6WfrBjISP8n1dbZ/qtG1HblaXevdvH3trGcw1HEr8
H3PoXw2B5JFJwEQHr8LqwHqFZ41jghnPOiWh8VdEGmH47m4TAP5pa1ITdU1g+0UE
G087njqCa/uGEbgWBYpjh3kW1uEuu0AQRVnEp/WFNQkN2v0IMK7ymBKrBhGg9+4+
DIh2ybIN2Hufwyg9y9T/gha+pe4keY0M1XmlxRURkfG/jwLGDP3e7y9LZuarzWz5
nRwk8Vi8dw3svmXTTneLrGuF0+8KB+M9bVagozXvDDtFyOyC5l1KToJgJewcAMYv
TtkMcV8CF9C48kOAeZq1bi2pwCPZkkf/0Bto43CfJyMILDdhfpKUfcmLitK9r7/e
QEg72SP0/kawR6Yi7izIySLiE9lWZ6YQImAJN3I0nzVkeJ95qeeEKKeICe7y8/vM
17YN0pJm22VDzFMYD+ie0zheNM0gAz2jJCShslSQhDe1kEbAO1sRkbeOuX6mHzpU
ES/eKoUsBRB1Xn23kmK7+5lraaz8cEoQJQ2bCP99J+VNMKfP6STsKAIDT+I5w+Mh
3JbzjMnC7KAlBNpKii/y7JV2nz9KvhBj7KMRLb6vpwZ+wzCJv/B+/EPvtHWVufLg
/eZaBEpCZKdR+Eksg6hihrGSaZt7677uowupaFYk1bUcs+xYUq7M8cStg8VEnqqq
SZFAwUJ13/WTkc8DNekBa1EzMwiQuvO5QXcvbvg2LrS5Xt9yvXxedkHk5l2NJHUC
H8BR7wA0rA6isirYtuuAVq9cjWNr4BlRYwR56nYTmDRj7VW3vrDw1Hl/ZTO6erTf
REvVnf3oa3InO++VCi6L7spMLtE3cQiML1SUEge+bWmFOA0CPS6SBEjLLF2PCG3M
WejE0w0Q988g13SVVm67J/kdqAEFKGR8Rc8eB5OXEnr0fy2jC5ri+khN+hHBK3D9
nwIvUhiimRzu+JiTMPdc+h1l+4cJes90QtiGgDYaj6E2D4YHOakw9MGqfPQE/a62
QQEMB6iq9AkKPXejX9fdHePcocoiy/glhjkD+NB2aqdWC09meri0dEcGGI66N3md
5nj9I+qO45ckHQtd6PDzAcGelkJOOonexHb5m9CO2RWMxgRH5WbgLBlqpoFuAGio
/0EmMFxGhJ2K8ejrvLrS38GYQiamErOm5nlGSKuZjyMwfAbrFY4pugRcbdG77gX5
zwdTzYfH1sQ/Vgv/W8NbdSX5K4f+WGzGJ/HyKSwsrl98CsVqG6U36l8NJLegv3/5
53q9QJhoBGR0abCklUOpVZXc7UM1MpLOPK2boOc0DGMzQqDS2meidt1G6cHV8VTE
D9RFuNwInLaYomkPUWEb+GCDbJfbC7LlTCnVGKdyVMjlkcDOzLGBLlJQWwWmeS7S
BbU49evYAOr6VugLnMmUDg+5mICZziVv3dhKVcRHpdiKfQkkuAVnP/bmBtGwyW71
9fhJaNEORe3zmZktUO+Hi6CqxWbcbRtxebBlpr4VJ+MygVKlpC5GFkOSs2W1HeW+
OXW5UBIYirEUTBdZZu1InHOVDYq3rLOUPk2/3Py5kURSSGvFbHeZLjSiLx0TEjkY
x4Qp5J8y7k5hPFP3ljNjQlj+KUnxYe5GzhGX/x1gD+O5xL3dORNVDhIWw+7AlOgn
7/49heDUFwc0M85kejna/wF04O0DBuIzv0nxZ3p/JqF9yNWMIOm1WE8fHUO0rOFx
xWGVOCGdEnS5ucus1z5m1V4/YzeOS1ruwfysKzJF0gCWck4SnqYrjrG0/tDrIpDa
OEbyQ+2ImunmfT6cusWl2P7Om9yghc3DO5iYRUJb3gMmHcYP9Kcfoigy+mMxDr32
DBUW0qxuSHIJUcf/gdcnM/J0IG2B/VszSU9FY6HRGQdIgQIWn0ED6xyK19mxI74n
l4Nutg7oXi58+6KDh501JMZzSXCjAeUB1CmwDP9aAm/Noyh67R0ZwGGJkjbDcKow
poBsF3ji32ctUbHKznQ9bt4q2zEAp3758/PsBYtVVdYnSxxC0k9lxy3QHmYAZwuF
QDyebOLoTyT7wkpemq5eCX9lPH3X8elErRfzxDrOBNRZr9/1dDcaGgfJjQynKQs1
5UUaVRGoLI7LbO+4XIUUl5D/zBPitac01KB0MzurfnhSBzglyMN0FQmlRplwYS1G
gFT1JItIOLf2HMGsdSTSFihPVKu2i9jNtWpjdPFn5IHI9IJHDXe+1h2d/PQ7wm+H
iw4q5ej9Yuxyo+pkJqMHB46Cvvb+yRNRF3Wrdt5GxY7t6WibiZeVSX6r+6CFKN4U
vl319fGXnzuj4LZ1Z27T1V80aRF8GrovkTEZBFaXJ0Go+Lu/ebWxWhXixPMuT505
MD+WwtHgGtRHRdcdPH0V3KbqXqSuMzhiK9lvdO7IaCr+OdWTpfUXFmK7vQ40AM+k
vpSmj/IVjhVA84JtrM7j14X3aOtFTu8rTJwephb9RLW1iR9lkQNGE+F91kNIVZSC
8ayOt1W2MyT8Frd0JyPdJ5c2z3RadwrUbDl6hKZ2PFj6rna5Ax1z631+8zCloXlp
reEPbLv+d4WUAaV6xNaftTlijpLKJNVpviPfakQ89ddV/03/iz86eatnknrrvvKR
YBhTQ8G4d/00QX/byZwnzKT989RKi6tCIYvUgSoDLdB9Rb8X38gwmLVgBo+tPA/4
AxBNTJs27Syw3SazWPuMQm69YJnBIs1dkRFh6TZprNFnY4+xwt0L0tyC5FSMG6FL
uM2qFtUzYQMFb0w35GZm0b1aKP9PcnaROLBgbmdYx5WPElenB33kfYVFCM9usR1c
hfjHJEK1/RtMG1OL2aAJH62pxArkNccc/zDVV41d0/wVEX8XWWq+KB3BbxyaytaW
VymNWF66yf6pilPFvcuEK6ybN9ze6e15cV9jeOF8OEh2w3p2ocsbTJLvTVqvmqBk
Y21ZCg4SrDBJI8wUQlB2jS5QOzQ8tV6DTF7dT4g9M0hs31feChsUNyBiWhcxpLza
gwk7PVLE8bex0y4d9Zw+AFSRVnOlX5vyi4afrG/VG1Zb4rJ+KDqApTsr9o+nzWG3
55QUBdiWksPNxiOEA+pvJLC4wkyQq9qQXP00glO103jqKGyb9jKJWaHgIw/CTH3v
8yPyQrQ9QT9BttCJcT1G0pEVp+P/7IC/sKmUpmObQYT/MKX9GjR8vOQi2Pe89nxP
dXNEv09HLoGXKJh9XH47v0bHxf/0RDQ8yBkQRc4pdmXS7g5VS8UKotEauJc1kX4r
NR5xTCY48YRNnTG/AFO+vh4G8P22L4hksbW/A0bqru2b6elYUjEvs+HfagirORrF
oKsLK6rdSpcuHk6n3G0hUYmxGsFp3VDheP9IyFycwPi5bAow+iuiyheqQ3+yQQUo
DbxdhNtKzpqyF4N6JinNpSyZ3N6Aq6Dg3wy9ChHM9Jn+T6glC2iLKANKsq/7Sy7W
4kwuNg7w5avweYSt5gafqDGKCJMRzS8nTMqHxSWtT3DlNdvaMY5ssrjNKj4ggAVO
r3iA4IpEYHs3Yy0btVdrw0N33M57ICnaqhcmTFJnhyPIHhKHVA25z3em+HD9zq+n
VzKc0BKWlGuTyo7OTDEldtvfJxOqjh6Rpm5zNBafWhki0PzcrO1UUPG2OrExG02f
fH5ztPI0VkrUkOsQhkwrdJKmsyPKEPLBcM73doKsUSEoWh8eeXEHTlBiwNveXIAp
IcRbmYkr1Z1AZnRMIyEY8RBusZNbmaMl7oheSN14m2jEOmBIVtv3BA2bpXvueYHu
YBDTTjkzjB0TwKKLsm+rJ0C/WNxcYC4JhxXwMQnafdS8pu8El0Xz0FLyTrOPUgDC
5vBJqwAuthC/EV03gIyAfQ3hPImXXxc3W/me0FEfgPsTfi2GbNQEmVRvhFrd3SJQ
sRRv7o1uHemcyN6rAtGOHNUlE5QSTePxTxAymBXGC2PAPmFT6GcmYVkzB3HAZ4vt
Vui2tqWTT7EuFK2aiTyHLlRzWwW3+Cx2ti7fau+D/56e0ZjNdLJ02pWr/pDAlxe8
eUprrGM8T4dtCQ2xbxkfMZ+hUMUOwYhXOtON0PBWU0H+k9Q5RXqsoIZpWQC15hJj
6VC9rNpHhvTnLKijkTMaKON/m+i+bdeahR4AZ8P5ADtQkp0uJEd/LI+4eG40KwaM
FPPa08FVPVFCSPqYFAsNTQWASrw4v6NHmVPGatFHPV4MD877SxlcunkElLbID/vu
HLPvskGg6uCYHEeOxdExFDc1jMsbMmn54OTgV2Givew+FtFztH1GeE9prxZTcdGJ
AJ4/LN454mbsEfDiEAmG7afH6lfHcYlA/Ogr+FDuVVZgO9EsfC/PPLbwOKtIAXz9
vwYT3y+MNVCBefcT4B7YufhRHrjzNAG39XqjdEqciNzhrgLYrBYQ1JkhnNlEGcs+
exfuqnMlWRXHXASSccqwYPCvizN+ydyIUqSSaKCs1hPZWOWPvnbe6K9j58B669qP
cbrvdrfpnspGmnaGU5XNoCeG3IYdH0IODgeZbTh9dxMsagrVZsX9WrJQ5uFhAWEz
/dBNl6tRNH8Qd+N1nbWL6qmpa46TsQ1SsDBDXDQJxazlkgeyd350MBp1mYxh/83G
T7Crg5Oq3eKshwm2zZx+vj1NaaKws1bKJQCGTEjDG5+OETC2F/IjqXRqoW5D461V
i3LBb5eooYlyyoLMORctGDMry1b5BRTaEk51FyKZjBrMd5acVf4nm9heW7XpAq+m
b5YG0qRUtUCW8T8jHCFheccUSrXSwDhzlt2PCIH8e+IzvGk6B8Fg38YS10hR66iT
SkSHNDT05k43C5p5/diQLLf7LPtu678yC782KGwC/zGDexRWX2WfVDlMZ2+o2BkK
X/Q61MUIvq22NcwIROp/ms+Of+JHFZlKxEO9jVMAhiTWFja4kw+rlHds3RVWuSoj
v/zPvfy66+EYSweRdlvZ/2OkpS+daL5dgLkgo/jqedcH2OJ5pYdFpMghSC3er2qs
Eusqn5u2FLbSr6DxhAwOxFhjbpebcpw7AlRPTH3KH9b5R8ZwdIa1El519ZMEyrr2
BiNyyusKpDsf3kRDlriYfZA2gPgkwNTURwGaoVJNVD8/Ba0qWVf/Pz24HBRdb2e3
cSvc3bUr/hlVZGi/qKCZ5ipMXFJPDGTCSzasfqsFugLHu+6N6ZvGkq3qfGEe5Uvw
1Tfz7X889U5ipQ1M1pH1a1mvRmn6U2u1s3ggAketGbPQhQ1pN2Gq81yrHJLjnP58
huUqvpKKXJK435C6rYJ50KtjGkdh99HFk4yokW2Nvs457akzEnlxLCVZhxKQgYiz
rui7D8W+Z2B6zkHgkD80ypT5fIIETLGkNz0jfF3lZG9XPdwHKUY+iomQBvrcIU2y
5kJNwFpl9Wcna8V9bhFfG7mqjq8Jvis/w3ZnGTLLi2JdIrwLfVQtl8fGlJUrPFgB
Z+Zm0TdK5f5oKwpB60VuXmoTE80yu9nGuNFps7YmiY6J0WCXu+WYfm8Rpiqdj5hW
Z3Ne14UJbhCsI9pLKP+N6qRmallvuGsU7MuTTo7EG+CMYA5/Y40WPaOe7m2rLB+H
cADtmbV5XP767qcEdifJYRIbI0XHanj6UvZzJd3jV7elEihCqZaKe6tvkyzwaTRn
pD+qkRZAkmVGQNodASwni8tnRFtYM1LYyi8c0HI6n82IS7zw87XfSYo9nN+LN0VB
1OQ1XXBIVHpQd9ap0zasR3zBS97F8s0NECZ4vn/dZx1nCdXSdlpzo/l4lWw+d0QO
6StwQBU9Kg5eJKF2cVpFNljTFfefkixP08m7/wRxMxou+jR19rJ5zMQ2HJ49Xcb1
eDUikSal+3U1mBD6GT7/JfKX0tTQz1xhwnbBGSf2MheHk25JF9vM3Bp/Nn6pHEhl
wQRzMRJbyif53q3pCTlF7sk3fybHAsBjV4Ps3/25sWvwGue0IraXGC5wEbrsXg/2
RXlS0glkZCOYOC4L4hRU5Q0SDBPJ8IHFH4/abJ37afkLCkM4Tpxqf6T1CMONiae+
r+f6Rsqc+tBkgEa58ym35dKtQr54hXSFwTwjRa7eqaoX9aihXigFpRzuMYoU4gpJ
Y9hppxxMBmeTc8JWyGQfsnFz489tNT89SU3Ptb2INANe2JRZ+IMJEbySM8I2p3+N
rv3IYCSAM4K31f8QRDj9QlRZepy6O2v8/Z5BK+53MEF+xMMTAK6iAmPFYNdsMMCc
ufURY3XvGYtt3mieCrccV6q2v9YObG7YXt/r2EOcnHUZcMduP3Y9y2gXy2Um6GX8
KvNdpwqYsvrGvPqMyKwLdkoDGOoj6NLfXcTM2DQoes1XSYa2S5fzQNfWdrjwBTD1
FroUicThC3Cm2F13hoaj5rh+atP8fYEKXgIGJ5lzywNITT4eucryLyHMHv+ABNdV
Yq+nu+BhuqYmlNviSOBEMYIQP4fwNQ+Ek5MDdkMPlQ+W1zmdZGaguGu9x8IJN7ce
QZDK5ADLGfGRxl79Wltd2JMH6FNusioQWEv5YJ5iNlz6j9mcLqg1QUjaueLRTkaX
JP9UJlNPiEcR9TmL9kffAMNmbVPg8WIk22MC5aZPcPFskBvAobdL2QHgMk24kGhM
Vh5s8kdqD5dgoaKCPY/wWZsIEbVC/KY607PqpiefUwUdvMBQtaUngPK0DUWfDgMq
J7JGUYAPQxt1aXKcarGBJ4dPprgEd973B9noevicjXvt8pZ6jqgcRLbEsS66Dszg
Y38skYOiZBuV+8CFaL/JlyeLeHZCNpGbH8YseoWZVH13LKk1OfOEDE5biqBfYyjT
ed8wksvhjT6vBpPMUqpLfDwYdX6t4CIB7+91kz2WGHqohyVzUZ0JC+tO2p0gP3Ei
5580hJ8swA2kdNzVbjAg3IfGhBYCoeT2rfYB6jT8EPGzbgtv+8M5xydTbs7H0bp3
hWp8DnqawbDNppNuF8eVevLsiXgE/TP1PcONqKT6jcHvJLz6y9l98DVIL8KVb6s6
GOx6J3dTsjQRhRDR6DYsOyEL0H4cKorlgHCZOIpIvO4eo3nq1sWXOKwfI7PHgrVI
oljOF2Ar/z5uQTED3qsZVhnTjU5x7g7vaHyy2yeyg9Vya3CuG94VExviWKZy4Usw
/ef68WGmhzBGDsdc1izco/shSDJA/hN/pMdS1LL1QoHO04nIPZXxozA5BzHjQPKk
pfn9UPHhpZpkrelRqw22HBDxJZlujSt8ZUzevYj9qGEYbn589TVvkE0eJ1QFzxdl
/AD9OkmhKeomQCJQubtGvDyUYHhiFiuABLuYsHNDT9EZwbPzjSoFLzooGf2Z7mku
z1v7j5yKG2HrXNOynCH5eEr00IaH7oCn/J/RMtsjb+gPiS5TXwQMaVNh/jQOsawA
D9YmEFq0pwauXxmT7Fozi4fWhGiiXc8wt3IhcbrsfxEgkxqLv8ziNtzEegHrpYle
IsvUUHS0K6C7kdchETJidLIICDVAcuaNvLaBpe+4WWI2GgVymo7jiMfdRhZclx9Z
RU+4Xwc72qwGaF3NAHIKndhPn6zYV03J52ox//HT2OmLImztgDY3MtUHjI/GyPvt
J+PR6FwBA62ANy0udr6JnQIZB53CwUf+swe4rM7QF/tXPSoSDP3Rl1pA1sEfbWI7
QPrBDUUz8qZPqRVRKBKTi5HbBRsk/Jy6emI256SvdJLk+Muyscw8hd6NLGs6oOb9
gnR4Q1TB8/RMl/+5rLSVRbgcNjuQCv1bPYEprCbRhAPKG7SHAAytMv7pwZ45ijzb
Z9ZNYqmLpw+SuzQiOp43hhqxDgv3BiGFD1N49E9/aQ2sPn3BaG8VKPs1wd9TMafO
HiMOjxaVjnVGXyUxN0ty5X2A7T3H8asMC4A4L6KgQzqvfcG76XWFtoj7MhK1hpS3
K1IYY22OBIRVCqtfXaj7yOzU76tOzNQIJAmdWzV+7YUuudCE2jephxCcudZqpNZZ
HytTymqRfh8sqDp5KPl9Q+X7zWbNlrLjL1jTS9NR3JjG7jKgF0krPC10Smo/kOl4
rxet8Ozbr0AH/fZZtSKE5sMBCoQ4P3osUCIWITkeKXB/S6pQky0I8BwLtrbZH6w5
DYqOG0YicydQYrdAcub0VtC6XE25oQIuBBHQdXZ75YVEYk+7kRAiDWihrL3WbmVN
C9pOmf/ipNMGb8RH2QKi9zpIVnLdeq/er8DwwQHMJuyBHLHqB2JzP0uL7r4MtLBs
j0obvMGAHuFKIn3ee1cRcS2vlw9dGe0BgLVXSx4+fppgPaO8X+LNAA2+yalftaQB
Azb/NkL9bRm7CLKWtY0Q+qrqLBb/7lJaL4ru22POlHZeiFizRtTfQbJq+6n5wHj2
gwVVxav4R/auFldckr9GF//hee/c4NWklmUMBg5+bzXwkyV2zq0SQhpFcxS+k/4s
rfQLUcxRStX+iNcmQG65+vn5Z5y31t5X437+fx8gooz+8g90RirzCoPmRz93Uivk
zSDqnleC1hocKoRvjeyneQNkswOfjxOjrtLfusVmuYg3Ud7NoKFx2qrXN95rWWJd
a9NrMZvlJeqLuZddGOvMoS1nh5yo/HR6p644XWntd+R1fb/qI/YebN0wJ3qndGGo
TQxpkY+YwgwO7O7vn/+RjMDQngD00w8EL1tSfT4i29Wy2kUdTqVu9Qo9+OuLELqn
9kmUl9vI1hLAHOIKxt9t1I9+6B5+J/8zoHPvc0mHvhA+FK86630+oocGADWZ+utT
45XNECKb1fS0DqhacY9V4kTLqiBmgoqLrcZdcLIK//ZxSXjOZH27mnLTF11Nnn2L
za9k732Jm7FfzXPhkQmC2AtSmfdKdD+ON2kQqtvobMMZ9DX1zbCdHO10w+DM4s1f
5kLxD7MU2MFYsSoBQIU5U/EGxLhz2kzJcvW6BevG3BCunYHRUmYq8agOQQYOM39I
SFiJbrNG8qpJqGtOpZhd2vXEItXjKrfQ4lJgUPQex9inagVwq8WrFEUDX98ukSlu
IGiU0xP7Bx7r5U6P3JBUs8Q6Bo/qLcADJbr024Z2BOh2Luiryn95FwsCMMCOkPKM
ZO5l9mXmCVmrbjorMwHj29T62q2v4ZGwzSaVuDMxThTQVjEtBUG3hPJzahiV7BCW
TtnbMgoXQtlHKc5A6nSdmMWTe3AoybuB0yzlRyvLayMOkkOhxdqquv+ejdCiRcPg
iHbLFnxmHqdwdISJDjtFP6fqgJgdc57xL13tdhjZAXgMr4n80R5lqoiEAVpS2ppG
F+lywELn5GteaDimIQbqKgDXvkHrB/eY586uGR0hMtvVECM2VunTFfre1h9xrwtz
PCZWwK0GRsIiqwmCqtnFfwb4N1hCNIqiuTZxHV43jUr0hjQPsse0EvAe4dPHKOsq
Eeh5Yu7WHSjTBMrviy0I02TgzXGOJ2SMiXhDwr/xrcAnlJQ12V4BXPQPuTKKGUiJ
k4c+TX30CSb/mOAqr537yfrtuCNISCiMCT5ckUH4W7+6aRKN0tMYbvi2C4eEbX2y
IBCTIMRCNHrTBLHEnEm9QaLUigVkkXHpzvJi96X/qbfHezQBmQ6uwnZCqePekVBN
Bx1L7wgN5hqf4NcIB/8rTyqGhN82pXa79XHcFXdNMdIJGWuLgu/HtbfV1Bb74cuE
zN6n8zkxpb8vm307WgtEw/B3YhspC1tZkV7MHCCWv3JvjPos4FO1d3fO1FiTvkL0
vUkdg5oHvMQIglu178HD+6n9D7Yj1liWlc0lv63PM0QcC/Pa3wgL0oSTu2XUTS+a
I81joEfa3E2C8reeBv0IyftAd0M3Rj0DSdCDfP1jGSN4wSLq2KqgojLYWdY6uFFx
qaCC/tdGAzl0eXa6pEzFcdEXwS18o2sX1j3u9pqSQCucJMyhZ51B2DBTGqVRJo9k
kD13C/6guYDjZS2/OJqKfANMY/X6ide8YlJq6XTnLAZ6ZfS8koSEXZvjA8l4mkvS
D4J+uU96IFWSl9oIpji6QrgjhY1GVUdQVu1Obz+jQaiimj3gf8TBY3uAj0dL5OIh
h994Gk+mr+BiqdhB7HEu7JGJFzdoQFjIcpvuwwy5RVS23cvkb67ckM8ObOpfewPM
jkiond07NNMwmMmDG6SQDujvYXjtNusvNG0A1AC69fVkm56RnsZ58QCuhzz9UBCM
Ct4bPSq1iU3PtVOv0iDzjOYLZ6k3/V/wW1TI9BidSvDjh10xKOj3ovRadPBbzoye
+b338V53TYAjrROWMAUGo7iCPe2DZs8EqR9p3YLX5bxVu8p3QV10utrx1+eyO10O
WJk0eq5hgRklGR27/s2bL/3blfn/br03hNUKM4OqTJllTpxjfh9dePouKHSqx+rC
xlOyoA73opzxWewn0FYt2zXLIQ+T8o1Kr8FPl/cSwKs4+AOzykg45nCQEsiOo0xe
/+5u+n9nczm6c4GPC3Lc9m2N4Vcpv0SxL4d9zf6YuOepbwYcTvLmp4zVj+JZU2qH
e4chf06a4qwFjrloOqXZ3gmo9sN3pbycc3NA8LOzYuonyH6ox9lHvPn0NrtCtBU0
Tp5qboEIN6CVbk2zXxl4Brq64YAkbajCWD66CgADzXgSD5HzWf5LwHtTowRccXMw
2454bd17qDGcV3DdZZBj1hyRPsRcnMVbNwmfbNuMXno85/KE9P1LJSWKP9VGgY3d
HBZPMtaGymArsDqKs6acsUmPZAVpoqNWpk50mof3l0l6BnFIa8EUiHc4zuIGSZ24
SZeOPL/654vzHR7S9qn+sX43zyXXPpj5TLS1iQYY9VNzDtXlQtweQJFAdwm368u/
v7v21gXV95tNAknyr+NuE1b+GYO4PAewA6o2exsTMYUEXd+mE9yFQ2kNVEK/1+l2
sWNi5Tf1ZiuwWVQFTsze3TwJgOVSzL7E09bdSPuSGt8wYjXVGdHWLRcJ/hPRhWMP
Bs2voFyVvSXfIVwILR0CNAUzAZtiZ7xOUQwTq4qVAO+YVhlWcgQZeCvpSToslgEZ
yOn4J9toXQkPVtf2AF1DmU+0mn1yHzRq6y39nF1mIo6vPrboNhM/vSbrmREri7YY
xEuyHuY7630PVimPezB7iyhclAOWl8LDOHCWxWWZAHxlQ2KbhwhRplpBO+OHQ/bi
+X5KyTvVi2RbRxR/eVUwi/G2zhiCrSCJsYi0zdkQe+bTVSqloQ2Xv2YrbBYYkO0s
ary2Le/+KB13KbUjmNJEJ7RwxESxrnS4bjfolQz1dCanNPNkijo6NNV4JJO2Oe5t
+l7uAgGT1UgXsD0q5aQn13ZtECUI19Ko6B8IuRDLh1Ue7jSiRTLrn1qczDXZG/NV
y4vuEVkojJa3Ia+ChZbpzrAC/tUe7FS7nu2KBwswtXNWPTTdTHA0fBBGOu49nvax
xy1pE8Drp7p/TXS/QrWzm5HvJWkYQXaryErOjoWsQ0Vp2lwprQ9frjOJyGkzAwK0
EIIYU+UksIYXHuH+f7fobYEtObHNvImczCiaceJvtHo+RlQxdIzQuWNAgby6urCX
UnrSpPpNVna4UPxShxlcmDBvQsCLT5/jyvX9s4OqjN7C8SlCdyygiUylJMScpFfb
EIzeGmfE93mtBIsMMFKNL061CvJvdTYkMOscPFmW/DC9p1Rnb17JXqSL/p0KvcWi
RhvDFp0Syd8uUJDSAILuNkLy0iw4KgVWhpn3oHuwewQxtE31cIxuYaCX6LTcs2kf
iQAvJHGvxh41OXqLwVXlVnp1n+4CFlmnj1sTBQZoXh6wjnxiT9xtlvxOhroEGPib
nr/2k8FnhDmu+WRKhdrACOuiD9VgxPcv5ltbcHOmxNerPr5lTXzoCwAc8n7v6kgE
CWxqR7jRXtDnXUf7482ZiU/zxgA3oDvT3UDxWlJ4zu7njj7uzQA5pWWVkovadAVg
f5/+zPvO5SjjACcflnCi8q5DwGqty+SI3JZfOWFr9SukLEpJB0uQ9kpStMHLgV39
myWYYVzWpXlsKEOdjovbeHzkdeamOkNvutVaMyaihWYuw12njOQ2olVFD0dfWfIw
hiSfB38eonz70IUw6/57IlKtG4NleUsdykY/aXdXZEklInLGsrXIJi9I7/RTBJ4i
K3w59yPu+LQ3YnQjgFKr3IKZ7jm08WwwzI71rFg5e/UbwCJC+BGa0FJXIt9NU6W2
5loS7+T5sNxrs75/SRpi5c1e2FtAvtmrCH9vIdIkGlhXBUXDg0gwIybc4p3UjSwC
uihoYxqYXxNT7cIWnToG0Ce4L7QKbPOjEhg3+eEgyKPI4wMzz2bneYIJBFvNWf0e
twD8tJQDf6hcDhplszRWON0Ic/DGOp2dMRE4QsfTR/Vf0IQgfFyBEjtAqicZRhRH
isMPyZOWnZK/Eq94M9waTSnzN9b02U2Yxfoe9QgSavIUhIFndSkgrI+uf8QwmC7Y
u3+TMKalVftj7KdmtKvO5PRe9cIs701uRCnwkecHHYjWp9chcb6LF0cMMzOfOpvG
xGtRwgxG18NKAFWiEYK/gK0uGPgRyHt/RspiTsQwW+t5sbq6ra6PRpTnbn67GSNY
+OX1FWU8MK/0DxzL2e1mc1JYYcAq53v4cjcS0aYmm6cpxAMj1SVhM9CZi4ApU1yX
3pyi2gaAKVBls4ZpnC5RTezqBD/NAxmZAFsnJQuceGsyMTy9mswlgT1hEc6c11Ru
7qv6spoQ6/4CkLplQ3Qq1/xOAYW3Lah/TqJLPENkPOlskPGmQku551SHivEkKoyf
bP3S/7sh7lAXbe2v2csr0E1L+a2hyJIf21C32KVsS582BSRZH6su+qrkFtDLdirj
QRMBYWjh5gGWMfOpNZhLZ9HjWgt/E3mUb2yFA5HSsmhHdpTRCEkYwKgojxOp06GS
1dGAeBnlhaq1jzRZ0RhaIU8pd6G/XaTbTTIvOxya8c/3d6axs5eCssiEW98jl8zh
5UhgQ7zjqMkOaV74mJYubp5f/UdWmOVlFof/L6hMckZF/A9whezRWRmhADDxIYmU
+lwCttmeZdqJGpcMTtXtekDDJmnUCVqsNyP/xZgzTyGSPJN8RuGt8axkJ2/BtX4o
yP7sNpxPlbfe3uuHJJgO8z54bVeKLbcTcgLWMhDEZG07TRj9cx//inwXcVt1EqEt
m7Q2eiH7V7e0YkxESZHWoecahtmnXBf4oFRx3SRNbEjmjYsn9thQcCsb4F53XQUD
cl0BIx/OG+eQZMmuSq4RbZQvVnYQGbbJ+BoQtGcuV0k0Lrr6Bi6tji9kgioxNdvT
Fs6sBwVC0t/h2IAZ42cAVrJiyJoo3mm4mcAMz6FJhEfNr6cRYZNf7uFRJZFIDI4C
TGpZeeXnDtNmMsUWhiT/wh+zzWofGntr9TNOjaxZLraGMJ15gVgGQ6Q5Q57y3MOh
FtpgAK4VH+d05Hi6DaNkeAuervwat45YU+4PtOPJWQlZqeMwgZYg7cQWxiUnjnrq
vXrlOEgA8WVd0ZMCqdThCN1hTm7en3qh0OTFvMsU9QEeq9FDqxu4brQ1GFWKfrm8
jI6fshWp9/vZ21p74VWDkosc8HWON0X3QguGqwb6KJ1FSXsllJvLQexY/HIkV+wk
5OPltuvQml67vVfwCIpSmMIfULcGq7slx6xNCNkQRyjG1y7qDQbZYYWrr4a1lFgm
2lYNnLAzBDguWMl/qwZuRpdC3NapY2l8raYsaFTY4wwx0HWWXFXEnHlWIvefnOS8
lrCKNwXHpYYPpReoKtAmMy4GJ6yQaHDRlNYEGUGUFupXgSyzyCamjpdENh83euc6
rrPhL+Vtmg7UeMqAsK/Dc2+TB46n4ifi02p5AsCyRNxnJYcDJG1qvYWlXODlddMp
/a+AaecLD8F2GCKqnXIsx6bsjVldkuSQ+U0UaavsrZvAbOddnRF/flnUN8wJSAwQ
6Hsxu9+G7Fsd9nlJSJBJaRJ0S2SF7iGFhJou9sfRdHTDidZ6jh5RRUcWXO3DmHH2
bROrzxIBO7f0rKnj31GuL1aOa5NUg+Apb3fEI3HcaGVz+oZ9vD500QmRc/EMCQpe
aszAA8EktTMOzmWLrn3okkJ9BhncZnDulhbzG7mPUWkKwIMjrLxCeqop2sj+yiJq
5k17CUH6Ll+lyRbEv0TI8odDKoj8DLHQ6eZ1cpzf0ZBlFkHolWwTJJTSB2c6u420
j45jzEhnKB1BThWoK9OCu5KkfVIm27QFuU1s1OklyNPF+De713X4IIhNV8xvL5bI
q9eR28Z/1JM59Oc4ZmTlDp0kzAayScZVOllNA1b5M0mXjA6b91dKvnVgtuLnj5/S
YGqXeWOOdau+PNOWRiJktFd7U5k8ybXeVISQpi8hvhrKsOPGzdMne8saxYjJJ+Eo
9ejnNLVpgRCvDR6cpZKXG/fsx5HFqhtGytiw85WvMneL3qx4K/xKfqkpzsXcz60b
TsOawn/nT49vl/GsqB7kIMntxn2QSq5m34sVNaYSR4elS1spV0ioHtSIkHUMDNra
8nSG6eBD7U6jbmxdoS/sg3i1MPLEkAB37i8vX1GrYsXDLd5jQFL9OHGGzRa8y/d+
sxXA1k2Bv7F4VHqhjV9s4X1tp3dbokRNOWLWBGI0LoNOrKvpB8nyo3BspNdm1OUX
E6RLzCfB+4Hhf3vAR6m1EYmTQ6fmJBdVsVmcf8sQ1Ik5etSQAWSV2AAw6yV0/5TI
y2U9ZYbUWaWqU+kQgIy0/E3t8HLwzvlTJ3UWiP0d1Oq+45YYstqQx15KmGotKfy3
De23rGLNwrn1m2Pa9m0OejD4Nv+YdI8R9iVfvfgjCOtXEL8WoAU91juYaU+4+X2f
d6YHdVsNWvTILwEBCV1swyFqhmtQgB0hwGoyRTAgqZd8rrpmkFo7OmNKU5JZAdhJ
cw1/EbENjl6ttiMBjeJbXxbxMsQVZ1sAFaUXgNZQqbAEztTP5iKHDuWBbqsQx0zJ
9LVJ0nWnFor5tAvk984trJMX8I7GwwDF5DIczFnXr9q6JdpPy75vuGU4owCSVdFr
jErgAozdP00zfaVhRrsqvENlIwkJEajEqqv/R4rQnNcCIg7VcJONhYhVBQz9gcu5
HJ5I24Tc7ND7RQtJBskbhlSXYAiCgWBJI17Eaka30y2NUcEdw8KXXsXR9c6c7O0I
aQepsABxwTPmlCgozExchFybiB5JP/xfhGqe7ZeGYhgtXqny00oqPpAzUHIKQpPo
7x58hIrcZBNZnxyqVGIfMTPfS5BbmeuhHDyl6zPE3jVe5qXbm4xpCTJ3MLOzkJrN
Mokh/14876bybwHtXTVC7QZ7nhEz4HB58zDc7XmkqJuHe3hCeBS3eTUX0yW9dc1k
0mxIq5rIkQEBzW0C2KAkgXB6fKtlgO83daJr1NMfVf1Erbzhsmpkt8R8Y7XLGgWw
HjynXzj5Z52H5L4m1NBiLl7/b+1PcMTWC7P8ZETa4fOH4AVf17bnjkX/WNV+Ii7D
I5YWil/076D4dRS3N37Z8gaO+0u+dZKUtxz3/t0+MKXYyRLTGhjIeqS0zC6OLncg
lhsF0GStQ21c4T8d5XtZJPZhjf28XbI5qvsf7eWl8kEDWvVvpR3EgVoeH91L9J4k
NqPFWacsaGmoAlk7YDLvn7jN2WmUJG2yBs+t3WqcdVQxxD9dIb5vqf9rv8d9yY3l
YEbQiGl3l/b5kZR0o7NgT1DMqFvsJlDtZBZ+ZkjNEZpJl4zcEODrgctiuszm/zzU
oNooj/TTaDHkFI2j+JYjP+1n1TOeCDfpdHr5vsgS02Zn/8iBlLXpt/Lq1nigx2AU
PWBS/PDyb6eAiNycl90TJzCjktJ2QE6FzAlDjJg8y01qBUgUMHPC26ogJKrcK9Th
uFHiy9+NoLAeb2nuGr3naHCb7FYKWH+0+3QYeXF9wy0iwMFNn+Rjlq/HdXIBeT6I
v97UemrwSFHm5Fzo9/xxm054dc5egLDXFKnl5gY0oXir9i/AMqHulcZmArWYFPkz
XtJsP3FwZAzxzJ6zYUR1p9iSIqNstK2s377t5Oe+QUNqzReCHfE7gQBAaFf5R007
mE9M2AF07ehM4CcdN65gnK8uI8BbUdBKoAv7je8Hn/Sxf7rilWQb6QHidFE+xBRB
lrZGqBXiWz1wmxg650Bcx6+oCI51vEnM3g/65cZfKFNYCJGjYGY7TzRCGh5U2p04
iEn3P7qBfNjQXsmKRkWaq4ZMjonGHoqieikbCS0c05s1uncOyJ/No0AmAwZ6j3o+
xLSv8Z4Ti22zzJAYjK7RoRNF3Ozj4edU84IEhke13yBmB6YMu9W02oxfzwAkuQ/K
pfxC9J3HtTb1nOrBX1N6uL2HBeC7LnX4vKLp7peB8Lk0Vxvr/ebw/RDOywP59p3u
4DSz/tO9GBE4SxJStH906rDIvK3JIUojPuZkJk5eQkImqK/JSV+LEEb+i9gn8eXK
5zG5AuIk4PVLzZ6y1Q/hN7gjcCZBpMBHjCCBDhOpy3Sh79nTcu0cqY6yLbSFYqie
BJwynyLn9og/cSgvyeMD+PTtr3NgdFYhh/28X2jntTiaV9ouceTNPezElT9J8TUg
ESaJgcmujfkS/l4TI7lRaQB0PO/yb7lr7Bt+nEVMUvKb1CMn5H7sBwS36fe0rZyA
SeS4SnySCH2OqFgaJsFOJYElyzSw8pzmOtAEjGpb+58w/xwXjuZ0Vab2r/0ATYCQ
nM1MV70AQRyQYZhR3ydl/FbSmOG7/Kir+kpJuTb7FSpf1bcnwY4YLs37bDKgYAfb
MzQddinEhOxQghGX3hGryIuCLYoNJQ7mFymQqiqXl4cJ8P37tKdG3185/KESt30H
UAanD7goCVonmtlCDlijUURIUtXiQyH8mz2hLtskAsQaq/AEaQsD+PUTnHNNMoVh
AGUz4qeMwj37uS2zPHMx5SjFmn8HG03WC6aIN17Iq/YnQB5SZi8hNtdTuXeqk4MS
dzZr2JKkZvrzzx7nRNeLH97XzxFNDKHOp6sb+mVlYMdwK90TkCHbLQrubkOhOakK
ZlTsLhR2mHuCfAEeQXfVJSBa0aFN0fdmZjcdZV2Jvbj3RhDJ9p9gVnMC3aj0svev
+rJXEk8BofvIUICjZV6NzMiZ3/yeCuHOTGdDM2Lq0GTPlIjfSlmxnyDP5nomFKjP
2Q6/RFFTmzq3ASijmTcgzoKZR3H9kQpaTjq1J7F77pIAd1Z1x/V/sQafaoWtiWzL
B1qild/VuXk25qauTGcwcMX+BKW+hHcEFyeDQCOV5paK0uLrIwGTvlRXJOrFssjo
GKWdoDBXGxjvFEogkqmTxlX+JV6gGOC6cNnAUTpBX8xAiT2sROplRi7AtKrwN6Cf
X+1r/xLny6uEIr3vcuxL05kZz4P0m9VSqzm4uU7eyxw1m24VlVFBQxKsZ+nUywwS
+BQww5u3pY661hdg5vejpu0OFTKWskZkn/uN++cYB8bLqIlujpHIy77fiWbgVQJE
hOZ3HFpGciN5TiJNaZXGfv0Mb6LWgIp7NyyR2RTvjY0fp5kQig4loXYT+WfFI33q
4TLYlbJ/yDZNiFmnINBt5VoMklHvNPY8adq/itM0GP9y4iK3y0HmXs03jNnV6RYl
LsoheRRwGtZULoVDG0OSo2QjMbB5+4dW/KbFhCHYavp7N03uxPDPkmA0g03CC4Kj
4gjD4tjNIaFXMDDjNA65t/iPYn16pbujqKPUVyOu0hKVQSNhuzFFTCBiQjv6+guq
Ivopy4SFtR9wZmD/EdmQaaxnpO/69d7Uxgo+DpnOnrU3NF65EEYhHK9Pyq5yiOvp
wmNYdpCzFouaDyd7AGsKHWPTQJ6OtKEAe7SQWfmKFRFl/SqV17bFiODntXv0R+sp
/vrglolbeO8+ZjoIXyvjxSiosX0BqjhWTwq0k2OXJq5ZGwWInFEvdxDaw3xpSQwy
SfxSQSPia3FMbPvDYBFRD5VuiXQiyKNw5GUl56SrIrCXWFLzYOHjxyuOMwRcVJtv
C+5/oCck+JzFSO4/oqipDxu6DaUVBmhyhUZn/+ZlzXW8gk8aPZ2QRqFkdCp/brKq
urp1OVaqR6fKuo+WEgP8OkZXyOTBoEiznKJ43W3o9izvjHGTlz591kepgZ1Ds69O
pe+SwTlk/2b1Sloh5BJJUe9wnLB60EoPQnF/1XUR5u2VpGxYdQka076kaDGXY+vb
qkcvU9kgCNWUZKnlzT2/SrCBttY/jep4lzFaDKCLott0aB6Vs/lo82ozujRdFdJ+
e6NCN7RDIzZEDwsnEjdviOETTizZ0+bkCBpUdXoZY0VBsrqUsNIpn1rERzCY1nkG
/8cnoW8PIucCIdQsBFoMunSIc3bfx4Y4BkS2RiDvPFGdSgRfKV0zLMixd6l6dQYV
j1oZ3yJ6B5ophLS7R1rHc/eL+7DNJQg9yeLugquaDMGErvtje23GRDdop979RAaq
qo2ubtSckmTsx8Vz4oepomiCCrV60gNd8IGoorBMzfF779M8enWy6UsWO7+yLyL1
Z+qomkp0tI17As0KZhqQraeEqW2LM/5HubPxePasLIe/jtlhno/fHj7pXYkQv2g/
u9cfJd4cJZC7DuGCHyQTg+KlEejYdiYgfpKBavHE4buyBVZ2UPEsloX/LG9x4GrO
y+XVrXnVlpfp7z0C7nK2LGsYNAmTvTLUIlVV4r+Gx6JXqbpse2VwMehW372B6BvU
HaU2epDFHJKYTWDhCofDLyTZ1/RxE2wuCCw8g9YU0gQWOYejUR2Ah7MB2OJDNX+O
+2RoeOq4MZo3vZCUe94lTbpi+kbo/Xqa8v62/vDG56Nsrw/KaUG31iDPSkIFX0z3
DxbBbjyKIYzNykxaLf4AdOqCLGAEw/z17+LgaQ5VOLQ40g4wWu0Qx6H3+HxiQ2DB
GNPp7KzJO0WD/i/O/984oJTB6Rb2T7wWycfJT5Du2/OzsPAHEUYEwEuSALEETCUh
dNVfAC910d63vdtuvtIArFCzpE8H0hCDGuyXyNy1788vD5wMY7nyHS8YtsGYOnuV
FxN1XHC1JiOtefnOgza1/qy0dgA1eeJI2SqmHveleOojzPEFK8db7mq/6gPUPGmw
2ZstSjA0eNDpw+zEWPyigonGRHe5SBYDTr9bhKLzOQR0a287hI1TDRXt7Fj+Uey0
Ea/WROKxvuRy5hmRvKjIOdvaDFhAvLzE0VK0IHg4ey08MHa8Ydby6vBvyvXHMJBx
po5ExZuZ2zL4pFRDv4qXm8/DZnJC9JxHhRiVRxzzOoLlkj9fX8Fb/J27q7lBhan7
maFQlyf/hlf1uCrykCi/XP1e373vmh2H+Q5qZY2uhE9fwzg0+smnVlsnC5NqTkgv
+sUZZK+3EbZo6ihD6avrnJxoVSlYXb7d+XTFuTBPlUw7FHo0eN5e+4kf0Bz2gG9u
VnxE7kpTmXcYkyF6pACcGxmPnhsEtlLOg+fdlXPwPyOoicy3VaLVRm3GkNrbrd+m
cnFm+Bai/pADnqySV88RYdoAoy1OzKA46+VqbnrgGGHn6/GygoOvY5whbBfhEb8u
ffkxbvw/V+ak0lLuo8earxO4EHmDj7k477xnr9VbhXDb0hr9DOjHD0fYNntpalOC
MwIi+lPzGGQsg/dLscnuZA87stf2JiRZPvXctf34pANZK2B3L32tTAfiM4yNfPJK
xs0s2D+f+GZo0bkJado1EkVMCbwgOkQpFp14yBhPbX0umo5ddSl+Lj3w14C6HLft
Yay5v+ITGwVc+i5As5cl+VmTegqUXRK5utI51V50PE8SmpLWvok0+Fv9x0zSsI+m
hzAdPcIsrj5+9Lu91xafT+EbxlzxvplI9gOtHOh8jHuAKN0tQzvwHeHSrIqQ0EtP
cBPFHhkdExR02J/McjOQomzN1Xx6yYBtPhKu2/nunyOuiBa2epYw/MX5eJ84Y7QC
v2f675bfPQW74JmhV5fi90sZQz2cHOLiBqQ29SnvZy1woLt38UX2vabn25pBwgYX
MrE7dca8FDLuk2CGqPgiNEzyPYn+rnSv4a1Gp9sQLMUmbg098LdWiM+7ZIj7/ngQ
7n1NwrEdskgY0bcOJYSgO1Yi40N9hgkwePtkQSe/f+mt9tzwoU5BgGFbocVeWZ8T
lb79RilO84DROdgkDn33R4Bd7om79lxQzL2SeH3+IYbKey5JAmQcL51WRacCCWlK
puJaGJZQ5oyElxlnxUi+ukSI2VKHINMPf6/EVAGJcoUfvBZQDPsTDD++w1aNaipV
wnGJ4e5tGOQMa9lCOw/vaRdGRKv96tsuI1+38/EXtrNip2+XafgErF05inxuPyl+
p9IgQhyyNQUk5ha6snKloyMTLzp/aKyrT8nxAIthHxBKm8g0AygDQpKh5M9RsYrS
mcd5TfQKrU2RIHZI0z1b2aWOnXtsNEehHIc+rNmKKLGADTqSc/obq+oLs+XKx9gz
G/iK47c/awYP7jfIghK1Oez0XgtVu4aadlP139QB63E8cO1CEeu9PoSULeKAcgZt
nVjeOidWLFToIDhddLA2tafqNK+26KlUTU7RMfPtsH92qah8uHBeYLCpALCfGVmg
LHJFFW16tKMVKXYsptOWbxCu+8jb2FqLVgluaWDDITJpuv7gaAfoXJ77OIo2hZGa
RzJPKCa4jgBYX1+ycDeUQt/MkWYkWULU6imn4jqw3FYnaN1nsrcVpfxlDyWk9CLG
Ta9J7FZGEKOJoXvncb3anKzcFRqRvI8yeNDDnom2aDQ9uyCMCdW5rW0SP8jCUXt0
U8Bx70yzcIKrPLGaJ8dlO8+vZjMJgcIi+DbOmilzY44xhA1UUHQmzzuPi4aHr8xc
Z7+m0EeJSNuvGx/XIuGKI/Cyi5jpDMzs32yy54JdmPLHvw5LFaa31z+kgFYaFKj5
qTdkC80BpMHh946uv5RnrIJK0WGcpVXbpTxWto/OSL2mM8dz2CGytxG/dzQez9Zm
qvcEVn91ERMIKpdZHBhEBfPsmrpDXueP8TjkZwznQjbhdNlfjfGQ/Vnq3GEWKpBx
2E2hXL7TGq2mWgIaKnJXzsARtLT/FvpUIoArPLAlK9RpXwFTZYqDWQ/U3+gsEP/6
jqF/Lg8mQX7ejv+7XmTjE1A1O6ugoz1PlhlU0Eo5GwINyeGEgiAtV1RbGB5uizFt
rz67DKKEGTxXiR/sVLPIq3c2I/ixw/e5Ll362qvXPH6hXNV4GqI2/5yjwBPYZZZl
L31tMo8FrT1Wc6V6A6oMjxlL+51mDuzIH78JOhcUwSqjq2pirJp5rKkzKdjMir3U
CJsCSJigwosR9Yvhl43zN8cz2c+grKbLk4mCrVGHGvS8xroOg5ztqeSt5PnGuvEH
rbLtwIab3OCaOINc7/XXczUucTcpDttHy/dpNaiorH6dtGseNquWCwwqzrQMavnF
wpDVRgu2tekjvAMmCEk0/CqWD7+Nj4+TezVGpb52+z+iyZ20SQsvIDTImqMQZHkg
8WWwYRGwb2LCFXbabKuLWIZbqiiYjTjUq3eiNVuDi2xJD44D5epXce9KTHOKeade
uZLe1UfgkX+d7ZxdZiI/zwuS2pXv0WqHOkgYgSgLjv6dWjz7/KjsvYoio+4QAfe7
uFA1/0vBbsUL6GoD95rOMtiYU1O5RqawJWAtg8j9CSnJkBbK+iHmHGqVazZo9J+S
D7aQ3Eop7vkCpvrdAsDXofoMVCll+9yJ/2D12s645pj1k4jli+Ealw8JZcdNYNuo
lXqdmY51SbDnM7ZMwEmdtZqGSqe8hC8IWJNhkg9DUcGioZ9OAcrGbArDixnhh15y
IEkEB8b+eCRIEjkPCSiFk9Nwt1OAd/LDv+gG2KTYzzXpVfk37QMMS60cokKgYWZX
Y8KsovuZXvitcXUQsgnx/ywb5sKMXUQwEsyC77j/x+ORHcTCdBEx0I1FF/XnOF0h
D8qL2M5uu8kMpWDwaFzw43fI9jiHJmQVe2HvhKaFEUXe7LI0sIIDSMcqqBvU/j+f
TVvmYo6VZAeEBexgeQZWwMWHKy3wOGVhaiUka91gM41b1IVKOZWBaByUHW1bzA8H
P343rdErijv4oirEIo/jWsJn8KDU/n/jEYUOMoVnG7UpWRbZSeYrd36jTur73Z59
4XTOKM2/p0KKm2VT9R3pbJsKrAhQAzYvwQOO8Jgj68kVDKx8oi3AwC37vz2OjEfM
EOwFzdYMxRHz36hnu+xbKkpf1WLQkFiQxeNbeoKIUhPN0/ni/T76pNKatGndq1ML
XTO/iffCgCUh0YHVxY1LH7rEI/LTCOn/pvU+nvn9It7+5/5ep1kQIX7qsAU2KsRi
Jo1nsCw27/tDjld8G0NKv2jorS/89IOPPBsl9uJ9a5f3L1lh2gSaS+fe4gkQ7Plr
xwnn33vX/uhLXkXPhNPW+1Z6is7EoLsarhqxSb5d8y+9oGPO1de+bF73qKoVAhep
Q8aWofWs7AwSp68yr7YEhZOZnXQjBSYC2t647xH99vR/NHX7kRbZCaTk+9R3S7Ba
2Uc+OpyulYZ7V5phGr+ruqOUwjLE8qhQ8L7c+MUqXpHfiCfjUkslc2Bpi+OD5dR7
/O2bLxCLpZBbHRPiBJHh30I+rEp7K2P0KWzEBxTNB6o5v1I1n+px+p4yH55e9kQ6
0X4tdHCR2D7lkVQovixD0VJnDlAbIRki0GO26k61KsJwTIKLIOZWMg5C0N1jTsNn
baIYgw0FJTZa+WneeiZ6bLzAf2fl2fUxVlH5QvLtDQNbn+TDdRfbaArwg8VE0Mzq
E9zY+lB+L3oV5vkUdP4tvKdBvs0Eaj884A6vbXhMt69//gk9aPLs+vsB+51w14SJ
Jnis4DXxdkJU3A4Ow1gAunjM/5WMcK0jEcK01Wn+dccejkIA4FBIPF/x7jncZ5ox
8+ftVGTxx+5z0kMMJT+ows5GbIXchaaPfjkTDQPqwClRf435i1nCTFi/m7ERTorp
YPhud3rkDSAyWqAGOrMTCEdotKxnAdxRvWOmfy0FqyVr6tytIOKM2y0PSCtSU3ma
gZW8Dxpy8xzD0yQaES9btVWBjXGt50/81kZRNo4DvwFhvhNfSvzfu5VrIfSQ0yO5
03+hqkbbeUQZgaBD275xASwSfpHQuvjROiAYUPG8gaa1t4lFU/n4fkKku5xElwIl
PRgMvRq1HwBA3jLe+oC0pDxTMz2L3yV5p45Pf6aPDI6xAIPoemGsHIH6WiGkHdwZ
nx4xe3S7NwFUmu9vSg4ptLrJzVUv6ZOkHsZ8dB+cfG2wIdPumPdooMRK+9JE0+Rz
QL7DGfRZQnblFx1GE8RtzcTBEIdFmvynp3o3O4DFQOLlwdOcHeKSSfPZJ9N1hnpz
RSpFgjKlEGW0bsNj0mM8wXFQTnhciNuPcYNUUpZMFUTN7YXpDkJKjs2MxvgueJLf
LOchu2ZXW82Nr1bzzfvK9sW5H1qVChQwfqRDAPrvyzJIJOGtu6QnHtFNFcKGyYCk
hH9hT/qK/xkDzwp0z0bnwyVCRkhK3L4XAdZIZluTZLaz2HzUGmpgPq52ZlPyGlN9
iK+2oyxrAvhFiU8OuAK3Y2HwgZcp8iW4WJFA7fM7JY6m2MvhzG4jPu0F1kQc1FuD
ma/lIGLPT/feAl+jY4EOp+G5YZaq0+r1TRj0PxjPonnU5nM1DcgBK0VmiB3k6zHb
MN+RLvE0A171SEE94Ey925zRCw7BhS+jv/Y+6gkarmRL26PU5h+Hwc2GjUq1TzWx
B93rqSkDFoGgccq9IMHpoJD5CgfEgPhXjC+/Wmc/7xytJ9cfUIO93OB5wg88RFpE
cHdoFOYtTpzuRDXFAiJjRZONCfRg2VDQ2sLH2bO0rw08XbEek7kiUYzk1xC/lnBI
fyx7fh185l+aAshaCU2ERRfdHgYoyWEhLVZJ1ZaRkC+/KAklPnrZEK+Vy4YK5h5w
m7Ex4JCYOVKoGFwA8W+f6gNK1XU9Y3Bynl9HHXwHugscj2oVcTugs+HLQl1p35L6
1EwSutOPmwQIU4CX8ZjaIGWIrr8rKNRfszHMysBIquImOKD5KPi0Xk2IvDObgb0K
0MpT5SmBGY1DaB/xoMQQBesC+7Y1u4QtOFhm+oaqJnD7Qeyb7QFLBwU7yKQcc14t
w7l84Poh3mKsF7XqpAAkzXwolOw9fOCyP9iyKd98sSvZ/lGx8goDpjsgu4ptWL21
51elCKBdLTZaiq5ekHMfgmyUAZKi4+jWC33SzB+58hpGRUfs9Gat7Tgc9Om63t2m
yJRNitOETpi7XWqLXnnslrArSgEvVLqPzw8dUT+HBaVdj+QP9LLXcbAT/+gRFtDA
Ho7023eIrkzBcfHA4k1fCEL798pg3DHIOpuoz3LZqGr5k4SlZiLhUbDZqC5kiP5B
hEiPgLswUO2Zx0/k56cibQeNwijlWb4HmWU2vPuxsOF53mBf7zusmkDcDDwByWfn
qjSuAMmaJwqgwRCP7Ur3LyYmpaETUhxD5nnJUKD3eD2or1sz5yPyhNYy0aW8A1Ei
TRF1Zrpz6iDZ3om2LTXGo5etbNDGMEicaevCxob/ehQP5Wp6U0M8dc8yFASOgzKC
RY0yCCCTOnznObK6Ekc20CynVRX9/UUSKhIM2DsZgtBwWmLOVAiFTevLcEqjzB25
KYQBZmWU0TKCRjZB8957oCtbqR5QJ34PAltbsh5Yoe7mOfgay84BKQbum1gAEkjE
LsMqBOS1jAcGCmOEiomKaF5zUz8CguSKcZdM4EaVE8mMcEs7nSnz7Ptb+b68Aj6Y
/agjq90NQe9DitnMkNZJdJ8ZH7zWbqypijo9Bvc64nqxFHnFaPX6uOCUDn7OAu9j
FZD3MHPR1cphCiXIehz8ps32vnD69NtDHp+FvlC9SN6QoDJCR96dcNBwJZT+8aZH
ElfLwHybMnc4k5aJicKJjANFGngxFKjbzlO3e/a2QO4pFJISI+iWkLeV4r6tAmdW
8lYkIRmiAcha8KT3wlbkFneYLPMj/aSc08NZPCL2T3G3PLOgmDK05GBFhykb3qBd
wh58cCD1intRUdIb+ICArzBh7iqY+vIOP7FtY2CbMSGALkvMt73HhzXYD9qT3ssG
Kc05QQdgpDInaIPlQW3I8IYVbRT+5GTOtLc/v9byOPHarnKQFQkBty05YH27QgVs
RXc5o28SN/JgosJsnomvzkvtUd22fAJeW8PIXMypkFA0ei6fu1F5na8jz+/c8Iqi
Snz/rjb/DkUQCQQHFDQIPGhvQfdCqWUK1yw8EB3AG2QzSt3MT/TjIOQZTebiDfO7
6jpR8jTX4fIFLSj6hX1pnD6Jw1jRfdsOJvsHbtGno1M3qqle05MDB4lzsRSIdRka
80wxnKaypAplY51sEZ3VuPLlKdJSRzkJjOzndGIrAUkCmJGWhjcQUcopP/OqNLJu
AMa3maY7Q0vqrshUXVQpdxFzmIXa6HNICg8bCnR0/1AROe7bzLUkC6pfc31C353B
CHWMjdnlBBcP6yJhhVV7APKcDrNj5ySqLt7Eo+eyLCHFfFiCswzom4JVGbC1rlUa
JYABxQz+Vo6BMKh+23QRAe9Nuii/ZUA1eivQ8/h8MghD/GIXZm5vNHr0+xkvEdBr
wBbYEudVPWRwyfLMMWj1PZl3NkHPX3YRhlNGg+lBTma5Cjqt1NMJC3amA/3UuXWz
JFFmb58+0163Jk1yu6JzMKkASLwphI/BhcgyrlBzTb8AtePBA5nBz9Nxi9ejRcwr
/UyU9UEKHW7S0nYbkqqo24OLmAV2xzxXb+Qab69mTE2KQ/KwFPbtm59UsaAyUKIW
fKLoKOUvhNxGmSOEqV6UsRQz/6N5/P/hzE/M6WXPPWHf4E6tPo6vjuTbr/BT5iWw
yHqgFSn0IGxD8rSeRYanWZv3GIwd+KZkLN2//HHcQyXOhedNQjum5euvo2qN7+RV
OCzsy/m3I+vESZkpSL9dL6Q+hO4bWfMicb1RoHi08zYDnTU1Q4Uk8US+nfzR2tcf
tLnGbc6AjcukRXbwM0WjSngUAFQRNL7JjwYMSFiRXapMckUeKiO2l2epeKMiwYtk
JbMl0wiv1uytjgEyAnvLYS5Lva2f3RzLZ9xU8QQDWLVOnITUvMDblw8ZaqASABr8
P645Yh0YT/uKjz5f5HU8LFCbQekjdUR/ArjdGyp2Esqgyj3AvHMeczZhB9sVX8X7
LpJMMivzSgs8sFySwRxA62ej0qBjOQDEHxqUY3RCyBbB94A5Z+KliA5sMzvPj1Tb
Nex90EQ8bCWl2BeKLkAryR65p+dAMBb8xDc1KufSpvzu4W6urUgXfW2ujyWB9dDJ
Bh46+zCpOvC3sqtNzvz84p9IYPwI+Tb/31cbum65t0roM707pwVrlCBulirYAs/1
SPqd1loOw+/yoBq0lnCk/4SeOPqk2FuO2aNx3mZPagnvFWB6xrh+47+HMseRzlyz
dvkx0a3wq/IQbBO2dF5nzQyukSP4W3R1FeWu7EhZ7ktk0mgdN7JaZxLYdJu8OHAi
a9x8+7b1+b5QdQ68Z5U4ZLe6asOSANg1L9EQguZF/KkBmI16pULHhJVJAmAn/JwE
BOJQNWy002Drm3zH/HQ07gdVPZG4HdgkTHK7i7TVlMnvriUyLUyay7spE37gPJMJ
MIZpdzRJzpXUddP2ISKhXdwHXn4Hj2WLUu9cEatge7Vunrqla4BtHi1DBkugO5/2
eY8AFCrFRQqL21rMmfB/qiawcF1M+gwS1jb2YtRyvchDvLkMgtT1qbX5eWMDUUNE
YycZFgJ+XGlERyh8PH33IWHpb0igi4IVJYXwE5tpX9G7HtutuOshPA6maMg/TrC8
uddS/vW2chekbcOkWdoFfCQLq46SHOzTZEkunW4xUBftqy/Ix1y32vaXU4OE2bPX
kTTnYx7tPn3SZY24t7y4TWobIRrQLF6T3VEONZZ69lHPFf5ShmjpLLPjAfu3MDPS
DhsYx0U7ma5hY1H+dB2ujRQhR978/Te5rpYKQjPOi7aDFXaDJgGXbsCNGzEU9lV0
axnGqriuidYHTmwcjZcG0vdUehx9dQX4Hz0V9ouU5MqkEXUBTALOdHM8AzdX5tkn
urfJ2p3aHkm9TQxXhFvLUJ8jCjpB1Ew7JydoMA3hJDFFcXAJumPjRKO9a15sF3ZW
RhfY+TVUetHznVOW/OfjB6DV2rkw9IOv8cEQy4KQBnSQXUo66nALg0Zbfg4uP3tr
0RqmcgIBIka1f6C7HiNk2aVaww0EVtvJ7PH+1dAZknQC9pQh1w8Aixvuw9PRbZjZ
iIf3q/2l2J3iEAmjUPjmtiEkHxcAFIgWRMf0tnuMtOn9DMIgv/idC9BfyuXZdATf
1xMEgFeroRh8ru+VxGb/wu8HfLFaCOjUMFGiSrPevcNCbuFE0lstRw6k71QmCcg2
lL1M782jrtJQVaUiWE5xvTJx5Re/HkOT6ONjGRWKPkUgvrzqZ7WdsZGk9bJM77D9
S0ict3gJriGHhM7+AIaep+V3GrIwdGdbUXzAh1rZ4ejfWwp06jSj0fqvyg6u0QtC
23Nod9bIOOmCX2M7iyYICE0YjF0DUwzvXBtOm9aTPOdwn4/F3xTkbxE6coF9Dt5s
VceyWdxMi/+Qt+w7il7FlUNexhOBvOicAI5U9kQ/hmR+x48TEFDtRdkTIgq4VxWS
CxT59alu4ElNYA2lS0154I2+kVVVQ+cVKWvN9o0WZ+iNsw9AHayXCbMe0Y4Vi3FI
OZ+8IFAS7yKrNo4FinDQdCNLnobjTjB0E78GEaE4PCBeGOv8mSFKqzMyFvfVkAOW
OeHjcjIaPOtXD0cnQ2XdWMMS3Ue0YciZGeKQWTWGws0e/UlvFVCBnfDYMPpBGe0Y
Ya/Rj5pbthuFn0zbEmg7yGfeeGZbHmhjzuR9Gttng/HiSKhtrRQU7otzEJ/hpj6r
0iQGVAQCBjq34GRJ9Uij3n6QD+J47R3nOtHpNnLYe/o4zPIjc6/Vh1MofGxNrnuY
9k9mYWBWPPqHvcHCgPVxdvbrBjScBKrR+SQXDvKz27OGI4Yb9NyRGtv1ayUXeGHi
datskhjhvSoI9oTHRIfpm1fKUY+oKyU9h423wV5MgTrqhBJqUFY4Au/FH/0NlWMs
rghRe39Yz3eJpcnfrCmulg9Rdbl2kXUtX/tDchmsCTcpAjHYS4TZ/16rQu0Sn717
nuccpAJldiInlski7BofSlIPxlJ7xuTCdyb58IfKflG0gQFuwsNdMAWTVt5DGHfB
odM6Det7gjb+S+uTdBxvzWnhAWQ1EXwaUETXNAy2rSwt9XQKAitBWLg/sF/96Aqg
oLH1gi6/YdEhjxzJ1cPbevyjE9fnuttdzCR3FZRhreGA6U8vYroUCouRElfiKhvR
YPeXm4KAJJie+VKRTSXRnCfnEcysESb1szUScVy653vufyJRcVOMaX+kXXQfvc8k
bBDXYtZU9bprYhxMQxD1LxpyWukTCvFsfckOoWJ3Ck1lWCJHcf9qLjZzbSII+wNK
8yWtladFbfP4/WnVmPo9nX2G99Lc9HKcdbjJ+glQ5FMXoReD0ksjA2FnUWYc4l1A
DG7ZkFbqMG+1h540C1d/49KU6E8l//jBIGeRmJsGVHcq5qlV1koeUqWHg0XlHe9F
TO5oeqCbEXHL3QEv6jsey4YX1+qHznVYVoHDyzVA0uOPaiseUKUaJZwbM262kPca
k23y0JB7Lq4TZ0ii2EDrmSgtItRYV0wZWUsSl5EJJJMJio19VM5CwXpu1RRnsoFe
bQao64frcklZkLRCYeEmFKi4gve1+EJ0HgS+INHBJEblP0LJgvvUtn38MHmUjHF7
qwyOfTWsjIaMH0QjnfU52wD3YnAaU0UVkXpaYE7gDjqXaf5pjwZzQn3V+q7iacyU
7GOCMvdJySZDIbU2ErS3m+HQq1/OvoCw3Hic4IGSdAMVULVhs9FTiypzLlJRxunL
xksYY6RR1scfKiuD72K1iceZ6VcftgG+jKXwJyHQEVEDUXLvie0fY+tUodmh1N7d
ob4WZ+FZOzBYIbOj9arbGoc0fw3oxnYCrN3KPgLY1HkviB7FpIor427dBl0sBJpS
Qx0hnXIl7ugPTag6taMtSzrm+a4HsirVow7/9FVYxJihfEYCTGqTRjSWCqGmMFLf
38ZLI0bpgEcxmpJUwPhrIU2Zxk65i7CQbsO70mfd2sLhx6U/OHxlsLvhLZYqCWOZ
1TsYiMyGijpfTwkdyoZ/JqoL4v97et3tezDWNd3pZy6JiRgVjFKPDQVw7v6sBE4h
dSGqtQOICw0LUxptES7rjTVkmCrpR8vUj764m+cUb5nVEsxs2ZtLf0RThKmz3c2H
dWTMnrK6UwnwJbF8xI8E8pmZAsO4aIro6Ht6EXGcDYrsbYF+1OUvT0cGbI9TfSb/
FQ+UFyACbsK1nrHE7P86Y3jYM/LxPU1RVnzJLikNlXmd1tAhfGkpyM1av8M0msHE
k1f+e+6Jc7MYNBAAqquyYWQF0CbZ6lJ/0WPiUDhyXFSk7wlMSsZMwdLlzC6h4+ML
X2bpJ86Ii7bo/Roc1NL+9Lb39nXJKKmLi4VxZiv7T5sgxkkj4Il3rLZUk4FKq63P
F2wLEFsnDcXbj821c6WPHXvscLEyeQF0HRH6JQ6bTIjk+XD0vBfpuE1phybm7wo4
0bJmtslOH1A8a3Wo1r42vyz8b/kl6cnala5siUfi3D/7TOzODj6h59DyMVhjw51B
xZlst5cwocOpWBSgXSTcmFOm1Y3AJOY320Q4i2Z6LbGZc/HBbYP5v2nj6FaH64Pl
lOUWEiH2CXpyibKC5Xa53dk7tFWx/LjdABBaPDSJECep6kZ7R3hU2vZrl5o8JPMM
OF634DEDrf6MSFfm85uwhmy85ROx3x0D3JY4ncEMWcUx9kHEMNas6szo0bM2DfoJ
sadzP5GO7w2kKIAtN9PslUxKoJ4FZ04iM4s+g2LzoWhDNOs4YbdnkRsRGOIq/9hI
gFKvAczhN2dt7PPTVgvjRrIVl8l8kaPXQ2DD9DmLzXEtW85yNUZX14FIh0iLkSBe
VSpki237lvqlBNcCeUcI30xYlA5ZiqA0zjNQCX5V27DDjOxZOxW2mtwMIh9kAT27
RiYeaOdVVfwUF7HSEQgIQ6UFdpi6YaAqOd/tUcCOQURGModF6nvGlDIjmkDU7z2o
3rgatsr+ZvyKKvD0+vmVELyPHKY78SUJ0LM26G/Mmp/BKu038/G5kTLDgFIebOC3
rwNS/phuGkC1imiHJGF9xiz4/S2ajKbMobc/dWXAYlgeWUI07VIo0N378fk2sfB0
GLMpR9iEHuSr1SOEAy8ZXKmVKc/9a+eDHdsBnAfWs1ul9ql+QbThTdrh1lEMDS5x
O9B3D1H9Nxy+VAzHO7HKipG/5RtvSrVUykNs+B5r3MdWm4IrHN7HZe0E5W6KAJhd
LEgGrYiGoz1Jmn/0Q49HxkHg9C77FM/nlMnPIkPIOrFscI8gPD3kQgTq3ARDhlwu
cnm6QFqkV2lVor15NqweXQcVJ6YGkau4b2V80qEjqfhXBn8VfMaMY+yWmC4eLNOC
HyfTnUCQQ04f1NTdmFQFKjDDVEajtgCC7+JwTVn9wp1J6+NYGGwtzHuBq5YAvsrn
7oSq+yYRuCXmzCe6SLAV38gB6+cnZxiKVIq2XlR7zzM3p9WeRiwh0ekARygYOUli
msh8liBvm2nSTYJGJ31F1fgTDnsnvlv2YrRlt6nBrF0ecaQewpfyn/2S0MXzM6sI
cW738Kwqd+bnNgIsUMOpgEmOq+2wwBdgdtBrlfxCX5jpQ1T4rDsSvxCd6X/tJl8Z
iNSN9eFM8JorHzSmFr2TCKa5jYRqMAajCFsW6bArewmUE3KWWZiTPyUcluOPXq9N
DJ+8XXt3TFmnJakuY6acJ1BwtpUDQbXWY4P5I5U8lFPdEq5GrzGdoU5UJVtwmYsj
o7/SPXLuh2iDpoC+E7QwBPtcPVMKamt3/wmxLoG88mzHEJ2RAg8XxcsIkDdMoPT1
IGIle3tDqnN7YI/UNib7p/fFQN2x2/w1YsqKegdOOKH/6Lk3a88O0n0nmqYVGRPO
62u7RyR7kcJgg3h0rTjQ0OE7x34tuBS/FCRbjLxBE68g0M5LKc3hZ6oaEyMLUBl0
gHvyu2zKwZjsucHyLxjtNfyhmKsZ25xKRZdfQRuEv1Nx26g3xK+R3jlMt1EX+M35
91wPKYrF5RkSfNRrYG3F84v2e5TVeGEHdinm2bJ55lgvi3lyl6nvsyKUqoGnr/Ss
EG6IYRmMB5RIOr59W7GcPLF2vMUjQKVlzdE3iN1aemGWYwNX+7hQ20P6RRDcPcRf
i+zl2a+iJspKEyk2bcecV/5y57VIEPu0VHkpn7tpzzgHX9smKn1nBTlBidzUJyLZ
SX9Mtdj/BlHxG7ldoDdMYRbKjvUPq+9vtIeEls1o4Qzffpy6RDlRL4z9NIJg4YuL
unwMPV+oqGftekJpU+W7BEzloplnYMs4gNuZvc5rMT1E3lzRVYMZUFbOZW1nWEen
GfgpFfL/505xIR6QnORzAi+FV7/6DHpTu/tl5Lo1WOjPEFKs/+2QGtfAtU6VlMDD
zAGmkwYKSQnbTs5Rgcs1hK+nskaH7C7r18yej2mHKKlT1F0hy6AdHgk1MGyxM46+
gGivYxOwGvYkzQa8G+AlWgvbALSlph9GI1/kctMMOyhj1DalCjW1PwmqA1Mf/T76
dTbTrRHCBtbfKH+N9MG8mIl3+crukDTkTxFymNsG+Rpk8nAKQMCNphvrum9BKe9L
Yw2slPB2K8WQvNTnSPOcVJ6lpwBQmq7bvMwlLwKQpjEl4bvw1plofL7A7aqg9ehw
H9glATjd+lS+zVOwX1VJ6fHj3ZYKCGJWtYSnDhZ+T8+c6mW+AqJUnQZvNYOzA09N
pT+ubtLYaQ+SsUtqK93wt8PdSERutT5nCe/VtXztnCfLcGlpfdUIqfHGu6bkO9SJ
HpWyPe76tR5cNknVAMoDa8eL/4mMkNkHEfjjzMCVWB8e8UyT5HGwmG9LcvJdkS5Z
bjTfVx1zHBjErzu8oxvr08fV8P/mPm819V7+7/7kqpNDCDLh/QIc53GK7pdqED8i
l84QrAUb9judd/xT8jW1iexSN2/ZT2bbqqGFX7p+2JYzfKn1WLzLxf2pRepPfhnJ
YlW58DpHiHd5Fo7vtUZ60V7ZoVBx+zuDGa0F1ffyo9eDD+GW6CtG62yzwlb+zz0h
KrqLziDtrKSCZnsYklwLhrA5oCAI/Mj8UW84LVqwhSUgsaq6YeUHXubn56cOEri6
beoJCjwuqMV+/DlA962R9OaN5XPFoi5ArtY8ySl80hLtty5INF5t547AxjSgL81l
4vL3RZn5qxXfgPVNQUbReWywZ34XRv+GF2OQwtT4KrGQmIv3gyB7FuyyZ7hmd9Oc
v/ixuT6QVYUGhT33IvpO1DcucLs+Tm5s4h3KJy10ke07LgYluUOqCmoFWEA+uKQU
5/+odJOuiuUGVveu1q0wGVNpDVfZK8sRTLU64Fs/42CUa7+aIOj+65wKZqT5OPI5
P6EOjHrdWJmk5yBIcbKzccorfHMehk76UUg5klADJkcdIxPpRCijjKzDztorim+B
0CXSCcrmy24NxNJulYqGuJaqz55RHT/kQgP0C/1zHHz7oZBFnHLafatdP6iOgvHs
th+oRPFkJgEGlFcjJEzHNlH1KYlEyfQ8PwgwDX3YEFi1VyuEX2jil3sJVczz1Nt8
bJrKS5qBaPubKYZZcP+dg6okj0xRF/O1gQe0CIFV23JXiwC87q6nZdN1cQlUaeQe
Z2hNfcyINhJ9DV0IEz77VnNvMgbNQigNfNOQdHZZAOdO+mgzO2Qyk9T9VLwszxyk
+8z7TGmyPr+VoREARby6BNouTqkDtHmH4znyGylB9tVp0pxxETrBwVaYFRLt9RM0
xdSHxMjGYmgcdZgPvk0eiDwpEO9TXaFjJcIdiS6GTC2cmYsIczCtYtvB6JgfJwL8
ocLlg0kQRDy7WZjDYvpQsyaSIHHv1keZ3rEIWLlaQQkaq9GeDEYPJ066y30148CI
pvjzKhif1iVGnGMIPcVfiovOOt2sZ0SOXLLGhZpHHBeWVVB2PzgOmrVUqBWs5rd2
YKAjRFlQSB/GVGo2Ms7HvUGUTcRN0EP9b9ccR5HovhcVvXVsfUdm25YMdtjZMYj2
hrap65MS+Kyt1txRty1aOsOofsxPt6G3KxzvbSjWyDuixH6qEeALsFr4jPtE95wQ
GD6919PAI2XE32YlbhRQczwy6SVOcJTli13KSRH18QQtCe3q+2ngFO9gkXE603o+
9//rrSZY/Ll/8PDCnOEtBSy685A5Xit+vwYEbAribGwnu8wHBg5H9FhikTVtX/qG
yEiKqhfQQNOwnK7JoSFfRWmUXxBp/147WTaSULl9yuxD7DRITtGk1bhTtY8kh7g3
ImCzKwY3UN8sNn+Jag+4NLxjGvDFCTky3dZdCokmGcWUsLQaloonrpauD0v92SG+
0/Te47hDoU7lQWfnYZWBqCEOsJwKJMnCx7yud6Qk18IkEPi2qnwlRRNCTKBF5l6V
IgF+Qpt4bq1IYv/ye8uQNKURNhgSdTfxk8Y6VSe+t6Xvv7mu4OXo1i75E38JSobz
OFYVipkbpiS8665RRVIYBYs8hV3vULsEPv8xFlnv/rOzYDiluAZBFpIDWkKpCCfJ
o58su5TEH5+ppVSfoCouRzoBaukfb7T1Ft+rVpZVwSrkIzR3R58ZZ1/+PP0gNz7x
cBdUSmlJyebN0cNpx1/F9uo8S1tDUJ9lhfFizk7ybupgTJUWiAqhAesi0LPx1lHH
+YZk9KJVphwuSuEDJgLCsrwBUNGZcSYtQvWoE5c6gyVh8fOSLmpegzkwpYSmd6gN
TNfkGsHRfHHAr/59jt5EgFxhby7woyBeOSo4X1GI+7v8Urc2qFpqaqcz9oXY5ER/
8otaZmmqAaCCCDOJ6c8RKd6aKL2Dv/T73w1j7rBVow818y6mTTUTf0EGGS4QGpsS
i2no/uITxNaAh//IeZ3JrOJZFEG6tFZVPaRa3bWI4vlJBR2HOY9VTIA+BZL1+0wM
i6uvo4YCgF0UHs6Czw+HxaFDjBJrN8JIueh6bU1piwyUbgeiT2AqJ8Mf9OfB3tn/
uPzkPMpvbYS9GDAL5l9ZDwzU7eOMYGYTEndIv3jiaZkTFOZAXtJdJtfXA/+fU1Kh
8Cf7QAayBwnbgjH9cpfxY+ldr5CutDzZkggYkkU3hoPtY4QSOKcwNgYYGZXbmY0E
Lg6LRpYNc6FszsseVB/gvyp2s0IIyemZBwOGELS7kPbDlYn7f+DWADTII2r/BtwJ
uSWT72E/hcFQ135Irh3w9HFHeycf75oKX7BJT81i5GNCY/iDKzxEQxlfXXM9L5Kj
MxWQ8MTmrZW0NKTvGdOc/NGxRZfZQjwsE+FaM0lz5HB4RL2MMcC1wiU/SdvWHFAc
YogFxqceSNM6y7Ju0L1molEnNqG3BuDnsMzUSTTLZW59aQI0au6gxJobBEEakEW+
YQh9guA9LrTopWF6LdJDbg9+lQq/w8ekPTM2L3grvuT178X++IW+p9x5wHzoY00o
S6+9nLi3YKReOVUUdav+Dxm7WBxXsv4FKOyqOp9x6FL1hspyx8MYRZ5yZCNTqqc1
DPU19kfhKMfhUpXQjUs4ldCWlENy4ibBDVVjC/QuMwo/e+U6WWVmGnh8a+SCCFWf
U3DyyeLi58KyWgJoSiyt2Ei5qI87Z/3qR9YbMwDPjune433Er614gZlGEiPRKwuA
niO9TkK6Yn3JYGqk/V3blYI45ycX1Kdg74t6rIgvSBB9xF9zCLXDI6HmN07htsOl
bHA3Dxhjlo7MqmxHhSV70XkEvdYQc7qYL9PiKXWKVwdfaqHBtkN+nQk3FW4f7mtM
+EMudKhPpk+Ae8pkgE+haoBfgeAoM1sypOm4evdGTDd8jtZakeQpXmw1mHSYD36H
Y6TcA/lntNNy5AhkJztDQje4KYTsA4CKtHXdjuKFEnRxIs9cnjqRcxBAX1PUVzf3
TzaGMH+3bfgWyFhgNsJ4NjVt9iNesDBP0WTFeQDwElgBwHYET+w/MgahsdBDv9vB
sm4hVrCFcJpUHPGWv5Y7aPjFxoekl12bhAD+iw2mEC5QH21sTkf+oZJs5zShvdrp
GCnG67AsmFELEMVaRfEuMLZhiA2OzVFIFd7EOAKAjgOk8ka/Jr5drqz/BY1WIyxV
+pYbNM+7QM0dwUpuXHjZTrmYjjT3XMDLfQfumk21OJYxSHP3iEuPRVGWqSlaNf+J
6cs/TFkLEbaPt91UoYnLe/BW5F+uzKVXb7KWEAKJ/0O/40fA5AN5mMU94yNI5f5w
YWCO0z3jM2ZbVxlxJQ0xedxUb7Q0+ClxMrhiaFvloNzRxC8vEtuTz4EZW/r2M2mR
55z/YNUejIzSyYpI2MfEgrN00iiE333kNAJcLw1O7nO1kag7vbDcaRfPyNINjv0W
BoXLYnrSHOhnphD2nCzhP0AlqUO0NZaD8gkT2PfDYsWzEhUHRAaQWSRWgfQoKtaq
DZS0PsP93jId26jhJNqy/5QcGocNUN4aLu7siOhkj6EUVjsUgEWGn9qAgjDH0VWU
zvUc2719YGzJGMR02aiFO1WOQuWBO2zQTAZkauRIPP4TDH5HRhHicMwHjkZL9LPs
jhvs6mwxoAgaekrmvPOcsxoT5uFfiVladQ8IU2oFDReHGbxvseyBK7wDI8yhh6xU
sZGB9DEM6RcZ9vsVXVW6rcVqH+RsMxD+43x6R6+PXPnPsznYSnmXQgSnk+QUszjV
fvk3HNq0+x7RIHkS73INpi2ZS4HF0lyKqszyTBRV2uJhUZyd5v/yyjJ0rqSahH2v
5Ug1FEdlmHMDWhnTEPFUZXrV3ioiErZL+1ZuKHjh67e48nQJpQZGGfsirJ1TSpKC
BqIXde8fFl2yTInc96Pr5HhJY0wQCBxXOa3KaS3ddIGj1PgzabDbpUbalm5Us+bm
OtqccakIdNvHPd4WvM6neKGkZwxyAtkIGTxQeZKs87g9UMRr7O77NYPb1rqxS+rJ
V1ufLTDju11t+GjEB5TcjY9NaR2700Vwd7frNk/do11gvO6JDOgKTKuZno+caa24
5XEpam27GiEAVNC58rYi1XEEkI29eLI9ouZvNrRpdo65gQCk9dA5asE0YWRYh4Og
Wfo67fwvjJoUX1rc6Py5IReNaKAZ2fTP6fWkSr5h6AV9gJbO3EiVUA/OpvaYG+BN
FkwRESTyCHMu03C8iVoxWArKc/d5D04U+Uf9d0caBXlcy6CIB4/wCwZme9mlLhT3
qq62v38GHL6NhtGxmMa2pO4WZFg6iZeLnUJss2jPRhXwFsIDy18vkLOszfvumXvt
Kpjn2O3UJZLqVoP6W70BRoasNZgu9pJm7BRYQF81lrm9MMCr88pBumnOVpBgRsO/
PoXAibI8Ic9rwZEur4kfrqimrPXxoatLBSQzPpAWyyqeFQ4F+to4sZ1xocmh2E4p
3VxtPIFkpkvvHvWDY+bt8Vwg0Zlf/A4HssHQowuJUcUBq/ogvzx/OEcYUdczQ3Pc
o2Zhrnv+4PYxUzzoiR/+BeleCtUAaJ7bxjwfbE5qxeJLMzOynrQjRWd2zjk9L3C0
CviC/SBHP6NPreQ2FC2db5JsvYseFAQ+yXzPIsSh22ksr3KfKQDDBrkx2WOEfJ3b
3x8Bb8OSk+RpH8v30IKrl/y81Qt9YUeehSnIq1q/ezF30HKsCva+MnXEr62tsxv+
zhoJnhnJ1qXzBJkpAnpH/h1s20vnkNyP+WYIuIFsXN8/Bc6F0iOdhRBCP7/Pzf80
FRz1CrZ61YXmACvb5jqB1F7pj3vQWXVoCWEeFFkTC/XPvfWpZm6ieIcb0HkXv3T6
CHFDC4+FeiOeps6aor/nQYMVwrIIdUnGHWMJhJpE7OyR7obzZyLuQaMbr8MFU0VH
krX/Jabuld/kk5IYPKhQG2ztCKuu3gsc6WaMAG9OG1i0uwRK0ulvYfEvwO4YMs0L
VajVnuPT41zDxFfwhgyDXVjf+4lQwtCLFnzHRtWWVsOUMAaFD4+kxBKDRIjVawN5
cQy4rpZc/XAZlMrNTwe+RnwxsXY6tR6J3/F6QDy34JLEU8h9pXzroOeeaYUXVNGP
xDQXHzvHdf/zs25oR5n2POHUhN5ic03pKSUW2MKzGgoFuooYFxDRLyTNC+d2+Ust
mDX+Ts/Zt4KHID54ooKNEwGfZva6v5s/TVBdYj7KGlB/jQD/qtw57AM8U1QfZbGy
DAOrki6CIZ0+ro3a+sCgbPZuHBVqWoLAH346TOzpGzoyHMALh191LDxRqiRn5w7s
evDNo7RRHqTcIj5Ohq9a2e6QhpCuNuH5aA0npx1nbxBTM0UvNoA0nlSybrZUfLi/
RbRNMU7K/mrMxSSIHsqXGQTMvS1Mn90ynBY2irPz9Kj0zkkigTkQsiknyia+IcmP
gcNpcxGM5WSGNulO/4AE8LTT0vxZaZK+FNkk3IJTHSmoPJLbbd9qDP7wskAk2QoZ
dq++dnPVRW1hrCN/WlN7dU3U1jZsh02N20SaLBb5Sb2ZDnPBeSw87G8+ZK0/8YfF
3MtMX9U8liG9LllfR/zzeCdEG6xRMx9San6T/k1oHcuIuRe5GMmOjnHo5tY3bQKd
kykAOpRbFLAbGayUSF55yMPnQsiBUrMGfrsmzYbQ8E2WdY2iQZSZ2eMtAUOgiQXa
EgzCOmMhJQAnwjguSpVN/qQLrTIbb7mJ3UOq/SmcFSvGiezAEZ3GRiD6sW9m5eB9
/bfFv4sc7ktlJlDMEDDvqJd1WBDcNKsmKd7Nnf7exp9brs4s/KOssHZGim57gdzV
h/5Ayve3Nz58F1VRErGNU33fKLlm2avmvl8/Iki76CpQmwap63odrcySvgrYdHjQ
GDI2UU8jhNjGp5i+c9bN9Cba6af/gJwfkL36F+TtiM9Vb9hve/LQhaVFzLxGqbZD
GNNutkXLHB69MqICn2FjBn9UMqPgherc5B62/Z26+k2671Dx5vKNCwYU1wrpncqs
pAmYgH3KZ8ykmma/PeVU+35H0xZiC8R7aFtEgqbGRH4zFS1DuQj73tgpYY1HsAHx
f0LSppbgaZvS0zwwTJq3FGkJ16w/UsaWMWHvHgOt9U5Dnv3BksEUoUCiaA/37GbZ
2amBTg7GHBHmzgRziOho0nj6M4C9Rwj2B7qa3fyXiBxgtcmheFPXxUbFAfMw1zL3
E3mbNc7WyMXsZzB7X7Wuhn0cPQPF1j2i73+Mgmqly/kE1kny8oA1XTDUG3j4obw3
8SNmm20o8boNYtFcE98SF74eOcmC34/3NLbdCSmr5RTSk8VSZk15ijhBKn7WXCbt
sy8fafiqcCQfVAKVUbUDVmTTimH/7xsQSITr2BoxDIU2gQxd2LyobBa4fuUW5mG3
JaELiheoeBf9mL9haZhlQTKzDD0ctVjlWu7ZN9p8+a7fnctvYdqZFX9Q1Z1m93EY
ut/GjwqHqelJ3+Kr0ci8ob8rlO41RpwrmSXiqcl5F3PDLTTNFFHstJLk3TENDQcS
ypk5MCORjXNaOiymjhTOsN5YKH01lO6BMGVrSfAI/ZC1r/q0GJ6F++YFXj6jWjrh
QAEBMwda768jLGr08wewWa/o+rD4zbYIJdbJrPFCvPgO4NeXtrptLMXVV16KbUGe
7nCWJexePkFGbLM3pKF8Qrp2eLbherAqPwpkv3AkYovu5MJ7jMPfFLTEtRb4iRuf
tOO9HW0iYnmguESFETvSv7vXGucazzgW8Duo41XgJ6tLH7t9d1I+Qk65BZuxdiAd
kO8AMydT+Y/wE/KXs1DcgQA3LMvfyGbVl2XWh6XGWmxIzRP5ipXRKySkyr15o20j
th7mxUs6tvIHgQwC1S6/+99mhPGqyTAQMyCL4LkI/qnhZKZIvikvWjXUX9xbQ+q0
VzCmIyOX7+3dmRN6zCLrfxIs5P3inhNz5CN4kSEwikgKrVIjNs7B8B8mkxNnVvT9
sGbOVUU7EOdxZpIT8Am5hdaQTcnGAsZrVHXMfyAswW8IR8Wz4XdX60R5iFSJ1ib/
aie2KMvotmFTi843Uwh9Qa4UtmJE2DFrVnklQxUeXNF8Oi8nMklmL/4Yt50vDB4S
1kavc2o3QXQGqAmQnmdMS6qwTY3V98bK6h7zuEFAgupshEvQtXJ7IZsexuRTb/GR
fBaO1gtdy3YgmHFgg0cLNU/9tYFbKnFaj6VgeSVSXZUhvMSGRHNbrdFxaykPxp4M
B0NpX10QxbmxfyL+8hz7bmKBCS3+0+D+IfFvrgjG0unjS+eZ6hP2zH/tc2iyaC7k
kRqHEnv36SmDNTKw8Tqa05ZpT7zSGKicAFrNpC/FAr/I545y0rl8HVh9E5E/fZgp
9LAeLhNCoQrTPXluhJtvWdfHqpObAv+EBbcn89hBMFWcpN8wzW0uc9gOOMSirrlc
klrL/uoVuPHWMO+YO9HUCcQAjcyAWYK2GpwxW6Xgd8zZLB3X0QmYDcFj1AD+/4lW
vcjHBK+JC7VZJNeOH5NmZhomjwicZYezMfTrwDAu+ziXB9j8i8BqeOsp6NhEIayp
Qh5L6f+KlxiOvKDnI1m2kirME64lmooo2RlDephPGk0wgVNZG75qDmqUwMxyZtpn
bI4SvfbymqgNNIodM7ThVXmODiWZr8G27WzhWYf5K9hUTBpWjYQBATqLbjBzmhoA
OzreOBABNr5Qsfp3z6JXkDVzSmx1OfWxb2Tlqe5vXgkobhmYpAyifsM+P3FLi4aC
LE8gR0uBFQ8wZ5qDwI4eTltUZfn87/Lh3k98A0aljXO1tgYABnBOx11F2TtzzAYL
5iGU6K4+t035BfwDQyt4yTyoMFdLKVmaQ4mXQZkFPx0mDI24cnvo0xP5FQN0BoCO
hnjIlwnOEHJMiHeXFaVPIhf466Vi+LWaD2K2Co4f8h4B//G4516HYNXH1mrSE6kT
2d5rkJ2RDp3mbIXXE0gRb22luWelzOOTnRDSmx5dI+w70szn2+YFTXfSf88w2Uwi
ZQP8JqwjNy8daUxZFkQVwaocuF+xIea0Xqab1FL+JM6k8Qa8uVaeGIASdSau9RmV
dp8ChU3AwVfITugEV6g9CPxNz6sU2mOwm/NIeS7/A+trFn1uOMKmjZ+V7Hq0K9eJ
lTiYK6xioAnGa8DryDm81DleDqwNpI8zjivFIF0g8JMT0x5mybdhHoVqMLYQYpKn
m9FUiCshav97I5/mE/UAEPRSbd1Rz0XxVaXx2GgrrfXPdf9SScKyvE7qoYtx9FzI
lism08Krf5pgMsvF6PzJ8xXUu6t54fRj9+wMiQV+rl439gKcKPNWjsRb/Lteee+O
/TziG+/oKwsxVm1xNIHTcf2nrEHMwBlm22diN8QaG7oOm9iQH1duVLD8L9nED+/s
Qc3uy2YYuiXCDpd5TUYapUEARa7nHUf4k/FmAXLRUmJV0pSVQx2cAEhXsbDPtHSX
ffRhzWr+hi+7AKTHsUp72AeQbzd53tZvpAjMm+qYPLhI1kgzBlyvu4g9WSDiP3o7
YDlj+sj5xpGQbnHRvjrOSD1mSlrd+X7Da5kjcclYMmYhR3UHbs9MTEpsbQwP2WXE
uqPEJEjzU71iKzegtD/cO6jSt59QceJ4oTRD8sm3I35m+LuJ+U4xb088O3kRPL18
6Jwop2heO2bv1rOqvqxyxjrB+HvpQm3NKekiBZ5otiQwk8J57dthbAEsisgSZmlV
rdwHJe4Zs7ErbZoxT1ZX0esugmxDWPIkDZPUFCaRqYEqqjMEhfqSr/SsfzcKKozn
FmUZotJLfACLJFOTD3Ex8H+YFTvKi2WucBScGyo6j6ihyU0gNFaLESSzmjHjKS1P
px70mj6U1PBWDYD5a4QwjlJkXpsX8V5KWHgs0ddsnwh++S3+gjkJdByRFaw1J3lM
Km7oud3lOlUH1+QED/0jsRuJ76ZZuLAAhDOpKgnRaMOOr4Iv91f6w3QsVSwfb+a0
b/TdK2jx8RnNb/auLy53f9bedIMvkXglt2x0HhvpN1UGCibrYFrtiwRqUWJ1Sd0+
9L2kt/c/MAjEP8YQaJrOOGq2iYyRc+IBYnVYjQP4paoa5lN9rC+2iM355U/Y6Tom
3RkJ1QVC3r9su0/kgVnMyPpGWrbc2Ft2msbJDenQ0E8E2uaMdXns8yGuJNw/lFQo
j7fyfzheQnQeGUXhHEyFBODBeXpn1wmD+Yxp4C0UNFo+asHIw6rar4fPgWeDV8MX
bgfaPbeIHFs9dwGVe14O51KP7KBgF1GvViWGraBzMrqZwTluIYSCUNVdL8u1htBH
0o3rypFB4xcRabjjQki4T/IjuNRv3bXjp2UKl7OJRwaol/moWY/c7K2vHA+DnNto
kgmzJK5O3wbG6J6QGV2Vtt15Z1B2XTGlcJY5LdKGLEmz76eObLFXrXgCpUnMrnoZ
euWQLEdPYY3u92oM8Y0lpadjn/4YvYpPRyW/Fk158DdF/Kvitil9BW2KQiL5P3FZ
jzMqAhI0Nm3azIo/dR1dvaLnubKk7ZeHGnf1mNPeqEmLOi6WhURn09td9aoqeH3q
SwRf0PtwWTMTvfnzaqW305/OoD9aBonmSkMiJZ9+UXtfrPxRNF3ZnqEQ5q8kYqX9
T8M41l8tjluCjFLecVrVptoZFGgSYc0447w5fFINf2S2h+0Z2UTeinV9O6+8iDEi
YaXBWl3HhGw6OtTft5wXgJ1r5Dt7qVlzDoJZFWx/yovRO+xzcu+BVNoUDAbXZSDO
u8ZcebU9zhN4P8ls/jTN5vKsz0uuReMnozw8QxTMjvjCsfqCRQngtGsSZC8enuLI
5x2TbPEHUsu0A7cUPH2cE8n11HCARoj8DKLH/VB2+53zGLKxqtZi+PD8akMTiWg9
1iEIM9mm2gc65t7IEYCBuyw8mQ0104C4C6myqqW9IlixJSAQpGX09X865nr+8Zaa
O/7TSfRmdRhk281H6FsTzoKDZVq6xZvUBiZZYBLr5PozQ8U+tXS3jncyqtyyw6cX
eGHqgS2QKICFvDKjlf8mFZXRcuF8KazeWjvLYHVh7BtMBaOsa1oCADhSfPPyso9I
GYOY5oWLRL3TTzBGSlsOVEDDJYN79s8VsV5u+HlZN/ld74Rj4UH2abzwL2zMHagZ
2d9vChG9zZixyQe8jzKl36eokOzE1xGubyZ6MSrC0zblOK1PZuTgLjXvAJCnZmTU
xCHariv9gm0itPF+eQ3fdsad5G5STxZwBhYzdC4MAcZNVjnPERJduanSoUWGSzsi
Ckt1PLAv2C19yCKh1SxoOVf8PQyZuGVft1szsD2c69OH/Cm1D+BaV9XTtbGUElpR
UfjLq8/y55XluLPXIG9kvXB2a2RgpYgtMEBWJ25ANCpqT2/pP61BH77c9XG+ackq
SxTlSYxuLrvlMQ+uBX5Flvmczp2F8O7suqMJTfKju7MaZrvqsKqrGCn2E+gBhaRn
PM07IQMqBTmt30QTHWBFIhYjwnIWYDV4aRS3J9E/aMtoGCgppPCQI7+mxsHG4Ykj
GF645mDk5PDoeAlgS+jon3a+6LnHPKdX9mmmlLB5GS9tY3ikXnsJGVExIiy6gTAg
+4RWhhm4wI90CI0Mr322cZ42E19+69fDtkbo+efF6WuoYNfiqFVj2OJ9tYRQXQ8r
o8gV46wguGcYMAXcKjq22Fkq04uTrlHQwxk0dNppjqL0HZupcFXwz8V4xVjLovCz
yYvOiQWS6KuR8NwuHRbEuqoWLy270vlhxjQyMs6H4xrylG5XPjBmu/clrqCQnLgV
yeLh1i+v0rTEgmqeOzbAmrIT3fY7lTowEo4x4Jym+bLIzwWTKBCOHRCtbG2E7Bm/
ubMeo7yBXfvWMmQ6JEpNftd0C6vCqUpVF0BTUTNacOLWDiRCqW1CNP1AOkymMWUa
oO0CbWsn/NlONOhM1NAoX569LgQtoGskH+87ybEfjDaom4fcDw4K44hIdfx6fsp/
PFJlD2oSpKrHyenp5a1ZZpR/1mizs2ci+CwiXbWBTwtxGD9Z6Gk/wajyG63whYIq
xlQ2rgEWvOPRk+G0KjJYkHgXeM5mrNBM9EAy5QSG0j3esgNIab3wIheXTqGE/tku
unXiLI7k0Cvh5Qs86DQt/vhanxQUlLw5Czg7mbFXsU+m3lohwFb3xJ0O6YM3JPUr
5ml9SvZY7Z20HzJ/LIt2UcI3qUweOLblXnaq00JAro1qP4NOxuWBti36FbOJLtCG
BB/KbTY8oyBOhsNN2+sRwj84ncs2bFq2N8r1hc7OmgeklE+4FJiPveaYQNXTxWcz
m1xB7NchfQbeXVFf52fW3c+JkG4NIH+6u6Hlg7V1oneQC0b4Pmhk7jhv7xwrwcV9
9KH4NMo9BpAGSA3G+uqiDo6hETuyJofulXP3PEH9Rf8f7ylnCRA3UZXZhMmLPJmL
Gac+4VV4dKDJSFg6di886RX2wgoD2AgHczOG45Fa+o6MpITdw9zQmbaPEcRv92IP
sDkaWzrrb4H73k1AjgWnKF+6pg8FtkJhoj6hKk8LjQOhHBZyP9Tqw0TWVlj0vzE2
mZzFofCgwZUTc4w+55P/ZwE+1Ym1ptw3IG0tCNjTVtwBXYLctJPYQKNIwN0schmf
+Rg3xjNlzgAlZf+lGc3YieUj3hpxpl/NzEHskfcBybTQat0WBwDO0A2e+6Fnrhf/
Mq0jJ66GqMWag6XdF9GRMIBqD1DOn7Jpe5e6CYf3rx5MhK+1XtI7gXIcSY1J8ich
BQBneDbox4UNbjh3EoxU1ff0rkRbgs7RwJqaacOtQQ2s5oivPSV0nEYouKmPqaEZ
BzKNhkJY2T/hJ/dBkWks2fXFMUD6w91z4nK9Pvsw5yI1WVm5RDcTfmTkjyTMCX1q
E0hBvxZro+JCKTk+f1AFBWRVrR/uWAzxH7pENfz/8Iwi4hpAoFyhwXuvx9e5o4Hs
ZBJ/s9h5jhyQLcolyw1SgvJCUe4QqEMoyq0+dwDdPLRASg5K29xyIo+61ObCqbPz
9A39IyK6xc//lfyZWZrI9QaUmSeMlDrEvOATadqQMseHrmHm0Dm9T6ofPdS7mq2i
7Y83IIdgxhyX5ui1mbePsUk3a19yW2yXwORWrvdBdyGkPoGSK78uqDSyPvlzVzzD
B2HFlTHn15TZlqBqU313edQyrR2JCpbup4QuL+62CUC8kY0yrx9ugk3UgJH3EwPh
8O/Uu5pXLoffRyE/2I7XbYcZT2R6SRkEEnlcyIGcjSmfTtC1QeqcDtSdu+osOdxm
T/Hwd2VaZmF8zay7n9tAnhHQnBraLd9U2WPlm4exAhA7qKsjOIocCxK/SdSJPTos
Q00G1aygy8tOFn1mClHjXn9OaXrE1G8a4VXWFMhhaR3AWdDaKhi1+mRchqQFJGIa
f7DiN9EKGZnKZkipK39v42FwW2E/vw6tgTzGWRccveDueDnpoSmDgWGwwdlSlDTr
KcAoALiQYXyK30xqqCvlq5eYFiy2WEKfgmuiauZQTMSqy/qirnYZKcpA5mlf+M+J
Xw+EtcI8kq5GLzhdf8mwdNHSgpbYHvuP2U00Ce8FZY9l3VIWhBvIvGaExfrFPogi
zeNFdysiFIGqLn3PRiO7tcDf2XZ9XOtOFEitxhXU7GWWoVUM/UTFkgn9DOUwcx9h
Aiql7T6jDvHVMOR/Ga7lA8DSSFtFG3PrzPUF85qJGXG2SJipel1UQT2a7ORBvC6C
unuXkfW4xJtrMpuSHs4NYKwYsBK9fhEGIGMN1zBAwEQWZpEVA6sC71K4rKpior+b
qCThXsES4cfmq8tja4eazroyQ4syLEU7QVZ0hUg9WGGE/LXT3KMEb5IGUto7fReC
PD/z5ld3+n8ckG4aZzvmaGPIo1E9czZRvZtAIOj09YeMuDEafhNWhctx5WoMs5MD
JSwA3JaZ34JMklV4qG4oL8AUFbXZEcmOjB5mkksrws61TgUDHY0pkls7qQROIUsm
hk67+nU7Eey5Q9QlsbDFj54g2iuro6B75ExQa2E+0bzgCoqypsPAD9z6n1vudTR/
HEQwNMkkJJxcKD+CNL7VG1w+2w1ZV9Y6tmhUvhFZjY3pyO6dwjde5+J0HfAriT2W
5p1VhCGvATFvU07prC+oZKdE66WB1hkjN5WmNiA4ty9sC8aNRFvwzYH+e5PFslQx
6Vb77CH3JcunY8neAjgca5kaqoREY8IrtnJ2d7OUO5jX8h4cY2d17clEcGIg0+og
BCty7y3Hxbmktd581NGjbDPpl/VMFFj9CUFeKmvnj7dmCwQmKV8TUnn/lJ5agioZ
ahyUxfwfFPJBV6qccrT2Ldx3jGi4WShGmb/QyqDRuOnXN7zg2Y+nEOwM8V5k8JwJ
3JzisQr48kGTJBInA6C/wJMDGHfxBwd27hc+bJENY1ws/bUbV5wnklNrw+2cfFPW
PcK7dQHAPBViDk1mhbpHrAV16W+OJLoYow7Ccg8DFXzHzCd8P2MDMnfNTk9pTqdg
dOGXd8qWczbYWmX5Xqvya9VBP/176H1yfIb9oGRYv9IeMCBJvkW0/k7kG8OAuX3w
I2yQEA1K0h83vN01QOr/KxdSzWTt7vQZoxQo8WNGg19PCM9Zne4QIcxWSYXZ7rUX
sCHd1UQ8qxpXl+PWSZ4o9l0Pr+AjaOeRYMod/Jnm04k4oXfqFOtI4FuZhcaYKRsH
5ytLtDSm+vE6QTi77v1fouF8Ctd52pz5Q9jW93jh02VUrLW0UQ3viRA0RbtY/d0n
qBqg8sA1suD7J2ptZCxK2xRjroZUgtGfxr7tqD7NWgD3JexUZjybIAWhmjO0nGc/
MFr5/5JQzUTMQuqvKewGtKDL18susCYpIQRtIVmSbylxmXXktCsADJE4YbzXmjTK
ue5a1Cfliwsrp1GGKsepepoIb8xYrHpgRO6AsID3qGewVy9RETgMoqWroK2RRT9L
w8GFwTSvt3hzeefXM7NKPoL8UFV5xEB105A5bv3na6TxEthIoGArso7ci3T/pupk
T8gY65amze5Fk2Y1wtutP/zF4RfucM2/d0av9kPmIS++vyKobGH8yDAuKwSDMmYr
RgC32XXYY3TPdXS4T93/ZwlQyDVuEEVb9VrISgIiCdEtPBguyu/JdPGl6yy2mdO6
WyJ7gDUSHpqyGdVUlhUmxRs1nuzMOjMJoI6BsrpvXwlN+kdBKyX2dmBeTgYCgnZx
sXWDVk2bn5V7Vc25ZuST3WyFJKxvoEx8b7qm5DQVQZotktrRy6vKFzw/9QLUDOdF
97A4SpQhRyJyX34bk8rIJfg6En4oD8K4dXf0o9s5nnxq4AHVZqDtWXTE2xFaSFNi
fi94wrLRFWu6s4SZOoVvwSIYLZuig6mCr+qqIWK+AvWSbsmZteKbuqdxY+Dydl3Y
b1QfZiJIqd0dYVnp0nMzOsPnOQZV69fHnv7jPVjff/IHb9xyC6PVzT5plk/OqCCj
LCVJIXlRevTJaOK5wD0+wE63nZ8TsPLV5okxUhBsmO7cFmwdtf3lPX63jsH1e8jt
Mrj27z16Xwa8XAsvGtoA6wVmvZbgeObJUBlQDcENfRdN9LbA7+8IHWgib9Giki2V
FqW5tdC824sZK4WDjMCnwgkBjim0ad3I+CJfUspeHg5eALREq+OszXN6zLWkk9X5
I5lRKrwIZjdnIaOfU6vkZzNwb2JApJXj4oZKoozX3/Pa1RrkN4scUSTsqzPcvlYa
fSDJNgr0gK/sTqNu6UmHHZ3Kf9lv0252Kah7v+L9uNW/7i0OHM3OYidRIkAva08+
eZzFcTKBNRXX75mphs6GZmycY9u3UBtlafHh5V/7srhDkCOWeGVvYSPRMqEttP+3
cMph0+rePqI/JK8xzq4jQtXlyIvHetdT7WovzgVbgJ4tzHXqlEI72VR5S2nKNVt1
4Y1YFvgeELpJCjsjqoWFCt/ksHmIuo2k0XScLdMMvx1C5m4vMIEVpduLK4kUiMek
zLZrhhStPk7AvAiz3j2s/bp7hsbJkhQikbt8+I2DlcJgRy5F8tUeClJwVoPP5EuH
ee5zEoIW8xVum7QxOJJW9ptc6u0u9LJJq9Rk9AprO/fbQEzqe+6P/qGVqX7UnkUf
Flmc7KfnvT3XUGxtNUXOXiXP61sFcv8VP0K8ajzed59GDxtWtkCl8m6e1ER1r0BJ
S5kQKsRDb98C+DCg07DOcV9YUnQo9f5TQI3s2Zr4HfLFsS9gWoUJhHFQVmEiqR3x
VIQTpNCuSzAWgCusI0cICNPJejfL9OOJJaF6zNJKpZjWVmkVPiCxyPbjdJLiYIkP
UVyAXFDoCNy9cglIWtlujx+uGdG24/viSrI8NfkmdEdl5EWyVbLqycGQRiZWu0Hi
5W8DHxnBSBgdNBxwblxvOk+Ytf6maPVvewLZtpdxm34+TN2cO1RDfrdH/xkDOw+3
sUJFjGg9H2u6rgq/bT2kPbtaofuCmf9G0FrZ0Pt9bj4sK6Tn+BPR1Z5Yh/j4y32e
eAbtycTdN2txx4eXVunAvLZw3u4yGbf4xq1dxIZimQYp0XhpSNMdvj/3Ki1/gCZN
UiyCVyZpu9bY0UrIjR0HqDJGyCNKEX7Lh9N/0BoLfz8dLCrSiqD6JcyutC23JKUj
t+Zf+OZ/ytzMYarMlm9SOK4JFLiEwiTLnfKfRnhpzevKoCHkyHarQbMTQZkBHYhj
dwEVNbbodTHEWoOTh5pV1TLkCC1AIGG0tyfEXF7ctb/WLKLulkdt5ZtIXZRfCeRR
Nn5WpbrEzV+Knh+N4iLMazMezrXgG0opQPO4/RwEEbkxkCB9ka+SuyKU2bBkpYaz
yh12EEIb+N5dkypJ+jyfPyM5/zYzcizioIbWCQqBtuHDImuIlqyMLh3WO5i4pvK9
dYoNqWuJohrr8dcRcMKpjOyJp1G6JlcKMT4Ts7i+SPaVjdDMBQ9wv8eljX4dgfCO
UQoK0K1hSpmHkXSVRtNXmCVFN/TthyTYMJv5r7BqTzVPee237Iz35aZwbb4Nrsnz
7FxQHpZjyar1ux4yWww/bCzMjYOu7o4ToTN6XMuQACTvwuD2WhF5N/qHrrgPJFv/
pD3DcZhpmiAn3PADTo5XMbePdFPXuCUWaeojcblGMUfoct1EY45JdoqPj7MKz1cB
IyZxH5iIMPL4dU7oNTuWz8/q8aDExREIIkhuMpPGUVsE7BCvCBznF73ZxUoZ4wSm
UwnXFOsjtX6Iu8afn1NIqxTOZp66jfafpZ9SdezQEJe9PeweQTqIP1UrMmqnM4fa
IxyY88pzwPt20K6VSb/eGRXVUZJvc4m6p5t1Es2WeTc3wD82QXiPNpl/JeN+ZCFl
EXBcrYO63/QaMxv+lZn6xHTzo90buhz0niX4TOCFesEAs4ugiBGP8vXC31hL2kfC
AqARt3c9YYcJKbUCN7utLf7Cure3xfMKMByvf5kKVeLhtDbYSqRk31UZcpkQM4Pi
8mtTcu2V4J/4qcEFIVSZQ2OL04hYXPd0ZJadia+4/trts2QGQwsyNTBlE/xNjV1b
mt8mYM9xTQmI4swQk1Jzi3LpyasyetiDZFL8YV+OxmXhmFZ2jn0ZAblZni24NBHJ
2GNo9k/VFcD6XJ8njj1Bgdg2r0XypGPwvdh3gl27ccefjp6ssdROfccscPlgfcoS
d8HIgJT1y1CECGy2IkHQeI4X++wTDszA2cVKRT9WJCbgsqszDUQnozI2SG8BBMXB
YiGvqSLJcPw+nTLI4ITbIcbyRlYhlY7XZmjjmoCVGJAQvWqQutKCoRKB9S/nNWS3
NSYf94WCT5SubbLfWHKJ9X75olBn1JVsDty2bc0zJ8GaeQPslOWEcFOJZvNYTyOy
6iH2k9IiEDbT8rtfb8ypklthzptnokeFOXOvmwma+CvMSeHrlMgDGfxQHGWY6Yme
nlJIQfiEin0YtJV0BHCKTJBzNwaxcj2cYrxeywxkbgIgrAJt5WdcFA+vMwpbvoIT
mdECt73+YK/8FhfShqIVPr4r/0i8BxDcBNXnLgF49nlWNcVyyKxeWpfJO7BZyYaC
87EH+dHWf9mm8tNPQi+5nN6O0P8W6gHe0joPDRIfD/+5lDS2bvro6CqBw0Wzf3oB
IP7TWqXnwtAAzCbhw2lo1l05jgdpHgE7W21sdLJMWuSvTll4c+Bzd2e24lX4fF/+
LPEGAEOw3Rz2TmmNDO6LRIb/rgzq77p1+KQ6UY2dojGk+JuDzL77h/H6OqWVcve/
8jynAT4R3HRdYxDIdEKWat1Na23F/wBf+u4ZpggBXgjnnwDdjvSxvyPFNqno/ZCF
b2/ODljyeZZbWl03ewFeH1VrqJUOYSBTxYyM6sI95G8A0gKJ5hrmmnaGyo+NccaE
7QhepBXTGlr5w4QZ/IL6Qbj/0sa9b7sG9Qj0C+sB4aXqDjIUmr3Q3otk9FzUJubm
MaPTNH7xT5nLyAzrD9yhJD3hpBYRMJ7rspDoYjNMpY42UrLgXXEn8RWg7eqfY7zB
/QMpQZtyej3P1pZ8PmMJsd3K739z3J0zBOeg3cYuEFFRz/YQOl/jXVuzhm7NKMNg
EyVAfnmEcPxDQbzcsxeJDdfv6tGL7eiZXZVKyQwTzsvcfOZSyvF178qUZCCv91+4
EFnqG2CYvVwhXA3XOXeqIyIoPhrQQ7KaHKV3SWevF14su2KsBSuLwcnlqAImrKM7
cLmefj9N16SQZG16+t2o8lesrh68SbBx9AbjNW75esUPsvqVwvPmwvznhnH7VdUR
b+ErEkCiWVpAccc1ijucmb41uyAr9EVW8HtYiN5sTEFndY1QapNeyBAsv+qzwaRB
mEG/QFl2JikkPC/rQqPTGSKMPJM/PdFjzejeU+ZfNyHzBrOq3Gnbx11kU0qFwWFY
5eA4vXMUzSN17J5puVZYvsyW+saXZ6RTPZHu4fB95xfASLzCBhM04yMDKAtHetfV
FJPGiObsw6WmURqcHbSBRQ6VM2uccOTnjhWZcNtB9C3W4xm/skTe5b3EZvE/f1sg
YRiUFTdxjT2IN48aX98duPhz1ZijGcVmvuKzLy2HFjyNeA2cnxwvSrAmwH9qIJjA
DP+fyNKiclXgz1+gyF9/XXI1M73DkbBK5AYVR+MjmggQacRbH7J6mUT9m8MgrMmO
Zd7Qo0rnRf65y14/IRVWNqfEre06mwKn9+LbSed9TSvjmUujtQKKOR5qrOQTqI56
i+b8NyjZ/EdQ8y7AxSpJxOqTsKCXaijFxQniwzVTatk3bLAAare+cIqKAuAFUZM+
Q/ILbiCY9pG2cJ9OuR30HvLiOEpT2EU7gJ/Jvho5TvA5Y4XwzqH74qb7Bvl/6SwY
oLHIqREkQ8/1ToK86zVjfjvBWgm4hqhAAUm9L8xsnMN0X2hdAsMXoVsqfO/rKFyv
m/27vThCtHR1dzDwt+ObEUErsJfdjWIexPB6O30QGQkS7Rb+f+YjPfpPNUiICqa4
XpmRT6g78DMJ4mmrjvDbrfxlnBp8iWp3DwXHXP8oquAwwsdPmWxb7qHXaUATqpvj
QMiP7EVwSGDKDB0MwBQ/gscPCrphe7HH3IuqYxc/vJ/bB2nlnFLWEIsfbrBxM+GK
GgAzwQh9LDypgd6QegK7jBIKZFRoGw/7BuVfNXjNU9DFGuhBxFDWWB/brktmO8mM
g+61JZAaGMmmCgOiDJuim+kTwft/QL2rcU9XUJ2w9kE1G+ufJVReUQZEYoqwFd+R
rcdfVKJs8A75YZ5dMYU0tWT2q9pyIy7SRzQpby3SKHlMDS2KLOJLrDyiFc9nBa1s
JsWHseLpn3NiZOQWZCJWHPceiqMQborMExxhWl7yUnSC5uK1KoSfgIw122D0/Y0G
YdErra40dp4j5ejXOefxL66GRLlEzug3i50ZWzdIJcJgpVD5bYcWBhsRhDABdcXt
46U0I00CTyCKcKe4q+hPj6z+J2cTtJ5UfI3bNdG8PBoL1++iPs3H75sSLe1TWFTy
XErsKQpsvcy/kc1Ni/i4RCuXmgP5bT1eGn7TYzQX6rRPFbVKsSWL3CyJmmJsY76b
qk1qYHySgbjatrbYFdi2oqC8f//dMsYJbnirF8oUUW5NXlA94KHlf5RHgntnAZMD
csnCx9dk73MLntwTG3lVqipgFpVs+FjSaF8HnpcqwJBjwy39B1saKhOc/nXuw6/N
U1bYRVhbaycDQ9HnlY4jFcevRFj9NHPN7qjmm4usQKkMw7yF3LmbWe176mbuuJjv
LVEUMcsA4x68mhJeFqWYwE5C2d8Bj/UnKaT+AnydJTejp+WY04jAtIZiNkvDegOA
rXHFTLcYkF6fdtjrp68Cnj2yp+u3vTLEvVrbVhFog3RuU9b2iHChgyQ+m0f92Ojp
yDwZp3bZ5UkwzOhfaiG2PCQnMLN1CCa5qNHICxj2hWhfeAQ4lidphKP7n6WD02Wx
K81qlntSt0mXy4RFuLQBdt3j0Ct8Sk4E1mJIx2SxZ8FJ+ED4dTdEcLeaa2m+WiNC
6yBmJCn67If8ene/s5YHQer13VrwiwcUu0t/F5HCU8dhg6HioTTQwVSwFMFr595e
bBPjRczuA1HFnnUX5JOz6ulFhXdmUF0NYTcPI6doDXVSichkDOI+urNqbXdrkNlJ
JoqdHX7YeuqwRgLjk3/K4jUIoOTNXtqkhbP6zeRpHtpu2+3HMlwKHqwPgCSvnQsm
Bqn1o4xk17vVflsWdQ+4Z4ILZWZmvxdyObCX7K+dFl5QwEQwDfRsV6hBWs4MiSpv
uGEL8VBe6kg7CiPe1uwW88YFCMWuQApa1HHeZxuin8M03vDk0IT/HQHzMVp2+Tz5
sQ3gyCU4zMBXvH1OT06K5b1xch82QaVX7ySQ6qxq05zv9nPOP8wXPldva9n+fveO
yfCOAoifRzHMt4gKspIxOpb800la3UEoNSvtmMAv2pOKfsDhi5G3+InTcnbCn1nU
vJVjyIubKbmGTvLcCeCyaCwBHez1Xne2HLbAhLCgF0cRejGAG6QrVK4tpsnQv4XN
2Ji2LmGg0s9xFzBa9BqZe0JLiWL2Y+rcjhe99LLPsgazycjYwpnzmzB8jOhia1KJ
6h79TEyuklf8OsdNe4Xdn+NAeeqHMfJ10krloROeRZq0M7JW9RLis1HrVZfuBsQO
fVyRQJjpSWxknaXfSS7THhbDE1N+sFe/+WbkH00Pj8ViUDyx7TQnI1zdwrSW4FSR
sTBiineJ1eRnEo7aSPk++GMUPWfch3T3R/8JwHsPwRzXnJDUbzJzmziyvpbaA02M
9/ob5dbhnKhTOv4dQ6lp437dQef9fLjwThzlRSZtcuNoooPmi6uXkbaaYCJAmmv3
eIFwLX2SjaWbuZVeNc37dIHP9t8LkeWCB50enK7npCZmNS+R+Epfr1oRd0QBfEL5
3iDaEKW0alwIsTjEmJdj/iM8TLCnxIkywgZ/+Y98qb9SA8W1D2lU1TGiAM6bVhS0
SI1bpauQ0sdQ2LBonmGc0z3RvZ6Z5H4Ir7LOleIBnk1LqouPGTz7TOkm/IpYpWr9
VpT6XFDudW0OAj8Awq2QIsSTTIj6UDt0dVZ/4u0L6mFaoHv5411+uc5HWVCDfkeU
03w78pWoqYU9R/9aJz9W3v0TijVloFN+qwytejHfM8LkkCG5Dz1nbuyXbjFUXfO1
YydlxeGKKf52AqdnFdgl9ucBzBQdtMySUxp2IRJ/vfXKK2DiQzAsZckxS1yGtWL8
1w+5xFTwTS83/iIxvnDQIvc8YHzQxaHgW7EswZ/gT/3xXaJqnWcAUUyEtjBe7Yry
HKsVlX+H+Tv1m0aHBxv106W9jiX6LXUZZKRUSOQZQ3UlEB69i1Ts+YMPD4cG9ydl
WeSPDf4yEAU37chKlVUXpBwHUKdTIOUyerCpYzxedVaThj0XgZpKbhPiPLtytRS9
+rPXy0xlXjtDfneLmZM+Ly6GxkLp7lMOLrbRl1w4kgb26w+BrRmEpBTCPozXsO/G
+3VxGJuCJhfsiZpS3bIRxqDYQr/+v276rA5CamiE4hlXzv07rRwilkUhEXbgsl3t
WRd6lWFAA0sOseRbPj+wmZgJh78e5mjwjrq54ie4p8MzmSLI57d88lDCmvA+Bjko
oXN2ZbZDow3QhTXnZ034Vah6p+W+5eKJXx7dgkzxa8WjAZmoL4CW8XsGjGSRf+/9
/D5E4WmvtGweKe2BllkrqWa1+EyNU37ogfG5QYL9b3JYeGv/9LTIadRFIWr6owSv
x3Z74aZi9TdYa/nwIW/lmfMn8kdLiYfbVVxtJHZXAsSwIW66c0H1oUkyVgo1raDK
O4WKli71D8QZ5iGIrrKVLIxNdLldV7oQrfiDjsgia0mkpY9dsLdpBBEpJTKPlWsu
NhsQv83QjuVudOjpM1jEw0ZNnO2HbaKzoKJqg2p4AtO5aXJ/cMuv0WyurUWm22Dc
JPNG5jDPJjgpoPDHirlTyr6rueIyrnMQDvuZ6VHOgjgkETeW8mfeG8IVANMY0hDB
0DONX4DLitwYVIRnyZjEZ616GQz92ftBJcnDE4Lx0vtZalVfJ29j4Z0gGooOPSTb
nAe9i6P7SjDpUowQxLXU0DLch2Hs7MmKvWWlRGTknouMWeLI0+5UZsr+LoQe6k7Q
Boj9Fx3CVvAw1vfAxHT2jjqVJZi18fhaLDI8wCLFXRbhvPM+FlQlTKSAxPkq1+Wm
UjWT3TbvAfQH/HLNcXNIjmJoe9lw+7ogcFRSzhKOJsrO1bNQULfGccleCo/m0wqY
Y6VF2wyIsLcr5wJ9mAQL1UTgtINPeb0W8FjdKynOSwVa+e7PbeVEggl3HlclDPk1
VYVX6taDioGDBre7y5456qHn7MS9Jo+nxH+fV4DTILmoobGZGvYns4b3s3qdtXCv
wBp5Y+/zpezIn6MmYmxspyNqJTp/paqw5Z2zJ8+U/NSJ9b8GM6SB3h5ctaa7eJh3
K/qUSVfVZKLWNZdYpf/KwYqziittE8F1anxKirgZcqoiy0w03H3m9dfbVKJKqtFu
1q7DC4lI1KLgJNgx5pjEtLYEjnlPNhceCjnAU2npK+j1uan9dZHLZ1LXDtpgxs6V
uzaaZXPGKPwGUmUp4aBQbG15AccnHIf2FxhJNDMG8mLkhNhA1F++BwYKXcATNbkQ
fWPF6eAa1DP5ExQM6hdUZlwersQxjUgTEjMwOZ9S+fH1fklvTct1vi3nMD6ffh7w
bKgWwSiKxbZBm8/u6WiQSbE+HPGLvE5EhDnsvg11UF0z84mqFf3NBtnty0vNvgOn
1ztVaNnHwi2UoMzN4zLt5jI8dnTxexjkqX+imETWpJb3eR3ky26nUHXS5m8PJRhJ
0paocEyh2srHA1S8yXfPCqve03lhTFZb6S+eEiKaqDZK7AmaTZdF8/f1RHC6R5BP
J/koZZHai+aK8YIeXfhboU/0r3tAyX/ggmuIiYqzEPRb7Y2vdwgKx+5BvpvAO8hG
Upkgt+sCwv1DfLCHdimZ/uGkIwvzjQbBFZpjHV6/7dFfchy0nvKCckZe8Q45IVhX
c08y05xfkmoyBb8YeC84PAwSJFbzZABB453SUQjVGcZZ6Thq9zrT4PsEz/zgL7y4
b8k5oE990BD7eZYHkxWI8b/eeQ1rtlZv5pXwpVHyDPTFloZcQPbJDDOcWoovwlI3
NUFjfRhxcciwhjFb3EwLYF6puDbsnx0bEbeDrvjDm3rIXsfYnp7l4D2pcx8OyQB+
aEa+trzUfJQ9CUXfCHuyeIapNy0TcRg1JGWZw0qHe8ALsaeFD7rr2k+HjImEK1eM
Psw3q9LNpZoZjHNDJ+LETlvRRp7B93jLPLYPHqLtLAg10wWhS2VhJ4yWihblWM4q
OXA6PVbXwXiWbIiMSppK2sEkIJCrLVR2XxdY967w1TKuLEIrXUmsPzjGgNqGKQhC
gPxqGQdvPd7jf/laeN9m2T+reLtZzIxk2l+EQL04YnOXgl9EMv/DNor5BUW8oSzO
bpncuJlRuKnRV3TtQXSzHy+5BhFg/bgxT/a08YaZTbPA75wDSR/bPeUVluexdOmT
VSXrSzdy0zmRi0KKxFAi+T+/W1zdM00cgVXNsPqZyal+RMujWdqrOpH37v4ZMMp0
M7qxU1XHZvGEk0XmYJ1r5ukr1NR4TJU6FelfHEgsxkpDAMd6KIUaiyV/xLS0ietq
/n9I5Fx3sCU+RNz08mQ+7XgONpg7lC3aY0J8Hv8hij+inY3e9QhaDp+b395dyWWI
GYhZclUqBpSrvmjnOkVbwcFMWBiad2YkpspSgj5AwSAAsP9DSZ9HPMQnFzmvzQlH
5eYFvZT7mUkM7eTRcOD965iS7x3wVt6bzc4/pwIiPNmSmhfdHzEWAjQiiHUsIJk+
w3CvlZWCmz3YBWbGUxjVAK7fWssURzjbLDES2AsOAq4LvxTuSfcsqTFXRk8oWc+2
K0dPDMp8sYKdjA5InjIkoFlPraAAtIetHXJ0UhlHtOV8CAy0OLp/IIoBIOLHUfCS
XxGO2Hj4G7Vz0AV7K4HXdfgzvWSpLEi9o61C7sl50SIKJiIFrMdty6duWIp8Cn3L
0Fz3aP3rogikifOz4MZ10FVsOO0xeHDv4CXxOx+9WUJo84YQGZst4slKXVjwG8Py
H5eXRMqKTALwhvVoVrDHyO58U1iAs29rIcT5wOklhrSogMvuOJ2ZNDUrXLiitgxi
uX4miOB8wtEJi9lQS88gHU+fht+a3InIY3KRvEH7ts7JvsPWSYn2gSH/TR0ofZGR
QvEXXdq8PBzoDlYZh7SsntN/CW9vsPbyukCLF5TgYQlHYXxk8GsFsadmVDpNjgJW
D41TnhgkEMypNENUZNVkxxWKx+J0YlmmbgyOo5LqqS16ljsPcnwH4qOTz0lkI254
dvrMBWOKuuKg1pX0XgVS/dg/iNak8T9aVLYuP9EwdWkth3TXqJpsfpN8aRzrDLzS
Un0Bd6w7O4wGv7VujDB1WttGGyBLEeMGIieL3eBfi1MDf5zM8wxQVW3RqfGQDpU3
GjrUbddupEFbBo2DoJpitMTnJx84iE7OG7qgvxDT4cgU1/GAIdD2UKCVwt4TWYHq
B5gvSU5VGVl/Ru3V90peDaI9c3G8WLYFeUks4azydxBsvNnEv5gq6Bf/PdjIc4jl
Uha4z8YzDkA8YFkMmEUxnLq8KXhaLckrq+gvBmYsx5pESWy1BKdGXXiMUtuP41en
jl/dqqKY4tLGEvim8p3M3CAhevuoPvci47VTFy9ISXqdao5TwaJZ0wdzpo1xITJh
5OFBSfszlqsF2EbC+nzj/rX4Z50O9JGAPkVRkFWUu6wUOMxYfcJU1GgyVASvqMRv
y+FytQZOZuamNT58NqxyWMj9vl7q09j6aC3gsCneoAyq5nO2n9nSeTqtohUp67wk
GVzUxeTvGUtR2FHqZhKB+O6DPcejBqkLg0/qldIhoid1NF6tn8uHDYuuWA6oEa0+
f15KrrCYGrlmCbBVr7PXfUazHNXO2UFYg9aSLx9TzIBrT3RFedkGhwFZhep/Mopr
6cNYk1qLW3nS177t8qIr5lhi+hxWi/a7yUv5gZpmEuNdUaRSPp8vm9oseZ6bzyTW
uLScHtTy+MTQtI+C35zN8BZvQj5dN0Ea+3FEYDRIjALMimsi9XB/ndeDWIzpLtRt
5DeH1AhIqXStK8GJbQeJpJOsXk07XaSDwSNQTSTJfHJEFsbAnwX2KxBk24N+zr6W
38/8ujiIje0iuOzG4OC8i50PfWZGdjEne+uLHukIQ5T485Z7sXci4eR02odzTDqb
YdWerE6dWd8wbi6OA+029G4Js162phixw71eZGpnZNxhO4bST5ZqO4P0+I4uUpAJ
eB3G6iK686b5Xd8GpX7h0b3uacIt+7gmtSj3UHmdh84hLWf0g7MVoAVEM8s055rr
GnxpTamgEtLoQJ2SLKzidiOoz4zm3kt0hcV1K/BcW7w01pPFqtSWZb4vNCJ2vPb3
DQqHst8veaIU9ystFukrUrZt7aj4H70rZsfGnILOFYGN+WHklX6tCNlhXAfNsWWG
ucPEbl3MaSJEuPMsMhLoKSI/2uXP9lkuJ4trG3eJDpJWB/VbIezIPdFw6UUDhk9s
ZEDdvRpz1qdy09KFHJ3uAdTVLBl6CX2yyj1KQMr9hFIYiOnSpPhZfSn+5cOxhlm9
f8jiT34SyCHq9t9Pczd68ZM/CJ44Cmxr90MFKCLxYEtWFtP9SocI9dTOJCaIuXfq
LMhSdyYHXbpTLL2elRwxwMRP9P8YFaGBrtK6pjvq8fX0g8mrrd+mQkbRXd0AKSQX
3PsgenmDqtWUc/6dh30j8i3ijF1+tOFZLXX8v2COdiFUJDEaUia+SG4YjF2xgBZs
G9Sxj7qnqTXMkKYkK0q1dln6MfCWbJBoxjNPQnxQC0jlj4099NTh1hVKUTGT8MOd
3dVLd8XQRJSKcv+1IEQjxj9nAJu0r/FmU/pi0FNIxbnykNFJbiixj/CNJqnoXdu+
ddezQ0igKvZ8HmiX/0yvcISHwYCumaInT4o3ZnhLhNCmaA96iLFUFhCFl/R2tqsK
YuOMcjhv5f3o1utxPYucAvJ/EtK9nOWkKnQ3XIZl5DITL2uvuMPhrDNLM+YKiyLQ
qRl3mk79wZzrR0iVTGbubYdJ65/iBP1i+4EHHXWXnn5WTrSPovbb6DFsRKav4w7z
CqaIxk05+VHsXK0N8DX/F49RrYILFPxAdW7ThGii3sAwyi88pWsjTup9tHJCN2+y
2pFvAGFVfacv6Zl41b5BcJ4J0W4WxgOs8+qdNq4/oQBAhBJd21+3zyeMEYe00WXv
znH6ld9iJCiwnj9ZN9/s2oKtvc1LUPvMMVfEVprxHxw9Rs8TtuF154CFDx5tAeLq
p4+lR1ZpwplcI4DDfbmJKMkK7zRhuQ/QUiMEmjyp6eDo2WpK7W4gZTUbE0wGdrZ0
v3xtXtMqgFcteCEZlSXqv8u09/3uqMEmwOLrjSKiH7Y2DNC3OPC6hdEFKd/YzyME
FVYVRAP5xo6iPGZmh6+g73pVChUrt8NTfUCw5/uzSCNkCd8UxNv3FketyMsqOGAa
vQ4Nzz9gyLBEWWWX94NOUX4g0izGhMQ7DKF5AM+yiFPQaUxObcZWUqxKDxTh74Au
h/b/0fY/4iS7gm+08cCyplAZu2ybdfbSQI5E0TNyy5e57JZY8LGjG1QefCBR27nV
GU5o2OOOYIEs5yEdoZOeOSTRE0+aER7VbGHH4RwHluY/sqwXap9zYX56EOLn7MiX
3coWGdeAaOFK06fl24tAIr4wsPm8qPOlTp1DVSY2+TVE32F8md7BX24Dxjbc4GWF
vvdBFj0RgkRljctLR6Eq+R8YglfWM42UteCA/Xnw2iCkEinliUMCUJ1+y2jQm7Wv
YscUed69mZ1ahkkSLQcpG2k9GY521pDV2ifaol7CGSq4xJPnNJdKyP1GsyjiudRe
B8URqgxjke4mSu0XZbV1JZvqOmTY6eA1B6NwfmgFRZzqOT/L8/IVU+Tp5onELFDE
/3p6dmYFMq5fgnuME6z9+MMpU5Z90ztDDKrWMFkvcQ+4bnbl3M6VVW0FxYhJHIPt
sBBU7sPfFMBZbGBd55AUZ8IjR0XlJz6ItJbVaLTnoU9+KdXHFsjHHj6ZogijAoDu
xB3EPFkaM2XQT+br0joq0UcKOE1ToL4Nf723qfnRKYxABH3fyP42ENvcRWRxFRun
KbypQVk0ToMqshx5Dn/SHPGfZlWefCNT/cgpY5v+WchrBLibOJImd9ZIR+0x1rBp
7LSoK0JiSG6Wro8Zsao9g8m4DiIAqFLXSUD+WNIeTwXMuS/OZrRsB3PDbAjb71CH
mlmI489iqA+6JMU/xXoos1sof0CJD7lFEcgOdyNnSq/Ib56D9DUmqLfyvmKKnbYR
UdNHjEGPLMQGuCn43bD5BztS7nOSG1kWOdaawedKVFy9XbzLOH3TbG8fPsKBGnHf
TyJoorISqEd+C8Q/KFYJX02Hvqe5e8E5e4mkqMe06UfJSpk8WWnjU5ytY3BQlrgo
G7qZ26P1JsDRMkX8vY7SEec9xA3RHzDLLV6mHDf5gKMhQoOIhE+ysD5iAi9xBq7e
sesWo7SaXY3vH96PRAOeuuFN8Vu4JRmKuMNyF8KeVYps10hwq+LKqyaik/U8mBbw
Wxy5WX1DBSmF5NP2jrWigvM7q4nBzBwpKmkUsrPuDp6YHIRtJ4vf39ufNj7SiFie
V6vV/iKTk8cM/Ng6RggPVLRbA36wDyI54xnrPhVenjENkBqoZZgia0eKvkv0ar8M
M9d+2g5mdUC/O17Lmy0pgk3WgDXFhUv4TREbwUlVQQuWZENba3QhviqMW5/6ULYW
Gtx/I2Cne9VYk2nFxsSNA6H9EticJgXicihutIigRgLuNQEV2AOmCSqsz+Phcz5z
/UNjxiFQysIfxd8jgCldsE2/QYa7ANkKMgBunceAfvEAb/l/hHrf1uWAgaKGMuxO
CL29/YdBwX0qbx4P5X8xgdt2kkybp6SRYQEU/IXWhoapGTQmgAEGa/cqoQKletBB
DvR70LQsT5i4bnRIBx7m73GT4u7SfbAIXbnJfIJ9JhRRwCwKOzymfsNzrnCqXCgE
yPl9ICN5M3kPSZSBQGb6NVTJ2GE0faQ8PoUbQT2n8gQRk0IrhzIcwWK+jbrr+LlC
ZPz0YMJfpeY2QQDCeaaYthknD25JlC0Bfc9VTgx6ae1WDX+miQcPvzqTlLIobjKf
mSAl/vJui35wiUPBotOK8YKdUFchv4g1cOtXR2sGaOp5ToI8u7SsgcK27FprPg2V
hCeOwq6aqvsEWXejVHDFRCLUKVEPt/xAhj0FXJPK3QIAj7VeeLS0hjgkRmlnebx0
fWhUGRU+EB7O0nrL11HUAfOZJx1Mqgibz+zm7kDIAgmlU2aqpQEovcea7BOFXH5G
d9bZ17RrcR7GkxuNFLveZOvMqFOmDdyIrAogFJtO7UUTuMMxdFvhWIT92DxNKr6r
vJbJolo6stu95rjIbcdJ85OYTIKJuYeKVDsM1KiLJwCdCg0SJnzb4HSf6KjiOXY0
dYN1bbE58LCkE0hdLpMrGTWehARRlWVE8N2AJvxzZ8rO4BSgcyii5+F3bR6fC4La
G2EVWmMzNWpFo+n9ighFfsDQweXA7qWJmT4aoSeJ/MHyFccNpVbamXLys/LKL+6I
3/GFitgOnrnW+jH9i8EWX0nS2exN+1/hxn0G8Pxza1G82r3yg4gzrYFaiFIOtQG5
NG+ihvBX4AJzV+s7v0O+FifqPr1yXC/+W3Y1MEwUXA2HwX5niMssjnKKTI/tyT1d
tmNvbFWEikdNqjvaDvgxwJMQsM8niytd+NJE1fQ1nsZ3LxWvXdTDE5ycN2UFMnl5
dJWk9rJ2Yc8P5qqbSBwm6H7lCFInJ+PoQD1Ou7BX8g+KxQtgEidcPYu0L2MPjURC
gt7U6Sj3ETJ3+jAazCkim1dB1x9LxjBL1WNGEHcknhNOhFlRzvpU0Haoa/FxWnKp
zsynDOEcTuFjtQ25H3+ejrlU2rjEaLt2X62GrllwCs00jZROZH5U2RLUScwVDpgK
kWjP8FDbYT4cNvOFRfQB6hDwRvVCz+YCTWEJ08sfvlPT0djqrGHIs3XcnMUQYP0n
k69N+11BNZDsUnhJtYOVXc7fZjjK+xUM3IQgiwhiOkJyUx4gsSpr/4H9pIJRoTdo
qJ/nQEClZgclIL8Bh+vvhrXPnRoYrqqox+avgXBYY76QA59h9IG78c4vPCR9BxM/
a/Ekrq+ubRVqCs0DrLyQ+jJsYhQLCfScwkXqLicVj/8o6S+7DRZG5fr8RYbTNWkp
kHWMhXUZtiJ0oBkD4aP6/+sFRjAPkGJTcDfYSxqwkj0Ht8RtOBptSvMl/G55plzq
RGMOPlS6EpwrBPCtaF7WIpdQ7xuSdyNCapV8QappQq+Xn5yX2zXSNaSelZPKEUsI
WuTfrpju61xGHKbfonzb5ZYlULoqFdAnEnIVKgnBOVJJeeDu17uQTSMPYVvhfpv+
+BtGTPhMX5uDsZWuBkMSx4Q9OD+SsqOYBdrWccUFvJxPNCuzyWGo/YqTW98OzUeQ
2F8Sy9L/SiLLos4iFIELwe9pQDfoqsXaYw8sBnTE+kJICiaZ0W44l1V23TC9XA3s
5YsKJqS6Ooh33NytVWD4qfo3VnStYOsudNlQqg/l2cGR0q+mvKPl0s+UnWCT1wFu
jjEsafaXeXCHRG0E2i5eW7Q6VpKRq1ZnIzurRMwDfF0F3yzPib820vi2f/DOrFWG
5gIya98GRV5DRjmW/thJ2mulXsrqqYXAwN9i5pAy4lK0gQhT0jm1qIKrsmU/GoJM
bbI4hLWfP7SgdTCrOkGg6YBo19ENNP5x3jiIfOvRPax6e7Nog9ngkcN3VbetQvcE
w/cQvsBy9uot3jA+HX5Deg8hwRZFi05hjoxUjHdL8/AWFpfL2klnSl1ryT7l64P1
MtlPkxWjHeWwyo75i16Wpde1X8QUsNjWe/a1o62Q4jBLPqE+7E69aIewv7dsQkzZ
ixCGFojfdxPHbelu53ZhnluN/u8EQ3l96yTJLq7JUfvGIoevqNO2mETK1xjCMonF
YpxExltFFrmvuknUiBD5VoNB31nP1OmVYK6FzCq1SqvRloHnvdk9Wl5qMw4clhTA
oBLl/fLCBsb5P0IOL5j6ErHbl1APm+QcFp0HXjtbQ93sSmgsg+7huDgiNgIFoJ1H
CUPDyFZfcW/6irVu7wjtkwm3wBICjCtVcybAjjOxS6OkZuYBdwF1Ogm/bWn2s44r
8JUEgx3GftEfEFDNbzs9S0ijYp4LpUPs122rUycY1XV4sVeP1x3EI54XR3OZVERi
ExGmDn9Jl+JitZ9LHDr9mIthvVi05OD1QQIQdYDVD7GourdulpoWI5SxCB2SzEFw
QcH/ENhwK75EeywAqp6J3QyCpqqbS9VkhinK77ufUy+srzyw1ccmPVs38zL7cPv4
w69HyV+VXm7xHtWba0DptnYFweDQaYJsylFuSJDq+T17t4PGW+8tQBgB469arSDQ
d2eP44bUEUTXL68oYsPANSkmFK5m8MjXD2vTPXWcq0YuZmFdpYlVze0cJXACxOjp
aVxFtertVVCnUUFWFOT/DBRn7zEBtFRFt0WEIbpn8VjTzWVcLeUnAnpDoE3LxbZY
6UFWYnOF+kjP+RLjzjOrKkNHCgDDny8GzV0MIdljs+ABsH5O5dtlrLCzq8EcjsPU
SOt4Ai8UB4V0wAEMKF+JVaaswmZkScVwTAUQweRtHsh4DXrEAoNiGdkFobH11cCb
D9ioHe96hkAk00pxRnuW7llrBezLcas7qwPERWOWhZ+GgZERc8xb12eAtqkjVexN
Agyp8tIo6LiWb3tugN1RMOHl6/c8X1avcAH5Yv4pW2/XHKhX9oSM3cAXIfu76NOn
0jaEU9ZIcUG0nF2lMEwYDF2nUdgMF8SY+7jui7ezuQTwqItGhXcsgzdPAs+gb5wv
NeQ7NxhrHey5REORMyD4DKkan71S6nWDGDPMIJiAGtKbbbSNMbt2egbD7NCgonhK
OCo7frtjOB/0vcqJBJF+e7MvHE1kNE6mXWOzuoP48LQsr/6pBUavd2HT2AeyEuIt
D9E5j7/MCAVc4kvKJgRrX1l0kyEqNfv0kgbTc7srfLzka8V6w+aggOgwROrVG/j2
OhSsf756KyN9FmmuWar6ZA+xsD3R1H1jopnFThyDc+/IsNO9FaqO3i2kZQMyZxBQ
yIG3Ou5VHwdFvw8q7Sc62sXgkqaDnOtY5Y6W8FHwDX6pf317NcE0zjhMBluHfJk7
/N1s9654e5xgm2cFKpI3Zlvl19Nn5AHJvGk8Q3qmAaZfTEk5ULrHr9iJqhbGtV3w
AohOMKnxC6qb7BKev3+xP+4ZsQGhYFIKWnF/FA88cWgV7TiS8TqPZIELjgdOygGU
DvKkXYtw4jTWDRzw/IDadV4VKMRdV2/YtKL+px3DzH7y/QF38etBcH26HY6uqjJj
JKXt+OiMl7WVWpWUxsMWUfxSrsFGv64sIxK+b+/G0jS/ES0MdN0madJW7xlfPzGw
X5BOTG2D4dgpku3tXJvVklaqcKdYXEkODW0Bg7JelJGlN+0b1GbJBg9p0+S8CTs7
/YfP7TjkTn86f3EeYvEURf4m6YdjilcKT8CSksX5WQY5XNTC2ZaRrSuDZDLAXb7C
6c9QDurf5MTpIg3bsY3ZvpSe17VGuFLtLCx6/1Nr6ywd5qT4KJGhVSbioNsSlFdM
ZPYySNPru+8AhRKVr60H71SngYuRwC3i8wfC3B3dISQBj9T0MOYkj++sTUUiHsrE
ZoAzXj36AF7sdYt8HBP7Jn34ypzbqVitArZA28s7Zckafa5Ytjpb3UYUh4fstnhw
TC/WRkY5wqXDIoeQDQb7iIK4VNlKcz5kvqqKKGDrCWyF8lanAsJw/cm7xTjmoE01
dUj4E9Vqo7PhNDnBKLOTDMCAvKWV3VWo4oPfiI18KE31gh2PrgSY9KoHZ/666o3y
vMVywASRPaSNOxkbsE8gk0bVG2EYJe7nq5YG9PChZk/7x1H/jmrx9ud+HcjrFbH0
wqNF2USrt1mS7JzF4lNVR5xXbbeXuWQFL+jHpwFe66HfNJntDpF5PV1OFcPF+IhL
dj0VLlAAH4eqZRkY83nBPYVeDkBxbh23TYHVOGYR0rvBepp5ekwldPPDlcrx2L6V
vfLPXPQVDyThTtKxETprxQ4bo+0/t005Tz0mYXGP2cH74WtzT7HBtTBjLv7906YC
rAzoos27GF37VKdSQwTSPyAyUjkYmeK4gnAte3jgLu8SYST9GkhX5EM35XJm72ui
GVOGkDIsv7dlzC/nIFejaey7OOPtHJdAxkHgyB9kPAu19FqQRpFk2uqSEk+/uDec
SUERyIeoo8IZBaGHeaDIA+ifBwRxomh0PFYGectyGTevsV2rhV8EDXHEC2P+ic1l
Ej/AYp0AtbID7K2p03nTbb5VH3RdgOWxdaOAMEEo2qlkVuAHhEJiigasUF2kStmF
RjoCL+YzHWobutb4DDDrsuopxIEbEAFOqSw0ECteD5FQgxKWPLt2gUCzTQWBiD4K
iVQUKTaevrasaVkLpxq5mUYzAa+SlaXedLHj0taMNNEFc0Tt0BS5ovk69K+O1BRB
RtKKjyiZILRfFZbM/2OiXY/MBGgS3/NrvcX54OHvhUXYwbrxHPuPoV0/oms4w/Ne
eDkumabJ9OJFEVzOOkZY9jFJ2NBKXMnVsosETDyJ5/MxroEwjnm5/8JKPhY+RNoj
pcGuwg1a/k77ObhnvKEdoIiAgnjUHu4PSx2bmJ3ly0R8N9h2FBEJ9XO9HCo4t5BX
6AmvwB7r8NaW3SUgH7HyuXsdjRKkp5TRgq5MIEhSNXrAtMarU1YQeXRScj+YX6m+
b+KTVfcgyS9viMmv6re9L7YIH/z155dOYnUyMG3O8AOweHYHGWlbCaWEVx+HLmdo
s2Pi9DipypI9FM5OBbT0bkTirePjjyAEU4ZrN/2RfN7a6YfWzt28GAuneFc8B9Ma
t8cURxrFtA1ui/jw8TaOWYFRPscaH1HpZZb4klXSmhSLLyg689ECbqf8Y3jrYBuF
8QySQM+C0Ak7J7HdeD+nDhGBdhskY1SYEWzSTCF9X6P1RvMjzb9LdY5YTDZubSOA
4AVVmb8VTw+J+JFhF5J1V9wOk79Pu+GcROa1j63H5KqjMNHtySV7g2C+Vr+eCJac
acwPqeA30LJx9kXRkRPuGqsi9JevNSubexdcvLfzNpIcB07lgXyo85ruSS+wyfF7
nZwtI4wBSEko6GA7DuY4XtPrShiAigZVVYtgkvC5r0AXqQhMGILaiomMjQYGySje
hgAxKd/vG+Ak4XRWqGahR+IS0ogbhcMnspkAD3StMqqacVc0YUY7yOz/JYRNX59O
RvQO3wL1EmlvBzIwkxMl/C75L+HoTtAovMl2bs3xingnvYgQ+m7IDR+F7cAVxC8U
4iKTK8uT9mn32e56BrzZiHkpOcQeG12StztduOt2xQcfUcMufPBRLRBLPGtZLOny
RY2gWnqXUNScHpZUCxJPfNrA6yI0LnRYMMV0iS7AI28g3ymD8yeUYHeh92v7PdNX
B5dZOVpujDMd6HsLBVuzI6C4hXrk1uTzH2buISfhXu17w8PjkFP8fQ4MmMTEeRM/
v0sr/5DGariDZkm83fixxz/aa0SB2UWoAB8kgisucToDYXx4lQ7qwWuttfg+tgpw
e+FZeXv9OPLgkcAxAy0Dx1uq+24CcqcnMNbpvK7lga/NH2XKXub10+gX9myQNidj
mrzd1KUkdAg2k6mfOTj/TKFFECHIG7pkBd/pKG0UXryT/8a685tnasuAwamDBGqo
D2POEWzNkEosHFvt644ukqbiLLSFB4NkqMEgDYpQXyJO8Gn2yfqef0j7yvCbA/gc
a6BSuaxR/Yq6TBEHjRU8+vjaBMzTLgZXQA1hp7W6KAx5UHeTRQ0lP0giZJEVz9hr
6N3ne8SqJBChh+qmT8XZYgf/oLfiBg+QBMRP+ab4IrvEDvh8jSsgRiwNjBdTECCC
zus7ci0BW8izfBvW4/YI1JwFUF5meMx/tBSAxJ39DnH139hBfzx3OzPsvaK8Isnt
a+ucfWqDpRhsH6EHdghizSGYvyB76PTnHSXwv8jllsYoyDR2GlNPiQBWqS7Mi0dQ
0dHgsSR621QSnKr1Uh4SKh0slqjEmZwjlGhJQT4tWH6K0ztp3/aN1oNauV5GSVmO
YNwVymZf4Iyx3mifku9XE1Qdt55oVKF8mDzDB7oH7vNHayxtAy8QM0I1xzfqI5uZ
FYzG6FmcfTvsTVZuSMNHVPWqlcb5krjXSK4LC7wUeCMrX0/vlnU5c2jl8bvqe0g1
4tJvUMRV67U1iYu1DMAcgFK/qOQAiNsrwaiqWYNwu2Q964s+pDUrgIqNICkSeCK2
F6Fv83c0lsjT67vM29xXQ+yzst4nSFrojFTx8JFI1XK4EhoYjmquWHPv4egOthNv
uBNlMQPHOtzEerynJrrBGOmVUcyLQUruniqgYlNuimcclqIIsxO9G+8EobY/GsVY
ChzMUgsPjbokUNqY2hTZ3fqK1d+JBmOlWFq9i1PI9+r6s9n91c0haYnCdHrNIdhk
GIWI5YYe/ZBFuTC3ocJmeWcurBvkTCN4edQh9sXOGOwdSUpivKN71IcNpWRGUiCn
AUv4GOwcsTfBSBO6kahlSp7FehuuEvRs6qb5tZZHLU1BFGpCkm9Jzufufvp9+T9h
aHIBJs1mdU4cr/Dkp6NiMmhqWoCzwahi2/8UoEIWpEIsYR5pEw9uTv80azKdGAac
PKnctZeT7AIMLz2sFxtjc23qkoXRns6oXqDdK0CVq+cPzkoX3D4TMsfHXC5o2LHn
mO5FDp7Nv1ZH7qDra7VYRuZFwSnNQCRVZsVSGz7E1GOHLuuhY/YtolcXeyXDy1MV
MEHn1pRqDUOlLQxUNPAyD4d9dCd2orsEfhUb366KaiKsWwMtIJRjU455peA4OEod
3MRvX6iWpJ8QfJ/xYu+iLtZa13pXrXV9RX4mB4rhZitc85T3yFLBpJY3/yW7q89A
53U0xUqj5Scykw0q6NUCeME6Y4aMRLj4TTWeG/+Svb0bPLuhZNswQePgMQfz40Ef
qj3ss2X6R69TR35R1eSN3WbHvBubbrBDKJcifGeGY7xu6Ldvwkg+hWQS3Rtv0vFS
V0AvST1WkBJBRk2Gtgynk5MaLsMv1UAZAXYJDnEIXaql3060shoR7/MQZTBh6xnD
fCYZXA5fJLjv1sCGhScUdd/xmBfoCRidraX1QApAyT2alq43CAgJr719PaaJ8Upa
64G62LkLFuO+tp0uM0pjkchhDdQUTZrzyhMoIzHMhvHu1yrM7gvp2zMYoJH9k8oc
9SYlGE40Q8oH0r3HD8lTMbPENapKk5vyMcHRiFgwGY8HBGS3sLSDms4/0o5QJq42
NmU6julxu/s9mIIETe+uxSJl9ehSAEFfjqOy1GXVcxCu3TmNLt5ZYi65e+J6PJiY
/rRHH9ErF6U3/BPervgW8ez4pZ+mFWAl9F1v0Jk/EldLKydtOm1p7Etgzfc6gITv
14IGMczzpW79DkcPxBOAq2artEaMKfB5sEQFE/dz7/O0D0nhZVYT1xipWQDbQ48l
Zptw7ites1qXYiob/iXIelepNXBgN9rvATgMBD4iabroxCKt9KklecuQrNbJz6I4
K0W+RQ0owucjcTv43MEvWE9PeY5kUUiTJDK1BkjWS7AO4eWiwKYrcfB7d5kidknL
kmy0qhxiWXE0H0GATQ2YzIFr+9wQKEUO8Ww3goMbwvrZu2AyQtHlY/Wx2E2qW/Tu
uN3Hu8984xmFUJkA43Jw4JVZo5P2gTtLtxY8TFbsvSdQ5C1JhuFLVWxG4Rd2cHvE
0Py/Tm9A/P67cDyd1SuwNr2g/dJJIU8vep2NMsyweNLVJrpLDTvN7AFW2dM7Sou/
kYCxrzkAD+5Iq2LYDnumU3TqqSXFmAMWDObWa4TgYq8DKdMD5DuVsOlq5Xbc2U8W
mpwOHmk7gPHjpWaj3FKOkbiuswdIMCOpnMDtRYl64D5BfMnEj31ZZIURNWEO12nd
QPkwlwHbAy+FTdPSEjCdp+iOlVUks24DCTyBh0fx+hiMK80TCa03bQoBUOyl5XXu
hPTOaQYH8rCof95FlPvQgsjtHiIweQh/p5JhCV38EJvdXaDTlQ+n6QN9v457C+4m
j5GQ3uIUJLyNrUxjaIZq+q/ne/Bse/bL9gk65nWpZ4Y0/aCLKho/Ky84L+HVRcEr
lRqUyU7gbMxClTkk4hxHYEjYXVCwnmApZ3ylHGo1UiVDHjcDh4OPA2eEnE2sKV5/
EaaW0V7ac0wGSAXn9jry7RK4pwSfJyALlcym/kIxfS7bowGzyVhKM85H7b+yys9n
/pSu6sIfxNUu+UA0E06nWMS53ttH/NvH8oC4ISb+XAd1A0oYAbbezZlXKusE9Zwk
TKLNFxZKoiomxgkhlZTyCQOWcrrE23illPxmA9ymhZm6qv2o4JGFw6TBsHdQBOZf
Ubrm1w5gXBZlXJJDgwNqcV4JCNHLcqFJz2TqbNRwxpEuQe5iy7OP15KMpidTmhm1
UGJ+m1Veqq05/TC3Qbs/CqzaeHDPNiXjNvuKaY/Oi51MUtgniXjj40Bn8Sgxobnj
Y8T0fUV4DRHxOUYn70cWLILsIEa6bRkvUdu/HY5pNBQSu/HMPSaeacNavB4sDLvy
2AKgyKnXAX4ZddCHBHuHZlqo0CDVmJsNqFk+apDx2IxxDv4fn7G5UqcYoQMcp7Bx
7QJer7gz5A6QWSGIdHxWbZhccPJ6j4490JwtjWbWlIvDIQ2yP00S8IC1JcGktaGu
wvltERSRQN16BBHHfeEH8Wr7Cic6PhvAN681bcOodHd1XTRqWNwjSNUf6FwVWeFT
Opz0cFiEGTE6J5xAQLRTWR13CPgqaOfjFqnAlVs8kI9TAO6TSSiq/dHvaRnrma1g
i5/6I1+sqJJIxiDygk6E55X7i9731kjUMLwsFSVt22hybXk4xQP9LDJBLZ2Qktyz
XrwIMeNjZaoAO5Gr4DQLH24B0d5c4ejIER3zp3LwYtby9X0j9moY/c00Y8bC50ou
Vy+CDnmXjRSS5lAgcLREYnm90Cvyt/wyR80XV0/NoTGPtFdozkTEze200uEKax1J
q3VuGH0T+r4tw4ObfrwJsro+1GqPA8c9ubrWzNipJhwPRv83hqo8lzvSZdjznFoc
I6uUNpHSFt1XHYFNpTq5Kh5QhbTynLNQgyo+aDo6WYhv4FW7PNnN6cD/4lZjpr4s
+sTtu5T+e9Y0YjStyqNSpxzI/QezZZbTsZmG1rD2H0aYxBqGyj8vlJKWaCvu3jKB
gcw6/ZT4R69Q2b/4xGGAZSZE5z3xj09TBQvBegcnh+3gQYtQbl2phtWqb09lu50P
NwEJCEj2sKW0TGfLmpdaWgGT/cCKacbCwCGKLHfKVjs3reiJxQiVK2DrQ0DLMIvB
iLfNy5sm2z+sq9/f54D1/1xZITXbJjuuOLqUWHT/W31mIdSwxZK3E0yMMnwhzVte
E80zKlHX7ogxTrIT/mOyXUWIpmUzvfdu3A5jaKpcC9/9P3zgp95QCiu8enosnHFF
RHtkWzQRkFIllH7ZYv+xHWjGrwWSvliRlhdvGESfCExWpZRFVXovRXy9KqG+rm61
Y4VY7htIw62dZ03tnHUkS9roY/aE9ZS50B14kInpizizPKEeQ8MBLp2OCE7NIQxG
Kxw2m3Q44X8W4bwD0HE2vfuzw3+icYFKZg7iJmHVAvkCORsGKNB3yywrvlWoZEY/
N7I2lj21paih9YQG6syQivVMpQ2QJVNOpiLcEI7N54JwE73O9lExTm2x1eA9MMyy
Y4a/L+DyxVhbpybL9vI+u7B+p8R8EHlI4u4nBnkhp4TeZ+LPds+eSP5uECIP9CvS
bAf23IpvDExTLdskwTNHvaUUCwvcaxUgd4ECq/GUAzN/F9zMiNXcFTfOBa+dglDT
w/TUS7Dnf36SyRGD9v2+2ziTn98U0uEOGve5CVXeHqVDMWw+5tlgqNxFKMxBfHG5
DRxMF8mtrdOuZx0lsGHI6MKSs/PAZI7YzE4Zi2F58GDAfi/RD9GjrqWankgTpLsf
8bAYDOpoCb1RSDQrviYsHcgxD/T7Ze05aZX+OFEfrA8PHoFdXlquQ5tOoakFlgqu
7Y6DMQwnlyIvwyAmkhU72yaY3bg38aPWQBT+35qe+X+SIx3qcyHc5atV1Zu+hgnn
Z3IqTkDNxoOqtMnnO0eYbn86rU5oEHBT7BjMjxdZxyvph0+sHJsoC5QatTdaZvEY
liS0TmRL/rDfS5W+QWputlgXGDuO2Znlj056NhpdpW+7hOM3VDUobk4rLr1T9kbW
tT5U7wOSgwFeel+8Fgr/ZtkKAVUjmyXTDrwkciIajX58RUQifh91YMWm8VXK3GGu
2OeWSj7fxjkVd1Hmt+xjAAk9wwhWndYQxMnsHKYRnmPxL2Nw5VAb9rn+opyEAUZr
IqKeDW4cI8adRryIk95quJpk9C9c4RpWyJ60PhlAhqTyo6qc5kLP8TjgVM0KHX6P
JPhWqUUNmcpxLC+xbg0BaaG2NavUqYjYlppY6wJGPM3Lu1WbobeqfcwHQgU1lEsw
3W/c8EqghyZqceRipuuhexF8rXzc7fQGCQz29kCJkO/2tYsATrviIjkgnyY23ib2
gMzCBOJEa02iexB0Y4ZL8azP2ywCDavSB6eLPa8A4QjV2nrYZ505k6F/OLkrmym1
UksTorMsfo/PifvGkt00TKUrLjtUtRRj4iFNG5SiKr2TS5+FyT7JbPeRwGTinB6i
lrl0lijBuRqc27LcfMztgavEHWdYsThHu6HGpvEBwOLjjFl4m+dhIA4vRCKsxmX0
H3hZMvyCWSrxi8fOJfXWOb4PtG5slE7YirJhU8O/PQOljA5Axu7GXMY5ASlLQwUr
OZWXDldbd886/pN/938zU6zzewbL6t9IHZfAHuaMal3bW4+yrmHI7oJdjxQEzewl
+yNDvBZ7Wg35ZJroNehEpIH8OHzHT4MEe+OYy57UdOwyTIX0cO3BYcNLD+hVy4xM
NnlJ76soWOwCn/VMBO1+8SM0gc/mIYuM0c5ImKXSlQd+lS0hi3l3TjsjdNhH/YP3
6krolUKWBEvH/K1peh0MEgPsdTvKbiK4QrXJ6FsI3pr8ipaFRs0U2yYdUQYSHzT9
dh39g3I870lHEwYvg8u/RCuKpgzTb25jcESRZaB54HldCfm3UKDm5zMyv4MW1hi4
hc39eVLWoUI/szL3WMl7RX+oooibi7qItAAL4JR7gyvbS3Z5DU5+63LN+wGIOmlq
ZT2iptfE3XYhmeLdgCF1JqgZsZtFN+rfrANQDEJhzle8yDCoqqLlPgZTiOqM/DDu
cCE3fOrdSN1ped9lNl84CbLkyQahvioVFt8XXW94sLP7bcLLtSpRB5LZdQtzME97
yWA+800IYqmlONxE953iAqs2rrIbamfulQOxluRjDQOLLEw24aoIhI8OF3KcLi9y
T20WyAyOawSmy5Rhwl35Mp6ouBV4geX21dPY2z6KR1PagcF0dmFqxVmbwQNeGRxG
djildsTmqKVU2OyJ6qQeCvbfufc79YLCiJIKPpPlcvlNtcMKMNvtOdjGqsoMjm78
bIFZ4XuM8fCgoxH/8uVyzPHqjvQFFUIo2ayg8qoWwWV9/r7lGnTAPSUB7FFiFlWi
9Zkr1wDgX4pCs0EZ6NMhpZTCUHloxDledilyaF+n08Pcb3qZaxbLx/1HLgK+hezI
Ul15vDQC6guhOcXC99z9YHldoaaRqPUhYSos33sQQ4X0L7J+lzV9UE5QPU2lfECb
5H8ZhRK9yzGjidLee6FufXgVsrGwj8YxdQhPWf69939MPcJE6x0a+ejiodolKmtc
sl75CRg/9WkqMREEF6Zpx5HcyK55aA3EKZEHEdMCAYfkuSBCVMSlikaIHyw7mkil
uCZxpwU8fvqemVgcBRElWiId/jxOldj+gaqLmazlR0Mu/oSFkpyYWLl9fMZtcRdL
emJ9iRb8bzd4/zC0+cwoNuhfFF+lhwXZuxLS1idasLo9ms3ZP/DeUh+Nyk1+IEo5
UvYn0i/GxG+EQ/gco96v5d0lFwfRP6NSLBnZwaTcB/lI0bIATfe86vRIZH7kYMg8
ZBg5wIBzkGVuzP3p3T6H5d0DfSyhdl3UJEQhovM5a2QubXQkGbnz0hBiKqw+gX/x
pSrXaQNILZY+biAXKZDvcRIRvCX3Io3xKx3/nHiRoFHBB2Rv53a+8b9RRsvyK1Us
Vuq0a8IgLnTnLwzixcIOoHCwlmWrk2zcrY68OZtveSdewGtXbwAfrRkfJdcKch3I
h8PY67AhZGe6WQczRjmkesh36h1rPWRG/TXYD4xPF6NYSiTURQ3QSlZkzKgzu426
y6mTNkIShvcFbXnKOGVGRNg9Ph5AFQa4O8x/ld1enB6r+wsAR46eGEMYfmak60il
OxzP2Wmn4r5L7gax79ufIfEWH1sDKh6t5AiiL3ajQa5wV+eSE9AbRlyc1h1eGebr
pUzPls5teHrSADnDLVtwzjX067s7DytuDBa/CHDWNl2h6X+nhrvJKBsyLiz7iSd0
N3oYF2i+kqGC1taoXEB171KnfI+GzCV1OswCyFLvPHDphYHQ77/965J8QIEW2oO0
VkeIAsSBI31f4xjUlzmo00f2swkAQ4s6SsEtXCfiaDawh/8H78f/0MZ1BeOejbUD
DZJou+ezao0ha2ADPj11o+wGcPye8wETWIf+VvMjHRBfmoypvcEgDSgtXsoz8C+2
teJ7LJfDhqRicSHNb4M1htgAnsnbtPO809TjWpA1Gq3Q73cMoyXf5ULGJJEi4ifb
egm7cTo1N6LJZQUapDlVAaAggW4e8qKovleO54A2uKUZ3n/YouzSLFsKML0t5hma
Hh7vpb1zo0qPgvLHtO1UIrHRrkjP9rBsl2zor3GtCfvE2MW91RY+MVUctT/t32Q2
Binh0Mce4DEg1BGJRmNZixgjeBjFWet76IanfB+yIzgFo8zozhrZ1t2V7MGGwuP8
ep5JxlW5++3cC7ht/rKW1KeyFSACH4Q2SDzAfbS9BCXD29Yq9Wt75ntCLqdAQmgh
rt73bAV3uuITa5cJyKi7Fw8ZUJM72qeXW799Yaf05jVjqYpRbaxi+ObyAjfpiT/+
8yhI2nMuLor/jpIpRaosX5oytsVB2BdUmfGjy38sWqE4VySplPIoQZcpArXgFSmh
/fYSYwzu5UPwVmfBPMVi7FhgqN7gZILT0QGUvYVav8w3Q5vaL1aPlEmREoEDXS90
fppHegnSx9DeeVH0gaMb26dkkRqj88qdPAJBe66EliYFTD8lscJYpuVxGyDNxsfd
f6u8Loe0kPtaVoXCPZjiILy0CmFHVPYmG5kSuWiseuDIOmZHCQmp2BThsTyDdUqZ
0pYJP7ecii5h8h7kaMOP3vOSk5omiPpVI5CNH+bhKGrSjhlCk2cqB+yYLeghUpWt
tDsxHrtyZrwWZHxOD95LSUnzM7wiMLGiE46KWA7m7KTqYk36w8R0238RzNGiWyv+
dPzA4mvc/POTeZAE0FZvdxJ1qA3HKoAq2lObeWb9pjT/wtLDi5R4R0u53TpyUHnb
/TbKHw4/pLy+d54PYhq9IBHyZfJkQ4ztC9DxufkaJfxmQTjMkCe+GQdW7lloFvgR
M8BOnUZq6phuyRt9upWHC5TgpLNqVQy2NNI4k+Vk+uG+CgRWstRVZdxBh08A6tzc
9uTczFxqkf7a+wVP5q5JxWOrzjY/s5Fjm9cxNxoHYPxyw2gAPnqgQTlzZiFAsIXE
c/jRoOnVvGUw5avL4cSL6/3qvkqykLaNVXN+lWHjYA+ISSvpw7mMK+KGPf7unIpE
8sGROkRI6pfQ03MUjmD6x0JnhrPH5d1njnnolxZq5TjwHyAuK4pEMc9XwHyBJz/S
7g4MlXigvYxABcgD2uS9DzjH4SFws4oNdb295UcKCdiIeSPUeriFwLrys//bOiud
stg4ZeSLObS2phccWlTImNdIYoUqP2j/kpfZBxHK+/uaWf6UPGQOdVLEHCZ//Gt6
PoECahfOUv3+3RNM55oPBVKjoHMGdnbbiKEU66rZzxCVzWZWe5QOhl9+ox3pNiGa
xh+a/DZkdi/v6jlbTjDCAJLF+FLkqwOZ+dSUdYShqlHcNC//0LZ3KlJK3t3kigIR
CiOb9M369o/gabVtvNoOAJ0HF5ppE/KiyTNnVggilDbrrR2DA00UdTfuYxFOw5nr
vio4b+erMorFCPTqgSmcCHCI/f8Xz2zZ9MHK/CwauFD6S/oJyFm6Kqb/+IzZFDl1
06eOrIWLdueSWMV3ymCyJHjRJQwc+pLjR+W8O5qly7p+a7msxg3T3lkmM6VJCr5J
84H++D8es9s+q5Y4/dtrBbEhHA7wbm3rI7kLCThjDgQiKCt6jOR7q0fSlhPQbOq6
5gHKf4bPJ4jA2M4SFaSgIa01OjuYslFD3b/CVbUmdkLT3xsYKSDbbJIXuYRvBmCL
k/7A96ibpwaFHvmq0Ws9lo1f4HnRDEH0/nqGL3CCe5ZxHo1iIOuSqPRkmLsV64qW
OID4lk2i/UUKhF9fzlbMfPKA4afm1p+UGvKsuzNSjRIGT+0XyF4vY1xI/jQ8toxO
P9rGViQolbPLGS/VFBN19UbyZfuW7GxTcdDwY8XYypxE4y/A4flVI8/0FJy8tj6Y
5G3yd2NytAfj3OkOfzt7MrWPxYXR1h8ywIinyxbHqNMQMtZO36zV7e7U9hr0hifI
VJtoDN6QL4dgIeUmWLjpKKdwjfgl9V54J8f3Ix35iZcE/5slVQx8sDOizb14L37C
EVTTyzJ3A9TQuFHDqqrA3h/LskRMSuOqpotx5sgxa2xLKhkeMp2K0/gWFdspxxtk
2pcCQ/YckX9zfVkyARBv7ifgBGA48210XbcwGQlUOs3TeIXo5kuyEjqIracMw6sz
HaE1hDaPAdv7b6Fh+lG9V4k558MRjvgTo4WTVwuedaohZ5On9POCD+i4kJHNpeo2
P0mQdrCaid/BMf8ZzLev/XtZxV8PF7eTaSyr2fICBTrbekJcLfm3EghcKaLQmSau
XZvE23tOjOeJCBu+1kcgnf7TXFltPcCEX44n0GbLyL9wXywNKAVQ6nTmaa0+l3ph
iNoCOnbERjRT6o8sqJXk3WD+tVP7+ZiFeUkwu1YzOMaWxDw6w/6bdQ6maAtG3O1C
ZHzqawniDo0L5XetcBBc6n+8npFb3GwP8VzLCzadnu2+Ng1MvxBH0EKS4jvV3Vew
BMBvh2niAK6Ky0DSRtha6SkCcGjXdveRwqjaYwZ4jb+jNjgxgCHCkNEAOCAeM5yy
5f8bDvtod58j99l+pODyo2gZCBaaOe2eT1Z7vcp3YuT9ox+WK0hL1kz4wa2z3ZQ/
UVl0zRJx81FHm5V9uAwCug6hHN4n9EG6RnPko3ecns0lguFtHLGLNmqGuKkxhJuM
J+RKtQ/XevXMNX87xPtT1pUgoarvVAx1sktrf3IKRoIerVlGu+UJHXf4bnHNqS/Y
UtMXmCIGrq5/pZN3dnyReJD5mI/lOL0vPtz30lRX2tS9X5PEeoiIi6huImrsnfiW
UzBmnj88b07BDtQkoPRGfPbOr9basvLjDAyMhIHlEn0/A0omSykEW+mCGgpisgPY
49J9t1R0QrSq+BDktWd8Wp4kZlOorsc9CBPY9GjFeLztCdgHffg8mfuQuzZX6RHd
czVOWwiq4a+yednp0Ge9Ib2VDK7G72IlaAIMoHbzYb6xw0ezB75FiMKURtcvgGV/
/SrwcMoKGX2Xh/ArQ7kv1lqdob/QoiieHYE/FembPMY4ff/SLdlybFIELZCxClPL
VBRhRvm8KSEkU7iYsVh/nmEZGUNi/IUJonixZ8RY9S4Sa+cjFOplN0KfKZ69juAZ
18Yaoo+V/ApzJyrlNYhOhIfqbDiMmK6Y5k8cTG4XadFuIGRX1/kUQ6WkUrXLiPMw
QCcoaIOoOmveHIy+1LJFtkhNHTilOg/Eobn2NUsCleY4dfmAJMXR5JniFb4F38IP
rQQLhQWdmeS8ukaLThR9CNDcmT/qArTOf6ACNX0KI7nUjHJd7me2N/YtWGpWNLQX
MeXA5RM001giLCkP7WL2enZqH1mPAfSiMo8f6OEnFw6DEngRNelFRc/JjTH5Q4pe
gAoc2Euz6rgjDfY7xu38js4BNqujbjqrw/+pZSjw8DWc65vVUiegshb6rmdMHZqR
QPqu6tnTKbfhkDgiRF8frsJDikbFosl0z8RJ9NNE3qpGjI2aw9QFDGVLe597duDS
Bu3IMoFPv115jXhSfzOI2k7/ZrPgYiPonx4aRKRpvl27+b0iDM7AqGVzN9AWzYrL
bXSFNPWKjy9tW/Lmf43No7x15OZSnLMieFXXSBDA6hOkc45MMQLIR0ipQJx69cQy
YWkokc2Fj1MZx3MFvmI9LBu7YypTXdQbh14OAS0ckx07cDYCfDTUF1z7qv3otk64
ugKlAvW6OQ82higQOJMph9ou7D3Xz+riPZWW9zW80nLaBerByTV+Hx6/fNCV1pcp
3/72PF+bikowFrYsQIq8gVcbmVROXo+qFjqwWaPI9A20YyNVROM6xKe0n5m7+u8l
tUfjPp+KC72WuqHUQVOwVrfAEfB7xAIYgMEp1WWvZIWfdd1sRbRIlfQ6wEYSLyIr
WZQGElIxDJMOFjhcIgn/2jSuGX+aX6OeAFswlJzhClbNDCmG5BHeYKY6K3e0DJDZ
Im2CzL8G5lOuVI8d8HA9I1exso0Hr4AKn8OaVQuYQ3Aowv7Sdx4KlygVwDiB6jCR
Xh76UEHKJ3ZyImDpi6IasG8ZIg6d6OrObH87HDYjKBJp5mikoKI2QGNuXsa8ZxNn
zfAD35hOOc+2KVkjwsEfx2af0Nj8v+3HzcJsWlEnFpRVpAXDP+CyGH9GbJdVWOdd
bwWTW8NO884fdraGxAexNhADqmbqqYy0gtZN1QY+x0xBFHszaYwP8UHiAkYkvOv5
URggKn4wDImIcKTQ8n4+VBazfgAe5TEK6jWD8GQvXUvE0d25BiynMxUfFMZ9ebL3
3rlAPFtVfuRKhlU0cWj3S9k29tDI3GsUzuZns8HIdO2QyVmqqSttbkORH3JppV6J
kUhBCKvYZ7aoVmuSRjtth9a3udZd/nNWhToU1PuQ8fQuD5WrExhJ2tziHKXDAR4h
bEEuCuRk3NKkdkMTRgeTxSX1JlPA1PqxQIdbfGj8LMdSYIV5+tc/VL2bQ+uef4Yi
BcoTo2DD1e21QSIXP+8Tk0VqckVkT4YUtW5LyAyQIu9i1MI1T4CA6fkbYRdY+2W4
YfHzLM8vGB5JkYItg5sxfpdGMLJgEDHFOl2PInNvvDeZAZIQnJAfmElgmNt15nMN
2FmNRTUOoViMmNes0sMeTXvwgWqmfywflUnoHuSPjPIRJk7UabwqVqFyGq9JEoLs
HOEbCWBFpgVWD+Hf2tpiz9Msdy7BtGJGO5jGRAJvfjIvJxUgrAZdE1TQcusa5+ek
VbmxjqyZbMtUwk2EZSKF871TN0UViuz6GekWwpLGji+f0qKKWsRuxLHPbl6LIaOU
l4kI7C76avgyuD78YtId6f5nHcuh4f+tp/QMBOSBDmtrq3s1NrEo8GinKTUvBPA+
cVT8r3uFFAzvKysjfkWkNxGF1q5xV72HbfbTjXgWZQugrSr/cFU/U0DivjlnWlGC
c7LCREYVtmyy9vo802Chb+iwTlnd4Gkz6iT8R5Y/vh7L/oFc+PqSWvc7kOuN7aaM
ugfcBJOE9S6sQfcrPnYsmjwHhYYA4VCxpyv+oFButpybY6TA10UmKP/cGr8fz3w/
1/kfcoWDoHiJzrMZnVDgxyWVVTp28GKso4nm4EqvQ53NEx480lWQk3dw+qGHKAsy
E3jfM8MIbrHyDoRZMlW+ySW6KXaA5X1cJqJfxyfZnO+y2GdxKaZv1JeKG7tS48gT
Q6Hw5zZ2WX+N8dNFM+hg3coNnMdC9TdLyASZZQISX6UuC0hBsQuo8byKszn0hGmO
o0lgSQ3pRYcfO+Gcu7hVdkPUQiLimk2QPYFLItExn30cjuRciWFWjaH5aIMogpWd
AXzwtvKCBbDY8QPeyvyFXi2qh8Ccr3MpDojeI4UshWJrhCiIemWUxR2u8DUjQEn9
7oMfe7tyi9PTLGcNVDEDfmXXZh++Q/UppmYppFayKtitBgl5rXFgVV1ItBcGlhap
GmaismxZxelocleBELWBwk4z+liABscN/0f+3kyZFDvUcyK37dcjOu34g9D1b+C4
+aRexiB2fye/lTEfdCNm7fLbd3a5jhDOn4HUBjbcZZ7HTLwJobIUUTKsPXEcfSaI
/EvbsCmc1Uoo8fAKNR3QOcJElWNS6Ug+Md69pupDAFQUlF1xNO399u9KsJBUexnr
JXNc6pCWdGB7Sud62fkfOb5JpUElJsQoePhKJHJhFaLAgUXioCzbxtw2BVwqzVtl
Cq9A0zNcVOauFyt2Shb81YxupYPJbvlkkWYlBEY/f2SsozXzNC/F6q5lPvTFOjPw
m81OqETz/tPctQwgXqH1B15Rr2ie9gNeeLkHcDEC9y5VDm0Rtb8EkeYn8dHlG1cl
1xvKh6zvrFNcfh/AbuW8Zq3kvaUYgdQ0TUxNG8LuY6sVkTr8Q22kdNFpoBbuE4Nh
xgGgE2HwHdXa4KBTmS2oMq4mWtP2qiAGEs7GYbvtZEUr0UZpu6iRtZSp6pYa5fhF
khesonx7xCDcF9uF1+at5kd3DHXru/HCL6RO6d2UTI57+/yO2TB/adTCpAjj6xVs
mduWcDLItjCmhM1y3igtPzu+xwT9oNChRfnNGZtzCUscrY0FrWEi+UvWuMC1ZTYW
BMuWGucycj6DccjrMivd6uHUDewcNpmi3St8j/CnAfWvV6UmfOm398wME2PEUCQO
1v3lzJyyhKMQQ0epPKPSL98OO1g5N8KWgnhUpE95gnRTdwfviOTSZYNQ9kUQfXix
8aZXo/JgR8QcmX85Oz1Tn4aDiWZrc8u3T0I6KqWxQokKXB+eJLUdmwQcnkjqDJgO
8Osb4NIP0QSGigwI4+BPceyTiXQbPwz5pCa5QQDwcfSG9QgNwlatHpAw3iiNEVzr
DZDnNsvj24eSlTn+N7h+uBpOxZj5FffozIpMIVYJjHANQwYppjei21bUXWziqSYi
qqYhPvBoDDx/YUIAMln7WC2AKtnUva/XwBx9j+z2gTBMsCynL88DaONcbMgv0+bO
8j+/VWqPA7YNoADbzJVxNXjGloDWXdbmcBDbAebk/ucFA8m0qCI6FnpGT86+ZwT7
p09FN+AyNbrErNc2R8i700p3CU60b+YPbLCBw9b864JrSOGyE0wKmpJ9orVkG1Yy
ZgsihsRvqMwfOa0I3OiIrwBKeF4xQBXO/EzXuImZNajp21DERD+CrSG2PVG2HiP7
K7Dp1tZCcz22qfE+W25MS+wW2fshHgtVncLUVddZ9ZaZBBfHsE3YLKSn0ramWftj
NJfh0SKABC6VEF5spvmlp2rthruxiwmbs8U+UN6AjvqrxbNDDg1B9z8vuXrSokQP
QuhAmIPtJpMNp/JIcduyMJGP3aihjf3U8mFkxv/aZbLjmshxNSyEZQGVZRySi/7H
UNnGP3f62jhfk8cz9mXUjAB6+RTEDPyNKzHj37KPrSItJKlZriivLn+8gYGdGDWe
kuIckVqPkTbdYg/GdVL4RRkthf6/jhQKM91MoFOerPVhQVDhwQEIAo3OdQGFn4xR
JbCdQ7YkQKzXQ2J2gke9cw9YFzYxLxNh0sGX+B2U/n+AjRm87/UtiH/BS1Hu+egX
Eldfh1QErJ/Jmsf4EboBo7vohMKZo0beO0hnGs0eO3KugfFM8GED1etD5P41iKl4
FSnWJv7detCUN82zRJUDqycTY9o0qrk9M8tWwAfSio/tQZ850MlW+srFYDGWAJ6e
eDG3XID37rjnGZxlyY1bqxhTk/YMrAZsp7DftCfwBNiJed6z6WFOpJkP5IRca0h8
lEJtMTfnARQoPsiy2bF6Ny5/00ZorIQyAv2hrEROVthn/ALpw4BW5FXdXUPmcUcp
+G9ujimVhOXceVftOn0nJ9k20b2u/x7OswO+Q3XwllP3T5P6cFZfiUpwci7N0BRO
NpGnX7/nQcUuNT8UfgXIQDUgPKoXQ5s7yVaeGs/OqyX8TmMnadHmW4jniNDhF969
XaDmPCTvT65cJ3MgX4T+Mij9u1fejjdgqhHj7uoJ6j3GPGiEU6lRl9eZfwUF8NIN
mQfj3uh+xWsWDrzPUhRwkHufkw9qnZkwxCPAGW44hSyvF+BMwaX1s6bARV0CVuJ7
vBEXTPX7rJHtSHuIPUeb40BkIALYetE1fdgEjig8muAFb4I4PrX8cR6M/1amFK33
ik92TitktegdqspD+J7M2EK6i5i0F5Gx2uDdgLDJ3GRUiH/rdhlWabbD20K7R9VV
Xu0Myh9TlckyW66g+qgATqzu0wUzFmnhearOW7VsVZM7rK3lOUSOCn9EAV9SeV3r
RiFK/9A3/76aVZg2IAjjJMVOX+nikncCabJh9HgBFTn8VCFCholy0EbwWaVJmHxT
gCnVMhDmi0nNMNZwcNx3UqvLm3G9M1FyJJaf/73WwUoHLZEwQDL/19gJ6QUbTYY9
URclc963sVugNsZ2yyoyL5nvZ8K6u8hU3TvXWmrMqayiXAAgymXGhMFXAPNEN8Ku
NogfQ+KBMx9+CwgLbdQGf6VVwykgIaNWA3+BH5E4+bwkXZtvclyXLvLhWneSCTBq
WBEVFj6qnTBF7QkmQi62SKUeGqtBCemGJ88HYc/I8HL/LAN0dBZPzwlOUSz4xFw+
+pAaTNFlkKJNoKlburZ6wJGCZXfv5/lVD/Zm9bZ3A7oY6gVGJFQH7up5TyNOXD8J
KiU3SbXxkFQhDtfLkzcw6duCo8seCDlCzeREYvxYnsOUb9bTE8qxtRM9EH1aAF8Y
JLLUwYma3D5Cu65PG3jionkQokqs33CCDFKGVob0Qt3SOOWHKaoSEsmr0vUHWJJz
OByW7VjxJuQhRrQnVTVOd8sWNJvFiGT2gt6OS/Yv0BuJQFWWfmZ8yPCQyhLK7q4/
ef/GwXq7CaJ1UoalhXxRzQk/Gvq3cLFcf3rDQxOKP0x9eHKo4czfBNPMV0DNI70P
xpdRhO+ZNCumsiIFkaVao3aorUFCSyKBtjLU9/KuLB9xRR7zV9QJFdnjqcUjO7P7
WBYBo/gCQm904fcDt5XFW45z8/+kDDQYOCEfIRIyWWaN+GbUJroafTfDANySuFb0
EHayHL/MpU58mGMzHg573r05Y8RV7tMVwtCNqC/sVzyq3+W3jJDixV8pkPOUW5k0
yT1UL+pX1ayIh+x0KVzuy/knebIDueUyOvZQ/qgyJ3WE3ER71lQye/lHEpCM6B1F
sIJqMPdv0tCwFSrzgMhE4b1N0eqv3dP4lEawUlEx7euXNhfrL6vrs7ue3JeWHkaz
BjvGT57q3dwdP6YqxGXARSsDM5ONDx1masvdwmKuw/p8gG2YVJdeDnuFfbvUcuBT
h2C6SjsZyIFy1COTxXZvXOleSMwNDl22/tQmCPfYkz0r/BCn2BwFZiR6OBnJPtgP
CDM9JSIa7iPtAzEOUvDqdbqIKHMUmqjtD7j++Gf1OqrxU4SSKK1QT0ySgvkrmPcT
fgQOtCEnvr7VMZ6N5hou8eQdVAJLPtWNF228qpAXXQ7IMPX2nLHONWgfkhUjzxrE
f+CGofOURAQkZy5f/Tg+hrFaprUVb3tTlcoK+MJL7yk5CAloWV1zQKwTL0fKIkcN
FrcIbID47+YmnkMOYU6G5MtjQy161NC47TDxq6+hBuyjPgtK8i29UAB04cXgMZi7
vlT9AIWs+37BBCjClo7vPHK1kWyzPAPpvpVl5wOxPHdOUfn4MoE+bajy5sgoGqid
zzvGHs3QGSSMrBajTN7cOVt5b244KTBd1xpziaIZpgl3vthuODnJCnqjnPAtO9dS
5A1q6SPIogDr0R3vIbG93VAbsHg8v/GME79wziLjpkth8XGDOHbZr8ELVqCk0oFJ
UEueqmOBcDEpuv5wWn2se2V0I9RVwMwAF/K2MlHKCQZNiDhgFEHOmxYqIDKZBFRS
z6w2xjq8RLGQVEnv08TqsGOCys60M3RZFC0ZQJEer3jiKJFz4BEzVpltBCb+3NIk
yb/jDqSijMKYmgTR55bvTkh/HRkvhuN0sBLW0jJin/JTscoSBJ7ne4N52ckHPc6c
G06nQp13AhrPJBkv9p3fgkFdU9dgpmXmqqfA1sR3+UA/dPL1f4mPuwiYQA3Z9ytU
q28pdoG9b4+GZwRt5zuR7vSDVL9i7Xlhcj6tYFaH+LF92sW/zF/E0LTODabVGvnp
TzwIo2QUMB4BTYYDljRM+qeQi0IaBjDxwpP1DPo2s/PRowMso82VCWEIM7b1YiRR
2nK/+FvSrh0mmYY8enrFSQw3GZ5CbLELahEkKC/g4IAWk7rL0NdOBbO/LVc447bO
ijTOeDVs9qU1RzrqIdMPWc+wYOEIKN/GgC9lR7qUgPSM8gL9ZgztdCSheQM0VRzb
eyrVpvvGgT6LobEfJlQsL2cL1QpAIB1hsd5hHQqz3/4gS/72KaCaymsjI8f/z7J4
wzH1VRhQ/biME39r5o8kyUvWCI9QBOpowxsk1HHQYVCASyvIOXVaYzqC3dJPzzBc
5FCKfkzSF4ImG/wFLwujQdqW8imJIoRcOkNrSR5f8fqYZ59Keu47OwT+tpBJi9hh
ieXifZocdjHTqpNg0U+TTEYXOXQSisgM8TObw4n+JOLG7dDHLpS7h2ajrpi6y3hc
oozd+iq2M/Tu3Th+OvDeBnxZFL5QeR+ukaUgrI4+vFmktAhnb2aUszt0i0FzrFZ7
SKgdnXjr21Wkp4rYGc4v7mQ+EPVRYVWx9MvEwciKqPrxmBb2SxHrABk82hzPDelw
s7AUG2kBIRHcWJ1WgON1dMNYtXJlhUPR6BEL375y+sxKtk1Cw2sh1unjxnJMnqhO
CZgwf9J4l/ABppxxUHthKMNFCsskTAbtAMibmHUMgqx9+k5/njtiLLkSjZRaUO+6
JC14ZfOA2bl5fHlkkjF/ibpUmnYMIy/1FfCJ5bPIRNHDL7Vf8p+I/UosxWzlWsiJ
ms8Hc75weaXi5SFBIEF4mLMVisb8Q+uRmSQynYu3NmRj17araXh6gr1+dWw1LMQ3
sf8oHNJCyNsXt3yAyJk21AKHqAxYyl9e3cwHDTJgRcSu+hXxGirh/jdPxUeNEEsB
hVCz2SjBan+Kn9CmHOF6JpCjW0Ca1H0yMlxYJOwt3lVNw9Ut0WYZxTgVQ71i2Jkx
wdWc8TX6vFM4V2jljHMtrUku9+gswCp7mgjESoaJj8HoefPgo7DWMTlhxpOcRbKa
in6xE1/gifupheyoo5rXgtiwXmjfl6NCEdw4TsXvW0I2Iy6atUOcjVIvMV2d6LnM
P1zPyt2HqQs95iQAbsRliA36nVwIL3DAIdOSHfDiWBEn7mRH80V8votceMSuOqHT
sW97qvei3Ok4kZJHsk2NoisrGhtPGT3sTElbHvZFpxmCTJu7kHkTdKZO8CjI7s5k
Gp4qy+y9EHfJVimZ22wsz/BzL9BR6v9OAZaLX7T2sKt09KrFUJqWVdQ87Kf08Vs5
o9KD+KwWwHCivbIPQhfrQECwlfhg14VKhcwYmhfTdhfXj9WD46/1tu/lfFQWVOq7
NtGuDpAwxrXbSFGnoZTJ7bHMnC4Ym4IRulICc2+U8GwSRG5dkJPVO2Jy/5JD/GLk
RyahHQhM6rq5i6gtbbe6xZMBa9LoiU129Nx3UVGqJiYPXVfJ0Fhc32SBProE4idJ
WSZAe6rsmPLOQePDvkiU734ZdAyk/fU4raCNc9086/SE6qmUmCDdfX+36R0kTOQv
B91Ol+7lDqUxasJCRUcILwr1/CcqcUlezZCaBzfHxi7L+dTRRokSomTD6LSuhr5d
EdoQ4sZJUIaF9gosMzWZnDEQeFGBROwd8KA3MQe8T/wBhjw1oFEHYhFhO0tlNW2f
vDSLTLXZrBpDFqtz9Iwp8dzUbAgdwZDkDwafGojkonGuDd726Oh/V1Nj9FLNL8kG
v0ht1XOgwEkrOLxECBjxdechjWznm/NAdvp2p9v9BvZZChOBsBv/PaFN/U0S9dRm
n5U2GEBYYrmFcqTJ/eC49c+Rih4ie0fEzGJLQ38EiB3i9aHIBKmvj54aQKFUrCKL
U0yHZyVDlVNL91pbV2Y4DDFa30ufwXIIYHylpcesgjJcVCqvxLKG/nlNE66d8atN
WWx2+0MjVvaQHtXpiUmleF+kVqMRHzvM0fJq9XjZPUAhd90LnGfEYTecFIkuuyXd
qvKgFVLJ6Xf8udyxbIPHneRy2WDiW5eUafOIiwRY8fRf2+X1AOGGytmYxTAgWlWp
wM1But8FPjHimM1W4us4SJVrcMml2OKr5Wkt/RcaGpWQmMXCyT1Q9/wVO94Wp/Sr
GQR3Jl3jSWHFo8OYQZELh9P3iYREf0w9V1l8a6rwt8//aclw6s5ZMK15uEWC7H1V
GFtQ1nXUc2+kr6HP5AFlqOHqVIqBUPU6/75ngWofJ6jg6W7l+u1Nkb+Z3XcTIbx2
6F1eZ0lsjqdESi1LpwXPDiMgA2H7eLMMf9LnuObEu1HfJoHuJhLmGh8XSpOXbKMF
bYmD9xDmHL8J1rK+Mgv1FCqYGwnpUoTp3mq2glAai9MtrNRx+zDmAe2jzZ6f56yp
xWJvTA9Ss5hw0SfDa/CCrajlRHxTvWYyPvi8HLklF2+87sslpT+8wsCz2ScbyhG0
8JcIhH6MXmQqwdeF6siR/C4ECgfkBkHpjChQKbsINfoTzTWJAMgXjJkIFxUhKdwI
oaVOy7ur7PdrdskkR5yEXImZttRUvDD4plZsg+mJiN7154Qmr9wMEAuP1kRzW2nG
Ab9QMM5LiyPi2mXSBTwdVXNbCHFEgc9mHIljdThVV/7bfCth1N/7yg0actEWk+YI
vg5WIT8+H6VXZ7/mI/jLgM4inlet5g5QX7j6x3lctIu37JU86dRo2Wwr2GMe41Df
nbAP3vjwr4oyUXPr7bV7GVQRBsBbRFBe5OdP8KDR8ENZ12aeA09/y7vmSf65AvpP
UaCHZ3QYut07rb9bDJhGCyuPAsLJaO0Ovarb8lAhETrOLH9C8GRwjCyEDFUznTpZ
5g3+WeNVl54Lnb6333uptKvFpxgKNEDQFcpNF9rTC5ksjlz9wDmdICN1IS0cGq39
xyslri5SHb+U0Y7zWErgU7oX2o3OJ1YGGtUlrsJZnTrHe3GRspx9xYc8V5lRS2bv
wiiADOok4EQdM8gCpfm2il/AIghTe9r5hUu4RjVU0nD3ozdkXlRJTJDtIEGzwL/O
rrCfGxM/ZleB8+0Y/mSPvwnAhcSwB7p3IraWs/MumSj5pbMqVhwYhyPy8En9rAtH
rUUstrKCic/b/zQ7zWJQpKUvziRKNdxWWlQZsN5pQTMO3b7gGhIPKC2zVyLcWYbk
ONgsdR9qkH2Av7U3zSoJe6iCtFYb4RXD94zEBhSbPGgvVdp2pObmmwlGl6Nz5p02
EOzHM0BDoT0NR/tLKNpWtyqbMkXRIOYkwG4oMXda4URKLiGHNNhkogaKKToVKwOp
pXAGtAF/UzrkJfOJjz5OPnmcoVlh0Il+AMiD50dC2YBeKPtWyF7lqQFEK251IbwU
wX2a7fBpQMxciHHxCQG8+wws6c2qu0e8yYnZsYBRlrt0CpRMzdukSRmzqQ2CCou4
NE/fuRKJKuj49xzPuV38rTVDnloRaoDqfbBBMkw6Zk4Xw4bEtd3HViJyvPV2ajZ/
iPDrNoQlMPP6bFnz2XU+M+MMRqJyEDkGGqzlTd0ZGS7vbOtnih/E3nsmCrryFu3E
fipA/Kl/qCsrMjxm4Y3H+fbpVwBQkdDqkhvMCz8Q0nWJx4rFOfiRF3xODwWklJ/U
AsiNJ/j9ztv6MKsVPT7hcm7myusTAd9T6BGksE2AuWQ3nHKDvIBe+qZKciUmsWfH
HmXSH0uq71hyaCe83JPWp/zSWLbAfq/784dHRrC4ccNYBYAe6jOPgGbnV3aezcLh
tci85oPBkxDBS2bpLMB/XmLXEsaGQgDbpYPy083dPo4A/VRaKz2uiipNg4ic/+3+
mu7aU9mW25o5PZ3d1L8TbgQ9yzcLT7iHLHRWn4YwTt590+kJbIn5XqLSGU5i/NnE
YfzauiYI8K/ln4rFhrgr54CL+czv5D7cgrOi4XGKdUrZ4crqT2o4BPD2dtZDhcZf
7fwXXqBnAg3/BzXhyvogoe0c7Dd3h454TwDFPinrNMnXfaAuJ10Zm9LYDruLq5Is
mLDFMe4ap69pyIb6iK2Cnj5o4W/Nr/6KgguY793RGKO0N61f3/I0br5pSPu72Y3d
Ouf9jTpPQKrQ3cZ7O6ZzxB08b9w9UF39u2aydB9giS87b317EieFUT2qUCLvlM+b
Rwu87pa3N1qo6YD+okgfVBkV3lLzNHOmjsJwZ4GFYfIi5/WQtgjxhJHvabu7BpRd
GRLqP7nngIrQDFjFogTHzT0QimTyse4pSAF4PwDwzEfQTBw9ZO+LhmtUKord/myG
Uj/MveS62NuNxM3mNahJ0YF54j3WyNydSp7Bh3od/+amuJNtFsbMZMqNiESfzp1Q
l39GEGym/XViZCfo8GvSM1TqzEzbczbY5fqnAnvop5gjusDuaGRMoXD2uFJJdHor
e9frL3JcLdEGjXa1rGrFPPK6Ss/L9JYD1yUfUyekRo0mli5sjewcXjsCnQF6NNwW
DsyHq01N7s2FzB2DeZnWB1oOGkgJnE7E6KWYgAg4wo/0Zq27TzlJ1HRO2f3732Gn
ZTWVdD59zcl939qYiDtlIMHGr8wnnV4RynoHZjIIFchOB6nDXHGhA6roKQQejw1Q
k06fbwDVPwu2mV7DrR/MaRAe6myPS57bxTNzOinTs3ZwnE80uKCYTwQi3XsyLpZb
uaoGarQaLcdh2YweYYup3QV+rnpfqzfFRYGBA+r8bxFN+VTcE8ko/mJNs8ribT9K
VAUZevEeY4swqw3Yo1RV0eCh1rKZCa3NU2uvdkzaaN24EM3WdZRV3REJB8xAwaOb
UUFYvfQOd21JW3du2qpbVeZ4rKPGiMiLwlgkdVXDg6K/whMPnrtBlNfdCugGOon1
pofjXs3UjMrpDtkSr9K5duLqecFEBLmvDGL57NcH92ezYbrOVqK7shK+IfykCJjW
k0vzHbLexeyTFyEC0+hefhD7ynK9i0LNHmMU/qVCYrWYO+qL28Q9otCvkhLC/EzR
HIMESg51tL/Y3q/XSxqtXcaT4HqN6BdoBw3PWxU8oC4fjDeBDmAkv9fPBlb7GGCz
q8BlwrptgBWH0nh7M93NZWgA+B9AANrBB6Pr/BMoLc3BMKeScOEmLdyF+ThFDlfJ
GRMMQP0M9e05lixZJvCAgp2bYJ3/TAlC5vm6PeHUJ0wrjUEOhtzmj0Rg4QPN27Jj
I67iudwa3kbZ7JT6jdKYGNSUmnnA2vCGygYJ+g/yf0Tr3h8EXlayP2CpG3Dt6/Hb
NBK4I7IfkPO/1+Hs/b8azzzW6paIQgF07p+qw0zRwsT2xYFkiRkUnY0jgpzSQBKM
CarjorYWe3nmueBz+Pbku+D9/C60FfSk6e434XMhVePvyewvj4WaC6PalFEMknsj
rOkrtaP0aInpbdPRMWz25A+9Kf6pBsMpZlzk29cG27L2PGc3oxI/1NNHe2mY8FXm
P7DzCmcf8HGkKfs0XKou68xsAhW7rZF6VQCVpCSzDRwByozxUPuf/YJh8D+Ga/jN
5jrJqYGF1PvaC/+q0QlGHSaWdw3IGAgIIK/5QvVrRUPriRTOtgl0VVIXxhhQ3Aa/
/Hn81n3BrrkxRxptW7SdH215dcETtpTjhhOrHG5rrs5uTgaIDpVFc3iPDpWyrGEm
0wscOwqPxZ7pX6/X/zvw6IUFkKU4hYSuYRPKpXd9ADqLKNRQevbvgNhd4M/hoATe
40uzIZ0hDtttPv+++JILTaKYJ7h8iVFFaGjK1h439hrkZrEhk+xE4T+9AWdAmCtC
fBbH/l0pRv7UiIe/JE+F51ZPCx6fTmpkyZydoaKN1/8mfBZWE+kDIWaY4DhovYrs
hUerr65cetIQ8WkDkoWp/7MhAFDi117X+FSkoIfUP7U0F5AYAXItZ2aXLD5mXy+F
R8VvbQPNkbaWiBbMjforO5zKvGu5SlwZjy2I3dBk9fUR81CKdbUQUrvPEzaPNLIb
MHT67FGzPEA246+nHo6GW4tAA3sSB6yoG5n3pgBRCxCzKXCjs8SG5i2hPeIbSLX/
DPK7ZCyPThAx+mNjFr2GI2KsVcDwL3EOwKcBLKfSyzbiafB8dTnQJBMVhijYrhId
o11WRmpxmXNb4N0sv5eKtixVEa0Yxjbf65uMGOEIDpH2oDUNLphaTPnRhtrMtvGD
mUP1o+oZ9z30t/ClVtClgNyFVJijqlfGr/qG+wtcwQjCMTg9QT2dXO1ITTQMTBHl
F3yFD4kn6/4mWTfK8ymSG7mVvrcw3UggSi0BGlceq4lM2DuigqiohcnwUkZmqwLt
R6dSFzH0X0idfrqJDFjW5vBlXTT9lEEHHseWuZ7ALiiVI+Oxbrd3QmU6Tl0HGMHD
LnnnAcpKXjnga+moH9hRDu/UOePhAJyfUZOEcHgjz5pQ6fS1oWuYuK6nK6e8wIpW
/qpaGHmY75DreLvpGMKRfLofnD33Uynus3omaVMSVZUJwOFxQVIh99PZq+E7uPfU
PVPw/aGjvTo8zc24lHEOnFZkFvIYI5SBlsv2qsCjbalObsSegs+cQjQ3jmUs5e3b
8hHnTx0EvqFNY+lVhsJfhaSWFDRy1t8Qp2Ts9kXp9GIDGt4hBE4g9LnTj+3D8Ado
HJDCylJErbaUtTOlKZtH+eT9uEemasW64bwsq0o+E0ise7VnGVtrsNfETYSt4gqZ
6JvzH59BzWor8bMrifciG2yIH3DB7PN8SmkqbI5Q3a5hHUm9kh9oVm+aNfd3+fRB
HHkjm+l5GaYB3nkouENFQnKajYfKt4QF/LrImasULtkYIXVAya7PVsQFLellrTYN
3Bsa46ryYkEzT7T2XithSn6fZSVHPe+EchRC5jwH31X9doJoNnI1FwdMtNgipE6q
1mM1nvJ0ikN5ZL7lcQIck9FhiMXH9gbjrEH3J8AcT73repBgjA65HvcddtX866z/
TCQUjs5X0mVAjlIp6d9d0J9P3/430DC7hIgS0MpsyTSEvqXLl4hdbL5DVmpFuGZq
Q0+8r3Tp3K37bjMNIMfaUa3PoibnCQnnufM+8sXiU1BHIdV8mAvclo7iOmgoP1cG
o50ed7a2enRoA1NNk7UOfm7vSFu3DVMyI7l6ag4f1FWLZifvkI/C+WAHYNSdytp4
AsSjhMSfx1+rIQQfJWfYkHGHR24NAAhyPwSTvk4V12R3HM4t3J7bDTUUK0m0D4Ac
aEhKkHUqvutBX3I1djla05Q/bNWisPLrennoKAR4+vFpJj011yVtTQqAcS7dSzAo
kwGG2axON6aodXhe//KKpVxyRbTQSo4vEKRHlgdOu/PkWpvGa5YseCH0YJTQWTvK
mbeuruF/1/BDN/HbBDCdHZkZ/jZ0q7d3oreF+n6mHiJdTnuWUNe/kRyUmoosX7hz
Z2i/ZpNGZJu0C0HgD+XB4V/aTQHyUh2gv4JL4mx6AjLBegw/Cg3laCypXtcSmeJP
aqz3wSKyggvRmPxzOKM/rGp33UpXgQF1aoZW9AkMWjTYLkDWKnUSn/GAm7pT5so8
HZV7/013gnF1GmSQiIa0l2YF7vWp4tzCGuDfhf5/+UK7HevzrBNut3n/5rQ82raz
6v8CKB/IeCa9KYNLYRSuEjKDwzWkTbuu6dUS+/GJ6uvNUPCL3uXpdhcN2x941qqz
xzDyGR45USbzX3+WZNjtOKSb/YV23FKls4ASco+T58ViguNWxtRz5UlMOM7dtsdD
QQTZO/os1H/iLDNhj8WlQ/97THotz7H2Q0x0yf/N8gRv2we2fo7seQ9qwaDEhETg
DnTVg+lB3KCIVQxv9KZf0FFaO/9wu5IWtM/C0B7uedRKWoWW8wIRZeEg6rn2A0g9
MFbKdhnsYtfo6rotFJUuBdYqsNKsq+nvRGyN4JPJ7g57NoVWipCnA6qveCRJ+J1D
HfmRMqOQtAlOZ3fqjhjooEmi9CVc9RYpUPKlLt0tPufUlJS+qFyQioqMtrNyA6+1
Wcc0MxjVqMNGoKEghdHFqSiC2X8t9MFFLAWb8djKBzBnrwa5SgETjbSzDFEHOWLQ
tibIYu6spDZMcXSs9WSjmYUZMmiQUq4mX9msPVYT/WjBMwi5JN/5DoA6ffUJA3lk
nqDq0R4wZNf1TpaY0TCcXB+3oN8Omg1rHpV6fb7swMj/DFUvu20mjj2m3zTKNLBh
Uh7CeAw/A+c39fLugD1L2uK5EqOlrlmjBzZ72ayL3yzEKsK1pbQZETkKKaFrMq13
fkRphh0qW7KwfNuGwhmNVEHaIkGwWZneE79DXvU/2tfH2ilh7FAldxL5Uvonj47r
tcuap8O6HD4sLOd9Ddf86ISHYn72VIibZngT9TKkUkdiD3Zzc85XlT8u389yNO1b
yNA82kC+fFqwHPutngWEV/9WhYEV8MYcjqbnuqCLpox4bEHGHP0aldZ7Ud4PqKuz
wOss+0YgW9tOM4ezhZBXgOAMhKKScbhap8eTJWbmXLX+ZP36I66iTp0NMiXOlBG9
qkNQZhBVRY7IKypJoCJWXSRmwDGno8hCEGFJkULC52/v6j1RkshJxvO7M1eC0NNn
8wi+9OCEfbBPVfTrVRHrUsGnn658MZkv5SyDhRSaq/bXlW7YXA9e2ZiwH1TQUiTw
1l+QwEIIgeyz1igGeb7dDgilhyAc4/KgSuhfPwnCysvWmL/oozO9tr5bBiFFNafB
IJ4ZkZV96cNYHCDEpd8uo5xAChl3P5CVasMNb5azNXdEhPZvghKV0bZVe9P7uEO0
xrEMQEAfDPPIjBI+xcw5HDO9xsPMXMbhhX/DxzOlnMU01XPRKORhJ9uCYMNTy2ot
XRyQ/83a2/RxCsd05w6xkxKAt/q74neEFhoEUpIQEQnN5359IbGaREhEIkQMx5R3
v+s6TqyWVkmWo6wrUfuvhs9WEoc/Uz4drFoxloO37jTkpyxy+ITXkQexjqw1y8Ix
bmCjNscBpKBoDVQS1flb6ZAwt24yadl8DmTjW+BCz+GomFbDwcFwQqLRkyKmF5Pq
O92BgOt8zJ6fOAz40zJkVVy/gywL03JNQGTC80IwSdpai3vyN+4PBuBvPbWcIEny
ulVLrlQmv/ueFtZv6wbl+wBX1crVg3KnLXa2l4+rIvWYebC0+9yb2HYmUcOTBuGY
Y5DDd2S2/j7UgZx8GRstqIM8ILkDtUUwDba5FmebJwVYNWwak1PD8HgcpfGjUn6y
3OVCMwvQsmRhfve7IVotw5RPEyPr9ZwfRh/OyUC3sTTvrYMVKDNexDr908FWTxgJ
48wZFH5tZezOFlA7QC3wskX9uk1KLFvYnEMgE89x6quD0/gocmSpL1yqLHv6ey1R
hdSvFI00DTBstBGiNaDdVl2VtquK9Vzy7vjBwwxowckAZVzf+X3jN+zGS/w/hHcV
jdRl4v+BRoMP077tkOGh+NqRkPScrrOZo2Iebwm9gBAGaVE7EhX120JKBeUF5P21
y4hKq7v3YvP08svHbfH0LwG/vNb9WFu7Y/LGuMXvNymUik5SX9mKKCOCwmhcmHXi
N/aZmDfniDpARsnMLWvH+C+NgQMFJOWc91yfOiCarqgh7QM94Wjg3GIKCXZ1MNK/
gopvqzwec9VnjPD0xIDSsy5z8HPm2ApIpi3Piv5G3QalMJhb3UbnwhjlzvVqhyjM
VgwJ3x4FU1cMBivxtmeXP+YeJRg3m+fcRkMBVXAxVlu1kOwYPTYN7RGSYaNux10e
60E0oWrdTVSTUephC+ixesxDFzlnmQ4EpQtXhe8Z2ILPTINKY0a2vgFIT1hpLlWV
TyD5U+WuGVfNF68I900KYoY3eRQZMZyjfwxA/9r/qu0XhI5xwVaQoTsRqUxvGRNJ
y6xNMzdEylbn8eoAUgGJMcEBUuzjLtXYoZMyeE9cUGLgZZuodi+wAFTpA1J2Ay8F
7WvqEd4jDzWbKiKLwskrNSCjNV+5brdZ67GwLmoDS71jstwHSPonYo7HxpD7Em97
rNqVzVMiZALLftfSq72mk7KFel4pfAIR2i2aW3vwPVl7+Y+32S9uLl8KuCyxiLk0
aW8QMoB64ckwky68pNxMkhBnCzDFMABvXV5y5NjpCpdVgGSkOqsZIeg87/hlYJbk
feqMDKgNJmhe8IyW83aKuwSKL27yCoP0pch6n7ElDUafcR1IEgpHbNu5e+V29fMY
YAuRIEwsbt8d80fERH9oTKSn5gzPl5jV5xUmZaw6pNhMhOs7B0S8tyRxK1UTRrXG
tN41Ti0ZGBI9vBtjaI9jUbogv48xW7l+s/MZpr2rChZMme7FtUJPz6kbzVlLLTfi
OTBmiSCtOlUr0QWcCcm8uGVmaxDsrJUVuYL+wwRQ0FAksUTA8ZgQGJ9RvDMJxFyC
ks8XBeQsjw2aIjfsSo85H5JqmgLaTpB4fAM7BEvCB288rpyjTZMhVgY2unRHTmPM
5yZFZ4lj0P3hYC6QHo5hJdNVaTW6SppncpKBnAAAteBFslbCWcPfuhr6wIU2KZJB
cYbIm+gMRdl356nkdPKxQYeUqn2iLTdAavQUJNoE7MxzSJabDSG8dAXc0KJvvo3X
jm7tko5b3F9Q1LVgAtpklI5P9tansl2jpx5n8KnqeV9u7EN0ozm3rWp8+YKCzOeJ
qTbpMD1Js5ndvEr06K61G4hk44np2foFMQeYfHF/jFUsZ5587RaygkcxaUhjwXz+
reE2xVzVNUvoG41jJ1bndHzgGy/T8sr5cn7AEY2QYgbjHKEDi2fuhG6/PP87C85d
e9afUzvFqi6Bm7mDc+DYqRZ9w6WXLXNqCpUaCrTTWW0F3JS0th0cAFe16OWIZ3hB
1huKUCFPBuAzQ7Dpw75gc+7jwHuSgKTuRY1UCp/NcPSLlAEbQpA5sh7AShfGl4SB
BW1VII1aVT2Qa1QuD+e+3r5T6P5nmyCZ87zAbqVyU6L6Z7D+31Gm3uTmrn6CDdNL
7ogoWBOIIXIEYWCjfWi9a687jEOrOK5Z1muW+rSjK+rrRC8ocB5du3fLeJUCbp4Z
8vcGwm2vz47T/0h5ritDrihBSUg7fy7bkBqo+JhxiN1SDxosu353kLceywQreMEs
vfSRIyCa0x0VIzwNCCPixik5+Z4vwO1eRmypw2MqjtocC7VxLG1ssfsdriyvnCbV
2tTVcbMX1e1ntb9Qqa7EN9hYX+h5rJXIvkj8WAybXpewW+BJ/fZjVQyvaYRcOzG0
xyMevWC6u7Hiur3LZdehCcuBI4ZDEwuAvFsOOWA8hvP/Mabh2YP1xluWrKORlQ7W
OpAPNcFK2ik1KFzxC4hmUHUonXxZjnh63y2GV5OeGSdE8koxS4nrWvE6ii6quNDw
/KzQBJ9xq3XHQTU44AVc+NcoWHQWt5i3ZW1AID8tAIxoeh564q/Wrs7g1Sqm5MJ9
AzX5duDOLLjjCm5KEqEmzUGf0hjZZgayRDl7OPFJCUY/eptilNAPI8uHcyJGB5M6
DrFumNdaQlBFwdLpz5FdcCp+aWApjUm3ifESkg2uRbu9c300AgvnVMx7qh/lyDQa
ELgpOhIOa5GnjHJ8X54fhjQppIKhvePiyNlgljOJCPQNnxTGJPex0vyn3/l0PRS1
cPJhvb7mM3b14jQ1Fqav4sZyQbxtc5yNvBFbJPEh1AxutAe4B3Z8djHImLkKN3af
8rm3b4ePp8D2Jk63GoqfC/kgCcw4nk9UKHk/q8t7cjcgQOKFh3bZNS7kABM/3Um9
jiWQ4G+GeFUE8QuEXSEUb7fsn2ucPah3s09FiMTHasCB5bs3g3iCxeEcNiRvGOSa
4YjhYNiRhcvLzTJla4KJIgc572/AF5bWlXoBC+w8A0GUjWny5nagrwqn7BFXZKnK
kR2cmT/dTSLx0p3Ph+p33X0pubwSnVQhU2GpxxvtPR3BoC+J7TY9eSjig7ioN5GT
vIt7O+RPAxiOinIG0gwlwfV0wlE8mdaxCDqV2zbVKPr7NRxsviPOj0wckQ7gMED8
NepavKFi++7Td3ZnnhxGmC+ttxGKmwPgGkv/f+s1cc6g6m/FLCP/c1GALntP5HhY
OqUXGLEmzR6Yr4Mwa/LTBWom2RlEbNYPzbWbkk37VezHtu9hs4agMFB9va7H4m4c
dnq4//nCcMDv52EnO8yu5l6O7xg2Y1vo1ZhRWjcTz+l6kPKp9lC282aDODnFoFSa
MF61jQHAjRixlajq+6zxZqmCNinIRnZHPCNAgm78yD/EswHFhryi/0V6CtDz3psn
7iMwtT4bFOb1yAVxPraECKEqNYk2zarMfIukMGzOcJHk2FBlmp8TyUeEdMHiEmQQ
Qdw0nlhxGNO2/SCqHx9N+ZYaOfxAn6A9whax4xThVTtFljh5WmsyaQib7FrMq7hO
5yojK6DyfF4HOO5MPQIilVJCDyRyPw6PnItjln99yw00qCOGF5IRxwU2hohbSZHp
CeiQR9oTf7seqbs4bZjX7gPP0r3stlBmZiP19Cur4bqL0/fkRlw7YjXgcpa/YTqn
1VqXfDg7KgHNYtFm7orDT1Stny3QByP4A+exiAS1kGndrk8xYqwbczucmyX/AToq
XwFv2CeZvo1R89t7dMZTzW1MT8oTXMampHryl9D5c+vM2hL8ygF1rcIrqSugBBh+
g4BSQvF7ET2UMz9ysN/V9q0SdIDui1wSbiRJtWlCKcAx5DrVz55hqKJ9ISV+vmyJ
znnu+yspYFDsWYw9hchOklIydU8I4Oq+dz8LydKHbPQ7kaWq3b7/4FJQ4oxnNox/
Pm5TMEZHYMZI/TeUJuv/saOL0vJpd16EDXI1cHg5TybTXccFXNxo4GKZPKx92BSu
crM7FXjWVwWhi62UbKnHVWVuL3mJW8QL1zs5Bbrb/N5v5C8ozgrvkq+NYUDfFcRR
V7TSbMwsoIy2lK/ZcxgPWDwRbCJol+rmoFFmUxQUJW3rCMCrzIB0BMZ4I6EmN4Ng
1oJqirgQ88/aeVw56IZMf/MGOQxNjqSgGrzZTTq3zZ28Z1oO2mrQMiTedCYUYXm+
VSnX5PeW0E26ge0sglJXERGwK3aNOlEeE/Z5K+XstPJaW6+3bkfjwgb5nLy03Er6
IsL1RlDjRZa5JPP2Fz4kgS8923Yaw9e5AcztID2zWetN5bKQREgJMlGiMz675T4Q
H6BpvLmhWOBM/jcdVEj9Sx4bqmWKhDhYkqUWPsREIZkHljnOqoQbrk5jOIk6fE8S
pVGay/N8awGVjBHL5JwB3u/MD/eRw2A5icGEtB5c1DNYAC4yfW5QpRdzWN9sHVXA
1w0iYJ8dgZfy1OWZU/fUaheEcm2AomlgkyEaa8VnA9tzl0GV6xDfFPbYMvLGd/1a
yMRbpoZioH8rcubwDIAZkuItX/RrmZn8nXl0SOYXS7eiLPRARhHo9hjVsWAIBXHM
LebhXD9jhF2hije++Zvss5JWf9h/OUj5WSm25+pWc+Q+nWnZjm9BwOjSMazYdwm4
9WyPIiOY1GVTaIgIb9eL7smmYL04jqpPFu+HvB9Ygr6+xBsKeOZFtRVagIq0qSpI
0WahYV2FwctcPwtNZZqIgaEyDvW09cZIb9qpwOfOMCLwgrmlb3AWiCjVQvLiNkRS
6TK3QxyzuLRlzlxEmRk9C9v5OecZ91/4ern6OBgZ3MS0KOvUjH8X0D/ogO+wuVWV
hudncwl6/nJ0cYUvkraOJRWiz4zHZzMznWT/aE/lvd07XeK4mIcYKDyVUxjvDpJJ
frh2JT943J6MaLKk2UBKzsXhZe4UI7uJdwr2qDndZI4FVJpCtIbxeMKgS7S634nX
k1LyhYXIu/9ePa69qpSDaV93J+Mh+v0EbHMC/fiU4XP5V60BvUPep9u/QaHl37RZ
4taLqa30WBx1Qo860em/6FygK4f9+Xb6FC2GM7BfdMUZLlP9+BdlZlVDqc1P2CDs
WZTw/D+relBv5XKqcQcpYhaYLMFOe5YNKgl+dFbeQTQBDWrihr5Onk2CZjHvV1MB
WC8dfgUuUMTGcBcMvM8xAAowT2J5TiUIAxkn5wMWhJ5hyZFBrWebYQo209pgu8nK
5Cp3HwwSFUWMDSf1Y5jopcKo88mWhBPR4dFKC1Q6a/40kYLcP0W3FHAvCpAdxI8w
AG1ktPFFTc4PoCnv4K6SWMpuREjDeBHrbvObzo91h73EoquXzYU8VtPFZ8Ebzz6I
lrxDGMrKROwenyQa9pnsJHnTSwumme+iW33iFIkM9dxgz6aS/mZ4sWOfWN36bf6S
28Wl7SnF4gfiaw/IDIDv72uWDxMg/6yxNrYU7e59xE5EHDFacD+F7yh0uccv8I/O
YRvCJzg8tchb75vUiG0SKJH164vIRik3R/jrtovEA017cwyd/LVmLSnN2xu3cgZS
po6J/PNjI6XV25mGGN49gSdh3eg/CW2E56IpYtPx788bo7FCO73kCFzciO4QJgwv
8rdfWlrzPW8cnu3kpyeduZr+RaxkIwRgQ7ltXYBgWO09048xkN6WVnrlYJDMPSdT
+OmT5akfDFKg4QOWAmBaozHSTdSiYKFu04F8J+SNjyMwNRBjii5KvGAGLYeNvaKI
kXoeAfXK36dvD1p93ZTV9TbbAMw3a261DB9bKJEZ2su21Bb9sAl/UcsYPPv4sVoO
UHs6eyBbw80EHCll9b7VsFAAcuz5yKs9I8VcgEHknFkeYAI5c5oeApDiXMOMjGO8
rev7MG+4+7TDl9VYqZpFKATGd+up6C7LHl6jn3gLeTchKZPVC2XXn20/8tmbFbmJ
hSHXOvqry4RvjZUJ67mNseYU3vfInFXhDl15T8bp7eim8n0iSE67qICDawW+lrhI
6DUnXgjnv2Gkr0GGVxNwuWJW6jDoEoC8abnYnf46KxW+rMiX7Vrbl4MQ8fmxyZW+
+6VZ64J9wyA8QTEX+CYq67zXP7liF1OBguXE1qPjs7HVojPPdeZ5KGIGhDE5S2/b
Ms4B11MUWmjfMq9I8uwUi1nRuqkCXsaocOy9cIiuc5DS1DCTDroI4qP2d7SXq4yt
ZM2Q+4FILYr0jPu9X2Rh6p2BtXGZ4kcWD8GIoq5zDufU6z8dYvRwSQFXJDok4LAE
2y5Lk/jbYxzZApQ2LPYduRqmTXvYzqPdtehjHNHr/5kMqUOryd25cNXzFT4CwDSz
kB3dHzOuA1yN6i4c2LfC0LzuWPoaAsPy8ZY0/lL4FnxxIBs6IaQ/SWp34IYOsAYA
hUXbpT+Y8Od8wwr1KhCK+2JcsJKkWCduN07vYcC5CBRBSvV4qnw+sNwcGDe8v1dW
2lNHO4STTVQxEtnBCom0tXOYhZ3lMT3aLzE/8WVfEgIYUR8A/X/G13TtnkL5hITY
nUO/TWK2qT1/Im04XntOcFZDipQPzaUS2+zkiNTwjovNpMaaTfX+7+MlCb8m2oQ4
v1eh5VU1pku0qIIfAa8kLVrM/dAU9XS9cvcwjTmU2MTLFUezLxcWirnFoiHZGQrA
+O82vSDG9dZoXRzZ1oHABbtvq9O4pVdrETQVJILahiWsWQFDvOlZIolWnjZ4LBRW
Ev2Pn91Ak0zZj60rFqxBcHEs7jQeRcdvTPCxowkR049gPyZFs+NCnMuI1G15/Hrv
5NzoPkB/DSiLINnlA9G0yceYmZBWamk/70f+Dhfa1g1MRtaZUM6SLpl+n8jS4sUE
sGa/X7J8hQDmednwikohYw9a7SxgeqwiUf5IpTbsazlaJQDXs32UCq3p2ULmAT0Q
k5BdGqS7we8vfBr4g9UIXi/AwRtAv0KcfrqcKqDfYLJcKoOJ6u35kbCT1lzN88NI
2P6wPnzo5anf+6f92qgCXhvJhFyOWhxzlmib1wkS/Uai0Ll5s2Utb+pGLzCsopN1
NaKsZxkPnrI2WKzE41ofP/1A6d8XTFe0kLPKefZZkfJ0im+S6F3M3NoVeoP0umNG
yxFghdO0tKLKvhuj78o+JcFDxdEEdB9IoZLSCGlzTJcbZcXINbG5tT9IyT8yuqY6
SBbQvaB8wO6xAdzgIwGcWB4F9+Cclz15GCYdqwNoMgDnsEA8X3wZECBUFY+HTwCq
P9jNBH2nEx3Yl9PDxV1tuKLgQba0L8m+mH8vQSpSKhe+xeBidtONReThubpbo0Da
QAvzRmVXUiaTzht913ylK7aPg+t9DelItRp8QI1pRZCXDCaFYgJwstkTEmMMgQRK
Phr2vfvfSFQrZ0bHuOR9Ugo1QwbKfqtrao1ADxsU8/Lm/ys2D7EFUjF2ceNxO2JE
frp3jt9CLLjVOc2FvRV8dBfKGoNO/DJXxCBKXxajXef+xZkA7Bw/LvgLFD+3fhbs
eKVgUtMfBnBfY9on1HtaWQSAytvzcqO36D7RigJVmAvqhlxZVCAohnumhlylws/H
O6E/RfD5JXAgY3++MQNFB6sMddZFiQCZbzvoGFpvzB/CQTNH/FyoKMdqjc6bgfeK
cYNjY38cOhEuOyDEyAW+mxypKQ/uwBXzAneJKfg9gU/2NjX1UiPCdd4CbiNJ7zq4
aEpdZQpeXGr8g2717BWMzSDNLeTJ2qRn8ftEb6QT6A+UOeRjzrRYNaiNo1vVrKB/
y1m2nWQsVYVd3SBjWrTL6HGzL5b1EAtqFOyunuHpIsAdym+t9XoA2BbsdTPNZc8h
vwqPTHduVn8LXhlEBUQa0TK0NvEnlKVJ+EUanOHtlvR3knoJpfYITLovgtmTck9N
fRCTJwP6qnHDa2BWUMEpewtiihF0WftXApcNXOq6Ma6cos5GfkCDCWAKM8n8WPWm
LVsgIJQPd88Cz/g2pi8bdtnirah3X5iHwgSgZKIsCGzVDonwhn0iah8VTOQsBOJm
gPa8jDDYsr9TDfjWLF3JfPGRp2vWeZWfaJKxJ/rWsEMZMcpBTQTKz1chJQzGsWXR
+GuIWt/u4SB6Q2Gz1nE2ThMGqNBNjet0Jyuj+iUPXc+mpYwg1+HgpIXR1rKF4EoL
OckfIN5R47+MybvRg0kjyGkdizgoPTTtdfZd6uTM3nPLWbefDPmDmrqsj5EqPaDd
UmqFaB3sq7E44nO2aldS7/W0yj0bRKExSi8vn39rTCSc9JhA5ZPkWBTpiMqiWbsz
9FaP9f0tTKvN5ojUA4yf61PsZyIETcffsOfda0AggtxsfcHaSdKnnerBw2SAIL/0
IzGJ7K8bbX/f8jTQAlE4vfKNCaQiaHAHolNGNXaDJV12ZOSG6NmRCwzkEO7C0FS/
DYg2huwChyqRpyyMaC6zYnDHEOOJn6TaksBorJ++M99J5ywOdIzVte9zfeh2iNpx
rMAb5DBOyNW3/cGSLGbm/k68WWvGFgAYSj85dIjdbCD+xw0mhvmguGNQMd1So5lF
bXwVzO+4bmopQgLs3po66X78zUeYKsMtGCIkj2yXvcKzo4PPsHul32jKm6Y8dahj
Xwl/UbYm2RdYWzSyh+rxmpgcUyVQS7aXyL6uzPB+PGcqSaTO6ziomw0WOKz53dFG
xJg3XPYMJESCroQQc85Kbx+h2Oatk63Cr5ae0icA8lyGwldjaq6L7yAp18Ha6yVf
4hYn4Rjd4iSACSjGkVYgo4dAa0wzdcyjTlIltYOHFQ5ikJYmp8fXWIsxHKIVXIh9
bcIqF9eW/JzOzT2qHAygX3/rCHN1xD1g44LddbcX1wH1WC7bxdydqX3PfBeUD4wK
VUWvp1SVVljuZlFSs2KvZSaZqm459EIvdTFH/NLHDppp467kKc0NcTnh4nD7JRyl
2E56Zn9c+PuY5bd2LQIOeI4ZTOnVP+dAG78vY4+p0Cac90jHkbFiyvYSV8gpP7hs
SSrzLeHdHcyXTCBkifRkj2ulM7lK9s5qKQow7/o4BIGtAePO3rRxTH1uUJNU9m6m
z3tTSYVlL2um7ktamWXafdjHR2TBd/k9V07dVvvzSvEhi66D2jKtp1gIBQBGtv8E
nOp1wYzKrgNCU9h3/XoRq+b+DitlC8LpbE9utpUvE+KOC5iuGcs5KwNrh8j9S5P/
zN0ODXsTC83tF7JRjceLW0sse/IAO2F5mZoUrR3giJSrB12UdGq1atXcfVrIA7G8
4CuVLZ9gmwQyBsCwHa/WBqhDRXP+pH4jQuTpYwOEbScq97BPefd+lfMhA8LdeHE3
tO6+CWSf1oUEgDVQt7S/eMJQiqJc4RpoLgd7AUilsBcoYZJjHh1CUFCX28Lp3pbz
h/3hhWQHPE2Mid9DkJuzWManqOKnhgj80TFuKoqcMoUclxW+orLneNZSLBfWDr8V
g2Pr8vH9Tx9rRK5w90xGvmX6J4+Kyit/b8aXURe3Z+S1dN9n7xCc0Nksw2UuYapw
uqYI0NRmdEHC6xMpqCaVgRAuSLcJASG9rAuU/HpvHbiHWfan/ph6rBCWr5dRlwrv
l6PGsJd/0CfWgniM86n3rjcGW8wIsVx5v5fRZ9TbfZSUFNkUT3M2DH73zePfwdqY
TGvyXzvBDLTBsF6nhAIxh4mf0I0l6ngBguLtYgjaW5bO0C+Hj2ZabJsRKpqfZM9W
b+cyi1JV43n/Z0umQjWWu4C7r7QXEIdFEXk5XZoCRMszLBEwAWZYe+pIWSpVTtOI
smnOoCNwKP2N96nJeEQTf67bMyURlM879eQBHmzoVqrNQD1Ro709/doH9+RSPeWK
k8z4mefdxLShsPbwN2nxixmJ1jDDIkgR0imFXlnxK3qGsAwpvluZH/H05cnLJ/Z+
8dAgdl20Y0nVh2b0gaxIMOX11Q44lNdM4Jc2R7goJNf5K2d169W2yCgldCBga4gr
2siK8ku+UNqbPArkzVmROqspq+5PHloFsin7mxQ4NRCFsS6oboyPcKGO/CPGGGoy
2mNkyewfQB/F4qKgFyI4iwsfCMLQa1Syc5jOh6AOcO9Li2vQHF0Q0SPWqR/pdrSi
zDlV2o2809tydYBWt5lOssVo5E6f0IQ/D2dpsE9laSK2+qYubI0VglCFY94G8zAy
RAzL4VQnAd4M0+ztuWgFiTe9nfhLQVCusPhCwg4U/NdSFrdC0ikCLazbIrZMHngr
SeMpr3ugwjdeCecq+KgshRi+FqCGc1fc8eoGxHo3wfwYZ3xdvNaQGptdHYlNI5oQ
pKgZtlOYbcHLlP3ASO/GJySuvf/B1abWWB3F712dw6epFVqz44W77kx0vAlp/3FY
hOz040r6+yTBlfuubaGE1/UM0DGHi0zlOA7ML94McAOwXouf2YO0ci/myGHHKHjs
tN4gt2PnX24h6V90ZsfhH4+1ySMlQ9S21s87l/gpOzWWq7zMLgcif/zZLS01gYs6
k3MgCa+d+nIeGub6T1cg6fBYizMoFzitQiuZfvavMylntXxDoAEQMn4srP/dflIH
Ylusz8IvOyynSnCy5hzP+8wlz0xqFGzQLZcL4PcgkC7W0VdMqy6t39AhzDYTefkT
yIbcXvmAdOch3F6lBBzo+gUed2zFFQ1dFKqsovslDe+/80Dd4n7EDdBbIdzNQRrC
AvFHod27wHBZnQIjDnycXxT4sG3DLj3hHWrZaaMSJFe0ROTyE/T0+qAhKqtHRQ57
xtNTbj2dD801Kth2BNB0Id3bqmKQyeHh1fTKrKHgxGh8tBlfZEDruhdPfqFhb/k3
1luq8pxA144U5YhO9Kipzg1alcURKWWyftp/rDv/OM4CtaPq/vppseAqHPDnRu0Y
J/HuX7+OoDhR72LkvNdLWctnbe77sF5gpgsxJccPTq3UDHYdsWVtBWVu0ztPzjZv
orwjPM1cM6AUTKyR9vZtk9ASQsV6Mm8pLoQs/J8E/zcrLSERKu0Grw226KEX6h4N
nr8Rn3XzRtFcAT9mku7sU1N8tXLZqVnbaq8DhH3U6S7KioIbw9Lmkfhw64nal3pK
4hZLnv5lvtSF8mbtobWxDxVYa9sXCCFZCvG4NkT+C4VWq9Mwd/EdsikdN3/1BNVS
8T5pkO1KH2XbxA5COqgB5pgCBkFlbR6epwbCpDXrfeUzdjjfpoVHcfh3J5bow4mg
oULBdd0Zae3uvj5YmY2mfZ48IZnnT2wXlkglI1l+4CvwOCymGdOOYtQM72TNhjTD
clhSDQdqC0uWCA97Y5ofrNQ/3lSfQkx/haT1tGkkgf4c8KroJkKltR2Vx1qZcUq+
hF0RTv52w3M8QaS1XGmjG5vcd8pznOBqQL6MEVE2h6Yfdd8Pi1j0usTOsNZiMDR1
X5/fD1F4ew0npmXBbPpWA6wVD4qqeLUtv4B5gwft29ajMw9dk7pT3BkMCcSebFys
2hn4THmQQpD+e8x4SxknxbPStLgRpEM/qK347nhFaHXRKApc1pDQy4GEqUaxwval
/uYuK4O+m//HGqq3p2eTU61Kazow/zv3veAimHDiBjSgk3FHsKpa/g6MVfx3HFz1
xRdy/RyWL2AZNF3ngesbk3JpYjlIxEVQd7KOjjdCcYThx7TT5WeM6EkCazhmNRxh
B3+uwn8LzI2edwa7oN5Gxu3qNPPoyvgsQVOzj2seZ0o98VSvMTP+MgMBiHqsx0fh
AzFA/LzabPyGi/Emy6MWX1PCCklwmGXDGs+s+/gUklbn9ls9ltl7hBkLDGiVfs2R
BS77MUJ0SJBmRVk8Ot1txsC36fxNadm7u2eWdzzbfbio9RRWG/DtafYzVR5zZFB+
98FmvjyPik7Oa4uxbc7KLBbq1RTHNyUR6I/XWFvGEG1f9USLSusEbYPAa8cvwbxf
HQZBM+aFwSVoE0KipbvgtFFKcBWqfLTxpZMOR4D1CLhoEWb4Nd464UP4mioAekgO
1l+jzkVjfw73FgLhcPesDSzHlnCF0UwqLRPiLdDHlnedRfewJPVtnOCshxmn7MSD
DuRLmBPow2BKEfUhj0qd9yMrVSV6pjQRuuqyGmVG43bVPigO5lnAv7q6rd9VDlnw
nv+ZsyiUEfA8GoZGuX31TrjWcrOpHM+A/ppnW1B/tSMjEGIrnm64O75JuZhVarci
Wl5m/uSCFl24Dj9Pmw0KkYdUo7i5fIm6nTRojtflp+iYsK9nj9BENM715/5L9FY3
6SjtjYIF3kVQ7PjrdSFCrDrJ09HoMxtdmYsQzBEKPFH7HMGNmk+TbNo27Bvlq/Uh
3Q8EoP8GdxZ+eA1UXflEWdmJQV86mZEghwZjR76TyFZOQdYd0kGzK1Lf2nmGKuoj
g7E4y7uRc7/3OqLAaYRRup4HO3nQeGppOZQXrpYv1aFF6B/Th0RuF6wkXWWD/0yk
XfpqtusPnRWoHtPPLUOym6OWxM9pCdCgHxWW8gR1iZQhhpOy9DHRxPS+IsANNi9e
z5VFwq3BXLdr45Qol/uYrQ/eMyiIjEqZGKyQwTfmTP/kM2gepw9VUvX3hCQr8a7w
qNunQsW9CsOWr87a76Euh2GMN6SijGlpTAPFdTn7ayNyeudESAvNUCzmrAjrmly3
LFEUn0C6NdoAl5nObd8S6F7V0mPbA4WRqLr9f0RE9xzKBTbVPHcrHNf7K5kN1AdY
S78RS1QY+mlJ2Dqh/Y6YkMXK0BC/wcJCGNBPCT6Uh9ogXawaVclvco2N+6Vm5xQ7
YPGMsnphWYrbHHJP2LLztZWLxdU3Ea/2XnZuai7LhzMuKCiRx/C11C6n7SmYN3ME
l8qov3mOoISG94KLB0H3hU/WThcmD0rOpY3fg7UKl31LcfTO6PN+RK0/OsXz44UT
yx9Gzn2AJjHVvijsWAHpdN+IfzlqeHKJIFOP6mu/Uu1HK5wpW8p2w1Y7NycQo7F0
eAy5DoEYe/kMdvZ3fzG78OvioZxinkaIBb2bN80usVOfXrVtqFxEz+8RxzBpHzSz
dkrk8jGt+sWyAydqkb03KQqfu3Claks93/LHefJwYaehIi2+NRP4hcoITVVjWvk1
vE7bHMYNOvQuVwp3FBMTuu97H8tA780MCNVTsBCosHoVzQkyAyWyJ4xBq0DJIXfL
eaDIiXQKCH8Mg1jZ8HbMaLF0Sz2O0R/tBCFxO1aKKGJr7QrEV9ihl3msIl6IanEQ
89aQ8q4hVZaRt/bnAsCq1YKdk4lPhcdsDTcwjFolFy+uxAQrn22GdTl6xPwwOEQR
npu1gGG04k1Sp1bmAO4c7/u/aDlgwozLQqpD0Cp9z/OGvvthMb6XWFsUqu/muf+/
zSuWabeqp1tU3yp9OqJhv0k6TG14eHD9bnWm1ZAvoiTUztvsMvat1lO6wncf9uk/
Z4PS7zvVrG2fI0aHhjuGkc3ku9hFa7Hi/x4YO9g4/1/oXXEHLxs9lAY069y2y9G4
ZwhAi0fWI8kXsG+xw4I6gGzrh00gOaJHYMfrAiuajDWesRY+WgpQvjAMS+/98g3Q
VMgJ3qYvxpIv21wL1y3DJNkccq3aV0ZYSEWb8xW9o24XxdX4rhq/6rAHwFfD7Mi5
ayYzyCLQuRn8mfQKMu5aFJlI7Oyre1EaJSk2ajoTilbleGM/utEbI8e+YZIOOPfo
hwV4kO3QuukD5GYagZOvpQfCJBiu7dF5BiGXATl2qU3Yl3ISomg2cDSrH8euDIWO
+qZZ9gNSo3inHcJV8ugLjltyyAKLDFCbobgVOprO04kuNXw2Zi+CTQFoQKTJTE7G
zF+Lw/w8//QlzRlnOXOWuRoOiMEaQMetpITBUCWRPybodS4vSN+INkGemiwOj7hY
tLGAf8Ak13JD4osYD+4viU02Xy4w0uMY2AGbmsrYW0Z30FXBV7Hd+XOgh+cFelSp
kYluuIyMqO8lepKY/icqOQFP8Z2qXwSRj6eQ+6oGXc3U1zV3qhseAgCdHUE4zY1j
LX3c5in40o7QXEPbJS/bbZJ5piHRWDgVMikz7xCs8TRzpWoZmH+o/kSgaY8Q0uhe
G5pbuYrHu7s0TVeSf2Vo0Hp++rNvrJYeFZYRkFNJ2f3nipS9z0uuM+pinFhcyhJY
lS/ng1PBtP0GehB3IjAZ9pOC9aDzC/38rEbeXFOit+Bq+CM61odFsnEtO3Xqxohz
jKHa3n0amniIfRCL3jUgKYsoy468ksPLe5hh0Z8CCGa3VI7Ht/s+eHmr2dn3IAC7
qcnrpZUByBtWMclIe8fKROCLK7wTQG9Xeh59jCvCBA/KP7Rd8Z11Iaz0ddfnWaZV
I7dwJDeRJvzJ9v9WD3Ls2pmUJ8vK6I7c7esB10Lx5iXTDK/8sL1E7m08csUL6nky
uVbrJ3xqB5pGCHKSf5XkNQVuXoQRJNOQblgURhzUAzIFOEWxJ3//+pMSiBKbeDzI
mS66OrUYNeRAjdXy0CNNlYD4F+2bi5MP+tzzdnAV8OChbyONq7uUCoQxcV3zk3cp
gQSvttA2WzwTQnxoijs4EReHYcSiIh8vVRe5+MoCKbczU4JDyXDXDl6jNuBffqOi
ZGllKV8nx5AGGlNbZg9fMJF7Sm+tdRljGMfA4s5xBGSloEWoA/wBkwZH+mVh7fTS
vZTBxfIWN9RsuS/tqTzNqNPcWVvFkIyRxsbe7Mdx7XSGz8HKqY6uR9yTMgNfN2ar
JFG43q2r4T1jLGLANYc74ppkyY6t0MrdmEMiS1Kn4zlj6wsIIvFU8qvnyieZkqgV
/4qu6pjbPyQs4bloYKzQsYfZqat9eLh6PLIzP9a4P9nDcEPJWZd9fC+c3I+DCNel
SABn24NSn6Fd9N4k364EiXer+1zZ8bme5ztvB6Gykm42Psdmh40Hs75LULkvPWEE
0N1/hGCWzDp9Xw+wMbAAW0z0v0wl2Y7YKxmq+zPbw2Sge+EE77XFKkgtxe1+ZTVU
yngXfjG+razDI9jABxONPCSsL16+723ux4rhQ2VkAlLIrvHKwtjH+d1p5hkYjrKw
h8MbJCSVHd2nvG1hc4w5FRoJy5jOGC+HpVuHzX4KUtM4eGGcrRy/xiqFYx3592x9
UZRQhPfqOdfvxhOe4YMYerDCmyqzQ7FcbNUVBCQPJ2OsJwm+AN5RdqeKoCnC4tML
Nm6YJzpIpp2gizk4qPquoi1ZV8L2m3Sb7OAxiB2ZIL+XveKPmgzm57/o0y69zIYZ
84YQIQ7iKGYT7eKMJsoltNQQthX+TavVmo+QEZJ6HQCGJ1mSKj1CEIsgtq3gIBzV
8d+ydDnTB3x5D0j03SSzbBnAAlx9Jdelvu0IU0MlEWA7ZiHsNLkdVoqjn21PUzL2
IgiYM8RUhxU9lr1l1EJn0SDv/MdEEm8JR/oHiA7fAl6ty1kA21uRKBp5LfSPZyv8
fkp/SCAIvtTDNA4s6/B+BC6hix6DQ6EBwh/LELf8XCgm/54fVERxU2E33JIblNhG
sL54kjsKtiT8F9vk6hh0Gz79b3ibt8aYO0dS0PoM3ReJ+93j1VWit5JPxB0pAP7f
OKRoevCYEmGDAFTmVb63Mnw0CCX7NbeA2rvi9tAIsjjxu2gCmlg2QKLTZQnWEMD3
gnEHjvkad+Ptn18RucYp1bs4DXWWWnor8sJf1UGcPu5JpxOgnk8yK1P1QoykqtEj
3Uj2nHELlvK5Wppi1zZvJ+1AJzCBTnYF6h46WLIJQqG5yJRmila7e/yGSNuFMeGs
OgLuY5bUI06vL1o1xv3A68VG2ba29jRma63OehSDMZYUrt/uMkpCTJ9bMRsNIQYv
iMKvYROdr6QutEif09D7lR97aNmNjhMq4DEFnXuiQa2eUgAPnZ0EDACwa1/v+UHw
SDMJ2toJA6OQchLye44VkyVOPUbOBp/GezoqHa/qEf5YTQg+VZhCFEWv8LIKgNiB
wKr1PhkHX6vnoJhQ/WZq8kd/PNAi4eMw0NQe7hcqYK2q6heUIEhepCTqZWxQ8g80
obt7j6F0abOoExAGv87JSg3NG1nyI3yCOFfiSqYmlo7/f3OsYV14mkMOCGuyNiMN
NPN7pZyA0cAAiuhnX8Ndt5ceuZ+X3RDpA6r81N+lnBJy1yP5kCiV4P62iTLozKi2
zjqx7sgR3mobhdzAl44NbIcaIRK2CmL9dqdFC+4spAuvJJD/peBKX0d9272BRdrl
yz8rnJQQtNUrT8aQGCCxu1w5YRzk3fM6p3yCAJEAjpIaJ6GOqfXbQWL6zxy8Fra1
NMiDF5LouOpzkCmbXTL1uOmWUvQHRFxgoi5bbXFC7qbF3cbcxLyY2fkXWopFxtTZ
q/sJntPcX24bCVa8B3NX62pqMk2tYAa1nmDfXWxkvBjoiwwPIywTSUrvQWYhtUn9
0aWCMHyMPh+7nQuKAcSPY96uZCAR+YbHfnDOdTy6uiPOhtJw18CHFdWPb7pP+SMK
AUdse51Zcmw/CMmZPxPInf5p28iBSubxpmJTZuGlqdTxft4pFsLARsX2MAZJp9tt
r4DtEPAhlWiGvrwDmx8Zq8qd2iti4oPAZzUP0a6eK+U5NEyKQSdIFZE9/CQaJvJz
vspFinj6fYp+e+k7A4lS69YlW6+2AHvMhSzmohIuco41yHzh2h4fHSI+ZHDX2ljC
xympz1ekDR69J+EBueKbvEGycUMdEz+LyEe1P+CN8FSwt2hFsWT7gPT4QwThTPCL
xZvlz7SFEKwH+7pmT95hxMGglAwm2bVBBo+dzVo/3Up2feV8bC/RqqiKqYDIuh4O
7rGqgeg2uC3ngmBMdGP0FuWTqR3O6mrRkU8nQDeIj0zDduEA+q5TYtbRJBi+80VB
d7X9KFiOuqRwEwqwDqEQ24yDDl68dpprVjZKDHw6TL4vIc7X2iTcsOkRfy/QiVkF
mEKlVeqZU+q6W3KbmRKjsqZhmPhoZ3nqe2+9gHtZWOuCnqYGndoAKG7zq6XaOqxP
pUQviMNnUojSqAKH76dkGZ5UJGmf9hDSDN7VFxbwTrg+HUuj+w6DdjcDb7C7MJjR
FTDKV7dx6K2bJJdn2GbCYu7ZOOBk6QtQJH2usOQ37I/XA8TKkFIfK9hkgfLBi4ax
dB76qAMIXqJJGpcJL5OBKSxJ5NjcoNdQOj+vKUDVnuUi7tOLBeV6JBQPT+cRABRs
2t+u9bcyJjqR/wrrGQyUpxY6CvTEERWqaRPM8UvDtFHrWlaNXMXqlQIwAkPnVXtB
Y891JduaCvZv62FsVcLG+HUKtqM6PT9DJUG5O6YtFD0JgkE9MUZi1c/jARzZ2JCd
NQ4YsSGF2DuyY6y+gTQTLi7tPdjLXS9bT/0844zWx7llws9aZNcnPbi3Bbi+mpbB
7XjTLOK3Mvi96xA4JQaSC+6Opn+IxX1JQy7NRnoeqisvhg9aU/CT5fx0SHfKVisB
4JugdkvC4MCXZE4KTxoC7virw2Qb16y+0AV4a1jT6+O1HXz+Eez6LbiPVGEFffFL
uZQiQmfyMmvBoQ+Ki35fkeWS0JJfXPbOT2VeJiKJwPqllnx0bLWJH10MPy1lGyyw
s9yNpiR2uAXm8EgsA3TS0jaXHH5ZoEMRihAuMtxU3DcX+BWFfiwzYbMxcc6LhXkL
Ift/txo2i9Gxp9LT3vTg6YD6pPnWUgyE845sYArlwZfS+5FuZhrCSkUOIEoaiGCx
0ImfyxnKBaUBwYz/dOqe3K1wQhO7y+CtNcM+xPIHtbgN5H/lNsueOElp+9x3oA2f
qE0OrdcVTSqXS0M/decfGo3tZbzIKwS/A6nPcasKKGCbz3rnJDVgam/phWzUabO6
EU/D8AEZni7jWkpm/9SwuseSNNY/fyC+aP2yFv7Y/Iwk3p/8SKNt+kdy/FWwqgXv
+DYtXYhjPxxrRbTiFzxGbIfMReNXeTK1Ky/FBs2IaQARX8T7n6JvKXG0VBzfsIug
bNepDi9xQdiERcb0wtpOOvv80BgwcEkE1wHi4f0B2WrMykMApXuDUL9CAF452OHz
ZbPsA7QqZxoc/vBeKc+1QZZTnJ54wfI5USLQ9cekJG8Hvkp1PJJ15hdxfM6aBEgT
n87f9jxe0g7zFEta31d2/eIzYsETsR0ed76KuY5zmT9TVmX6AWpIRXmWUzgJGejJ
8JEpVwDyGvxoQgvWEGp8ob1NwxZ3CTcGenVFR72kZcsvKLuf06mLWBkqyNXzMRL/
sX9B5xNKXt2e2DYSLk83GaqGNN/b0q8Yx/OcR/ZNj0jymQXQLGFW39ArSRMBGyna
wW9iKtCAPp3cJgBR6sfa8+m5o8w6Tg+3UXkV2q1/ULOgC/eEZbvh5HxU9v+1HGTq
arJuyMISff9xA75tmMIgR9y533AvzK2sYpYZ5nrxk8IJeyMhsMyzefHurIaF5xqT
aYUnkPJyd56fuxqrWSEix5IP/8Bz49bEzZhOmdjlMdVSSqzrGNtgg3clBcCSX1sm
/S5aIouFF6LxyethBaG2mIBmZApSUD6B6zQppyq3+GQ1IOzdPfG6O4NJHdVsmmUa
0bUra1waxBl3lXahl8h3z6echzztbg2qXM1Bc0h+FBEP9jp1hjT9oQknMoMH7ANv
3howZP0iur0lUnlXRv8QjsMMoDcgiiZjttVQtgwy39LHvfqJvEuGXOMgPFe68WSU
g+zIL0sbXrj2HnuXqRqHL/mnIXk56fMF0ykssRkvELt55hkyRpiS39+HY7JUPVrk
UFdxVg5vaSwauTjD2s05ulOM2JAMVOdqvcTnmpXYuxaAObHHiUZRHSGVKsnAWaNA
kTGb71BiWw19X4rbRl0RvkgLn2c7AbHPXjxngYEy9P8maljM5SN0gDivkib5ZsjB
fsqECFWPpuVFK8hxlJMNEU8Q6DDYXvpJM60O7pIBiJzLjk+N9ncGwLsa5mZvQr3J
LE3DvavB+IntVbeRqLSNGLSiHsqVqUBaZaT5Nz0nxvJnw3BGQkiHlihbz2Y/Gxmj
uiNH0JAxcCpK9bmhyOz9rEth9AL6ZErToTIj7Sn7LbguBgrFQHhdzLVFdmf8wrP7
ERcdiw2aoweeeXy1RgEXjviya2ep1jamwflfxDhKM2jtkWwUNgw5Nb5stBDfCia6
AG9oFGvbQ2LEIAn5nyeu2XXdwAI7jAcnQvdxANKNQpOb3k2yPsK/ndaq2NCvnaIT
eRlbAnA+V4O3kXTZSVhwBkCjvkVfVCraf0JpCSmSF/m4U0COJujL5IK8/agZ1NL8
CIvZl2838BxWV0l+o8z7S1ohSsSM2Diqz21MD7WrshK09RGuUA646+/daKW4G6SM
Jjo8BrUFGsOd69DO3faGReuymYPtiKjqhf2mqZkILuLcvP3mCoY/J/YqQ5q3Kzgl
d6a+lDdWvI566sTm9Wgxfc5Kqu8AJg0SVuzBDC5ouZc99Kl9UImAUaWIdKOGhaHk
pgsesybAQKl+Ksypn7/7I7TQ5mHUEGkcCFCscxYRMQEayLJCP0lIGA0TFjA6jUke
q43rl4mRzU3e+hLytrPZXAtmUCLx4FA6Xl+gJFf+wNMA9mN6R91sYENSdxPCd4N+
lt2+9bC6e6wVjM8yvLjQG1ugl2JOg+R2Md0ZkVAaObM27svDZNzVhEiPGvH41Jm/
1r7DPNIHTHz5DK3+H8IyGcfCntiTXEjra9JYFLPZc68fkJMAlp9ODR+9r44SRbOn
MPPqtbDt7qth7r/+C4+WUomjwo7186+1HkB06qLm3C7HRahRefCveRjuG6/hogyC
wBD5ft8mbz8C9XS30idcVEo+yNAY0xCpwv4KaLLFNi3mAjpYBv1PuL4TozVWRmVk
dtauw1dMAVRjyy4ly+A34k5F6+9zlZV0N+UJFQU2ACG956fq68MrQKWHjeFIABT0
P7fmYu0jPnZb4CTokSKkRbqnsXWdGF1HCHThE7X2qSlSikIv7/VgGPCEF9kI0pYR
m/UXiPfDH2zqcKtnKdKcp13wZvJ9qLARMcUGZFrEhSYagvWnigbTuEzhQYXhsH55
WATYT2Zm/ynqxlWj6E1qQ55QG8Xx/uPEnzDvTjbOfKMbcfGCLLbF+va/lzIgt7WA
S60iev24R1pO3ffh07cG0exMg8FXyRnKP1oYPNuGWb8IfqQyKdxe6aaFgB9tBvo6
bluXdK0lE5wq7Bso1fMZdIVCGM2cbZ1rEWyKExN5DY+PtOuNGYe0sHmDurqGfw2E
WtGtfVT9W3doGFKDVptfsu3sSR5w4rHMlhHyXm6bNNYyBBujj3cdv5zFVUgRN05U
yMIH3RERwJdBeR7asu2RSlSs12tXbc3OUiivhJmDuUeym6bv9Dg39hd4HKQq4WTW
/UYGfpBkRGfYWZ6FweLpv8Au9JjAja6iPCA8jguwQEqLZuISVEO2HGNY7ywY5sj/
FBwJn2P44moYth2uD/5TimL81r+TyL/pqXwBixQcNHFfm15pmU3yeP+o7NlhwkRt
kH/OirSjVMMgBLapBcwgf+RWVZPDDvlzdRDfCVlaebUGzIHclm4nnpRJwcneUTTG
GbLBq8PbLfRiXfTNbnabtt3+tWMWSzgzcolP5e/QSDCqRmuMPIPU3sr+xcPsiNEA
oyHgf4UZo2i1s9OlJoXsPXAR67rNdrjN3H4fuia+70PDcLzh7qSe3BdmcN3lYEmX
l2QJEMWTtWdVkjJ2Bhmu0XSyCQ7iVHV9iWoxAUcoGgTxx2xY4EW6itWZOFCObT8h
b0fUO2n/MfXgAgjso36O/L9BdIdKDj5zx07bzmhU7JeyM5YiHNpr5ZDHsqb4bCo1
0YC1dcUoJxYX985NUcdVZ3+NrJQI5VFJSpN5To7tqhi1NN9qkIxsJ5U7IvUVIxjV
Wzjg8JdZg4zMKUTCmIU0U32tcvFRNmzLLeCCHYI21o290KaH/XB7l2N9pgJzjsmA
Y/hsiKf3k9bqdG2sEJMLQMiM3A8ayNMFB0ENntXSanUvbJ6B3HajD1m7frciTWfr
rS+vwOAJ+1+YXG8BAgekYsqHxtmFih03IqPbbBAXBOYypE6JEUvwjni9eESVfgo2
DXT0jrU6KYkL7XfDsjRf3ZhWopHJemlepKp2YMAtw70f76OQv6RkA82SmeG0MHpK
RTRM5VyCdsX6ddjm3DXPwJPKWrpyFE8tWgCFYiiDzQuocZHbCkbeLIA2YP9OIUvn
EnhaXcrVwHvb40uDE80nfXbgCgEHU55L4gK/koFpIymkQvSDXB8xNgX6h8EEG8Y+
9zFFfvs6S4xH1b7b2xiAcUkQ2IBcZonyX6q0WCJUZXdNX17bHEfIuWSGY00XJt9s
DDGjwxI/byuH3eNNZEFmiTA5EhfC0xL8A//L95ZbLcFA4SNBABSd7RPELf4K4kex
FdBknaxvV4qCE2FFRFedocRCuYhEsbDXR9x8uT6uhBhCy2W4/s+X4ztdzyiNmp+1
2d0gyqtjaVJ+9xqjqSYvEaRpwezcBHEBjKMS3rxtCrJcRyCfH/21sC6aVHUEBloG
Q9JIbQC/eyUEG9VlMDICYS2YwarYfROw1A7JEQSoTBaxhNoBwEDQ8Y/1qrcrJQjn
5+dVhOG9MZGMFl7osw9y8+aSroiuEnqF8yjS1+w+Yvce6bl0XCVchtG76jUVV3gn
I7KaSx4bmwEqU+fYEVgEuZPWyKmQzX3iXCi38AHtYgYAdy7aNTuHFUmQFWmx4Fe0
WeKsll6ZMY6qa8CLMbb0guwSJXNe/vWnbq+NR/3HxHWdIbIAaAe8JAxxrJKKSlZ7
Gye0NOx9yPI4uI00T8pJI0ei4MsdJHQ4IlEyEIv3x+RjFuwwargFGnsurvnU7pEM
42b/+hyNToJghViYk2m9egG5K09UIqjpErp1rm3/Hw0gvqC4VCkyHzAm/TdYtQUH
92iWkkSt5z0HylDj6XGrtoSILyijU78AewgE5iyS+MPpJCUEWTW8Etyxq7SYx0qV
ZhP05C3h3EEeYDAAqv1/+LBA7Lx26sXT8pBWF4ObVLq+TQoP3zRqmZUg18m/qREq
gEhTqM5cHSsLn5v10FcWF9eO+Vayt4m82TanTGx1xSzZ636A7JCil1gU5A8s7ZiF
G93GtkTUOLwjXkNJQEQ43qyI4aFMTmJQ11dBgTAXyoTY6pj6bp4GPGFyN6+leWLw
mxMQMqYBTGAxZIUrlHDWr+YiaeGS4ewBj79++y6j8dcA+gZ2Gk+riOB2a6M3q5G9
IHXTMg0hSPO54RaYkc6jzbp3ov1SwNUi915i+22dqJRzh8/Wo9xdjSaWAfzUte6M
IG2yy9oqWU3g1xhCmBQXUXiZEFlxK9aTHBDMTsv7FFRtN9gjTpYUqnDz16FkpRuD
DcNjWOK6puRBM/J/rdI6VCLhqTPCC9EMg7+2QrDUXBz91Tbk2MHpd+TqEEqxt9ht
xrD/FaAEHrb2kVWuOpaegKrwZ791cuZmEakX+KdZNoKaYbyvKbR+Lxbv6B5LOxdW
Yq/QHoWPUn1Os286ap076WbQELUipj+zgauGLx/qU34GUltrRulQDufJTfstPiPm
8oa9ekh4s8OQjxVEkDJ47M1yPzs5PJGjhSIr1pS2xfIUnL4EaF8+M//sVkR6qdAc
mvSxhalMXuWwUWMP/floJbfvLB/+cq5VtHgeocaKK2eG1Ih1X1BO3jaoUC2E6FTp
p/IsXN68POOcohdw27KdDw9WoRITdviD3ip+liUjSpGVtXP+PXkUoBqWnHmiQgrQ
eU2VSXfOUj+GWNEQGglawISG/QtejF7+hixk6wU/YSuuYyl/uacBLLMhuLgonpF5
vIwv6jGsdXj9/BpTJcFy0pSw82+hhL/GtwS232cGmbMKEpmtySxGNxSSl6aSvZSi
QtaUJiNm56Rfe3ezeJy9ulQtZRv4oo0CRJIKfygv2761ps1k1HKBXx2W9FLt+8K8
DNn43NMM+8j+OEirTUkcjDCPvsDwBQ73JtvJhN9GrxLz+2644coD0iyhXJmn4BR5
w81CPLe8ClTTGCxKb51IOOc1CPdCduV7kacrvfwV/aW0TH4cwq3rZwviA5vsEi64
Ysj6sMakDG9Z0fUSJ3uLpKhLbPnQo/nF01JD6vJMT55u4rl8TzZg9W+zRvCJB7dB
6c7E+92mAGZLVVbIL2XrXqvIdIMlVhKDss4SiNcnk4nt5o+V5xlR4OwIkHbqXR/o
0TbWnan50lwy9H//0sjBxKevc9aJfxZy+GF8ddFOu+kyvfeE87FP5KsBDsssLBfB
A/MtSGSWXyH4p0iBkrqSEq2pzVIJBNCgm3mnrHekK0XnnNQzFYb58ulE52uKWkbG
PIAjCLzVMmuKST15HTNZGBaR1kNYV71Av9rkSZvrygEoYucOxibzNlvfx5TOIcsh
wu95Vr5OnJKGnpMKTWbQX8dxYKLmY6Eix2mIji9B0him0xVheYkfz053kt/yo6Ld
nYkVBp3utbARv2SVJaZo/4hp2iPQHFYBjLl3GRvNLyBQVZtnaBAvjRKaNoX2AB+r
ig9kCH4h9Zg26sd7cW4u6+9Ikj3R0WqIHlo36cCZ+kcr/riB/rBiJmusovv+mzeQ
dqrTINkKWOwrkfAXG1O0orui9mKCD67OcqSEyWBMEUJVSIjVeDXCcaUMh5pQO4mk
txwfbIPD9bSlJtnDMZqk23XJhsnbDc9JpwwoYvZgEfSqsBPJEIvp/XVw30C2nd1u
mRiqeDuCWQ+4aTwAe5mMhjgADUefea6jngQbeZNYZXMpfKFtgKmeHrQcorNvtN6q
o0P1mVJGHtb/DTWz8hLLLBIEkq/v6kpz0Y6CFiMElMg7tieT+7hhWd8gxKqhL+Z+
X9IZn5mjyrKq8wIt/oswmOHu1JnkroLT2eJ7SD3ZmdWjMhYC+Ik+k7YO6sI1Z0Pe
LMvuhMoBXPyNhZwGMpc+zlYKNvpK5RAD7ReTeNgNEPqD6XCYjSqIjqpRMODc+nY3
MVPwwfgl2g7Byl/d7xV2H7f9YUjKG2eL8vYyS5lTeCqlZyrjFs8poPBS//c5vXQQ
X0fpV0sTWWPJNW63xqSkrdvdbpbBes5zrmSDY+bXQ7UmQ8L+YTpV8kzaJYjKqaBO
Y+a0wrdKOJU6bvCZgVx8emWEIdtoNHCpsUq4UGhgZJi+Ztq3nWn7u6civjVRq0oZ
o9ZUehB9CCtkNfGuSfKljoW6g0sTP+7C9pLXx4kYkHY33tvfHTuxPHaTUYRvpQ6h
CH1abkhe3XqrC8j//NroLXPIhJJK2VMRDppMhcIQbfZ8sFSP0tai8Ut7eCJ8A8Ap
EvfwZIxMwuE/Dd4xdWvwR8fuZaT3MUtI09hxEQdzyZ+ArrMROcriymh/xhC5V4ne
12g3kQyHdPNKXaWtqxrjnApd+g3ooNzKOme9jL2lteBLkjqjc/s55Ad4/BtA0keg
Oqf3pKtYe0lmQ8KFO7AZPRjxS1sdLf+SNqQFyRoTkrCzzMXiararOrBA0pngGZZT
GbWRtkatLnP8KaUDvabHUejVy+OVKyFV1jP5TB27K/TaVdPE1S1LFKYQ25ekN0t1
1/b+CP892NYU4fl/5jR6jOgbYTO5kfhOsJObI7lkrznoAhbj2HhF4ZmnuPJlpQ5u
Tk0aS9TcXVNRAR2BBYy6hr0aPfPhSWXR84BQGBlmYs6Y4F5sTRarMN1oxamerBoR
KuM+SEuG39zjf42GsSHSU/kskHXHrXKGTF8gbiMHmiYBXrXIrDti9UPMi0mr6Z/9
goEfbsum4Wla7m33LocYbQ0VjR2xpYzPYR9kQviFfwQgsy6LZAFQS5TxBt0/4KEg
RHO2mEqJdO+/0mhuZb64hb3/tJF4gRPvGV46hzMM2cGs+OY9xaoApP4oGA4vm+q9
0lpQWb6qjSGK9mZ2rZYgPc0YFc5tIiMHE3+SNxmrMxQ8kELLFFgC3jd5IO/XNdlk
as691y97KmLgcScSeS1IDSPHsXp8mnrz0kD+mWiQxCbnw81IQ7f40TNBTRjWyPHV
IuEdTERMb66WUJIB1y52z2D2XxoQPuHVOVtotYc65RUGVVcKfLKN0SxQQH5kiq18
wiR3jCbPIY9Vl06ad9NciMP+QY1jRx6+iX4rrds6rOe0LQ4NAE76NPQh/ko52QfR
zXoLERBdfeWADh6k2hJ8UK5cFPJ062wPEs0SnjepjE8Tm7NSCpUzvjlIwPmkvaS9
h08w0WIRglQRSMpB8IkKGsRqs/PXT3J2uUE7/ZixxV2NxqmwMab9eOLOiwhQO37C
k5MQymTj/Tr/Lzn0cNeIVNIdpMW+78sg7HCZ+kIq60S4GE/78q0qrnH6VgJWdCiI
P+rjv0mPlez1AIKb2hP7Iij6/0wpr6b4PguarEofiDRYp2Ir98r8QSJG3WDe3+KQ
Bb8NTGKb+dTsaC0M5oJw/X6gyctsxOliYzRF32N0BHM+ae+jykNxlR/eYeAoVw1N
4cZRnWzyHPPnZAJtH2O26Ug1M2QvqTtYyDtQmUDs3Mmg8NAFd8i+sEnzBQOkbqKw
d9YBho0PhcPA9PFLpZMEHbUu6OLTSyLPV7aKEPje1xjxtEWaX81x6mpzWIRM0/LA
9AUAYndNpO9ftN8fmQZG6fniHRSzPTTUHyPFrqgKzolqMHJT3QmocloMVTezx4Ln
ak3ZrEyQ0imF2B0KckAk+2TtsRCnsrYZXpQAcv1IrSFYb9mFxoZgSAjnyM+0ELFE
yzChd7OMML97Mq6v7U/CfhFxWjhJ1W8I8G567p91Z8c2yrmFasHWTQyJf6Bse2Jl
vWxrlZS3RqiwBteSTMqgE3ZonQCtmJXONj1Ca7JgAybFjtXO6KjD0gu3IaO0u8as
d/+1x6yyXknsk//BiQceLqMwUp3Q7s7Jjxiu6gDz6Fe3Xq1PmbWFzh43bltqOJKm
EUqafL8tDRp31ZVdEpXg9U8jZwMzkamgX2vtVnT8rNjeq+lyzWibeFbm3s1mDkc6
9JnxAn8hJh4qFEJ8pVStbvswTx0HMEQFNzTkZDsHDTw3jVUMAOLWVUGhreArnwVv
e9te03+9NNa+T1eb5hk1ExK1Eq3zRk4ecxPAUy9c6Bj3CNQHNcTY36E19ZDHZM74
beRP3ZZmVYT9nPp6mW0AnAnNvuTQJQrlUWD0ILvx15+ljeLviU+lLxCualVus1/K
iQK/mnIvFwDYgy6L85fFRUIQuYxss/4K8IZUMXqGYVlCeFSMrVqJWnfagPZ9z1EZ
9d8nNpVhXAWkkfXNFrIOzHdPvjEY2Cx7t5dOtVneEBQ0KCRTgW/qD2P97nRyDlFn
u7ym6AEPyRTOTLGa+oQBieBqMRR2FQTN5CpQqQwrdNZqFYJic0SqXfZvgUlDOO2r
wi+8KGqk6pq+D8R1Fhptf53/NtYuuGrEaBjS+56xXj7tw3bHfRMgjotNq7qqrStv
jfLkt8owcS1TXwC0715YYal74lQNCCwohHhi/nrN9wbx4yb6jU8BJVOhK9Jc7nEx
qU2NRgECEM/bbPuxsOMVyF3nxD+U3XVI9Cz6NrHPzoVxQCj4ykXZfAOUBIZeV+3H
cuop6KVObmh+zhLJiYAnOqV7w2XK0AmKl4QpHSpYnTknynMY4XEkTxZRJJIuK/gb
vG3RAssPI6cYxLxJRJX0PKdVmFYfQaTULF9P+HXacRA2dfbptaOEEvI0lNzv72hL
EkX+W275gFVyerP+dHloaFvRqzqbr30ZyC79iMjW9mpiX0DxIoxpvRH8TkPMdgCA
hraBXyZYzW+w6yAQ/LjlQL80Y/QrNmjbZhEFaBeoVKLsp7RxTTYF0sY5xH2JpBQS
5o2BWfv9QlNwZPQUT1b5RmPGwgm/0y/7lHruQvHJIGsyYf8CLnAzJafsEjPGxCC1
jV3ushCYn8f9xc50YYozLI1hGg+nt0pLs6NnDurIcj0yvwq9Xwqlv06I5G0H+1dY
dsLvseEl+pquIyJwKiUe/jQUTMiajy4EKZPKp7N+dtW87I0k/UpYVbrppUggMBFm
XrItflfZ55NvG49N7R2l4zzTHtysdL28XNGp+sYimg6e2jIFxn1Kx42kw8V+G/7F
szAJf9vGqbrguLQRpr9y/J0A9EMCKQwDGQqyQ5KxAO0I4muMnGBnhK7IS5gSNBne
GfMxG58bLJA+HPaqm29ii//bE9JbeEe0nsBoWNH9BIQWz8uwksHos32Mf5ynJQ+U
Bf5CXESDB/wJiSDgGko9TvOXbtfeFSCb5tDl/KXC5TkVzwoXh52EcFHMPbXWgPiy
BEKTw44qTpIfZV2MIzs4Tt2cXoSFE+wjxHQ0yS4YUIp6HrXwlkg44kWKLUG1SEcx
tMo6eCVe+0gEfihAuUudyvG9Z3rklqjOSyhW8wisWaY+okLlScKfi8jaaFnzyzEM
OzPlPJIN2/tcyWW74wT+IzqxaqDnMXBCg7n2eg3ZhZm4LQkC10whRBopmE9Ptb0w
8GSxXCk1cPQM0du2uJMPmoB9fBwUcaqBC1BMb0nogH8fBGRr10HzZ/IW6srj52Iq
u0BQ5sm/f60w2YrlPxoxrVFaWYILEQkZJ0k2bHepbyZIG7TLO8dUzGTKlkb8Ej6x
IxhkRJg1DwZmRr/+nFalgGEmQH33k2LAimOdbHcH2tR8N5INJwRaxO0G6SKc2lTt
EpcyjoWefiGEg5Td7NYiJTl7HWx6br0DVYRo5XvfWxJujhU3WVXrinL8gymG56Ae
eqInaa4S3Zh27b68BQoy/lU6xqrIVZ31oPetla9XPr6iHXE2obgGrzWWPuygblrW
K1fqpzGoqlszum8ZV+AfBZhNcQy4BPL6M9tNDEedGSFXZJrmcNjW+9mR9e8wpjv9
zTHs/bkXci/uhcAIfijP+JJGc/1XQuywLJA3eG2VsCC87lX8dWkEgQleQdWedIir
4P53Tct6BiVAAH6LO/QXBO8E+SOv2KTallLtoBugcDhEpL+AhVwfG1TvingJhe2t
ET+XcslqHdrrr+ODsto29zVSvCJZYmEnTTxYPM3vFb3hRkMyf/U9ovkB9l7CaKFv
TwtVwMuWYFMkwtPdtUvbPIlEj7sMHoHECh/oaDJDYbhu4Xp17rMJjPl6Yzi6qLO7
RBDJn8pTU+AZDthgVPLmtCpACcf0NwJmGcF5UIbGJZ6NBx/Veye4zOeIK/xmIq3d
BSLdM3goUsGfyGA1HkDZhjzfsG14mmC0+TZAehDsUogXoS6tpVOVxoeaHE5R7YOP
KDjp76yAp3fCqhLl+Tq/cVxjBEEBc+dBBPucHQlewuejf85diCmwXhkrQabKiO6U
jQgTpFLZQu565jsvyzZHZzX0HYIX2HLEetAjOvFg2Gd0uWLFQGUkOeKI8EK1uXkE
vwvMNnBdiLNxEQD1q4Qa9UET83IVwdfsEqUTEXcl6uFIBozEPGzT4HauSXaioE/4
Ojponwg4HaFbpienaa7VhMO8CkzZroKIUGv4+Y32URtN+fM2/FBJ1CiTUblZ1Enj
uxMFyptUZKppxBxfhn8iTG8EwM3JYB6fUMXubw33+itMD92XHAhcjaLwgJid/beF
eU8UWaqQDETheJ8xsBhl+SFhM6knLqsrfhGQToSdGhsmZ3WPI8w3o5GHvxfo98he
xE3beG+MajQkzyBHGifBwxcgo7NrfwD3c3ZVOLM9m+DjsCjE00A39agZytzTIaLF
ZvuGuqEfam+wytUBhAqZQyiBaxvqBIrfcTh0ySs3UVDKX2KT/7/EBT+/oukKtEWt
/dRFkLmKESGZaT5DNX7usd7ZOIey1EVhrL2ufR32+qN+IknUORxuJWFgC/WKC2kR
hM/2dx7z7fpKkF/j+73IW08SqlIBF6uF/N8DEKUgvqjrWCBBA2ZxRi0Xj+I5zXfJ
9SE6mX+KIMIf3MnJO5cJgzGplrHK9ZkazZJE2D7O6FfxGu/k6rOAGDzjJDs837bz
Jjxa9NuTB+9wnUfiRibYq5OkY6slttv172gq7Ycut4ycmK6OIWx2ouCEauh2xshr
4HIeErT12/mSh0JGuk3C2NyADFXm9sy+7bDTKrefWyhXIZreO4FQZeRjw603mNpS
XNlnFcGpjhu//sEbsPjE6h4/SbehWiVHcC5GVZJ7cPNm6AasYybQDAh8rUDpswmN
k+qUEm9rMn6idmO6wMJzGeGy2J6xE9C038yUKbWTItBblYU6H2KfA9CVzigNbAqM
FodTmRcSAaKfMnxH3sk33a60ZKernb7DCcWNUreXvDy8i7sdgdZheAuOCoeLYzDq
MT22kdjJNmhck3jYLS8+lvWsJizfDPSY2pNOfbd6XAHQotcnsBd2dHBICAVzkw0W
cciQSF0DSro99C1ptU63obabeX9BuurN/18tlnmXQNJJAv7uP2L9mZrtZZwL/d01
6lfqk9i3P6l0NqpQLN44Vm8GaBqCP0tP+rh/qgthKvJi3glyhOMh8rI6+AfsGwIG
efKLTMyGGjgmhPVVPSMzWjUUSN379AuXukIGuQi+Kh9r1wTJISo3ioecCCJMXTPY
MDrrxotNCsimfKCEXbzRLJT6bhR+6/MRh9Hn9rzZDUWcXG7KZFDPKWkk/YDKERcv
BomqArDcCV4Sqy4wxAMZyU0nHGChBwNrmzb4XKWs97v2AVAv8Oqt1vuzg9dzzXGp
6U6VgtIjpiJgyQ1Zksgm5gca59qoGm6eRhBcXoWhEnoGhJi6CoBqIXFQdFB8Ow3h
9DjObBVWKGilgSvOhCElIBbt1T8tEu3g11cZafAxDF99j0gc2QDqMSTGYvFr9vZ1
f0Np6oiUsreqgcMeZ8/YQiHpS3ozhj3uWplyAh9tIKkSZTn8cRJsbUajLVa27iR/
Z6hTiRVbH41YlusmKdqekqYvI4VlncW8O+Wxvbh9oMTP1T8KVSCAMYWR88p3Ib5s
YIsLza3xk/VS3nz4cdVAVTR+VmiFvCLPD03Lv+s3R5uchAZgAg2GZgFFMGpAqQnM
bsCu4CcHhZd5/130nu2VDu4HDciefJEVjkZBpAUwgihwJEBYuuZIxZuWZS8vVT7/
lObEDy72iEZ6v07gEhokauMQMOWSNzzlrJL5noxK3DbHuDzmIY5FvcSIheSCVyvf
yWc9L4X/MK3ZcW+4kBqIG95kFqSJcPLnwDa1gw1Nfg2GkW6sDWqEi3GmG6wAzQUj
5JG1zXB7lNilry7tx1tl9uDYX+kY4RXyV0hSDxp1F1XlrcJ3hWRlRXVysN6i65+1
AHYbHAyGIWIA0peoYNV+nlijQIL8Rajffmwnb5iHgz4R487S779QhwCTFI78GBUy
yu7Xv2XJCV8wBQtjYTig5+Yi36zHwBYs9kXdp21Ybfyt1a1FQK1gxp583BYlrMcx
qni5Bt383WpXTqWTpj1WnrCe6f7y48F3p/UcYO0/AqO2MKS5UcHNbn58+szNd1LM
QIrBSL7YNxtBr1OVOuQhx9nc4qn6b5Wb6NHuTRanGYu02AhxOp64ji8ib2WDNJnw
yoXHBl4cYeg6ccPDt3nv58sifreJy+zHz/aK0KsaPU3DVaF08mkEPYlU7wEUa/Ls
OJYhnOEJ1maGub5GqvNnM3KEwvtjDk+O0wSJI69icUv8vr64To7BeEUzkryQpVU2
guWSmGFqBjwe071pNiXBmZygLxT7b+sekVRFJWQcasGOb8+oZ+/w+T9J0bxOBUoy
bv5S1Yf1XwyKIYJ0uRs9nwwT3sG5p/us9V+6lyZBq5M2syJGwgLwD7bckcidi+t2
eGQ0MVluN3ID90iWv9sBwHSHvQOrWcVCD1ZoH+Gla9SIVSr0c3wkgF57tmqq8pcX
X9tJilpV2N214FNqT1Vilsd3ePK2hyxpipVHZ1Vn4AtifPHij1IW0HjkwHgZXr8y
8oiahWMw+vS2OTl2zMT2OSOZWBocZ/10quiHlXHbOHJJaKEUBf3idXMN8BPyFL0a
yxPh/cCUj6Pl8+trmJfi7tA/T+iGKhmdHHxlY8+MblYjynigL9Yg4G0p5oDJsidH
uUHIBnEejWet6GoPuUpQIFYKTcLsQuaOa5vrOps4g+yJZOPpeuDxYUjhjB0ovSTf
Y9xf+SF6qX47xiGPbA2p2G1Y/Sr1nfQLGAnMEk0EVrmWj+KtkimtMpFA2XXFYZ+w
0+7+s1FAbeFQ5iBsK4UaGYr83v6b9Ywp1HaKYYrEvNp/AD3Mee/zlTfznx4N0nwV
XsxcmIm/TAoH3U/q8/d3tD13p+GsCZgtr0KzVFIVunYtxrYh7z8gkuSXUYILzgPj
YARdIEMsUaC9gnP39VMSPjHnSJn4qz1vk11Gxy8Rx//4IFU44C0aUuAAAu9qwdqD
Tgs2hySosLKUL1IOgPrp73VtFRLybiFRf9cQEq5KPy9Ydzqlg2MVVmj1li98U6JW
dLfpKJLXFq83Npdrk70oELLFYmtZ1p02ELOksORQJh3svZa7XgeLOvcRxnQ3/Nje
tevfb9h0UY1gpUfVKmis7KVe8PQlJ6HciuFBiI5lXT6iIzVvdFwVFytTspOuFbeI
LmASjxD8+8X98duLJIBJQOknNehs5+Ru7Pq9GhnNiUx+MFmjoUHcZem2PlIy4zTt
Go6nEnf2A7N5igm3D+2im8iY39uqRCQX1otWXIEcaxo6NvuGBRkrhCcWDi1dd3dZ
h9aVZu1y6ij2KGU3dqsMui/3mGGckE0UNXB0uiBYexCe9RsVcd5TsAR6wn0Zjl+y
1xj8nVdjDJJK0NpJY52ewv0nOtPKsOQDb4i/clLAr097BnoEdaqW7RxaVV0e+yGA
e+rXrbvjHly3wbv0MJ37MbhCq+5zhCn88FS3JgrrhSY2lf+QzWG1VmYvbwmstkX7
7BVV20z4ELDi77y90ByUahZYGYSCDsA0niUe+3X7miakjNYCCj6587NfxgPCjQ+d
k1K4gXIJn041a7SJv/1YDPYECJIAWG1hTzJXO5/kie5KBpV1Dj4cf5Rdb/lYaS9w
N8+uDsGFBSSBYS325YdmLYkH+gGGwhRZYRRyxzsVQwOd2JALqa0cS+VK1Yy2MwKQ
PvRsZx//Uqd9wP5588PmxGd5nI0BEIF7faqNxkiS+vBFOn+Z2cRCbbk8xRSO2gnp
S072SJwssF6A9083I4M4RQ8QVYkRsXbuzJxqTuMtFfGL1jIwgyKZUUAlJYehdaCr
eS3XSjKEHTqHx8UZnNcDjWKLy1NwfFNkzHLbyzcSpI4qtq4ovHBUNuU25H095Rin
F6e6/Ikp7IdBj37lcvWW/A8IwckUOj1JtA2jwtF/iXlQonBIr5bNRWYF6hdESuqc
DcAzgYdujzLbM66p8xkWdrlfLWvQScFXc9T6tRJrrhhN+vFdj+HBmW4EOZfcndyb
Y8eY79kG8QfikrgwioGwPdnDZXv7DiLxUDFKX9rhdtgn/4NBUhGQrSII1CXPstPl
1VSycYDyuGjesepDz/4m4zDwtil003GFuIwRiXaXTOKJYu5E+OnPKc0+euD3MkIX
NOhpuDMM9qQ4/SjzkiUohf8xSXUMwlkGNng3+LsA0Dk8m+W3T3LQFSmS72XLzgIv
YiQ7t30iDRx7+GWpUKn9aBkaLmAyTsPFcSwS8jPoC7s9EhwI0RvgfbEocbXuE67Q
wlV7E9sRXWQ1xmQ9cpxngJXURHccHwZ+GyHxOKJFmOOT8nLvan2uCZNLMW6x1OP6
BRj8qjcOQgrx+q1oOIrFhHnFCtBDWx91CXIIBWWLa28I/IOirLW/zyWj8eodWVW1
Rtfs+oEBpdMezp3xtz3MWgjkaKNewEjO9UmDykE9SxX67fy+2KI9JYk+06J2bIJq
g3arCN5sRBPApezB2RlqKI4KFAw3UR9ZyDVTVmvLFc5t+qqILiKe8Mmkuxw49E2g
gft5qcpr4XUXPd4W158IJttNOhSASYYc15vw5nvVTIKV81wgHx/1JYy03u27Lyi7
/unpeqbwud7LAKm/xG4XDULTHW2k740eEz3nt/mBSdIcBX4igXQvS73D/MHAMlOg
ZIdJ9Jt4NZAEJVGBzuN5oS6uaSO1d4g2Lf8zu352Ij/sWXIiLIGTgouzfenN839S
LdDO7h/H32vKNFnyeG/nqcwn9JczHCMUY3AXE0FtHzRRVxPEnZ1NJtmOJOo/yOYM
5uzbAzWu8ttWlAJroMq2djhNkstKx/O5iuLysK7/7ClI2NXPpLFARrnEyDSboUX9
qc3M/6+VytBlsvQGdAwkqsdr8zH4vZTWQm8QZTQEodqD/7bVUvYwPC91H5guNPzU
hPbThdbMGsxYdP+wnRIDHsrj/VeOKEVuMScPhenJdC61UOYp7UZaxcxN+Dw5PjkZ
pYbtSIWRHo/XFeHOl2/aEDrzEV82k74TFg7VnHuNaStlWyT4efPiUVA05FkJE0lQ
23onZ08XE8YdfZWqBzKd7/6iZ8u051Cop7jO36G2jEUF/K5ZLfm+LLuPbxIZ45q0
Rj+pnzbjuzDseGKVu8Hev7s7TVmcqdxMPbFai/9xRLJ8OXUG42+JIC/hBOGmjjYJ
TVXlon4952al4gFNSFWrTHDpQb0lPfMQ/QS/9kcZk1J699bFNhqe5n7SLmRjN6I8
LnZWP4wKisSibwRZmSqjXU2WQwTnqAzwjqhDlrStjboxlbD3RvyzoOpoucHiplZD
50jGNyeTLeeIAB3aFi/b8YVlhj1vz8voaA3g2sn9VhpOjTxZ1wBWRKUI4Tm2eYxq
NmuNJXOgyog5KxE/nujMpr2Eh3ZkGknuk4VXhqw9JLMjeR6Y5NY02RWqZsA/rGTY
+eTYx73HUwa0pwkzELuWIBC6xbqtkC8L9pIUb+dH+ulyFk1HzEH2ojELRkO6kceh
7S56n78x046dz4WwQJqbP0pH8pOeBWdqf681JRl3JZdviNbZFGYFHJ748aI6VQdn
wTMgWsrsPMmH9UGjZrzEBDQY0O16bjHkYdIo3NoHt1hcF4FIpLqQyWOhbtavY6y2
DfDj2flS7vbHYTllnWa7UckbWmxxDXZffqIvoRsTS9BYx8SY+PFXzQfdQawbk5OD
ObjhriL6P7F0BiCppx9inNyxivniExw6KB5NjfwAueS1IvMSCgApSGxDaRDy8z8f
Hp9Kr7scj38g7IGVX0YMjIDMBIFaCYwXxC83v6vYGVIYXZqu9nfPUlJjqhnW1h/3
xKNrH+MQ0OyN4FKUrFsAckXVZuDHo0vGNxZmbJTg+fIV759K/fYjdezpdL6u8IJ3
TNLwhOvGv+VaZF3vo+NwwLa4UNJq2rUKf3U/wgitxotWeRv6HGEmaK8vYkBvO3Nl
vU4jkbvkVCR8WalO9/A6bRa/VUi0v/pS1Os3jO4fw/0CnrMrsrahv5tzMJ7jp88Q
SZ1UGBxPDYjG3XwUNFraSKsj6XJkRFEjxwxE//9HSaZKlEC8YPRTaVmxhRJCPWjV
AyRgg4TnfReRRDHdHTC4IupHOQjYp2c+BkGcxNGTBnzJUnYX8b9LyOrw83WFmVJv
LoZkyE+BS6kMc0YiCW0/V3kgiueNeM8WNKQmvbTINhcjTCAmxbpAbJlF7dsglIIC
caQyez2S+5Qpnwo4ZcmeV1ugVuwKR+lB1C3/jtBGgZhpWvlQKP3ABYKCYgTxxtJ9
M19W2QfXvwPpIevsZ3AOSonc/3X3IJdCBJc2XVLG06PeA9B96EBUFMQyy4wsmv9D
XBnH9mUcs5HMSgFtMPJGjYvyZ/PwFvuRIXoCBsrZEy0udZsNNXZbTaZI3KuIT4eC
Yc3w0lw+GucHOMViHVtEO4rApI/MuGw1W8ZdHBbF91dnp8CPn+vR0m+zvsBKZN1C
D2Ktl0LFwiA1M1j901hKusNSwHRaYWcvHOfLIQnpUWqKVqwPI3WEysZ174dwDdCK
rHZ2LTyQwG4FTFScrFOwOazBOKBIBqZ8Yv9M5HiAQDR5DWBl1Urri2KBPwVCc/Eg
QOu8qChaWNqRHh9s82vQqGEQh2JAmDF+OiGcFlsINviaCBnl9E5DtgZGt32o6oz2
+EkTaeQ1EbKdYOspwxVNCSMyRqEpdhIQrmXlJAljtlIGUZs308s6rf36vhnZVfka
siAOkKXU/eu3YPOOWU6W0N7s/pUPFB6t6P+zS7H0PSEkyGmnvszmwzTUsGAyGocR
yRQwyx+2m399ssyMmXoNuPjqr9sNRfRn+yV8go0movCF97aIJsqUM16XKDGmgri+
BtpZzzXGGuzILOpY6uMnluVJ6raddnOu5NieLyiI3JsmwEmHE2L3BKe9BQY2d7mE
FKorirQmcLvEBiMbEHHYPi636nyi/WNlmQX2lgpdtUnyWzNKxY+Y9KNEtbLX84zF
0cLfqzFgIxikght1tuJQgK3fQiXNnduc/ptcd5HffHYWu+T+3LnbyGy8Rvl0Vot8
Hhe/GEfQxL2KBZXOMzT27AHQSFT3fJ4b//6mdUjAhQ+NW7vcgSYc1KxbQqWtaybK
erMHnMbsRVJ+mN6p96tq8l4jRlMnqaEWFtmH2aCYsadgRZf4nsH5P8LJkgDJ8wz3
hytRT66jRAJBWZY34sPDgkDyx9IDt0isFgcf8BvZ0/vvh5imhXa7ddAo/n4VOPhC
z/CjMHqrEwawx/WX+1ay7hi2pSf3jayDycRRZYjmCoPBY/sk+n4S27w58LYzcTYZ
FA6XtQkDW0kqyo7m9/uwkaVaNeB502dVePGUjlmRkQ4Im1NWJKOnjF/kEkcy744o
vBjtgRABvM18tqtHRwy+lWfETBXuHzuNz1LVLawzMQ/B1sGMrgD3gyOX3H2UjaV0
8gxJiDSYHkuwkQluw3wr0RXi2dPaIzZuDPGH9CyRwC249OqloQDRY/uYQbhtmGWY
WIZLWE7WxiXdSsaZyrs0rRtxFWEF88vC4iHqqyfXrb818z4yNMo7OxW5yHKQPEN5
23phmCo2CNuOJMXpZtzIlN9EhEc7sD9yE2rEcuK+uofSzg6v3QFD5bfJck0IwWzD
+VnZaOZtID2NkmkGFUxyzgwHwD0uiF5Zd0056tSd2Px2fdZNb+HgckQIGJALxtTJ
cAz7rzb1pHt9SK/EvwTQIOb5BdTLNC5mz4m2WbPHdCcw6IAPQwANjaf3e+TQewcY
TrsZIinVa2dOiKnn4vi5gnAq0gOe1JUIKuXKb24wLmG+3I6EKgkimhfX4I00n3pA
YvJRxNIM8Jo4htWmWZidcCjm8mU9t0IOexQ6PGEnlszDDgiMo9cHy37P3Uxdi/RY
4M9g3Rn4p7qcbmbPqvEFgxFyy/WTjna7y/6EDIpWrv6wqmru5WChmbWcp0NhA/Bn
AiKW5zU8tuKeZdToi1PRyze52Mnmfulv07tU/MCg8CHmgX+sH50JCOaKincpu7pw
LCpEKhQtx910QowykR1rReqZ1FRUSpWRB59UoeBFd+XcXO/Ga7QNf5nrRq08EfzS
vPp/0shkyFon+ZuPv1s3tJ5ioo9J7nfrCbMIrfcIwCzUDbDT2FBESEi4/UwPuxZF
MKKYgpcTw2cB4d1CQ6Xss5QxGUIuore5+9BHhs32iUuezBto2gXeStPWp0JT3/tf
GLriRA0mKak/+W26coARcCOFjTCEwcNH3S4ytNcfEBtDecH5tUZUH/kcJfNlwwnI
Efxmo2zkgnXzHmmvepJeOQMydEOm2FajaZ0T3L6Sd1fQ+B1toK18DeCCPm+2kRBt
wbrInorSUVGJjwVF0fLaDof2gybgf5Vjtr+yosjbpqJx9sjEBrrI1jCQl0vqpyMA
p6cxN5N95T85bO67VmpQaTesnXeq2X074n58HkzoPGb70fB4fom8QygkG7L2bGUI
Roixg5FAAHni6WCY1z6ndxskKdWUeSuG1BIIAhs494XbEZg8EAf8/QgxaiYLQie4
uD6r4QUoRVPOwysqv5QJ/V8KXWwSKw2eJyKV4pbIVJ5D4sZSGFMbsC93dSWmRCi7
OsajFG08TnG/qTcukjk0L7WKUGvDMSFHXM2OKRSkTatJmGNeCFNkEssOB8lSqvrn
TV4P2zU22X2XeiC2tD16IZ+qgzmp2KRKmzgL33MTjZ+e1sWKQzQWAX8CsqrfdhbD
i6pciX+SP+qkfu980SEGLBCFeofh3CiqhxNKNWgnc1qI4OyA41Lm/MvtJyoNV3SY
NPLpZ5MP189y/0lLZiccwUeGEqMyqMCXgo5ucMg619H/1EnKyGWjogqP72WE0qHP
1fJ17gHHyG2zqEVd/8cuI60no459UaG78LicS4jtKFggtReoyJGhKWgCFm9ePndt
N+PMOQtP3bP4D9Tv3qIdo05kP8zodUVF2z86OFAzOobFGZ6TW9x0OvE/jqFca6jm
W2rCsfcxfCgkq1kG+5GKhlCWcooVq5AGOVSj8GCMLIDcIxjg9NaYiqhpey++U2lO
AH6y08FzEdfNIDeNDi3g9yEVcXeCCRBNiwrUK7KtPOFUYQNIgMV7JlllVMTF4Q7C
Q/dRmzein/r0jF+X4XOx3Vpn6kcu8AEAFQfYDHWJsV4l9wfrIwU5kbax12eU1GQ4
wHvjZDnQ44BSPYeRtKdP86188DGAGfkYho7XHEzJb06MnT2t5G/GzB2xh5FHdNkJ
AyWH0wYMlsYB6/HGZhSqlIROO1GDrEwpGPaFVRwBfachEaNuZbCsjGZ5Nd01Fdkq
4isheYkaZOXo0iaKvG10QizTZIgEALz364SzKxGs4yNKkBSEB0HpH+ZB6C6Rkod0
M48wDIVFRF6wt3hlIXSIkE4Q7rtTWdarc4bll94x4LpMtSnBdmizPvwJ/YDhNZ2t
UFfzbWVcxJ3tqqv3MlPOBkGYppnaO0hbEh1G41vB9ZTc+7Hp8j06bRn+3U9R4nUF
9wWkplTrmu+YSUuQT8BmIBw62xHRtrKyihyzxmVzdnh35RFjlITxjNJmfYkKmtCF
BbmgwBvlK5ALF6tk9LwZ2OFaN49srolAKCPuQatVcvGv8M4fle+Adtj3GPbc9S3U
bQI+Ex9xCPFa7CmA+B2jyE+gZB/KRp+uEg0/xC4o0Bf7Jfiy3ld2ek7P1bvPKHpM
Cy0Oh4Ufqk0Pl+eeMxBPq/zfDttOP613PuqlBvgEoP9e8bK2og2xyWez7yNP/vp+
4PzF7QjVEEqvtEmO8NJOixfCFXiBJV6jjVBnkD2uEfabU+6804ITYCx7S4MQxUbi
kAoU/xf6hNaJqPAECfgLkPeQ+RGG6ikfDrPOWLjPwhqFWGLVva9ZuuBpeyO7L9w6
6A//4JABck11VWKuw/Rsfr9YMa8are166sWbvzSiAAFJN7F/mI6ijbBqxL5a2O/o
aoz9R5F/tvZec/ZYZ/Z5NP6y95QMGWBpS30CTVo7jsGZyWmFZjTlm/YLZ0SNg0b+
OKS6AJyser9tXDZdKAql/3xF+rdCh2w5Pli9rxJel5zwqVd7EC2qbiRKZ8jvRUZt
Xildpkx1eq4upmmVuYjcuz1SqD9ANUfI7Hckjr4/Lw6QVxccg/w47yw4MXTFNl1x
tPJQESA1x1Rk7nBYOSpviFDxRNGASwcIz8rPoS/deopJyriKO4rMr2jnKY51Lwjg
+j+QrAVjF6Z0ASbekFtgM51Fmv9EE5juuwCFT/WsMrP1DFOxj29zq0aiVCR2lRoA
1zNhMQjpaHK4mQReWLIlo4lxWxHuvU2Ft9oWyJ849iK2T1fTkq95iJxackBlJQMc
oe2ZFoOhfLgXOO53iQZj+L5KGuK9tskHWppxgzfzKJ/zFnAIxZusNTdmlktNlA3m
p2Gu4Z61HMSYxnJrPI31JgKMV+x5HxvAKZk4QDM4PsPSpyw+Zoml3/5Cb3m9rt8e
5PV+CqoVkMWNWHVnCEHM+e1WW1bCubMD63NWbwpMebuCpT7BIE2KfzM7BvdIQSsb
T+r4L5h8aGt9Y+qA8upoooNvqx4m6QSV3JXmxPU/3uKL1hdnqoKHimvQS1ikQH04
+b4tUmAYWM+fbJNesi8k2rl37C35dWsXmfS0NxRnVNPSfEwH8HD8KcclXd3IAdAP
iTK2x3W/ihFGDZ5pjtJL/MrHmN5z3VH/pG9v+xSJczvEdVpCkvY7T4YsO4qVg3Kc
CVCL+yANrM3CkjANbfwHhjuDb9+HktLr+iLl3TLfPsY0NAHlsJn7BNuMxAoDCkex
4uCJo7hww81e+OHaP9hYsXwpEevM92K3x0Ji1OYHFTENYDWMXVHAyoahGgFJ3q7H
QLTY4jxWNd1epWmVkQv0nrjmamzBQ80a4gaQAfvV1lgly9m2INyMPQcjrGQSdGjE
XNV4N1treS+SQ5baLb6leg3DLYQXsYc5CWf1ubvX55GvGKoXbXHgrIgOi9bozv/l
j061z5ZhoeXvwddfM9F2KDBFr3ubG1psbCOcrVvl6Yzq7WMO/rbMyN/V3Xvx5YE5
mxUhZ0sJkMuGeS3BTzwKNkY094dC9+dc7ZnpZAJON61COET1gxLS+gir40P7lbA/
V+j6pEnBTd9Lbv8FtD4acApPYclvV7fH3AF2TnIov2sMbbmGefQAx4TuCJJeByW5
+p16cAcf6RSnYnOjUa9smqy4PTajYGxtRRWrsSpbwbLc+0MxUlNezumh1c4WARPY
N3vQCua2yP0uIcbJP61zhpOpblZrCEj9Q/opLaja3ai+UFTgfcceMN5Jtb29HFu7
6mq/YvhSzb7CN0usAfE6AZvJJyf9fjjSpsSW/UaCEkDAn+qSkOcc1DPK9tW2is1A
0K5M35fbkslRM8uuykUICkBlOuCHYxcL0AD6ocd6aXb2V7eoB/G6PK2Hi9vj8pvd
0hcAgXblLAboWg9J2GmVxEG/69LFzfClGIRDqAaJtgn64iAj22P3zdoOh+xJFCQA
NVj9V4t2RUbKKFuGhO+lq71dr7QLIrIWZE48qq2F0+0+XyqiRg1CGDACH8aqko8F
k9qPAFngNygdvvNQiggNdq5C+uN9OIvrqAEhQZK7DVxbYzZASKk3KJDaRUS/Mqfn
JzcsHJlqsE+JNrevN6WqEAegbIJbdN3k26sGNS6oD+Qzb9mDfI+4cWJ9NZqBzV4U
plKUzKxoI3Qn8rBCYMY3JvYTkYO23QTssbExDRpaa0szfR1PTVYFSzK+NvxWoi4X
gpOQXIZOwFa5RKJ94x85spaPkkVmsB56AiTqG+9tw8HIQ8Rf88mtFdY+qk6TLbfX
en6gN4zWed59OlVuUt/BLtaDXLHsrNWeaVk/lzhLjX79agbM9zLe3gxBDCtf8v6a
KTRsqGxBPIlHph6j33RgN94WJfdVOAqqDPnarhXl2HlbaELa+7XBqSk/G3nAOMuW
7asjkxWl6gbtRvNsWlAqVFHDPsxKxrluHcSugiM6bABjV1WqaFXTFS6aXxYWMkry
G9vgYavkF0hUA8SWOZEsVmUm9PCTTpX29oIHOqKROh7ZZvF1+7Q7WU/jE/qWeeNM
DhhZlHNruJoFRsYu+0IcRCG96PCkfKqwgZANvWq9q42i7HgVLAx2kcy+Pan1878M
YwljE/Ry2F5sW3EOtMC5tVVZ5pNvVm91o2J5/YB+hdQKvgRFMn3yUsZQlyRXaKMW
FUF+Vqm/5a51dE1UmzVKFunE07ovv07OzQowcNn5XcYj4mqbCxRT0jPLWgFZAzDu
5DJWj4iBHXyRFdUx0XFw3DEopaV06yOxZnffJHkaUO7IIWjdmyHpThL1m6ueAnW3
wiQUd+H1jpeEy0bF2FjQnD10S90nrpBOkTqTJSuzORqpM+S5DcUj6JjWEpFokSHD
q/hJL7uSHt0J9igZKv/mr8lB0SaFYTXkUWqrybm9OYzshtA+YGiQKkAzZl1rBBw4
msw1lV/Zosq42E2LNmPF5bPsxtK579ClSqTzqaV+3ziARA9CPl8gLsSWFOFK7Rf/
74zna4X3zliAWbRXkvfIyVtRBtjxYZ0if6wbXSwyOtaePi4kPRa+FbE/+0wmFhjE
INiJb1bun6RS1A21oAshMHW5KRXBlGF61LFQ/M4Bjl40cC2RIqfsaEuVZ+/BMN4D
rL/PnXqGH6IbrcRMMBKkQhG3UxEFBdnU+CZTGE1lEFgRsoUEi7YagEqowun843Tz
1bNRMerrNE3Opqp0K0oPGnor+9IfJYwM8rGSRQOE9RLHJAK/d8pXGESHHqyfCusf
TbTGJ/NvAWpJHR/ELJDGeyTmY2TXFfBR3pGEmaQW7lfBP2wKJYkWZo/Yb9PYt2jO
4FKba6T5E55sWlT3AWzesIunr51R608p9OxaNp7rFzTfYYaUwDfJyBIH3TpwkYeI
82568WuQ6ycFcBI3wvIsK7Gkv8Kenkww9ohqyA7FofdTxZs3hQYEZYbAXjSoFs4w
alXHpmdYCZks9Ez6GjmHq4hrPBwpddzt4mWDSW059ZUOyAqis+JH8Q3UBnw6vFC0
aIFAfe3TLylQM2XrLGagBHI2VLXNBtEulem735f84csSwpcngcqvN8v8Pm5a5+HW
C1XPuYqEVEqP1ubXg8l6dX9RRou9xhxgXIUuZpAxsDKj3FRXxiG8zJGdVxnCVLnd
KaMTmwdmGklSJGN/Fa957Uq7EZTNTaVLuKqtN/CXgIvF4F2rQ6rIdyRX3Nwl0yNh
/1uPLSMvicN21sHUqiLa1zP/XSep+OKRe2ov85Y+Tym8tkK/RkZJOqfkR2Pi7VXC
AVoVNJZQ4C/AiPjvRkovobhTAwp3ZdlVpBHBw5+CNNbe6BW/z9KaQt8kHxilnnLG
UMeYRBxC3G5TuzoBlM8WHxeCIgYSlt4D0s1RXYLGFf6wiVrBjWvUKwkcXewaz4c0
1Zo3nLhPTfSohRg0rstlm9VyhjFSuH90SCcUD4BdNTvso7Y10uzXfGt8Z+O2/BlV
poZTMALkynrsrS8JPcerNW78OuKyH3rKFjYizHPfp9hliFDaDoGGfHfICi68EvMS
pNvgytRsK434oYnms6gf6erZpvZkBrhS/gLCkphjqth/tY96COWKVc68l62GfMo3
hMayFJQHSxrTmpQ/2m77HV4Xx/PAGyU+bftXgp4wNZo5L6CiuKvAU+NBfqN6lk9V
xCSZzTWYdrbh1x/zJHXgupMZXbR47Gj73HXD8e/XkwHZY9F8ShcjjaRyOQG5QJRW
JobXWKcjBz8qllmYK26VfzJUxxoDPGhBbdwaOuw3WCT3m5UN/GXCbOnQ7ZQzdSCe
A2ChZY+HB00Oj0uHfs9Mg/ZyTO8JWOlJiURCSEuB73WKQtQ2Eggr616xPnDDPUTl
6oieAYLN6yuseS/ZQbocM7LCd414n01iffj4ph2lNL4WmYQyTAsPwEc6hahy07Y2
GG1xRFIbLYwJVB5MFSgAiZpDMEnrJfn8L4FlfNd/NPivU+l0Mpqcm4dzdb89MNta
l+UiHTRampu3GyHvVnir/jt1yjm/chc6P9pH3qYu2n1/sGYO1WFuNu0k+RhBY9fP
A1Mauv8Zc1kxOSl/mMTlDmeZZPLlSAFNbhiNsLC8nEiS2+X0Y1KAvqst4cpoSXxC
oEfW9fflRIDlVZ5goer5jqRVaQxCU38I9sGWZFvsfYk0zWv9p+/bxfOyio1uDW3w
cztZ56M/ie8s8Dgp9sZkSNnow9W60060f3dvercGspojJ6g38jpj6OTSdKbo0haF
LvkXEy/iZvbcvkclyMr6ZlEn/+H3CtwIWKOy+fAgVhgo7vMWkJOZa+zs/ubE9xkJ
q7I6aT3r9w2AqZ2p6iPki5Blpa5id8sBr/5XM6tN29HEVEdBKTfFJLGkoRjgbpP1
EmPv9B9II48ckfynbdhuLsWLTgE4/7gVWHBdsPPXmvA1Gy2jJ6EwuBB9KSGZl1pA
HVs7lVdxJk2TiLX8o96VJcX8rdyAHNZatWrVVxtQ2TR5kjJLBGaz3skV3D/DN8Dt
bjwXKS219p0DYue2RebSO3pEZhFSUT36tYSv7X5H6n9VgaZtiWnin1fXq8GVDdl0
fE9BxLT9W8eAaWGfgAeiEK0p1CyKbglExqKZr2SbRDKkG/WRbm7Bfxuk0BcJcpKl
wJw4Rwu6L9SbY77fNiPcj72QU1OJJsmrvzj/UXPbmtzHwlOws6iBszjGasYtoIl4
L835glvPNZ7PKqL6MQcct5QpIcsI0XgQUHqtqWb8kzaEs1C0nNE6jJI9FCqToHfN
4gbCk413A/mOOtQttDMtmE7NECHAljLt3DLMUKkPkKQEGZ5BkY75ADKOEijbBu2w
Ks+q5pbKCJBx+b8qxUis+aNLSDcrWSpZps5Cotk3Ki9F6wvIEKMF4MiKu91QMObp
VvyrWPhXfG0mx33VSw2uJq3wm+FuTNFnunUutt5omvRS7c11+FLrNSgbOKeA8/AD
4+WTaM/+MrO68m8Mji6AHYay8OSSTARc1alkwCMDRPMH3rkaFscWpXqYmjfzmaLC
o1kJv6QjB7tvleVZBBzdqPxKGFVr1letkshvW2WjDYxzmy2Ner1nTFNzOzloWwYA
OTdddHoEbvDNoGrfU79sJZXVfZ1/cM5ABcYymxq3hvsGX4TfByQ9mhukyKX/q/51
W7BnEBcEr9BqXFkC9gM1m6abkN+OIn8Mf3Phc43OV0LY/wkL/LpVOiaG8jJfXyKB
VK0Sw9SLBfT+ip64qgO2Si1Ocl+Y4KCw86JOJo1Z+JCZZ0kA0M8gCi4zMnteSyUg
CXcoIjooRD58o+5dc7bG/BcKnYY695gBIGVfjbqgm8Ysm3zyYe/nHCahDjDImv9D
GtpmnGvI/xo62OPe63cuEX3Qambn9DhnjGI4/u6IS/0OxYRHJl0O5C3XnejufEqx
LeGz73FPZAsaBakxErb4MYZVZGFp7Lr446KnXH7wUP1n67GR+DRd/9Q9NO9bcjIC
nxK6CmJGzcb4owMJZ8xEZR60JbFopWG85yG4qg3d9GjRi67wYz3zHkBMHHx6oaEc
+2OPZePlF+6C3kwlDpnUFKAkyoRv5PoDF7/rMoKRY9ETqUrnF2eN8cTKyL1BGeby
L0hrhrz5WFvPY2FvY1LYXr4nv9eWFBLBMiCwG6rLJ0VP3G2GoQwRVNFF1w/jbL3O
lE8FyXx2ncra9OXsdBbEV9poj2JALZnX9tHCveJXAQhVDf3Oy0pkyNocC0f0Vysw
XjHfFJXArLSCwiiV3YfwIQAAyq9cdWk3oZhuiH81AWuhpMAf8oA6FtdnTqWmZu4W
B9pMYXT3geiG5LmbCvFO7o6sK6QM81E9CnJy5Ek1qkX6nxjg7EZoJ0tqP1rfloAS
9JHzrXYOSKfJhJ+6KI3L/y4qsqZOkkc6hqjNzrG+M9mXsq7g2y28uVZ+f5gvHxMS
GD5px41YTwZC/ddz51MhIXDTntyi+6jBruhqc5nvzYVivHbBsEReJ4n/4fyyJmRW
uu7ELRrrBy91wByrFO9GDx9/tTZtgENK0EIldSoBvBQwn2qeCkPcxdgFTh5irXPs
lnd7c3WxxXGd74pFdj4cuu69j3ybtTrPTzLQpqPrVBKYSaN7AsDDfj+RBil+G/Su
ObMwxkiZE/xosCSVprxuNQh0erqLEzd2SmPYuG1lWJs9rdnRqwX5flxsQgnMXiv9
PA05a4UAUa6HUfWFDU0Zl52VL/X8D6LdY303vew+cekoW241oAvicL4T3+q3KggJ
Jjwi2h3ygdxu2XitIxRQtiu1bWtldUR7iKyU5FfI6xXR3b/lTTTCPH+DsWHigXch
NLIbYIrl+FP4jakhCojPYXfplcTJZbsAox2vz2jw0Z5o9AHW7svCkCtmMzQnXSHM
c3kh6h4qJR810TSRFcwZFvMLtnXViQ+qr30HXyXzDTdQrnjHBrha4s4mXt5/oECS
dlrqiWmMkJqIH1hAIz+yMmn4sqB4rKZD4EfNJgovdduSUtYwcPm17fpZEBwj5C0V
V9bzi6W6rDd3tFSoJ8TZrgk2LNXpvBTrsjNrS3idf3b0tGIVWmNzHZjk55LzMklb
2wGjPQNHBIYKmTrJqzu5LvdRxVZyqRTtUztzVoMJG3GjWBIDSUjNUhjpKw1393+t
6qSm6d96jR2/LQAe70vm7yXlNRe93iqGiHjmIN/dZw7uzBMY6Mm5p2rQgNgpOHf5
8XeCoXvXf6qoFXFpuwBHZWzPdSNy05nCTIcDcoztb0Btr0vRgCma08GjJYQKjosu
TgClwRh9HzuxamBG+MnT8NEKY855CISoY52e0hgf/c0tWaC3BxoXPnOn6jOIUdfp
zw7CNLiMeiyz6bHjZLJvSaTu+foOv/t/aaIfyTZCg3ZUd0+2wdHbHmAuIjJN71P5
ERr5i8rcL3+82dHB5eTtODoeo/QyIGsIzPtHOQJZIaoFjQeQ4WokvtvA7tYoFoF9
gs0f4xZPNByuA77h+Nd9PVW0qHkMQmOhlHgZ3eSG/LJ2cXvYfQoiSFaB5TDqDhUV
S1MfhQW1PxpZS3T0a1zmjyvYJOQ9uaiIiczQ30ZIkar7emyPkaeJ9RQw11WYyLAp
1JywhH4mn3fOeP9gOCAtNJMxMmTPVonJj2reO6didbcSgk+La+zbiNoTkt2bUUyI
CdrT1p9ryXnX8KPN1KfA//kVLONRoDBGS0pL8fXJfDy2YQtyiqV/W6gZ7q+nb8fH
elDHDuwK+szHM8oC5IaxzRxwLjBpJ6NWoQ9DpuaqXHH/K8u6HyCiYrbh/2Elcwm/
wc0lTnnSpGaYjwNZ6A4ZqqZtN/AldD/fjFlCqA7PkkYKgYetJWktjBNZsqd4At8w
osHG/h2AkxaOnuoiY54z8zwaXxWpE81V7F8aI5zV9/BKHoBGWYE675RK9yagI/HW
qnUPI1k5BXQbvAwNgKbL1xG4MSWyeZNwOIiJ9Lm8LB+paI7fHpJcGhyB6zcOE7lB
4UseBwmzqfXW7mOCLWK+9sqHPmKQAO88cBz8lwhPepHdf7/wf8+/ry3YPviE7gxW
fuAtWxWOgEsZBFSzjKIFUFjmcCMEbqWsc6Qbtr8DdqJilu1bUomZiUVQYzVRzzWw
zUCJojohsLUZdzuVa1E3gA1q3FxKy7XlxiS9sY8PzccmItoPkZiHBknA0WouWxMV
KLPMUhBLdpUn232mv2wOMK69RqYUbMbq5m3nyNH7WjHnD8I8nLQ1BD1zYsDSIQu8
tmjpkShpBK7XNPNavLj9nlyl/xoGU7n6gibto8qVw8/W2UmKo2C54rb5RE4ZH7nw
I7CYBCdWzMHWSG+PjLD1ZxqVZ/kBGd0vxEVs1FysK1sB4JpSMxGsn3aca6vLh9wJ
WRtVMkeiaDMVAeoutDp+Ny5uS9rIlKGz6DgWXE++vwFwvgf48bHiaZSWwmKP64th
XOBeEmaO6CCM7cl0RXG7jtkeSeB1aSkG7w4ILih5+TGa03ApZAi7wdwFSnh2NgjV
XpheV1323y3rpMfE4pxDoAYjClXuNfNdE8RxEzkHWYQnhaYoUAmZHdpiTNfNondH
rww+FKuVxrV5GSipPLgcDFaB2xXdEkDopifU3yLxzVdIku6RfJ94mbIuNDsuRmfU
yvaGJh1lciFWro2fvoRhjJjlE7tzKKzPY4uSGrfbhi0LXicjrKVCtdXbNdyP8cef
kIym2Wb8Vq+FiiYMvOi06YmJ5pGnENEQ6fHMNElxFVBcaNpdoAcnQ1gqKs69ORSV
/MeNhKUJIuP1o9i84BG2TNwLs77JGF+5JE/e0+Yd5TSe1l8Qa1cMSvJdcAT42omc
854UWs2io07WloEYuY8WZYPUuA1crpwrn2aeS2jf9fx3SHbTF3Wi0e+vCmXdptc9
CEGEdzXUrtCb7g4+SlsHCwLN9I4tsZDMKsV6M6V4qAI/1EPZRuReBQNKnKEVhmIU
yTKGbwGAV/ARP65DW6oBHdCMnGXiX/eMQReIuueiEV+e05P9iN37FHic/jnAb5De
t4maZlpyzJrBljMNgOSjZIMOU6i19gRlSMIEWWn5Ky8Qc0atDNloYoC0x1pAekzW
39/mCE5pK433U/c/PzkeGSfUih2WPdxvWkYsweYkPCZUjDSmaWTq7mtgMu18VbPJ
7Z1G8MZyj9+11wec9Y/Pe076v+nejktvMEW9dfa7JyrrhqVGr86a0tKMGii20IGs
1Lmpc2TydnWxsQW87Yan5E0I+2Qo6GBl4r9zVhZJEEFTH7fuiuibDCRTPJtWpsds
FJIo49QS39YSkBBMP06GZ41Er0croFefdvdTFQZwofZO5u5qBbi+QBh7xqB3vnwE
UgkZIuB3Y9wsJBLnOncu7EbF9j1+bcNIYa0lQsvtzWySdgPic05B9j0mEHwClavy
qa1ZADsUuaHAj2T+x1+J3olZe3F/3BPInhGWsIp5+eJHIMNpa6egohlN1A17b7DZ
aQBN4JMsm5dwkhT32OwM2P/8+6M38gKChss45x2bz9BUcUShS6Br/XAtvmHzO2mD
G80YBEuCtShIm6rnek5FED36kxeTjVWVp7y603B6/wjCgYEF47P+R1L2KoqFubRi
w7S8VS+fwyMa8xZVyHg6iZ0Weco6mQE2EOtDwy29AQma41PrBgxpz8vMtGrGehAF
BDyA9JW2jaWr+Wyf82cWPpiQndhmYymjE5xJA0V+bwKdaLeHLPsBZeurpPWkMw7J
rsh3x7QkeRjHOXd7pZv9l89IJQc2htolZuf1UNqfl9gUGgU43LsPTQLVcHEOz0vi
7Pnv8oIn3UGtHCLhTey3TsHDlB2KdPStSjWqBzk5gAJegSpS5SLdrJRwFCVuGkjF
9ecm3a+KN2wRYNsP1pf3I6E+RrMWFhw/r9xNWEULUo4NVE889N3dphmXxMiTHlVE
BvZ9j39wFSzoFLK40Gi6FTHvfOOuZJE2AgMiO2+Rh7cfnO+0ZJG4CDWMt8+1LUzx
5EhwKG3JuICVhzGzho+1vBC1XnyFslEcq0yIQZIxKvyhdlpUUYHkcA7YqR2huCe2
EyTv7Hy092zVdwRdAIasIvOAfwQQfnSyuyBD+WU2TiXMkTtuPlETLL/ffnaTKAqT
mmvvd/fISV2K2vHlupfZXbN7Wdfa0r7sU7k2cKjsoKOrZto73OyhH3siyJiLFrFj
9S/2FBo+UmLbd9yaJKwkygCZubotNcnxxXhetogvmwuvpMk0+E82lmf5rEvPy09a
KXK3Dbz0D+J2enmjBB6FHXWudLxYjlAaFzaohpc2MD7OubCB18fS2QScurCl/38v
xqD8P8igljB3IrgLgz/S24xmzMYv+zbp9RgOl/TqtLfP7hRx5nRO2YEEqxv6tAYy
AXBDnuEBKTubKOGCfcu1TwGTIg4lSvfZ7sOzU8eIKG8Oas6jVyHGlvpY7rkdePme
YAIx95MIKkf7bYwOHUZf22BSDUGGJ5ohVJnM4Kjy2fz6qKBE1A0H81Xq7tGCS6X8
JWvnI9Of/pHB48tyDQ8k21ka215QgcHke9ZJxDItJoWFu4ltYN/mzdqoTOhJBUE3
5EQL1hvyq2oHjt0GoboeOjhv2rvpqNM8JGOVIuTkAvsV7edMgYyf0croe81pocc5
SCKxUvwo4lQ3pWI67rcHEbb3I+LczbOw2WJnjHYrS29Z4j6wkfq6QAw1aehMVbtr
otBGOqJnUTQQ8NWKOpbhRzxQlYzNeo4GMfQNxeMl0MuEMqf1t5a0m/KwWM9mnjM7
HaLxHrcrVC93Udr0erDweb4804VbohD/FWa81oSPLhgOJQ2heSpvvCUOTn/0tk4X
gAWCwDMhwVXnZxf3zTpP4ut04s//WwLwsldGE3hfxaGUOKiLamjhdOpxelnFpqBm
WTrbfPcQhIsYROtqMTflvinPAcwVtwRwmSBj1/qTMO1mAf8noyD+1ZBG4+5FhOYQ
WTCbimTSzqR7FJFPdMOM69hrO7VpqjHgoywwAOGVKuYSOHeo83qf2Tk/BIXmylDo
wa2YuJR2e2m4HT8LxA2EGIu32k5bsnXrwsfJv4/7523Xk4mjdkAK8YpK3iih2wWr
Azl+L5miSnFMcy2r85qH1keZL+6hjXziPloff2iD6CAMpqUFj1nxWEu+BdvcaeOC
qJ3/Lp7i+KNw5xXMcmeDOTs/7gnv5C4DORcubZ1G6T1L25VpsHsMQR094o6g5myR
mbdrconU1aju54U2kaLU1vlhAkpPtbhXnb0otLClGeicKx/dRkKrFBDdGxz8d4Gh
W1y/vZ76JyjFl8aWLAv7wVNoQVpxFR7xIrJetoyQihIktWgXY+zKHASMwDD76wKj
oHWqEbrvwJN71aF1Luq2DSHFrlIok8KFu29yKu3JhmFT/Fj8DmtBjTzL7X0JfSPx
IR4WCj+9LQnR/Vd97sN5N7c4+Ml9eVxP1/oCcRjwUgWvV98AlhNQuFpSs+UOfVd6
duYuV9A3i4ZFvCD5uciEi3XAM5j57npD8YpQu+RoDHZYjYFMljdETiKLn3vrxOl1
73Beny96mLDqDG1+RBXl0hepR7y4H+LksC5zHIMgys4iyVN3jYwhIjlz9nMTLIty
25Me9tbe/RI9iZG6vl8xTj0Jraaa0HliCJD3raczaDJVsknXBv6pwhM4p3cuxgk2
dH4Z+4TQOCT+ZRAzPNZsCjer4YfM4jT8TAzHQzueUVU5wzsGX8QhKo0MzS3t1mi7
3Eot1+VVhQJFVNXdxfB5Kz26FE88ouMzNwzRohHbc9PsyA4f1dXIfSW9KuGEqG8i
29fInrp+kHiVaDiFz1M78eOW+SzAYd9syYtF+dz/0b7eXZ6Iz0AlCBBqQE/xoRRG
SawEBMVRNOZaC1clRr3/V9NQ0w+QCpgV3w+42sjHHyhlAoB3n4zuvJnW9ecQjFW1
e6DZcAD8hvCDYDuXkO2htDG1XnP0rDuQr1hjbjx7bODOwK7c4A4c9yQpqlHHxrF2
nX9wd7cK9+LO85SNmimaE+bMaJjfXVA/BFT5pgMNnDMvFnTSoalcyE6iOwnOiQRZ
GfDd86abLxmlttz4j5AVwpMHvn0rDPzM7qRzmcfjsIlR8qBQkMXYcdvIf3j0Tkx8
PX1+eFwWWuJcUBA8WKaUFbCP/k4tDPfYGAxvWKdcbt2O2hXmmGGNOAACWUJOcytk
UWlkPRMZh924/wNKEaP6ZtUfLUMc2PdAVqHbuqMrHXUEMm8BB+muC0DC6/+jf5a6
rQUe1xSPLPbg2RdJ9GUyVwKYjGaOqfpctadAxs9rYQuRlGkKxsfbR1tCMqErvHtO
vkAnUBIPEusJnbpsTGv+rRR2gMHHHE6tO3NfY6HbH2pe8aVO0GEVbeUXaMTzeWAY
40X9Dr1v4cS61Av5UTjEfXRkomrkxx/BDKWszoV1InTeUvM1clZ6rL2uVwKtcwk1
BgZHQOT1KdxYDw6/EidXDIQ1ShIJ9Hy8/n3OLNM5odLZHFu4jWEM+WxjPQvPBldx
GVZ8mznXf3tVRS6ht8vTjGTMyDWObsqbeL5ZbHoEkjNQswgl2AHnYxiI2MD+TWe/
5T0mKBgF6p5f3W/uKUNZQ8/dZFUcdtFgqVaB27+LK7NAMTl0++4A5Tum4IiK+/BG
aPadouGYCSADb8wT3xR4G55YlIPlfDvpzM0GkAbM3fR/IAhFmADytf8QIGUn2hll
wTsVQOFfUtbYeuZ5K3QHLI4sYZE0jJ6SyQEA/C/ydjIaCugOlquq62bc75wzDPxD
feryX3XBo6W77BxD5CIfvai3PScXdvV7Tqfa2jaKxj1lLaQ1+q+x1p1YMbGUS2JY
NtbUqHH5tz3IJrO2Em0XBESw1NaBbSaL9mREmxughFL8ydJ5ycZqeHqTlnofOBbq
wMNw3GNIlmVgM1yNClObwcIHLlKMvsP2gpUK6XVniHtVvvXT0mLnAHd2bpbcfcKu
0ceV4Sc6Pam/0R4yR1EMGU05jejo75s7srqVTuC0JfM83ba6nK2yWcdzzZC9Vkwz
cdNBPkVrY+tse4Vjwbtr/s5/wIihL8VZVfNoJM0EDNjSiIXjSB3jMTnXFtY8HJMr
UvKqP2fcEmddH2MvS1onF+bMj2pzb8GAfLqROoquT0te4C8ICiGW9zKZhmGxFMiy
vi2IdreH8cOaECZu2E8FAV8E+edlNT7UDW3+0B+DEQeHxB9VNN5ANhE4wv9Edka8
kfIr11xXkK9MuKAtgbzWQJTjJPB2tkYSqiq1BLLk7XYhd6npTJPMTQeHxlcvRbL7
AZjFjvF6qDpuTnSv7M86YU7IO6bdIkCaZy6fd2VffplrzqOXVsSwMQyeDXD8A8JR
LlS2lsVgpzgjdCHgiJvC+YXYB0mvLxes/ztXWg1BWMB0YP4wmTvx+q0ILF+KIrNs
BcZWsLtwruJbPxHsyZL89hJR/hKfFHIugN5GJhLsU9tiezim12nN0VeAi4g31/7x
WSGgSzt/heZfkGsipbGNhXFAVMLTuFCjp4HlXhqWqLHofcK1KHqTmJMZWkgcceJj
sZbmQlzID+FpZDb36DdKiBi0Rk2Jkt5t1D8sD7l0bJZ2VqA8bfWJz9EceSslRC62
FVRco4yKod5rQ06/hRZCeRatNQ3G43zYEZtSQlovw1WQIWXALuXOwtYO7YOTznVz
gGwl+At0Czd3m9v+Ehb52TSvQDGehubB5Mxj7/f0YqvTHFDPcdtuRRrtILFshfrG
0gxsRlZtYXZL24uzUY1ldQT7+iuklTUo2WD+AgIYYAHs3r6je2jAEBCXuTWQNzCg
415k2zI1cvyNB5SIf4yhUPFz7r1gQI1ZfG2NJ0Qc1AG/FnQYbtGr/qeFNiknyqz0
YIAniIA+NM5wWP1yx2QL1CN30kPW+4FG7QSladT+4mnM4xLVpFPG5qK9eKA/NoEs
eTONufKIzxNuI7x6TlWt44cJqY4Y3CipaOqU7Nxe0AO96CH+nl17wh8bZfDmmIl3
EOAn3cyiTqqwKrH7j7DJOREbHtiAJO5cOnU+0GGiNZBLDpuXlfDOU1CZ804tQAMX
eyhmw2yKU6zmIM81ASnaw1LGJhbA+VmVzPysNy335qs1nLGfM5RjqBQ0RRoXiX9L
IPniP5kFAMT/QJHrei4t2Tz+FXr3tzzpFWXEcYwrb8AB6fjkzyvXGX8Ecmh5AGOs
a9jMOrDQI2Lf8QgfgvPLGzM4BuKEWjsmgIsRY2GGmhKhgMlWgnCLZa8jp6JBcByZ
G3lGYtV3pioNZRjyhBym5m/rLy950BDihIzg/TqudFR94lsWq2h6lsR0YZgtlqV+
taY+fIEJFX/QG97mbtOS1Il2eALm0/zr/xlfM/uXzz/GPKnjZHUdrKr/iQk1Hf3s
QHa2PFMIlM3c5idck7UsbU/ZBADTzOXu0Nx5a0g3Wlvq2jMr9yLJKlVOFH4w39vU
mjDxdEKU0jrKCZC9n6upNfwSQlmYDrMhZF5ffnMr5RIfDqzGp+K3Qtmg4enWru3G
1cgmO38rNmmQMSp2FX1s23BrSBMGVnN7OhYys6yRgoBREljo7PsWlg+56nVj2/d/
IOLdrAudSWg4dVVY0lhIVT6yLdiLJDytRykpalCxoPuygTyJk1f6jXy3FJdXxQRx
JPcoHNj/CA079936VKoDw/HhSqiZpniaSWlLcf/1wQj/VaSS9qjxWpxT2+qwVPDb
wBRJ2ykx/syrUZ+P0xu9Wn4Qtg1BxD7MzoqNhuIYnbtF2kPjno9yiD9AhVYBqDln
AdJ0glCte2UdGEc8NPXLPvWvGaVtrsfyO+1ed6bUAWyEtwaFLsLCqKSFnVYBtopI
QR32SmkpQnEQ3OYaYzAuSsXEQJS/PKgt912U+HW8xC1/dqzkW2WeAtuATeyNBf8b
cs1pHV38qWWM3O9b4AcItJUTBCqkQviprLZgPr0x3gPet7jm7lu2QewnzVi8s+ZZ
7+a70CDy7EgzA6N4cLuEI7QPBC+PPzrlE94DxdQDGs9HDDbaxl8xcVGllXgvOusr
7sjETjP4ZI25X747PEoTmSg8z+oSeurXw6J17OUOSF/JnLlPl6PeWz3MmEiWsgDm
nS2t0QQEnC/QhcGX8yynat4kFD8JGs4xcXdJZ3dd8nXrGsfegNVp8Z9nCc6kTf27
GdGGhpE70Q7AvV9u95BG0Kah9bf8PPzXuNeYP9bveaGoxKoHwO8nBMrE7z4JRmdm
4ACzjT0heAFB6uo9IBB75bapPeDjHeiiUD+VbP+BS4VAUi8hmphTzvEzro+wGvwp
AnxIKxg1HkwMQOpfXvRGN37J9YESLTmyrSceVJ/OydCfEB5eyTvcXN2N7hqjH4rJ
7vZQTm7V0NsC/zFPMFcuT1hEX1qpANBR6keoLUFEm+GrWsZCI+skthX9s/iCfGCF
PKIdIelRKG7Io0F4Vl5QrjlkznONlev09B4uDL8UIuwrPgPJ2f/ck8vOSxrq1I4o
PWVHdUcmphys66LY9a2w2S0a6C2cxH+YwiVS7CEjYZ6QWXTvqJZWEoDaJr+t3XsZ
HN5gFz9Ra/x0bFi92OaUChQXDy6iOZEQ/rl5Bgh8d31bGpyFaTyN/GfMRjS2IZi0
hKMK5s59+w79ptOtS3cSYYzZV/0Eu1jraCJYcBuuPMz8Ws1yfpy0t14Aoq+i3QFq
YAQk0G2HOyOnoJK8NVRvsIO1bcxn21UoxDmpB3AD+rCcoWRiWBYBQkaLQokhUtNn
h2/Wivq8UEdZmOwcneFdvnGPECshwaBuqpY/FyGerPhuwCbfd00496QSIM61ICX+
FY9AMuAO70lXmfma73m69NeC/0hlLHJP1eOcrYnkWNeS25PJC5T2f+kEAEOFTIGl
j0n2MWrCTQ7WZHGGs/blCzsqTpmGcE9Ih57J7Jixj7n1jwNE65B02Iud3DJRVN4S
BDH/zxI3teezeyWaWJvvELgg+48hMWrB3xWmbEnrISS7L1x7Xci8y4bagvQFVv3k
OcqWHCZoTu+Ym7MsGfxgx8e7JSOs7qmJ7Kwq8xXZ+zTLffzeGzTN8acbHlNJHGLj
exPjDGUVoXQ8lUBRkQdPj8uZkOxeezczvrhIIG3wSu7ywLvlnbnqiL8DEBLLJdgg
0GKihGMtw174zcs8/xr+f/965u+gExNA4uARTq7hKZ4TQlBL0oQ+I9e27zWlPfmy
ClsGyF/8R6V75tlIrxPdKBxczXvv0lc16ClwF0vQJKCoxTWD7yidb+k6MWSs5TiO
JksVL+VhXH+F0BPRLaNGacJ0Plosw2WcYY6TbbIDZlCzQlkXoHpvsATKdBc/A9VV
UymS+12WEcq+cWJcsywWyYZB0X59L4flTmh1CTIfA1+8cqhflKhkGNZtriOfApZE
/aG9BRL7XfQBaoHwha1ZfYR5Eo6ToNWHhe7LTqgRhHD1yXidLKVC+v1oZsrB+gSr
jKRnfsZ3u6jRQluFl06kTH3dm2YOIniQBWC3owlstobmm1O6koVlY1HNSCTKScMQ
z7DuWmYlm59UVPgp/lKe0Mi6nridZ1MVqjQSuY5TS1GeLxIkfay4sF7NWY8oIdl3
GDG0fGOHmSC0weEZDkmVo72KypyN9zT+Vt7loFaJiAdbSbsQhweXnOi1SXjtNyzn
kZWq1GNhuFmjPUwIRkSw0kOm+wPvKF3Lq7O4Vs+0cfmVggkGaMSyuEDLje18uZpW
qxiMYMs4QGs+tHkWHT/NzUSvocB6yYXrcp40DQX1+j4dF+wFUe/EEl8HbTqQU2QV
utWi5bkGNg+5YLromecK/ij5WwdcJXVKbnR17OTB1uJ41gJzpC5Ld10rfCmFgcm/
71Spc4bBLyKPCV02zFJeWzgL56827QIcMkVZO1C8yN19esuUdcJ6cV5NJiGDK79H
+I+3Tlh7dSJpWF61msRg3xd9jpSBpDCp7ejrOWBERWwSTLmwflmAaaTxvvFPKm6x
SJ5t+ySBpQcAvTIa4YYMu6cyXLr4eK5ldalzhg4LjhV60/s/N2R+lq1xLZoVsp4Q
6UorkbggwbUMxHrENMQ9rx1mYuIbbHVrcKAyDuqSSFRb7e5GgipZ+Mqy4P1G/cRE
4lEMMRIxvIJHTjRGWzOlqfgTRrEVM6d70AbpDvztHt5Pfnvm7L3VKTOnWEpQBSnN
yWSKw62KeAKF9DaNMa2uY9KYnw+PE+qmSLZ+rbqn9VAb40CFhHKcv5LfSHF95hGs
F7HNL0L2zY49sRsIBkzdijjGHQevvAJP30eyi+BbxWHdUGoFLLbIS/p8ZpGzLHYF
TbFA12r6W+OICoI+EzSc8I/xBkI51SFvlgKUQw7SH3PealIYAFQAHrs3CHOaqExu
VNMgm0oTViglfzPeILMc4qD2gsvLB6cwAWMUf7VznSAz03v998RTfyxCgagSzNve
cGbKJHVWX4CV76H/uCrooqSxv367CAgjrzZwsJxN2u+i3nF5wt2Fm3QWs/habgTE
iBDUGNHF3DFVKifp8+lLXO5gV2GQydxT+u+/fa85oys1ef0pvT65l7Y5S1fj0g34
OXv65J+JW+TwCOIAzF9hxNXQ/mrsX6LJ5/E+O44M+UAVh7KVDVcfwO6BW2C8xas6
BAmh0Ym5nOai4yQhUO+PPcW389Qqz2Gh6VBT2h3j5NgINYNuflAFq3GS8HHv0yiz
a4qT565oH49rHtsFKpGt3cMWZuKfjjrd91no1d40aC9uZpUMpXKWhMbWcueY+0EX
EkU51HXAArCPs1rXgudU8CqfTP90vQGqq6TItfnaZY+azyUqRJK05hXhcb7FkgAJ
yxsXgpyvmo2mxAszI2LIxHyXa5epsJxRgl9D2Pgn8taFbc7FbZK5QTBrckBbcJOC
LcSoTinaP0kjZVJyOz5fLAyrCWEvUoZkY9G4K2ntExj7g/YHEdB9esE90T7SH63d
lkG3804lI0VGPMx6fKmVqBuPlvD6u/5RR8CO1gLGP48gHW6LJPy65NkMN9lUmQNs
jAP7IrU88zYNjuzN/REhH9AmTvPaaysPOroRP2p3CflbZ00RbVRa+gvtUHN3t+jQ
KWlhyFdkAqL8v1FBV+y49F7VRH/aQGdIIoUFX0byvoUS5PGBclgozPCOAMRSayn5
PZa0yOug0hqghpQNz7k9L9Z9C5zhA8o83zQ10TfhrXIQvdUw84TgfphMyInJGlM4
SVszvv2NccPn5w7w1uRChVA/94xsVlMcJZE4UFuXyuhgmkHPElOHzgAiDyz3tNcd
XYkrgA4DvTeo6zoqRTYSHXZz0OoEHEjO9SAC86yA0FfBTXn10jttlCVDml6DTHxc
VrkYZ113sFXdnWwNaIj1PA/r2U26w+rb/PmnJXuY8+lLYLSe966qM3az0GYgDhNL
JgFWN/yUw2k/OyNXPAq0AXE4Vg2OpicGXr64camWrlh5WiIufnEVcseujwHGX7aZ
/l6MQx8RiEaBigABRqZrI9td7VexFpD3KhwzGQ2iUYLEM9XiVAWdPdszc1oEnu84
C0osn88buqoFXI7JtR+Pi6ZADuMD/FYBqIKx7hqUHyKoyyQvnSRTRS0t2ekW80KE
lRVyHPUEJNcjf5MS0QNE8gkkB85xQypDpMbB2nApGPwxJCYHWEO+XcUrOXNu9rWs
ISU+waUzxCW5j+Ig531EmYQQoMxekAtyDkI6MGQyG3ssuGndKu070hRd6bJ4qp3h
wd9MlBQTr3EM8+Xg+p6htBnn+nyFNXhZAizsYMJehKuBsrqZbtRt1Xy8D0taFhxX
uCBTY/b+WW9VBuc/jPmsSgO4liW90rrmaN+rjxe1miR62w+gbW4/ydsUf+/9YYk9
yDgpl7r27RjTlpcYrt/YsExXFqlP5r5UI+Z9kD+oUBXZBgq45nl5qPjRgQ/bEzZR
/kYHZRrcZkkPFH62AHQXYWbN2oXQ3EfO96c+X0urwxGgmVsgEkG9fFfatJNaNE57
dNYyEqfwxb0vF+vYf14DjWq0rqriykrDN9w7wwI+cdZmKRpPtKD4ua/Smp/A9MVk
aiS2XL9a9FG1sIofPqe4LJ7AEusldadyXeb0uAvCEJAP0GA1u+ZF6QXe2zbLK3JZ
stLPidMeva5/gNRJ16nW7T37qdvzMGXyhmSE6qkovU2aENHhq3nlLC3xgX6BrzOz
kT1neRusF8q5p1EVJolYnBaMDl32ZNJe3Zrc6wPtfW1metdQIkD0+1UgKLpuehQP
bjE6bgj1dopCWBNc2f8aTjZw9Kr9fDuYIot2h7ZsUvqe+OSVrokkM71HqhT5IV2J
m+4ygIaBWW4aJcWC41dl/OT2uS0vLqM2RJaC9fxgN9KdSzUJ3GBUSVGI5rjRcuPU
Axp8P/cIkbpEIHpK0A75471vd6LgCh3plZO0NEb10O4PacX1Cd5W78hfthN9C/Ng
SbHkE6Uzwgsgmrxtnrr67U4mJvEfBWSF0Sh7PzyVCQUxBHUTlrwiTs8XLc9KsOAs
3uM751rZl2vy3b23rmN6LJ306/sba7ncUnGQDHk3QBEt+7qSfraa25awHlYB1FJ0
LJDOtUJ3+XramE9MhEwaiW8VbWek1vSICEFPoMdQD3WSXSOqNxoiGto914cF/HMt
j5SudbMNMuck4r8OmdXLDzKOISjqWnIEGUhZfGJ0g+Rzc6HiSHncl7DQPdN6X4th
iuI9a3Ne1OB03CULot4R6999qXaB/zJDjqDp4Unvx3dSj1s+j32yBS9VjpdojGfB
VK7bFq/952kXGnS8Ukv4rSOvuphfk9DzgzXz1qqYWJJdK1XGKgXrVfQ096r0unzx
NH4Q9MVFwrm/J9zaKiM+Y2vWrYxKzUlu5Smg8sci7TdpKYb3Ue7gQwbG7HlDR9Sb
gq8frsNlKhG+YhMK0f34Pynj+SI57OejLsVgsWR9PTbeQwnKiEwpl1aA1u+SuEci
78aDJF8bU191LpaGHURHOfjAIJ8BzVwR7cwKDkoO2MnglfaAlDiq1J/muDxkD8LV
S4CFNvH6ZjAvZNhiGPiuEiJeZlYJQVJeajPl27jtvxm9F2bEeWm2OF3cRNsjcKr+
DPmEaCz0pj9aOTtXbOrw0JzsJHdDceSPI9Ij/QDNH+oACir/9V7bTJF8uo1PT/Ni
rdrlLLEZxz0RTHYzhvbvROG3GKOz0NdeT4Tcfo0N/UmIlXjNEqs2w/8eVa1WyaNh
HDg0g3dfSD+OL2m3tkcGPyyaeWlya/gGVAz42gix3jWr0O3nx0AVhCaqKduBxxIZ
QIWYO3TT+AF27n4cpoYiFEomZZtxCeb8qZixdgOIX4bC7DaQWxP3xt/nyeaACeLm
8MUBEfGDfw0TFSqpvaZNKUb5Wc3qs+g31ycCrJ/oBm3FjwB2M/dqajS1hN0wywQG
yZiVK9TBwfGJpR0oLrIvsZG8gaV/E5WmgxyeFgwINXcwa6zx+6oPRiqnQJsmyIiw
yLwdKkH+7yZ2HxuxiSj5ueRokrvG5SfKWXfCADR/iWzkL8MKdB6CIm+YOqjyJGZT
amIRxJpHG0Musvc6eV/hUq0Q7L1iPIVe7FoMp6qAa6tYTC6bN5NRcDX5KDSoHo+Y
dg4X64l8KuxAwuRvitRwtxaFAkUjJeHo/ah1djkDB0AJkmRMXfjQ+eproDbfFta3
tqa+A4qF+LDmT4cIouP7YM48nkdjPSRzvWr/jituZ9Qb5zv65fIFvm2BqaLm97r7
kFE9lxH96XVr+L8Fi4EnpFHY150zxeBLPUyEZPnuqEsuC2xrxL48ILZgL05p7hUD
52Rr+dvQhWwnj5r2YImB9IUv3ho3bexthenz36HN0sceWj9Lit7BP9Zc2RAQBMe/
vyNsH0Lq1jkHRq5IUibKSCjZ3uBOlt39ROUo01nh4fCQm+XCKAj7MzvZTVu9U889
x5FdPoQpIZtcDAgNMUG9GeUyaCrzzNtNcVgK0K27weeuqAOrDbUzLNcP7Qj5K7wW
FiiDNP/MZwfFQrTLDzj28NeH/cllNk6w5Q1z7pL2BGFQVYTDysG0valXlhGoqnzn
ZJ8CwE7REsCJwt6KW11d2rJiJJ56u1MSE5Y7/Z6Wj4SH2q1Y+hJEpcyXws+eELsc
0aT1Cg6/rUfmixxhFXT4Inq9ZU/iiDGKHeI4K2iZyGol3XeuFfalkjXGAj9QhIUy
uCDGq8CEjW8XremzkTFNsZIBUI680RhDmZ/mZHt4TP4ddJbbc01L3VJf7HUA8TP1
vrFCYdaLFID3oqdMaoskHA2xvroLkDqNScGS319VQGZQ95vD679Jmo9UYW4WDxje
RmrL+N2MfBproan2qXvQwZ/ED0KT8c0IarElYiJH/58kVS9fMLceYYnwrcBXGf2d
gFASaI8gfmxhw3HFnWMQtnNhnWpAVF8p+91R9elLAZo/OOFGmZ1+pfeTHa/YZ23D
VJJIi2pu02jqca/Sdx1fBiPK/d7yor5PcgFEOmYqZgTOJ7shF/pdh12oyDNgARmW
yVzXlG/5NPQxHig1/z3gOzFwJM88SV+uRvWZENAHs8Ouh3h+hitdYkPqSG8iyj/w
33muaEhz1/UBVzzcBpkrVa3RkWdii6Km95GywyDM5ljWCIP6Ch6AvwztJxdpbKVJ
pcMafdHP0xr/1mouuRMc+46Oz02kvwQAf1gqRHGZw50IO8fkAMk9PxmlFXMVSvRU
qr2iOUkFNq6ep3YkLhtBj46GLZ9ozTuEHGrwYHGxHzvhKnz0vz3c7ljfc1mWydtr
LyXzyr1NcA2ftjB7+ZcHwSc150A+/5MtV0wFn+IVVQ+94sBgYQC01qtqz/S7+ek1
HbNCVLFMTD4L1pmJBx4bOJeF8e6hfB74F7haYmZAPvecPzdWs85kGa0FuZyKAffE
pBR08r9p3mCOGZdYIas3vatgZln+/pzjF5g0PhhcsqrbZPpmorRXtjfZW4kkm6mk
vJ9dDyTwWe8kqk2oRKnhKXMQgeR78Zkl7zqaMVsxGIKlVjxFC6v0uwvUtJ7hCjkm
ooko3JjEhD6YDORacXob4xTC/ef1vaIOszRBx6eZo6z6Tf1A7eELLW9j1Q4SMFIp
tg5kvUtfu4WVPWiOgRcecCo+MS07Kc93UqIDxXqoRXXDtZmBt3biD/OgDektortR
IDWfFIjDAUI6ZSBF8gJVfNt8TYvsEmRqllEWVVK4OLv9hMUmw6VEQpl1kNxQMwtE
U5XtYQfoA9I35f0u4Bit7V0TbFAmxCKbZJU5TX2li6tfH7ObU+E/Jzx9zfe6HcWA
g12a3xeJzqKBZTYIQuwCqR4O5YfQnT67I3M7oY5Xk5uAXW/p7BmkW2QI31YVQ+lH
XTBgHvr7arcP/7n3W2Z24XvRwGWAo3mGDgVfh8Q9C7auW2Fxaf7TqiKd6mTsbWT4
/YTeKDTrxIrCSBLoxez+mURRHgy1m46bo2STHX1ViGAEAFn2Bf1DFwlK+BPzyv6Y
YNs3IfsswPor9RM/9szR9Twl4PsvvbXlSj/qEpnbikpEzQn6cAQVl9s8RsnS2Lyl
OY7YfhqmVVyHCd/76lQSvQaWsYM43KuvYr1mzk7LmLaHrvqGXIIqaz3vw2M/BgPy
/736Vzo2Ff+4mUlRjlu5FOkwHNz62u3MTfX10CglSiuadnK7w8oOUsDV1Wv+Lyq5
VKH5BHHbPP3qKC+Sb8TXnEMKxF4dg24dqRWImlssCV6z55xzWQVZf5GJBKYMPFQh
NzVojmmV2LoXDA/mKOqHEBssE1XNzUytjJGHZjO7q9sn6LxU/+mPSd0C8zbyrFPZ
6zR2h3HqcHJmWpOc9MMzvzhp1ZXoDLdgFLTOWqZSHtcXwHjsMhERSyvxUEiZffSn
vaJ/xmoTm/PFOgwV5kwGgkCH7NzeYHU2Pp4MXxzOo+8v5i5Db+reKE7MrxKAXW41
UrrBJLjFNN9Q8PJ7fRZE2r1XGLtcrco6zrGlF5ER6uyuQhXIFUqo4Rg1QnmoxWjs
D2Znb7DV5NaAVf6SuQu2r/74xbLcHvxEI2PU/veupF/o4PQ6/aAA8SE9277OT17m
5/3m97zv1t7Bja9Cz656LF+O5oYsP5E1HcL4Mcu+iwI/vjhx47jPiylA22XEGU0P
V7Yhb855r2RDRs8y6sfwADxtoM3IQz8r8DWTKYLR0WwQ9oGNtD9B0CfViCUE64N+
A//ty5ftjiI8ammdQInqNHHEEn2UFovHbupbxf76YSjVK+C7atRzHS20vSw/PLFr
/4G7BMBUxFnGkvW4V5YkBwT2mBSfrbQKaneW1NwgZxawCK/jQjt7OrW9mmE4RdhM
yOONm2Tsmni7Vz7O6Re+kEOpRoFoTACxwKgpNxBiVYRaZhAmkMNYp6OBvDfxEq9+
NK2nczG/tPHKkXCkK/HJN8REBtj+IuYV7ARbHWpY0ovES+RHaX4wy8f49yIbVSVU
8SdBImLCaFZR8p2EO+ODRNXsA5GzYsBeD1YN9hrMo/OP1JiRtLAX9r7XQy8AsU7a
t2FQk62qDHqbTKU8niH/K+9AQXJINFFuYv+5Vx3Spnog2HBEv0oFxIuBCAYt7dU1
UVaqRCCUwlFoau6Ypsa0esipPevf4pN9Ds4qfOJMAJc2SX3mdgD9vp+y82bcrbjs
G4aarnDJJqcPYLVsmNKpAA2hlSQRLdR/D3SLusXlG65g0x3mR/27iWT6fzuBETM7
Jse4FhfrYCDPfRQvHEWCDX6ZaSTraFDmyqVaD5DxAj/ByY/x2mYCkYTtx+A/eOO8
O5fwPCGn0DljOgP1/+p9WeATVnlvzzs/JupEWIPIiqf10E3422U05UX5rQJSYdkn
jiUPFkygB97nKWLNDig1IXiK4HZvCaJRCJzrzUhD4rS25Z6j9v7LYdZWnbgx+6fR
XyWFUaHQUXrc2+hudm7wlJQZ9DnHmLtH2JFxVtAI7wMBrKEntkW8PCKkSZCM0uiz
R6TzxcpJ/KXjVscjugwst7kN2KB1s5JkZAASmGTeesD696fIPSAEctRfRYyG+gNe
zuyUCjAxM0OALtngyLFw/OMfdcrDka7/1uXlzfrSFJm8SSH52tePVS6iSZgvgRjY
a2GK+zTamrY00+AdZYLCbDZvEku0lITDgq72Qa0cwvy1SKLTDQUHV7mVPLGneGe/
MehjrPUpT9BJ//tINZano4NUA6mMfqr2dboFPY6+Me4c5Bd7RuWLLTSzAGFZpwYB
xlFPrjy9JLaugNb0mZtZTHKm0s9YXY68h4f2q7KHIXDGHWucnINDx1+jskKr3XT0
vPTqQaj9dbztWuNLMTie03W4fI9o5PpPArWVyiTR+lQfI0g6msG0NgY8oPqBZexM
16NFjQtXnMlIJ0bXbTzrtXr+E+h2A3EkQIr08zLPsWWDNiYq2xYdwWUHYDcTGlZd
BGog5EvBqMSTL1XuwbdsuKWJxf9ru64zVk6rsSyxFMeUhnI1T71K0l8cTNGlHsvF
eumrXBkvi1Ai/bl3+ZlmTctUxXBkrBvotxECnUAGdDcPovfBy6/XmbSIyQ8/aFpj
3Km7wiNQbV5+JFMcMdYRltC2GgFWUDm8wAZ+T6aTGF3qZ83lhojehuQPtPQvH3dy
VNOVAmfPc9dr8E+6elOISPt9o365sOhRxY6F+nTe9z1s+iEgZ2M51TeMdKp4vaMQ
31+PHOVtySWgBHfAuAzzjPQr+lmjasUpUArVe6mY+FbvMiEnwH+KB2ykr8ts2N+U
bq/uCErMnCim/8F2kjmKNadpQV4JGv7VkcZZPEEXNwvJgongHUg2MUDF979h5ZrC
tQg2/zzLtkG6xZCe+4JF1n8KcBdK4rDclusOkIvGdxnFw0kGiZhemywHjUU8V0YY
4RuFNJpf4ytwPIx90C/Wz7AK0zKBpET0weCRE/8y84uE1OFhhkI2PoycqsMBVoXz
b0AMmBVX7ke93ow90Ew1/5ek5sBRSMT26kzlyQvEXq8GXgs0qJxDEAlGdGa/P9x9
RzuV2i4EaKuSYorQ8AZqFAUbxMGgRii2zkv++b+T8cVJW1kdQnl4LNXAHlx8MgnL
iQITPaQa1IC4gU0J1aePtgTy0QOufKKWhDuGpEuIp3aNg2acmtcbniMwsw0of9L+
a2J08wWXAz4Tt78mH5gQD6Z+xOlw09wFK2CYnwTNe/w1Q4Vpeer/UtQlO/hGKuAP
5Xq52D+OdlH9ZsPJRMMOMLYkKl9BjuHRGFpRRAcGB1g5t3geaPqYk1rFbi1zUsbc
B6lDSV1HSF3H2/ptk6ppbuHAF6fpCbBc2nRLhiRcOmf/w4mWTjzd+gkr538FknXl
O+8jRh5LfBaUF2wXKGHXg4jfLqDOTcDBDylqaBgMBFSA5qNLq6+dut8RnlRuelq3
27BhQ2Q4vIiawI3gouVbCiXszyD1En60vf9CwW2CwDOujabW6EDLMqNbnAR7HP2l
dHgKQ2cSsXuyghUjF4nRYSdaUPABGEhicbQ+VsW+an5rOwUPqr39HuisPUeKt47f
tVxuGDjVXDlgZLi5VLmzOKsEYNdBpTxJ97bzGIa1yaWxO71CJBvhd21MktKvDCwr
gJl33GnWb1SMcTDn31XqnHL4i8HQ2S6/+fBjOjsdobHEzKz/YsJG6snYixHqw6QS
V3EyFvYkbtcoXg6noKumVS5/4IQzRlyP1ZkVgq4hLGMblCiahoCDfUeKJ/BvajPd
F9S+NxNyjEBukiy+UJFJy6W7PhQEWp7VcHYN62jnGkcx+QlxHs3GnpgQOFLbf7MG
ouF0BLSWt1po53+StfuUA9cMuEQizlFn5Ebd+4DSI4fane5EZjbWmOpLnQ7qYKpc
qjxEe2EvrAYJepMiamgMVlw/VplTvGdrl5tA1zvKpo7bwfg5MBsHOKMLLGyajmua
eLZTVO+/PS12JaiP0CUNOk3nK2JkjMebGvow5UqK3ZGAVLHq7eRk/zvaWsNo6OZG
BoOG1upgyMl6i6kBhlzBeBix6T/SE0ikxlr7UR/4RKguw0hIPbahgDgcW09TvI6T
5avoE/drxDSMWm1y943VvOKUVEkY9EdpXTH1SFsQqXR5B9vilIBrX1BGdg4t9DiF
CKHhxFk1IhNOlyJm9dJ+qYQWIiEsd+JC0jEEYeRuQxzbKFM9svPWenVXPICI+mqX
17Y47R08e4sf3El7Ga+UarbOHrT8k9tnCykYarIpa/TYTjqv846XFl76bKpOevxp
WHOTO/77w25E/42WkhWSuDIElCdaFDP/lt/8a5no7boDVZ2tevuYWqzHZZuybk7c
fAGshb7Yq1bmLNY1Ru+5kEdUN/WPzvHItIt03/7WEPJTVJ2QPK75dxdV4ZZeqsvd
noCDTL63D0CrDrkpsvPnRcShdsBkOaxWVUYFOWfs66EtUklSsJvNZZoXODZwHlfl
oSzCU7fWBFIB+sO7ZGSbDDIqDH49uLLkMp4nyrwnRHaP09vA9vicgodjKqHjauJb
zhq4uk8R0Pa0sQ9/+Yn30xGnfZembvrCL9YJYedBljXKCUgBpC+EGeztlekYcVlu
j8nPkPZ3v9tm6F61xMx0LGw50z8KWn5vEnyAK+UbWG7gkSfn2jlkUxWtv/00jNQ9
gyEcge4eBuCgxWMB7NN0oqjWNIQI8yHa6EqDzsgfLCa80JqEgs04yUnkRkb5CUC7
Krni6XtaAZqXsHiuFpuOzw1g5+D61Nz+e0KRclYfdRL0Gy8dUZu3D2m/QtECfyb2
YJ/t0Kxcgju6wjI6XemFG4a4xNC1c37KlbBaZAMajsCkhnhEqkUZg4Gf3sSuI32C
FOEXmRGCEN+ch163xDVFI4TApJWyPj77uTj94LHXCJKk2lGaonKyM3OdxodipSOj
fh13nUBTLWsEQRNLFEhbmkQ2M2EaAi/hxZAWJ/3JSkAg1En3XUCRph00gRc4f7zF
B8bVNNrxU4EcohZN6aAeUpgGqR3mCWC1NjE79SzckigRxV5ofZrq9buwPx6L06+t
R146dVqLThXhTnRhsHifW3pvOHobtXTM+j6iFqez3xplqRoOf44J565r6xxMF6Al
vbFzawOR8FMpaPV1Jau/98OXBM9UsCxRsUho8VSdEymRwDDCAsEQ70cEaJvwPbPk
3piLepo+ZH2X4QPMAH3k+cTLWJCyj42vyxGhXshes/Jh+AAZoIeevz3qsbQsE8gi
ijzG3QIiAXOzcTmNZDJcUTMR98uLBVL4ZF6ig7ZzoeHPYvbZgFHjXg0E0vGcIbWY
Rg+M+aWU2JsfrzWY9AtNJKFeCwSp1C815o7aNoRxQLewK1ehUYAlEjSGIL0RXiT4
M4m22S2JSOIkmL7I7WQAIviOgmxUiCoFA0+Wn5L7fX/HzxCDXU/l0gOfHCFMWUjn
ANey4XNKYO3NnQS8An+8Dc/2ioaK57IaMAJwl5osAzGIXwWnxkt3SNtNyTFWDZmk
0/hAeVxBvJ26I04C02OIfUA7MYCnttYCjcG8uV2HnWd0XK9cx+Gn9wJfM+CtSUXU
4IJhUCqva42sOoMxHaeoxPgKSp77VHg3ZSP8n6ZJtmbq1GWXN+cdupIYMQ37JrPO
VC24Xu+to+F341U7zNAFbqxke04XheIfDxd4ZY4ABDvoL1W24bksHctLMBBA8hxW
Rdrx05OOT6gSAz/VyofEnORCsBTlGT0e+ZDg1sud8QGhGZEf9a7mjnqAO79ETwDV
Wd5D2KpbU5x/xVx3Ns8BV6hcgoQnXEQxek0LQv6+pMnFSnPI2n0Dp9kbW4Oi+djC
07ttOB2Hh6WzmRp80p7cQFyFiI217jhsiozb6cBtbqVF4y0MD+CjdGLg7dqN09YY
vQ9MkQ5QSJz0cZtxl47JNNioC4ti8swDuDObIXPC69gUPIdsMXDs3CK6S25xY7aY
7u92Zan798LMaFga8wBvaU/iyHWu7O2mBr4RFIRuCtlLQImnYqEDFCaDPrnKaZb+
nSB/JGuCmlCQhAUqYlAbxQwepYr8CUu9QIl6ppFMqo5oRS4z0yoIQ2ILXclwKjeQ
x4F0ENSzM/4V0DtlI2Ix7u5n6yZYwoGKevhK0+70SaXGpm2AHWOUEV5nhkL/j/lz
UFXdmVp3rF9EsZKAdMjLH71sc+G/JqsSIKawUFTTnz2qLcg7LTojnj72+9Sx1+v5
gOlsKKiAMeK/7ryaIJpIkdQigqbAqDoQPOhGju1NUETBo9GW43zsWL+CMKDOJQHt
t4o/1uZHfsgh9b0MWt6slf34mtjGdmU1icpKG0Mv1POwTmo6w93C6RoqqeA05St2
KkHlRlYxI1q1Cbpg7GatORJRCwPXFKqW70U0NSvSkDIq+LpsQI9FC/rTIdMWtupr
yHmWMY/FBu4rzO2By1Pm1mac7agr4+bzt0P0xZZF+zUggAbA75Lhsa1Kns7bLWVF
bh733wn0lCR0S7TLmzbLOpFY9DwvaX6d/uAcLQbfvEHiMHCCIb1JrRITr+WfpZpL
DqsQlFSh6w+XaLzKahtScHDPGcAyPZAztlfJohAHegsvPcTC4cgu2UG+BhsxO8SM
XSEvKyhP9vn9wEgy2m7l9E3+UEHz72yN0Ylel83ByzkNPlrxvvswJHDdqsJNtFDV
gs6uwavq1kT7ltDONSuv1o2Ba9j8Fd0Uo1GCfWdUZ9Sr7duYYSQHmui1Ndzgur6T
KWPBPo5pqocOxtjgFG9UHvLMkfnywu+FMNw9jLcINCM5hX/YfpioLbgoOgk/Z0pL
B6ip2jgOP2tlbJfR12YqN1RoOCFwGjqb5NiVWZDUjaNAGoJ7yNZNi6HiXUq9YJBT
/1fdut8E+EgrbJtFRWI8xPR+uSXrvJpeD3URab7kivA74R+ny/P4jmNmo342PvSf
0ilCsnOFkGLc6skAXz22X39MsfskhHsyaiKykSOBMNzcAFK07cYdAEZe5/uJ+MnJ
6mPK26//r6bcbjB5N31Q+sKDxSDYDx6PSTaU6SEpFJ4D0DIPg8MSTypkhRA6t6E0
L3cLliTHIxpiaIvOWfmpea2NMD40xvMo1M2XSVVmVqH2lwarQ6X/sTf6/fgbfCXI
XAINo1aJ0iC5/Yg8MevEf03n/1iJhtvHXRlTiwOPhjHkqqOUPAMm1IZYB35SM8w4
JiZOR4y7oMiOcV7v8qShLFyLMkNRVSHTHl1jQyvQOjWeFG4gMjcNyBNUpCGyqxiO
MSPiwD8zU+72G3UGtXmfLWjmU0JNOOq8B2uthKY1HYgqqHEBAVqv+d0ZSJPHT8jc
SKmN5JrZeHg+LRiGroDixAMRN0bd1Wsrp46zygER4XfxcKcTi93ZctpSHtWrD0Xr
Iv6rQPgxH+C93xGzPrr4pyX2uH8DEAc2C38N6Vr3Ox/rG18DMo4AInxvKxLAHmac
wVc2N/Ay1L74V1zsepBruUz1bS3GZ8F30QUBPDPGNMElGaS4TbsstC+CpDWtC/xg
1kOEhCK5piANvC6kIy6R2/9lP63pPtAF0oIb/NFJzM3H/xS7nvnw5uXEW3Ps+2Bu
Wx1ZFClN4kUbXvxUeb1DX/xMSOHRtwWcc9JtpAAk7F8g76ITYY4dsAdbRywwoz8c
1qd29ju+A1VgEw/CWpWgvXOHf1bT9JOS58NEfQ2NmTd9NpPZBF4w7n0Zvsi9orPl
U+jEPcXX24dBFyYt9g366SKYPvAEH+Zvfq7N9ovXKU55tB0YTYPdIFmh9AoRZjOZ
+0L4EiMoDoY8G8nVEajEsEcjMezRl75k1Z6ruR30s/8+IrFhsS5zBfCkM2lqgk2p
MkMaIYNodEE4Johcza2pSlIisAuY0J9YwjzhtzteJaDqmcIQSGK72W6sFp6ZxQ5U
KZplXebDsFWUisigaAvm8SRiKmOo0lMgKlkJps79+wcSoQzEzEdS6C0JDJ1Efp7j
CKx1ABYZCgcSPo84A1iwW6sFQuieN5EXLWP0VuEeNxx5JMXskz5RmaT4zSBJiNyr
uWUDcInvCE9oQJULMIDj2kmY44HR/pLvzmQrSlmH1xMgw+ogeLGLuZ7molBW9/Yj
5w0Ow4trZynOEsfMeM1d0r3Mbn/o1wQI01unKptb/U59Z/ggm3GQMlZA+5kgqrhE
62QMorOyvNtzX8R58jde5WIIjRh2TtVD7P3oBV5gkCXmQZn8NWNEFUfVgwKXBU87
lZRDvM+I4M+ca6eTycCwKQdM2Zk4gYrKyosrJgWv1GORZ3c/vkZm4c8npqNv1urn
5GaSvzSwnE4YS4g4gnNALAqxCmmhTuRIE02p0Dh5t67aKqQHiljCfjaBbAK2HLRY
fAZuz7zhqftgZg7jXVRAknMjqS0h3Do5UOasr/GIOf/LqZQe/RPGIR+y+IG2GjI8
nqQ5+rEPSXbet+SQZH8UFLOn5/dE3U8vVHqUlceI/Jmaqm+y94/8A7BD5PxLq8Ib
kcdlO22250lCLplzWlIMEprEs7Z73OENeHo3fYmqJR4wL+Zq1DsQKQ41Ah+IFAAs
EFOP55dBZ3zgQZmTEsZgtHyg56pNoX1OFcq6yn9vLmuvTn7EFewznoi2ZYO88aWn
Rmc13gzFTUHb3MTfOxUgBJPEpq4omRKR/ttqFAJDj7l6SyYqnDV2TgFPphbG9FK2
5XvnCXY0RD6TPSVQFBAnbpN+BR2adN0dOOnRjvEz73BXeep+nPJqNG0ps+Wc01kK
zf1jk6Htnj2O9aIM74s5GShIXy/fmnLVgi/lyLln41yVQfICrtbkJvDmxDrDJt9V
pCHfFOVUOibNrcBmztAGB7L2LOxwLRHcy/y+RCiuKglKBOhNDsVlxlnpT/nYdHdi
5HV7X2vb+0jsVcEfuAoOEKMLTMwQTfCjQzC3WCapowrHzJ5PfmXYMr599AWpdfHR
uMSNUTN01/URpdKrO/0Ac3rKm4T5lz0M9nVF+oqnQAEmbanK8VbTK0SJtKVsO3kQ
QJMJ1y4yU1noLX/XFWpCViXpvSJxU6x2njYaYNlJciCiMKPilgsqbHEwmVqpZ3KC
ZaGzKojv/y3xwWjIpMGFBB4iNnAi18UbX7nu0Dif0VjNv8VWOm0fsXs35jLl8jJk
l8TNNkYVN9VeRj/6PRIpjmL4+m9HZ0F3azOG4neSzkrN+G/dqTeq3AuTCim4Sd5o
l9OZKXBcI7k/JDXTidNjGM9iOInBG4jjKAOcxA6zaN6CQqKwCjI3V0Ts1XhyY5ze
xaw+ZJQ5HP7h9uyV1VD2OMHZU30OAcwqHLWZ0uvUeAQYkAE5GfPwJVmXW+4dlxkI
bswCWCcWMTsKwea923kjtyU8Nhv0k9wOYAhr3Z0OLsFm8c1UENRijCrEQzpEvXrH
PElasT8L+8xQrGA7aiJW30Xkxo6MGvsIl7UBHJ/8cX9keJtJzbL58SqVnjh3QxkL
POp9wVCdN3xd7Amco+iA8lONL7cMFpu7z67zMISejZJNX3xD8fcDKsgqdM5sBMWy
Bl/5GbRAh1lGDK1Kh0YWM+ItGgs1v+8v1yaO2GOG9herfBAhsZlmJhGY85BjTL2w
IAj9U1aQThe5No8aupY94VAH+GxDT02E3hUxdkoNgJYl/3euXbeEz9DkHbaGLvoS
+1VcPOBU4OmtkBPjF9johrIaiNEGAksO5/ukI3LWN8HQ/prP37gu66+oMRTijIkC
aQXO46RtiKXBSm8E4FuPChuqs/0AoNzaCgbcV57+6bskWISSKxcsAqu5WVU24A5L
8BDd80f/51Oj3UGb92GBGd4SKx6pag162XgrxxMgVMUs15OfogzOTOKubwe6Eyfv
SeY56aPVQPcf0g1kwpuKx14NpTnKRn4ED/qvY42tGygxelvSI3V6zFY/gzAkp7xZ
8qfUtlVLMYUUvKPtOCnyWdmugF4v7zxLDNkqqHp6btPG3+oq+PW8SQaUyqfcMfZY
6KXHkTGe8veP8/lgHHigfr+qz1vZ5UDixs1JJocQ94E1EejhkI39iYR+TYmdoPMj
RIVVBVKfUmC7jOYfKcLODPI9oXCPNhdNN+Pe23NZrBieDS9rrEz2Hv5AlJmGLbuI
ITAWg/Am/HQXDNOJ++8mNjcbUbkQDwiZeNZMiXP937l+sagQ9DrkaUZRU3lPLKmW
OulZOVHyrE4gZHNHIIaEMYmug/oDIEjzCdn1G5siRjW/k1zEC4qWTq4HPyKz+Qqj
IdEg9001VxUIIgYTBIpQ9L//FJeHh56a37EWh0Wcge7LZP+n3p6lb32jPkJJ6+gm
UY5Dyr09cLNKdzx5c23AHDaqrN2mhJJEdjQ7A3U8utgLl08WQ9mcX0CTKacpxlTO
+NXRHrnDDx/nLrUsQ4xXzBXx0ksYh31v0JqlpCoxnJtrAr0droYT4gDn9GCn6L3u
hS7nQyXQFWFM48C8P7yazOZXij1yD2NH3TRBIFitw9DlO2o57mgR/2h03h15TPjZ
apRgMM/vOC4qjferB3oP+UUHj5z+yCKFhj3xVrocgT39B7Si/g/Xkfv24wnsnqQz
V28v7/KAbKt3gRs6FhlWt2nFhpBHFEhfpxlVNl9BKObYsyTVO10C4FZZaHBVmSBg
8IBbsGYIuyybF/UtF+yr7opsE2x6LPPoZ6cfHkFoQPRvPUt5Vvyf6wPkgoFSvQGQ
hDs3hWl0wHVsTuxEBa1ORix0bAQwUL6UHDH9DcM7olefRkYbiWzyWldKPPaoG9Am
RKqVgCF5nZMsujWJ0ZDgYdLCG5DNCSCmAP5IBOOtQZ8VJhjPxiEQ7qC7dXlOwOdQ
ePPfXJBu9gEzJ0dIgl7yrRBJbF3wrPP8z+jD/clepptrPrTTitnTHdutTezFbd9Q
GSMt79WuDw2xfiLffRV3HqZWvczAlTL8NZX5qVaajUnlleB4ZEG7NOQO/36cux68
5cH26RkNj5k4b1qoaxtKbpG+Out7Vn5vLGXgR7gkDRr29aB5oFfEQ17uBce6iNDJ
UaTbhHbAxXh3l9/vDU+MhY9wRGEf3m6RyJn6nYcsbW0YFxphmlgSSsfNj1J6AvKx
nvqkGy2ZT6QHQEajbR2c7851V9qU2mGlVl9rwG4x3DbkDmlWRUTkb2r64UV1FFaG
P/8fe+GTzoq6N4ir1VGdsRYgB+zDT0DtqU4MDLw7Xxs+dj5UwY16GEz48neMczBz
UeOubm6jmGFj9LepKnlOTDWg6eCOe51cki/Iuhw/E8U2qiXecSt9sAuuC5yqVwuf
ALUPr90jOVFdrITWpsZstPKmyj6ERhYuX/yHwYTZ0Y9OINCKoW7Rcp803QXmoD+c
1N0OF7+r0IPgPvJ01jbe64vyO5NE8SXxP3LaJbRgBlGvNzH+eBG1m62V43VKjp3B
SZ1kjw4MOXDowVy95kUOrtcIKVXV98MM1OJ4SPzj0vgVM/HkkQlT0ckqjGLXLmlu
4vlFDoVzQ176K7DUFEn8AJMfitZYve5xffLQVIR67hf1J5ytxoTrA2s7wYCuflYt
A8aBGxK82LMgNpxcIVK/baDEN0B+fAqfIYKTwec+h5Kbf1udnYV8MMspvgrfFHea
ava9rs7HRDHseWTZN7AFdqUF1sbtA9fJ/eFdnxGGCj45DNTo7aPQM+50/60UHRjO
hTHbpuWU1UqEGV2lGoCx3gtdpJeh5j/0oDIvz1sdLwmCWNzvoW23HIFybSJ1SP/l
SfiJzXx0X1fyH0ECCsH0iewkqCs3HTYZ9JQSNnp9+/Cq+aD/0DD47pjc0X8hGBbO
+gzcFTnBRLLW4e+Ko4WZKhlsDfBW6zl0hluw9TcAB+TnWfxvdCg7F2RloTXi+/oh
X85tiD1zs3XvpFgYOWVv3fxYbdkd03cMsItjKztpFzwc3uuFiF6aHxJcWEhxSc3b
BwGultg/Y0F2AON9ekA8t/ymFMPAKIY20Hn7GEO97kTlb9Prp0yikZqPp47C0WNS
gPbPSrNZ3krg0FGRQiBZlqL+gZ8w0vBoFwvAAHE0eMsN4+c2jEa35EShFHQ5IUql
YzJjelxeLqDt/FOGKeecdTXHcOStopwDPqlgCrw7c8kz7MPWnIGakw8SoATZd6ak
v0+iIxF+kE++WZRRYlGpeIp/mgmrP/tPaFgjCQpLGZ7krhQ79j5B8LIPuONcjCKe
Ed51INU/VmQjeoDRBdbSLPrEoaQwx6BI22c5kjaCHaW/F8I/1CIEpYlmEsFKjAa9
+/eNB7s1e00/+azmwqoFtE8+tHwwAZPSVnh4oAx+PdRv5soV12JEg9tEdmYZ6gOB
Blq/sEDCisjKLzTOocadpxOaNuRN5D/Fh4hsdGtx3ybmRJqVsH0xUzFiMgsS00gX
umGz70X9stRxNETqiF5ZI4B0J7PhTDOEaZnuzN1NSkTY2A9lqX7aNwe4CCGQzhKR
msG9tTLem73Zmy4NHwbkItVqL/luOTzzh1qabM5T/JdcqByQbzPViMxE7jafM+f1
VzxpemIXGV5veTyeyJj1oaU0ClO5pqTnnz9K5tWanpq+lmoW4gTNPciYFcMrQVa+
1L4fyUUEjSFNn6eFmd9adaRy0LAKQ7f9BOsI6ZPaJtvjdBzOxNbMyzwyDvo8bYUK
FMir6wnU+ZvaPKakYTHITGzVuJkFD6VWkDiehP0XaId/D95iapyVmZpg6vxKr0zz
eB7d19ulh2fXXbbwj2LICG1ykIpXEQFm9esWfhuh1YvKJEQN1ANNLRq6Px2phLOT
0giSE0XuhzHiIWklCkOx6Rli2vPMH6+SF8xg3ub9gSYWM2kzMIG8a3rxOsysTIfe
psyWGduJOAnqcOUg39Ti+sSl/X0PnJ1WeV8hj6km0u2DypylmGkxtH0bhTMtBqm7
zAVczp+KiY80vieGgCHlfyLuhpHVDX6LE0hg3+gMwCvEUJrgmudLH9Tuh/z8dSv6
ZB7HbpMLYpZF4qJemg/EqTqm0T8BkLI1uatx7Q6v3N1L1dkx1TL484as/M2z6Yfc
6Zfndr+VztowUGR8cPEPCpZ2O3IGkpJ0WCMVkbsIQEbC4mIo/PwFuEE/obRQ0HIV
0iBSU2BQK0+bAOwZ2qYqN7ZXQpBKr5b3Uv0Jp+1d921KXEF1c/C0HWvF6C8Z6ytE
uuOGk3v41OdwCGBoseynFA5xLWFJ8fxnTHomLH0aPpZ11ffnoq1JpbGj6EAVA2sK
Z/DaNIdoee/qyILqELi1gr4fY46wMKjWELe1WnWBfGcS8SHdUhgYgzwMQE+nNk2m
bLTuWB1zTaBDCmNpYx14uXTrZdn9okbAJCPHe80dhLuJAraSQqssKDdVqPRYWTNI
PK5tUnT2uN88peZ7a8mBfedl8lWf2KnWQBB26wtyKyqWABs3lHopNKVCbsbo7n3w
bEY93mD9EFf3z9ygRsaJ3tyzpDqhKfOC1mL3EVdiv43EK16AJcULEF7ng+N49sZq
9rT1udcAre+vlPISBGq54domJQp5R5NdA6AqqZFFcK4TNuqVpJJ+WyxKFT0MfgxD
9yUjA5qgk3eVXZ8VJqe98jyRUq5eVt02iJUNtgcJEp/pheJxyD+rChhJLIcWjmWN
5IV4E8dRpUjBhQvJoXK9ya9fCBlQvsRAequUgSPsDNpxY09wXU8POtmP8O/j474S
rEOuZy31KlDEDveQLD02ZGUXVZ72cBZ98iYC4PyTsQWFQfAu0Cch5Wgq/1NdBPCF
HrKaXLwhldzKgp4aR7UsZ1trV/0+aILzQnXlICmsPH0VDOTrIywB9dIhvIAr9J5z
n0gQW5WgJtNeZIaZjXTX84qJPzN9ze+Kpcg3aCCU+VvT4eJsewyQ/8lcrBw443/8
PGkzHebHpy50Ix5O6MrE7wKbwU7CT/UyaeBwwPLcnslcLcnShMs72eD32TGzW1yP
eywyB3PzaqoMTntUHS3WouCdRi7W/8lifZlkSz7qw2DBccEqRv3JMxNbtRMH44nm
M4FxCKRkkfB4y0bnUgNI3hJqZBV5d8tOGLb/Xb2wMjHK0Vuoqm3kiP4XthM5d75f
1raTlv9+h2FOhmGKWnXX/Tswrzz9TcYd9J1wu5ClLURRhr6gr461mqtFn27IKIIs
qDWfcCSWgB6JpH81WDAqFHQ4TMVhcrD2OOYdmuUkA/gEB9JAnkHcexnPgKdhtzL6
mAKRgShSpPT9Cx8S+7ofwgBesnpfcLFyfnHJ8QIrQ4RFbpjADhtXqaCf65YIJNrQ
fBigfM79RVRkye5DaHu0OFAGurjsw5dDY3ohYG7+JNcbdfAlUodBCWUhQ7P6ZQvH
9h2NVCoEPrd9Cge1IAFU5xCdOtn9MoXYA+pDknuU1HpO0IhamMbxbLuDaAXwS9Kz
c3mjkvFIts7i83ogjFuu6x4HZaADnX/GIqx8bcgICWTFO8Wt4Y60PpVylIV1J3Sp
avGdEtjZUG3y4Psvv3+Y+pSx4ZfjDRe5AzX1P46VzxMi0O7YIfNB2awVwZExNRe6
aTaP9/O4Y6zVtc3qz1HYKCOAe6/qF6+mrs0iUtqPevuAhA03EOL6/EBmnRfnjH7T
eOqyG1iKaGKvCkknkvAW1rtijsbNlTV+q6zIB9mVVpNtWPzfWMpNreFhjowtLZEY
kClNZWsw0wD31alWDkrkShtYe9ymxug0/E9uR5PcF0v/poSyP0YFLEY+vZ0RuLlk
tUo8Mb5QmEm/ZVsV3cQY5Bg5dkI2xrTq3v2680B41p4CX51av4EM3jLxC3hoWRVj
tizLdQywAEcTkbsphsQUmpoejRP36axOZiDWDyPcYsj4ZEM6pruVoI6JOrxjPDgi
o99PLqkKY+Kcl0fK/rcFymGSlSjzcZLFfhMye84MAVNKImpPHcUkO91UD8Utp9Jm
B64Um2NFhN7a1NVT8y8APGWJa1gkVwXY4mQRZjH5R3U2rFf5M89qS45Sj0pKxQf8
Y/EruwlAhAICdulbcXCUFa3++SP3exS4JsfR0gkBIG1pPGDfEMrDjWhYUbw6SVC1
2KjHdDissrxrc1GmMKTwZ3dlmvwdHAjLczZXlGQO53eWzNXXiIpNpKm3bj0MIOqj
Mahk5nkqkfQNEWOtdMyWt89S5lAW3cGx5x7a+odd2L4FRAzGQbBsrBz6+qTvfZrG
A6wNuDC5hvq7CYnBjih1MibPAwrUkehHNDSLKAuDHaIOpav9WnsPb8DYXmViPANH
fwwE6Q/qmADzxFHTuczioxYV7jSr4GM4hRpbmWjZXszn7w6IBDk1TK1wjoAIecho
YcBsKjp3jRqq4Fb8v6ydycyQzpkiRMFIQD90U47s5tmd2Qtux9GlBRayTYMxe3EI
PhRvMCeP+ydz3D2wkvREyt3LexRy6/edqRlPtYvfcZ87ZD1Jdb/pKsTFI4iOrabB
e3FsjYnYq09mcscUc5V+Fmr5tNVc6/o7G51KW3Pm91TjVCWq11U1QKi8G0/6In7V
2a6hwcUQ04YZAGfS5X9ja5RogGd6jf7GdJX6H10mcdsP/SS3HoA82pZaqhMevdNe
dEkj/7cKfDWeoq3EnQgPlZ/sQgBczpCFIror+nhMblbBNZo5CKtiuPlcaujncPyD
3Uk6kUseuDx0UQ4PITsM4rGzcMTslUuWr1FROJH4JyyIoXH28hkgbvPSMmYodeS2
11Zsbw4Q/RWBInkjimfOMWY5X8gLbbi4EmM8ZrPZqD/XKXIYBJHIny5poSMEsTrT
aIWybKZQk4WNYKuaoP6KBZn3nvikBdnRFNWOi+8wZuPPzmxCmv+uWDWQ15qbbVRz
0pRIhaisrnvOvaKsE7u9dAP4vcaTL5nO3r91813sTLGPFXar6btZV5sW31kkiuk7
lEqAjgYovNqd4AfV6a2iXVaaJQfmhYGR8Qv6uY6/EKyuNeWZFQRIZKaON96UCW/B
O8ba6jg70KUHqXWkMNffdKHpOm4ms3uGCCQyvL4tih8bTcVk9ZYyTy2BJU1AjBmT
LOE/JEb7u2IqfhQSvqZF39LNvwNxDnhCCbBzMm20fOcaDCFABohFrOhHLhWQ1hDk
Ph/2x4EmMJqDSU1TtaniEL2zpm4Tf1vXIssb05Jf5o4v8wTVlihLO/Ygta78YOTS
mzLRbwJ336+1u1BrhWLgXP3abY7C+wi0W4DLANrrJgSHkmpzlyOu/ytNzJwxTEgp
D3ImEQR+gqSvozWXe+EgSmOkl82HaEq9ZxpcId/fGP38cCFFI29B25b1vAu1Qn/2
zKLqJEAvrYAKkfcqqPlWEhqW54aLiHv7CbPtkyurrFq+zj5UfF0Oj7ITwT+aWfPT
KLp4J7bhPpeM6ev4wLIDLoUxvsKi0z0oUGZg9nyWQC4pEThjz8O1GHvNCOTmVk+9
AjrSflH1iXke/TUoBPNNIjBt1+r8Ukox7g1qTUaqfDuDIwWy5387u57JPohghzyX
QtRzcieCuSZt9+pCcpiotNPHnXEpjngvHX+YRffW9aHmcK8FsPIG48jhEGEOBbvX
2EoYOIFMVwOLMIKUEpA/K5x6f0XMza1Ji9XvKHLN8DgUk9D+scFkRA6XQhcXHYdD
Ge5OXGtrxNk2w74Stfl2r+jCGzH+kN+rwH+nLJiJjRAsb/hvyjO5omMVMONAiMwf
FTId5Ef8nM5iio6P7HOiZNCLPlDYRrpLFtoozgjKCW12LUssmnrXs7HuTEsw05yj
SYDuyxIQYgseZZjCzrd++z3IQF69Xm6xBl3PjPg04c1KSGvSDcb/g+qizo+X95xI
8nPkm1ChMeLO15/8wkmDHuLkCMH3nZckg6nZvezy/ss+SxMDut39svEBCRgvvaCC
C3tOCjgLf4Jtsv5G5y8YxT5NqD9nN8N1MSTM6IJxwkXbTiREH/C16lWScNOXSQ5K
8QeHuQsomiI1vF68Rqn/MivV+W8EtWMi4e3GlIJk4F5N/S5DGLy7IsJ4iRrNsLSG
YpYFEHVDGqwQugAf8nJoD+Y9kTe8cwx0+BomBEW7uQ0oJCZepqHKRToPR1zUj0P+
rfslRgSu4+igMi/tGfYqE/imHhtPTvfWR0TUNjhqiBerNP8FQRB8JgV5quOJ07aO
F7JuHhBHw49UQX2XAnd2V2fetEZhGn72Vx3NT6q/Yt3T49Y1NJdTILXijbCADmHf
0EvvqETwjdhMfBk2eJKY6ZOYI7XNtyB7HE2A2CoiL81n/CLVWrgew2dzzpJKZ1Rr
0gdygRCg2+bOzDLqqYVaVA4CzISPdTPW1zBMZd+qPkD3ufig2bHLZnC428pZVr4v
FMV5HdrOXZPlblEjY7+RquYTnsV/UYzY4IdvNGWiBEBFnwCaEI0OzqvCT45JH35O
tZzEeYs4oRH0aAxm/WLYdW+MwU5SG4SeW/Jv2/zOOsU1LdMFUKoqlRqtZf3sWLlu
xAgID5QOY75VM6SgiwqURiPI4Vkt3xPkIVMIonKeRAG3dZUO4AEsaudMxAdwAm8C
CwVCI74SHa4jaAQ2xOBrVSL+EiO8kERiKqe4eUiCxRqdnDbB8hi+yI6w7iR8F1f7
DWR/26QfXnBm1pCtVs2AQzYvxfkA0jKCU924d9nExuVxwwruJq3tJMegJ1Voemlj
TRS2V1y/2HqIf5pEjsXa6u+du9nT2xU/9UgLEQltlHr+co0ALdwoixZFEXBtg3fx
rHQGRqRSPgF3FFxzIkchrFc5LyugsfPKHIvsI8+woYtHo+JUMKCHIjCA41QOnZZS
DqIK2HCq5yFezHZOhW+1uUflqKedJ/nPCUttxrjA+0n0tWiUYt2Qjsf0WEXs+V0v
42we8vHgF67ziATnwC/IV91sWsViHu15J82qtGmLXEPygBYsWYhFocCTo4HO5Ps0
epsXcrIcS9U1DAqUHEb2N670TVYOFtKbcJABNd6HB81xSmkXoRkGR3r+A69Z5nAv
Tm5nfEzjriSRXKx7AHvQ9aQ8ELhqGKd5H+KG66e9lJrpu31ZGzkuQR6+QWHuF+tV
8VX4fYimb/Qmolsy3H5OHpV3igG45r8FCMVmyI6wqKgE2fugjvl05tI22nJrM05i
b+dZT/6YSaFpQ6FG97QaubMA+/E2y9rfjOY+CJ0/gdewt0umFz8uMiyyR99nNHX0
8qT1NXKsOd3Qf53gXTglWE/fvJH9Z3G9nYCdkmg8C4ArTK2joemKXN5mGeXdwmuo
wNt55aSGyiszUH4dAUhPa0x6kJGH+0ac28dRiSOdEa4+9Fite/w4edUvheDMbsEZ
Aub3vw32RTVmKrJpgfNTUVhTiaoM3Yyk5vNDMNri7A0+Dh/TLYtYzVD85XsXR0TQ
Aiybx18gwrebDOLPFcFcMnCFOBmLRMDBM+v/DkS4Qnro7BksrH9uJ8PmNnsUuMbD
aWTLW57vx/DIyrvW6sH+EwpQVaFEtFmgpCCGI6CeuVgEQ+na/JWvM5JY43/Yy6ZJ
TLQB2DgqRKuhBa3BR57qfPJyvIiaCSJ2p7Nlh2p77p8Zb8qhmBiQ6PtqKeGr/UQn
4VSqme9CsQ6WvB+aw7LMPCgXjp2YYfOGhcWjSTRGS2+k36PG6bPjQw9D4nR0PHMx
ft1KTJ+ElQnBocQKtZQey/nbNGn037VuXsnkbzpC6lMkiy2TD17IwIzRERrE4Ky3
tvYvhG6YslTmQXKTk40U4HcLfKAbcb+kBtoJwAfH0ZxeL8N4/dnQ1zSx1pqmwWwi
QCkNs9lY7RaM09uQmXuIzoXU88OnFoR/f1HT4hkbXN1YsMKUwDIp9TfWVjcp9CQh
fzquq0hlYukVmijWHHcjcM8JcFbiulUCONbxChr0G9vSoIJeAIq0kxPNYVaG+YgM
0Os0JERFbjmugli9o1fJ9APvh9LFv0i7+/exQ/QcXo6WkW6W5QdE1XkkpzImqBUk
xCai4gSwm0fDzjwDBehAVNKCmfaTzzxrNC48EG06jR7G3F8pbjIS6OcggwbQpVwx
BGpEaOnNEIcgZqJ+AexgjHvmh/OtBcFDrxXopZj7vBNsBrSfT8aX4XWzNXHvWpJy
Z4Jn17QdL00SVaaq+he+D0GDp1W/lypRbB6Cs4uBO1bWzn2fkSH0jefip04KaeVp
oKh0y3WkLtGYB0utO4aw8svA7ifgg6iJZShbWZDGkmbL71LWU046yV6xJdwtueSz
V2gzSFRuzutG6XgEq3eyEqaJ7lQrW7gpK7TTVQ4BR5vWJ3ewS9OGha1DdHu+Z1qq
sDhSZzAWx+ZqmQI43N1zaor32QCD9qo1xK5DK5sb3A5rBd/YxnoR6WDh2iIKZYVh
/FXEgdSBIZqYjorrLc3jg4yvXjXGBWdT6/YV/YjmIwq5u7WgHC7FbvkDKlTg2Cex
EIEz8wt7fFF3dKoSwxXOwhdHaGjTV2RtyKiPtbOnjLbXIHMoe6W/tzvTRQbxw8xq
L9AkqZpkr7WxGu9db8jLuuJJJrEU2biWeXOvVfjP0v8/9uEqG7buMpQlYcfQYDBh
9Ps4bRAIGU/7J+a/MVWybxca4s0nvWsybTwaj5nY1FfYeMvtEZx/fiO47UQQYdG5
oBtMT9SO3prhtfSF0Zj3daw0cPBU0/oVs2d/n1TlBhyd21zUpXkllhX+bpXh2RQy
H/kYmz4sVnf4OPtwugHda4Sc6rOeoNsVekN1x+WZkWqwQyBbOe8w0nuNZWVNytpX
TI1CVzlDshBVFFp9LtcfNTWl/UGpg4cPsy+JmmylUA08qaBU22AIEX4xsa0j8hy1
hoHk32a6I2wtfcxbJ5zYtNmjCrDmfc+RrXn1vkt/e3Yj54knU8g2gh44ekVI1m1Z
Itc6dxpQHvjeAH1ZjlOkVxYYg5M2cakmIaxg6QdEznxlw+1USC/BSL0vmkzHCEcL
YTB/h32vdmadXVKPFQlWxxL4ktUQQZkU/OfSAGcVqMp1mPbOxvWQR0KScepqpVGm
+OSltCrVEYGDMKsAOA+6x/45VD12NCiZ6MqB4+6TzBwqWBamRzkc9MT08/yJaJF4
9kosJ45tgbWrI7EyVHR0XxQ9/UMbHD1IQPLtxLEWbPQ3Z0UYPxPs+15HE0s/tSRK
csSz6Lph7HTWLzQwn2WMiTrLU8CCyMqzm9Nz8skbxQ8xITFHF/KNVZ5Pzwb3efN8
KEnSmZvbGC3PnRAICFm8EJifAeaLemra/J1zwI8zbD+bfmr0sncxEpowgDlliZ8z
gEATpRBgqLHutdfCy5Pcyy090HjNxhx3v57XBR2G/gEku05plj0cbXIn+hW9ddMl
FjEAz33U3yBRC6+jAp3dKdGQZucNwpJ0TLl3SmSSgUmMNwHeTaxdEQCA/yzOri8C
XHy8niHhFeMejErvYp8JY9er997KR4/VNXLwIT7aaZWgJENJhHA5AOCVTRe2l7Lx
bd96nlcg4ucWz55xNJVRMkdhsv/9c+4AG678HnAuKZ9ycH0sXpwnVF/rCtKt4eOS
/iLa4J8m5DVRcLrlNnZihTo4ckFMxkr5q/lArmfe2sBaDbbhkum6NV+2LdeHHGLG
FJLdj24BrgqoY+GUF4fbof3xcMxYM6OgXEvEJHhIACXLyvw3IpB4aYWHx94ddtbj
wLF7AkXPo1gKh6h0rBPBhjiB1RBH22fhZ96CplaKJwKq/939YJoR24cwPFfILTdP
ay9x7GYdb7FbVMW/44DxGChhChCJTvkeycwYTbO56gmQDVNtEtHbsp2rFVD3mIyZ
QeFGn0VHgGu2DSM7ECUOrZXjO7b5iL+PxOBUdVJaxq8vi2LGhksy2VQ3f3nfJv/N
cv9ErTEVgz9qk4sjxBhjwA09vd+UfzyMYRpX/OP5+Aj0YwEwiw3dzCdOwmyyQ7sS
XXTl3lmzS2S2upk8fUoSn09icljMW+S5XZSbL0dzA8nd60quWK9E1iDwH1KUcDgj
gCmfP1xeUu8R8vVbWi78jwnYD3IMzZyOT7AP/ZAzULPNindV9UAx5veCxAn4dWY8
1+x6+X66eap7yzYopL+OOlr2LflQeuWwUugYzkWyFUrroXXZtQkF0JPk1cTt1Bvk
WRDOjwR11kxv+ZimP72QyIq4AvJ33SMFZb3T1Vp62cjEA4REKgPtK3yufN/tSR6/
i2GV2EtjPtwGx+6ELcEM3X+uBLvA0JLa5zwNe5qxepiZkIZnbSFCmcULXCaEqyQH
Nmc9bPzqS+EZ+V6xCnXIvasgleJPAWtrIEny1luOiuV7DuJP77mRAOsns91PZIdU
+r0yqpB8kag76hW0AVKTsLpKbTqKD3Y1TPOZBNQdNTiflBbdlNcOrWnenmu9fY7C
2T9CUVbR3cJ6QThE4XyyCel5s+PMruyV44PS68QA/4T0j5igckCZ61I7JKLID0mD
8l2rB+d2SmkRE70lftZZcBKQAxarLqx6UHNh7ErAOW6RF4fEOjkd2Phx2FVE53xO
1GBcOZBP8qnueoORXNyHKEM3XH5I170vNzEYQqDlO8QffeZC0P5xzf7Lm93Y3vHA
tq4JMEJwAY/CaSbbEeuKB3yViELQkaghAq9xDRy+bms6nJPhlURtSjeJ7JqtUKAe
aKu86OjQb9ZvrZDnpMGw5+ioAMK3EHk/+CvaTsXcgSGb3aycHcgeh4uD1iQ8w3kn
TU8/L2RQQ4kFr1YjldjxchHI8DSZPq7K8WzzrCXqKAoaESZkK4NDf84cZ2TqUYoC
iqtqVAmZi4mrKJ7SnSE9CvV2QhhaKcD28iLe7+3kcH6ouRMf6+t6HODLpmECARKi
kAJbxt20dS1iWiWMgDmkmWvpReWwqQlwzhf8jwqz3xBfnz98figA65iuDjrzcS2+
3el0dJJGyDBIWwzxNE8JKa3RDzari9MYltLGb4PZYRwviw2VnQdVNO+eYNnQjOVu
YE9vwTi8z46E9SCcn4BO00vd9ioFW8OeNtjYsn2pEv3awP9B67kjlSLmwyv6QQo6
5bwUo0ufAoRnGRXMyiTSacGNWc+cWO9SYOZNs/wB7kV3excAAHuUS7Nr5f02nvLw
Kf2i3hCZ3rBiDqa5DqQy7Qxj+DfYHt94Trbg7XBT+FsxCvg6s2z/YzbXYsFFQi+w
c9UKGyT3gxs3dpU2KIoFKSJRpa1KBqlPtuJeowSukm8nf84Ei6fmENwOJcbVy6Vv
cIBLU9jWOtY8e9dOYJhhyoUAcwq7sLZQ/26/vYHd0leW+sZcy8nSa3i4tfXsme8v
7EDSqqcH0KwKUck1A5aon6kkQcfJV3DFdVSmpzJeD+XK9CqMWZiJ/2qjxTH/omH/
f8HJ8O6MKjn7AUYE3rcKsol95N5EvKLfaCSdTRWcsouLhg0aE7fZ+gQhY7SfStiw
XRIUQ/ipelFTyobjr2HM7LM3E5vJV/9N65X3qMejKu+cDfnah5+fCZEEwD+zEMPb
XEwOj96DuBYfSnsRdb302fdXCJyo098jks/34BHZcswasn2MfTnQ0Bc2JmbhlzJ+
+KZdElvEeuYzWk0NR4wPxokld8a5owospxWEA+YGrYJwB/Y3lASiltS4c5rHIiJ1
7gW2HTIQAj7A1oPVOCm4wJBJarrsH5ooajPv0AikbVzD6z0WgNHIK3Y5IftY8sqa
XDaqQolrh56np92yToYmEHnyJU7B9FpVlMRak/1bFX/S31s+ivrIV6ghAry8bjb1
2uFHFnDTC8p6+sJ5pPmRWigABGBF4Lr4mLuEr7IhXw6kwv1gKe+aVkDeVjmUcN4b
X9iD3HP9BR57MV48WnaLx12CLBV0rBDPpgi1qFsfluEjbtYW1kOc4kQz3DqJzyPy
jFgEBhszIBmqzK/7ixtzcH+tTYLAl6sZj2tc9Sb8U7Lo+OSD0yp9qr3aL7DIuOXn
B63tuTwdfwFybWVFQ9nGDMOGR6zba3KqnbyP3IlO8xbfeLlYW27eFqlKWBWY1R4V
VxnNbIeee9LiR/hb4KRy9zG988JbYjGmWv9SQojHlRJh/3COZolisKbSG9mFPPBt
iiv4lEXBXOqawg7riKSLOz7RfW+f3oJ0XW15xQahjlqvzD//ZzsXfV9Mq+n+6REy
KKERM92Y+HVvCB9Bu4B4ao28VXAcFdIIvqgzncHXvcWEvQujzj8zlAUillAs4hBd
T5pFIxnLck92ZAqQQaC/MjetyHiQD7QgHva+ERUgC7Q8utc/TV7qtKBFikmWMdv0
w3nOkzWmqnamZ8/JlfRC1WGPPtQ/8NOTo1Adgf+ODEThuMXws+x5sNlTG2aJb/mm
oublp+CFp/9wBIkbUjCNBI0GRegebwOgP2zypNlgVtJRzc9cY0gD7J1Faz86d6sZ
wVgaMeobVvurfgumZp5u4zg0ZYvS0E/Un18w/Da46xZK06nv3syQHF4Wp/+pV1qa
AhsRW3SCW0HlDzY/q/fj8i2gwcjJLYXFzY5DukaPFc6Re9dZh6Lkv/tJWebq+n/c
Cr1P0AetVQN7mpHlcRQAdPDHMEHsiWApg9qiBOWIYu2Kpiz+N9M3wSIp7HqeAYu9
bj85WNiducX6WmPt6waVgEhAUKxiHnqffVkAcGaT2cZdEytj8LVS3wPh819jtPZ3
PyIjF2oJ64f1QEt2Nuwhg2CeTp3sd23wnMsQLj6aXiUkiRQ1KDVKa7B2ZDLD/XAP
Ul4Mzu75OJQ1J5MP9Z84VcxCdS6oQQ1E95UwX/EPSz9NVun4KMQ1ximzCcMGIfaA
zuqC1XvX2yoQpbNBn3smuzMki+fXcU8XW9Z66BpgciiN+yigmVZeknxTAB7H1lpc
Pu9R1sXRQ8Qog4lYBXW/MXkLKKWsE9QOsjPlwlwTqFK7v0k4gb20T0L63MepFV2t
Z8V3N0krMsENrK16rQ9Bb6/XXZzKlK/Sfut7Cxnht5g8CmXD2M+eIe+kgtZ5xrU7
+4txdemXhJn6fNyLkfEsBfum6abwSS3SgRxFvosF1s2Cd5zTKHS3636kwfi3ohHG
TzO7x074jjz5NcW0IfOs4IlWjzKzb37WuNY9PuDf/EkMRSZImVpkX2YPrWrOBoO0
/LVapBgyfY5GypzGSNU8/kf+DZ6Sa8Ht3phkbhl76WPaOYMwrVa7Euaq5kHOCrzl
KAipvTBYZqi2qKjspjO6eX0UmnfAkzy0kYk8oE9TYRiWm8B7MN1mdJRRVnB5cpZ+
2qmDrsaCHesDYdODPSR2jIYVyjrCkqaqjyCwSuMQXEmD/vyHXYJ3WfdBw6qOmgHc
LM5wFx9w43B857G13qMmUjNgM61NI5xSvC30dNkiPhD9kTBD19GHvRO3TeHEUStv
brfw4KBBVfDeY4ymGoY1Z+ZWSOFX+DWMmy//Ce62pNg/a8aRZWhU10vrAzOZ4swx
Z4idIogH1AelLsi4lF75vmJ5XID39od/BkQs1zy1EpXLlBtsVfcK1lhKfNdnVbJC
j3j7uRVhXbzJHtDS0BwJuWtGzq9KnwUNHAMWUg0hu44/D5tSgkkwpIbTQBNZppOX
AASpmZCC5GULCwpRaWYYDHlWPW0IBCjEVykkTbGD2u1xOW/MhB3Ou6ZxNh96fLlj
tFVDGyY+r0oR+zRtXDRMoXj+2ehYPnm14+Ov885RbkdmKLnpeasC1twiNpMLr5c5
IBjOununQBaqLTAfVVOdZkNAsDsgx3uBvxnltV1BR/+FYJDwp7R3yrHmruI9krRV
y3Soh2/7jYkOGBl0OaozMBpIaO0/u8vlHOCaE5AGfRTOF9w4rq7YsDqFpav9NXZs
BSSjBpe4xZWd/KrBRL8NqNiAZIktmwKSdW4exdRATjRS8FW+whVHS3tevG1ATYuu
v/ov76OHjAAl18dXS0AN6irOWjJCyAoGHb9fsEo40NSyNZVIDbdK06kUSp2bfWh8
RAw/fhMhn75PaubHwAVO6XvWTwqJ19X6u4Dmpii6b2VexLne4rb9iiirR6Npiy6F
PXipqEGXOC+VLrVVz3bhKsHUf4NDIg3dlvYYq+f2pkwfPB7I27Tu+0LPtaL1NTpE
T5B/+qnKfH7seYG5YXL39Tq1nB4JDxZ2m6elhxUjtR9L/LY1V5OLuDXVcgNVT6AZ
Ipv8cDgVUtqgZavGRww0kTfUGYOz+PQH/VlYg7ehkqHE+lNDQ3IoEWZmLiizSBDQ
OYA077OGsjA6kIzYw8/R6vmc3yJV5QxbTa++3VU9p/c7C+EY522zVIrRipJg+zEs
KrfREuh8Kzl/+hiwDWYKcjmonb6UWAaEGzsJbG3T8L0zj9U54VaIPgjsln4YBiPB
HEvty6LSm+QXU82sQbhvrFYfcZUZU3w76nvSNhtb9WbVBx3xa/o0f6SgebCYMg3W
3vlPD1uHrCK+IWDpMsnxy7vhvL5LA82++m3oW4lIXQW15EN52cQuS4F6kUwFXiU+
ePAiujAkykElNNQI+T2y64CLTsdPDPq4E5DAJy1qyZEnE42nCrvepzPOoWUaL7zb
nQcOhrukc46sS/xQmzbWfOms7pFnrweGZmaoDmu8Mg0cLZYOm0YdEMbQiVC5mYow
RBZJ2e23BX4VYYfV18OrDEek8A/byYzuXAb1Sm5s4fhFkSeJA5lK/gQ4OidrD6PB
iVpHVO1HLwCNk50zUiz/heyISqXAn3LWkUG08AiH9cuqqN1kOnOiHEdZDSmKU2d7
eARjWP9R2Vg0nRK39UN9XG2kLoIiaF9hPnb3EoSQ4JwX/TP7fsfd9O8NZj2Fzwki
kW4JjK5dRTigLqwn7kcXSohW9tUbJ0s9DVGnrAlUPo1GhoczkbMWwi4h5UsGJLx+
Y23ZpxAYut8E1+YlJhmraj8U/gZHyuFNaVC6PgLgnpChhxEuylzrrkXDjPqFRQW4
xCMIU1T6VUQWC1VF4bnMXZRqbkn3zUxYgAB3RLNCMjdvDznzaRlgRjIAxIfqdEru
Bs/kUKgI5OwgWcIOcjW+Oh30Uf3WOPY8s8trYjaGUUf/vTIu3zxWlBaRQZKs0Zso
dFO9+nOYLv/uFbue4tQTEJQwhoJKFkiZ11sug77mP1JLp15zYJaA+kdOStv3iWzh
syj3I6A+DqYa62ZG/WfUXWgiptQROAw7yw9L2iedbXuOKMa4814Jhl13x4eVahRq
fN/VBBMbEMQjYd6T4onX5eGZxPZsjAECcQzADVzWCQY/JEbB4Qct9F8/kxT1PGJA
akf88OzFwwsCTepl/4NsLW6OLE0BNHdQsuP/jRXs/oK+STGRQYSjyM3juidGv7mP
JzCvXdRDPV6z6gIhZ7EuRSrpTiFm7mEqpJ7b/3aeuCypc1O2AFmXU1sCKNOrz4DL
3EYUBLv20VdiAR3r9kc6BM+cwxo8MtexGTp6fD/Gu+i1IbhgZe/1MaeaZAFMGY7b
4Q2380S7s5QOu35YpQgGFrfvd3b4by6bY5aG7Wsq9nHS6s2GArgtx/uTKfcKyRby
fFPVnbDlkuA15qkZASNjlNxyEcc2Pu6OU11lhKOCB9tYCaTSVYxGH7rCn3lrCNKa
C8scwnUnJudpzzeN29YHODAvzuGfFo5lyr8OCgG2UY0ry+r1Njp6HDWfBwaJe4z6
PjyLVc9hpELbrqbdxit7YI4Hz9zwnP+3mMZ7uHWG+FmZoigLzrIlyt2ekYzJuQRE
9afvQYFrQso3xiYiM996NlG7umXIFgug7qppaYrKi7dVhuHCv2DIbKTLH8On8bR9
hjR6npQX4PtkY3hNMY6xsLALpku3SVRISEGKarBgLXwDq7aYfAAYcvw3wL8+zvFA
OdX0MOWxg0uJfrYZICnD0Jc58rlB681cAfHPW71ckV4Pd84AgmT/CqhpgoNhK45W
fpJtku2XiczesS8suJQMtZeLJlYpG5ZFrhorWYnr5zd4H0oLbXVYTS282AqYe+u9
36r+zvsz7SM1nP+NdrrzLwDDqV+wactgSx+TNRt2N69X0PjMm3Y+PevSjFVQkrCI
chma0XjuFnD5ueIOxt6u6zhk6ZptZxJ1ugpJuKUZFkWtcK7tJumxIe/Erk91Sqbv
2p8Cs6CHjml785csOltjkf9k1gmoSk/VUNyVP0LV6GxfZloccJj+d7ncexwToU5r
xneP1+my7oMT5WcSty3F13Dd67E8TNM9zZpnLXfvc6HuULNsxYlDgIrEcVlLFigT
HjCWbxVHsdiMntSRtAm2wW/P2UIeP2NH0jruiZduYgmiZTP24lZ46HTXT2DTneCa
DyrZpCVjzl5RTQ3r8F37WwCWfldAow42QrTS2jhJiF8BfGTYaT3q8f8yUK+0TRsj
YwpLZYp5tAf3ZoBiaMlOcgKawZFgoBn2qLK4fkI5hWfI3wQYN869ecvANdAB/q9s
XUjMX0jYEN2kyyTwYqQwEYZtoOWkUQQZ6oAeN/WlKVOu1NvFdZWRySerdPmoYV0D
TRk4jVzaPrmEKzazfnPhmHnCUVy2s95cDfYRU9O6EICZV1LwluJNm9Kgw+pLazK2
gqQS/UQi9o0ZLloymU4TH982Dr50poGfZrV5SjrhVJrzBUfSJ3HAM6/M3079d0au
XT45VkQhbw46dzTmOT7Oyh+/LiX8aSXyKIUBf3FNyuMRFWvNLRNbZMx4wp3ufThm
F66kpHYXEZPT3hBinCYxBWFAw5cCaV3chNHor9qOnSimAcHueU7Z1Hdxpaj5dPrq
RW45Cs331wTaZV+g3VljR1imibqrAdhJi9702fNIJPYT2IUcwflCp3TD6HtwT/jQ
Y0yurFduIN6/ok9TjlgB7FRdS3lZavph6TkNlX/TIRdubU53qmIhAxRoPc9hDlJR
u5XfWzAAkfEJJZ+rHhlyAhSBw+gfVRFoIUaMDwkkxUkFMPZcHoDMQRpn5fxBlabk
fwWS2wx+cN0G+za3TMxBzbaqgie0sIXEvyy4kuNkPXq1M+o3PKp4F7cB+TEi/HN6
NwzNoddKRLxLY44ccvEZkg4cNrkYpwqRvkOYWGU9OkOQvp0a2tA76rMdAZh+vVcc
PBVhUsKcPGCJP7QEYvNu+3AJhhOjf4M4JUPS/uxRKT6pkWgMf9GFaBTTIvDxU6lz
lTW68FMfxyDdkiofjVdWey/tQYcFFk3+CCyWeTkIeO3P8Pi/oaqRMZrdUNzlcJRu
tpaI7Oe+enTqK6/VGeKdXuZzYhtav999RejvPOAMFvgpjLWUGsU9U2KxWhm8Dc6e
YhuZCTuW+FWV2bcWwCuU27/IeknOPhvN/ZtLb+hcRR89jQo6HRtcRrKiBFPTRPbR
9R68bUU/vgm7sJI1k6JbS/NGmWVZpx20jNDXSX8EsGuN6vRjcqQOW9CijtaPzlRQ
g5bz7KHC5bLaUXuEo2YJBM0XOjt4Z1lWWokr4vHu41SCa82uSnmxK5/7wHFNsHz9
w9W2ULAiRlMFgYyZb2M284wgL84GqFeWlBljCaRoxfPct2mHmzygmw9DR/ak6iec
n9La0XJ2Dm9gVmNjhgqyO6G1xYqnjaj/A1xaFTljBDGzZ9FWxi9hdFA7RoW1U/e8
C04JBilKzLswheFQfYHFLWDrXOj/spKMn2hBsV5cZKNBlSqNkYAn4/DAh/2gVRpM
vtgeHlEqAnqelt/2TPgvjFcUbuZXTOMfi+J0elunIEuX0KS8uOo1xAhSCVs3zq7O
+P76VeI/couuozS/vwL511iq6lipMlZMmvCaiZRG9FxyEfG9KWOQHsJOPcA7bc7p
/S2NehoBM+hoVxOs83/x8pMM2VDCt5wFDLN2RLo7PAACRmZ8CoEfpvmJZRGnjBMZ
MJOC0VmXEuEBdow3kvl0so1Iw7nwmeLh2D+8lL4uLxEdt5btMqb3uHKG+cpZ9W5J
y1+c3Cyj59E0Mmnn0ag464lcfpr+WhpXJgaM/U5AZFil32uu0y/HZuyz3py0y2k+
hlQgtFazDKp9UGUDGWfnUq7y/Iznyo72LAeuNLI32C9eC0Zxbffo0TS71rYFmb/9
fKHpoJR/X27rqfOxPwKB1QzCTdNx4g4ArtKGgtvGroWFrUNxEV1PPvymr3SotswG
cintJ2LvOdbwe30VvBfj/0XUbm+h2Ya++Aqs36W8BUqCBj0/2R/MSMzTXXG8qZSN
Z+GwY0EpANoGCTZdl/4gxAbIwf0/1j3b/MDfNn0/lIB5NOc1k3kjdph/jYb/FM5w
pYQrrEGCq7bFKI6Qxcdv1DaZG2h1nOHDPULLfKrnruTFQFqOJDR0FdFXM1VlEhEF
V0Zo8FCiVFsvDU82osrg58HPFR5OU1F6nnpWLno2kORVzmGvH55iVs9+G3suw7W6
n2JZO393QhY411lsKECRHgK72omwOhxIcKYcPkKg1VI8b7OzFrP8ICKknrk9DaiQ
KGrj4QiNx/UvhwTz5H0niQSjKN2ev4kT0Nc9tAQNkz0EqEJWMYiRSgLtI6Wl0C1e
DFQvmKJ/VdLh3t4AfyaGyObiMUDtT4ba/kIvJGHGMGEn+TqN+RxuwOnwAcShXcAX
IHB9qInx4OVEUriyTBemVNZz8k8kuOwHT+n9/mws3MHXd8uqHP1Ov8GTKjmyxdbT
eeYn96XzeNQsRW0wm/UHfCvgFvD98a1jRQyPt7CSYdGGbj2g4BxZ5lq7YnN0z26t
pNuICQzQ/0Dwh+SK9M9U1+nT/NXYbKe8sd4NRF+UX5Took1rrLG3MCM02a2NVapF
Cva8BebTwHmDz4R1CAy1erfvCov8oSBty8A66evsiqBOGdsFuWGcviFufis/pMtU
pLHeghsTaM1kBbFOAyQBXmZIrNcgg3dpZB4i2dfxvEKWgU/sqw412Mqrwy2+4aQf
4s1Zs2icVmx3QjTWfJNvKzyOsPv6o1V6r4D8ArVX60McHp5sWKmQ4i37Ij6qT3/s
3EFj1GJuaRqpdrgRc/F0QbdPlede3ZSijYW68IWD4fmEvwbeJiO8GFFTS7rN9P+P
y1/p2T1LN4/r57yC3V7lx0UQz+gHgy6hzkgaKD6zfodoCu8VA0RDqXHr3YgWnwC1
Tg05LUZH96cx3bLar3fnrbWZ92kfhS4jtzP2wE4TTVD6tVQDKu7x91uamNBzcTEA
XAAYCZtpCXDN3Xx1Wi2pHrmjsBB77NmiiAWX3+iM5CkGVAvzPlhHt8rcZu8QQBOY
VxDfpSJbo9jTDboa8c1IPKLn+1OvI3YX6lNFyZaLiS0tdBjtrK4XDLga79/yP3I6
E2ARu7Xa/mwFNV7bXVihLNmPozDHVdh+lESDKzTXTGvqbYjXgnJTnPWRBZ0x4pmy
U+OntHEcf6tXFbHX56UEvNE6hUQjnSdj85c7R27MtpXcWBB0HIIpmbx3aoI3lpeF
vzivdzyyLL2T5cPfuhiLjiT5tQpHe/hEq8NdeOjFjeyDyxSFZlQoSQQSoHuOklU6
BKKdaRaLhr04uEin3Rc0672atDbyfYxmAYIMDBYH66fiuLKsH0b1mwyd9cT+vy6X
6y7Wvsk4KONpVluutdoV/RFQN0Wca16nHTwQWVKwZ6NDWO5ZVraf9RYILR7TQimd
/cL3FWEEe3gjl1Rr/rxvj1LvSi5DiLai9eZWNgWV2S9YJf0VR/E3FaUZ3HQjhXOH
yJHpDJGWXPGzPP2IvSNCx3sx7HGMYPzdazg5OWv6lFL7Fn/GZVRRU2PRULoh2y5e
LFCBga1otR/1I/gUe7Rq/Vb5Y1Z7irX4m+J+0Y4XIILfOVfB+mTtS5G6wQd1WAw4
mVBcrU+LAbhWFJjV89mDryb+O811lo9sEQ6XZkSSZDJG5lmXoOpVef7zM02Nw+TZ
CvGUo+gTDC/1hatu3D4M0Kzrn7bG/ObQVxQG+hCBznhSd9I1ileO6PoxVuVzRhOS
lUKIRO/zLmiJ/OiJyAAwQ75JmOxF07Fr7uQ2hPYBoteFuDX8yrLpmOX9SOO5sdJY
kIREsBykpBbEWouFnYh9QW+8S+ldLXiWOtBXfZsfC8wzQkp5STXQjJhBbJomy77j
JR7kchJLdlpMOKno33/4l8nBjK7ll6t6HlT0Oc3rtkrKJRRBeRImBNYnQX7nBi3h
dTuiHdYGrZ3l+EhEjoD2Drt3ekdf6rG9IOEiqpW6ykpWEPM9VPs44U9PUQb1jgjD
4th8JyoNGzPxjoVQmlkCFT8/SDTM85sDEvbpEik0qIM8/CHAdHQzYu+YNUpU5B75
LdpTrTWm6DxrOF0gQqLGeF5hPdRrQBsdlFaLphaNZ6urUstOr1RFm/SqormIKt+F
Pm4hWjitu+cWl/7RcJEhP3uGRIUe2vMD0NuGhsGsIQpnXg7fzsjOfQC0omaKWNmC
6NBAnY/lT7lqLKnKxGhvjXX35IM7PIy+Ew4hqlmKDUmYcf/dJIA/cdW1EL4Uvvvm
99X8GcByvJgQXMzUh2AfbLnISEj4syiBw9uAMyhtX9FQQYwmTIebk/uPplGDpjd2
SXQQMVNa+lOxQviN89HJ2PCqDHKbD6Wge5cvNXitmlQsZPSzZCyyMOnuY75gGxgA
GotJfgIu0a4yZfRUr97ftjLNOFYcFTfl1Lzj3psMLwql6bro1FYFIwJf7ANtrf5b
sVG3movOVIF0Xid9z0OidlFbP30TXkBKeUPf7zmuUlJAtZC9Fn5WNic+5lLOLfxJ
Qa3KBnYJTKnWVNwQYZF+vvdE+qNNRrEB2xywal7cd6C9EUqgzGKKdiza0bjNV9Ph
F1i95oVtTsA33OANTlQCVF/3St7KtBYIQf3RfwU3nZNHD75qRCOhqkuN5W36zLe+
qIK+dt2aqh+MsrwHZrxNB68up//CsmEicUDdZMGV8e8sF7LCMOLloKvo/VB3il4h
2dqfJG+WYYmHnKoyKZasY35oBdzk4iE/1ro0QyvvpPyT7ZrQgxFGcqqt4Qaq0/Bq
DxzvWdhCQegaU5KUgb1bJSrXxfnceH1RF108sLWOKv8lBLIEai4i4KjM9jKZ8Zou
372CZa6Z1Eg4BEmHhnlo7eijnM/ebe141J6W4FnhKo9jWdbB8x8iZb/bGlcqwMP6
6HcG5ddtllxRrq5wgzLC9d4CE29uUCRjMhpS64iVuhvQs+nUHZdBCBI/YDiaClI7
TFLXBo4BGXeWYqSS89H0QV4K3rjPLBkHWaD7Pt3PYxNjpUtdRrKbkNysXCsEKAI8
hjZZl2NZRTELVdxCMqqSNxAxt3icNflqdL1I5CDtLpCi46oL8zaLVjl7s2Jc3h7b
RL1q2s+Z7+DilV6OzUo8pd3PmDENIupp3sT2yhjYHG6yMN/hCi1v8RyR8Iv9yRqE
OS8cEEIkOnbfQfLlaL8JDEA3kcNvPdoXHmp3cyBmfoTRItLG2bd5iA4x8Vph0sPv
bRRiRc+4B2OVLvJQN9khbs/OJtw+4+vosDCXR/6cNYi6Gro4ZxCZzK+XOUU+7K6S
wlUXVLyKYDV1qr5KsS9lV22lC+DchffXMQr75xk2G3nI9hOJ/Wtvd1NQmHlPpBum
t7WIA4EHlnlraGewJtfSd/yrmGM4aM2zphtcBen9f/WRNavu1JjXwm+qa28/U1/l
YjXjxFFEW1HzmteBtZF0bqzoipygHbXA9wmM0WGjviD11SnaXJA/bmUPHhiDMtRG
aMBOlmR28kerBBTQWCUMQDP/QQLQ6DMpHjobQzqroEX3bHD4SSEfoXQ7SvhBMkgL
kY/ZLzWoVjrft2l/3lD2mXiBif2wcLzl9duXP6wnfnp0M5ml+VdKloO0mcKgX4/E
sDULt4O6NWKCBUavcDVnzja359Jnx3G5HRGzxp3Yif1ib9TvsFd0tWyeNRSHU52Q
KWZ/tL6WQBT7A2324mr0ClicaGkcqUQljyH8Txe4pzQxPHs756xYA7veiF8C2hIc
dGhOXcVyKBoJ0GXFJQVKhRW+VE//3hVTzTpr+GEGEXLsRYEDnbDNKBe74/s1L18h
q8mE/WOolKcFlXplg+hnmCfMiuTSL8XF1AIkNFgj3YRd0dWkdkHro2iJP2lTTESk
bCnPc7W1XzP/bpuSoZ/P0kSY3pWJJl6xH8bVfnsrkwAkpV7Nw3mcfcYV6r+/3jVu
0R/Gt173TY2WLZlDQ/cuHe5kD0/d3xP16Tz4zSGoH/7ynxXJZBqIeeZu5BVxi2Sj
R4DCXstT/478iUoPyv7V7mKQIvCzS2aHn8C0dWk/emuv+9e4Wv29dPTkvHZCDqET
BPkTcG5Gv5oWiHjIY/ReZ/SQGCnwikUhs/0bK86LrOM0baIgUARxijJnfCrNFdf3
ad19CxwIsOlPD42IKP6tJcb/v/vDaDKmff0P5hqgnPu+ei3q++WnF5KekLTtAk2U
YSoF6Ls1F5+ZMzGAn5593mI1JntKlF5JIHN4eQvJfarQ5gm6TYQFVbw64BwUfKNU
7yx0eReDUkYyYF/CiK45LNMmuvAtPqFLknzA2+PR+Fvf661tk8GKs/PW1Ffr0DvW
BjTnNth9sZWjhL+ZsFzEAvAwmYqzErahNGq2y9ItfEG4vfUFknLUEZ6whwKbgZUv
lEmjlHHm67PKWZ1XrFnOIjttstBN/bJ0z6ytU+/fltJcgqt3BQJ/PTiI2ltRXqn9
u885aYRjHICLbR/QNUBGkKRgN5Mbf6uHzyaWrY2V0zALiqrXFSN94Xz8u8suppB3
mgQzeM4a83JXO93whvLswn3MnCzDMJvpNoelMzYLUIqCscA72tuFH+70Bsp7/ibw
y33EkwfRObSKLvD/5bnRYy7oaJOpxPDE9P0zjpnl4lMlPeO4szBy+nFWJgIgYji1
eGAwg/2V3uFbfIgtn8ZeZ75DAPn8rdVOtU6DNVZfb84PC27sOeu3SuE8TTF8bl7B
W1+XmuUXpUALdS61hrmmbVnb/cBgWSDkT1BiPhVvYnAkLOIwcwTabU4N8BpSPhKk
AVHGGgotK9ny8Md7UJhPHQWdhwi/Tz6Jgfx8T8xsnj4d0/8lwJHNjE889U6ByOFy
Jus2sOhQVyCsyXRow/N3bChN14c9x2ReHILp9mAQofURNAs+QVtsgoHY66xRS673
syNjI53uf468NALrufa0AvKJjEBmQumInGlaqn6DLYIG+jDknX9gFIk+5ictauRw
sEMO0A8mInqvphdeb1c/TkN3j5tKc3mpVqm74IvOxeI6/uVw5QTQAUGfNgysk0la
zuRPqcSsIF2GlNz0/z5HoN415k5X4eKlv/l6veQErFWD2xuLe1r/JXejXJznP11h
mmkDKcB+joD97mPw1hx3MIO9YZe1E0BG293Ly1YmTw8a2J5802yoK+jM6b/zM034
ZS9Jt8pGx6o83uiq2Ybu6jLmCjujYp6RnNxh13Yi3rmR5RQHUQLeM5m+LUgdh0e2
N2qiUzdLzgHG2S/q3FObCJiesYAiWA8gFW9lOqk0f34ahEeosFCAwc0WTxBysh+a
0Z7pxYsB0SATVHcblD0jXnYAKHyuK0cdmXFFvTWnyz2z8bRKDGoqjHn3SxKmddfo
cXx/evnAntqJLxaAptqVdV/KLvFquIAYbhvPtuW1vLnJZzoX9DNnCUfpP7Pcfwud
vZVpa6ktL+Sfw1uSlMRPcasIQzBmjuKhcZavBDcy4X7D1BnHJZl+q2kLz+Tp78hA
WIfmTEwPH+WXtBDreM+lxxgdt8bRMwYwRYsDOWIDyxIALJRUe/cAitlYTpnQgQzd
srFf3FaUDkPxW2s3nyGVtvd5wMhTYaYko7OYiV6eXWAu8eIvXCbaRl21qb7Js6zF
VTf7Ywga4u0iJqt6V8dQO2P70R46mLzIvEC4racn3FnQUFwDOgbkkxrGhzkiyqko
4K8dPmZN9q1CU/tr2YZ5Unb8qObxXIRtdcQKn+BAErctIHMx5eRWVH0kr4aLxtSz
F4DckUify1NI8d35C+71wqIZ+r6cgtt6LjL+iEvFTepPpX1K4eDU17KRIAOw+P4c
zTkoEfKWFi+WDqxwjksIfmbozwPOPaSTOVG+wuTYz4nvJKS8UKPuF934pveep5vL
z7UX2HTiz+jNkPc/molfwJl2W1ndCF9kH5VK68pP2oUMKLBCUOVhwn84GqIPe6IJ
1Kr3cTbefUuNgyxhvhkksCfK0XQMFBJT/UALw3mOyE+6NRNW9mt/86wSTPzKI5yi
I5S7Wkd/yd5oG4LgA+jKjmILlXHl34LlGi+97CW8aL1iKCUkhtv4/7p7VhI9QGJJ
KzuUOzCk3ESbqG4nNpeAz9/20HEuY2tq992H3gvzDayC/5bLi8kzge78YfCX+HUV
nob/0Yieal5o4JXbFbFRm1l3yvns0amsWJUgALHFYUOVWnjAAOHI2uGvo0E8QmlW
F337sIIEyTD+X3kmfE04gzy1jQDsOrtujkM5KGL7HxUphNUmq9+Tq6+veVmA4Aay
BTvgM1avPqcnIceHMofm1JRnHPVPxY3EX1VfEiU3ugkRHH0xrxNsWdxS9gbWkCpJ
o22uhqlPRd8iOxvn3YY5UK7Ar/rXxBrAqUID7wbsTHS1QKloHEtzJErDgchg9BJ9
QZPZlV2oqJ0lAICL+e3VZCkUY/EjxbX1P1GbbfACl0tUUBUXJwbwjvJradjDMqp2
OGTK5R6i//f1QBIuArWVh+g6uFdMl8KZGGXAHNLVDmR5CSOm3TjG5FvuQX6rPxdL
pr2deL9LYdLn4Htf2ASm7P8qmnGjcH+JWgxDCx6Gs11RbI5XlA4FmbVDfAQhZA4Y
Ep0cpQqEcz6x8wUok/m29TusR3cJMjbPi4zOsaNpppvKxqlR5Klb9FD7rYJ5CiTH
tcwLlWP6aCXaAWx9aSrmKs7N4a5+uhXEu1WeyTbf7WJ5XDYOXS7k9ZTjMgy3Njxu
kf4GvnXTcIP4T3kH68St/ClgTHjo62ouLbQWErg964Z0aPuURyYGMV1YzZ+qktyV
+KLqxCg4GHQz0KAjyiiQl4hPv1iac0I5v/FcOuV0YM12e71cSRpFsRmjPp3WkBBZ
Ukmu5GjMyvMOidDFN9WIB1z6x7qPtnd6ilVthBmYDPsRAhzijnwvwjzhhsc/zMfc
2K9kNa/U+TYY5WvcCKUAmDqvjjwmK1BbM2TnlmQ2J1+V11pysr2lObeinmPvAzF1
3/4BjcjeXym7nli7tMH9aV8Vx6wfmPZffrHZ7i3at1Gi3uDHIjjjh16EJzfM7eVQ
SrVxpaWTFwZRIKA1tICKIWsmiX5ovVGTiwtzlTOxkHGFSdJCYEied8B0GTvNPqM5
2wyivi2QXR/uYKUOXP/vZFZo+7YD4vSnqgVV3526n4vvJn4cZuAbwhsFupfYaF10
jcR2mVi8GJZGhisfllr8ZrqP/kIH5qbHpiPYQcgXdaRR51LvJ71VJ0LZTl5Px+Ug
Sh0zu1qClYFUZcLDKMKYXX/bJjCRkRyxUwIP1GOa9pKrq6Ln52TWtmHGJvihykQJ
UpXYKr76JM5WWygt4T2BbVTbYeYb0lckbK1EdwiR50hhTLydAB9/kQtMb1EVhz5S
pF7YymHwRW49x73i8F1e6tl6LivJl30cMzxv1LEE54aKipUOucZZ0ex+a0FkbH4Y
GYpVsdQY3xqeNNOpB1bmoAh8lqYfw/7ClIwIcmVnN2c6uBVMia91VT7/7xMh6ykr
qAKhqZqe1XLSN+LzYgsiG4hm+BTFsXt3lFat4RasR7qMRqPXImK9g0UhcqrECbsi
cBvj7THEF78KzAy1236Kf1bHaSuBtjJXIu1HrC2UvmvGIwc+Hp6KURrOq6Avb5x0
crvDXdrlv6p01gPvM5sxarb7aHdBzkhKgkYfO4m59z8xbWwzKkVHdq8/eypnC+Xb
Gn8iyfSdcRzcPZXRZiw7Ng77fmJHGC/vIzACkj4zBNUlK2gWxS1rTrcsW1OJd6jQ
cIDrrOivnEmsbb5k6+BeuuVcq+9LxV2hgAdKqVEIKmg6p+zLuZuujPHSXp18/IuB
FlFa0urLd0A2gfAscM3VebyUh9KHmzqmv3idryMMW8YcPuTO2l3CTPqh0Lw8Jqg7
+zVX0bBqsGbeYUa5wvRTSQYKcGooQ8fkqbwhlJc2WAq02t8BhgC3Rq4H+cpMmVO6
+i1om7x1xXDxE3F44sqw8BraWN/6ECGsYqTxvV1Fltxrnwbo9eLany+UMq3uqp0q
ctZPlB4il7jHq7YUjyooCV8haziuVVNRaNLtD+pc4minkxJdLsRRNi4hUvOh1yiD
MhUv13NR7qD9Qed7obRNsgnRlFUOEWYssXM3V4KDvoh2zqOsACeYzrjKdldDiTo8
Lr3mQi+rSvouLMbQyD8spojWKGP3cf0/b58m8m0YjayTfaBpeFNbfleW0bkrR5Nh
3pgDrKv1tcLamoesyHfNSW3RIbLqUppzntaMjAzRSluZ2aOt1Br0dUd2CEouyZCf
OgGrDRdF17+58WrpelXQF+DxYxQp4D0BtKOCddyEtQaeZ9YO2wqk569HZLcV9Bes
hUUvREHbHcFfUJ7gDpOkuSKvKD3wGBRMebgRQxAESmCs3YBqSAXx/2qJ2VHr9OzU
FxTSkXkPF+H1+7eMlkfemNzcBQaftLfLNRGy7/YJoPnKzvL1WDZbBG3mhXNXh9al
vsyfPdAPxVyCWwc1IsgoyTzs/PLA1pyFOMr8yphctSAW97ErUFMIVgUqIynOe4j2
cfq0HdrtminCaDqUWRF4rRUVirI0R9ytNwAejMOjG3kCfFrA7BMvbid47K0L43L0
dBRfOdy33p+ZBWv6JM2+m/jWBvKicWfMVCWBt4MCHpc9eLdM9tVpa73CxlPWXXC/
5x4MCUlQOL4gVQ+t1BSq3Zv2e64cWja8vx5Xox/nf9CVX+7t+bMr5V9kT4RelFG/
gWXtb2aZ/ZBWKWCQjnCRN3TteS8u9lYr+P4EkIENFtM3FJqCtVWgvo2nwo+LP5RL
QdIEhgU1loCi4dRjpbT7IT0jfx1WPmUOd77fAGNQAlsv2G+gzHUrMs8Z2UQqucaJ
vcrujGLyDLsX4rrwGy2o0FT0BMCtn6/uxruCSPPJvwgYsnL8LbH+hYh5f97bx1IR
1PCIMlG/DwaW0rOrSLhPrCQpogp5bemskqcghKiJGVB6/nBgGjCmLQFTVPfOsV+w
7Sex73j7oNIJ6HXfw3MzU38VGii3Ktd6lEDeFobzcfh+sdJLRw1Vrs1spEgu5HVR
25IfOIpjufXoK70rRm5a0Ui3e7bYQvpHTW4P0b4HRjwBvrJs15+G+svQlDVBLto1
YN/96E4u3f+h2oqZOwXp5IjxteS+99niFBAPeaF6nYPB0grWS2FphW4CxLcqTi8o
gGsDVOyUHuRIdQvIPGztcyiZ6w9bk+rd6P4wH0q7926XdOFPJ6LxxR+nDCWYQZMC
dnED3pSkmuKFp6xWefG1d4D17fYLUeV6lxL+VUcvjH/bilDNBAsq6uoILoi5qB5Y
+74Z5oKnRZdk45blz5WFVr9lUksgZMaG5RkVhEhK3wjJV08+6IJT6UBwR6l6yhKL
cU3Hkg+mwH8Wv+Zj/JfashLn8S0JAZf7L6pIEJl6SOER58/1w5ex1rhnoS45ZWhk
+x+T+PQloIeAjQz5mAwZUgERrQkAeFTcsyxKkXk704+yOX2NjQ4ziL8khiAkgsdc
mlndIM/tjsa2q4afEg59xfOLB/yfPjA3tg3VlzaVHSbALJYVWNwcwk/kh3dMeuSE
a5lGHcmHOfikqO+v6+I25CxBnbpDYBZt6I6eWgXPnT7Y1H28Rmm+mklUyjGIn2Mx
M1GlJ8a8cGIo00GGpEkEXmjkSON0M7XXbk+/O90ZFIBwKwaGCiWvXkAuGbQt3RK0
1MWYpJljLmeBoF0uzbuxJBIz3600sfA/uFMj/x07WRK6LDw/BYlXzfkgrzBmfkUC
dacdeJNusEjg9lg0DmwJ4mnMSzhrjIu12XUQkL6Nyj2bMXMRRqHFO66tA1qpJsku
8IgFfViVu6WrHKY4d8uqyIZu+F+ibZVB2LlsobU1Vra7OWkAErUADweqrBmAhNQJ
3j+oeEWOCTZ7/eszH8MLJJQbfk/J0YzyzaEHdtRY7TQ1QTzaRpR5lm6ZpGZXV424
LT2BJ+qQvTNEEQvnBlYeq9xud8F8KWe7obshLAMpHBsJHNaSJRSmMWqyL+kYdi4p
HIE1X3kBl/OVRiTfCdMJ89xWgGbkWcZ7bB4IxdDibNtgcvjw3CLhgQjyFPMJfkxJ
lQKhUDLmfIqjNTSezhfvtyk5flpIucjjxfzdEeDMp/MAQ9YfS089ji89EVP9aUjG
b2zaoF1iMpah3LIJLudCTwh8ONCUXpuk5DSZ8jqxEp3fbIhfuboYJrDNuDWuVgeF
w2W8GijY2zqJ3odR2AI+Bc/KhVsX1Tyx9epIfgMRElK1bFIXvwwaGoRPspeASPXr
J4oq1CkKlQEGj/zVHDD8VspL7d3uug47OElIKkC8Uf+tC7bP9mrGZ8igK4Nv6zD3
Pr/q+gqZs+rW/qQk8d5KRamn1ptsnnjk3sSGylblsjTU3B4AMiin6O3sQG2bVpH7
Zo98cwnZCbiEcs5jJPt/wpm0SrdpDRlt8Bgc+YatdHHSpZU72kLHJzYmPpAqnt1+
agl4eQbWCczDcXpQIu7P9bbjgQmx5VHEt9VfBOwxP0aOmf53nhYheIqybvbCg8LD
i5dtUIq4Elm86NPx8fjkFpg1fA529eOEtq7yDFn8NIX02CFuvIA93caCOxO1AZLO
KZq8EtaGLUDLCCn2Mk1AMqgsdzAbeff6JKOwgJkN+LAtEygRAVhl4ilVtS9w5yAe
4KeFISf3HIk3icHQyCTl5MMc5i6VblOPKn+hIDDpzoTT0Baw/1uQ3eqKov8BBWTe
kbwxh6VyaOkp9dFuPnK+AIXHTuCFi1QPX0U3ML6diuhpiY/ZKpsqXYkO3Q3FFQTd
NUKgNv31ikIWJBFLYlYr9zCB9Rfv77vzdADdYRQmSRL7oyQ5zEgrwSddelioPaV6
H8s6HCSJeS10+qABojJB49qsAe1/aMjT2fDwdPfWyflLs4kLQjXMzfdtAxn9Bk3+
gtzYv4ptzZKf2cyhMSfdYMQXJ+sjEmmKauM2KplQixMQwIxX6Fs/lGRobjDTXTHQ
QX+kSlfCxyPHOK9ljXQ3z9O6Mre4+FSeWS5ELhf2dKwReX6CxkuvltjnX9qM60uF
//aGi8nrw/R6vZccUTmz3cApt/5F98kAaT2uIicsN1njkkPNvm/ruoor3frGE2ZQ
fEc4MyI+EOsrIjn4U9pjPst/6hKzu1XqgQcVn5IlWZ7qeOqpUjTz00UKn0UixEW9
mQ1VKgVfebQq3w6kQOBkvsbwxFO0w59W3F4H8IasK2Jte4MgdRuTmZ8GadubJMGY
IX85HYKvhOh5wS6ilRCWnUCihTsKjKhsf3ncJoAxQAaBlNw5E+1r+N09CBvh7UXx
Qmn+xxF2d+x7lsyYaSUx5+/jnRMEmOes/2ftiSnrs9TNI3DgJbKASX7CkTUdtVyw
xOdWONiaWm6zjmAyuHDQe3ERyjHcm3mixpO3e190MRKYeAOBEZNZ/SQcKqmeksBg
LQd3C9gqd0OHI7fUkifbjEYUoa/YhFovE8yseoG4VBOs/15IZPEvi2mdXPEhgtCq
uL4y1E4ZcnvJDqKh0lheY2hAOCNXT9ymUL0WvBF1y9ID9Vos6CYl9513moVVPKBG
dl/uM9vJMM8TTokzWTjagZsl1tmCCr1BE4LwZ8Rb7Qa0hfh7yYucgvCV4uCaEo/J
GvPzMaDBt7SAi4S0UL7Eq+FMicwW+YOcF4FSCVUsjcZsNFRVd2S306n7ZqOxxkfa
l4Le/VqamyEfLCP83EXyrGQFeWCKiq7bvgBL1Ain5Rof5PXT+eHHfEqVeTJMuGem
MBL8EsqZKbkp7U6wwnw6MLgQBEsO32g7JfnmpI7isMqiyqeChMh3S5hqRUHN/a0I
OquPfKAIzlB/j7EkpYj1jnnCu4SkvRyuMiCjotzNlOHjw47V7j997w3/3PCSiGu5
+91F9cTWoIWrFKQI8dm3SvR4/NPoKp/2CikVVM5bb7IwFhqjEJWIcd/cx8QjtARo
dQI326FvLveQTw48e8QEGItWQVAalHFxh3z6Q3yXeIW3/0jwAeh2yhdB+A4gskwd
07mfsibJM7k1zy6ovXDN2LJVT/pqrpeWQP7cZLo4d14M8woECTUFMM3sNy9tNbl0
vhQhKEkZgzGX9dciiBszl2MySvanqDP0z7zw15FivR6XQ767FMqNQpi/ZuLWWXT0
84M+iIYh0Pfbgeiz94QS6hAxkCvAxsSFg8ppgEkjOGtAJD4RbVMDHvg5zeQn96FL
EsdpwaXSK07dpaYEaN4aeK2D00x6eB1EUVbv/+MXkd46uwgNzzuqmE+6NAQbkJ4d
xTZpxNyP9TBFwTVwkfFSd4sgXuIrcj8QIG40RlJDBxy8+/ev6eyC0Xc5EuKwFixv
ME0QKzTxOC2sXLLkt81aW8IOol1wz8ih6+WoQeoXwygMmdx6xB+p2RJ39KbvFH/s
TkmNblJG7Nf7mRZB3dxgOO3sUtDxOny23XaTKjX1uDiJDqAt/lFIZMO5RsUlA5KE
GjM8Aj6xwLAFUakUsZRGqIBSQ9KiTXoqg09Iokzj3Bgue8rbflbI3vCZe95LmP8z
VEgXe+KfIZNp39md7EC46EidFOp1xU7+lCfaxMCPNpn0V/+u/DDfRDmknhIf8lHb
+mTODu2oIyykX5k0w3KTeZeEhRBXLwbOxGF1XRhow9xSerk3+dY3dpoPro8G2JVN
E8MBhGtTao1FNU9C+pi/IefvQZQMx5g0c49hB7+Li0zlHIQlZUQp8emGgFnSKCbx
3cV77RcYktEL2zrYwDq0TfQRyRpDhQyLVROGIFZvJSh9niwXnwQxOFP5KzYHr9/1
hCm8IIUba8KnQZ09+l4stEDqD81Gbh5N5qET9A/ThnXHBfPKgfKOw48jzkptwRaw
YDVwP2EPch8YKTL/L4TIeBSs3UySmna6VcTq119LLQkPkAUlHuH48NYEVN2kqfxn
E8qyp4yyo1d/upR57Y5fzDx9yj04+Px4JLX0VlzMxRE+k0K2KpY53Jkp3E8rGgcm
dMMgTv+aERDNHlUwYjYmVVCo0xAoZypwnxGbG6FhBcgXWKx5U0IyGifjMiOHB9ge
UEH5sRuZiq3LYEVUn4WcsZNoRAT8Uf8bt328RPKT2zT6nCd+XI8n+RA/83vspsOy
OOVW/LDvMvgEIkIBiuTcr/4YKQpo8TTM84ewfbiveDLEnyIllEwf9ZxT2Tlhc3zP
8HSgWT/DJ15EGe4UZn50ccBifLpZUDRbTiRAQzwk0LpQuspxthvHFUF/SZQvsWUx
wiC93Kx+JkuCT4D4O/fZjDHEDwj9ZM9zNdl2jaikocFDGfEp92D2eVtOCWV4imAY
ALDnbTeXQ/V9Bah5aETRQ5onmDppbAhEb3/t8ORAwG4DuYEHFrmNycn9mdQwC7zc
uDAd/LoHDJ31rvGc+yz7brbIrPLXCjGRRluTuKNriksznpmVMJtMJr+TxUajLH/G
lRMcU5dc7XcdryDmKP1WnZyxqOrzB4qsJZEDy12QFzxl6M2YUWCJJFfIaaR/2cIS
0Z17dEnfgxLh0xqaqQtP0G5Fly9I60THjMHc9uYVGHkuUnw9koTzRLnlMYbl4jEA
/msn96m0TQlbWhZMHxMhTB+TeH6BVbl/AV6Vje+M6H4f/3WCQx7E3OTkDjH3Hxg6
mVJy6RSUIqKKgDHQyooto+zsO/3+arFJznKrr0fh1BshZRSyoxKVTUYCJqfcOf0q
93UULoMTVmQSQdrcr2kpZTmdGCyLbTAU46IkTfTPnMhZ467Hkbq9P41djqnwpjy9
F31niDVO9tFW6wqiIlhT7G/oCNrxVKcvao5A/vtT3qizjPQEw7Nt3T9CvcnAHshd
kPr/tzJ4vkqHakrc+Ls6kuisnOX6ESccFudtH7gj2WlzG/omLKETtRuWe+mU0e/m
zKBMbodT3usqyY3bH2gG2uyNixlwPgG6m2kbVjoiNum2jk7tEqfl+O4LnXJLMIAu
meNH9r2dGvicpndRMz2yFeuiHlZMgKbG+9RUUAj13f9OCyZ0fKciNbAeT0+hh6UU
E72wWrZY3ItpYjbcHedhLFs+yQbXaE8bHPcmhZXL40zWlLCQG7lNve8a5nf15DWc
AKf+vBVNB7szimiGFThRiqgu6IiAhugkpmtoE89Wb4g4j2j+nj7jrs63KKtkDjvc
KLSiYZNfC3A0neAhvelVCss8RyQbwSfjjEq538hl35xZItMJnwJT+Bc38fpIE2H/
Z1q2F5kmqdy39BdtRdyXfigp4EzcE0Hkjc6NujRLuTVAF7oRMXk7iTw+vJUqHx/p
P5X3wutyrSvquIFaS5zfJV4PKu6YzlOPUZrZ4ZgGcsaQ42xnmEXDdEDp7VlEFgcJ
TDo6DFp0ISbnmVDgzPJ7WjcAhHEnXXSiUHehz/8grpPOFr50Mr2D95Sq5LW10i96
CzRJZUOeIw9RNp/Jgo8UFf9fu0gZ2ZCpFr3n6ISMTEPDHdw9akmZWhj3dFXuNk/1
saJbK13g6jSR3X5uaWprPR73YEnj/MFaQWpxVJ0+0cBw130qouDHL2KVNmzguI9N
1jpnBfAGoo/zSUWH9ZRmgNK8IpQNIcZOEuPM7j3OQvMZwTGmYpHRuygvmXD7bEd4
DVZjeseS+dJj7jgUnWC+cNEJ5hVOueetInNyucybspoKOcCh4tFsoRUJqrzbuz+Y
8H+TVFSKJ0zi4LJigslcXUEfOPqdDS9yQ6z0zYppbiO3NMktW1LSrmAZ2wi98jD5
LuZmK0f9eFeE+V3Ycjoougo9PB6ZxQyKm56E8RTmrZ3m9DfZc2OQaND76AgRLgIA
SZgdzvjPf4rvIzUy7AdqzYPXOaA43+5ZxxRxGxnsqdYkA96C2oyRpLx0dq8LBG7o
4DC8NIwaIWgEZXzZtgKwprb+CCwJLgh73bTGRZcQ7ByKQ8xSvfjpNAH3jZ4l7F50
XDJmF1qmBJCNPX+WC8KxnBSwBA3tyzW1xwXdOe4M95Y3kzb1lDN+wTajnPGz9WRB
5ASzKnoZH2K7frBTWiSIz7fjU3y86Qaz1ruSM3jcipySoiJxApATmn5iXfXBRWWX
XpklIauKTHIO+rLzX3KTirn0RXQuaYHjKctri6CkVFMdJO2wilcj+IxVoZ4jQLL8
w4ZAK6oL5teM63YioSuCprtsc0F3zrl93jyULqTadeiqlGkYIYR+/AhrTN0cN12K
vexRnSKYDrAcS65EQAtER/ckSGtxdtqWyfcyH8ho0OA079cCsEtwJ6EtYKeI/m/K
T4e2vF5VKyzhw37Xod993aPX6LCtmQhouizIPtztVl3+XAVNtncSt8u1jH9fUHRh
SATGLHwVQEfUjShbzbdaQPo7BsZJIrNqTXcE4zWvC4XzPmmjr4cNUodHOgjfyD6v
A6eKoanT6c05xs5ePCeqVNtu33ADmuNljivmV30qtL8KmjRtDpGg1aAFT+yisf2x
J4Do9WIUEC0GQb9F21Clo8+nysb2Abppl85pj6IUu23MpGyxh5lSFjAEFrzdhukF
Y+/8zWYb0IzwtuktDSPWIWAHn/0VMKW5aJDjT9YBqQM7p4kM5fIRp5Rq0sGBhtdB
wk93UU6/4hunuZfoCmWNx8ELEEtntSBgf14swgLZJlPneljs1Lxq2Z2VdK0C+s8S
oH5vtwOafC5qWNikiU6XCnqw3ImPigM+5LSpzFvIOgGZ4dTMKXEWdOU3OTeyVTz7
ZBxxIAxr9d92AUdhoKbt/QHHfd8Sha98/pYZNAtVEXpMEIlOVH4PyhZ7an377aCr
0WhjrvJqktWPliE3MZ6Rmv+IjOI5o93fdK3ivk3GKSnTp+Plsq270731gsjFTDO1
RM6nIDSvNH8rpN1dMt0R5YsBrcX720lt8uiFmA2PFeoQxEXbSW2MfotOCRFYhnzP
zhYLFKJnq3DrA9U8BprYxCKwqjfY1bxaAj9zRhmOXpT2G2/0g4g6DFKW/NU18+gv
HjSdUVvzU4mZakXI9+T8em04ARBRizqZkpdH+KFQ6dEfYBfKhduUwOOhBQJ1g5wh
jeJ0lxtt3VbEIcjHd0im9y629Blqy2Bx3NwIYsQq+zlJo9abqz4ndYAIEyHozAtz
StIIzMyD2eJTKOVBr9JQBKde8HdvyOaLs1FO8u/gfIQY6WQFgnh9CxcsA3JYAD4f
Mt56Ble9f5SwZuZ3ST5wpffdxYyGsGFC9x0v0vU+2zildyYCHGTegGNZAdqEk31o
Q2YBpjwTHMvRqib4l83ZAzLWbs8gglaFHwggXUaErJ6IOqMrLNzH4hQhFhi/9/E+
cbjBZgxVzKYFIcWNKgEHA6WakCjyfOoADiPUNtGg/JfCKscqSIG4B0MRHCFepB0F
+M+UQdEyohKv8UszUCqfGVbkN5e3rf4A+TubicoFVViBcX/vXR79uixaCyBZbZlY
G4UODP6NQU2sWd2kOHOnFZUMAv9teLLu6waZXpaFh2CeEwC4y3Yrg6hoxYaKuRSX
UjeLKfBLFMowBw6ms5yVvGMsKU8n7Szdd1mEZ2t8kKOTTaqrLRyRBOmXpva2X8lU
GYqz0YA3sQt+mJb10Kq9+jsGTcFMssSXTSr5MQiSB5/5pEZvlyKuR77kcabs1G/K
jhayg/rgB26uRpfNj7Z9TFd014PS6ET93j0fgQff/H5g5PrD25n8irCMayZeZWDX
js47EgdQW6dPJkQSxnr+GDvDhz4F8R5f2t7X+88Axh5ZKnjhrulM62y/Jr39SSd4
5J6VQoCXxpnrsXzm04z0nrG4FU/cXCrKqrvDNHreT9v5AX9kqxndrMO/BQBj/IRP
0OjbZy61vfjKZ4US91wwwAOXXK+OaQdjsiz5vARh8TTeS8G8OQs5ikaJcJ5fmRew
EMLNHLufdDoDfu6X41GTJP2KoTgwJ63xrOJ+NV2Y74GJYAlyTorCd/iksRFdQjV/
BnIO1pT3oailItiyFeam6lUA6cTYd7VTIR3iLUkLCk8lzx2s29rP0Yq2plFYVvcZ
jxizU1CPksM55BCUjrQSlnHXdiwuoyE1uaUPXfcxBWdbcZzuBFKJv02+v+BMG7Pl
gQDR6p93Q8Vuf7E/uuM9nl9MmDsEAF/djmDFzgUtH+XOxpd1smp0Dz3oXZ40PQO2
9hpO8yQ3butnMaFLbS7WS206tS8yxRJu4SpOAFcrV6c7yfy18wMdixMdx+3f9Is0
myB+bX9SxsWclfWiPMuu8ju0PZVhl6jGuUFjlb9G2ThvgZfB58fIjMhxsrUcJGmE
KypFUZHM1TkpMD5exHEtbWN0gdjd9QeoXi5qEzr4S4b5jI8AeihLgwrtInKa+4XQ
4jXoDmX6OwDW7KnvmbOKWVJRZc1dsWqYFKk6Mjjj5IE3I+pCKnIGM4W6BERks5cN
EzEIAa4bT3J+g9djyhBDnkpMpkPUlL5RD9PCSEYVx0l3pTZzZ/r0yAWlD71MKFHf
has2vaPnAaGNWQkHYrmP77RHrggN90iEmb4ThUnddkj9CpwFMo/BpwR55PVuyu9B
A2W+ZcgNt6TDy/6AtUuHPp/UKnLnHUPZn64pOb8ZQ/rDlDkuQfO4UCP5+ZakmpLU
QwCT9K4klCfTgQE69hzpBZQVrg+bsEa8yM/FrkHquZvxQS+H6ZBroooPS11leTp1
3QmkADsZRsc5sTcNeNGbnLLc5tHYnZ8gsk05QGg0iRAoaOp4wcfHX9OQ9gR6riBq
iptJ2hRRwCvFqZE2xBn10d0RajkNyl6gS3G22aLRXRsU0YIkpZ2HrIugFDmGu0Du
Iytmc7RJA3IPum2sOOXwcg2ZZH3U4CqzM5d99jCcjXi7euLXZIPmSn1GWXhmWk2K
EY/w3uvA+5q6O79zgVON8dUmIxA76oLYxfiMArhqKabdS/O5OmPUhq7ilb6WKGsP
9Jangy90Q+uhQfWXWfiyxwVtlzVpot3OrQY7LH5wjwlCVbq14fpPhvxTgXrfqsJi
ScmvuH07nI/WV06vMTLfPYQhTW8wM/IbgyLh6LHmW7/2Pdzz5iVcFPuJ6sbAwPnf
LiqDFPpBCspLJ1pkLJG815jv6Sb/wX8Ysfr1v1ul7UuNWnILbZHjscCrhpQW00t3
2c886peHh4+iGgEpuw0xUux7YeOPVHNNv52YXDl/GtdxaJ2WkPF4sRD+RhrgH9PI
EDTnPbUVNID9QKbr9imM+j1i95jNZUdHn3BYx1KbeUkjP3noOBJL6jnb3psEGQng
CjdGxtv6ujPo/qSThojU9MieQvuL+ljVrjpNAUdQ8RmXLFqLy6IDNHJtyEEsKMIB
PSAW/f+3wBvVMyE0+7P0Y5dzUFGmOjSXCuAP+ivuL/oB0IkHhyeY/DQw3ZCgu6Pr
O6MepaylttB/LbgFlabkCJFqybiFCOqHzSaDN6nkSl+vJvSLnzDrUZKgUfLlMBIY
cPGII7tKbMRXtDOyRQbIJv8sK+vy/SaJ+1iN32wMQ/yTNdTAJtUV9+QpS4GVupv3
j/zu0K8TjYawwbByazDP3JZmvWwL6TRH4xBEOqDLuQBmY6kt046XmBddIuQiyw2b
7GncAqDOBowUGse9b2CH6UvLJ8XABbowvU76i9mGW+IAJnIci8WrRH1pxdvDISX9
RWnDc1T8H5GvnUeQxDO5Ng6g5G/VLmEWaNS08URYzyydnAtKtcK2xwiLbMj/KCLm
JLIgG3oxiDu+lpp0eYPTjNdOJ8nYtBnIFbCCQ9rybzuair90bZJ0xKLrFnZ4SpL4
aoCeMs8w6G2/JKizD6IgghLcoML8eFRF+Avl1J7KT3XZ7ySYgkwZ4JScr9xBYDwP
FwkN8RZ3lCvhvtBD5uLrwF1DqPNIKaOnwTnWlRf+9t85nUqUon8mZX4myXW9BvRO
svufEdnlN+zYE8ZehX/JJf4M/Lq5EhUZiW/rO0TizdO84JnL79UevOwJPpSCp3lj
Ll2UgtWgpk+geqa2LNhqARqCbc4Abh5QzfZhU/IaKH8ybwsSbaVsN5CM3jPMKbXA
O9+S8nxTgVE5iF10E1SfiZovrld8WIiY+J6Tr3MnOJ+JUqhrxdY8JwDwn4JTxJZa
TKM17/SwqtR+/V32kdSSlrIv3TC6g9YO4P82JPkpPcUNyCQE36wx/CFLUw1/ibMY
ffbQ/us+YW7Zqlh6Z2Bjbnj0NYVI90BHajCOJcojlgLL17sbcxIFJ3dif2ryK8lp
d7AUIwy+AG7WQCtL0uGVxzl2mNVkjCiNKh+GudK2oMm2/40eUSszEvE4eVAV30Cn
+nKnGAvEkLOgyHfZsY48kV8hK83aL8Vxg/E0l0w/UZT9/dS5r2QIz/3HfMvy2aG6
mFgmCP+ZlmZk7TSLxL3ux+oPUky4N/Bl7qRR8vSWAF8nq981hUZBAZH77GzVVgrK
pkx/Ff93b8qOPSuYzBkCEOtxc02C4gGV0KO5YD5BhyLnJBMypW9MvUFPCu/9oQjl
oM0uqbHpf5zDbQC3RpvRtRkZ5o82ahDLohEOP1CFkLBK8Ctm1G0G0O3lOjnWj/hR
s/y1qGiNJmZbEZMuxoyEoL5zL4m2dC6KjgMM3JVIgA1ha70GEj61aBRnt8ajGlvn
vPi5howoV5MV6aVxWFfq4LWwChUra7hBlo7GKsLXK2TNYMg7Qry2FNDgdDTt25O2
dijURtq2mgIxJDR8bJVYAHlbhvbXhXaNUZYguKzse/xiJi/ECGz06crbZt6IanEY
+ijYvZtorb3RYb4wPXbznRaocnEnQYkTaTDAHSsaLP1jZb381N1qtdAv9ZRanSQa
1kh3JOCXrt1kcarKtoFa5ZDIvHeIa3qErzInM9dsWOkG0TK4WjWb9oJql5i2TDAq
O600xNLFnHBSOJHT20rHJJyyZczjOmHywQs8TC2q5ytHkKupfKTUbzmKSvXvL44H
6Sz7R2VZNweb6j9ZvqDRfSgRuCinDGYn8Ey6HMVFtC9xSRXTOU7Nr155a65jWxIK
jC0SQf8keTDAq8CdgG6kMZqTJ/w5g12G44t7q+kpkYYXvC/io56hjNS/j+GYXctr
np5TVGYiWGSWQdQrCk6y9i0khbD/9uHppDOoldijXVsdb9KG+MlvnWpkIjt+obU2
BCrsoa/HpIgzH9VaGcBughbWc86UEJ4TYBEXXdJAaSM8RHX8C/BA+ijuVGZyAOaw
K5UP/KGQrE1l8HXm4t4YgnJYU31Nak/Y2iSUK2K2rJfXX7qIP8j2syREUQYapfZW
ynZ7I+pL0+e0GQBNicph9DXIwQ0hCVGf7FytWM0rEeGVnd2HQoj2uhJucT/1oCeX
31tc0avw4afmCXsecqklz5PJj+WsmN0rQspjaDVS7FBhw3A7ETPJtOZw44sI0rrV
Ib8Y+YEyUjmjgfGuABBqXWU9HfMFfbjKGOtYr5ezPPEJVmc4no9t6OteROJMHI3g
PJisyK7rC3IMzLKbTJ4h6BEGt4sK/Lb+lWM6qJJ1rm3y6XF78hMesKTzZn8LUahZ
CHelLJ1Y0X9qFHhP/DrF4AnM1G6QvPABWQYir/Pzvdhv8VTQr5H3bGX0/TuI/KcO
RxTNoLIvXx6kNm5fm9VyD/OKHFRg8UqeQOYxTiaHq8REecQFpy2GIW8dlaQEZJ1R
tIEXBhsO8UtyrIxACTXNR8MZnWbKKrlkkAU2AAhXbk1ZEvPrkww6stERLzfZkV/B
ZVFPrGTzDUyApgGuaRjB6jUNDPN+pfEUHV1BMt36h7QhR7nGjkqRfPWbVHEBWy6j
toO7SiV69Pwdr4BBv6o/M539Ymbl5AFdIdBPkt0BFuA8L+u9JJZI4otqKaG5Tcut
hwySH5gEhXCBgNimpaSL2dtsI64tfFAzVMEbkm94+1cGLFzdOPZnRYvPUkmFtKvo
HhxUbEhOGI/bNuUjXLFfM9s9TftjC/MrN4RauABHrWFXTjc4ClG1Fl5NBYMUS0h7
v6FfJCo+SpFHg4Juzuyy6snKzJFwxu7H/hSfu9jVfN1Ep3VX1O2yCHe7bNTF6pIY
8/GsPn3I1PQogkx7vdgEQtw9eCIWfzwKO33xt/a3gD5RiFouXRT0MD7U5PWjEy9R
JcxyxrpT80RWytoYNEOcj7pQaGuE+ciYZC3Go/dwxhuq08RhgOpWccipVjUgkSq9
Y0X2qmJw6sJHm6XHzMn5yWQBoHNen41nsnnwkWc6j4KgMgWJtQrq6SYa2f9PCOIO
w3/lwU/6uidYjASKPbFgns78SwYlYxIynPokCZYj+abng1M3CM1R+po20jHdMMOd
cwxNZ3lTfLq/x7MZfPVa7IVz3hBliLZ+b63AwdQG0qnG+S2fya4rFAM1PGbNHlCp
71F7UKnwF/HiatdwrMIdNRkyH0XQcbBU4wTmtS0Uqr7Y/T2yj1QahPPrzr7I01Rj
ok5dv7smjpKDdlfYwHIesKfdO93Jb/VgXkJSuu4NXcWp2Bflh3uh6k4qLaYbDlPc
406zF0qCZsUlAjjcufA740Sy0G7+GzNpdOQv43vJAty5p0BXr374mXXc0jOeeA2t
9fu+Dq7AeH49grd6/FHou3Hsds6HaJoo4KLcGyALgY97QpZuDzSduXC2ktQyeNCC
4CcVdtErrHLwaZGYCr5PhIwL5aDrLQqCCf0ZNcyYwy+F4fKF3OerAOUoX7UevmWY
cCtHj8C+ujnPC7NlE3DJtukBqlmBIXVFcBFEE5o3Fh/M1/YCp+CerkxB28BzQOwM
OotOFyLG0FBKixTC1RvrMovpaDCNs4LbIhT7HTHKTUoc9/l7wRb6MpETGsx6ZSKY
5fulgXPbtsX289krYfKEcGyBQ/InDx1WB4dumP6i3jpigm/kBvM7qPgblkXBrm5C
wXtOURkaT3n1BoW8AtI3p6XqkZEKFDTIL4gheJqF4GnvuzuI781AXengrxMoQejP
JvTFAB3v7g1pTTQhDuZV/1HTFgWDsXF/9T+eEN7ijHW5l83pSwg7H8EbA0VMAm9X
auymx386yLbs26lJ67DQTc2rl/fUQdUPZ7rjYTVxvTB/qkkpKWigiHqMCf5bIREw
sd1rUzBlMdtKm3Ftn4BmOX1TAtv7KIBPS+yJNaVC2nIT5u3Y/xtla/6weSoxZQ4E
5E3H/2j4EjNOgFmF52CDB4Hy5+PtHK5AR4nS9PJaexhX0PNzGh1nQ/5fvZ94Kb81
1BIt5ARZzJCMMWNinB+aDx2W2kjVUiNDqE0GpKl1g/gWwE4uESWWU4IRkskDayIl
9BIUFaUHt53b2zk+gkJ1XS9HDaQ/5lluRhjpOZ5Vz6qHdtmE7UEiJeX+Qi6vCBxi
VAjG1Us/yOxaqwdvaIoWY8CubOmd+aovy6aRzaWy3ge0clsePBhIKNerRrRtWEnP
pNCqLhzjcwcK6hIj3ALk33WYNiPMDihalvres5JZi84JQGrxdHsurlnGrbz0hrg8
rEu1tN/nXZ0aRhVgPoptlSLd00jQrsZTmwYNl2GAQr7DNcrfw8ekMayaG3hRB6LU
86qbLsk1D9WREhwoSkO+bQdafWDwrcb+frpLDX0WuxmRE4gKEW3e5+sRP4oY77W6
dywKdxMaacCveSzVYdCidy8pQvifiSw4+cDZ5kDx8puS7tJG9eVoYB9zfz0H2JKn
uqz3Mb7ly1O5XrVxmkLWqahvtPNTlMnt4uFbwNtgxl3CUcQ+RNiS6hQZIWnauc0o
hFxV49WmxpPSyZ3S3rg4NbRFMiF7Sds6qdoaeObV3jPj8cmDnMO/Neo7k3jKDnmD
YXQ3pF+7+3MwynfrXUf/4fmh09R8vhBxKQROglAeIT4Xu7QPAY2mRTxsrGXicD7K
P2MRjgipiLF5tx89W4BkcvDh62dNmFUtZinIpCBtuWhF2WRliH/zsXiQ2EQQs2GB
3Ro/kIrCoYAdQtP593VG/cMkM9c0ZMGID/t1pMeDhwBc04CGCsyI7+iNZkmH9ew9
/NiiT/F8cJnc5hHTFxVgScYuBBTYL/qcOFhGIoYfUPOquSYA3/OpDlM33ZjWPU9g
QJYEi+RKUT2upfemsQKT2aDwFCDk95HXK2uj/k66lckrPaWYVTwB8yQdcehDs9o9
ke3BJiAi/heACpWmyuB+wPzGFCRl8o9tKBzECnAlajOu5gFCIncwUfGbyJawsF0M
TDOIBX6fctYy0JMGST+SomfhG2b1JABUymthi3AHSNjsFrZozatz0rV92cCw6+qB
+TStqKNqUSEzMIexxaQr/cDXysZeSncqiXLhcPFNQ0040cw4dVGn1Kb7uWAv+PTc
E41IEgrH/GwoWExOKJbdQl5H4Qrr343X7LvfTu4hHc+KNmaRu8AduhseRQam2IeI
N4lzew/qgQTOQ1yoi2bHhQvwgqf63ooZeISX77IS0JD6tT+p7tVR8ndi61VYd/Rf
S4WWtPKhIJpi6VUr/wGgA20YSpYqIVyTC3pg/epzq3xImVT02502UttFaXk9FD02
cpXAefdOKS72ufg0xUgvEIhma5MtChAHMYQiDIJoO3P2mdJuhA7NpATuM6dXjcU9
za5RJ+42wzPV4HFafAIwwlqYMZR5PUnBlRQPBSs0tNnW3wJHTEjWfAtxu7FhjCcc
oxf+cBkKE0cG0GwnUod0UfCa2JNwkue7NXM6whMri0ygrDnw8p7oHeQAosf8/Lw2
FonSjdtE+1oM/gt4zcENfrUmCZ3buSTWsHZ/uJ1YJxvRCecVp/Aj4UmauryNZQdl
Cr46pn65Z3chHc7AhYSXUqAUlky1isHfsa38eLRPtWYex9ChpBRCdsohkDQMYUvQ
PNm0hGAmk25bZqsV6p4stmUkMAlxzB0fLAAgu7q+Ao4ThYbJbWkCrXswCTOhmAH8
jL8a0G+j0b8X11VmTookcL84StY+1b8qevNm32er033PVbhctGtkO3AV1ONeL7c5
uF+nHGb++hQ5+M5FLeJbVHYY+f+KJbG206JuMoOjK0bvQeQGsTZ76tpW865cmWJv
GlJSY3wPeakZ+QAze1SwQ8YzC7wH3MhjiXNb0R/ZEdiNY9h3pFaFkNStDA1zpKw3
udCn32+ccZVIr+CVZMih5MIhTc7s0cswMgX67a/dYRpyaFqD+lzx5QwRSc+eF2SE
nL4drAPliE1ZgpzssM9kf/Y4+jrDeNfQAwTPG86lguZGnJvrvrDD7F6h/cMw4Zjy
rG95V72Ek34jq3xMKu4mCOykjI83M6sz9wzKlC7IfjdvgPThnXcSOKjIOaFsx5Sx
++WNgadIkgqhRBZvCBdUMibKKWPjp5bAuZLmDZoL53kDYRlnTOWrziAg/RujNQiq
t7WcSmRt/kXrwfqrEfZQKIdq3d++KPXPSmyfrhrBmTW5fJRhF/Rduv6WZKx3RX1+
FKuvtYfjgQIcStWZ9Re1JJE4pRzcjFxI2IVfRK68A27fJEU/6prmL6JJAfOKDjt1
mm5Co3Itx1vF24At/9WMIteLQBWY4RuA1LeTUr6JcJfJsoOTgCp5tG68ajIDuOJC
omc8OjjUgrCoGI0iopKQ1XyfZHgFwVAP2JBdIc8mjo4S1uJ1JQ7UnoKlbvT/Ts+m
O6qt52r5raz1OtbIgFMHjkKDZNYmp1pBNGaA8l1lNqFECF7yv36rJm3pyUqKMYou
y47XR4+URzYkbveGPUGK7myHKGboKWSmvTSD2bATsBFS5izA+U9MscxNo5DlHfXQ
MJ8EyciF0rl6IcMmkAKZEaBL9Om1KY/0FvMWnAyYUXZaEu5TS/JWOSHu//M2f40S
ee7IBP05XL+zOTb1rCbEOvTB9/psS0KI1w8KLrxPa31lyvgExjAu3KfLccO4TGXe
gQ/6viaar7azx5OPvVEE9uUNpKsC7ohGS4KiNpNS/Hzg517YJrbYxcbK1qG9YGeL
S3RerDs6nN1LgYMk5mqRcopzOiRu/KIzk77ow/O5p0ox6IzNzk+ApV2rpcAe8kOm
4HoROcba3VO/s+4ZobOTWknhURhCIc+BfjbwAgxLp6UOZPqWVh3dbu7tCxwFS8+x
KSawbT3KIjtVBezoC74OeiwojroOJc9M6RT8fGw2DJnOlULYKd4yu0T6P23Ye5I9
/FbOpKSWAZiJlaOe5fbjsZslY7n6p7spnc9FIJzni+3rGu/bPI/zXDHdiLIXXiWe
RAv6Xb2mmNCbOWpCApElriGY8aEx9K/RmW/ARKgPReJHZA99MBCe0ooKXb6vcbMZ
yqz+fLnjTNpXy8DOqm86ZsFJE9ZICJvHj/Dp4Scrz74rAlZ3EVOEkBdnf46MoNlF
GoqaBKYYoOBtFRe41aIIwiunBw36Uzq+CjKuNkS/kkRbNvW6h/q86ml73V3s5P7M
AZSYcx4MwUHRHPOzBdqTdo9wFhNgy3Q2R+Pk2iXFCL1Q0JYcFcvv68WVqv3jRNfO
ZF+BznUmuy5YYHmS9Bjafh/8Xwa+WYHhAiovj7KNl/oeEQj7Bw10Q49jh6TqzYRt
WqvKbFXmCotRidokVTxyR+9t4qpSF52sB2bomLe7mYDEuKf2+RX/Gpl1U+Vq4+Yx
nj0+Lgo/lC1Dps75POIJRvDUxGcRUxlKx50M43cp+3B01eQ2vTaFtW5cp4/qaWyX
n3cC+hbdDVOd94d+qfC946obxcJU72Nnu8aGSKgmLG2/vpFXSnYFwMe+N5VzX2Eq
jcO2qxSkvcZC/I4a1o5T/rHoy+lHphSlt8e9MrJYPljiaG4mg4qj0zS8Ua0bHTZR
T3fNzyk6vES2En/v7EdhVKQY+jDdSur1b4uqzJqQ8Y4E+0OG05+Xd/I9tDsGDPaX
f/DSq730ju6d1tJuY+dX6SwKZjWiyBjHkvtFcNYnVjZJXuaP2jOS9YdwNVd9jSOC
LjmIGIDDQtMzEIZ8MKgzvo82AYzYCzkXN7kGXsNWJo6RYTdSqENCmpjzPBdx2J3F
t1A3+B3eAX9SnIjrROk6S3jHlGvq12AqzAaXfEHg+ORnSY3sCCR81z3x2Bjq5bx5
i6uexX5qqRyt+aa1hp3TkRDkf1YbqFsmnCt8QP0siozjamnfqcYnvZ/LMu/hBAEs
tNtHr8m9Z63yThpsrKudrGh5WBCnV/xcx2YE2FrEtETHymqmF7I2ulv90qUL4uTc
4Ai6MFHBSwPMsgNXQDsdIpEb+EsmlpNY8/BhlSPgbMYKlj+C56YcZHMbDE2GBVTS
5fRI8Q1xNyzVa4jMAVKgWFiXV10enmSKpffRZcboWOn3Mk1ldB7xRI7UJOX7/LZD
CZDa23zj7len/vx2ow8cZZ3LKO0I3wa5QVfKHKWaho+FGDnGNpMPJYHtrxHFOQjk
sEbD1zy4jYs2nudJxSbCQ9m340CLUgRPOfTBkUxrIpz3bobTFtTZOn6/CUHlwGvY
9dORfzikPWLSIAzcsZqWR2CVs8xmiB9RhM3Y17U7rAGEKQ3F2q2zFpooxgVLNqtP
CJtP5lA5FLxuAmK9qLfjDBT/PyMuPDXTvB4Zo3Q0Uq4qI0q5T+Re1hrqt3Og2+UU
zLWv+5y5etW9t8gIaP6/wMKmyiBktyYCpJ9QfcUFQiCifrQDG089prYy5b3I/4QS
aIUxO2ziRHF4bR7GcM+tNr53A0wes2j2hoE3Zb2MNK71JS1PXhbelKKHhGaJYjnt
phJDLo9emG0j1FoITQ3V2L1IiZQCKku4bPpo5EmeDrPk8vxxJgSAI4RyB0YdCBmD
FsJtlHA1t6QLDYcxLEs0msmHTSmbU0okXHmUaHacGVo3XKyOCSrOnYB9aig4IK7E
QXUhxO71yWYJsBh642kdBGE+R2Vn1oy37X0tUiE6kBbkZG/XNZeCx3Zst+QQ4pAd
v9GYovY4rNT2jSVTPdyq3mCieXS1K4YjmxX/7ITdqfLa6dGaIq/jahvnkMOOp7CR
+Gx8lZyxP+MzBbU8dT2H+CQuw3mbvcg0eDq/XvaqY46yHBvcXgt3eWVPUMZK5FJP
6q6na19XZwxkx2m/iTsNW7oqpqnXt1mLBtwpFlWsMdBOfjZ5Y51ZJ/TvWto3p9mQ
C7hrFeYfniV4JrUv7nfXxXR3ruBW5rEw1b36Jb1HiTD6lForA4VRIsn1zsD5IztW
pYdB/wRKHqSvbncPZhkDKpqcisW9d1PKNZB7kAF5/wHdCQZgYthvGQzt8afjJ/Va
D2BYNeEv7PI1xPjaxVCrCuF6IdFgLSEcC8z6BwY3fCa7pHSGqAWATYqvrsOmWaWr
EFHt3Oc9BABDgP3wU91Pcg6CXwqGbQKhTjmHLn+T0YWOPZAoN4eaCIR//sju7eej
3phrh1m5uqI6p/idvIy0ydK51Z937QiKNqULeymgRjdxCNnHBE6zkYTl4eOkwEix
lJX+Kp1aIWqVBrcYWIUQvyvAyIu7aUZL0p/CwwVdPafcjjqBXCdWJacuOuPVrTkJ
Ze68qKA04FFESUl61Ag0+feNHAh6RG5WR4upgXlMO+Pz4LvwhcLi6Oa0EhOrhJUf
NFdKldATQnQZq3TU150Cc0aE7/cEd4ehEELZ411Qk0cR/gPyfgMJ89OO0n6IO6oR
d6hAsHY/5oeffdmGPG7afQNXYZwLTX3SYc0w9X84UtG4Od7GzPlf3q1H8lB64RPI
YQGpzFm0Aqmvv0I8XkzSpG18jIg+ms11Et7mis3WpW7cnqh0MFi00fe1eaaBy3Nn
LiCFunvuHJV/qKcsmLzbkFlRWXgmxXvgQB1l36vjZZwmsQumSmPWZak0sggp3aPm
H8W3AW5vi1/G+npCQxNZAbVMDip9jp33d4K9lEmoMKTqXA2SIC2Cf6U3zKYMGPkU
BY5jS20IA7VwWux7H4k8DMiFU1tWg4ifdLJftqyl/A3bCRm4lPQ0xZprlox7JKHQ
Gyfg9FMzH3icFg0i+1gV9bzDiSkk7DruYmF2U9kK2DDtcb+E13y5C+7sdMt2Jxlz
sus29AjngcrQDnxhKwv+ahD6fGtnLgUlp+lMTr4tEq64z40WoeC3w2zoRzHrst8Y
ylyJQ20/c0jT7ouZWtup3AvwXZrEBM59CJeBKFaCJTZ4vFHCOaSQnV2PhC+9Dt0I
4ArYKjS+/TU46GJHv+aCheHyrb45C1FhCJDGqRru02PsA26hOXP8062yUUFxqDOx
IHWJVxsxT5ePw4N6bXgR5TQKaJxVnk34ham6Zt7/lQHYibrA2+FmNEh9DQ8g3Elj
RUCN0M5svOTa57n/fmn+27z7RLUB2tT6vqqKNMqyawOLPR1Xf9IDs5x6bwBw3dzD
+F/m8ZR2hqWKl9ihm/7bHONJUkriJ/14FR6QYcTEVeqkC59rg+iMQfkQoyphXEhA
tu3Ti1QSIkUYbEoWWkRB08npAOMV/PPtokfE3aiN6sr6KLNhyNu3FzxGGO9Y4sDF
HvLrsxolOytcvasyLdb7vRxlrO68S1MsS8V22eJs1CpqvrNpLBDkX6MZIMDpT+E3
A4mVNPqU2KLXuXa0o2J2KiCmOYDGRvq8BYk1cnazqaRSU5hKAbSEpcaA1A4lWZIx
0zrFN6z5Ar2b+wizw/gcVQYIjvAOoP62RfEwtEnVQe9zABb8lh9vqmZAIraFzqVl
HZwnbAtpjHghQ+06qJxBHuS5mpj5kbIuyKIfP45k0711D/69t6SpZJ1tqRYFzd98
GOByk/XNz7480jML8uekw+vNG5rTsvLdcbCUAgYWySkS/wZB4D/NW8YkACotcSZo
WzXzp31Y/krb/AiiEPrl9jFDu34z3NFvJbHtRkc2VweO9qZPIn5yZo01cWJqxfOg
MfLkxoc67mchzllAvJ7q54PU8kfJa9LztV8r529yXro/PIqRBNFXzRxXKK88pKNv
q0Qvfifza5Pp0LJUX72b+hmtb5vZlj2Jwdu0t8VyAyFg/BsFedkMAL0YQ0NDfNUZ
J2gf1sjaKx74FlHDmCib293cR3Z42aVoZQ0Gu/ScRnjJnjXuJtZbudY0unEL+1rv
XHvg4zA8FXRa7r+zVB6BpUzkvi1JGK7LxQtEcJyr2SdmgajpWSRRvGQU350zxQ3l
KkB8eGlJBE+18R68yGwxAy1RyZxAQTdU/+HVmOce05mq5xyri5i++ZyPA5CqD9EL
Ozglk2Ktez61CZayUYXq66dkuqkuMJ4AtzatVpECYEm9hSsoZ1dkaUT9zcoHEGfU
6wdbLE+W8zUj+yHK7mBV0sfNiFgG9nweATgEgnxBhAgWg2uL/KuUMCjyxF6uyV9K
xbwDQ+IOED4mNPoaeRlk41VlEpDu+18GGIeR63zHEDr4ghYRLUAnPhS9DttEYXuj
Z1zf9aTZV3YOALFu6vF4LAQ7fcVZACUxkFTMVOvHF8YCa0ybEEFmIcJu6OgydQAR
pCkVBdgUFHEcOMkARmDOafUq20+dGfbq5Uuvmcc7sUVPl1rYKm7/lEJtoy0ZtHIn
nfztNd3fzh67zcauxB/D70QR2+8SV5tjsRmojQDHGGz5tbp/wyMXrBy2yN/HvboC
xQVQ/b3zp2/1eLVDPft5hSrwG+rGWvCqao1Q5z1fhek09BFPNfhs8xTXaoEnan2c
6FlOkQfp/vurrMIwTwdwd2kmna0GPTF2yR0AfTKK3b6/qLV4iTGch8d8J0nG4gY9
OsKvdWlgJ72OaBQf55YRuUan2OSaZDmwpEqf5N0E+kDVBTt0Nm57sPR6zcTmCMlD
Gy04mO0gZSvodzDuLWxvw7sRvmYRoMtM4LBioTTsZJGyUzz3hGoUB3rGD1EJ6yKG
wh0ssZ4/nlVrDw7qBg/MooxAcGPUDfQmgXqdnfzUZVjPKKh+OAzdYbn2v7eRvFsi
eI2jbi7q/h2hEknehMoNAN5MVg9g6bHSSz4HZ2kt8ziHXtDSkzt23KAX2cqG1sJL
ZlM98HTs341b/pIUbkU3d+ZjpmajdoKAFMFZSLXzVTsoqZr6KhUSpj+f4Zzl7mTH
+619wx/LDx/goFzb73fwdY5UWYsNlaptMAnCfB0xZ15VMO8dKzRDUJSVM0YIkN5O
je6mM2R5SQT9gnnHcSNOwZ6dkIWf8R51EsFjB+4miM41ubjCrlDyEOHw/uKsTpoB
ZQ7zxmGQxbHHlLSlogvsYDou+g8h7AZ82G/CVurIQRtswA15XHAp13JkzYLVtTjk
/2dSFOntM8Mc88FpJS97qSG4zdfCmiK96eiI5KpIkmg190+bHZ0WEFOIw2JVzuun
gI4vRldX0oAvLbuRMptJjQLpD9RSgpAs31JVVG7O+mCvVcIlBB/2reOeGy8d8aRL
XPDuOzAZ9mhamm4JdC9MgwAdybFMN5AoXPnvUi3omQuBJ/FNRLQCYMYt+KGkzc6Y
Z0+7xuZWM7/oXC6KN53H60KhtB289GVdQCFMTXfsrotA59/wxFpiDZ02LXyuxta0
b+Gz08INPbmBzXEhJxsLYLxSkcvX+Lyxr1CdNgQnF3m/EbMwx5NB656XcFZmWCXU
q6eJKgGFdv+GMknm+kNcozlRGaHvkYXclVinrm32IQ6v1cu/HCNhgDgwf+br3Jn7
RzOsFrCOo0DEg6rK/9XV8asI4Q6HbG+ZI21wQBQfEevR94OCx2FChVHJjiopIoFI
W+cOe/11wLhQOZeVrg3BXaPgxUD3lEqgw8LkEan06CuORukUjmNgBk+kzZ3mnCIZ
MXgkPb/kn5H22sEawGu59PPVSuyrbdhYZ+ryirJV1n8vWCX/7FKtTz5mczKLM79o
QufkCFK6qIOPiLSWxxqjzhrzszpPihLH6Xp06N/kDfvk8+ayqc9ZPJm9NWiXh/mc
3oMUvzSx3TAKn0yH1ItjVAReao+xdHJDxcxJFjaStV0QCZe8nO/vG8vAkrskHgti
k9b1IDv4K0NHfDihYZG/oxe+8Nj6/Ql2qZ+l75skYWBE6lv8CU7HaYGdGgww4U6R
oWfhP3nvlAWsK+mEY11xSGyxlcs6rM/Ia1j0xLAaBQ7M18S9m+0P+Z5qUsSwA5cb
Q8YG4xTUeaqTJj24QGn7bltL7rRgsJqGijTs5WH1HjxznuIdYyoBTAHpP446Cbdp
BxLxMjFA/fLN4HjoHgpQu2PQDnZjIhHVKSwUSKSNb6Xsi+o04iRSXKty8GujFmGH
zmBScP107HhJdLTXKdATB2YdZl4Hst/vbgCSSMQ/9D+FW+C4vyVfj2b1+UQr3jKi
y0s9dpH2MBd79jPDhubi987ED78nW1MxyvwQ8cYRljKA1upTtgB6Xa/fIWElcyCE
85jcFaQG9t9KBLtPOf6vAxeDGxsWxeUBoMkXKeLcmz4aePwGnFisHDWym98fSQB9
A35/B7QOS5pqc454Wi1bj0o//cVId/JyD/wxm7gnCkHrpxcrz3iczMoyNV5o1T7T
oqE8XtlE3aqXBUA+c6jG57sa5ouaZb+YEai1yCunQuavIGiZpqHemmUjJLjvltck
A5XRGaclL7GW4XVK/DpK9f7GUHRQiVg+qKJTcwkLLZUf2c94S3rXogdwSlFRo+9D
ycDeKy16XWmi1hcMmYbIRTZZRD1XN6p8rP5VMFxKb5vVY1cimou5+u67vIWbahCG
XH43TSnsbRcI3JP6aTVpyl+lNvx2mtoOx/kLb5epjy73+o+lShi5qu9YYstU0RIi
kywmsOyvUuYNNA3R0GCK251K7mxhcKAjQwip7xi1Ae8fiPoGAOrofgQBoqe6+4j2
BzQ/RjHz/BQV+sa/qazgbxnaB80wid5fFekzY6GUDz3mMTgAHf2mPMBvru02yW3Q
cib/LvVjgBQs5OvDzORCtnJ6/zDXTbq/eWRuclSJsIziAIX+JAOaHzvkDQyx3yxi
KJI4LHBonsp8vukARcxl3vx9rVfpPmVnCR5ohDeLQ2dWFmz/2KnNIUZ7JRLmV4m0
15qdRFal9LLeIBTphoEun0FG+fG4pY+n+NXIzB6/pVfKWxb5gPifPS47msF+7GhF
AXEtZXMjmpVWVbzpXwmX2DGf6I64v8v/GdHulVqxl8wKZpMjK52y5lui2Ac4+o6c
9X/x33E5ZpbBmd3FhgZcHDCP9RbpJwiLbqZeJAmnNtHrswRINvEOXFNIxQBEzPBD
X0pNZl7syOY6NTS9+sm7tfFbG+FORIxLG+3Qoy+xea3ymQWy+rvXUTmbZfu3IYsY
RKGWu3Wvoiq6XlC0NTIArfTXTdM/vxAj0elbKqtNwgG5l/3ItBFwoxfLq6cuzjOr
14M2zB6kwAPoWgK3cQMY5qdl+w+kweqgGT7atZB/dLjERtRoXRdiSsrT+HtENKXu
19bLNFVKGd6tugqaZkDtwTLLaDYrnr8B9lw7BxVeAqppOb84eAVqlSIH0g/YBbty
uKczpW6xYJnwE7Kl5H5wxjK64tE0mKESVVTK7s13PA9jDnhZzEDBz6MkciXtBCU9
Mbp6Xwo9YNIr2S3QerGuRU66JC8Tutnl0Y9t0YuYy2lAlkvyWq9muEYzVFyc1LbJ
aje913N6OzJXFkI7OIkmi1kKHAkryzhl6iapAq9U6e6ZpY2pp46q+t4snZZuG/mD
hCIGV/WCY+Kz15eVlqOOQgMIpBLVq0zMuWuLraniMiLCSXwfZOv3gSlFqhUEVweX
wwnUnZNZ9XF7RzZgMc97XCBuHR6Nlb/X5ShI2Kx6/ZRsKrgqH+SWUmK5cfsvud1h
IAfhiPzFiOqzlyfPZJYLkqtInrN9lQ9z1izMTSf/A36l+jZntgfCFTOwSpOnKdnB
lr2mkjWnc9GV5NKKexhI96+d3bhtyDnhUUimJSLLWsCQBi4z45h5Uirht1A39qW3
pF0E0kdaOpBufQrFr02Bo7s0jIlFxOvA1fQQLyODy0AbT4XT+5CNowM4SiXhLiGZ
oghEUZ6ffg0gmxccVH3eDiVGXvdj4aZq2i+7sUrjSproayWpaloZzDVUTceiCpOT
/oJcheA1mty8AS5yYWnz83uAeR21T7IDFp+W6PBwAJMYGHAyZNjx6XX4+BvcCvTf
nQoGqzL5Orsrz7x/ucSY4zp3Ekp9u8ca3fkhNP53vcEGJI1+m/lI632vbczz1uSL
B/EQAUwHRclBH1gWPpYBWhBwPQgs08bYv6L06fRt6+k0/WXY5sLMQBL7cQGMP75m
98BmsaJZIQJDKAWkbPRox24yJVp6WzzXn6Qh4LsGXZDJMoz+8XMqXjSm08ZIpkeH
YKaDshbpNLiznmsmAV36n1JjJxhpOD/zCYBlV14avh6xx0wCUPX90yyCqqtcaI1O
GRiv06PPIjcYPLfSM86fNTszHRtSrh91/kZDi6WhRCeEOeZbHsHCWGZV11UZE7oI
/iPojiwwmfEdMUaEIapRhvP9FhCJURXQJN9ZDO8P66G+oRsP2eXLLflzEgHNBDGA
XSk1hEuYHc/GhVO2fAkmrXCpAqlvMvPvA2m1iLGMa0eZgwGadS2dhC2BNxqJBLgT
wTC2a3o3OCdU5sUoBuQ5PUlLGeHGuz7pIPrPNLqIMdpvkOh0Unqem8fNevBP2E+e
UL1VG75bifZIHtFTO+WyBmE1OjiChlRqKby45rtSF5y22PEPnI6ShsaZ3vKQsPgT
/lWEsrMV+iyTKG/m/ZXk21HvjI/gvZZcAiu/v9z1P/5W/Q7OVtn20STtohzA6hmc
O0qrVskD2FgucPRnZEu2EXRQ8wHcSkaxkDIxpgZkNS2cnN0ki9AMpar1svho40bS
qp4v1O0TqI85gqlRHaWbQl1z0MXIfIXbH8Tx8Y7l57wR2YJq1zIz8zEipTRnb32q
LSp0jDG8OhHz72lnuD067gFkrG3jYv5aVXBUVrFbhgLxLMmXQ/N4+3P4KCE52djs
VvdTBQDVnkprE0OcnHZjz+soeC+4eE4TuCXKm8fL9vLQZZ7ut3dXKR9WntIf9Z8R
WVXNodjb5Z6w2lHrRrVWx5LHxHVkOjQ6jYVMywJJTSgXt+B9WmDbrNxUUrGpVnFL
OiIUhxZO0hkvAxpRl/1SP6s/NY48HO3syQYQlRo2tQ6B4025rWvFcxOwwZe3B5uI
DHni10lBml0Z6ckS4SibXxws7xR700Y7wuegFYDgjCCYomZPLLPgInYO3qeOT+/c
LkZAe9LPVL2WdOpBy2/EsF5d2aJLcRCDfs9RjTnj2WfaPrV9eN8/aAu0oTJeBwkx
R7+0pQCFttUsL5mdEJdEvPWsph5nWtIHl/JWZGiozDSD+tXV7N8+dRODsrnzmC37
jokpqsXoDXDEL2rDBd4ApwJkS4KMcVRdK17Yk8suZ1680+WjydmPaobh4wNsHaHm
hb0CHzEZ1QbrkgcjoR39sILTE/kP0BMh63WKTe/xKp6gxfgE7JqzP97rt2z3pzSN
uxJ8asfg5v/mgdqz6aqOpLMnB7kT45zmH43+sL/Yc3aq8OCWELvQ7on0pAVIhmVx
tA5hKr9fqBkHPM/aZlACaWjF/SFsjM4aSPYIAeZApl68CelBqCFJJ5xwjk+H6ZHz
jXIBW7PKrIp3i6+ZKrOt56pxKnyWbvNhVxtcmhwYWou2zXUMetd98ehfgMIy8Q1b
9nm1hVSuyd6HZLwNLjbgZ9e0yljPi7DzKv8TRYUMnmvr2lNHhdKojKYoZt+9Oxtt
k2yAuWMuVvatdU0aRyqKG7bwnXI2kWvynpDQBNPcVSi0ZACd2L4wcyUcK90Xhbtj
ISa/PWVGIbhBtoyEr3rgEmAECcKECUDNBeMS9C8r50pL9lcDe/9oPw8hC1SBjoz4
ppg0z3HgaYyuBjTsdbXCt4YUTQDCIojAEzDye3pcGWYmTy2q+/jxxrBLS7ygUniH
nnbc7V3Zxy+acqxmYM+EkDV1awfaHEC42lTBPTndadMYrsTUoabCXhSuFpkpCtS3
60P6V75SO3J1aECHEJTyXyu9sS092Jqdg18Kyi9jTdCJFlqhEEfzt6/IH/oqFeAj
aQ9CEiyzWUVg6Z3TAMhwpiyjwcwaL+5Hcxd4uSffMx8eJ8e94MDIJf0jVMixTSvX
v73ej3keUq9LlQSOv9cZNiX3pPi2vpU7JYoViKIdOVtkdeq9ArEaZlVOY2rYKDvZ
fj3Jag/S7HCCA9S127ZQ6pUfML1sRxZ/RWrnLjjPQMdNLO3ZfXiXw06wnjMNBUJf
o5I1ii9k1yquLQUNQZt8QPLQQ21IqyyK6pXBje4GMk1QyNKXzVGNc7KJEQRyp0X/
AaYHt2OqHyvm7ahE/2NIFGkz12JYQUrk0V5D0VJYd4BLmUrtZtTf6h9VavkRFDwi
9FTEgOel4RiP6VAjqKbaSjamKuYvDSw3/0Gtu7fwHCOOC2VA6lvIruypLH3uw8LU
Ap9BAEAGEGX5my5JCMyujkq7zySQM2Sov/nmrOd/ybXufBQmrKmakdb1x6TIcbF1
0aAh77KUbQ39T0w48Voneau0xidkeQxGaCGPzLoN5rW9M25S0c0xmLxyyy9NgEma
wd4FQyWTxlulQuruCrcQcPYJZGRI2znF+GpskoW3QWsQWR+dMEfTttZcc4JqmZNE
FLY7T1eAT3PSjlrsGwa9/XDwABiIZERfkQ5BW5p0mGY6z7kPmEzTMAlRsrkqvN0U
H/W9WLMKwFCTS1N70sZONQMhyxx6OJjAwd0Tubz7L53zHX+s2yrUcSD9jBfAIwMg
r3UG4EoqthzA2BU5eqEKg2NxeDI27bgix0eB6RHf/NGjbR6eYKtEs1YaiUXfMnQr
GQVc3B1QYMq4/TCW1T/5o4gKYI/WHMELIDVfUnWikF8kyA0Nndiv2CW412fc30U5
vJTz+7DjIMj3RjE7IhufnCWRr8GJDj/DT7IyXTnlJyHSTKb26lP/wTO4XAAYkp6x
ba07RSjPLJIRU/qoY7yYv5BtPzi7CTbzfn3AJ/gz6vCmaX+r0caF9RrsScyPXdeZ
OWqVhK7J16g/TaW5hByFLESk4Ffs0uaLh0R0SE6+dUQmSTFL9VYYJ8t0tyIYzqfn
wZufpTrFjl/TPTfJK9r1A/f9/KokX8cd4S68veL83hF0qXtfmJc53i3pvMdlQd7N
gc03eJNakwm6a/+2F4gPQtYgCqtkQ8zbLfTnzi+DrqAr10i4nM/WoyS0It2IkP1L
oCskDwUdo5Kttt/qnOiT9zddXwV9dN3UKT3WcpCQ3BRFrYXnQru2Sdj/JT1WQWjG
hf794HYn8iXAdOndy0rOU8a0+djreUfUVS1V7lNMuc3SKKy5laPwKy8Kz6B8UxVb
nf4fre77bPXZTaGBRaGSIGfbrUXKdvDEeyssn4F/mD9EH9osT7MebtI6wbz8fubI
LOdgEA/XgmZan1vWEQF9wda+RdDZYetXkKH89qjUKTjniJHGALWWQAUIoH88XkXk
aUjOlBM34E8HvDMLUcdHvlHKHuCof36u7nwQwjMBR3J8ztvRFzhWURCxZVL7PYWW
a7AWUfaw93P3RK44ukMbG8Idi+j42FhJcs6b6r6ORWnWZ1wSd7wmDheMQ0dB/dVS
vJjUst+LitRhi6/Vjb8Af7RzO0aW/NmG3AKN/NcYt20/BZHP+QSbKUTLPFL6H8NF
5mGEdvytupZOVlKpBuE6FdPB4jCfOdNNJTCvUTvwjpXJFcPrIjtwyRI1VufttpFf
hcJ3NysgYTUBeg5TdlvZZkxP6duUSV2d2PSOKXCpRoquJBmnFkogbhmVPDBRn/dh
ULqOTTUtZRSMlQxdEizeKQOrBE/DbauGjeUmo8QYwXmzZXBQ7NZ5SrzPEOXdjgnU
ydgZv8v9uAnzTQloGcOZrfWHTmdTVuLYfhCIkEPBfEVDWJeupc1W56iINiLjcQmv
QR5sp/tIN9YvNeredrSvQf4Q72SyqgGpUMFwNPhjcfslfpDNZzilF57oVaZniY8X
Rvw13PRK9cG/dfTpdsaOOGEaurSEzgb5f2ULhN4STVI+8iICZL8PMVWW8j4+m4r1
HiR0XeiP3WW6q2326Jz1wzxDhWhfsjSvJFW2L/2nIzvdRZibKjf1jVSpcVCqSl1W
hTrmIS16CWTl68Q9mMX1SaAXYR2wcPSoOtTz8uk2PhzY1OF7SCfJwFoofKD4sPBv
gmbd8eXbfzryQ2t8hbOPPuCkJZnBcDO8hDv/i5JO+y/igRwhNhBG82IVp65tjtEd
Z/94fIu9Qe1V3z/hGmUlds66NhAJrCGSuaQdtruWJXyhdpUHMbDWSNaGUUSEuEk7
CqyKfV3jaOMVsgQ/a2kmDdsUDKEwTMRRqY0CZTSSCg3jtLLCX946gRDveJSpy7NJ
YHQHJaJXLHTNRNAMhcJUk92CKiGMgA+IPjuZaGdLjotLjHv44koMS50YY/6KbZ6s
zv89Hd/nm986mSt0IFth/Gudl9D7eJS16mYZ9CP/qkhRXGuux7EN3uLyVOA/aY+C
c5Y1e/0+IDKr+afBhtTKX37qMLB52cPPBYL3JCQo2An/6xC1XbM9gkhDa/2gMWbn
xx5E/8Z3liB7nxu6QBJr6vDATacHUf1R+RcMAeVDldJ/nfwyi7qFCemNCTkZcK45
CY9AUApln2ke+JZ5+azXECVbXR77/1qvDJZ4ewSadONHx1JbRXFsv810guVPp1uw
MDc3MvkXgA3pVt6N/sb0ZRPtaYcPrzcS5q3Ft9R5CpEF8H0oEA8UNuTJMFdxEINt
d02geTxmu0wjQVrl0eQJOgdYMM48NwhpmO4sprHsAIAAjPo7e7kvrt/fS8F+09jL
JU/OU8HCpZVe2uDIFV6Hf/BQRKbc4IKKSFqEWTdVJrX126kKCNQL5aBgj7iG46xZ
UtzOYuRlPkddRkTYkl60vMIz6B2wyVD8QgVwyEOsIbMF1Hc+qPAZLcjc0PTmGiZo
B5pGJ8PhXhBhB1Qs15kY27PJmb94bgf9gp+DxtlY0GeFr3T0ReeA3gM1QfuVj1AR
1Lo62fmrusLga5MMPkXeRUlAo98lZ2DmStKTkywePqTGElg9i7WwM6zgxaTtJbqK
2g60YXAkRv5R5SCzHTAqhF01ZtZpDXTngzC3STnJYpxUyUnW2I7MFUpS2zRb48AU
VBZL9HrlpYQQ9spC7YVb5jhAH6+vHZBlYocv7w+9t784uEQiMKMc9AGcKjQdLEZG
MmgSalCM9X7ljaMm+uDIMNHkc3j1eAJHIXkxsoPWGDkw+nRpihWnIgUosGSsn/tF
6rBdNxotJBUrbPWNZj//AYfGOY3Onvf7TavZzLSCqOurY09pF86lZbISJTLJ/03V
+SO1yxkuipl9a2tlLL7k/OGrAKdutD/Kgg3ruMWuS1w0w9pZgAptCrOKYGXqtq3k
xDUtyBGX74PraTHX+qa/wkbG31UYMWu6RKMP1eYWeJmeT1eYPxzvjDqJoPkW820/
IG63DJI8uPNzi7+eJm54YCqjRu02m4EPMdYao5ARH5uLcB0PNKcUodBQGFMQRlu5
860TDyPxi7I+aWSq89MF8yK4T0/qBni7GOwkAv9CJub7DK4/ORKzwfsEsRktfkuc
7T/tv6t0WsidlejpMYbM5bRHAIWDO9egt6Um34Hag5tM+gmhdujNZ5eSuN/LqnRq
eNRYr2kKEwZJchpaWHlsJe9MbCP7hcpHxgT9ZSLWZal44ThswgpizdUj4z+rlbiN
5beEMlD9PqIA0MI/wO5t75J89XnfxypsAlFDhIxerYe6hYHHx7lU0Cs+Sznba8Mi
46smyA0cxQPZNCd6jGrkXfihwl+lAy35pUhu957xsrZlsb5E4/SZCbFkHvfGdMDJ
pyJ6gNMe8BmOKKuQlgUAWSLD+bCE2Lv+LtQ3SnKazewDrmlWPCO2v4uKTha8kdwh
hnFpROOO1Rd3MPYeJPSV/dVNQZu0Pv3vfcunUVYLpW/wrDpGHeU2QQ/IgMUFUa+Z
wfuGiUttgErJpULlksZa3KOpLcpQWOv4/+xxM40EInFGBc2DnAoQJ9+ZcyxefOSw
SR3+9M/EWy/fucW/8noXHK4tBnyuYd0mU8gHaOMbHAcs29NiWO//PNtBtrtOE5D6
V8zl9yORjpJw4nMPlNfMOeWhSXzPshFu/8SN7FxYEP4EWxO+RCfT2aIEEAgQUOoY
drqGkqzzJhmWzFC/a3EI56ZDXo3+CQiJYwAVm4a23RQxoSlIfn5nq1uCDnfAuDGe
CcoalLwfe/T5Ckeu4EQl34YYCsXCeOaTyogV9aUMp6LcVFBer94tV/R/XrPSDZmn
TL8e+++qts896XLuHxJbVNwetYhcnUy/0QcjiTBkf1apRWa3hKTFVZIVcRc3W9rt
nVo2CjOaDzfeOL+8P7PnAs7IeJmq8dQ9Fo50Mtmw/2/XsXUqN07jSnwSVp5pXJN4
mMAK7UpFqAGV/EAw1XQVDt8rDmTnvXQAwfZy0cjLb0FWRovLvRjHy36Kan9+pEtc
aJ3ldj59J3oFyf+DUXWR2s7//Ra1ZtJdZtMYGIqOHCF62tDv9fI+ssMHjTTzajB9
VQfjptUQKVNSPnLQ65GUANjweEiOZtgZiHB9Yc/5oHHiKCr10pEftmslO6tKX33F
G2c6pVNyhWU6YOyxTVQBDmZRmVx8KyhS2G+ZyYedv+NELjCuV/jRqtuOSLHv7sa2
Nl7v1DMbDJS68sAt/ITwB0dXVFk/SOY9+2a6Sal6ruVYEImoARIj+fcqocAlMbYi
5zu6MSXzQn/99wJXyNA5mqni5JAP7odevprWKHgerqOAr4QIKkyUIcdpEeZ5h118
AeWp+qFKc3GjmcQ1kaJKlMQ3TfPk6BhxQFrl53FOhtKvFeBmed9j/EjlX1syOHoi
uaI2Li/x0jLCznw63afm1sFkN8rOVEs3axz+oTiERqe2MRCTv4bC/fHFjfmZFiyV
9+5mUxTF1+pk5yaod+OlRjEuZxjxDmcL2pNzo2cthaCCnGivzoWRSW9uByHz3bNY
7i6BnVhHmsz4+5C5KrMYREyZYK7HRmioAl1SOHIzSlKgSdk1s+bK8yhpcbc0jlZY
SfQYZLXkbVC2wFio2/YC3GtoeV1xd6ITvaC2v2BhXqsPhhgtaFUOHrIbt5sfFndj
mmh625j4jOk+89ybltryfGvgPxaSRY954eQKJAwQOQHhvRhOaZQDsBseymuxFMQA
1r6rrm2+j4JywueTq3hRqX+BJl1Um2cipLYfPNip4+sFu5YBW4eDDBjIxnGJun7Z
oXqsBaWq1MF374Et64KqCF5b1aWiWLZHOfIfqgXoRBAjLNnQJmNxCuf9d68IbfG8
Sjs3RwzpJ1X/Wcn+WjadFNXjvQf0yM6EECs+AI5Z7WoZydy9ESgCxzSXwU8IzAzq
A2dR7af6Ju2/f8CfuzdgLsjIq2DTss/Tua+yd2/DmIITP6/YvlWOpDuDaCGpuwJX
f9wWqOYB+52fHr45Xt2tuU9r3wFiyCGRPaPXW98UQDedlpgYHQ3T2BZzZ0EBewaa
8PxDZo9/Vj8SU5lMogCXUliRwFVnbPf5Ow6VXH6RZIr+cXv+YuRSDB6JXarZMgqw
dkJidpV1sTx8TVUROjZF/gvPdUt8K+wMzNS6zm5XLks026M6V+j0f0eFsfv7qCk+
kelVrHJeptIJjMpTD+oh8/sbH9zPZgpG6++8YVnpfl86ppFybY8aDjO3PU5OYQ8O
NAET3+ZJaL7ZB4AgO5mVzHOPyrGUGOWc9R5fLoXinfQjsxE03P6AvovoWlbbeCCv
pSmSDPXDuT6hwDIaQ7LBSp8z9K3XHhC1UCH3/eXZdQQo/XDlmuOp64fq2F8yxenj
3qOe2s6toO2jceQIMFQnqTgkmx6tDGKVL+wHzxGRXnyD424c0nCVOx84b8sGG3QV
bEYRvoNzAXBANkKxXWNaICBZJr16Vx+iOzVSAWxZ+Po6xlWE4sgx5TvFWJndILAA
tEsnb4eKbuZG5gePgmJG7DlvX+ipsRtxStiOOeQLvJtK/AxI5dW2vMtF1vVgYZQO
l57bRMeQNefMPalzt8V23TbAFnKab+fIvuCIirwk+9TcChtXqAhUy1t+J2m/+tnl
lG4xkO8u9pv4yb/W2btocpFkn0pRXVp1CCoWifUi1u/ZZlykA40upWH+hLR9BCtS
Pz4PH07FvvRdkGttn09i1fDnzZLHEtdrZirUijoWA8gxPpG9HOZF19Cbdc8XBaMT
KDmRdMjpM2AYlv0dNT7C9pHrNwWtzQ//3WXuAKs3Gub7sNfY6Z/q/xbnVtdiz6TN
nzvf6+FVTWvJcSPhAcK4MyDbKNEPBWnhEOnLVlDBnyIS8dkSGI1RWhbfq4wA8uQ7
mqK+xNd3eNRy3bzF4xARWooS0/1jUygJX1V3T1bqfW5cCnTYkcPrCInBv0uVL9Yw
YRqti64uKU9Jma5tWTBLBftijWW6PIwVKvwBX4UszgpmBqCIFk4tsXzdz/FzsueA
quilJgoAPtpJlWq4zYZ2lcJ0YmcHtuklgWoDeILqb03/iKx/xmBfkAV825YtWjAU
TamTqGDzr3gYdWRPMyW94GWUX1B+89P28O7Sk+VzepjVbXslpvLfmKWMCD6mQd86
QL82li40Q8p2BzkTw7wLCynRFDukPDK74VjigqeaAELItj1XZemBGeQqEYxRSKl1
JLL5NGyNEv1LA1TbjkP66C0uyf4ady8wFcQRm3sN4z31H0z9esDdkM9/RgpjFnWZ
YRftw8PT0U4HWG9Vcx4Yl/zAke4gcv2NEmRQ5Ue9BD30dpYkQ7kOtpz3d0MI4t9k
0F6nf/usFhW+wvs1pvOxoEO7KhOPPr3DvExGfJeTXSqkGWejhYz8hs4EEMFN7RPC
L2H0PZu31B74atOY5y9h/rhoEeB09Q/OgXGdDILScMwtAzpM0xFB/Z0VP6aY4jEF
4j7B4OhwKHaK9T7LoZ51bssUiIfPLLMwChtCLqjkIBlrRpoyRT9vaQJ93PsX3Bsy
rNP2dkP7v5TD0Q6hWpMuFci9KbZgRZax35ITR062FFXFFRcA5o3g5GjDXC/+/Sfo
zz4rs2JJeLZrbxkGQHopehOwgicb8VD6Fh45mVNIEwrSdUP1KmSFjSB8Bq6L2ZL/
k8BF5JKSxpy+2SmWdCNqNRnMx0kcuPVXhTCxyngIbi7YX8ZUxrFDuey8XbMIB7wR
eFcBf1Hn+omyh6+D/rnVjz2LO7l+Qrr1qE7scXafX56Txz/FSmZvUzV57Uh+OesY
YDhpszFuqMATJu8CDUKBTfNTpLkXMBamv/xDv2/1IShfAh/8n4m0saVt1MiIMyKN
H0l11xETU6bbHuEOMK69BYbzDEQR55LyRIeu9aogtWNl+NVhqcNHsc2XCU1QQ8Te
4ByiDhSsU9nq5VF5efFUivGUytJg8vmYU+c9qapGgvy+x4WDAL6gqKW7LqxFe6gN
hyNOAfBuvDTlJs/9eGfaymqdDUpt2KrtapunHTl1hWfun32PsSlUcCE0G3Yta/7b
c8QGPlAnFw/x8KBwmmMMHDTLwz/UhTH1ItnKrlDt80rssi4GqQn0MAVsHL2y1kwI
+4Uidt2sMYrrqXQYKMDc0v2OOHKqobvPFljOxFmyTYQ6O8drGXEeDabhR44OZHpJ
aigplF+CuJHxQDlFBkYqbg63pLY7vf5J8EgGeSLZEMO7ZYvYH3/eJ4Tu09HQdDFx
yPc50Q3qAJ2/h4L+iQClPdLDPqVk3/NeiOLDU2/TVUGY4VC8ibQTfTa0hwgNWi8o
q2xev78dUtHuSmqXM2GA1nfLIZ2LUkaD/u67tmdSMe3LjbHRXLY72PV9r1mXyD4G
rVDQ99Jo3mjzhVR3fLuUDUpFBkuCKyTo1koyURevEJKd8cVV1fd1ytgr94D8xQMt
mutJCGErT9q1HOwgOS7F1En1ExZAiAtF6NFW+ZRKmdVhJLnGrPp3Vxp2qbbIfPMb
BD0v6+oiwGFfFB8OupTz/iHfkPZI01b8BH6B5JeA3sD3GHRjBnEkFeMHkBLNQoXE
RbHRIaXnGCQGJLPyGnsFmlOxlw4HN0dYI0G8pEEGaraSwQAfBA0bHRvwccQmFTG+
aduWq6gqbQlf/iklojl/LIr+zh3dyNqxTIutmgEzOS5UFFb0H/ggomi8HCVkWKHm
jOV/fDR3dRLuKfwY1SJPD+oVVfnu5eIL24VGSlDguwh9LNIYp4lkhmYAmwND0pBP
z9MV5FcIPrM94k9qrO0GYSYQPNM712V2MIzWq7+H01+suW+xXrixie6Pm7WpAa4y
ccC1faF3iZgpGFrdkREoZGHLIvhDRVSeEZlpWiKrZzE4CB6W9F9OqaK7uE9aLR4T
E5r0vkOh+bRmcxHc+JpRn53KCZFQqr/1gJhLxTDd+YE3iSImj/1QTJiBuT2d9Yn+
8SMPPXWtiRzDQWPVzGc0YTc83bpmUQwEXvkmkOxf5iCbJYnv1ZCwreI6V6Xx7uEE
aWeHIYYYMtkZtHfOsD4L2djhggEPqqd6qHMkCh3duJHjqRnYOxGZ92P101pkdpq5
QhECsFbzADxnoSlgP59c+he/qHZfHHQluPhX1uxodln4Stm/NWOA3TuonhUlXYRG
wkmeR7mJw9wU0RrdLBCbOHtWJ4Imjnwa5Mw1Vl1r4JuO20ZplAIU544/5MJ4YzwF
AywjT7dJFhSEnug/8vfefZ+6Bkkb+zA7DbicgDHaLzgOxAH3s6cemQkfOCK6PFnk
k8VGSOyGOpxN9zpMHKkC37RHdOGKQG2zSBezgHhDQVyPeLCKfXQtW9yRVjRDrs5+
yC0AwOyq5Y8rMTf3fzXxxonJ55qB6ryb32aJsHAQ/wjOQVydsFbwIRuS9IEldXqH
wzh/mSoSlg1tvOevYVa5B3lVIzwEUE9A8BG7YibRqEH8Y0y9jl9lWERGsZ02aivO
4wtqmDEO3ulye966y5zJbNUvfKIWrwDNQ/hAjRwnX8s8loYcW9irgWXI5lz6j6WT
yXhBnMk9jDFBJP7PT7xvh6YRoP69puKsWl0Q7Uj70iAm9t2HutRjLCyaTyw+hU11
zSuqsKJ6rpQaZV1XwxvkYXvrix5Xu0vP2rSKw/JCpIfwRjeAaYqnqdNC3SuITz88
OlatLmO8uj7OuSTB09p4X6jibiQB/NinLPWhyxx4unDQ8Ki7aL77KnZM3rGrcSbe
RmmNPRXhaF96og/x5wBMidszfTZtOm3ZouiABefLA4uNyGUBPfSLvA2rPh2JaQGF
4wqADZgVSZ6L623rrB5AhyEOReXgE1HskQhZHeB6NG1EJHrTCqHgS6D4H2sSD0JN
ieGP9lnohnfvqug4tXh1WMCAY1VK/gg+gLZHjYhzdlnE0AsF+p2MxW9YQkWKURQA
fMsc+npZpPij+6xaJe7/CFWupFMIkbP0LlRXwj3mOl19mq+bD7ht243msH0MwVs9
6D30wx8Womb34Fu++BDTuOk52QW7ycJXJ72Zq/x9l41tMUd6m6/dz1RTQW8uCudr
eozQm/FKDaFzLKVz38ZQ640Pyne2alEGbpE/HWeLWMParWBp1WZlDKnZQVvFKtpz
c3GpFxvDIcwnOipuM7Lnq/YXLdYlqYfjAVnlBT/S+C80ntTv8SjOmZbyXyS3TyKx
bqMI/qebUqRNnNiebvSwG+zpGxWLTsR13lrgtrOFlyqiqhCcyXlFUIw7sCaixvpw
XZPunaepvVmh0d3pjhI4Cc8jUojwfnVmDI4gYVYMdy7vPdATJ0Uxjymlzwl8RQOc
II36EDBphBVcwc2jZXUBuj5kkfOi5CoTEsC9kURuf60LfmBFQxa4BFotS3WKOupd
YeAglrwsNOolhsg6LmjGCogFS2GEp0j1jjZ+nwfSEilaq/xpYLyY31s505v3wffc
aEAMHg4J9j/4mlJqIW7mDX+SkpxQyaZnX10i1WrSGCErbw1a5+iB/VZnPC8vTTPW
hffJmN6RhXNghWwqY39uDJd26W6Nb9itTCmKVHQhNeGPdyQdQb+4C/HanNbN7ia7
TV1itH7HYPdaGK0VxQMgsvuA5lgsgY5eNhvF3me+JY+qr55wrm2kvjeVIC5BaP11
waC6uVAmyyNsMRBbD2slYM32JT5r5KRr2z+XiSXWnt/Xrz6thnfB5KuqEg0L/KMY
sr3i39/69McfMts7rSn0zVA1BaXzxBfuDmM8Utip51ytVW+ZE/YB48K7l/GT2+R4
44OijVIjXkklG26ww4mU6RbROoDdXk8Eosw77CXuR10tH1WhxsHUpC2oaX02vcXQ
LLetl+KCXdPD4OmYRnUNAxSKhMse5vsYZ/VqAa+tHqX2Ng43lRUNX8tMF0jRK/Oj
qkkuLkdIuN1bsF1z7hq2VptiDlh1qG7S37rG0iXYrnZoLAG/EtAbXTRyzZNegSKv
Vgjwhdlblst15UXEorQAZs6lkCl1bxezNJQJV1vOd/7Oe7GgVI5QlORdOw/PLTF9
sqSULuPCQtaeVLQRoP6ytYVohWsVGdO59uaMCFNvWChoaDp087Ici8CGBO9Wevua
RAqJ1QzUFTLen9OP8UY/qW0TcoLyLPCPTn+CEhmDfBfmnDq2hKvYfZmitmS3NnL6
gr7tMMs7JgxMmDzYCbxl/cFAG5o1ZjDBpVF7c7Rb9YNzw9oJwy+XP9UmMIjwVz9M
wN9y4Z5v1CEPHCFG1rr67JmiOhUgkmQsCA0zaoPbVKu67jYC21fcdH+wRqpAHqY5
xsgdSHB4KAnnXNtU91uVzJ0hKnvluy5B1PWG4YNt3DfCGPGWYvRzniKApTTI3MQk
iClnt8JIejZtDAbPlqYCMQN0G9imal5LSttGxDO2NK3nT2A2j/QYCLR8Df9j+FK7
3vzkBVCaQ/IKKYwYnIlO8FzG+uZZHoFu0ULLoxZxkl/vVj+nB6xeK0mPqqt8vFC6
y3CODtWtmXmdfPup7rYtGgXwUPPLci6QfuTx+H9IMzVu6CqOkpLZyWos98VcA+4u
+8MIwNNM5fTG4t3FUldy7OPLKpQjL/ZIacF+criYo/+a5Vjz/U8sywtI7AOHd/kL
ybNL0f3PnS2IWG4TvX18VopajvqNoSlQdclP6YLjAdSZQlY4euiW6DdOLak1pJVv
Xftv6xoq42pQ9s9rMtZESXZibqUoPxNIgCsiMy/3pAHokH14AhIGew7jcroHl67e
gCJhPV8T0ycqVhCKKcIR6nxGY+4w8XLkx4YS5JbFIgPmwyPvOLD1CuENyO6SJVYr
Ok5wDqvjx1zUQQVg/JSV4sGhSDWe4GUgfeDt5GvIlsBJF9+FpnDvesFVl+q+rVt7
sRau2Sx2wh9AafjGyBSgkCjZo2uTy+obUR7wJ4vAuURGCU6J9zqGSOqcRez8uWvx
9WQJlXtRTqW956A5MjQBFmeSXoaHdNoT9gHqu8J3gsWz/N9TOKgWYKG69sdj04o1
GsDRyRgoq73gtNnW99V2WtV6y/7hCGHww5+b+9ZeUq/qMM/NK50KKRc88mTEO1IH
Yfsa81j+a7YeEvvwYZQVyw8gNbX/lAEJfBZO0m4pVQg79iSzUOK7wsPbzogbjFbk
CFD7DDlCl1IHbcYx15Obux2KHUqbXf+JEG/xQ/lS0e+vGjc6rLLzCzkNQTHLJA6I
Q/wb/LT00+untmgN61Ogs4NcqY3Thd2dJXML9Li6FyE6QVF0Zuk9wd09UfdbagmJ
O/UZaWJbGhNxdU/XF64xf07y/JseaYfWEkDKjNfna3pH50hCFAXU5nk7e7oNjZ3T
Ytune2c5Bwrx/wKeGh6ND/YS31a2BHpcr+JFB1k+DGpEzl31+fQTwC45KZlSvnox
knenkzyamXxQmiaYMNKQbDZTSBD44UBPLObacGehEp5t3omvsezS1dZGLDbEYaj4
mcRQixNQzvMr7+pCtKoBCvoZBhMMXWeOftLFtt7pcivX1Xyl1IOCPr4wuA9rOxT4
ZGFJi/ULkZJMoIJcXvUAHoI+XBn427+XnWi2WLMI720CKRDc/54w/lqsfu4ljMeB
4NxVdGBOf2H3LtTTKAuTQSHP1auUbNchg3koDHX6VuQTJQlcjUdpIt9EdBN6ryGG
gZqIBOvVMLa0guIlgvRa5AS/mwrD6jZ9j0h0gQZDTghwcjIK0E7rb41vbP3Rs6p0
SfvHAiGLc6Gi36sch4ziHuSBQ7xcrA1KrptVxH6gOLqW7Tdwqu1/VG75nwpeLT8R
AQmg49pesSKt9pwh/MntVytEBu96rn2e2iWPNCJ1YEmYRrgW9NrwiRzDNGSIkaaJ
1U/DGcaLTwSOVP9ziH2ykYNOqsiwzYhyzAQc7jjC63pv1cGk732Vohzr3OZ2Fm0w
KBqH5tNj+1L06SC8bCDDnagGKXg3mk6AKapGbl4lLmiwiaN+oG9TKmxk/ivG/IAw
WVDdgorZc+5SCpYsEnrp4kz3hD8335f8bk/lkHUd5mStNfbaiRaQxoIQ48O9y+lS
BiS/MOtSRHb9vY78C41W2PULUC4CcYdmdxEqD4XI9pIrSIK7m6LXCcYk+v9yCUTy
RhxJ6epEOOPX8x8ojlMd02gKS51vV1cCVVGcFPI8IUHAlsX61BwBfmTuXWp+T0lD
PF/6R8O+mRjQnIWDzY+zLnxcXUUjLxIS6O1I0cSyFKNoI/a8/BhbnE50/GG7tA5j
fN/2vk6CoDOvyBxQ8a812sargYhwMZmyCyuw4c1VAFz/+w1FqyDdxDX5zezsAvac
rYyG1IZHszrdpvv1GZkOF6lldgilQRiC9vK5svGFiFNhmXMAUGp37veT8HQEU5K9
gcSqo7VqQaoyj8rNj0AYxBzVEMS/QlYoNYl1NFmfyN6dR0PYyxHY9ZNvx9BJ3PIW
91U7QK288LCYib2EIz+JLctXgv4635wlVKcoa/lNqnKRA99jGdvpPbhGPylqI4MU
zc6W/gc04BD1YeLxPnqx5oEiXBRN4zuEo8e+EPgMC61COhuMmow/kiPE9Fk9acuY
zVu4ZKr/8AlzPQKN8UsvM0S5ObfhlNIE+1FMDdsfGujbq6It7pV+Cl84lEumI+wP
aKOPnA+tTMry4udxyjB2WAP7f7M2rJn7VtZhP96U5VKUk5UQatxeNO+C6peZquQD
Vtm8ehAotk1nkLepbBz4zursS56x5f4kKB3ah2K7PrLLI2qgnQCwnCTqMJVxwsFq
mrGQ4J1tzoV2nSKi4IV7n0Y4+zVWMZlykHTMtYJH1vT2XEnHE0VXfU0siMdgICBF
3e8+hkiNQlkp0XGyVOwCh2vePASaezJ6OHeRZGkVMSn4z59QcsC81bYnUULCjl2Z
Wf1mEIdesakGvKqN0ud8644rdBAWdXp+gC5amE727dBDmdX94eh2X0iz1iohmyAr
DV6/KqcEQoHQNciKGl4dZ2GNT1iRPZEVIsbSdHuOMlt7LvJ8Ehts9H4FUfc15qkZ
5bhyWzbQ6bpP6TYF/0LIvTmXk5wG3Yjy6maO/iRLmgyLE/v3OMfUsc5QEQgfdQ/f
rBJGLVX8QXaze0lObzjjJ2vk7hHJnsVe/Kq14ZQRmox6wQPvIXhadWvJl+ioboKG
XHaI6p3cqYI9CgcaBCtBL0romlHJq2VJbp3cTNeNzPmXyzcvVLc8bNl9lejjy6xi
95KjK+gmq+cvRx55lUif975D7igWytqrNZCaPdokxLFwo/cJBBObL0VuwSTA8q29
MaR63ZqyD5jbW5uu/Zqg3EX6kQabxlRoAixhqVNGFvMLC1sEKJt+u1w7NiERbxpH
Z6+VYY3093xpnN3q6RHvACiTjTDTRoUdyfpoT4B+bHbTwApXWyX6r4MYO3dLxWkV
MT/Y5BzjZZ+9FuAOMfduvx4TC6Nzm06vRBY+FhQGNMtfGg/Lqva/bxhdSSE7lsn0
wdY0aE+qZMOMh8ZNhltAB00csaCeWi+c6bZn3aWOJ+lnfKgZTX+FMlUwUEXvXntR
2tSM/160pXKydrEVkrfQnVGKXkuhvYnGRfa0egJgkBtHIENhUF179VxqBPKVOUgT
mjIlPr8JjXR7ClFqBVzthe6y9qrxNYL8633JekStygMkebOXKhk8nWVAoHOcJOgv
k0NUUaTMZInkRXh91y2DQSDWwS80wPdjC902kkX1GiFxazMHxtHj8/gtdWUW16EY
SX5uUITOGQmAW6yz9Lp/x8bBjYneyEhaMY+em24pHa9hxCKVpeqw9sOGuk69FQvk
UOjBprCBwXO+WK32nLSoRWj/pEQX918ZPca5VQhb1y46ufN79ZFqaLqAMMA7lZgo
+O0Fr+ivF2844QvIp0Zov8IgBZcmKbFYq5xH0ukfjBwMqiyZxud8hSVIeqiMt/hl
6xk9lbbFzVegU6HsCP6AV84CTcBstKP1tc3XE4R7CX8bSUkjZtyDIoHps4oGldm6
kg3o2F0QEHd32ldOj42mBUDME6KqxdGJIoaM2+CQpLHnalZd8ZhffTLoIx4C6Md8
jBnD3tudJI8b6UDHJ+Bov7vjQZD99IG3U2NXTllhW2R1O8urtDweFuZs5TYDwKDh
S/MJZ0nxdjLwrYIIEjBoFnMBvfi+n5BCcQ9o+gIp1jv/vGCyZcJ2/Me6baVZyq1Q
vNfPNE5cH3MVtn9BAU/+Q85RF2ylnWtVvTWYuQ+hpuB5DBi2DnJcC3JkeTzCwfFH
GZJes02y5C0Al2wjM0YqKw115DEyPWHkcdmaLoEXzXzCm3mTD2Zp3LGvFnAbw9ch
kbD9bJ6pOUb3JSZftMBeTGyCOaUq1Rt/h9pHAc9DdDjEfEpIruG+IuJvqUTDUqD3
2tlUYXFsUA9nPtVJTePmWwkGvBqFqPCJZ89saHp6AKwDEmua2xcPLZZWI8M84EFI
TcV/y1qDEBNp8OX6YSQAATiwiVPGaxm/nDaz6ZzXRTyomiT+MBhQswstbZSfFLf9
HZp02u9vCpZmeaHeCtyR3ui5RYj0Xbt4I5q+yLYJJoYyo3QtDMsgtq5t8uI5kDye
1mR/O1EPiTBk739NLpIVs65/RX1TLIlXeIh4RCC0n2wNEJgNx2pQURfG9AxGtGKN
d2wykqYicUd53E5ftV6Ev12qyMRcTzMrDrra5+yhZthmr3hXz1X97j/uMlxpioG7
JX740BDXbstzP5GiQ0i5JgOMbFfKGtlS6qwpm4JvSEvIBk8fCkR7M8ATCmadC7hR
DM65I2QQZkuwnYBPHGDMkJj5uxSGxhGHodL+BxxGs+xJ6RO8ifmEIfaCSHV+V8oZ
bMyqKOv55WpKSPBDtbFUUyp+Yao6fpcwMVjhDdKgcyXEmwR5rU7H0HpgPd+sNHII
Wfz8vWLODR2eE1nt8xniLJZ0C//vzm7oNjL4gY5sE7tMYvJPwfcvNEtb7Watl3Ny
5ZYI5MTKPocUwGJ+SdWKLX8/is1UT1uc4+2F0YAia0e88nxdawl4WA9Mc5FxSXc6
69jzT1ELmJvMVFByznuRO2UyPW+S60k8lY+PgNsCEK2yLz/qUpf5YXwevx1ogmO9
XlyUT/TtdhRuBbjjn3CdJuSr9EqS1wwn5bAdPwOUms5SVe17kdDMBBUxb+drGhIM
5/lUxrtc49909MjjRdQ8ABVTWxPqO/IOQxpieYS8DF4hW09PXK4d8WnrGiCQsw8t
oqdfW9kYiwnFChyN3tvcPFsXBxfDgdli/TRPRdAFmhbn5QvJeiIfky24q6WUKq1V
0Pr7taLZNasj0zCd455qizU00dUbA5X8TJcquBnFPPY7mhoi7+fkqA/6xkIkZZ/N
QS7WY5XuiekhmGScit5RIOoy1TlAgpzXTlRZ/GRA6O137oFds7ZZXZNn6hAncOFC
CLrj2CImNhbSXdHucmP3yQ9F1WyFEy4avPVhalX/ZgpRcixdKDyXSWGzpMWOmfRm
36bI29LKLdL8Yv7q01hMgiZpXnHpvK9SwPlN5WJg6CfiwZfa8v+lV9UGrMBEFlUq
VwlXe3McHfHZU4RQnt0ViSOUZiKNdZyG7ebz956JBrZGKY4s3/nbmJV463vEgUE4
8IBPTFkr5nunL9CK4mCG8jISboN3JT0VZPR2Y7XoRWz4uYO+vXYQlpsQelm81DWk
8EljJ/C+6pX5/UxtishZxL54e1qMiY3JIefMjHJCEh/A+jm1u3ibR6jF6JONkVaq
wrPjOvfPBqEZ2u+tbLA0hhpQQiyNf9LI3ZUNLN75k6QYUxVN6C63gsrG+hWv1+eB
SMgDmUtrTSuYkfsUdGGHA+vqbhyUQ6z2Dqnja2Vje8qtZ5Cw/0Xv42kT0jS8dmha
zLddcNFgvE8pXgxAx39GbJ8OfFfdqjzRVv/IBn7CD+LQOltV2KlH2zkAEOEFXN5H
TgdcAtCOlLBUxn3qJmzr8BeBpjJtcO21fgUqqcOL+SicU4cuIaUbyfpCOWK72Rhv
RtHhIc9wZSwlaO0uUvYLO+9pfeuhlYWOiUk7hEWTEWNxvhLUMKmA12SGUYBxZYJf
sfofIx7KZIokvNVyIqHf1vSh4UT10mpIFJCgYGbGCuTA64bCpDbzy0vOiFCBx6UB
YR7NoUFGahQ6bV2CAvYd/VNR7PyqY6I2GZ/SS0xGT3KBgQI4QVFqwX3BYTxLsTsj
ULyvUHefQ1EuQ/ADzPnEuVVXMCSG8RC2u1fQmm1loiqe/DF9x0bebL7EgMfZks4X
UKGKxvk7Aozgp51YD2pSvnCridS2kCCNGXxsrVIuYv/pLfvdU6vkwJzH57Rmix5n
Sb0vUzEm4RMqwJdz5S9PHc9eSN/mXJK/FD0iGwiadOwtmTjwHkyK1SpBk7Zm5oJ4
HNGeF05Ot828ZuGVtUTAfZieIvtu0Za3ZKhmuUfUGm7ATrj9r50qSoqiVh6qSJag
/LqCmBdhILQC6X5x8WeoUhl4//xlHiuP3xtOONgW4Ec9hjwiFppkfUHdhrygLKHa
cL+P2OkYtz+/a3aN1rxAQn1uKKSwBpLC0fIE/R3y1uzDClbS8K6MFoC5bLnTnfyZ
sG0uEpJIfFg8FRHkFpFDtprlArDMcXhJmlPGq5s9aEdD2bshK4SYh2yYlZ4Kbu/j
XceFPRHgoP6yuMHdo3avZGRwwtEacn+iBNfYD+aa4ilO/SkLNgEyWNK54pAn84LJ
CL94imhsvPJfdCGRDe80inOHmyiR8EiXZUaoADEFRIO8DSNlZisnRxiJ3OOETFHU
N5h5Z4gc+5cGaxpymP6/Zy5u185YyQwDgaK7A4Wdg73pzrupGvkYgH7cDCM8ReaQ
U3Q8e1qzPz11Z+OqwNUR4sVxva4oZPmIGALMpozRlcrl1F0LBb2gVB7fnZn2zQHO
X0D0OtdCxaBi/G3j4zBgxkXCGR9jygAKKdCS6Mx2ApMnzgdwwm6H8WQ/0dc0kkb5
iuYqDCs1ZD9a76FWaH77WjuzmqMWt5/SRnBdHE6P2uy+iLzD+2K4bntEQ1hJTVSq
sAcMGE34nIZIuDiSLHDJq/8J5BqUawDKbur/sGCoZ7eg81RKnCjtuadxkB9xSi4v
fJ9qvOU5fi3UlmzSmGqxq3en9EnOFsc3U+Bc/Fh71VA/Dvp6EG5DHkHcEbtELFIt
56Tn4Qx17bjQzOx6nZQtL/5J2Ayo4pFgN1hmQlkG5krLQuO/ivBeyif0x5TzF1DE
HjPWSecugHW4tf3GckWwxwldpnBHDalz6QuryFjWI9qol0PyNdAsANr1lyWMrQjI
rBDEPfDsdCT4dAGizT6sOxyqNyHwhO+4ruBtZlB81YxF0c2L2EotUvQ2CXeOczUK
Bp8/GUDQjqW/8pe8rqeBVqwJS5w30lEmd98lUZQyd4ZchxFWkjZx2KhgeZhchKSQ
LOLdzcZ0xoaXBmz+RQ3gl1qumBCzUSNMbKyvWjbDK1lJo0fUw4qVA0pU9+K0LWyB
1YkRhaeA69KdjLjezrg+Vt2gxzL5Bz+j/WhyLcLK7vT52hIGCzT1hvqTc/QFdKTP
wZ9vOf3dnCn9xYQSRqPNRtSI1v2LnmcVLzFeIBXsMYQ7SCf1ceYumeYUZHcqlh0p
xnXJMAGQTQ7KKnxvCiyhyXE432Z+Jvm468iDRd11+KmFeSgpMv1qCU5uBx6/P7Zy
h6QLlodJn/fVjbulUZyndQ/b1TgHYag/xtKPA8fcYwJV2rbXyMDVgqw/8YZ8kTvZ
V/p7IZarjunNu8VwLgLMKs06uEjmJiej6nN8S2cnx+Qbo+4Cs0AZJdLteplb0u2V
SLYtJprqhN5veFWq+E12Evajm8Y4RDcj6G/byino+ECuwUB2XBMYrxIWm50V2o3i
NBKDuKXRfGzMMC9iK9BJ+WytSBWSJdHCDOmCSwzhe1H4YZ4oSt+k9tiI0AJwpIUV
2pS+Ln6xf1gG8JFYxRwhIsrlt8vRRr+uDGFR5X9jogPxCGswmGLEvfa44OI2QNzp
fEZ1YCy8wHruRmItKFqWeLVub7iFtI8FGcyqvp8SdDhuWIqKH82PzQE0E15rx1JL
T5oWlTtWxtvNGrMfzBY5lJ4qnyFgY8+Hndn5zTPsPy11d9SMmOdyd68wF2WN6WZq
2qLOjmVkDRPpkrILAbZYJCP1oZh4QMTxjgdAaLM3qowDaMcVCJd59lLhd0WQAbna
NcbQdd5HbxOuL9PADxoy7znEYDpaa8ZRGk2o6bLfLhLea1hOFzMw0HQXWJt9Xwyv
oeKBTdfWzIP167dpUJ26EBcpdDlm+VnZZyRnWyOvW880CMA3P6zHlKg6oReyUK7n
peyutNWLVH7wudHgWk/qsJe4j24oCNnAOD14ELrPg5DQysZM8KrJilj6K1HNT3Kh
ejpmhG0IF9JpJwnprm+rbPaRy53gSgB3EaCmwUtjCyMFSky5EJ6ioafSgUZQ6sH2
lQyZ1+dYK7Tgkoy3+lcZc3pCfwuA62ckjeCLSEDoBV0jNVccFveVp80enNFT6GCS
Qe8uv/rPikIkKa12hij8vP20rhnbXSRli0JvkZiyjkiTi1RbZWxoMBfXrTk30MlW
odXXfQzbMz76r3zFW9azSGTxHgJfXmM8LDsP/746wPiBjEBj9PR64gU8m6UQ/Nmt
gfKFsgJs0ZGnzbaP8CPm9xrbpZxpCpAqcUdbiNc3HHqdOh6S4d/GXetyq7T1A0i/
e1gPJpi866w3W2A+bW1F7mieUNuehiHpGhVy7AF0/Kj/OGV5W6rIwR+mScaBx2Xj
RaJtOft+oiXLh+w6TG9I3EVcyDqX8y4Ovfyz0YD2IxcK5ULrvtrS93NgrM2KDZsj
yKWNs42pOWXlNrFyZiRreTnbg0rNsn1krbC9kIfsjUvf5jzC+YOJpPwM+vlM0lh6
8pNMShDSqKKa9SPkNWvGQXnPRZtWqVBTVNTAVvoEnlHyXWlksKlM92b8S7sw5KWK
gCexyH3f1EXgvtdJfoVvFPiDvLkVOxuTnAZ6Gz1JflAWPznyMGSkaoX4ozu+H7Mc
t8guzAWO5mvnE0duK8vWzJUTvB5ZzXKx+mSOwJgKtO/VoA+vsCnxW51+sgoCkImy
Bn3LmYQ2Zk5dLJDQIiXWdUZ2UGG6WBGCbQQ2Z85J5hnVKBefyHGveEW/vbzc+g4N
me4pb5QqVQn0ufNcAzN5k65vvfialltgnn9vj2g5jja1g9GNisxKa9Qkuttl5BIu
SAty447FqahWTCJHUAvtaFXHoDihaEwQ1RnioObjz2GghmpR8QV5P/fMNnGATO0+
eR/rL8lKZEG7kH5CRfiiLu7CFb8IGs1Bl5H97y5jb58GXnpAhw3KYniIpfzN5lZL
NOwq4Da1CJbuyxWYvKjZDkujix55+egApWBXakJDDtRtVaJkksemPdELhPd+h584
21ysYQIJU/bvHWHv6Dl7NGUMSqT6aW6xrYrcppyXGLJTC+mniC6VGKRzVMwTJBqf
w7zOOCyQW7c36EAnS9FcOWuE7qygNAgzOlqOrXzYyf3JsoCJPz+nYEI1g3QD+6Wf
Ugsi+R743tYRXUXNInYzJZP2txkqeg0rw5nxheRNiFZONzMq2Xn9Lz8Y4mfWVndO
uwztdUt01vzyxXh8nXOholr3JVUNhLZS/B6BVhE0u8Y1oNsf7kXS6P34P628uCRQ
Trz5y1xmD6Z2D6bFNmlgynEKAMHjvtBRJUvEYcQhV+23Sa7uwPt26GxfhiYitCtA
eBW/QINnyuhEOiJvdCbz5qr1wY3gRaOZReLJsus/WgeVpvQ95x+fsONWYB2HhF/0
eNnRschqQwR8R5HsdlfMuHmUvRk4ivT4ZWxPyN2+fLEVeD4/jjvjjKzSpOrhV6dJ
pjcwXWucq3MlwUFqDhC+n0aMhq5O9Xxbw1ds31QA19iiG/t0YP5wRV2HadY2It34
YPke1YFLGSVyhUR8Vnr2cLsGb1ZsiIWpPHAec5J8coPgJnt3sfVy0b1dFRaDDtt2
wU8FoaT2/7aqpb3Ygi8+Oe+5xSjRMezd5fXBbdCpyNpVz33NpfCgwpJDi+OR2Tmc
YugmCblNhsmKoNRx+GuBfNB89Xf3lvDAPlmBSRNDc7s+qJDxyuzTGSLn1MOIgedp
mRqDsLUtrl/IW4HMN6BJVdWXVOM6gCwMPhS6g0f8wog893c7u3ed3xp/69HmFK+b
o2IoBuWWVNpPeIE13asS7U8mEiekoguNagWv3GcvcFwrHmk2vliexu3c8SA913qh
8JBbdOTHUprPHxZNxx7UXkmdvAQ2/5fLeKteMm1gDMzOVViL9BxvTaYCozllBx6L
86gf15k18d3opY+1zrMFdMBjqmnUaz9+iu2IQcXWtfk43/p5fMmOKMH7soozBboT
HOEp8m4myAnWXNl91Eo0jZz/p0cOZAylmhrj+/axtwtjOWPX6jYzunc23rtfTCYP
EgIfPu2d25XtSj6jk4bNqroUIY51xhMgwVVhDonYyU5qZFUo9HZgDxyQRyvZkw+F
IrfFq1du8YXR1xi+gaWX4kp3iGZWOXUSSY105YwetX0dCqsBHFKtq/QG57koV/9d
x8mZ+V4NBjwish481GjqwkJore37hOLo65lkU7K6EAnie+LY0yH3+Y8Uo9LD/Oo0
wN1z0vbrt2ZKXrfPGXW+bl6sOZjmgcMS2es30NNH9WjH3TDx7otstZOAIIOMvSqZ
Vkpzoa1lgnMhDVGVHf1kZ0SnFaCE82oknZrVRqUPoHNkjYsndo4i4QT3MudUKDj5
gZ28vrC1vAJ+Pv1mu8lcwOcFhbxNJPJ/VbQosOf2q50980iOz2ZcuahLHiI7yC5p
pUVHw5C93PAP62NVTcwXaCAFxavwIMyGIPOFORBHvCeReGtN755xog1idK8/jRMX
I6HeUOShXYv/qNMrLYfJHfGILNlZ6hdAIPSz1qmPMT4rNe5SR/xN6oRdM+ZndF6A
cKvcqAXaIvmIlywL4cwbTWOX9IfLioUgBmlfp1kA25Oqn3BdUJxlDc2M1qzS1gya
pJPQblcrvW4Jo3NUmmEbJsSgqJ+VMNP0HQdrEAlXwbyYsnx7Hr8/8DJPMKlngkKG
oSqCnzP6WIk7lJ3kEkiksEYDV4+ulBwkBTR71x313OUhngTkZemnp3XdXSCe5jp8
tSpFapB1EDKGnGJNR2c/WRVoJN3bcUFCuYqkXG2W5UedG5RumV33jJGJIWbP/2Nu
Uk5pi00Thl4trmtLslrFTBGczw4II7T7tOU5ZWiZ/VSonztHKL8zgpLq9PvCUsj4
zqLndogZ7NF2EOw9h5mqT8PAVpmpLQQwEGOVR4Ov14t8KQN30UdIrM+Twt9O17QN
h4fJX9WPBlF1wDHryTto322I8O6LojQYewDLq9+297Jd0gJ1Opfg5lt+fUtJXyHt
pjQiSb8yqIH9cCw9UdaRiAHp9ENkHIYLyYhmm1eNG4zCJYthFSUHEk/Q0AFBkmcu
WXcIwfRndoZhih4GukPda97r/jAT6dqySe4ooLFaHnh6DiWGX8yCXu5G0gvidpuq
lQE0ERcBG4dimAVzXIMUx+iOnwpzWz3u8Nx86uoXQnQiZ5oxweWzCHLmL8Twtw48
I93+VY1ZFjZ53hLE4baisCeArYAhBlsDuVapMjkPURTu6TKe7vHRwsCe6TTr87kN
itEt2xKaG9H6nxxQ9tK97hKl5GnniBO/Pno2S6ab+Wmaewzb2DXpYh2SqUwDWpNv
rgjzoqbTxX9FWJrePw69Yi6Esuaz3TfbpztTpvH1ecWoRjfZnaIOWPS0C7xZpYz4
ua9tgO3o1BBBvbOad2Fc/jjJeeJdYSoT4qohSzsSnIlIhHbDaqvhq/IxMsZ50xjW
8lSA3xkTWu/NzCS8W+CiPPSYOCA+CzLvM2z39WGxEybqH2pFggrrfLDXCZdOudb0
ZBOUQH1McQjwEzXuvjgJul3LpuyIjTEAbe5vz2Rxhj+udfpRa24eScXHx+CDsUho
UrKmrXPGlYoj07XMkCd7fw+PfrMVZqMuPsnocasyLRMIjepfSFczFzVW1Eo9TPrp
bYxmDVS8qM1/H6/eALbl/jNheY6PiWvwQ5G7KyTcnn2aHkbBaYhpr5pbpZDM+3qm
SsmYL3lw/NUldy/DOsmWw4cP6Bwy9N4IUX+r5uvwN6xmTbkR4fbk1gq1RsTRdteX
obe7EDuFgAnmXKF8DteZuo8kNsMZZK47QhItxSoENZv2hxtt/NMQqm5LiaIGyoPz
J+Q1HM6q+aBHD69J22bBSgX0UnUaLeqhlJcl1DoKliR5CVo83srfThP4fLX+UR4u
EfP8/7ZmWwjS+snIC2ACxp3tjPsYDA0ySeKYZY/x2Th/SPtm/QooKu7zOQ5RKYFk
RVltgcCRLNka/Dvaib+7GEJeL3RlFBKAnYtupEhVDbI2RrlEjbOPDlzeW1n3f/Nc
chfuPIGNnGzX4e/h2x2sCWETyFmYquHkluk3LVU9/oUvs5e5eI1Ya/FMEDNf0vcb
eOV3UgwH6Y8qEfmvi6anFfBtX6pxrzch5dKR1r7d+IziqggA+Zl24ADqpa2cn+49
bmeHHU3aVc1KQAHxhoVdhnn4p4RCSsuA2BUyVIansH372WiszG8vE0wl2r4dq+nu
lsQF+8TJfNWBJy+Hpi6jVnRbLbML6Eeb3PgZ4j5X/QyBfI+tohgDRco+TNGxp2L7
HIl5h8uVq7n/fVDyNeeET4zeTK1rnpncRxEcza+N7w6p8PC8llE1hwRKTJJDAPVz
rwLt5F27dhLLBlJ9QT6ZyfKoCs4rKH+z3LHjmqURxjl2K7wKsYrNTDX1//pnRW6M
SzqsmtiP/NsfQ2M4uYe1f7NO+ZuRInhUgmWMfo4TPchfOVYaeXiUnCBqMLQuEuj1
r9oqbRWZOB6Km1z3zq8WIMbDtHkBjEyTZy809UOCg+0olhr5ewl2BCHM0Bxiwbpb
cUkWGHA4lWyGas0JWXHSpf34dzCSCJnczO2++A9Cc1a4LdS8ncs9rLl57DeEOfmM
biQKGX307c4MhndNR8c1QBIRJGO8EftNVT1W6tgF38WfmV+2OJev+0krMorit2fv
TbSXksl3DFtXJr2v7ol8ZHHeB/F60o2bsm4mP85FKOxjevzSEHumzJPvc3unW3C+
Lqa5B6iy29+UM+mABVVAw6IaJGl4+SWb+dbBGy0kyoNIFnBftjyNfX6cn+cGo5UW
2bgAEckboj1tc5Luwz+DxcNgMIDCrIClv4tsFgooQArmgR4wWgxDuEOThtQcgASk
fiHfwUvH+zotwKe5UK/5z2J1ZuBXv2wHkBya54dqTUEYHfH0df4R58QDneUx2Tei
obYY2XKWs+axNLGcmIv8/RkvSBmMrOcZsjk/mkxSCvG81PkkNhHF7b531efIRwYf
7kyQTwv0xseibyunU+AYzq8wvZ15jDy5y6Qk4kgOLdp8VWGPfpIlxmQIlovBYh/u
jRDZZJuit14/VhMcldT4jLWUJRCuCXbZY6xLPcN6jSOLhFeiIKu1gfPFeS63ZOa2
NEyd92y3baU7iM6sSvmvUmtt0SspmbMIGFH1n9FJXnfkpJqmB6qdg3ovCwnzfW9J
LuvgD4mSZc77d6j9oKDIC9bPETiAr7oo+S+0DgPozewxIi6+dCmAmvHkcQa3sD55
dFfSYIx/YJD0krowe8AzWqmsat0T0YtiSPP5P4EvThffeDtdTY0kNmHAg3Kt6IJD
lWDG+zuQbykcgx7Ie3N0sL8wUXy88R+LlHnJzX0hylIA6FODyzdAfJrA9wN/TL/3
nIRgDt9+o2xVzpJm56UZJnJ5jvFTeChCPMiAjDOLsuZojgdz88yul52wbc4k8QCv
JNYO1SbJEgtf9dXCyg+ifyma60SCgL/1FYHLGPO5Zr8EEC6ryiWOUFNHfl3VnATc
ONYxAK0SRfTsoe8tVn18q9s9n97V1sOzbRbQoJbhM9lkGvOsg0xphWpInPTmU6ko
L8M/ggPxIAJLm3s+zdNeu8nmrT0ZXQ8KoOe40WW0sM7h6SmGIyioGwRaeICrNIDa
5WdmfMGrch3TgRgpxDOPlFNdZxCu3JODqdwezNjvu5a6K7gLVe+NgEvwL921Hs15
wqjiqwWVYpa8Jy4POHxe/7eiefATtImaIZVKeU6DoqmD6HHajjG+WwESStNUqfdU
ZqO92PnDg1XINepbxCkJiXiTU64Bx8yESCLOgB91CBz7NWDCTTS4NU0iWQxyeJKM
glqOuO29gwijKcw8CxxM2hG0YJy7SP3ahvd6Q1v+LFssKsLQA6K0dRp2U0mJ3DEJ
kavndYYnMOgI3mF7+KBmDQQhhDoPm/SGAL2a86JNnXNEalOixeRQeNrtmyRa07ww
06z8/2Y7bBN7jnNX04YFwZdrcR8iA5F/qlMis7wiw5xnDSrMBIH6FHSWPwxUrjTN
dgJjsv2NvsommA04uT5SwEcOK8sw1e0ISsoFDT6YR3xFktw1jDci9eq1UbTfPuML
ClmJ3erik0i86cVGewr/AQI115TqGR4D985XTkmbrMEYMRTenJJpZx0/NIZljdYL
E7PU4egD9GycO5pBwwmxO9AHMvMRXW1T85fOdRxX4jybJowfw5J7o0lrvFOxUoFp
/WWVUtpK9hiSrYcUyuWadlQ1FJigq/GiqS06RSi1FTfWWxL/wZ2tQRxus58qXaSk
JJz+/rvp4z74Qjj8qxrOz+Id6wFVPMZ5s56pLJI7AHoNs0cPlvxzjDcoVkBstxp1
a3cGOyI9wwWXxK37iWLoCFlpjougK+r2/RiG0npHx18OYxlycdKXD6Rji9cFuqIF
ee8bipUUkEupmnGB4SJYDiXSI3+bOW5Q36yBgRjh7Biok3OmH88NpET6uvFKsg1O
kD5Fu2GEK7DupL69JCtIr7asWoZbC3YkJTTzJ6TlMTZqoCTm7xF0cYt9WlNpEjOq
SRY6LR4xMDo6CRHOMP5SiONUgdHlL/kesBZWgy7gezACqYRSwO5MFzUbbdPx5/yP
hbjVCpW78fDB/4RNPN53BZIOjlwIIXtijKYEeyDIyH1nU8lZ3MZ1ve02M3mSCNgj
esF93OMlMBxHd/AV3AlR2pMm1q4aih2p2AIgDplUFWtYJblCyYo0vB/YJ9sywIMz
Hk+Z4yh9pI4RvTE5Y8P4d7YgiB5ovkA21ozMeLHuE3zN3FiHfIZI2l8vPuJGrulY
hadOD5D8w1rSY4t2pzSnKdD+svTPbZa1Tgyqnzr/897ymK49KWNYYZ4PcMqjDNcM
8OWdJcn5R1xXUy/BisIFVnV+sSNO3srMOK8rsVblFlb8ZzRx6/sMkhqsWm+jFpAh
dpwU97Hk8FlKor3r+Z/0OaTRVCKi8SnAwGnlMMGu4VVD4S7Zc5AFCOXuLXb0SlIw
A+4v/dsJImh4iSnw8I3ewnxKoPkEj9s3AKRHVW+ebKT3nz2rhsX/3rwqp24/bWyx
yWaD7eGy9rdnrbNwTrdVlaYwvTHhNXI4LGhJlPzgQR47tUafK0Nbvlamof6J19Rt
REi7GYaX6DaOomrNxCsArnCkst5FiQ3eK/o0yO2/esWXio4K+ObElYGgYRGBtyd3
KesN6JOJ5SVHnHCNlJA8Ngh05gWRGottc+20kfhum2Tb0fNHHjoCpdW+xpt17I7D
HD9IT04wyISXZWDy5oKXLYy8taKJNnfWnadyBpEyE039Wc+8JFD7Rtkm9RnWtqez
AMuX0FnKO74xj8CDWtB79OZIuRMcWZllvdK/dmqHa3gQIEYTL86CvvYBf1+3zH4m
mpbjFSTKRVJbqW0z6emCQSIcC+ijikJi0ivBN1gkdoFyamaABp6wzQIRb7HNZdhw
3ciO0QSVueSlYF/+VYclMyNzoqKBDbOumhM4N81eENoPhxsLIhBkKq/wdHUjw5LO
N18I2MuFE6PT0HI4m6Fd0vDWOKgUahmYzhziNlh/FVa50+o7RvQsrT+r09z7z3JO
b1gINqnjJZ4BPfQefcDSftXxs4zMbi3pgT8ZUTe7LG3s3zi9Cs0n83akwCU/ILG9
NtTR+yhHgsN6s9tuE+IB4+rqHUbOnIchDhUR3bxPVt1s1HNY+OQA4Zmp9okblPpG
/iWNC74mxf3I5dUNfIECHnwiTg/7q5eWPj3fzoy4oVgB1C70kVffI9Ix3ICAllK5
HQzYYnR2Oj7vn1EeBy6m/9h/vooKXvPi9Tw2NRaFyTEjEe7653z9Jjl/nDAqBTqW
qj6AB5gsmypNDKUBABp5ApXunvxnTt7nYTL+XqMjGXWQi7ktw060bslM8g4CKTKc
FTYyatcU6/5syJesdv8Q0sz/dNmNUptcfNSICBFHfbTk8WOLlwTHZLI22ORiwsIr
Zyuw+phR9LE9AFHgaASy24wMlhp+q0Ho/834BzP/1H6C0K3Gzt1u1umSoOLdLbXf
vZk/DnvdWlQ3Fvk1S6RY6UFItz9tgG2/NoxnRTfytJSFLJAGt7CR/yYES50hov2P
ZyC+eAOzCViY9qFoW3DpLghN+zkIoLnyaVARRZ8mZgv2s98edMXjavrj4KwXLhIF
B/jxS5onJ7N1dMhoaOQmo5jKD3r5vA0beKd3VWib0ezFJ/wgBYJmh7YF4bRVBGro
zomeDPZWYoAJVQLWmSOWhWEMwfMpuxYRY/wAEhbwpiVesjHsBGTZMoJlSESuNW/x
HNFac3/ojq9vFNwQjNmo9I7eCgfSnveOjUZNxCb8mxgT3l7E7v7THV/QORziCJ7i
uLOMhjHS6Uym/uwCbVmmuBKrH+N94kAirPSaUhI5Oro8OMOEQZ7TwFme7aGyOcrL
eYDW6gkxZ5msFZuhkMrympLnMkUiL8d8MMGQJEd9+kDqu/gzh6N3y79TtDDEJKsT
0CKrjgqtuXFelOkBwoJzVvN5BOcSmE2YEQ6IsfmZjgCDUyyAGp/lkE+GeL5GoxVA
m5e8TiSW46FM1IqEijwdh++10xmz3e+qFmrrLa+UsCbd8+5YkbgDCugMeKAp+fDR
m+X8Hdk1KpNIKiHEzXKyiK6JelMsZ6cOfdoH60XSm/1Prlqxr2Y5rCJChS/0mVfW
B9hdSaJS9LL9basnsrQ7JVCgeb6RkVkKwzcNLnpOYwDXEiO91oxiPBRT1b7pYJhg
xkEUk+1OaiHqqw7G+oSZS8B9FaVlyAOzBP9D0+mPDOf+N1MXofv6HbUtEyN6kmGW
ItqtRfE9SLJNfyQMkrDllZqKwIDmSx4ipSmwY7L/vqixiwOUEfFyDCz/VSrBtXMT
nVBxmmXSDZm4Yz+MQdHWDoQrCVp1CMYv0YqnVWaIXhIzA13HTiqJ1if2cJ4LafVS
W1Ss5mD0uPtcwhWskk29PCgU77NviDMDeQOtAaB9hLuLhKMtciXxO0/QvUdzzQMT
3FHJ4RTLxBIdDyusMmDN+8IH5EeaNwN1fI8KF1UHnSafIfzAK3YnrbtEzJLYUzBD
NVLMzYBgr+CHRQaEymPHYwS4NOyue/gUoIHCKzZtkGOgychrw0jLe0AyN68aD5QZ
Z+MTfNz8tp9eWQie6yfv0HYUTGHDPs+2yGzZ9QgkJ9O0Ll6KpjH72yLaAHlXA9qE
gn7B634J1mr7SG4JDlKTH1MjQrSE3vbcJjGqlz4inuGa3s86LN5iuTfwGODvIqNQ
TLTHPVXWmwYlEnM61eBVKgDATZRvOBmuVA91OR/bXiELaLwQdZzoLvyQCr8ug0+8
Vn1PVdlKeyzZt3RQ61XrJE03A6YwBGG3Jmfp2j8LoZb60Mb01u4scCDFTDMs34Za
nZRtu9T51XDLvjUCwNucFbzBP4+zvsKCOCh6V4qIBvfsAnYN+UGJ533gVBMLEFs1
4KzZFq9jXT/zs2himOLOAAo4JVIF2T3Vb6jQwb166AaGrZc+NnPoeF6O0ZJgnQi/
6BO82yAUHcJA7W9iTE7dkg4MHEeJg14NRWJSzp66zGiUiAL2dZHYkrCNDQlDupkZ
hRw6hKEZ3N6Sr+7Jp0CJe63A7BlPKN5XUpENp8QOitUf+fC3M8YC4ujavKKWD/ib
ptkl/LsQdSGuBwoEQiswYlBEkUmy4MnXbwqxjb9wPtn67EpIShholx152wD+Q8nN
GLPXLQVTkNB22w35OFTZd3Gp2LUFDZP6C65wEb4oOmhYOmBxrvfER4dqgYB37RDY
nknF07W34IS9jF5/oBsVzn3DOyb0iSqbdx5n7P6UzjVJr4fYzpeqXAkUegqCkWCw
G4FQnVBILgGHuANdh41lO22bW1T1iesC/1StIGuSEk/HhFvfmHvc7wNq5sx59XpN
DfN1xqo2G0iFbtOhyv3OJfhosHZuKNE5kcd+QD7ogDXI56Mp0rffZaNfyItjSbjl
qzI9vjyokVAz3JCTPDmhvTuOQNGzJAOVXaQn+lo1BWpntXH5N2NntE0AM+BDhiaF
YA95LI9QtmrhhZL06tNLrhw/Tv39MgoEubeRGBqQruvKdWQQCfcFoDSg7sxoF1wT
jAFX5zv+eDVlIw3BJz3XD2Xddvxeg0AVOXfulxEI7K/q36ooSxuSP0nCU9HCn/Hq
1Lb9xVyM56gNPIqNgCkwNK0IkYcXVlE8x0gsMw+QmNthIzBeL4NkSrNj2zKeNC3v
uO9h5AskgIf7ic3Ah0Fyc1voWJJOR+pQq1b2VOegD3v592sZyJS/BHku8CT/9Uf+
1OcSsyutOHWtQqZRwSoSk4QF4soUGFz3MlIgaJ9J/ccx2odm6yrsl0l+E4LlNN8m
w7HO401vYpXBhuYMad4byyIjJX6f1Fh0YKxOdras7RXO5TP7OniCkVzqe2n3rOR2
uNpO97t3xZ20Z2mVFvwyFbK3cpAnWAQ2zwZH8qKK3WX9OA8SMuLq0fmLacJQ+1CF
5gYV8ih5H3NLinO4/2vhZFr8DFUQOjSOkRs5vMusq0/jz4fib7tmi8Z+/4irxJfQ
wnGo57KKqVVYpTNapVniQlf86nAGgQFjkOyQCNEYffYdrtqj9SiFqhSDHyJJPq10
itYvNhzTk/y6C0kl5u6MYIUMgbiYWazwiTBAnrX9MmtK2oozOymprvT2nS3MUBUi
W+4T7WXSoDfXvAKq7oxPRfl4II+GaT/qBn1tEDwrfmqOCEGRRcPkt75YPj1wLwY9
iysoHf8qLN07JtFwbtw37R34CIvE0ei36HkU5ONI5qv87wLFB5BSk6smCdjkaCLi
VFiyZlatny3he+0YjDieZEONafTcXFeTqayL/qMwJaDmIw4t7QVl4bTohOA1OGq2
2/ujqMLs+R3qTMkNzjYcyHwY/L//nnP+hkp5ISyX2KyJJL080brpcTpF5gGURYYR
mSc2K3rAA34QnovMgGpXQQ/j5MjYhr6v9BSrX08HAyFKWKBIv/Hem2zyqT6YhzQN
kSqtga0bMkMVVW7dQJc71naVkF7RT9s9BWm+H4RJU5gQsEcBHu+MXWykLLOIGJYK
hQjG0RQU2CPO1KcRtl+b761lkP57QPKTozIKOWYk8pl8dNpe3ryvOY+hOA8dcKrj
0aPbXaAsccbB8MXDz0B85RW/6/gaB1QpnnWKyCUw5cfwyVrq5KAWXmaywKGGiT5x
0TE01LNlwhPsxMIhb7vZlPcJvcsPwKS9TkVXyEJR5l3HOAOufJAMn6BqYX8mhJbi
Fz/5dLecaBB2WHjnwVIbsFSoxJP2YFSReWgscgFOX51SUgsq3CWfpURlDQssRAJ+
OMwEbIJ4xQ//sT9hCx7cPwzI2t5tcqr+Knk4cIDZrZzebI/u1RkBemfIJOi3lkwW
plgGKPGOQqpumGX69d7fZQj4t4KpB8cDFEP7L1ZD5FRJS3C28ganQCaDbnypogt+
ODKXNz1Ovd2leyqRuPE81UXIZEOhZ2DQ1acj0Cw/rRx/Ed72mY8PkIJAWyrKFT8K
OoimvD4hLFjWiPwo+tMA3SBb429nb1sVdJmmmRwy8AlmYx9m98A+t/hPEkQIxlly
+sISMMNrQfTf+i6rS604HjM8vMVb/gap1UN6zD0z/J4YFHgApmLrIuhFDotueTCr
KBuWejsbvQ/FwojJgRW2qYj5Ecz+WFCo6b5OOEYeWnQCTOm6SHXUoYUsODNBuL8Q
vbEecu84bGh3IF3dkyjkQTwlRHwhdu8MDWWtcr58Iw/B5QZ6HcBwxnQDC6XHX+3b
/liZElM/yCVfL/eLnQ9A7yKtqs0YcEh28OOIeYTbGCPfjvCNwamu/ydSi+WGwOxB
GRY//z6oT/FuyeYW37kDw00p2Nr6/xq/lFUZdJlbKYCapBkUpXLWJOLWDe4bQjUD
M5cMwRTlQIXGx9ZQhrmg38NzoYIefZVEeGZyD9/ESzkGmsn8fefFpiQl7Bd6lNlL
NpkskhtLiqk9xWNTjSiK1CISO8/YwQJIlA8x/atd4vLx28vnV6vxMtb8/Vwmf2xM
jtRWR2GR19s3lWLCUtrnoeOftxrJKD2rV5LTg6c8lH4mKdoaULz9S2H94KV5AKE9
cR1Vyx2YrEN7ojiITLOk8IgfxFbuPOruhtD1XH86UkkzFfmUoextl7vyj1rGKmBe
2ziCQ+8qNGJunyEfaQ+vly57++PrUTW91p/DMJKs1bPqasmm4t/sL8JkRO1l5xA7
rpqTsGUDI6WbNy9u8pbFnxu3PtkeY4+W3WnXZFamganniGCiMitCTh5I4JxzOAXS
bia/agC8iNyWoTfkRjNC6+ln2Wd3AlxvWJ3Kg1qlocVQIrX1TNqyUKVhqNgCRzO5
UhQYeW8EGXxvYItSJpZKuigxX6dq+n86Si5swVDWVd3kkjZim7JPMLSP2vexhYJA
/lPkyIr2ibVCwgzqKeWoJVzIpOVmdlLArWUSwVh/t6pKJmvNK2aJaPJWv4gDigR5
dCeLZfIfMjNf8Qk/MSgxRTBySjpIPwe89wgXvtPfz+lYG3FQGyo440Cl/yQ2wp2I
4gtu5fComxNtmOSGZ3RlGciq8x3f0s7Vsp0v55Lgy0J24V03XicVXhxfBbdrb9qM
t0Rkg2ZpJ8CYHf3x+4kTdGtvTpm5WAQ5NdQNkP6l9ITlwUqUqyf5UKogsIlhxEzR
9hzLz5rv1yrZAI+qvniRakH88V8NE7u9QacK2LrTlqgypHb/nLYpq9op+W6zAcQ2
Un2Mooe0RaB9y5zd4vBqopUeVJ4bwAtS5iQoYVa/rkF+EKd/hEMiBEnjGVp7+Xzv
rDWD55sQZh8NjhV/wkf9NEqIoZLwU1i8DeRn9LpsZFtzk90xDRzBq5Jft6eyfdAl
RfOfY6v6DBtZUrzEAf+fLYqkgdfNLLzCmMKAwYBs5Yk/ig6HnRV546uP4E/RRKYK
cGwynwmi9HJrNuDPgN+XR7+nKamzv5qUeUtun/L0JPtXMcUTd8/smvQ00Sqhj5iF
gfzW1l79SdQJCnUjVw2mp+/Hm1TMc9Oo6gCmbpy8XgAPcD1n0tx3Dw3P2qzj4cMy
kG7PDgXOjxVad1ERuda84VQIQczH7fz1mE9flcnGpUsYSgEDumOeRrVRkAWx7Sho
oldWrJFZxBjWsgnrjt0z+YNcnxFZwhJkVtf5XUkCcGSh2Sj9/cMlpqVrBVob0d1L
FktrM50nvwlktTAFcLs4bv0lUN8gZ0B7vfY7dbx0PPH5NNq48whlMXBrft1Mgvua
NRvcRXtM1sJrxCfLY5YEMIXCDSGDl/sr7sMR8QbtuUbm5rhiTCQVxtzA5cBnT8p0
U5N4xiatoiHzAvYyyR/6U+emRVKZd76LDDl/WAAF5ce5PFYLNf+P9wkvP3LONExx
Tatolo9U8Zqbpoye/vNUepl2vNpscz5KHav/2aCUIZldOhhL0k1baQ+2d74rnciN
NEMTu4FhUXhBpdNgQiumDoELxDD+cYe8Hl44+Y4Tx06EFJAHVufkeW/ICw66gMlX
6bCmUBu+iPqO8YifgOGXoEzIvzJgS6fWluv/8BoHg6JQucDo5m8ybk36hDMKh8pF
qsN5wKWkOZYUbw8l9FNj3WXC9nASJprhZhoc9BhEs5BG79iBGgGVKoCI2suUD2aA
mjQTRcXTAfgmHMaHFJom4yA52mVrXDcqhVDp7w/UY8pwJtfkelFsfyB8eYTkM8Cl
hy46JrjZv0QD1jBXfSzIA752qkSJ69fPARtMIgJv4UOZRDXomWIxdi8NGpCWuoe0
q0uFxPW1LB9a3pvOkHHZRVgQym3R9M12Lh58eNfI7F2nxgq+FuBT1r7OlialsFGw
PJzPJO1xCy2nP0Bd0qphnVyk13KpgwXsUFZ1OGFkUYabxHTM1W7rottXtXYviKwN
83Z6jBpoEYnPrcpe1Hi0KuG6oZXElvE69tPYRXFkbBi9BY5vfRdBF1Cox6tF7CUd
9xW6lcChfPLSrB3sS8MKHnnEy2l5iLchzUsHh+CUDvp/eX/4nZcK/Opk6a99iV7B
o7mLHZNEse0D1ZOzlsOtosLBQ7soFz7q+xmXm26z2heWatelKEBfXuET05hE/TGo
iEoC50svBmVIu3X3wbL3xhIlxSaL6oEV5yWj0OMi6JKJ96y8eVK4U3v4Mu2YI4L5
ych2wAx6GDTJsuDV0pY5VhvI6JUUm8GjauTKVT0K3G22tf1hpCbETr0KkjD7IOpx
ZHvyfqENoCNzAx2e7uQTnHjR+zQk09eqJZMVfUQ7wWMdoytMbCD/N2O2cE5jiswz
GkpC5EQeTWR2LC1LDfHnVxx/w0t3yhYhClEeWlzjWpHA/JnubDGsZqJpH7B6MgXs
fgg+KW5qxIxVewcVfgXGCQ0iam517l94aK3Ee3UGZ4DxQrFgoUhok+Vv5R0dgzJi
+6Ftu+XmcqhcKp+aEXkrQoZh7DLUlj2DnFUwTFdhoK5P56BoWBY+d+UGOoM+/w7P
U0ZbZ0bLm4BMc22YIymv5fE1chm0UVssPdRoOOoqCa/K7q7tEvsIAMlIuQqRmgE0
JpacdEzoNxitn59zL/mc2GBI+z8dN5il6UYWETwNBW+gGbEFQmZlGcLWoDocHt1c
7rmFJv/vgIRoAJ5xEperCDc1YLazENzZTv8tQC5opGHoH8OZo8BsMJQwmH3aE3ON
CavOZkT9TaTDoLyqzEvtmtRpx0fGyuU6Rrphehqv6qH9h9LCKSAEBpyN1y//OrJR
c5WtGWLCPJ00S/WwNcKPrihwrepvJUyxjn+QzcWNwT4Ec29PDEObD2QTJKIRp1/X
i0+pl634HBitCsMhzHTS+no6Kj2ZJuzRKiBjLO4yxHeup7iPW7+CPt6Lg6n0bW8D
YxUGfco7jZPimMHRmWeQlnsUdwSa4IPcYer+I5omjElv5BQTz7wglsNQupW5UvvD
xEMPLx+pEa2a2bQ/pcNk9gzile/RrCYbd+JsiZ0/ansG5AQ6Hf9tmqA4CFQEjlQh
QILH7jcmLVsD7urTEKFhU/LfFE/OYuPHuVtzzgcitE7LrK7sTCdmsYbGm9zH2A/g
zvdyBiW0IWV6nHSZtp8ODWvMR6+ZqG+NSfxHuHr4hFpyc5DNDZ8v/hAd5RZprosA
T4MT3ZyqxWgAENhr1FG667Lg3bta+4Nld0dQ0HNj0NozZFdpgUETn7W21o0PGe/D
aZtukgJIjpFT2+tiAQfhPNMpFN+tCj2GA39lMG/ukbiSGvdjvT3eIrlYNm84AN2U
9NjgbcZypFGnz6FwOsq5VSkFqWSq2a0OYJWtFhBFM/P/+82OiBt+0Klk/+OsnfIb
52j7eMgRihVucBIxb30V+ruXUZtWpfm2OrUrpRJrfNWKq9u5v2+p8IhTymL/p162
0pSGJx7curcZeHRARjoRFNT3fJe7UGLR82taxszd2foamtxxu5afPwxszrJpO3wR
I7gssCiUsXq6N4D2YmLHt7+qcltsBCv/WqdRiIRTCloVz8Zy6dsVWp7c5OQjRSkh
zw/66fIhVxxgto8Dn16Y/SpdH5QHlx0KDhYjXBfVRKRNhZG9Vhzn7npU5DW/N/8m
vx0VGldPH5DugNo+aOIYZrBwxneoWONufk2y2LdHKUlql19CGoEAgrU8R61s+2vJ
7WBLN0iuhYgYq2O2vLiPa/S1tdCmYb74of+qzCSNs3+4hr9aOwjgAiAOcNMDYDT9
96yCxVlFQ444xsKwtnp940kZ9qBOM7Ml6mMlGMqSXo87LTxvvE7Bd6xco8WjxA+V
CgerDoS9TmNV6XD19CO/1/2daIXc9173d26cNjS3XxYHbees/fOYZYb/ix/aRoSH
U09XyPy06aBsOdwmUk8Wk0NUa92o7e39+/2l2087tWjrM6v42c1b31+cYPYockXK
xdmcJuau5N67jX5bAQgpHq0PI26yr6BmxwPDFYa19X5FPyQYqfEiTRXcsNBD1tuZ
hUIFUkpoPfm7OP6Lsa8GrlZTcQSWNfEN1OEvbB9+FjlMykI7Vbe3aAjpQfCbQFaQ
iEAKunIXbmH6S1HliOJKqY6kyikCJEOk5Fh3Yx2qUsgDioaxK7u+AiYMLyLrmaUz
ZXlXtxX3UfGseGJ4JtZ2GrHyxu2Ng9D+Tu2XUjUVbjVae9CNQXqRD0pmlme2DMXa
HGDutkdMxLyfWl3Fo+JhEoNjndXHqRXtWSy1fm3VK8zkb8I3RWR50jIOQXlU/WzH
a3iGGIq5/XjqUjyZn/vmfnMJyXeZfnuwhlBvWUFRlYd/95FcFS7urFTGD8RIRDnw
9IY6Tyrimed6IJ8Jnzgnc72Bhpqqen/Whrxwka3cpqyhVEuesKuWXB+5fUSCymt0
5s0oVjLtVgE5D9XuBOBPF09M6kJvZiiG3ad3P04PEAIbvQUB0JxauZz2pIqnd9EY
TQE0b5TFcCJOV68qpDgr2Xm+k7svrO6UUOyOWDFm3p+Lis/qpvrFpxH0Jmvc17H2
3iN63OV3KJVO21CJfjFSSkYRINBHXLpILV+YFGpHixn1DRwzCcGTerRdYDgqWESt
G+wt6e0nOeaK1VfxUozuU62sNRXp8zClt1wdpGfbdPIZJaA5qop77ODwA3QLtbKM
5zjk0kRCG1WyGuB0TcpJSvlL9MrRAWK0934CeTc2CiWkua/N4GoLPmqsLFfYwA5N
Bq16NopiEM6bftpNnd8zr3+I4eeR6xB4isB4lf+DVlHAu53Ne78+dFkTiPaxy9MB
3paIxiBWPGjAefUyR4glil0pIsYCWqklaZ1+5E5sqlBBhuppM32bqxtFx6McIKJj
MEuyCrJInNGgItEjeUboS08sVOS4tpMxIIRqjmHy5Heh/KIzDa4rZafzIY1RdX5t
Cw3NkNAIoGGI5tdUqdlGVN3gsmaAPUSysM1323CuLevS2SaHEDiBGFmBv0FUTufC
M7TO9zX7C5AI0HoPwynfAwLLamQ7+Kh26VLJBTjsNoI87fbGkwWyU1siSzXK35rm
65WxixKXcwPXJ2jNgN1awfscykyQvs3qf+R6tb3KLz1Kt3gXIuEo7L2hOf3Mkraq
Uc7pIYoKczxMWQQWgzpvL4yanCbz8hFB9UFkCvYb8rFzstlW84/ffNQre+F0WlaA
2PW1TEuD7CttaMnHElnnz55VqbX3jLU9lR/UQBHSXX36sXAMUn/eS9J8tR14KJgv
a5ZzhvooYWdlnL9kvXQdoCFkuIDNkthzQNfHBMMhIX06tQWqcZOv1UUbl8O4MECd
ScbPLRCAYpCZJQ/FZsJsZu/gp5M3cWSWZr8Xp2/E2br9FX+JSwNGRaPRTwmL5oOm
IdRlvoSK8dvT5gxX+IgjQHKCFvnyzeuVdP5jHkNuRh8tEurB0Bp1bWqnkPME7k+M
QGdkbJGtlSFUNAZRN6zbYz6/zsuKfunUfj0jOZdbX0OTvdQ7fh74vs8NX2KYrw0n
YATJLYdKvbLJIs7K685nOlTxw3wN+bIbV9g3B4dC/4XtWO4ivdRZsbRxpKJB/9aA
qk5zlDJhkwfP93XL7jKPztDMhV22AzOwSOioPWkKjDEUwSGKUrXOiMJkaGADJ0Vi
mKh3K1qKVgWTobU9CvWT4qjFevLMN0dpf0iDMiJbGyzN2y7UJCjO6uMhTfZfYQqA
tgDIMw6dHzj5dcf6V/qu+bw8zGTP1lup42j+jRU29LVfSUD+2VA2eNOa4XYP/xNB
IHMZhQAecJusB9YMnYzr8+jGiZOcMlFPvGvWEEH4LqUDLp2nchMz8ST+dDVcW35L
MLvsamL/Rc73R6dl8Fss1nJIcP0MOAKuAWz5NWPx4OQ1HNinSA7bgU3LHjhswrlh
WV8VU0LR+/4Y9ZuVSW9/k/q5RqgKklzD5Pj8XKCVhTDsC/UWhvYH0C3bqV0T9UAZ
QVCZXBnfLWf0GlvhVAbSiNlS+8c0AOWNoPODh4aQup43QM8HuK9UgwJ0ZFjGlNY6
qN6yhXrApjrd7UVZs01/tg/MS4lU3jIkrYCD7msR4sj+RPeXfNCRl9OoC6o+f99A
8c33Jmj5QKTMBGqsBt4uII2LITcjuwRNr4flna5uKBQjmbj1XTeGW4/2l2YlcT6k
cZQOzNDj2G87vK4wyanz9mHZwuxkkLQMt5JDBAb7wSZvpJpVbemvzrYP4IJ9RosA
jVdbIvvb3irTX/1aY20HTkLUHJ4DQ9klhqbPI6r4NevC0p5UIXY307v3keaC7Qtd
3WnWjVKoeVsJiEzFLCVKlAsd7/84R96ZttStZ+q84kNoOrpsUgKlk16cICtn8mXG
OT+p3PYxEVLlNi6i5YC97MJhOzLWdcprrtAIM6OnYmr8arv/Whg9dsDL6LfDz+Ne
s9FVupZTsxJm4RNqPjd+B9vo9F5k9x+fa+qZDmSLSDfasoAX4+/U9oqeMuCZJn59
fuVALvqfLoyLiF3bulzj1rVSodE639uW8eIoWmJNHHRZkGRzLPP0SLnWJjpnEHhK
0szJX6Nd+y8bFPpLC+NskkT8uT8vJU93bLfAEO/YNwjs5LetEIsYgIUukzjsLhRs
W4zifz7fq0P0oUfh/4BMc1Kw/lLlhaanPqy9UDYBUERp5SQ7Eabg+F4BA4BN5oZ9
oKU+m28SdDd5fKpHvE7w/DWp+SpZBOatK5zvyoMg4RhHYpWV3MT7M0ACZcflPJyd
nSkL2J+RY/cuRGrLUVnUUkePj265O1QRuGRUf2nIpGa6UdHQ38ggWhyzOTihJ3JM
e3hpng8KSy8oTSoLxBOlGDy1wCyj5YSu1hoza+LqOKtfCNPaURKJn1etl8cCjQHa
vAx24LNttRjBizK0BA7FEisqqBGNrRLZwhh7dYorx+b6/ZJq+gHfQnVbmPQ9ldLc
NB4W2Ua9yCa9O8DYNf5nuiIKegqZemVAYxVI16X7MuYkzu6dmwMNjeRTpHHu44vm
gfFyXndzF6zvX3gFvZOtXnv84zLzb+13+a7Aj8WpccujezgYYZA3WS4lyxplqie6
j2Rp+7JKdzj5nl8WEv6fhP9F926EMSpBg29b7zB/8wtU8086L7t85MNLN3HiCeWe
1r6iB/DguTXHf8A7BdkrH/JT2a1PKYTANdOExYNcBsQLS5tWpQk9xxQvf0mfISCi
rxcHTubAnXK4uNjqT7qfzS+FUez8wUk+fwayMYrzfRaJEGhTOmH16AU7mQcxTr2c
1G1IMrP815VFUegs99VZGyXBUb4j8n3zVKrOEFE5QsewTO9XuHT2ctUfwEZAK0+r
4yfplqH4lYZrraFCVkjPU1l13I17NqXJCIXcYacuh6RXzQYddBshTzEauKhtSk3u
E9MaD3ClMKpwUkqHgDB7ABL0T66gZwoK435L29vpYxpTE0mprsv3YETYZNWKn0VF
aSwjzi62ah7T6qOpGzgExWt5lroaeoWjHWkMEt/lGPhruZDK5SkuNel+MVOmoSPy
2TQLTqgtmoqy8yqeQ+3SApn3M2e6w45EeVCukP3G1QGWJxk7ZIAV8BA7K+hRI5DX
j468UEjam8NammNpSYyQQgjh//CNqiUxLlGlPHKkTl+2c5uKH+Z9Jb1t9RGdmN/f
LeLCmbZn6LrK4iSL3wrftchZyEVgAjUNIglV3kjoO1chVkeksCaOrSSquPEqyxnJ
Q4pF21sZp1jPk/nOvE2WID7gkW3nQFz/0cptm9FWZf9zAk06LNdY5yQCSshJvqVs
xCXEH/sr9hJuEE85oxKxxgc4OQjrzJsiSDkcOxN+VvK6oeb6t/KFkwKAzzImmXIR
9GQ3D66y5xK0uhZNc99s4k+6KFK/06QMZkPp/zO9lhw+1iNNGgV7dPIz/T/b+dA0
tZz6bd2G8mB3L+9KEH2uIxEzV5uLr6t7CmIimhfTvWORYWtkBpMQwjAyHB6vG60S
RP7rp6KsDlUM5TMt0iipTNhr7nXKp2Y4Z/nWfHRayS0TlW1AboawSuCpJ8by2Byr
ULL614ciHXR6FG2Fr8OgKq3Nv/uB2/YjFTboUW4yG3JV3mMIQEJv9ntyz9wE/HRN
zSV/b2V6clfQn6rjAvlzLH4qi2zNon0wUN9F3njoQZiyWZoYLwkSiWwTrCx1ek3o
fM98RnMKvgNzAF8dsIKvQnBzwoWR0RosqzWRm24N4ZtM423rtj22npGN2x0tnf9X
6+ckb2x6765KaGWU5Raxkg6bVTAboeO9DfM4AD8Wy3780wpbZtvn29BGck9aWeKW
tjYnIzsksqI5mcZnCLPzHArtk7JNQFdzEQVgHlGQsNBew4ym+aYs/t/doWSdBbv4
NcmHRFhlGPNAltoHA6tCkiODAml3ur6tH4bx3tr7Ij5yN7HS9OtpuVqEdLbtxfW6
m0IN+W/W5ZxNfKhSm/ofcK7JAi9lfYiLD6gSKr0hhrvwhi4kWyNFlGPFTaqrVZ1u
lcqq1EKAcmZWVt2lKLlUZj6hxa3D2es7feM6PUIMeUIqxeKP734ChogtuRARAIK+
nQlXDZNccuiOWOYOaHCWSoxflrDaqRpDnSyDmPx1fqU0e3SE9uhuY+9Jf4i7Kj9Y
GiZA2eQu/Gm1KT2WwHZoN5/0DqSQCkyoov8yo1cuDdraUu/afgg9Q6PfzKLhCxCB
iOgZyQzPqEgtjo7DTf9itwKNBouk0C7SxpnwJ832anLUMh7d6ZkRAiiY1VyUHrQJ
yun51+GZfFmPGIZTmqMbNMplVXuZCSGd0qH5V6Tq4uZW0WWFvogQMHQAktc/bguY
UqpPAHngOZD5USPOagEibUrOR5s+4MPexQSI7Zx+YKz+nXjoG0SrQ2boZjVo7g+u
k7NgyanTDkWv4eEtTac4y2S2MU7xpAU6dD04xrwxRq11EnHiYf2p2RJ5XdfCt7pK
nM/3/nagD4Pn0m1bDL8r3vYMKQcfOS8DaM41vW9Skjj5Gur3WvC6Tod1MQ7JNoNH
V7ePeeAJ2GaLMxlQ1VZshMTnrVXTMpHs45upX9pV6LBm/F4Ql2E72gk2Y4PBXOI8
pIXXREaG9QoxNE37yyCj3OAPOQsj9VDy9ZGLO4cuJRSx+aH4kFUFF5XgbiTjlXBE
MxSrU99TwWsqWLk57yKqt0TLI5FApresueW8HzuB8MvczG9toBGYpZjh602lFo+j
YSWSncIGPqGaQ/ic92nMPAZlrn1FGx/UFBsoWw1wCWuKpXL4lY9Yu1FJaBJYX90B
GOcarrdQ0KOt9KEmjTsncmdDyQXiswAIR0X4TU604P1EUV4NpUT/edOVE1J/GCGU
0JzrU8KreqH9BTa1Q/9zLpeGKqop6zn9pPNS1pX6V14gKxhrDOKchnJzgWjUsA5a
ii2s2E4rkSE7vo4taKNT+I3FFcdTJevnkht+5QkayZUlI7OaiR1YtslXTeFLeVEj
2lsqM8uu0dX63xTE/4DaQTJLR8gSg60O9K/wR9y3g8zqwt3GfNZ9ndxq92IQTLA5
YA8gV0+Bj8ShckIjHU0+N4kIaLRZdbNpjF8Mbm4ZDILyoLFNR/9GqbtkGO17lqLM
kTeEFxlyfsJKuhwbfjemE8IeYNAllN1Ts1cKc5285K9DnrOWVHG4UXneErIYSC1i
xbABDdFRh26NirRPLLasmCRrynjn2bwvU8sSwEvfG669KZnQ0fOMlllb0z2a7Feo
nvnS5gjblYOOQmnEl0ZQ+MZyPGfFBUvOTLhNihH2ZJ3FQU3+fzYTBTt/RyBlZFkZ
GhAIZUeRCklqttDT2EGVw6zF0U349MjlQ/qgxDggtMK3K3ofACP4TxIMUyofNIcS
oqXsnOl/qsrzSagNChOpdyVPAUGI6vlNUPyedKW0GYKuF61ozHp+YRhRyiYFA/oy
OLsUAdDVqQ3DmMQ+GDHQfDdmgpPzsZfXtGf173s+ne+6KeL70eNSqB2julaTFoc7
TDkd7/FOP42Q5Kd446RXoefkbb3p2f3I0ELniJiw2pRviqdqIakp5260cxZLKNbe
BnSanwCwVEu8/G0o/KjrFzDS/R5+VBDVieOblT0N/vMBVnBflN1DlekusH46XtuX
C3Jyd3jyoBIdlaEU0q6DB3C9qghUz6KEJu2SPm17mnH0ds9OUvLMZO/PqwkEgGCt
m/rkTHFOOxqRlAL/gvLmq/K3vZzpMBJioAHBoywel1YtoEPdc5I48KuKQT1IKAPY
sX7rwliui/uSAVckizxUGXs4wKD2/PmwXLwaTU9EUngrJathZtVjMqwuAvgVda2c
2IgXypKCAtwquoID0O6KF6rHjSbxyTP88sZ5SQvGPYxO4oVVyR/+b6XVzvGGEcT/
sTrUtZ9vftVHRpiResdqdbqqAbHQ5E+bh5raIGV4ImaZH3lKgnUGEeTn20FwX6v2
7tzTG6xKhH9Xe4uyVpqUvfVYNjLQpBfbt3Kb24LdEGDWlt4xCu3iRjnus75Xn6lW
VNgPbohmDrUVS29VVlBSsn8Bf1TQd27PlSRYQ1/7E/Q8ByyjA1mzv/1xc1zBliiR
4Liu4RFhlEWeFWeHJN89givmgKQuzdGvaUNQNFRHU1ZOb9BEn1G/FwSByBuMkSiq
KbLq7qvkQVC2FVQH2jXC0d8fWKi1lYfNo3sEliW/+uFcPBVbaclZiVcnt0RNymkF
r1wf6WJRK+1/CRfCsL2Jh0ZkYhSdSzs4l56/ADd2t1Jy1mc/d489B/Inx9F2wKbA
zF4W5CBl4MJ7kiMOQLH+qvPpqTA9D7m4GGlLws1YNWD44qFPSgiOW0PVMZpSQEyD
lcJ4qrXMr8CcSJ3xYU4Uul67M271BrOv4VyPpBHFpCp6ACO6+keHld0DjydkSMsW
/cREDsdXoXfNdOMn4Oam9BQZ3tZq7TJNKXKyluz6pYRjeSQn88TsUEdpmfXWpjD1
fZjplVQlRmclwftUbpjhDEu60tMnnngrIDJAXfbiwOcKqi1nb+I/xwfGrZd255C9
DFTMxvwq0MbSvkjluynoOs0iR0mB4LYFp+uQfY006i9Ei+3VKxLDkmUWHQwbS5DU
wJqpuJSbzracSMK8KAqXoQOEc2lGKyChqv8W9ad2Yczb+AGefOeinZj03tq0UcQo
FxP8kgkkPp48oF/h1PLuj7f3P+cej+xUIPCY+p/gX6rx/7Jj70tI7u/Uh3IQW/Fb
sMssY4478gml1Nb84x7X3dBqvEnw0iE6phrisipJsB1HjdmGDHBVG/jLgalSMz1y
51dSiounCIsC9E1a1wjYifQ9bkk9nm2qOyAzNMv05f9FbkCMjPZ/cJIVlg/Hs/Ui
ARmr0E01kaPZtyxgRixt6JmD7oo5GiUan1URlXz02/hblxXvDj6Xoc/dWDIGuQXz
rtPDZ4ddiXyVF/Xs6MBkeQG4owLplKbjtbQN9gyLinDUTPk2NtQEPjgdH+HW2Uwt
t4btXgL7UjSOnhtZiV9iFvrK6rLYH0YZXUNw1q4JY3ZUopFvSCVH8os2SxMs6j8S
Ic9CpPDqU833xKEnJtXla6Edy4P6JOQN6NrGGVjRxNskYf5VbybSmHDV4G6Iic7n
tK1aeLajlG/nSETgcOYCoZF1nej9fS3BASmxe2o4Y3j0JyUf+Ddh5cVGEpLeWwxH
q4XPUO/2YQcE8q02zPSwWxeEqeWhEUTPa3LmKX4si5CSnSNn3xe9ZZTnQseZb7qA
2RtDKhLjozlDgutIZt4DGJJuqQjbcc+3wwdy21/qORNSYTcYe0PIEq1j03zBqiuL
6w+vaOlNM89BH+00NYvf32Pw8zHRlxr9gwUdQ8AG4n7jX0Dnvw4Q/WMGCDpIc3Qi
SUFOchR5lZL0G8RMxqXigPIcePayqpNrkgsavwIA9v62XNi5ud6V+EDfHP1wPEI3
pQzERIO26PxO9T93674U8bNxY1YOwr07/H2d/GkdiS0UkD3r+o4eE9dh5wO5G4E8
Yr01QCuPksBg0fEpsaOLdMRJ2Qz7yzmSN+TLZ5qNbtWunJgGPdCTSziEtS6E26mi
Ti4Wrhbj86RiFCnCq/qMINXRkscTzutnC5PKF9EfCBqJmVzXkOguHKTqKAB4xy/P
WGTxxaNhnTZS37M1Pp+b4I5TJo9jHmH10foVS07ow2c76T8qL2gEYeZoP+NN3TZS
Z6AdqWq3XqwCbnLBEXggumMyRFhmW46/PV/B90Y6p5jN0zOoutMX1ZdPPG9NIEZN
3FweeruHEOHP9eG9pgYs8qsw9/B1PyAUiOAdfQeobNI1E6gBVnAcTBJXO8vz3nxZ
tTxSXpBsBEujRbPfRzYqr2WQLSATpN5TI752wOsZpUahT2045/iyIHzlgR2UdD1P
7txjZN7i92FcDJQ+72/6i+j+LsLlqX6c1Ai3ywaR/9ZCkiACtDQn3IJ8NofruyLD
wTpzT6zNGzIjgIfvhts6ZMu6gD2aBceM8Kn6Xf0IzUIFQloJkzxzK/yzzmrbx/ph
P/SbHriaa62g10IESd6R2pN6RlMzUJh2J22GjBnoGoiTDAOQhTVBqNn4F4Dvl9g4
KLbQd+ehQ0BsTVblOhB4skV5SuK/gd+AWyGSIvgvs38jsBizKVy/EPSHtTR7xptT
B66hs2aWMgLob5EC7j0rAeGehzsQF07YX7jp7bZtn1d+v/kMW7s3PWmD4AMio1kb
kCS7XHJ+6BHWEBPEUnmeADhqGgsSjw9X7spa4NR1pqEh6UMXi+0MQWxxkLLPXOwm
lybjh3iHGfh5i+7/+4ngftplvU5ho0vlFkijBvOXpLU+OckuuMPLZswqX4E079Q+
IMCuA16c0k+hwdyhc/J78Zi8Xo9h8A7PReZFEPlF6s78swcmK9k4bTZkLJUgeSP8
/dSmkaVzdCA0v666EldNtxw6JO4elnxU75IJ9d2/f6U2oy1VwgTTsysK3xFamx2I
5gTVvSMkspUYwSRy/mQyXM911OMQ+SR8WnchtQTv1BM/yz3JsoIx5MqKGE4df0TA
OMwwYwihyVf4oitj8ioHHRNGnvKskcugvvc/fxk+y740EGCCe9bw1b3l6c8gMcE3
cDakZOyRXlRsxTgGJOknUpTGVy5uwCKVTdGU9GFn+z7SVo3fMF+QCJh+IgxQ3FJu
ld4WK0mtiCaC+8cU2kZmwpJPDOCgMsweYZdwQX7mc7/psaPvZCvvgqeBDYA96SMQ
h8YmtKd10eQsDo3N76CzVx5ttu0w7hGWmqSMcANotkzvvxTS1EZ8NlPl5UbwS6l7
UZUcSK80IV1fgRQWS58s8UGACd/O4a3LVBzumNOey1RhGNJI6nD8QY890pv1MIDV
AK+fnTTmZJqiflwXjPwCUv0mfw10lzc6CEGmjblqmlKi8h/dBZ3P+VE3O5PGUILe
V4B2/4GkOBCfF/PsZwmwROKp4+FI6MynID2in59QcohKpzjg12bsjLFswRDFpABU
F01IDbl4PbzJy6LrdYMdttpkK4Gm5crpSaQ+D42cCLo/UXiR2ad0ouVuDSrnNyxx
ASQOMO4hHJXbyIqK6QBCG/JZdKRxqpZyH/SsUPSpZJLSuw/zbNhUsJ+ZXIrgjYHW
nxbLnNsMgeLkoShBeySgCfrlHARWhsesG9IYV04y76bofrtBRtQl7nB6I2MGz5sJ
DIpJNbBTJrSLPcz31Oj6wY6Wwu2P2pK1+fJ/Bp4R+aKCThuS4A+pMyg7HNytrEZc
KRxCZi4nzdWPAiSkG1Av38ybTj9te/GOMBjiIOULai4k2EruqZP0TJGTGzdeMnBM
fJxXgQ/5Q1iPTmqXSyvok3PaGpMco++ljtZwlHYflivI2Limmfcp2cX/MjpWGDRw
dybuGe6w/tkMN2+AGqe9zvbRDOPrS7lpVAhU0L0mfV41JfF3SFnE+CcV0OcfHXI0
VltpIhXfuRcDWLxa/lGf4oomgBShKf8P9oM6PePFIfMhqytymN9Car72o8omuwF+
He95kUVBMT4+fMwSxa8WGn2b6VvlLaTi14yeoygXy8e6hCXlEmfjixGlJ1t65GUN
+rRmoBZ4qeNUMhczxNjdxbSiuUV5DctTS4hsRMApqLpD2RfUbTQPDFWYQTcxL83P
7bgzk8Til05rriJRm7DlUXAH6Yyz5pKwXMyKnX8p9B8gx4YpKfxpAu5ViluBwOzr
Krwv4oJ4/2wz3Ewk1Uc2Jc9Mfy+vuQBCRYtNvsOrFw0KsvX84WoNTd+pba0YcHnE
zB3nTBkR1Ou/p6CH/QNFT7nmlsHQFk7xElBzHybc7qNe/dg4EPqQJ7zS/B2gpwH8
rjr9w0iSJEWCu8kx9fSb90oOeNaYgMgJOM3TEstT1yD7sMOSQnmm0eZgKwjfIlsS
lzzmYvvgb3KsmAaBrlHO9kLfPP2r4aRjld5y5dKdA9X4noMJ3Jnm00vi6yV6YBOm
pLNcVUJ3eKT7RiDHks3Yulq2tD88WcKyP9fi4Ag1+WHWQ6eA5vERIqxxlRqCRDND
uvQMNxXP6rv43BgRBRhV6W0zHiHUmGymo3DSvPeKTDT0odkGR59x0EHfwMzLLQEH
wDEOjqdSJdJI0NTZKq8eAUHnxXUAi7AX8YXw5eirMXnb60/IWE3PEJ51WqWaBPkc
FsbPEsAqhvG0mqej+j6ykPuVjtooBLI3YYG1xOqFnKn8PW/tIMqDd1Dwe0CVlLYx
d7kd47dLkRG2GyLs4KcAME2OwK4+u9vkVYrCJQx6MVfajeQjfRVjwEDod4Q+Ybk3
lWyhDgBJG/y3tBv+PkBbYZs06dcgmC7xnxU3JASKnEfx+ujFq7cUCEpD09AQ68cU
DIXYisLZszJFNBB59Uk/ECrMl/rI5o7NQSrvjA/sFiVXJUfP3Y/SEM/Slme1cBTI
8HmMdOvhB2reEphqnKGUkppFcCt40d0sEL6PEYOw6R0zLuX86Y0q+aXJxOh+HMPA
SmaX8q4xcRwlnRyEide+WMw4iKKfjsI9IeDC0TFa7bLzq8BZGuooF5SXd6vMKS2d
rt7ssL2YLUk8c/bATnihjU4iEKwa17whRuiqn21Ls7//Nx3DBWxM5CAfCU0erWDa
Ok653uCTyP5CJNzM7tqdh09MW9/O289dUfvE/W3c9rRs15jPua7KqPJXtw/pNHU9
qxB5h0svc0EnmeiTOkMXNmcD/Yo/rtcPHzuFZn7ZV61ByQMeuREYeFkREouXDBaY
qhk2R4igwqqondYVY29zcnOsGulQGLpLZlcwyYG6uLMGsE2WUjCMRtLf8zK6sPD/
CSxR15XYrIhhiTesB3+DOJd7qb99WOCqU2fPr2tsZL/F4kwaDQE5RHhaSU7uAzsj
FxMFg464fb3I4MD4nwAOhMN1Eq5A/4gtC8cv/D5HOPo5nYyikdN8slbUS7SBgwcv
bIdJEBTD0uIDQSec8XnmZmVJ+eEVateP0XBvmUlqPp6KdLOQmr3xBl6uuybC8z5i
tum5u+ZZ5ntD0Zd2Xe8Al+vvJW0Plkjz4yPAmRj8e6UhIOOpS/B94EXAstVJNISN
+BNfhpPR8yfl3FLR2Gdk0Li8SLWpQHJux0x0vX5HaE6SOs6GKUlLG0HYeuqsQG8f
xTQCL00rR8/ipLSUWPC0V/3/n+hvuxASyj7gouedSI9MnlASqHLrMK6G/B1a++7N
RpuuGb0bRJ9uensieL5ChlK/NQbgZ50x59aiwdODyWdE9k1B+WYFgnUW2GIdWYbf
cywdbbK/WD9AAiAk/pGgktd5Og2K+sj4L8SAV4eWUKdQ0OoyoLvDRHSI/EaN03bv
g1RywfD2yOoAsR0aE86D9ftKotPHZ7qVU2XFMnWi7i8VgiucilhDRQAMv2dOciR9
Y2PtHKJj+d585v+yC3uTTa6XmibjRlVClA+MZXpBe8cgw/eE9rufvRHt+42YZRO9
HtJp42RPgQ7ELsoQrZ5i2xjw/A/3iw7omHNhiJg8vOmBay6iXTrmb1qQ+9ggaKuC
M7MlIDnPdwKjTBclmGH2r3VX6FbjRHooZfv9gUTVGxvA+tzp3pipGUjypSKP+ZoO
CWcnITsaWCTROZEISY2bJNrvfnT12kQAdMFwX/UMSOn2qDsBTr1rYOfdzW+dmhpz
PUe8HLuSU/ZjO0YI+FM3G7uayWFz8ZgwneVXAGuxEAEp8ZxOo80bVPmB/hoPWcSX
5CmUYhM0OUP9VGB7cNDRdTWSF8MrKLhsVgO2eXpUOdXtlSpiOzEfkB2pa1HCnSl7
bIarIYnJPVVUnpVFM3T0J4ppj/ipiD5n/FkQX36la4DT/GyaVLmHS3GSEMWOd3+A
fa+Boagu4uQ/P1EexLHe/tpzw68JUuwP7vYirUKwZbVusQytEEGZesrzzj5VjGY9
Z1VtCXMU3GeWx26cNt9VaO+5TaCC2sGhMtAOO8DIpPCIilN0jRuXsr/sIqhofvFx
wRqYSh9+zfdD0lOyPlUha4xnNBmA1mMLdphRl2vEQ8ckpfflhfX8csHO1LzG86wc
6iCBVvdFvXlm1QooIe0MPigKAB149cewszxyyKpGbWRu+3W8ZXnf7dCNIhZ/5om0
ZeqCccXSN056EN5FJ+LJEeJacDDLOX4DcKHWuhQxSlfOe+5U+JptauB5V3lnjaOd
so8dVHrv7uCsPzp5ICIEvY24cRKb/NZGQ5inUbXsBpl13WViMRUG7hX2ltOve2Y0
sE3G6CtvKqyAYUraJ70O57XFFxl8lyDlJcfGHxQyX4hyYQYLRwQGd6RbnQ3Yse0D
3qawRHix+CKlhM3iJiG0DjrdSfjIsR+eKBUKtchEjjcvI2FG7VC+GETH3xNq+wsy
pwJnX5XpI/2iON+Avaz1RMCAMAuStA0RBnc58IF8ieJJswnLlKrSgglREGW2IErI
ifdTHskwjdeMdfnmS6Wp6+dWro5TjUl0jt0Uc5r0QZBO+0SqhUNf1LZZcBHz+dgj
d7SyF0FzpUD8IZO/7+K3OfETalr1ZAXsGasBKwZTIb7Ts2B/wR2kx1HCCmikhUXa
2lpXrG1ExWbrCwaffkobVgZLWXhyLyAkCj0i56I0f1CJcMX5xdSeRC+CTk9cavcP
SlWVSa3zHl8TrzQ6ln9h/cxpVUDM1tqnf4jGYB4zDRvVQG/AiZ9qKRBRxPfouNnF
PETXMIqaCqgLcR8KTnaSH39FKlG4/P4RrMlvLcMzaKZN5fEZTm295WWvYpvry6bu
CTTdpZeNC1Ok1k9pDEoXI6gK0VEDNozF0RjkYd5N+9ME2voMhkqLS8vHUaP6JOiB
40PpR0nxImEQ6WkRYOxFIEWdkf6Fj6Qm6b1+6uMwNdJh2hXP389y1UWbe2ZQ/iO+
55ymf1+RuI8KvXA8PA9OG69Xm3mRJ9afZiza5LSwb/wd44IrBzFxtsrFHGir8+42
xg8AqxQDij+MrswlENT4X2i45g6E54zp36MV9Df8lzVZX9WCDbGYNzHxSRMuHD/T
DTntWD4fby/vYp8WyxFmwHKL8ZyiMAUDlKQvT2TR7LnjCHBGmUsT86PXmCksDDl9
agiOvGjCGZB05IpsFsWXjLj6kbwkRhdo0/E3657yhotow1DEBwtL6uM1F7Y5yUP5
P/BTtYyaV36jOdH+F4ztn2jHGNxu1XfCkOWyfOMChYbyG0jVsU05M4/LxquLnyxC
9uTijuZUxdr4BWOX0jAyZ+igIA9DgxWaGhpLp7/+u0rDNVmytOpqA40YZj/DDZtv
G+rz2Vb0DZshnt5bJgBkLYz55QV3TtZRfrCCuYLwdFP839qS7MbSiOZDoEnFxW6s
sUJDfOq3Poimh3T2MIW00kgUuUNVzdnjWJW5ZMLDG0a2Tc0IJ8qkew9ImEOQdjAe
Lo2Kzc4VBcZlpbKOiG8tUmxp6KVkIT7b9wJRTRkDwmISv7TYqsakdsKxGuWY6M4g
eF4j0OxP3ivQV4cLRNwLb3pTjzCkwAUjqW8MIo9qFhaCjcUiOGZwbc+dIVsyPDVR
lUKhNR3k0m88gwnNQuMO8FA4VVf5hUFPgWxjEJTJSlIRCiY2Jr2ta9Vl219LHtM6
+C+OfoYUwY5b3/HuWcbBydXLzx35WgmjrY+mXzkn0xbkKecGG45e2SSnR45MZqSL
C3byLUe9jmnAGD575h5BQIqOR3eMp6HEad1g7AKAhtjAhgTLMsXjgAskWZ0JEEnI
ZGZKOgHLJQSIw3V0XPmK3VXjZmSsoA7CrPeFk0ZS3c4558PkABNJO0Hb4r6O6B9Z
rXWl8TAza2dWaIrNyjWmaC8jWEx0dtTkBGSAco5IjqqQ1VMgE9i+KdYYWzFFRUdB
qM16T67HE4fwqoMz3EFd9rTUMgDGaBdLK4kUkQ45MSoZVIQkLBc0YSXVadHEaS8L
l62D1cor4sifGyr15+KI9UjODrwGofPMUKlxe3mToGs2C9XOSLZtfYk3JP04STQl
ubZ1+kk5qJmdqaWf8rIn/R5fI7uJa5BOpdXUntoAKsyHEXqZjo1zCtW/mgl97Uuo
GTNBmww7un0QFekD5r20ED7xAWpk6yKhDcKP1k1q/6PS+T/eVQvxHIljOSpv2ro3
2j64F7mp1vetZWLU55L5QS3BoDWqOLbWFSNpBFVk+srviVRqb00DsF2kYg1W/q7p
TWjWKXiplLyTZ9Zmef3JPh5xfm1e4hqo0JAdMK2148Y9Y4D7fRd+LwBGy+huY6fz
iP0+hQlApbnh9bwqIThydbejYcD8uRHnQ40mwVdVwh4baZyDTBZHxhON2yWu889g
JXo0qTFGQ2LbXs4nGv7ogrsBoj4EnRnB6A8JRh5Bny3g3DdZ79o6kQ7TmtOmC0b6
K4pYkDW0DlA9k1YC4Rqcq07lJb4EA1YfHlscyG1xgHULnG4LTA7sc18vOA0clxVv
sLa/37AOByki5nYacV+wUd8S6nksulW7Mq7Pt62I3gT80u3B7rilm644j8BZTduK
Ax2yjZFHIhDOl90sDffLreDcAcCeNCdqJ9LDOO07SeR0dN2iHKwlYosWaWgtYrnL
hZhjZQMgHAH10TG8MhSSisBCvlv1wJoIIYt6vS74ME4P84k26vg1tSYaIvIUUQel
yqGBJUJ7bwbMdvJutJ82NDNdM0ZuQ33a+Y2oFBBnOIo+sauyg2l779Mkv3OOsSzT
BKIjLV2EQUSeb/3pn5ous8Zk9mGi0uqZjPqFboVtdwcSovhDGqeU3sFw+PawABMt
Es6cSqoF04C3xzZ0glRSTrYcDb9ioxHreal6qYLLeOV2V77yoeoLgU6/ZD5h3gmd
7vOnrQCt6FYoYDsQcaWZYPzqmvp+Zc4p1aiEVxpXM5A6uClHxnZziqO0L6ZTRSZI
VNJUxoSFHOwA3PDvoIroaq+mU1iuBjOw/DzOsXoUOMFYAFxtWhjxyMmY9g1eQX8M
l09jXnBS+nnAVXVy/px77aARL+95tWMNJSBIlNLXqna4fkeU3z/gSnZnfnX2TYaL
NaPKjuAmDJ+SmsRfztLXiAWKcWxl1hbgA3WHXMD44J/1MdWmtrG1P5RS8gHQFBzb
mo6QusG0KAKnR78cZDs7SDVIryo8DbF5aEgoSKywgFf7h51fA6PC0dSoKhK5kCuz
fKMTlXYws74idesgboHN2ic/O1oKxjRedEIq2EXzEMPuHPewMVvYDvC7kXNvKbhe
r6lj9qF71EdVt0CccTRySvQBtE6cejG7527XdiRTpyGo3osBgQMvhGVOIUfgERyr
lAvYjzVqTcorfGostAp6OISJn8CTFRAH30xikTaLD1lPoB+HSE4FoRRgObKTgeEe
speQbWAiNk3vebhkxDJQkyyIPyxQiQGSxs4TFJ1Mptmj20Xn3JfVx0+Hr3Ex3CC1
DUZwjV3k3Q5X+gGfPcH7Bk+c2DEBcOGEL4g3AKMnyJOYWsznd6jdMGmDZkC1iZ71
EMQLYqh2IN4LVWobhX3wzcJX1vTe0ImtiyZ2Mo4LQl9L4QllkydBHeJRRpuAlFwS
LY+ozotAORr1L/DzLMozbwjzq032LzjxYBOk1Q10QR5/eu4AckCIG7VPyZdzfSn+
qANd3uFY6NMT5Ioo0vlW918AWkbms1Zf6Q/GVJiS0LGyaTIHIXLqQNtlakj30uup
/KMy/iCXbDsWrIT2cqT4rVp7wyCzoQrDwOEsd/D/G+Zjn09xB4xRmaK7MrR3KRIy
CECyOty0H771hO1Ex0NJo4J/W/9zsZis8Wuqxaq1/Z7WDBUZFlggeQdpXJBF3LK1
uCIeWu279c267ffStm4igxcOgIWVW8wcR8ri3un6Fgmbv/zkjoHUvfeKa269y5uT
gC4bInLPhdF8BtxW7U8Jgtz/vOxkb27Umyw5/jH1fgCxi6/1HT5gmC81mBREEUkt
93kpU+YBktf2z45z0kGxr5Z7pwPzUjtBdOOcAdSuIrRHC0hrIKircrQam0tH8mhN
kDO8Lmez9zeNvOnJpLH6fF5d3aqoSBXqpZTa0/2LFSSYbxVKC2cz4mGyGg79Wo+D
KxX8eTxHFlvt98HTjVMpj/wHBVLNfEviO3V3Gx2kf1KCQe9cL2XQ1sko45UgYOjN
b7/bYffY47x7oPoAJnLYQuR/7k74NqvP1OLToDCV8oQ4MlOdXsd608M1GHl66sKe
KmccvuXE1j28Rs43IsxoQSf7RDVEVTG+1vRyXFmYgoHwXD6K5o4UtsQiQ0ceUIVA
rWZJ1F/3ylOWeO2HiZSfB5AUAXCObzHlnZ2gEQDagAC1JVovxMLQoMm4FCZeLPeS
Ul2P9L2GBptpcyioPlyOlsGh/GagwJo9b9RWaQ6yLoMU4JqavOuQHuCfMgX97viX
2925ZyogG4+zUn2tp82xUCKXzFOlmaNju9/pofltxnNSVfo1knXFztpzWl/tR2ry
FMlSBvy20jRKK2uGrtjjoObWhvT5QwWcA2xKXhYgBaFYP0AlvHFv/IOBPSAJq+dW
9epAWKtjVwj6j7R3an1fmbOJYR+8AO2RfmC7olrsnWkE1w4jkBs39jFi0vXP/uyy
V2fhsdH7xQwBL6ywZj/SJ3WHnpGmi5QWsOecjk3oHXyKo5OVpFHFQr4h7J9aatcc
KtVLYPLifir3ayUYojKzLDt4knY/ZCoaYedVch+z1TpMcS0v2SWIMKC4YiOyQ2nq
v1vZDsCtjDldSJlUgZZCpfTCpX91oRaXpVRPfqTvEIAaz73Y8YgS+jsJ3yhj7T/e
9xFxaIGPLmdV4i6LICBFKUlfzCjgH/xlqeCUV+0EzxYC6Uvikzvl3vL3l1SNXznM
tuhpLSjAe5ub9+AJR9stCJoi7TUTqwsaZQFwi++zz9QT4MHv6Wfm6RL+kV3gspD0
DiqFDWbIrwOvSIbfhOOjFJG0RMANcTAFu5tMc5JCEEVuE0FY5KiI83DXM/nmSK/9
EuOoeOdK6hmixvTM1id3DPKPZ+TdmKe7xs3vD26juiIQtn/Dgd1CRDxRi79Qqg38
hHs1Tu1vBHVeJlLfOIqrrSnT3yFiQsogZfdqk0J/kG9oCr4BgiuDbFVTZmWIe+Sf
Q2lzMKgL/vmnVil0as4t9ArW4gDbFw7ipT+zJ2av+mtM0djbL9v2Nc026AfzYlVb
uVljkR7seQC0/7/Wk3CRtpHa/keOLhnMc5RI3kk9nDoA3bvezFU8JFkoAiPfUAuM
eZA73uC8QaNZFtkbdsC4743phEHodMDvuHtlOZAYtt+A4UKkuQzI7B/XQeAxvb6b
H8EY4d2skG3z0bGOZRmsWHxqbCzZNBya2Y0l8qKqn/HeEHVVkn1OsiKANUyVu4BU
31dGThxBA2nCxzA7hHhyeF/Wd0v3mqBPDZvav+w6PW3ZjsVAknI0gNsnoPg7ofMH
pFCfq1wUk47yKbOcKwAaxFCv6AKkMrMHMvTX+C3JHR6HoQ/49Fj0kemHbqXa98li
VS/hgpv6E/twXQqkCY9e01GV7ygieAe2E8VOYyKRl2MeP3IzTmpoBwau5sYgVJ+D
Yw13KD2Az1G0lKBPAMj5idqXSexUORNcix2ObKSl3r/S9Q9IbLY85f5W2aljzlF3
h8UnbgAXqxFq/AhuGfD5ysxtHHdiYln6XqIKTddZtcFQcBUA3YxyL082yYJKdG99
j7Gr71HWnU9mdTii4Eyb3NKa7PPeeqjHnN83K1ASAyw/N5Z3jZPWnlaFsXi6ZHgI
rH6BA43IM7oW0762Fl/Xoq54hMDoWP3NMM5xyBw13ydSCYurAo+9qnlC198yJLE7
HsLfj2D2mfBVZg04DMxBdOp7SilgO4Plk2S8W1Nd3D/ld17nq7OGlJFGQ/s3mWpe
Xlzc+NQQ9/GuLSzFf/TKK+PYb0Z+wyWJ4lSSTu4aLBp0UDSDcZJLLQNNLFCHnf5D
ZdTTx1piQTqHTZvLBDAmHA9Kcqt+FzFBqvOoTtWt4lUoq7xipcbfcGJwaeCJnPrw
SbzdKXQ05q7axDHt21z/S6oXOUTK09LkZbMV0mOQifLZ1HjpTSqoR988Z4FUkrx7
5/zOZu0JLXvu1nTYfDJDZDavHQkZdOgKHm8kHxwIlmRidOjUzoNeLsmw2U4SX5ea
V+2NwiEFqZgWqhz9fJCPZfxsDyi4eJmNiZ8rvT7P6RoJY/sxKAfzzMZHqTUEyCtc
oLny1a+9Es8gUUteA22ULNgHgyOkK3PLrV/gsV5kYzm+BlwQcy9KIv5dL6jDAf+Y
khPupvYF/8X0o3EIOSD3gs9mSmPzGHfNcGKQn4spqP8CDm/+CsHJ+F7xwkyv4NZc
lDRuJFA1P3yQajsj46gOn06L+Bptx4CLGeMPM8Jf5mm+cbSRtYlCOea4linSwvlY
S4EfRtxt8PDeYW4XRnkYEc/0VtcxPz7TEYi62WtdzjoO5LNVU7hahvizDG2Pm+zT
P8x1wuJDVcgFIFvNCv/8Y7lXzPFbGUwcc9c+BQlsjz4hX5/AR2xMVCUInEzM8l3y
LzoDGwoW5xQ075oPFWXapKpmzEchVHOnEQbSDeJdqSILbkujOe5vHRKBfCDk0fag
HKHXeX/x6DEXGiit6MS1v4LIR4KYXm+w4l8+MD17ZnG3Dz0gn9tJAW1E5Ww9o/5O
bnbaOv2fQohIO6yaesH3yRO1hcoPP+xYOw+5tz0HwFAui5nVS1hFiF98ghe9fb+2
sqCi7W6tfU5ImNaO79V9l9H6vrdkv7vB/sI6HZB2CGr6BGobqlzB/MDyHSjpG2Yc
mucPLKZfXpZfIsjo0YSdHzgcp5QzaLgbNDMtIT1aO0eV8L3zinX3SUIR9oawuXTb
PCxqSU2QYNjELI76TUVSKQq25RS4bcJ9V3BRL97pqSlwGXyPu85xUR9UbmGtGufw
ZVCeU/QwEkjocTkS/TQsdMzdg7yRjWlRqFllII0/ibFiKbusrYr/qPjsdqpzx/w7
uZP4kw4FYJjPE0dyqL54JPtPY9/pXHZQWOcLl50q2X3NODEse5wLEz9xYg5ecCVV
16+31pJZtfTPk1eCEG+wUix1tIJM1DmmFiqqriXG7rgq88NnhtZCaKbKTyzOlFNp
YZdgYQw8TPpHAYOVO7bknyAbHYVX6t6aDg8m9V9eQp3Xsv6kPH13htainICVqXYf
neraQ+LQZWJbsLlEqWrDh9hu9Np7nmuIiPoEJGB3nJrRMidC/8snvR/zfW7+bsCQ
XEw2esHgdPCfJJBkS2lc/Iu5HZNNiLnH5x4Oe2dBVZ/XVf7jHqud0faGob3f0QwG
Yd7EB3HVZzrQCJW4Riar+3k9VfhF+bVUI4QbcL8Z8aN7VD0dBqf70EQ1ULK7Q7QD
Rm078X0aSv7NLcjxzZcNS+Fqe/HWWnJy8PJqijty0tCsO4xBbiI/0+ZZ3y/Cmy5f
BXj8QW2i3wd7SyxZCAqJY36Ob4EkDSvUzvgOY5a5grZVtkeFe+At8uHJ9PAu7qtE
XKZJife2X1LKX2T3IN5fSXVXieyGW2+K0sM0v7VOYHd2/wdkTbsE/0UhtDDuMJ4b
kc8Gv1hK4Kav/UxRrWu6rPPp3AsZDbW1k6tpa0seYH5A7atRjDoEWRc6msoGyenB
IUB5YrhFS6OD/pr0F0PSSworm/Fh59iRncZrLU55x2WgLfWpqNTytWYzq51Sqsq8
Wu0GpLscbN6FyF9YhU6jEhrNJ8azsmfkrtlZteBDybnxLOOURrLuEeR0oYU9Q3bw
DD8Ob/rmQBVXyDFkpuNKMMP1nSoqMS29fjQ2dX+OH8F+y2OMRc5vrtlcpH1i6fz0
poj8Q674Ob8t9KeBjeBCuvE3Mib8qq16KQkiwnM/snMiMH3RnaFFB49e3paFGoa7
B/1+/ay+fniReBFT3UvKltW8f4QkE66Qv3XmHY/BJW9MfqyfLZDAJeM8Y1mF91F0
4l9WSvkvJwI8Jjfqo6eqhDNhBF+ZqiKO7iHgAl+Lh364ycKk34+JKcf3gW1OSl9Q
nBXzStzISqxpVyXr/+r8Cy2S9KIDgGx4Djeib4yg0HetCFOgBEIlxPsSIYwMNcra
HQC6BXsEZvbMoxxpiQ4cmUlcFz0/PgOhNDIFvlpWFGEUkgViQ/1SPawVtNkcIYY/
ZjHgx7iNYuIBplCMSue5hhZ6/poKg+E5ha7BSQYWGwg6rK8piasf2xXRJnW++Djl
MWt6PWX8Jgbo+ec56ucSsx54NyBUN5mfLJFRjiwQBC3I9iy7NbVAy5feGtN9YUFw
oc1MBaVwvGXyLZmCrey80TwjaLqFZH9e+UQWkhbPQPkOob7tTFpq0An1Lvcfgvhm
GepoAyXfAe0WZuqwdnemZpNvXDA+OZMJmIKf0pHY1C//UfJu8gSvGWDUMYscVsUS
Vh0QKlgnoR/cOkSj+cbKayHjUVXccmZEYJHXkkOBMKMqFg8SwQUOtBB2/ru2AuJo
3a1kZiwfPUTDzndDQEzpzhKk2hKT2oTEaWCOykJsvRF5bY5VUsC9HNcZf2aNt51p
XBOMjosxxp7S+ClFAfcoqW1K2ofE+nLDVOxG2qBqZAqNm8vfmiEqoFt5KJQtGqZo
LFdiX2ao0hDFGWWgZ12V7n9bjpUZ5Fm6BF6ecqXDbaBHneSal6sXavuN+OtcEe8h
daFIeUT/NEsibIp8fCJNRrCI6PeCiNsyOcRM0Dz4srXdetTmOOk2jpD7rsZxxkMb
uDKsyfKtT9xXinHCKOHBS1g17MqRy6tyJm7k8p+0UbG6VUtlwKReERGHPMeKPIIV
U1qGYsXqf6BJbOhAxq52BclxAc5d6dvjMOuJpL3FQRiTbAnuMmN1JJOFOZgmFxSI
/1Wm5iW4bByyFOEGDDMi6wcxhTiXkFXd0qzMTQX5mXezooUExL3alhNGV52vzHwv
1HLg49T29sahvZs8o7lPCcvISM+Qy397Zi2ZrztREdERJAR3nZWb1T9MvKSVRBV2
JwSUHJnQbJrWnXYl5H7zi95Psjv9yFgHE6KGHi6X0L0EhatqQ5BFNUr5ankFwXzR
bhyVpPgDc+cuDfwYV5pwfQFtSluO4KKJ2H43S4efcsBgSGLoCnnEJKQ0+omv0W8x
+AtklhbrV3/SuWyXsytXsDfFztO6/Rwz3jnIar1Sy8M55ByJ2APWZRU0QHExdBbx
HzqklNz8wU8Fne6TngWHquX3rn+icsevocRE2WBfttTc9BTSIetM2YBVtxMBFR4m
6pwu3HAuaguDMhUMrbEsmKZqaKOHReUgcpbzDuXwtAZWSnfi8EU0vULIzHkhM5po
VxxoIejWmTmRhXHKgigt/RXMPvobLV4i9XlUYy7fheYYl0Pp1QaUKy4JbWYzxKGM
Gei+/YTtBt0gM1PlJHCPNSJGk2k8EWqFQbEhlGPbWrsQBLz59XuGmyKoVfrv+wS2
2tb1HnBVrDvneAFu34cnPFq8WjpOUkdkKNjtWAUPY39I0Ao2w59gz5R87txSPchk
F4VaJ3OVkgu++o506rOJwLCpSHahn9EKdSDpSGF0QAPJoyj48C1pIELaGI++R7v/
AnK/genjdToMlz85KpZNi7jQ2GlXHM2fzOBW6jp+E/lBOFq/Os+8PRvnTo9GqR1D
0HsG/VSILzgjWXr2i9CZn9Lhs/wU3dzLtT6uOwD+dPCz4WOYonUIoN/vpaqXE1wb
tdl+p/pM8u2/fwwWmkcqaCc0TVL2AQI3N0N1RYYg0aV6D65C5BqV750c2cZhD7yj
vSO6wcWflreM9u5Hb+W+obYEcWtBXPeFiMTZoZJk2p55j06Rv/ce+ibENZVqplCj
2X/RPZbCYEF89dBUB1nPQtA4XCmDEKRyx+om2qZe3Uu8PoJ++TmVXqzLrJCIz9xy
tF3s3iBlvHY1c0V8iayEa2smaKUdu8lgSfqYLiwzPdi1TuKegmfKS/k9k68WN/nr
lK0nYdE5ZPPN3yJ00Ah32+f8RXLSba4xMieX+LTwuPa2eXfYI956mwqjq06MrbbJ
JTtUFedDLxG4zWLECDGzOvK68YbjICHcwp2oDxXdZrKP9R7UuFcn+obC8BMPNHKF
J4eDNesdT7TLVt6nZl/yf2dA8j2I6oO8Y6/oUgAsNsoIookDHLavPSukr13JZlDd
jMi+ZVGsdUHBE4Iznm/plG2yCCPZgb5XguFdrXAKjGpie4D41Q+xCR0G3eCNdcey
iQ4+IHRgUZQt8J2O/gzgnbsK4owZjx/59tA6f4VJwIVNRdhxw/NC53wkr84WM4h7
ve2m1/arbMF0xKzkV+OY6KkyjsbsQzOQsri2JHLtjW9QkRw0d7iJEhYy2lKldLzT
Ezy2/8adzkh/TF3qstyYYD27ug+KULpDScmniFwvOQETTu9PNAF7kmJ9n04Bhgm1
3kqo7aHhh2aYvy1gyEHKxzzonqaY1KlA1RQTVf35/38Fl8M2HiUHZwIGPNWDgFdJ
WiYQnUqZuZR4e8yt7b+prxEgOaaJ1ek5DsQt3ejC4PHxATVQEJdpOqynpg311QLl
K1dhdQqmHB2omZCzeT2dMAX47xN1cyraXhnXvMDCmSPxlsBV7m6Xw2upMA34meJ/
Mx41hCL4ahRdUy1Jq7xMvQ3vBVtjdsCRWKUFIYVHuYXH3pbqzlwr3gwXTMneFp6X
UPpmzxv0eNoybJKlaH/YgtJEvlgWinOxGK5S4IASY9OI1U9VaIWnRcH5/QcWyG4/
Q8J92falt0XR1vE09HD9q8J9M2JKkrRxjQ2exZraFBotAz+mXL9FjRk5VRcsPh9W
6M21pBnqsuKprWY/bWhNYKaLf7cdOp3auFFGyZBT4dQvZK+T8TZWi9K0qpduxIx5
HpsqLLra3Foqvti5uaEdWrBLQ9WZ4lKkqO5vfbgqqUsXNZdcPZZkITAxlxd8iyK1
e7TfiNS/3bi27/yoiEm4jiOUN6bcFVLuETiUT3CPLnw7HZs83Bn0nayNRHTmkZEa
mOnXFLu5NprPP7HX8Z3iw69TzN2wOdg6z8riyAo8WAdmr+M1OvmzGcUgmUncMRFv
axuvQdtmMvi9/ss/zXaptEioZ6FtbjZaKbl44kqYaN/2pPB0h601jRoOkzlmSuTB
zsMIBN/njc2a0uyiPrfJh46ab7kQEIjp6dBjReP/QKRrAN4qaHDCT+fU/FH/0Pid
ebPtgr3+nMrcr/LIDKL5CjW5kB9VXDoEek0KzjYRnW7SZOka/8nVxvdZUHeFn+sI
COw/4hlsspttCbCXpAX/7voPTnqta3rVnhAelW+dYUWNTVibp+kLMQ5LPEgLbQ4H
LHmADfsUcKxKswN2ka+dIg4wWOrr5VcPjoTpG267ZNFuSBU94YglZoxxDPDTcPvv
yH2AtPd5T4TeRLdmjE0wpGc/WPqe89xGT/AfJrfpH3NpO+ChXYZs1QKp526crPiX
JZIqEpfrnStexvEva3+nH4F9p0u8/WW80FHYfaogsAb3WQHfyTPCShv2I17BWXOy
AN6psUX3JUfiXtAEHoXa1J8oBLllnYXImzCkw3xAwbsfoeQGN5w4h0rBPIBAj8Up
2gRW3hKnSz2Gl5WbTsHYi2wJARmGj64DUQL+ioq5lPzGIJwF4BgAPvrKiHr+r+u+
y0iL5c2AjVuy3dgKM40xn2Q1vVuvbYG81/i/hUMglhe4zZFyoieB/ir22KneBpVB
JwpJVXOvV1l/nMS+2w00nbxk+u6BXSz37z97OvquXByHTPewiih4Z+5IiTV9QIms
07YQsJQ9lNhRBi0CL3Gxlq1H3esRHj6anBYkAYTdXNRplZZXSWY+6dA0kfl4eSWv
g/McD46dS/Fv5rIjjyhrlC5hN/r6Ely0TBs7QtywMjPqa885d2lVDTIoVBUEv6kf
j982PlDRsHUGGzx8P+VlwRDa14jr2EI3nNOnFYjSlmGoYIC4Grz/5tCo9DiVCaxN
QFUsHeqIIKspnffN6OTfBlH+CIlYIYZ28dtsI3ngervkUlDvUzH/kLRagUnJ4JGN
BvP9opPMQCxt+SR4mcc9Grzq4c8WoyGFa2lwjPHaTWClblWJ4d/r0YupAjJy/7Mp
5QMFsRzlwlCjD7QB/8gJgrTjP63EYCFZKFA9eXETC55Ozr7jYTBsMkNgiy4CXQcI
QlVIcE9SFooMNc9fkKkB19JG+ADLWbIwT60/mD/ElnMdVv1TBrb9J8HBeuG3sJHD
4UJB3ZrsNWZRXeJrFPlpmYibwnXozbcGyxgvZrX3iYdnkvyIDX9lM+AIUoh/aRzi
1uQCzy2mngC+8Z/BtfsS0KmPU9rq0lRQ4Ja2Xfi9QjXgY8PcxGcM9Dzf4ZCYbtOt
A0RpCafVqgB/N8s2uStm6ICS4TdfWP9Qc+E3V/GZHdj9WunADgSmA0ZEdUEWt7oq
q+LvttaSogCULpZNk8Jdu/M12CaAuY1jqi803PFzZXKtiP8adTVBf4mWOumdikY3
XaNRQqYEE0S52PTabvyF1C3WrhDCHBv45CxBVxatacYexpAHxXqC+hUzG4fqcJ60
Mqtm03ffSiNH9Rh0biZ5lqVEdozKtnbIFlkpvlVw/h04iToWTNNBUapmYtB4XDdF
80tCUsvuYOfWHnQzOBxfxVlGQiwoVvLzhMG5s46FMuMOa1mHhdf7pIfaAOZTMkiR
ZTVN3zxcSZOeu/hdiKib1DAIxZHJ/jCAU3hOu35UhZAJYsaXNUJsS7wI+Y8XF2Ov
1fTr1aDI10fPARZl+nbyWLYONOPqjapy/bt+pyxnEuCTP1vpIGwe4ish3yacGLLX
iyfM5/NpNxSpakQsfptuKfuz5IJ+KuQ2wX0B4BhCbPysONYIkX38PSbutqpBgczQ
At0ir+h3uCA77HhwexC7pDuQWNh8LMu952UhVAklBetRHHSk0EzEJMHsE0N+1eWY
Go+fKkTTj0GK6ikn7fS9r8028mBn0FhiaWWL9cN74PIgUslJTj27/3ejcAz6u2zN
jCq8F8gErI3bectZAt7p/cjNC682ZxGdlgsrsx0Zh287wEa2H7do1MkC5Qx70Tno
IuX7ZWnKhzMDazSACa+TGRAb6mZJyKOsNKQ/bmrh98fTuRW8vc9tsx1wMrOfVf6v
ucHa2bhH1sFOWkRHURFQwRHhaF3YC/LzSMZZQw20kIpsB+/nhDNLDRszrYX4EpQT
I9bH0SN6eYekSrgxV5btxYh3NvvXn64bPgyb1Vv59ylNAG+JiV5Kim3sT/L0qvKg
mNRVTVkf3FwnAyHqnmDGEQq0h4du3IFdkJi03YPZwoER54+KowoPDZcFlFKVvO1r
LqgCjxhxWFIPQsP8MISetcNxT/zgO390YJKfojphfxX13y78Xu0BDIi8tEYX9PFF
mLxbeNufRaQM1er5lM9aDk3Ezbufy/L0KEuJCsiPTkFZTUAGj1QSOUAXevgdpTPp
Hjrc2sYSvxdmG/N82J/GVtsVHO500KFD2GJfIhSBg1neETo+wlVBrV0SJGzuNcRr
ggpdsz5nB6kDX1AE3Y96wdP1ReZa8NTaCX0Vqo5BaeVZAsJDtEIPQ5fmqKKLyO+I
x/BQMwoRArgVP+v0W3GnlIwwTivZy1V5BiLVdqcg+4ByrwLVD6Acj0Vr0Nq9N/qc
leoqFauDb7eHejPyBhG+XYTvj42VAUGasrjS1BY5v2czaytqihq7q3SgEz74ViMW
Nh3ZxnKqDn5BLiwcSbA32c2CmCTh4bmRCQSJx/mBE8Hm5aJI/bgeCp+NORnq8qPo
3ePdwJDjHPFOiBSw69jiA2YdZTGTUVAKl1BuWQmtN4Ng/XWYFKckXHKb+jnay6op
6kaxdiVZyZuQBAF9kwnIpuZWTWVc+uepDyW9Fx2FjD66f4OaaP85Gr1D8RC44KMc
ohTd0o2Ie7uCsRi4eR8ohSoAgihJqiEk7mwS6pqm0Y5CUCueJYrRDMLQVBYgCYrU
ugr0ozOmlzz4LZTch4FBLwzWzJ22cxRXhueMyKfR2rok8DCKR68VcVJr1rFR2whL
C9P4Ll0345+fZoo4mTeM1HBY48uFBJ8h8gE0/DgUG3d7SqmvV3AmQ8F8pCgi9mCG
LJ5AeamOEwer/kTYk1tTgqksZt4KFSD8pPhST8GUJTvVGngJQyxWzde2ayrZlEY5
Qh8puc2RAAxu9SZkAH24uFTC4gfxXJ/KngbUVg1rY3XOORrgL/qR0ngLDWTRYadf
IW1rWbzKaN6wT8amJbOQySuQxHyM0+MddXZWilzkqK8+REjE8TcN9zkXariBM6Ym
3WKffXDO2nh2k5yZcuFlViFkeBRGJOEnKC5PdxPuS4qk9Dk2Eje4PLRFIAbxHm1T
WZgxPxAu8nURqM3TjRd2sjKAXtL/D6oJz1ecXmbz6MvXALNM5AUDvslJAXWM3Cus
gzyjYqIQi7M9vlFaLSoKTWdtKV9ryMAkssHsZrPhUjrd8y4iWBf38JxGm+vFQWSm
Kkrrdj7jQueheOhUmawq3nJMNFXpZiJZaaBBySswJkxXfOtn7iJJoGPhNKoQvwDo
ha0kNYSXDJhvnO2+zAuA8HSOWURduiHdJh9aFrfuBoGby+P5zYF5v+byeewvQDzq
APg7Vlk7tWNkw4eEo4sqIFDl0TRByBAJH2G28i9kNZonzB+HJDVdXf4lPLX0MnGn
yeejFvFpheRTLKaIng+oOvi79Tgkt9StWyRLNre0Xv/m5WaR0QQO16wAmk8blmTi
r3akgzFLIwPcOL864EQVfn1ptpwHFNDJdtncwRg/3BaE6LxdhyMgKn/iN4pgsUfa
Xcj7Ea0igjAZV8Z45YHzz+u+BHU0x8AfsZz4opWwBCoBBqdz79Qa5P/q4nn76APy
cf9EAmtgGBQvxgrqC18qBL+FaioLGtFPr/KCRdJwntNF6PPnYmxvDNyJwVFfV++N
Kinf7tNqB5R9+RLaiZ0qsP1FzAiJsR1Ly99/afj/D01010/PYwf/xJo/ie0UQcVd
B0v4uP2UKODNjHLuuAYkJA9fcGjjH1oNsqEmCzBsb5sU56sJkG8Ifu9OSTvKXUKy
qUsZHuPf/UCLsXEhI5QkBGXQaAFH9HnFC2gsdi/5ecoeh5/NEwryq4qkgRTqYZ8D
kYTJHePJIvxwXNVl/OYtt8pnzEMxSaLAMbW/ULqD5IC0+DK++wO/WRlwIfh7o0b8
vb7oYqgX2u8NCV3zsZGLeNj2n89TSEIUa6q29AYCPejwf4YkU42RcEfSCONJGK8Y
ZEqAu+nG9jvxrUd8v/L2JUyEAJepM9/Olj6nC8lxVPFgqA1RvSBCEfgYM+gzt0rL
QM5KKt9hGDwNFzxF6fI0rbWcMZTIOS/g5icfkEyrJQrUDrpgu634DsxxEF49aQJN
le141G+6QtiemNMmJ45hmPf/Y9EOesjVMzyuMnY7a4xpr+c5aZD8Y2ZkWuZ0X9WW
ZUasD/yk02ZGOz8iATtDKD5lS4q2GXk6lpzy04aYsnPBuNh+AuTwYNgMnuxGGHp+
H4yJbljV00h+8yNGqTZJnHKKWqn0AWTrBzmgXGEXAkwdIYkFMm+BTdqpwd6u7y2j
decvjCfoQH1x47rKgY7uHvKkuQsoOU/kZyBnEg15KWlVJW8mnGPb0WIrWZxOofrt
tYfGUE5rVlkWnU2edM3yYs24UdEy4sQHiDpUO3cMvOfdX8flvGd6PwcHmYbvbv2u
2xB1WWsmDlSliqWXZRSqKW6yxxZQ08uNkgL/kHnagVMC7uwWau7Z5HnLZ/pV70sc
o86xvdY10k82U4fWoKIAPJy4NYZ8ljBidPf+ZttEnPmiY+marmw4cZtAM6Ek2RVl
cy7zBpUHyws8oRlGcmio6s08Mg3hUELcMqXZnhy3fNTwmdZNxXqM2gazxO/bc5rv
wO1bE+U1mGQ4/jkmpiAaUwpSvwBMwF7/gtE6ePg2YKLgt6VSDfS2Rm0zYz2oLgUw
ZMN4kYyrSNz/3AMfvIXy8D1Kns/w5M2+X1dmysLrfkmHcZdCKFdcEP65SRLM9s+Y
8F2TTLMG3BXULwmHAeJkTdnBe1MVBT5JviBjmnS79z9a9jnytjr2U+mavWsAIMWi
UCIz/Cf3FANwx7y0p7o/HKeWXd4GS73YJHxm6bXOuIDncPSwPMxNxFz26Lb6SzeT
8IWXq4mzqZ+1KNTHbzrusbzuwWzWfkc9SmDGcZfDpdRAMBVtYFCdSF4g7OUha8R5
D4Ahicr5ne5kT6hThxOvt7myv2tlq1dboRFdlrgU4Ug2n82LUDF/K7xWUT/krEBl
bcxjAuVtWIDBi9lFU/kAYosG4mc4sEPUCxvX+nXqlYWgT8Z1vTCiQ28xCiiz/CBx
hNWMKlwJZ188wddUUkx4r5zsGJHeQss21It2pqMkJ3Poven/Cr7tx4ipQTtb3/gF
nbKvcTU2T5iFePXiU1R9bHdJmtt0uk43ZJS0xeuTn8DAOzBuYc7dK5mnK8p8zQh8
uEoGVf/FI0W1uCtFVz7n7u1yrXiOOqBjVB/CmboD5LF3pCCaI9Ej5fmzi9fTd19v
wQ1NK26kqNzeXVwa3HSs93SMXEEzCz3VKw+0CTUGGZNS0eo0/rSZz88STJQ8U6Lt
pMi66fV+lGhjsZ1B+JwmOA47yOzcmaNgRX8mWw0zBsbPlmb+MUdl3bM6TO/rY7ix
IyJAB+gCeQ2WUUgE2SqNwrZVj9nHhrdCAXJkMvnEB7TRvdB+RYzd13LQXwCHL2JB
4SZrYY3kViTfH7f5gGg3Jh0C5EMfZkUFMI6l1ChxdJZNbtm4OR9RQEdOFdSIYEo3
sjvf9dDqXK8PkRCg1AEo+kKXgS8qt6f6dYF8jWvR8TKwq/wnN1nE+cUugywIyxLY
XcH6JazhTvtI9I5tEYAN1X17YzmXnkKGkSCRq1LeWxFyLXisTiaLdL3OcM50XB1o
rGH2PohuBFC5IfGt4avCSdlFHWsH7r+uNqrwHRN4m+4v+kjm5rWn65Y3OBLvw4qq
QcZPf4SOs4qTdnee7B15ALJdNCu/DlBYLPra2kdgDuYwthY9ZQY0l8z84ZUl+aBR
C5ptTwX6DpJLMSWzACs3nMQI1MIYM9Dkv85k2jhFCHm3NBgAVosfqc0pP0BuimcM
jUKpJbMWoHyalh9eSs/Ry9ncm70MeBDXwvGpoZHkZ1fSVNmQwbxjUSHpK9Iy8r1G
kd/EWHMMVQW4Pc8Lq3SwePU/aUvCa2TUu2OF6Snn5NNInZhI+YQSRET7/PxaAXd/
K2K5UGbAFOwasX6UwGZ8DjtBBf3Ij2STgY1R1qTa9Lqkw5+LSJ7FcC6xdAax8ePR
0j389AqWm9rpfTCgpgKYorpIyhw24xHKV2QUCCumdKciTFNDeaezY7gkNcmXfAf9
ktVQbRjCb9QMkjQ+mKD1rlQazTI+xpzuXIt4q6keJToedzYvuPfRyLTwP7eRGyrJ
TLHJr0t2A6glM2mxw1CQWG3Aa4Fu2bAvYFDeoIT+RvdrNTBSx5jPXTNis2mEXC72
F3B9P81ilfn9tsyCi6aFoMUxXtCYK1NEsxATRGwZI9xs8Jt70z2iGCfVqiw8Ifun
+ojbjBLyueL/WFaCrPKiNQYuRTJp5nvbzJEq4LomxwIcGbWZk2k/OYd53W0XcBKv
yJyqBQ0O+tgYlHPhev1D90KYf+zqDvRF1gAbXlYA2ClzymMz4/tRtXvm6zNQzWCU
Sw+SI3YkrP6D/70+nBO5k7WxG1ajio0KDH1hyVG8DeSp07MT/6Ln499HjRzE4UqT
6kLlFBoO4oUsFzvISqhExwIyg2wc7h8o5MzeMe9fJkeTm7cgBBrFJtmGZzsgaaui
Nx6JC/d/29T9AEBPVagxT39mALToSdG2wfDkDSuIYZEGy96McS2gd1SNVboWzlLT
C8tWEiVLS6Sm8BywuKFQ1i8kXD19Ch61ZcbHkTFloTgkUpfnzLLG8SSfenrurwR+
P30ujYfF5XKUh93CfD8GJ2mSY2avxpAXn6ZidBmHU5oUx2awqPeVLRERvtA9WWdB
3Y6Gw0k+vKNjU9Q7g9Gs/IxywpyRI8x2KexJc2nJ1MgptCPTPCbup81yjfZYEqgp
YaRBDw0DAwBzUqJGySbFAWxMvFMQdFbrlQ4w9smf34EUo1dISADJHv6+k1+6C/CC
5UlE2WS52hLpmpey5FiCAnb9wGQJtjtHsGh+mhd7r8QpBGH/pneeiT71EpVKIy6g
CqIt4vQIArEZp5yiSiPsIyHMK4VF5upslIHHLesvlip28MBFld/bLTIB/DmwJFYq
kBfzdJ9jqRRFghljK/d08ExmCsDTTc6WFnuC1ibCessU8ChKnmnGxtbs7H3Zpz7Q
++9fk10r/ljNVqjsk9Gak8qusKlsyhaS+2xrhKOG90qykikTS8FAH/2Qt43eNyS3
1504ONWyb7wYwjmnMmkffNzMQsX3jn/L+RYUy8hynQ/6BusA6GuTSJOaDKl1aoG3
4V8RWw6/xqIBbJMigdl3SzAlaNj6s4cqVnHiAxENkeYi88+v5E4a4338cY9bY3Vj
cqLg3We2kkbXUFMe6UlJ1Y3nqvrPHs8QrWQIYIt8baPLvNEACF2YrliX6bchCkVz
fcl+9zn+wCw5SaSsNjEY7WHOzy+hhG87VXNoVITgK/tsrMwGWqauHsuissoX+tAP
4hEC4PVLPbHSbyHeeOHXmN0Su/rHESkF+NIvDlZUYgBvJ/zDuMtwJj5Esu0bK65z
IoVfrDqbD08HWsUcxbLH7a3HIv+jcwis2dtp77bR1Sso9S9Inf76w963C1VTf+4p
aEpITA2ryRiM7rkv0x69s5LRC9Rf9akCe4OVRhevLmPQeXn4NyZRuZSMAgusMjYO
CASv1LUhAF6nkBI/GPBE2jBZA8dSqlfkn6pZaYEX+NLJWXPLeojVVyYABMLhJctE
xfl0XbkecnLzXNJZqXhssAmBEqTxtmlYuUpnnysjcmv1wUuToOQOyT5cdSh+7BZc
/O6zVEignLrOrNb3l7G3m1ftbR9VZBZEt5q08Wi6War1t1W6zBgbzIqdWD/t6KtT
pdfoDNjJp9OQpUBfuIdoNTBHjmqX44pqgvO40ZnlU+kyPbWn09LSKkxGE+bGpLKa
jq7eSGRdegCsP1Wy4jLGjKdyK2jxUQ4mB/OfyUgJibsROdtJdHgrI8PQrLRLEPfA
XuSJlnP2q4CqaRj46Lf6m2JBgfyddKSc18NlQFs9dLUJrUDgpSQE2blrrO1AmdyZ
M1jSUlD+PxSkS4Uu9EP72tQyjJs03cAFD2rqmGVjyY2aDAb5/S4MbMRZ94Rgwv4p
x8FCNJs5ZMYACJnuaCfdWLw4V/8GvTrmfopCjM+3yaNdVJCiBLN93Z7nhu75UPYE
NtmuD+rA8Gp5BTqs8LKg37gO5DscbCEc/wL8dSVm5/5YtqcmIxf0mgcb1frn2n5a
RyJ2G8d44WBJeyBRT/CLVf4mWvUaLLdnvKnuOFfhHVEwWH5hyTfHcEy79hRJVCDf
eSz5MOpsei6xdtzatvufUqq+sTZeHGJZVebi2HXWzruXB63Gh7cEx01FUgCsQpFr
Ql2URrF2Gth3YKzrBsMtOIcWv79SBPA6bbXKR9CvykT/IRsAvCShnPAnD3l5sPU8
tbJ1WoXKxZXtLDxFU1ySZ4KFLW+5Ro5ST3RECLH3B6jhio5mDvjQiS6k+/6udXME
h41N61P740VS63Pa3bsm/anZ2BUV8wqP7AbdY04cpoamGJsKlawCJ1PZJw1A0UPw
Sm6sQ95nN1ss54tCbGvWI5d1uK7m3Mjj0AbnTHc1upr1cDfRjZknWremdoKLjgSZ
If/CdHF26dJleIPeT6dGK4Ey1yh7HTJKrPyyT/MWYADzrhaNpRyb2Y3J2RF4OZ0V
4xt3D/OqwlSbTTuhrd99EcYWC7kkSObVmBTblZdCO+klF/VJFVBpPwwKTARjGj0V
uMCWq+ND79rGjiXa9O43su+Y1SKWY/0pwE+xlo+mZ6YubkdrSrjHNB+Sa8hCFHDl
v6bcGvf9m9etIobexmBfiGBdr2snfMzlMahnuA3HBoYOlJUbjR9LHlePV08atSWq
SVvPoKb1u8azqqWklbXfKjg6clLol0HNe3N8kqCa7yGWO0V+bEFy1JEXqUGJI7w2
gMeRpmXUs9ulNDpWY9P1Hi0xfegY9qam+uADz+j41xMFD4HCh5OkPmQIdfm6SIJo
MDv+wTs9bT8wf2b3k3WzsdoIw6yex+SfE8Wq/TZHK8JJpTtIRUkfmpSDQyNVF4xx
ee82bprIOPcxLwk0OCkSe2doPbwPJ2qm3sHeVfdqgLlabHMosvmS7F0+K1SyaF0f
M1rDzxS5lgtvMK2pZr1oV3TjfG6a8zosoMQzO1eQfpP2gmR7nj3SEq501QT9JR3p
TG2XdeVv8DaonONxXuchDwBwkqKPURAMTzQJHq1NdIHwrOkAiA+esRUZXoT/VBDo
MizOffujlmGMDFIQs31U76ElgcSZQsVqxUMmJL4KMGjUghFnVqFWHAXmzVnYKlDb
lvJcJ/tFHJuYK8qTQZmaHFWXPOjkIRf4lnOv0cGuwyR3cQvWI7Vw1FnFJiDmL3o8
3xIALhvekrMSIi/3rB+AgsoCdsPjyQzP+cf+RVrO51kKDulGuBS1ihG/obUiAB/C
/JMkwD15wcQHS1mtRU2LGmRU1QXcpjW7oJsQg5sAQ+pjgUNtQHwKw2qTBN0+t+Vb
pwO72cEP5+rHH+67DREgNYkuODMBBeY9p9i/vHBsIMCRMXOt19XbBZb6ptrhmG+2
01GCAPAZPOZ3MgL7Y/8f3blxWDBOGMvJNcQEeQ5Gxcm6ypOXGXQ5qGQMRBurCBN/
1Cu+EsFP+zsXBSjW7LqgJ43acFSXmxXtVgmmIxhWlbC/RtQRGUF6gOnmvtHTmnud
nh5sAXqYD7cajPhQ2v+ICT5n5XdWWVXmYt9NRN1DVjZNVKhwnqSHESbHus9HHM8N
ULImDGJDwcmbOSDj9jWJvRxGAPs7ePbNZSNXsaGztbIP+EKeKVdzXORQaDLcdWc4
p2Psiug1CsDKvPbjXBGJSVvMn4sW6nQKU6UlXPjMCUb/GPCAG7aQt34KbiXbndf5
GqMG30ZU/Yd0YZZIVSGCZanH1Ruvk3ks4Vmqy5z3DeL8Cdix88hy4NkWtM1UnmX4
OH9SOQlefsnF0LcyxT56JaptU7IVqwYKCfaa1kl6fAbOgdbhUj9P4HfsovLBQVi6
Eh0lVVEjvUmEXMkrvvMzZOHcGd7VRGryt04henvwPTkXCOe4xvTsQj0LffX28uaT
9hPdCQfluytgsqFwn8IYUHKC8Ilb966cBTqkbEATD6imoeTiFEgTJUdTMgkxt2KS
iYutWRWVByVH7LXqJFLw9tk2pUVakeUjbBjy79MRh++8fDeeaP3XY9nbSQDwdFRL
HRswnbUUJySaDD8M2e0IGvrplgrQ+lLRTr9oYupRs610xAVhCHAjyKqLK3BY1jGm
uZJvY5wns890pOimh53S8I2fwfN+O7/g4VVrI9XDqcWucSdOf74MqUmX3mDrb32g
PyNwyscp1h9MPX3s1nn5mNb8gpeiP+ZbshGCnwXIZEjH+n5ihZem9rUW2co/7gA2
4Tv8tE5KaJ6Y5fg5Ces5WTvTvyw4AKhmSx5SEmN5TjZBcEiim/+QS+KVcW6EuYtx
V+wTWbVTICJvNixCpGnUo1gbuiJ4Rfwglz4+VoczhpJM2JSvyBmdi18G6EvlQdIl
u0v/WZPHO1zE4RZZxF3POSmp5mu/3b08dDcXJNITrUjnvLpCDRcw76EXdnfkY782
WjnRcgObpxthYP479UKxVZVLj8V75BWEFQX0o6zh8VcXwt+I3HfHBScQMLI2zZRv
N5MsGyahsnyQQvNe4gWmM9b1tKUoOz0kyXTqh97zpUTPZtychBRhQQcEBk7sl/vU
d21sUsLc0mD5oW5GFPLIIFQYHmQAXJNlsEllbThxR+/CyOGPZgqiLdIVHr866DZ7
1oGfu01Lq2j+tp+aSp1ZWp2gaGEvo0myKinFV3OJ8OnXPTNy9NyuO/mrQ/M1hLf7
1vNj207+Ma2GRvfBcjfzFY9FeoeTfXCdVYttM6l11CDo68kCLW1xBw9ITvG6RXFz
gqLDifGrlVLgPvlqjZ42SknF8YX9DfsDYqB/ovYnGSnxB8C6xY/7T8jyOJP4Wkzi
WhA92RhxemtSLZXrp4xHeLphIrh9ws87YchAP7w1xb8g5fiEXJ7GrOa1JsN/sQ23
LDuVO8TQKjJ/DdqNTziEMu8x0BDkcFvv2WZR22J1A6SIKECS+aC3GX/fquJtLU3X
aaNb4Irmte6O8IT6QthLvTqXWxGh0SafVo38BxHdmgKshqhdllvHCLDwQrcitfNf
CD0mcFyMQeRwOkpEgs+O1brhyg/MVCvtP7OWKWJhtc7nMJ16p2eisTTl9XT2KVXL
O/ez+YX6/QfSlUM0z3QDav/oztfixF26IhTDWf20BPlJAB9oOlzgPMvDpt+KcHfU
NPdHnda6PvESv0TQD/U89GX/8SxK8wEzH22J2gAyM7dO79MZ+gsdn+jTunBBwTwv
J3sTmpIh+b3HSlLYPmiJQM72OsmB1K2shcBKvzmFN8uZrhQ8d/96pzyrI4Rfc+gr
zICl8OewzpXDqD0Oae2Q0AFwfsqeN2oj9AnkzQEkOtrfFreehfQSCKTzW9yczhEu
Pj02RvV6GOhTlZZZ467VVCcKh5syW/6blQgL/wxwcsSqWjkzspqwkQ0I5Q1sZchp
kNwzWwXgAKJ97oQhxCeMxgHe5Lp5JhJWDBMT0ScE8xGnQUVGMtCaAX1ms3+KqzHW
dMWEltI6U2KMd1rqRaLzcQDFw1OOoa4UQe0dwXjLLxwNCKxUQucMOi1GqAETi/kM
FMhetyPVnz14CdpOBmaZUINMTfGfVb266J6QVkIizfe8PaSWxknclybPaqhNpuSd
EpzBmgXWkbRra6JgOdN/2gSvkInGbqsctdqE+BcxxYRe/REv2kKoFOw1qbDE7rAk
l29AY/F9auChkkM9mDxJYIkmqCgZJdzmM5ZwgBpf8mAVqNxJ9dE0e77HS0bFxE8h
65PsBLv5/1PcWv9qKp9j+0nUFFSZj4m5FnT7A7bswCquq50n/GnBz65/py4RVuNY
dvpOTd22CGJY/RmsojQ0B6pq7xE9SbVpvDoxI/MgUGPIP0a0Go/K926C4XRSLOlF
T1hk4PjpFq+8YER0VKZY10yp67379v7Vtmy2HNOAOz6EGFEKZye0TqGRGevId8E0
q9FJAhnhjQ1t4+bXo4sJE1g9Ixll3ctoq3fxf+ezpnfskNlkr4z1mP6X7l0ZRkyr
C7dnjvGAZWlU4nBPzqrltEVuVsglPe9980rbTapyOGByk465fnev1qFn4HIwSqvz
FyT8XwAbPdgWTiUJQJinuedjQGp+aAQ2ICZ3oSu7Thh2VLJEoYMNfd4UDJUjq0q0
ZpWRAU5NuIlvkmQyEz29Sm1oWXsgdTTRb3TFZd5G56m9QmoXsLfJEElcVY9p19QE
XbPhbuPOUMjLsNZLNGL47DQLqXEI9ClFD2NZPwVSFeOoMd5bcliplXdx8yppjbso
KGXBzdosvicQ0K5hH6D3sCd+sHuQ6k/PFVp+b6+V0S6kKEC+mWX7u8NG0z9oQKIc
me9m3n5I0l11wp2ACAH0e5levboGrfAVPSIRB/9HAHsC2ydBY5+ODi58yTrlVmKP
EvSXXKZaJ+kBzhp7fTURGwpfCl2tgNg8ILWuF3dln+7xRrNL/ZKWzO3OaSnRNJZy
/wFEOpP3gmHjjOpaWpUcF3aylt96PcMOlFPvj4k7wl9pYBJN4FVr1C73SUI8I7gm
95TnRgd+ATa/cPWvwNG1tLCQKpwm3n3zqnaj/pWqHGXmB2W0mnh4Ax5Iu647H5+G
yZ25U7goUw6EysKm06bMQ4dnKtOKROsKVCKinDG/K2OG0goa5blA0DXvaGncEzfz
6gaC5XH+WuEv7CTHPkFiXLGL+KNV85uPJcX8hl5wdTjwbGK7vuk++BaXDJtGo+CD
KNBN0aqCpQuuYfgdEnBaTWn6P8njkFPJrYx+FeiQM9pJ1NuteBvLZxyBI98ZyBWI
tfo+pZMszNVrZQUn2Qjm++nBA8jjo/s+LE0m8eTDAo6IQcEVUmlrY9tI5Dafrhja
cLGLExl6oKNG5rb+A1PdWiEvaEgmuFfcRfPxQkJWOWn/EumxWoYWCkQoBjcfi4td
ShfX52fwCYUz22iT2+SDPlvrplel8uZRfsuDquB3A8mm3bXu+7mucW0YdSWfxgQT
04grGeTTE9jYOQIN4Grp/tQDI7o0YDvmtUVp+X5tW5qxK5tjxBG+Gwy4CgOrVp30
dMtISnvWlpmGCzK2NTT5HgMJwfFASFniQmfdek2MLXwQIdsvDYiz9CrKA6Q/b1O4
DbzCIvrrBVuI9EyvTWvTsjq3PA8EyWgYWk2J2ZW2wMm5zwfdgVanetWEU0eXP5h7
1cLQgVooTrCUmGNtOELHDBNNMOzIG0i0eGAzomq9niJSlCmnSO35f7iNWy8FnHGk
jtw1ry+dFzjL5MtBPQOI4XBfOMZHWQEEbVpMDSwpKDgPOX1Q+F8zAKCPeHHLE/Vy
zXKvVbo/Ym6cuA/7nwQgi00/yBqSPNh2YTcQ6Kt8mIJCwn1WVu0qyP+COjY/L1Nh
ktG8wuKAJQPpJJu9zcOjsAVJLLO3YrrVHN7gVfjafi10rlSpMUD+mW1JegiywYCp
FOxjCjFXN2juWLkSblLNalYKnDj8vVftZkEBV3hSyqquEKacm8E5TW6BMdxzMRa+
eD4+YulPZL164DPey2P30NYPIU77idO+T1YWd7W/DXI5I7v6oDj9iKfEq7pHaJLz
ldK6Nm1UUFtHd6HqTO6C+biPjdfR07qXPbz+Qu3DzHWjjFTQwMMcP0ofwxp7Wvqe
ShJWYS27v92UsyAdEKc66UkKZ3FOsLa1E9vgqQ/T28ha190yqrjl5Sh+JkXASIrK
yl+F3a7NnoDpl5xON0opNmk200lHUlNV9x++NtDdefw5DAqkQnBaD0D0R9edlqFs
pb77dgkm9zlqr16I0P9IOzLTJKjm/5qI7dsly4wWMLZA+JAbToTu6Bj3EEskGILz
3faTLqUQRPpWJfuy0kHRC7hExbxZu58Udbty55TvMz++8u5TDvdr7g2lZi0NEPX7
u437NwWB/zwkG2w9tobHia2/0tXir76/qbaE8Trv4KyoVLFvy8ij9WNs2kIXbCOk
4byg1lbNjPavt5cvPBr2BgYAMdy1PIH7wJm8aFCGSiqhJw5oPbpIVe3nmsxI7GaU
17af+FgqZrjJLEJ6YH/Z0SEUpAb1Asyt7tg2N11jbLaTTWDYz0hF4y7LgbrcBpAm
HJVOCxUrVK/6fHwFq8bkXL/GLrC3ztJfS5J/wQHBIz9HXwqy3w/lIw6aV22npKtO
9/+m+pMviYGQ0mOhUvAt8othZSwFinjLKQw/zh8vsTFnfAKkib6AvGz+8CqaqqLr
K8M5tUtJQT4xniQJn7OFqqxgRIOIPwjasMOaCtuFl2hT1XTky8D7eVQYRwndnx9r
JzoX2wB5NPVobJLEofunBzATfPD9Qsv066RslHbfM66ADU5+UUvkE1y//cAT5iKd
v6fLoglIs6yvTgbkju+hkKWT+3xR9z2dJ2GpQ++9ljuGbaFaszrtfDHaJcDcC85Y
uBGntVJsfS/QdZwmv9x9hXW8RX1CNkagWnwhjqYbtvnp049PzXGuB2uTVbrSqTNf
ZRWVLrlrk8p0IN0lZZKmo3c692WQ+mY0Aa8fu/ON7TKvDXVUfHM8M5DaUa8FsqIx
XrWfkRVmdPCY+QIq/oZLasrTxq9uX7X69GyaWLqzF7HU12Wp8Jb5QSojlr+Sh/aK
ph96PU7CPIOnTCa4dqSKvUe0orVYEkXdhATiZWHsJ0EL1O4s186fmNbeClsUmgFx
XhShwWAOa0wiMJBz07+9e0ySlsFAeJoLaA9DMlPYgN/oYZMmRM0QzkMZYVTuMKod
Uc7z7mcSmNN574K4Osi1G0iGAbxYy8fnj+JDfn/ugXxc4U8wKyCDo3yU/4mc1B6Y
AtW5xUuiiIfN2hMaULASbvsL8kVqdK1NWQtGha9ljhKYyhWtFguhuVqfr+miL8nA
8uUtYmJFqKeVpi+55tyvlTGvAltcjCKpLmO2O/tHIpZGsXHbU+q5SbfanhSZAIaD
q6ffqxfhQNhKcyKH6oGZfI77OucstNGpqv4mTOseOpBPiHA1owfmJqjAT45Ss/4Z
6ls1M5CbcqHewOl49vl5xZJiWUtKkmvIH9s3aLIjpMvkp6/SwqFeLG0i+DIOqQnf
KG0lhJ2ziWaYeHH3x5D4MCH1BimGBbzwg6p+ymjwTjt90/o2CxLYtlqn491aMY1N
1PA0pduR2L3m7So25dShMbKo8rcROL8GozvepQpgFsrxDgQn4LmWL0Dvgx9MIgDU
FE6MJH9B9i9htBr4rQHggCaAEwrncx9x/1sWYL1vkiC1hD2o0D4XCSF9kh5JEZwf
zVYbBW1wJyp1Jy6RP3KgJpJ7jxTo9G8Sfe8MHK2gq9IroZWv6pKxt2vbf4noMVMb
nFwsFKp11OqNxpfrp5h3KsCZnMzzCKdt7WMgHSA/FgfhN+YjZBqschqo2hfichUF
k1t7mVABM+OvxLJMXdshl/sNUKslATsEBs04W4BHfx82W0YM/P0HlPeCn3AicxMo
Iyuhn65Vemg6RWr54C5fqV8SaOveNykpF2qHfCMU9FhiJ3m43EGLdR15ipFk9R7E
FLqfbmF2Rkr2rozATdnO1bJB6CIM/NSnm2l0mZ8AmZy282bu5s1/sO3TKcRFltIz
VDTk8x+6Qbzza6VjSNDGzexB3EOBmqSfQO3ywNlPwNVTv/X1bGNs+d52yCyIOGwk
BvAjWdJ/DnQUFlnX22j7qpgYHvKhSwsQXc2Jdp5fInC9uJ7MOx0sK7V39Vvr4UAG
cx7s0Mi80Ag89JIlBkPnzw4GgIR1QXmm8XIFsGaAH5J6m77nG232/fe098+qeEvG
6Fb4vj8/uZXPJjFMG5F1Hpu0MjAtFmsG4H3/tR+0Fw+FeKcKeddQ3DX3XAoKiGWv
wPTLyQzpficirjlnmSlXelPE3GJsJdlfHa7U9DIltgdJ6AvfJ1AykYyqeBHCXA08
pF5BiKZTKCc71L4+udjQZy73Cz83lqisTuEpjOHSAar4U0CCUp9AFMYNpsYfzso7
VqdbUjU9t1vLpH3veoMP07WT9us9kuRzisB8Yv4iw75vQOQ+G4SK6J0Vjs7Q3IJW
QGhAiKvaSnvb4ewV4l7fR3l4zM/5jk33jkcoYl1iphDzkiGbOiwBCvGgFqbgNWt1
bpsxUKnrvUu9SjHtKwAkLOiagkD9mx/WsdP/gVJ1G6im5BbUyKoxyrICtSUxb15j
+OGE6RsRdPcY3PWa8czM9naXdrAIh8Csq4zMHUgG3fP5DleMCr8C38Rwz95nSYR9
EkWu7oaXiQDMFBc58ICXWXlopCHQ4lA1DPf/HoUAFMVcJngg625B3ZxUn8XieaXF
crmxlmJpwR+GHVfi1Xkv+lnqvkYq6wRD4KmVXq48QsT/LPo6jVWXB+D0raDDbx5/
o8KtNEHBqO06Z6PNKbsfnKejyyyse8g/7ReY/kydaXeZXQT8GTg6PcV1cgjgHMUF
3/pJtmejXqQLpA2SdzgjFk/2XVOdPUXrvWtNdMBIgGRQwQNKSlcYoE4Chx+H9nsc
yY4wWlV7W4L57i9TXkw0ewKZYAV8Pv2A+8qBEMEBX3ZHobnidnB4PzsWPyUFY9yE
+6l1mTRWBX/49pvoHYxfe3skSTqmQiWc8Q/LF7ClOTXztObogDGzlLjWGA0brTY0
td4iifhLhFsurJpeY4OpXsLJGUH7a34Bz4BA1GAZb28BGv0xGrCsSYlnf3s6L6Th
p0UwDc49XnQkMt/3ITraXNEwMtNMFLmkVXYp14JHDMABK2Soz9M0ql3hilci6eRp
TZX5laufVNRqwCS8UomgZwSX0GJU8KcIiQCls+4t3MTat7JR+BMOb3T+V8A7Cmyh
Dp6iZK8s6fwFaSiVGJeynhor+8dIvMBr87HiKA5TEamDc8QAKXLAtCqkw5Lhob2f
yPsbtuZ9hmQ4jJBNU1meQt0pyp2bNzMSwbUzABt4u4bswsyCdHOMy0NczUSdkYLD
V1T90WL1F/1tdnmnrLtxS4ePtfdMQYiVKPhriJckR26hTzUxs6MfkHFyGf4bbe8R
bSYsDwqhWeA2s5YgMxuAd7idRDVNepLTAny6tvBv9uLP9efP6KRcsIxsqKzR4TYz
WtJxXy7adLWiqkJbhI/poraARa+wEJLR2CsOzP2onHnJeeDcV8aRzwXwrFHRQ15G
ygaBlMHU+iUVLLrZbE80HDgUtrPeoWgFN8YtXTmUDEXdIOxzo1kGX4Q90CX3VLus
aoqk2UFLiClBNfpHXaUyfYpLqjCeywYsSGmMOfFmWWAnARhMAQtLSKKypmFDoOLi
amUuL3wuhzXWx2NK5Uqta3qhkOBoe8vcGel2LuagB/hboVwjeRvW+hEm5zD6kelO
yBMEpf1TCiaCCA3n7O2PNbkeM9ppaltJTlkNH54o9fN7RyvxcV6Dxl7IFlxm/Aka
G/ITt7MpKpYQ2MMs4miCg99oLg0JZ5tQA/ppvvvPtf3M1rtoUZ8hwczrLDBpcpxy
FkU1s08C79Oryat0ytqih+wBEAIE4pNfaNrFqLrPs2pIoq1/zWY1v7ohLKfJWfzu
vmWQl7iQKiy78pHVBiNKXiaBYbi3zhVnfB4AMsfZm7hLIWcZmYT+5zEDzRSAH7OL
S4ZE4OmadQNeU7uivG8WmxOxAluHzi+Y951OQI7DZDzoogaFL3l3J+07RkIHLD3P
3KJUJFAScFOAMWJrmaaVeCMtU1pWMuWAxImOZX7tHyZNerFjLh/FTLEp67zSrRSs
eGy7rcqE4Z/HxSYW6AuopMBBSTwnOyZvIlN3RJdXt+xVr5bKRQVGwrd5G2liKe+Q
a1cuEeI2PiyEGMFoBEsSUapeeNdEftk4q1C0xNkVr39J2KVgWl2TwLJBhsSEE9Tn
3do4ZpyKhl1Z+4Ay1nfWCYHg52qm56GkZzvsQ0p5/YufBrg525hjJzy/noiUBa2P
v/p3I0E9TDBof95CnI5LtRnW5Qi4o6aa1iJ026L0zVOcURXZGUhRKWIiu/X94FE9
m20F5Ci7yF24Ean9r4ORq4+iIAzHFBVJjJ4Ae5Zo/waMFIU5mKRoPxlgl+lVipgR
lHrDCTvzjOQuNjqahTXQ834daEW/alonTJ98GOB1OTSCRPz9vmT8aW/EaeRtRdq/
SpE3O9knmPNGtot0ifPJtPzVARlO1CFm1oTf3TzQ+tG1ehhELUCNxTJ5LFOIRJnV
iMkHmEjto0t1j//5RmSzjIjdU25K9Xl1zRyOjfFpTs/cFL49H0zlQ1YSq3DjyJmp
JNpBtVXdW32ydXheqJNhuHFvLiMR95hy7paStlUGg+01bPFp3nZqx80UiJD01PZ3
63lt5uJfR+UG/CNaHDKKn6zNikhHNg295Q6CFUzjG4spWy25/sQNWg9IWALTmZTA
wdlzlM2HMtjt2ZeuNzE0L2IfWHuizwPNILAyu5aZENT9ez7ofNUMHg5imwtteyZe
sL1qu2MkmdvIlPPhroW0JR5c6L0aXP6aa+RRLD3QDqAt09/wUIEAxJZmNA8yWzcL
53eglLtDzKvW1frUhl2o/S40lpwHiP4PxrZ9C9bUBIP1Fwueg6fFHcaRlzMaPZIj
DrqYo/MtNKXzq2ThLZO6CxxBHJaUBQ+pJh5gMI2yqMOSoVm2ghpmM0ceutGBkiLT
LJBuo41x2jRKHME/aB5GkLD2RPI+wZE6VVcz/pkAKclKWFQA4f3c39ifig2qmPdB
6viRnIqsbi3r2GvPYH88yud1cRCVq0lPqG/zNseiyUVTWHpft1M2VijKv5HD2MbP
OfOiZNHMZn6Fj2lh/hGmqffHE8EMZYr2PKBynPdDjmKK25Bt1XSviXfh7MpgsYqZ
OEIgPtrAsVyc6wIOYlW3hnzReU1rs5QyVEdPpl/tB+VoNhITZK43rImJT4JFp62V
n3Xh0dLgxszwNipH+d8xWaje9qtt1ukTPF5iZgoU7oADMzRQWvLCjvlZGkIn/4wX
voph6R6UBlQeOQ58DqgFC6zlLM5baLFkExIcy2iSBKJOf6opy0HD2REddvT43S/c
CsEEBSBTYbEdJDhButHQia+zAkggmOHvofcmlGHWYGWzjAd7SRLFwri3Gk6ZNUQw
3RiQUePUfLPsuxRqBNcGUrKmmmyXMTxSw5tKGqchCcnRZGTAb7oHyKWTitYF3VrS
WwyfXgfvSCCTKLyq5Ftxl7HkPtk04sOyFdJELf1mAtYW2qIg1xxkYEfcsgmT8ws0
mMTlXPS7WGb2LcfqrzNJWaEkCO6wggOj3/Y22XsdEurzI1j1LVd6zeH8W4QUZ2Uk
wxYQaTB5hjTMtZHMwTbP8B/QnBGg+1g9NRFjrdjA6GRS3fxZwVBJ9Mwv7ESI4dPB
ROeYzPgHcWrjFnWoAAcQImz3ZZJbXlYxPlp7MKIT2wzX7pg8lrw85t249EM2ijpH
0sIBf8wHaxYUy1iFSbXkASp0HnDR+wzvrJZPFr5jFTuEseu1rw+mIi59lwb5kcag
KkZKgmSJP+YbngeIQwtEwJrIerCC+0YOeDyqxig/C/TqP1307IgV9e0AdKwF4qz1
dKS9S5qOn0a4GwvDwPbcQTgQtjG3YMmBLvDqC/gpy39NtO57/RQSr+67Nz9O9bTI
DiSNrm93ZU3YjqGOIe9oTVpG8nJ3O7ysOUI4t4koSd4ddfPipggRgwgm1OEpRgZ3
3JI4zeFCI7KDqzeiygCHb4xtVgz0b1ZTr0mog5o1ISI88wrxgCisuPjM0FGcIGV2
fEKOIC7nG8R2VNVqx+R/Kbop8D1YHWmU1xOa6jV1mUwnAHGJ19Mym+xBevv/M2J4
tn0T+KdsAsXbWg/sNY0qvcXeyupfkWCP1UM2nIw3FgUN+DFORYirSPbMq6mtIEct
ms9ywjXC4FW1+Qf42jYkSGupuoBi9t837Bg+gNSmWDJbNLuvQklYXGhHIy0tCIfI
664cGgjUWapHtS9xrIVdDND8hFnlvFoariqdOwgafBKjjZmicGg5PbwKJrFubIhc
70S0ImVtsI+RjeHOYqvEgj8ZwCZVFYAWp6slUlNiT4j3rX7ezCBt5jtkAgrI9gCW
1XiqlXAmcBdjxcu0ePYozqf92oJUw6bTqhalR0fEbn5a0AoSLUbD1cSZ9AXkJ+p1
Zy7h7ldbACEzE+iQIVBrIu/LLmjW1O10hsatRpD2rEVqFTWzzVT57Acb82IkGmLP
ZfZjYOYGxCdfB4TMVSaqycH52akhnmivcgKcZigXug9znJFirjXLXmbzEBNcZzKg
KpfmL0iYcRI2PoNeIsBRWHLjbPE28fN2433LEAxuIhMAzs7mGp0rM1pU7PSEN8i8
L9d8n0LbTglOpg7fkZXbumzH+Duzdmbw8stfrbeHUPoG0MNJ0r8Z1n1X1dnbiTZ7
aSH1wDz4TjCFwjSm0wau80rJ9bU/K4MmtEL4thmgQ71xJAW6pwReg3IEUZfTWcCh
hawajE10eeYjxravtAOfStsj2MzyNtTTvMsCmbvQ1Zm47HsVhU+gsD4P2czZNDXn
yvu+87baWGB4DWTEIsz24hsc/1bbKf2vgizfMETKa2bURK/ZCLyNA2zPAG329FKe
YFBoX7KQHMnE3nT7B4AqO0JoVG+P+msupaAc4X71glxy6iSAtGIt08fuQdQo+4DU
y2c50h5ZUYz8krQ/GlveefA52109LtiRVkFouIex51C++N4+FFT349e5fcL+HUxK
OknqyMyu8Lmt04RbpQpcpdK1Si017eiVPtjOM7dnj6sLiPJWtsx548Wz15Z9Eaoi
3akH0P36A6IzGlrE83EvhxkcllswFRIZKCKG2KoAyMwhIuEGgo9R6+F8AyzBLM1/
aNhx3FE9Dannprfqs95M6cXcdqLSqco4Z/w6xQPx/lZGD4sX1BuNSi/NOiO7aS80
SO7yGPCLnmj6HtH2xtGOdsgEgumwi/CILRKqj2mPaMfI6YAIMG8bg3emE4P/26N0
ccQozhK8C9r9Pefim65fhAyV0oFPFV6J1PQ9Aeub1TZRzE7jOdlBRhGuwRi538uL
oVMqCCV8LY8VHDLd+B2jziDhcNYSUV8l5YdDTAZas6tVqsZN2k7QnY5c8wDmlGLJ
jJ8PVR+NTgdUMifO0DmCKI6a+WZARY4smqK3zbCJas3FZxzgRFm/8Dbot4uszkVx
PCtksjszj0a1zHyKG+73Npr0PwJM29ASbzoqzYjyeAsnxNWYSn2u88Y71pUCdAO3
T4ZiN6sF5/nuvuDsLetB8B36n03Ca5njOd0FmJB3+gc/hPZmUcUxG2UAcNPLdoxn
h1qsxKIRjgy1ftwHTlrrN+LsrJYFsP2SwwtFqwIoqg7QJy1Ar8NRiC/PbGssQXUg
bjH0VnmSGMXHGeKmYuJZzK1EGbpQpiBCLIBGZeKtqgDJwhtmi2xOMk3g6wXob6dN
5GccNYNpe8sJrez70VY67SHioo3hu27rquWpD13FqkbG2+N12RcaogrIpcLaCdMS
0w7JIHWQYMAJfhJXabMKih7JExMKbo76iIx6hiSbCbNG+bE39CKS8BaDEjcmrbhZ
3wp46KMcpeE9CfEnYlmRKN7P33BU2vAz+18lAqL0Cxp62OdEbpXWn0mzYmncviyb
lB02MO2Lgek2+ifXdC9S1AM2LgWAjJ+mOxa5eyRvORtWDlEpemdE7BVJT/vL20fo
9CK6sTqd/zb7gdRMy395Yyd5KSlljHtpUtZw3mTyvvXXbVH1KcruY1n2I0KKmD94
ZV7wkOpjyXVfWze4X/WmMUE6RQKpsCphZl3QHxHsQZVu/yTu1djuGRwpCh8G+8Bp
IPeaIgfHGeeM6Lcw8ZHZ5TOEgNNDFGqmOCKaMxp+wbW8F9UncAplNMPPdcDNJmSa
k89LvM41riF7Ld0rwfnNCEbbAkx5r05m/foJnffCi9UCpt2eFhbnDdVCioG7zGCU
z6GOvwlyRI+CV5KAMa+bh0ujuRDdZQ0KyQDrSochi4gpnFiQoen8aR/6EoPEpcpM
T9aloMGYOPio467Bla6Zl3zQRAdWrC9mZdiMJlnZ0IJ/titEqb/mrRr2OlIqvGiP
IMrXRZHdpiWaVxnY0L7hH2IesfUPWifd2zJ+bhrARLcbURqiSLKLJum44Ia8t6sj
2hlmpxmUxbyWut47nbgT0qBAnuQVv9BL/bgKdehhOCuJUUBcDfv2VogPVkF8qjv+
N/w9NAI8eHf2wYpNmBu8fvLCdrUyMxM6BEw1zHvy9IoqbbRLrAE/YZFoDot6D9MN
SeNkhNfMfqNhEcPNnhLpk7HDcbNjY2N+SPjHqKsQV1oq+uGsLHe1viHmZzCkB/zE
HEXFXNZEY4ncdFz0uLdH0RNziEV7FIcc8GQpyDNBuPgJmwO3ph1C31lVUHL42tRl
vqcMMq6yTLIBE/RdfNCY6bkgdE9aOXJp2Nc4k8fZ4Sv7eIJuiqQ59UsbFVJDKcLB
IbzMOsnB+wf0zf3Yv0p5blr2ucLt13UNiFWoZ67M64tlQ7D4AOc19DCRg3sg2ZxP
LAVYjm0BP9gEtYG8afSgUX7qD5n/gnvMQ0Ki1HPitbHdrmOnoyhGElg0I66xXa7s
4gLrPuCc9auJold8PbPdXPXLot2qRIknF36189+klTZveCJz6DYvOmpveW4LgnZZ
/qLEkAwmX5VP9L/4vUBd/bLxjKmj8jXz40+fdKNo3wz6nLmanf8wYyTcU14Z9tRe
e8g4lmhUPLHyspcQhnHFRkQgWL+0MtYRoVto/zfavlSeTPbLA5MpICYdpRQYSq9b
T42PRd8lOWW/t8zutQFfwuXcOaZDw9jrkMrEqkeU1DWt5IMo4wCmE9IYy0G4up/i
N3Ju57nOiDFJqCNvtbdpAwa+5oUrcCQfJ+kREOiIzz4Asz6L44KYofdITnFwrt1B
9ypTeintvM4cDsoeCgLK51FoMhHKMJgJOkmX7bF4f8S+uL/1JBCREbQ6R1Z/tEFm
5xKWc9ZZphQTcDyre3tVtW/Ic1IlfLIqW0bGYUe5fs2heS0taVu+XmMVELaoz5H5
JqQ0c53uiVZVcABQoPitKufqzMR0eXRkQ5qX1rB4SkgO9eNWtHcMne95BZ3LHy1Z
U14hOOQwS3nGwbB58V5NmAFoLzzjWky/k8WkkKj8CnNq1TTTVbET5eW2Ufo6vZ10
y3tSwNXk/DtQVqhk6yBOfR+ewr2DTtPDi1Mes2wlsXbkKu8QSLseKVCs+7LIpNrU
n4m8TIVBTlsGGux7uE9sBxYkYncd7dWGcyI2q5+W0t+9gK7GUjDUGsAGOcKdt5UO
rfuY0gzgKsMSFaLam69RpGvG2xPb7uNsDtFME2qjUsMWovyyMBTHYuouxYqbpiTp
3H0IrbUDGqKXQ06kZf3bqJa/R/lDd89KsG8+VDJg/Rj01pHZlyBdGRL3tPM4Ewk7
bVitpoOld1FXJ9BXU7ZcugOyGaBC7XK3GU18UZdv50dV9ayvFdOgK8i6pkOb73xw
HcT2+5sT/W7/RjtCgihuBErb4t/o5efqEUbCMiH1I34M1nEkgDq3L5Rvamuh9/ya
YrXXRS8+7JHZtNn3NbXQ1aqhAurJSRQ4giEVNNdb6JoWtbAyes5VOqnaUFBe5e17
KnaJ9HauNRCdMr7TqnUy43GZqzJn/FO23l9l7mBesdyFLPWFreUnbB7j99UI6BQC
GC1x1//R4qI//187+TkqxjOrciWq43337/CWbddagMMmdLCQn6exYDlK9W6VZbCO
TVwQrtikPOG7Iqn4FTsjvEFEYktZfmeZwwFXs9B4G6AUEGeR75eyMSOsXHijv8uP
HF7CWb3sql5OTjgysU+y/z18yciM6luhzM66uP/QuluNh0/C1+KqUXQ4d1ADr4Va
pUKHlNFebTjnOXVqtAUF1OHALXBz74sYQb6N5Myb52KxSfF8tz0YjMDz51RIIgCz
WZeEcq1WreS7qVajnsR/OHsjSlNGMRytTatOCaSJTevA5SOrf1r7KX+g89zv37jM
wXzZRetNK/gi0eX9pbdKDb+J8+CBNd0Umz0ciNLoQ3cYmcB6dJJjnpoBLVLM4nt/
IuS915SqjscNKW/dMsX/TF/DlhrZ2s3qzDwvIohDM2HkRgK9QeNocuKlb3dBGwmf
Y3M5SggLy2yjF4c5QRMu7Kt7oQ5JO5RLLT7tQVuBWXBdlz588kfZYHxlvFp6MGCE
ZlMJGuNSFT269GV7PFSJbqQLwaItwI7iPR//0tUxU6XVy3XZhL7P4X9RzI2k4HhM
8VW7HKmLRgQ9yokywQS8wdjHhQdawzdVfVu71zQGpz6qzYPmMRLUnCy/OCqfsI8g
UPPLxvXfspMkyWufqUdkT0HTD7Dk5A5Jzih0Omb59epmWiJu79C6dd8/aEFppGuy
UF1gCCNF017sVVYAHQOxmzTOrg2vkZpD2YI44YImagvTC5Or+SJRFi04x/nUcQcT
yN1xCfeOlltScYYF3XF7eRq8WvbDfqQSa15lIvpng+vgwa7DG8I7KfXOKPJ2dhAY
79jilU51kxkJ/rvSm/FvVIs9xow81u5sLMfE4g7hq9PHJ6e/67NiwaQI2ed5RWin
DM5w6gvQkXsX4mxur3oBMfheiLNxSI61BkqQ5dFZU3W2vxv9B7G4Ifih15HBxTnu
XMw+vYXDD+HG7YYMEc4E5GFiuR33G9kuMwd12MXs7J/xtb0s2ysTh7Y0Wuo4n5tp
cBSzBhh7eJFg8hIWflFGCF5zncfriR42XnfGoPuWECQQN7bi+cUGOCMRYeh4a+lT
tJKR5X54jPftETjVnwlcKG2gFiqBK3Z7vGeGpN4SOqnpoJHj3TVgtKXe+U7bhNQn
cc/R/XqGKMIJPcG64FfkqReEc5AtzL66yS9yFK0CLNWgUu158lUxmtCxm8smnIM0
FIJTkwPL0WyhjbNOyaPg5bM5StwWiJ9pVmUUYPLz+TYyjnhd2AGQ8eIKCMFLz6M6
kPMKl/UCXk0WeHKKz2JNkQcRPtJAfymYC67puQl7z0/jKFOXfpxsR3zQfNqTKJyD
Rh3kl6izje4vvf1kGqkN2084czACY3OF4tCYJQvcKMCFPVAAPuUfj1vBz3ZNjnFu
3mobxeX2nhQ5NmT7APrrP7TPczjNcjQsTb30D2XwetHJgTRnVUKUVauiKgxsa2O8
uxg3kkmOIiX/pKyin+jJKOMPO9dsCnebXmwpxXtsVuQLFd1LJbf5mExPv/U9cK/q
GPLm1T/dyTlf4eeqW2+H28sn875KspwVttI3FcuNbxbs1bJo0IyPYIjK9e1O54Hf
B1NKUaZBDKClGNWwRtuWfayF4L7Fl5UNRXoCSRkZghLG3OO2Uwzk/Xd0cy3sN8aC
wiI9So3qwmcZPLC5hzZqdS5UvjyhoM03yA/kaDh7ZYhmx+w2Zhrk5LpgqCcQ10o1
JaqXSeJ8VvLxpHjr/PyzdXCjrGhscQsYybmzPqgKfRvX0JEajmfqZPkUha91Msw4
ZnLc5lBiGRUdeDpOMuKYw83vedFG4M3VZ816nMlYgL194jFOboxRiQ/9ZpOlM7mq
I5CZQei3+f6y6ok4CptDMh7DC2tBX6uHLbC5lbQ4AT2DO+QuwzRkVAfvxjwWMRtG
b1juhj7/2807ccXm33raMdkUoJrtrzN5Ym4YtIIQdYY5j2TMuuxw2rNzDxU3SGhW
5y26IkICCG+bKlp45ZXRdr8TI3MX9CzsonUwNnI9XER1MzdE06fEJ21uUfOTZ5fO
qIQmbOqq4BUTIJgrBQDF+9kMq0d13LPz8iIZWwI2p80ztFu322rIChahziROPhY+
1H1ITsqnmuRB0hyPJf1LjZNmp9ylMudeEocYrdK8LjV6zifHHcU+Ls6pPUkRYEjy
1N8vyLxfnvqgEecthJrDcbgeQoBxtKUAn8f2/nZGEKcaUBJd8d2sjrzd7Dheh9nV
uGoa+ZQwQGVxek9Ru6edr+0VLKOrJOrcPEEIPDN4hIUo5sfOMoblWtVhkOOkhtGO
u0mLw4suvjSQNzXaVlU/nBeoWJ3BgJNHH68DbTNY0wVkxo9lMabQWaOyhdndrLgh
4WlOsIU05hdBZXdHqSWzDNe9HMIBo2MkVgUN+w73e8YHPocScGB1dGdvWplOwWYI
6kQKAj/19FdX7bRj8OTPknAktps/dMrgAPqqEqYyvT+ASeADyCwIJTr+pAkoezVZ
gDtF0ubfMEny63TmS7fMxv2cBaYoyuj5BDUwMllHyBhIc9+c0uqfZAcwPGj6UxYD
ZfZlh1rzXZXeaUU2zuYplkIV41G06J9Sym0UFNcviY/iJMu0/egmSx8DwKK41Y72
0VhuID78FExXSGod0zhRcQyWkgr2PGa/eM5qFDE36k7i4SsEkH9H4wwIPkCzqLPU
32CQiFe26SPWh5hiNOGGuDjfEEvHA4TYtpJV7X0RRS3AbiXLjZIwDbmVup01gxpl
zmfNwd9uJphY6P9HkHTx99xkZvUyAc9wbXC/IsQ6xk4yoEJDv/hhVuIQyDNdh8Xp
L/FpUqSKDDaoq/Pv47jjbjIemKMIk4o1BZV/Z56XAOCZIICAqiUM1zH7t+tUXqag
MMzPQI09ROEAmQCEZesIoeucR3kmZOq8gKB30bE3RU0kJDr7lmjpt4NflLhvMobO
EwTmLwFHjeBL+xSGvqBfeA0U+x4GQnQemBFKJv4D3NvV9HubFeILcurNjPCIUsi5
SXKJk1pQtomZmTX8Sms1v5Ei10x8xmF8CfgOoh00Lr4M5g41knnf18TMsvmMWV17
jeBNygGGr3rs3XvcXAFJ4UmhbgveHTnjPadTrPkEUdRo2lxnCE5dXfx2qfEOEAIS
AfnEfPaqqJfo7ieihiI6+ivcq2rqn6gkJRwH5lK/k6f5wryDBiiM9k4h51yM5WSx
XpGbG7RQfQDLbSad6TQuARTaTgb6G1TOwBpcP1Y3oaUPt+5Zk6PO2HsqxD23n/Ql
mzrJSjNALSHPDnYMj7xs2WkjuoLdsYsJFtoktLu5fg4cVatJ3h823b1eCck//yHf
Ew7mz6x021TehklFV2kd/j91OsgdEi5vsJlWe7huPYFF4LNyPXAiLA7DzdaBzxy8
j78PANspfgYZ1fDv7hJTq8IH8c6txI37ibsbbP4GKrMGUlwl9SkAExxVvI1Ky2ET
ArtFFrTAUjA1YjxKM6HE0ou7kHvh+uM+POVILVdW6kdHNzWl5x04Ore6SE0SemSo
nPt6mPoC7GHMrKFvBc+MPditEQKig0LDG7XWHfT3AiMZ9T0RtCyhB2TsJwYc5TfU
NAHy/i8xc/P8eRlL6v2tvkNxFnYBqLwddYmW5ILwZlKssDL2YpYqGmI0ldc9i4gp
O3gKyZGoQgSDU8WcsMqI56c60ZepQmG1hzYcPILObeGfE2o7P/JJuhOmtv2TMWzz
XrcOtpgaaq2YDttrzwM/LVC4VodvSht+jnzrc+ikCkmJ2H8W3hWjeRalsG61/Eia
09A+Hmdg19cy54hOnpGHZt9i5eZc9IsmmR7ECSFIro5coF1p0AUcRzT9Uptb3/eY
Zo1fdlKIsA5sBq1MJaGjERSTTt+LBgxL7lZ+7N1uCH2GlRAGr1dhrnhTA2BKbi2P
FUqDXEj5baMIps/ZnyZtzX952z+NW7+9+UePVJ7oFLj/VtMIA1xuAk2Ok9LcKo1a
zOSVCGfm2nZNSc/UFcUSTv7ZqXOvDYHguK4KkjyQvIJJW5U2XBxjh44+ds7I1vQA
r+tU9PbGqXU7zYy+NyDQk55ZW87hPK5LGgkAbTPvpkk1+kFg/tKRJ3VLknteltwO
mvaasqQ04bQBgUaX+fzzOoRVuxgDiYCLKjtt5hBPAL47eQfgBmd2/H3GpgtYirEd
23aRD75sDYvM2wfeFx4lfAdaXRFTIwu8tGrqxzyYo6lpPfQgHrTRB53sTlEMlTWd
xOhUO5OW1I7slFVs+yiRn0BiyapQVhvXjdL8hsibswULoHgXo0SrP3qcOq0/jvaV
ehvYMjGCB+wDzRGrEey2QXDp9a+Z6XDciI0YfS3yMmVKt54VE+vdmoy8EeJV2Dxv
i1mibB2Da6e3iNQ1WDzXJrqV1yFZoiWT+NhSNfZH6uYr9qj70oGXmrZAvlrGrrR9
TxsUBPNDoy1p6btulzp85I9ojbYLTttcy7J6hNHdTmnsoT3iXUgZia4cGeuopN1t
3LyLad6QS+0SwJiDsDnadHTvRbES/Eh0/0Bvo7N8Lx/jcSWJYbgqgmMq5Vpz0a2W
MUvth5Felz9/MUNC9sQUaWTd2orha+m39hLAMYb/5nq6q/aPDetAq1mqhyqEjlEt
NYy0TcLx5QTcMsNGFknpI/ihpNj9OJvQishTki/sUHaohjGM1C3OqpmBF7Km6Hxw
wtBt3O4XRMNCOE5wvm+cz4I0e+9SWrxalp+IdAFZz8WAuN7YTwRY5paLhIZks6E4
ONgQ97X0w2ycakoEGuR9DfL675Xa5EyraWsqKy7I7SbT2B8kMxxw7pdEu0E3DO/k
rc/k2xPlsa590Mr9kZO4OtERiwy53eKCWTvD0J+1ud3qjBNBgSlu7GV2LzFVpuFo
+yXamslX0ZRvFeMyoM1OU5RCd72Lxz2IS9veNGFB+eiiBYp4h0Az97TKB7BfeFrG
ugJy4sO7L0fgA55EP72+TuSwIWA3pKeqXt0zHLrB2cfWIxO24PAmKm9I8LjPNRiz
4t/cstV6ZG8pVL892YtnB3pGTKpga1iyh7lF0zOZKVOcrEZOP15GiuZCS0oSOkKS
TYGPDHwnCcAnTE/Wh+6pW2sthofbs5BMd9V5b4LgOC5FHHqdYxMFtyJIy9zRLT81
aRHyYSZcFN7ri9lf1FsXj5ujKAXmUi7apaKzJA2hllMtT7i2j5uhMFkk96UUPcZp
PQwWKLrr45RrmKBOmq7Dxx6nsOpegpa9gxICxYKdgRlxNw7P0VHKpd3U/D7Srhp6
eDSjylatT1u5pw/Vx+4PddvDG69aY2SoYgsUwinqFDyVR4eYunm9Ca/P/OYRXOeT
ewAjXLAjrJz3OXQWUCHMGtGI6JOQIuTvOKzPz+mImzf33nWBMuNQI02R5TJFnIQB
uknqqu3yevuCoCT0Q9xearHY/Fgx5Q3CnAoW7xG3gT4p7WSTfpy3TzBHwo8xQzAY
sU9A7/WlxYXOnF4kTSBvz28JdQxUoDQFhJ3ttrVsCuAk4KVu8S6xoJ7Sqdqdqx0i
8eZzWGhhlVjuo3ELvojINUzzell/l8U83jrsuXyl0nOIRvziPbAIlTUEWFo7L69U
yDRTZy6nNckm68eQQ0bvbvyJ2/hFEwUy3FaZr5c8TUZFe2z0LzAkEiabE+5rPI3b
KhHumBkOLayMM+a9+P4zbAWVY+ct1vS46HVHmxvbPIY7adRu0MFbcvuwds3AZJTx
FY830VFMExXsgB+nhpY1cQqBeyFFMSFuXeHs89BU4xXoKiOQEQM2kGSffBsJl1Cm
HxlXSiZfl37k23FgqAN05YZ37dgcCBX/BHRktaD47+pfkXNGqTlEjiDj5+97kub7
34rKd9WtZbEpa51l2pTG0698jyK4glaMIWcosDLt48d0+J7z4Sr4rDcncXKwBcEr
c8KK+Jv+6PXkZp1Errfs/yn4AuoJeZGFGQ3tHkTq/x5ATwxkBuljSv7pxki91DcZ
Uip5SMebFi/Q3YM7ybfkGMGWzy4Jfd0mOb4sIyZTrFQLPmaQTdrhpoJf9QBsPrCy
JXHVpFkmJlIVQoVjgq5pTUhwLFHQLp8Osf9kWv4hKne37B8Un5PapW2CP55O1gHN
A5u/RIe+pv1OBnGsuWcEJmyG9+R3PEPvbLFWcn52xnNh/tiMqtHLZw73FKoqoou/
Vkpwf9xUy24glyBcZ1yVrwvfPM0J+NBC8AkuO4eB60arp18JgOoM/ERMB7InCC9q
s9/5E7vV6pJsbEgVtUJIrYPDm2g5QtzNeBTCH+I2qsOiKv4PiE4Mlz5rFub5yh5Q
AauY792a8pzHeVHNaqaMd1K8nLUotFYFJmsmsP0q9p+jGvcgEXrHNm6C+s4nixrQ
DMeiDDcOJW2rG2xwpiv+ddVoztRA2ye9xwRIwgazFu8GvGjl3+m8uhQOpwa1gRRf
781hgnMMACyI32iO32qI61/QHAQWXK5CdD4l/WjCXr/+eFSH5RFq8+JkMRxKdhgw
GJCUlm+X6ZOJQoIKhKyS3+JTw0vomnWZWD1roD4UNbXKbj0JAY77foxIljUE8X1w
n8coRhdvaUhn/hJL+81A/SKtKzUPLxFhFzehWZlrK9kJcF/51hCVOuQHkmXTR6si
GDcWxe6RKjIdvbM4IYf9YlmL7b8fx3PsDyTOok9QUhhbCyCcH2ztMprzcrh301Jo
OmQzgW2Rda0LKqNhh6EFI0MSIa0qPhbVmC+EFVkK5PqsxXwikuVNNz4AGI/eCYNN
OwLZLKDWyc0tg2lKHrdnn6r5NtUPK0M9h5t8dZWGDDgVb/LUyU7wv5ko2E8aXFg7
hRIfwRPtcDqpDoVlcmHepOSP1pPSehSrKwVkI1koQoHcfEwlSPVTgwclMlwHRhmX
TOKVAEDobRunepXkU6KqCuVCH1H0nnuH6BWPkLrPAwni92JGAGvWSJ4lFAFxHjkN
qjcQQvhLYoTd0Hh4iHvMFhDSBDWkEEFud4xAkgY599sbXnTnON+L3eo6Sqg3QcPk
cjGieJCJKLpkt+PCsGOyItoo06FtJnv0aqNadqVFH2lAzIkeCn8p5cFN3hxLiiTB
mjaAczIeOdhoEHj1xG8cJjlQwTkENbIaW7Toig+E7JvefaL211yB7Q4xb40hSzsj
zkvcOZB/YYl5pNKBqiB1RhB/pK3W4UaI3HQKQEWLk3UA2pgX51inYG+cbmkGeN4v
BSXMAcGTyurkCituc1nnW9p4+d/PBWQ+GzQvYX99tXJwOTwTJRtcJXEfdAtYi0z8
pMlB/GD8rtNvRD7BhtcNiWproefjkiX+Lr9lr/ADWicF7LAWS9qBu+hao2TTB2Me
MheAsNOO6BvoqhcejeH4FG0hFAxABZK4G5QTgPEXCtDdjWQwh5jQ65fRkEPgzCYM
Frd9bYjHCVF7IwNkaD8LDpwiW5zofm+JJPiCwRf/358TrFRt+8smhzuEkXdXw/uJ
/YgmB5lTqzMdmDUbMFUe5Hn/RJ5OMJ4TnmkEbqEfBECC9e2+anC28OB9PJhF85bz
Zq5lCTpI/Zz1VvOsXzTv2+gWVWp7EL5CTtrMVr0PfLG0VfkiwF7DVuX64awEneXH
cVaHDVCpdqFIdylHQ1AdX3vsXkPJxVJioprvRFLfd+wkQ0TPSa8rlllDN7qJMHYZ
nvQQbdOb6NxgYn/awQVIZ6e8i9+dZOr5Mrt9bXmdXngLeNDhQJsfIU8RVnTMu5gg
24iek2KJnCEjPP3k6tJy5EtbCk/Ln3zK7YNGa0G8tzYymSybdUCll5sEXztAkZx2
W7j6bNTE41PrxGCBHFLPuhT53Z7eDgaefM5M0Gnv0bBdYIgVdW/jziGbP05Nl8/5
iWr/PBdMjN5E2eJ1mZS1jTW57r+OIFpusu2WxozQe4r35SKrD+3zt19ZIyYvUEoI
z0eDPT6wYeGW/pvZJsb9TqUXDbrMyIaIlofvWN7Kstg9bM/GwjfGMFq6Fv0ZMll3
gqIyDGytgxFLu1NEEhF1RIFCnhIEFsVNa8SnA6X1Dl34150QGt9KZ2TsydkU1ji9
xSCQf75TBSFjcoUJfk9KGB0u6HB6/xW5CzaiyiWM2gxn2aq70KQhSuApZ7UDn1sy
fXhJBAkP4XLVvVYLYbyivqTjzbeH61cxeB2Ch1oT8lejSxOWPBOjnXamgrCFp71E
gkQVrr3azo5s1DrXYdyOupZEfl6HKbrhbU05eekr7Re+QlqvE1XGTiPETtBAU12V
Fr+pjEQcrVSUwb+IFD8MJrYoDGDpzrjQjBUBAkQCKDALTSwWJ5mrXokkfqRbQb4f
2boRgO5zflaiin4G/bWiToh2eVR6MWKsI4xMSXRCeh0y9272PSVZOKKOCLWphy3V
akxeAD3fR2HzslLggZhIS1otWMzP5vEmIxNN6toL3KnS/zp64EFdDdaqAc8oJSN4
Vhcq3+I0DuoZig8txV0EGGu/2jMuWoAi01EVZlnuoVErSsDtLlSIFMvuyzzPs7e3
sRAOw34fIUvMoRoiYogp9AAuqU23XFZaVYT6t4dlqRTpMesC6yJ4Me6S8vfHnHgA
wtUSECwFNoz2BXtuJ/a7TqymQQ8EyHKwIkKcGL1DqjUX96DSRD8qadXmE50UxSma
8EL8sC92Z31CKlLbMDqBO1id27DnZXbYsqMZrw5guYsReQ3xKlaSdaUikiagr7lt
DSHpNA/kXkUgKvHIijePXI3FYUsmfspx1JwWK/40zRp5FG0bpMqi5P8LxjtQZyqc
ureHWQATBfDbUxNoXWkseY/6iDy3+ia29HpiUMaw/uuMWCLhOthRxsI7gxNverPN
1r0lp2TM4pvvZi88uNhM4RVvm0/0ozSEuswCLEZl3AMAafj4RQlGx00LdSSkx1+z
A9SBgGoBZ3GHLQHIIMekpMX7rSxCTLGdEv+Y65eQDMagwNkrtL2+34vVnM5QpAre
u98Ibav/plMakS3Fh3vykizUTbegYz0G4yLaKQcmHrzY5BPbPRTs/C0O8SsbQdZh
m8JfEb1LYY6QkPajSjufd6zNjjrqNV2gATEtz/kDHPMDLo43Gxz1UvaRG9cMHBY0
Ip2ftEJBP+nijUAjgWMTno+3ix+RgmLu3SyxKLI3270II7UyxwO+FH2+AZv2OLVQ
o+sii4HmUb8yNTZtUFHWDO/9H/5PYAVgBMVEkaf16JKvZLDlQppZDW3BsBjh7CFQ
6dpjX++dpQkVJHTcIeNrgx211RCwC0X63x20cqbHeaU9GLY6W8WwkV6zDD2T6qj0
nEWGiYYcRWUdiF8LLe08rw7OFEz+D4KJdw/zW0PY+2JrPPbYGNB6e9k3a/CkUMqG
0NZQnet0DEH5dOZrb2XYsolt5D7Kg9VgPQHHUAGVSCPtY1tr9DeV+VyEcYEt5hTa
MqnwIRybOkYFIrtwyhexhqo3M3liXg9wc5c4aYtxGwtBhEMyeV6uxDhw2NtkorM1
/EMDJDl1/N8G1ZOUISTHXROoU+UiNgT1G+Q5mXNRwEY34H7sIoQMs2f6bS8WANMu
42um8AJI9pUSlR56CG+ZWiNbo8v6+V0sptgjVvdOn8HxevDAzGkTqz55AF5JVqnw
DuqWSTPTzsGey2WuKGtVlVRSDMydmQJB/qLrHGeUeFp44vGDgbcBzvi7o1PMO3/2
8mFYL6+JJrQ0P4HgmhY5iVh4T0F9JVJYqJuj3zXp23kMgIfskEG+CAf1XvOuCYim
tdIjOh022Vd9qcL6TwCEK8F0PqKhNILcxQQRr97ot0p7I3PXwHWaU2z6J8Gc0yZn
BCsqoYRApWNp5BESWo9CQFmyYtP9uhWN5vGBfiPpHu9EKRnldtIsu3q9TrJHEIg1
jIXQrsyyaKaLWqm5QVsipDltMQVyJpgHL5QppcBeeRnXNa65048TK9SbKoed9+YU
hhoXvkHWte18EKWlRGbdcAGW1bnDO5e0JuFesE2P7YWqvANOzzPc59Np3LX+HNBJ
MiMwnVQyfuzHjmKjvBdm5DsDW+9F0fCdsPbsn58r0YUS7TkFKgFY1RnwD1ooA3XG
Mh9JxC1Iy9RzmrJlGGPtZ4efnKUB4J9pYA3lHuxeYvj2BQdlv3hvuQ3IG0exbmjC
xisGu04AhSHN1RAAobyLXgHS8BIywL6VOY2KqDBaXh8ULiAe06SeP5kW/vkCNC1e
FBqlHEUnqx1J4Sc5p4VUO+Eda9VGh+iqOChYx8w93qbF27qMmptTREr+UyA79sEV
zjo/QgESSRM0nyHeyxVtEqydfVwNFNeXsJ+SnQfT3I+xgdjZxsN6ZKGhL9y8sGvO
RunACYkjkNx6l1iSXqLPqf46kU7iFPEc81Rh4Lix5RnwaJNbmbrPUHMhddXW/CAN
L6K6vjipdGBAyptEkIaXCxypJfNoHS/3hZFPP7CNdaDbji7Qif4TGu0RfW3lb2Ft
T2tUJuChYB0I39eqzlqXleLn1sGl2VASKNuvAoQqSWKxZWpQVGsXHzeTGqemm+9s
kr+0WzaOBUXnMeljEdrxuddLXIZOWlIbbALFhc062PvpqEjc29LqA8jvm/3n1Dap
6chJmA+Vz/mpOx8Tn7KX3px7D21e3TC3gAGRad8Mg2qcvjEoIMklht0xEYf7Nsk7
luT1Tw6etzyDb3Zlw0GBllh1SQBHwu63kAfIWncwfiumfNRCNS483bs8oLkMpi9E
sdPJ2iNM3QQ9SBGyF6bQC4NoauXi3/Mp3J6HyC/8qmkXfq3Xe9uAQxtYHspIAy79
UX385H3jWco3j9ib+lhLjmYzlDOBTZ7z8387dXV7VK9ykDN7/7hsxRmhChsIheda
XC6WLwBC8a/GTuYU+E8rl1Iio/jUVyKM3bLKV8mttUnqZexUFS9HkznOzXS0Mtha
GYwRC15e34/AbjezY1t0ktZV7FYfUw1sMxyJMpXCnByBxYwD55sIFxSTmTIGr66L
MSdqZCZGRSl81oWrWnYvvJuKv98LYMVmETvdMP+ylWzsbfk0L5iQxuH8JrE6mxYH
FPeS22l1DooaU6AMkYeZsNpP8h8RAkmwfMztNNJ/ZL7MG0mer6R267XwBYklTBUx
JZShxs6Vj4r+K1osqdEmRW40u+Mp2alk3XqWri6nXZ2C2iCL/7CizRw6eOoUXrIy
OWf3gM0rj2KyWHiWAbWJM7kEmtBUifAkAHIZRYc4wM7XnndarOhiYc+xbieYda9L
hXAe4kJ6SFO+8P6KD6Jv8mya5+YtlsmFAvgG/MImLZCGY8Pn8jv1IBoWPu9NURya
3POoZPa/56zcK3L0dYpCb4PfD3yufQrCJGpgGlOBia1ItLfsd4bfhI/jm7u+mPHo
8yKf9vNPLv+MWGrMrWk5LaPYoyV9ZWGWurDXDLFaeraHKrveWEcVAKXAssEx3CsX
I1srtkus++vDUSbEaxJ3mwn2P+hnzjk6cbQ+vyUf7NgMkBr4ak4kUvhndyNs8abV
eWTZpotm8Vjrhk1RuuLGvQo9uMN/kJHyShqtRM2fhcaIVGFykflXjBJFxP7iQ/nL
5F2zUDX4Q4P7sP7fgUpeSHqsuCUqm7rLiN72b6MClTSTozQjYxF33MtGC+tWs77c
NZNreI2MBDWPt6RigEuV0+XSHsPnFR6T771IUNGlGSZ3EKHP8yn4rTwzykH0pqWa
7SzSZid3/C3ZBnxkLP8iPW8ff3FnFn9XZt2D0lNmKOEYi7qdGyF87wXGb7QjAlkz
+ucDvO2K5lxkIykJYfvs2cq/flcS5Ebct5012Dvq8ZX2O4GGTmPNCALBwsDQjkAk
aduhSEfAC1utBhKoE1746DOCOFTvaIyrUmrVrOfslbZk087h/GyyGwtCqeUCm0u9
kkJ5RasFVsu88WMNs0iq5CGzw2+OYIjNWWMXokupq8cjfxd5aOl0VRaUQu1hQtUa
bPdua1tlnFz3FHYauWZ5IfptuFGVSKDrK1rdmg8qLG5+nqvTrp3lY7IgfcGATVBn
Jt+hlDX5EAYx571leexSSCC1T/Djr8ZWUO06mpGVssEq7eEnxJwOdPVhnnnUb7vz
a/bZFiHVVvM3TVDzFBd8h8luYIDcYOvCBWAk0v/SSEk/2gzPTrbqo2JXFiAyC9H5
Z5fim+JUWjCx9volb+NSRCqC7q/YSnp+1mfyK++8V6bWR8+o25iJGWaAcRaJr0k1
0EFN/x3mhZkCUNJ6mVgazKXLmrIu4ymSoS2KgTsOEw2PDE9MU6CyFI+jBbwJdS4J
S9M6sNZkQjTswHXuh9IvJGdcOc0PE9mCQHESuJhfQS9dnbkiiIAmCssLQplTk7Xs
Pf2Wa4Tl6F6+iUwci4bJRsVAD27tAsuyan6xZFdlibAVpCkVaFraPm8e3tHQ8AQa
eB8WolUJTjxDugkxCHVXx/l5uO9yciDu+W1iZlpnkgKxRVmnTRl4AsJYUClATcYq
oFMjdpf6loZhFXsKsIg/iYDPmfuCrubbwB07IbwAVcFu8HI+DL6NAjiAmx+EDA47
oIFmn7k7H/EkR/nWrSykKWyyBEMBt+C28YTXRUm4eXdGd0STCYMf4W7fYotYxvom
eAYemUNyRyaVDcmvo7ZW/lVfBBaJITy5Qyn+EpmlOoEzUmPm0NXBGybQ8nNzwm02
LP6PeBZPX9ZagvElqz6As9wKbVyZ+3X9VkPyEo61UnYPVHWYhgIl7tEbVm7HNVmo
FykqnCjuYgGOWyv+apigXdAc9nK6AFi+W2+Iuiifm7Zo5K0wdUsi662TX6I/fyyi
wPkhwr0I2fmV5DyRJyMAY6oY65qprJ+DoH5VWldaFWfQsN39eu74smJClzZOaoIu
xj3/QSlBr6p77sur89/GZtZN+JnowBRVS+ZlTuqgje+Xn9s3FnJ6yyuXjbxo/K2V
4rmDiby89aX7Bj1ry/eNLgSKukqXkqC7fKkt2araZyMSdfHnXSOkm0wGSwQgVfFf
6iRa5rfPbtOs+rd8n4BSgMaS4gaDP7mA8pHbDmZizBbHzqK4dsg5m8g331WeM1Rm
AeoMLH+BngiGAqaWWrWHaNHk9MA4i/W/liLbI9vxnadL1YCQ8Vsrq7g79t8lfOuO
SSD9WsZAi4rAxjiXG5fWlUQE5BM/LE3jmYPzb9us8qETOyIt92oICjBdHUQcqBd9
TEA/1dXSYGNTM2Jl3vcbdu77FO+tC8y6HPbRvHmBauo3B5YaxtzQf/7b3EhN6tJ0
bp30ImC8PWQWA1pFRzWqew+65zVLbeXxVy0+NdnplnmP4kzbJQHgZs5XVQ89zkad
tUsaVFuZwLOqJXB/fOWC+KrkwRIUCBc5ykSEbbpK1J7tBNgOvuYL0ZpDAdynkkXl
Rl4eAHBLcdkCQtu0AJR/TOEHewqIPB25hUqOqWzv12TKKpVF5XYAEBX7hldl87hA
Cf3oy8DRW3tY5wtYSqCrqKSTJLGa1yBn2qrRj8sZ64SRfRg2Xb0UKVqLk8zCqkLN
km574Nj+7P/BaLpNCRMUL9uqmOQu00HKasfATjNrXgdgjRr5Gsy7aHgrgg03Bohg
ejTiTHCH1nmNZjhJCjBd5RZlG834aJLQPekE3+C7L1sHPvOB41HmPGzseIbuz/ci
XiW2ibCJ3QK6tS2c4c+xCprniv0I7rGQcxyweX+Ohs7Ak63nYICPTo/lcCkpq5d6
1bJ2JCjeerRrkKzmISx55ythOcnR/mVMzx2gA11gBPp8+utZ5R6M0Kbsjgc4mYo9
BNImgmt+DAxJ3pIEurJCVrsC0iDaMnGffjkleMg++wrjJF791A5G2ZQ+xsgGaUrx
u8KsjWiqsdb44VoW9Iim0ZsifsoaY2VReVS/AbM5zHZTyWnuvVt1KiLvmwdkxS1d
lheEDjfQ86XstA1IGD1Ufkpwjv9PUEOmrAaxnVI1QvXEXMpZqgZeB/f8VvrsX3b+
IjgAsIEKuCkjwCuwRvmsQ7j9ltrCcZ1y3+brSi4c2KYS+wElBq9/Tpkfj5tHYZpu
tAISbvpLJi2EIrHPQQOCcd7/psm5rtM/xSQ3o8H0kKz7AqzW9sNOd+bDqUsLbqKF
B5tx8pR/pKADixi5V+Yjp2CC9b+YiyMM6KJInk6uUl3F2n3A4KCuRlymrTdoRxnZ
QEaZuBfeabodDywZ7X3E7xHfzG2ONq/wJ/LnALmRhTuzecp3nMi+bVGzo7tgbLsZ
k+ArMiTM42VdbS3f9+9yHoRTM6MSVKuSDpaA5LSAb1rdlGR7YB8M7Zu+AEV9Hevk
ahLTt9BtyE+YJmmKAR9sowkQNODsq4+PD7Iis0X+wKixPh7bUs/isnvZAew14QHU
uZMvF4O+iDpjdnnJe0Mls3dypR2JW5/4cHPm/Cg44Y2sXRQbP3UKuEUpmXh2bI4d
W7hiYxnbQ06QQXaK2nX5hhNg1fwJKhz5rfKcuSMmHy+Vtk4rKXYIHUw7gsz9LS7t
XO2d4XGMJTali7XFmT8D6htwkWmrhFJov1mo8y1hQpPGOIzIwLoSaw4yDSjFkiBI
XfDX3CsQp6ced1hyz3oJyR3BCId+ShmMQ0/W3ffkrhdOWiT+BjKrNVReFMW2vgVt
cnLP/HzHBYOMVQ30DHwdmJ7eGW6wScJRJ6++anT/o/Hpi5giecUbbutABEo8t3qt
XFZhN6yS2PnI+QossEx0hDbn0ZBv1sn59JIDkv9v3CdVxf3u+HOnZvA5lsQKB1zq
NgLuCXPpa/0vxxPjOq9JXOFWlbZLHZ/i2ufHCyQ7aqN6+vZyghtHrBJ/8DwKs3zA
sdDQHSxZ+QyS3QycrPGy0sGs3lV1ElA8Zqc85t6/7dtpuIEjAmp/JjhgAM5mYTCm
HUULD+t0z4Fk4lWLHB0XHqbjCUY4hDBqu1x8g1aqX1pjtBOMFPL8MnCz5FNe9rKJ
JOl31Y7JN2vclTOYboTaMIXhRQYAsMc3NuqrOq+eZWfuR7e/ekC2bCKnL7lZUIIM
34wIWr+scyLyP7H/wWbNMcRgzsve2yMn/bApnuseSpA/OFg1wWtWH5fYrjVRxpBU
tHqoQ1HAR972TuldP1JRonOM66EP5XpFHFpBnuCco4eAih6jjmhg8BBQI503Yisr
Gj1yLUcLVCPryLzyjpA+mF0VtxyjNm7/jzY0l33itAIaFPL7RpIuqr2cBHCDxU9R
DG8Sf6N8r38RPCUozTf/7Xp2g8JeeOD+dF5sFvdJRs61zk8588PZoVqYL21d333z
fzWEIeofCBriOOs1cVht4Q1uqolSwlTspJZB0SdQ1SXwDOYZToo1NsYNUkIWVfXX
txZTXYgmDkLPwjUsAWchHzWOkwPSD8XSgZgyYA9aiy5D5nOQ22jl40c8pzNgpsLN
PZQbc1uwHAxxWVVz0InXnOmjiwIYzW+1Apbxz3HUIenV7JAPPaVKzjfk7BKawydJ
aF+JN0E3/MbQ8U3vkzqD8CyV1RryKmwOjvI1Aw6ljqQ90N6h+4VemgsraMnwkWnd
BxTF9XVHQTCJQ9780ta5DN2sGcL2bSUABM4IgG2Ow4vf3HnJu6WBlN1nOcTSq56K
enXy5BVhZXPSkJ4Io86pbXdyQAuKmnQPqtJ1m7I1PBvO4DfSvK4SICeQIVQyGEJF
LVa07gRBJBBfDjzyR+sDF6Nuarcjc0C31BhEs7a7Z5CaGD3vQ3neXLvtcVLVjCaL
ZbktZk2IVqYLN3YDhvW1OdyH6op920cS9xWlTxXNM4DGQUMYgx6ih87/LfMvLMiV
kO6DP5UXZOKWaCU1VFHkTx/3MXt/xI6YwNTB0JmeQysviwPk0iBg+nwwh1cboohh
wrTV17aI8Gxfwu31y8rbE26rDQWSgoSFm5y/JpD5kBOil6dzyC6bc7mL+dUU4HtK
W3XKLz1qIh1tDLIHGtN8ZnFvoz5YueA7vUXSDfcL8zFjHbZzZx2t0hgpuYD9ar3S
rlQzOZc4/mhKBi6AOjQoysvPsX/0ZjBdP+ZFOt7KBUUhYvBGSnL2sO2aWmx7Xy35
iqHG27qJTRtO6AimwhxMtu2QTKXIRE/H+N+PjHVKHJZa3tcFlIm+RmWVxnQrep/w
`pragma protect end_protected
