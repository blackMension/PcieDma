`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D1//MA0K0jFX2W5r4YeMVtJ2Dxlb0oVU4AtGix2KGd026Xh1pwJZlK5R1gh0Mocf
oO6+3RejBQlUS9LyFeLEiS7+HLibdMOf+pLspmYbGwwziQjrWlXSYs1nTSoe+RMH
jtpnUwost9UB/KXcKBQXzzgqqeIfKY3db9+lhd+FgK4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
wAf26IeiBJFQmHPdTOpIRvZqdqfZji5HvBbDn/Imfyv3YCAFS8ncdkxG4WkgSWV5
ddCeQyKLCcV8TBKrz4dtyyN016C3vsKfEeV9SB3wOIWsHB8vHUs83CSHNG0E6nZS
RZWuu9XLVrlbPrYw0ZdX68vYMDMUJVwTXXqgIns41K1iueY5BJpmizqBE4yxi34x
au56l7jTTkO1E6PfML+4WI0lZha2jBg3/pGUVz65kq+FYUb1aOGQ2ZZx/OvR8c0v
+KRc2xFH+h0VtVYX7Q0n2+bRD5ZEk8Dc9pL1+u4Ew8zvIYXVTdzMgLfvJd0kTfbp
9SOv2LdXzrEL94y1oy6OsrNT/NVt0tpGwcCWHtYNaMAONabPxU457u0+JCgp4zHP
ubHWV9zfVA1ZiP1e2NZHunRmdmvYfZQBDtlHp1ZPWLiFzY/F6/mZDMa3xIn85MRW
Cog70nKL8PsAFNUDcBRt4FZzJonUmz44qGEq5QpWt6iZ+Lpl0DQDcy9RaP0oDGRt
mkufcCDnVMJV6199KlBHj6VNa89RmigP/JdQKUO9dCKqXTajt7dT2E7tsWDRGTHZ
Nt5xtD7zgG0Iyf5uS/kreNSqTT3wJGe45a2/NcLcQrxkh2XbN3P3LgjvHYtfLXh8
K6InbjFkO0o5ZcS+7pZwyvAF3tlmc5ruWUmfwkc76NAjaCfUKpEPEPUXa3JsyNxP
WEqah+mFWFiZCuHP3RhaxaQA1ub+R0rLnYPgQhs8CzPPb3LW20AStyrcCdAVexBM
xr+LgrGO87dSRwqcTj53nxALa0DApOi+Zw9ke23GC0Fm4popDOEUkk2gn/32bS7l
+R1A0KbeUkZ4rB+8c5O+yo40S3EciqniLN6YfE2fXpTxfhO/Zjlf8qJ92c1+MUoV
LOaO+bPbfymIpnaBxiMjx8W6OQ9vGg9YaHS72ViXbvCy/aJJcXOrOMLxKvgrGUK7
Fnd41gPpytCYWTwrnEXwcaS82XYIi8cUQGHxAJsDJrxFNxkw/Fjk5KWndYzsefYT
KBN9aIPgkPtbFeNWwj43Unzx11zcw2jPcmQuePqVszSdpYd9ypy3WRvgcIYubOow
vfe/fthTOg8Y9mVhzXov5JDCeK05t4UVC/AQZFdXXzIvYQoyklB+acYA/YnMOBLk
1jgDG/PwiHIoQbsddaT9yzY6NosUHN8izwsKYWl+kTp0f3cMOE+qMdPJiTeuIew4
YlwTtclcK6i6E7EvFUkk4Hn4VbrzeYe51ciJPOf7n5gsWxR0dKhpLLnEcBi7lHJr
3MrdDTDF3XenRR0LRM4qbsZdiTM1KdojX/2+5qycrObbbCVwNKc5MI0wns+/6Dqg
xAOWT67upGHShskYIOiemxX81ejUhfAu3Q3KTa+aBJK/SE7lnj9nOLk3m6p3fREs
DnOFifMHh5VDmSQacOJz8rX2KEnUXEdMinZgnRAwpTDfuh7ZnBKOpH+P+2rY+lrC
ye6Q/RQ1H2Qf8AFJIRUsFS6ngQxX0MNbWaeD1UTaPsJfBNgWIPgmCuRkwzPD2JOE
3zDNhYN2E0JS/z6fXfWC16YAECZkYoJ7EHyvt1YKe9RqNJ2PetKM3anz9BLOA2Gd
H4D/9BUW80kToj5VYBh4mhFcJ9R8qcHzMQzjBeITcszSGPwAGHHf5EiXdCojdW/f
VCuXKmZoxqVoCjA4OwEOgKHBvLH0H7vBv0qxVSkgPKAa99PSLi/8cVNrmHbXPw/Z
pkxRKI552u31KPC8+Gl7HMuK7aygB5gBI53eRmNB91cuSgJ3qAnpj5wtgzEI77UT
ZTCLxnjsF99YhVDznN9uQP+dBpu9mumlmU00y8LUOYTnYRiQv8kDi5t/Pqozq5Hc
oz9HwoAwvU5t5sPeKtCOJJO260piuOf/mzki/t5rVZ/Cg6Akibx7bazvl4tdMbm0
4otRT0pGG2jIRbBcsidY34leTTFq8oMWUINepZNt5t6Kwl1XfR+3PTsi2Zgrre7k
seD1orZ1Ctnta7LsRJucYhAAXP0yowELC3IA/H5nHnuNYKlNruWTtOP8EM6ET9gV
cJ60j1QE/V3JAHBwrZVBOKr8vADiYpoGzoX49hzvPEaOiRbjsdX3UMgeXhWwqr/+
2bV8DnKKrGunz+Q+NdTPuCWIb2XX/rO/uCnsa/croo66B4xNCzHZgkEb5FhzJM3k
PtQxrMUWw8zUwnvPNp76WQVfWTjbqaDwQCnab7xxBUj4S6eAlRLaVfk8wwxEF/be
mIzZImcICRzIC1zViSy8GSvdg2bwqRW+XURZKbGrrNMuKQAVdgvDhAwixyt1iA4G
DBZf7D0sP2k61DVlkADwYJiEMAjWUoB91WVXAbzPWTZ+xJfy2YNbj5irLrhBFrPV
3WYiV/wJWekgNTAosl2F/eIzAmhsRuVkpQE5fdlVC9X18FELD3Qsh3fisM7gtR/v
N8gF7aZOF3dzVcWUcGgoAO5MRqHlgbagZKzb8Dy/SGh7x5+vVbEEB/b6ntHN5l0k
vRgMK1GZY5/tFsNJt9rfSLjL3ulQ0drUqvcPWXW4l+87Q0RPdxKkHpARZiYm2Xos
KecNSD+FAeq02NQvfJz7MOMc4ZipfbQSALYes9nuUJLNGMbIARhZOp5Fjj7d7NbL
Q2OM3T7dJuWTxK+6MMovV8EDqCpueU9ddjfUIQw/M3yHJ5GYl20c6QiJ2+W0ZfBc
PPmKAhuTvNIDv5eox7nA8McCfkSGg1Gbw6YQK//uC92lMEeOsBQ8Ki+ZtLCTuljJ
Y384bz2c1CJ+ZtBXsMKJqFu5/kGkt5TQ71x9km6u7fdhkV7VNkifPT8W815A4L6m
ujlC88aj1DKdrKrmXASPMoXY4qsyZrkJMZ2Z+tBXPgB4wZ7uSjKHWQaf+2tVoaeW
g0mt8HvkRyj11AhlfutlrQ+gtyXaA0VmJU8NM17uuDIvqGvVyvlE0fHIT5+xXwgW
kOhOFlvjsu4JAuZHS+FNDDP2rb/ctutSXeLeLd+qZI3N8wHYT1lMvmIq4uuV/GEY
vZSJKk0jMZD31AYgYAxXG7XZXLPPWIQf0KY31WzTH3i0t+3w0eMlYkxNMOP5qBwI
vE0ac+PEip/Z9bQ8YOi4kAXAEiOhc56+TMVGBwKDcH4/yA9tSDRQz4JlyZZtU0Nm
FrdmXjB37ihOPcDMzlS6B1fRmkuv9rev9oC9AZw+NfOO1s4A8ZgcyAvt1ySq+cFj
162qwAwc5kORYTuGoNBKRPEDsfpKGhS36sMx2aG5r/fcz8FLtzEs4vOg+0f2zncq
5pZlbFAjusMtEkxmF3Fmt3BBO5fgeMTzU42gFpgKWDzorY7gRQO4sDp+P+dQSbMc
1YeXBlTLmr3e4CymAud/kirC1BjJ3ewQercmLhXatqyq+GqCEgZgMUUBUMa0zeSJ
nsMVRAbisqPJIl62hrxqil01cFtoVHSXfow5C14aNflxq6FudYKzi2RfmaMS5Kpl
xEO+DF4AO25KcZtXVNTr6SxPCMwRXoFWJW9fXZz5XyuszBregwWSAUkhtbX67Pc4
PBrfxmtRlBj9sjOjH0CZEVEtdJcfsf37yA6BJMuET4MyOX12sscz9/3fcvfjF2x+
EdaoO9ZAFru6Kr04lFbu9Zkw6Yyk4o5tYL1ouxe1veAfOWBXFwyftmipWHiNkxx7
cSz16iiu+C2ND5qdInldoN77AaYY0bOqXY8zjNWOBgeBRFdJbZWZee8l1YtkzNdc
IzqLST10kHcwa1k/h2++zNKBJpyng0Yxi3Il6bX249Cvcp3IhyJ2sQZSf6GCeyaA
+cqX6rThf+d4JD0USDRGuLZTw9ke6eE5UALxvYFXH/39cWp9z5YTVajWviTZ9Xe/
9Ns/dlc8NEDIXsfdM/pRTKo4EXOV9P09T3HzJ6E6lr1B/7aeB4BcH4aZ8i1R0JI6
IBbk9H3ffeHOvqGprPTyBj6ae5FBHsuwJnzdEZzeTdLylAbs5hJeKv2RmalH1mT/
zC/VT/oW3kRKp+inoJbJjX72I0K1tOnhbM+WSuZxaIf6n6j0m+C/EGpYMKHFeKLx
sesYYlLUEIXhxonfqcCnZl/Ujob01Ae8FiC73V7ly+BgaPVm1n2QjxI5njFYmvKp
GPoeMjDNIUn7qHgohmmNIOREaQjZKLZ+mvdnhHBdftQSS9Ve5eTZ7o5eq9Dsjynq
HjB2xxtqiVFiisVkVlBD/+CRvJM3YUzFPjN0Cc+EdTkPScRrPODi38NzsOKxMt32
8UEfFHyTQ6gMwww5ExyYOkLPW1g5VxERUQaJ9HeufpfRGHdQ3C5+z0VLfbOvOor8
e8PqyABtZg1UFJI771s4Uyub/PY2mD2tcJ8EQMvoBuS33rO/W072dQ3Jn7l/RF6e
EDWzFJKLOItcQMKm9jkcnOzveVfQT/KdhFr8ZWNZFtn7fA7RhKc89enDsmSkQV2a
y6XT8PEkarfr0jAsJpTQU/CB0ghlaf3WOHk7UwyZTe9me8sIpxOgPZMNm3LXtLMU
NVRY6EhE/7pVE/scSgFa5eLIeE64gBkzKLW8p7PmfFFpDRc+m7kkPnECuREhV2Bh
UA+hL6EYCyiZSS1W133vRlEdrqBzRw1zHKmGIi984bh+vPpgX+wx3PtKVRoRmmWf
+7MnuVOVamR3liF7HNmEd08k9CIOMgn4Z5mqa13tASzS0GDMZSy5xuq2EVkRDhRa
2A+A+PEc8eYXQXRcrTRFC2W6tdMa3mGeJg+lWQZz10Yzu/vRT0dn5wSW5mbuUftB
teTBHzOtmSUVo8dy4jHHuU/6bFrBtNS9G/nkl2LgqxbaIoCyrVVz9e2oOHrjU2ZQ
VlRa3OEmSTZyck7HVHWG2gCW3Jxhnyz6JgfcRe443SZkKMZ99wnIy9hay3pJTkD0
2bu8Lgcilr9cQDXLCePM+dktXiYBXmv1rqv8UK4F/2EmbhwzIUypGU8RXs4rhNYJ
4JZWmJzKcm4SNDowcNISeqxmTJHwAvPsEDsHkt2/ay202xkL4UfPE80N8OG+qkcR
Qy/z1t7W3f58QCIahU+HOi5oWJ+hBhnufPsp6SLR9UolBv1RTU2JKMniwP9cRhki
4qOSEqR+S5gw3aDYTx3xutmsiUK5+J+ol2v3+5WAuLONM+ZdseaQ6MA/c8QrZbtb
h1t5s3o1yrz9OgAITdFQjpuwRZjmdkXkvqLHZDQHkxwqhw5bXNymrSSuxd/wmxPv
3LumSElsXl80L8cHb9u1qiLt7Bw/EyjmlJE9GBQl3V76vF6LY5I9fRgXUxbRKhjY
U9l3MOpHKOYw1FJk8oGTdH/YSSSJF1xbMI5V5iGrGrpwOgRRTo/bdJYclJjzi2qJ
Em3u1WCidv3B+hT74MxZPYM9OIlcEd3NwLVaWeOg4a5ihUuiq/b0dM7eIwPIQZM6
fTQlhw2LV3669BAXmSHiqhPvghPcTrjF4i/B9Zsi0wgP49XO0QcODbjpdibPjU05
sWk9uB0lR9oCsgNPRdk/xHAw4PxfkCIVsqKWeip7TuoYHPXr3L6WV9/H19Qfc6HW
2J1BIBZ7oXWeIcusMtnGvNaYxZOEJnNxSHiLbNYaa6O61HqamvZXYKt5lHJk1c6H
PzInQEYi5xVzNldVgj3kGb3ZyRvP4fdNy9VfVQKVIry34n19hEa0Jg3+IyTE4vdh
U9rjBQ1eKRnGFnL/iUz4V4tqdLv9gz/1TbS6MVLmCqqOu17aFh1b0YIqawspATbf
H5rv0pEaobe9yIBfgPw41T9rfEQpvPLHQZ44TutH4kmk47yc6ywwZHPFwm6JZzuR
siqLt3Bm6e+uMVAqrVLHSd2m5r4OUBth+DV3SPeXgbRAaO4b9AeClvMsbot78Get
qPzyNhjLRlxRKncHjlQ8qDcx39UE4HQYljml8kdUtM95jEqjBa6EWQMKwOjRhNlo
DsniK1X2xVYrzoAa6sMaMGdWtrTXc8O/ls9iMhPzQC0hiIYkpDurHLrNsB3EYdEE
yQsutvM9keEjxV1uvwI6l/ft704Lyvj0OtCktP5oHXgZjDowA2FbxExnF3aIiE73
NXcVlBn0NDARXEjIn8IwynQ47LzEVmWLnJLoJbHY+Qzb1XdFgwP8t1IFLeTpkTml
itWkG/TgBbBT0erGsG56nGJT4eVMFmUyEqpnPGpomFbNGWzqZU6z7JhmMnSyzPOU
Mv0bBZ1w5XPZEltDWurq/Pjf2/8+H3JTfmPb6QmYIgLlnSf7/8OJXjqn8773Dc/q
m3m07csul2+Pikvs1p2C0XGndRUeI4bL2X+ofW8xnvnNnwx/tnOJ2trVLSA5V8wR
gTlxFEUzULSz5ikfDn83bH34Q3pYVWij/YrveVi2tiNQWRgdQyYHtGFzMr3y8gw0
NlHR+eyitS/HAwo9DY1iRiPjT93mF0QWXP/dOKVPdLt34EPgAq9KUrPFPvpdQe9g
LJ/F4RaOzBwQt4x//XWiJXTT9igTLR/vQZrZep/e1QfPgT+sen0Q1W2LfYMt7a9i
N76cKdcWMMDh+/kupzgZfiwSAWWqY+doHOthN578yEAENsiST1S0Hl1GmtAfMCWy
XCH7FngdyrP3Q/qDqSah9rv7s32RW1+KfH2vNULPbM0ZrU7tnbIT1t7Svjg1xP59
RR7HykUloA5QA7XAJqRmqc+oYxKovFKPR8oBS8QsrPH+oLvI4D19O7kfRjNFLZvk
hyMoO+JmliMfh1lljDxNa3rtVvXNtRJQ0sGeoSBJQBqauni9/RLfZK2/+ubxNHsc
XtxDObBPHFX8qProecp5IOWk72v1mlsevUzUSrpvccGWzdFMA37kPTp2DPaiFo49
OlA0WAgMZxF5FMrNgpMjXC0/yxFRIzCdAa5zKSeMtb88F2cdC0IRKM7aMK8QHaaH
UcdZ6XYpxIE2LnIHJk0IEgqwQ9sLrRJfugD8F520Srx7RV2s/Vzrlz4DS+y7pbL+
eoi8BLfFJBlMr7q5J3RouU3lhMwA1NTRIAm7F/q4pu8CBrE/y7mRWoQz7wLmqXPH
JwCxGfTZnqE5HOz6YPTamZsGgUz5czKGkuSMkLQFMhcZ2/Tnk7sjwDylxdzdC61l
cBfpJL43Bw2lRWefh7aQ8r8tOx2wQ9AOTzxjOX/2s58Xy6a9ziiB4+3fCI9WIkQ5
Z255WPajiST/ha/WLW5M6HRsCZ274KR4tIrzYQihZiJbNaWup3VUfQhz6CL4OdPX
CS2xHRFJb7e2bSk5Xc5xdEqtjs7WBFk+KZMTw1Sk9xqT7ItBl8Qv6lKOkRQVP+NB
3Af/bqNzj63IDd4uPMYWNcKdYkkjEIeGXHjNEaQvqZmsYq6f6ysCiySLLXj1mSRg
H9RTZll9J2RrmPRFXjnnXp02a5GiTR+RBIOEm09lfcYzueHU6zCRc1AfGlK2EyfA
oRkQ2G2yXHvo7W7dYK68gsfANUDqf0v0XNuRnUNo6qyUwcMN4vPeKtx2WmZ990r1
e8UnbDLB4KDMjeW/+9KxJhNKaY3jLjHgARuGijTrAK8HK1EWIbwmzUO9OtVEo1Ed
gZkic35Yy1PJdodLGy25Gzis+d06NPpTMiTNsOeL3FVJHLrct7XabC/RZPczjce3
VyO9kM+KKnMTWFFDDUQeuzAgbUTrhmWNwJGLb51SnaQEv4mZssXNRs0uFioNVrfu
wXa9NQkZcQcE5jihdQxkKsg1TCsgSIzhhuENskbycD0cykMm43IOCNbQr+egwuN8
z5Mj5wQo/bxwiTy/Kqm8e1UhaWp0rW+EMgvgTppbwEk+gIV6A0QWL3l39UEa41cx
YvkkeV5XHMX3LD0s2JUxh8NDazK0mfvXvwxwS+2IJksQxleNEt/sUpW3LLc0ILbO
k4l4u7qV84GDohALOq9cEwJyQyq368yXHW3eTTOoZvBzZTp4sc5WSBxh0qeHNS08
RDqrkUJr/Zu52Oy5uxMHTN7akf1cEtz0eUuNhLwyk2mig6Y8OYCSFcuRNZPOCOY8
2Duf04nOa9y9MseCGR/+yKc5T1bZO92bFkmuQ6kPkdhAye1+kPHQeXsCHoCVQqza
uOUdX7eCO0S3KprNZvmcqGVk2WLsMULrOpeIhYa0jYorubOZFtlKsQy/gGknsrO1
jAsmRz0/P0VwHfymoo7JvAo/pCNCzYCaPQx+pbAKCBDA4EFIRI3THCGh9217yG3K
/tpWR/LamImVncOWmxzJmJV9Dn6+RfAd6eIZYSalUNd0Memrk4cn/O/DKqUtTJRg
ta4wiDZZtNG5gqge1DP75C+NhVZS6F6M8EHQL1XFZXrZPx7wzwR3vSDoHuezSKOL
Z9juzadIJyhGGzl5Ff0tBS/ahznrU/yLw21G0+ZHfb34CuUABpyWyUzV+YXK48qa
bci+rd7OyzjGYQmyeO2PZHEONokfkfAnvZb0+keH/Rqzm1nIz89AI8/Dl6Nu1706
jnJ3RelWfMX+RoL0oTDDkzNM1Oqq9dG9WfXDg+w9ihHiEVZ0MIttu1y7ZSGnbN/u
7aGNfxES1iqzTlcYiH2Tx8rRMpPVoTse+wUHMl3GN4sU119LedPzPlIxhhC9XKXr
B+niWFnWlXi385zo/BchCa87ck/BDtxNvkiuriBQR5DjeCZ9JXykOVxtQ8z1SnAE
2tUHkM/vtc7xV+5bIWWTp1jG/+/Cllu2jYFIHfQY9ymOO/YMRfMOl/JA2YTzA1/3
R/DNgIoYE3pqDDP8Wi40wha4o5AC18YASuQUaYbr/avPLzu4ON5jzAvqBCaAcfQx
hC8yPuCFLKUFp17N9E8cWcaKTOJ7HEngebYm6yCwgeAvJw+zfWFIWpaHAsLDmBjv
lT0JiH3vhm66h5GjA21IOZEv9KDWSbOvGcz/+4HRAZWRDSwN84Sm6hRARMt75rA5
YhuQJOeI4Ip5LZnGl+EryqhKAofDVL4oWSf2vZr9j91H2SFIM5FKZ5wt2vx1iy+k
/cxORex//bfNDA34q9qDuudZuth1vdt8/cSUj/CnLtaTA4rGHQDf2DJ9m9tistU8
H+l6MRWf3ODVUJACuX9kxrjHTlSN1mxPMGt88+bZM5bsN5syKDctWPH1s9zHBRax
2H5ZG9k11jnztcWgBxRGuleoxwUQDqJKeWUHrYuDzmS/qO/EayqaotcLmKQY8dRE
WVcROrygPM9Yfr7/cSbcOF+3nfaJfEndxishazOtzPcz18aymKhr8pXxovd/EIFZ
O5CoBA0Xle5AWTXJ1PCxSPX/MEVQalvY2EShckTPF+/JiTdTvU6SqiXT/CSjqHIs
6nC2XosCnohC3L6C2aAqh6grQ07foY829dwIve4tVidNq6x1Nn2GxlR6Pq317fPg
ix/fZPdbMEI21IaIE5HvVwRHPe7NxvG6Ws17qb1kSub0xQlgmFnOQxegA6cntXKf
2I6ZQ+Qgs+IZm1HldziCcmkp8zC81M1CQwbGDeqxNHGU2TMtdPIjPIOGEMNLLtFu
0RiW6Zt/alA+8f/rZIYJyCg9+C0AIv3P4SCG2P0yB4JcyHuZZqImHMh/HneYn6Y2
C47obpj62WVhRzoXWffIHEF/+0xkiv52erjK4Oa1EFghUQnsjTidP11ZkbX+ICX+
KIFObBPffbQB6gO7N7iYaOcz9VOz/AeGxtIPWdgzaIWvFwAJaJAjZUChT/rY6+e5
wMO1nHM17kVEbvFqryqZcYFR75ZP3nNyUMxIrkB6BudsbLvjZvCc6VftQycyLw/B
lw65jIbIEDcuO1xfGSJl3K3k7l5Pi4aC943GXRwPfdJiY0+gRkXe2+oEzM08lTh1
hNOGKpP/DYQJ0u5K998Qyo1mQrLqXnIXT7z15mYnvR1nPE33TseqcXzPBtDzRLGC
vJQEUcPXXMophrpB/aZIM08Xwxk6YuC7Ww1sdQMTbDtpFO7i1CfliDe8J6If87ve
zVF7ARGyoN/TUZ3NCJlS0sSiCnG+QWYhmk72V3peL+aQF9crBcg7O3YJxmHUcPgx
OnOnqoYkYiVXuVGibQoCNhndXI5xyzTVGJ3UdqkDhg9n3q4OoARzbHjSuzSXvCQY
F83rabLZEMVvJziV58oxqh7Mc/ZKZMFiO/xlv8lcejHq4rmvfoooB8qvHq/1AUau
AWZdb+Ja6bdX3+8EmOOl8IzK1W911TL2OZeI+I/80CMcze0IUZwW6OmIBuOvkI4C
dIN44KUcH7RK3l544veKBG4L0/X8GbomLqWPr7yjNRLO759+8TtWUp4FGTIxeou4
kO+WeCVbCvcUeVfC8D24pugvZeIEwdAY06W4SMOTKz2drza4BkVRDUT7Ll3/uOth
f8mqTlCp8BSZm52/04T0rRI9qmJvahKoGtkRqYhEQSEpN/0y6n5Ys5zqjg3fy/qf
miptjLRulV8BSQAe5WLzRkgFldBQvHkTybDdd92rIGZuVNRKgkwFzK33t4FYKN5f
Oxas8lavDnT6ECtN0gsWxDoDWXJ1BxtU61Vi/Cx5DS/N0LCNIbaQcDJlqKlpVoON
ucjQmJ2mwgi3/nUKObRtOqFTRNeFLjnGNY+b6jB2wSXWbmLMlfaM8f7esdV8+q/U
2CCsljL9Ax9MYAh5Bi5C5SEg8BCrY+ZWkPBIOeqaQ/1aGXADzPREgaTQwPWGGqQT
zuXE5US+1sfUvhWnhb8wlVg9PE5FCpAC8P5WtrudSXHVNeazBUye8Fh/mMP0reKC
7y5+yw0SbcGEa7baheUaw1iInGdP17rMtq90j61FaXSR+xJDdxn3JK2rtjE8JFBG
aKYqSP37Iuny/l3sMBrG5hZBAKWjgEZnTA0l3IsM9lihYugz2gUSnVaedlRBOBPH
mEH5oV6tx6auVA1sbsVuo/m0M0DbUzVlEGAjMHx81y3ok7Dmw7OfNPQQ8XrPV4AU
6YyiZZDFx+3ioB3mW9bLXmwZ0LGDAbJR1WkvgipIuSgWM1ESW6hS/Wl21jTCY7MR
5parlfeT71N4f8bWPUUpFqZZjuFyvHzjKu0pdYsuwKKBZanu2pRkAPRDTvD5pVkd
9AqKMxza9MXgN4rFDgWMZViPHv3lp0nZBGn2qsKyHBiNuNXXijo/aUGZf2UqkYHX
b/HPtuv/JKTuEv2m8tZ5NUhIQsEJCQj8AHRkkmZQXjtyZYuDFn7DQ3eXi/9AhWpw
dcD4P/T8nXqLthnpGpCB7Scg21p4ucqbISTymQiqinvqBpWh5l9i6cvghnL6r4BL
oqoV5oFDDsHtpo2NwxLXsu3YHh4Ny/Q7TJ1AQOf8C19coBBV5m2gRfox24vi72XS
D9b/OkhpATJFWHcmAnBZfCXv1zlyHHj7ordiEg4RCivih17OKt3bT011jjrs0o2i
0Pu20WQEVwZR/rH0n742OvHDJrLQHgXZtOXMPCz/tN933jlxLlTbK4FKLHccNB4v
RntyZMQxm+1Xq4wy+kzrxye0GT2httTwCnLLJZhidthn443O4kjgmR+0hBBfz0Kr
rrBVJDSikSj23hb6Q53WZDlQm1iB/RcSLNsF378/Gzv9dhFfY9V+0EbkG1FCnL6D
AQyyN1/C9JHhHSEuOLQk+3PBgqXkIdXZgxWIOhBF005EL2n2l5+y+l6IvEUcoZmY
05GU39qn20dAxXPyT2bPKUDBemQR96TERMf9bxU9xJj82cdyT2N2yjOBOfARRDIc
bDlWqp5NAripOQbMWqG4f8l8NzkJKXZK9rph4zVLtzFlr2mEJmUnjV4B6kkkpILz
tgk/Wbg88l0rrI1rGWSLrU+Yd5zZhgUQw2a0YWYZJWYQl4PB2EqXH3RaCC3hgtDv
3hv/32ht6775JhVhYJaCusLcXnC+2yPCMt/DI320ZVZWEZdHz1wQB0/SaNnpc5T4
Hcdnyh77wU8ZisfElsjnxClCGm2P2wVf6Xoun9NhheUjjLIbquOg4u7kisZEwlky
VKecuWuEpGmBGLOKbc+ePVxr1qXBH46Hv8gdmnG1wFNZYNTYuRb+Bu9ooWaTUlyo
DndUhdPuTUjB3e9u7WT0qlo3vwYNCbDcs+wP1wA8JtlZ9Asy5NOFtj4i14eXyfTn
mRPcSsLFuVw4KI0m8EH1vE9ZDIV/8Jrj0fjKU7JeBbx8Ll+UAi9sKZYDVufplb6M
RTcHuYlgRQ/4LbNOStctVw6gT4Xrs4vh5zH2Yqvieq2aabIatOEzza8q5wIGLPhj
57K1rY3QCWuQvrYAbEQ8XiJVlv+oIXhK8pBo3Cz9rTzvBsopXC0x2NQ9MQ/k7l0c
w2ZAQlBGi1e9Pi7dKqmSicdAmSyiEmoX07hFOn7ScaU3fsZaIuEXajduoN5l89Jv
tasn6qYfMONxSFrJMjnC0B6lI9m2ldtZLqjrCI9D+Vd3WzXCDqtX/rlGUaw8SdnJ
ZlRjY/JF2QIg17SG2fdzx6UzO/z0Iy/1Om5grBU+QTryueCFn9AVmN7aIwmycoh+
1o1AqskB0M3vSfe+wj3+HEQu1SLvC9cszLzyBJDn9/9FkrodQyb7bXGduVaTtrsS
lE71X81rNeQ1RK14Uel7x/PM96m8FJVgIRPYy7aPJ+jYcb8ag9fYM2ODgGL4zApz
ljIebgeC1aawMZnFOPizhXIRNPeUBba5ms4o51P+xh2Ui4Sf42MGJzuQn5JAi0DD
oqBWm7LJu0h3sDNejTvBu92Vk0s2e3XVjwSs8JsYlyojtgAXKoJLiYNddZih3VmO
E6XkV0q2Df4b0A1q/l2cHmE2eAUJtP2kvUDVR4mL34tb6hmkyaftc5vw8dZvAPFb
GO1AUzkweGCDYILnw0C0vJlMGdZlWCjrXETi1TJ0Xdjtv+KV/O0o8z1IH/dBIRay
EPCZfZeNTFYzR54t3S7I6yGIic0wmYsH9xwhEOHPYTbCVOjJ3GWHM8Ozo1wWa50w
FIYkCfjLU8L2z8/7ArY8Zp2oW58y2PaDbGldyYSwtrJeSmpnKJSHSY/PBwqO9+rr
2uBnPXOOYvHL/fs8FdT4hYANjqKoVEnR4mSvUvT+77NKlX+1I9SxogHF5EZYGMYQ
adCD8w1LrX8GjGsgSZDIsPO0la8Vhr2PnsVzMaiZs/eIExuy4p3I4rFod4o81NQm
6l5L6OqkMbA44jlmsm+HXWn0DkDvQ5jefPlb983OZdxSr5wf7QYpxIQRfSRdbIpu
hNNib8vOseLLWgY9xhQzAxN2+Cleq2YlhnrXOkCoZ3P4Liyv3jRX9v10//NStitI
d3ogQvtltWqttQi24DfHlkM1BQlBf5Nu6L3pOCyu+r+sxe18044HX7gJxxSgR8xV
BaWtut9yRVY6Co1ysFH8ZjZzZYo7fLP9ko5qMWxT1BOmk+SSX1QIY4xGD9axgJ3y
f7llPF5rGCtRe4yknUTDQ7zHnBoQoEm36mG4WvNJZU2MhSNGUstKo6iafjyxc0vr
KC7KGps5TkDLfFp67AGF3HsKToE1//gWZW42TE6iWxrhaTyJlgq52zsegVtTsKmJ
cjwfZU44d/2UJDQGgUIQLQPIFszCi01uquNQz2eGYk3Q6Ctk8X7djKHqgdjT4vVn
Vdwz6Usdbpa9I1RSEZrgPRSnfN/cjN8WBNJ1sP3DkHS1kw+QUl2jJoilMx6nuxJd
W32I+GhOvpXcfkBCIBepVxvbB5OhMDvbB4H6MYvmwHndE77fKiSmL7g/HxIvJgEl
/3zFWFpAzA4L0ZKrbYtNx/GOkzMp3IHNNw4+M5/J3r/U3Eo0c5BWArpAvW0L9NXd
oXt3uVRqwUv6QKWeIUFx77LJnryDn64hAKs1xPggX0egFN6xBZON2695wdabeaaR
LGtan2fWWcTRyIa253cvszaz6e8XzFnZLgLNb6nPI9oOep5UoBI/SiUrCu64JFHQ
HoK2zUyPQDMRBtfxtJoSeGeegcghE0F3+o7ewpgerRfbgWmsmP7IBMfPdFZX7z79
wO45tYM99Bfixz/0D1ANJsNHQk0UhYgbJkQcdby6phvB/SSp90C2DlndLo0LubaU
lKDDRpEOfUxZ4qobNPfagPYfkEkLPKUYDiCzgxEvXDTsPh8lezQG8/yHwzpKXwRc
W9OBAtc05AzwV9fuwtjoFd6kqoWqqfQ2QStLlCKqkKjpgRaZwcdgH886bqx0S8w/
FfKLYqTp/azw5E3ynqj/bT7YNxxzpNmYSK1hD4NNCWtOP+qjyDshTP3hk4lf2Nqd
6+6zo0MDRqo4gTzm+WwUfvIt3rcmKNXHGKDSbgDmScy307lf/Dn9NXSduu1eZNef
y2oB7EoHYzmRM2XMwMB/7qp6rAdeiYBSRHqPdzZbduxbs8j0tkouKrlGQYl1BxtV
1CE5BLDSxQyijjHEt32193tAD7tRoiBQSfi2wG15qa25mOEKdTlVUpZmlOEqJsZC
YbLeEbMprxrLXxH9MOAKrmNKSwokhZy7xbEyxEFh/ER2Na5Z1EKV5egcJMLPHHF0
uaEpqL7LVHfzLgBRlvl31UFSNBUk9GLvyXXUtUEgexHKU7bdpKhMpaUIbseDE4YT
GzOf57nTNfarAhA1idDb9w3XkvEQJ1U6tjFOqGlltXRP3T+YptPT2qyP2vuznWSJ
v3QuQvSmNoMnwPX7r1Xjiq/tCpAqz+pk0UUCJwRBbMPi00GRsXDzL4Kaz+7vhR0+
jg0za+uYMGldUe+NT5aCfPgF45gtIgFBQ9vzy5C6SQgEOyy66kMb3PX10HiAkxf9
0JF//T3AkEH2PnLw5bQghtxxdxN8VH6Ekmkl3242K2adml9Gm6sdqAKX/3LH14VE
s2Ef9XcmpEEk6YBkaARnOX0nBSnI3yFFNIS8VN78DbX270moNfBJGJXqRDBOPsL0
/+53cBJwDrOOCjzHckPGmgXBi3nlwSzdM7B6Bc8Hi1zUH3e8AQb7s8bPDLOiUHr+
3FwfXkBansfAhwMf6My2BtWZiDNJL1bQL42w0ujGOd49G7OjDlGO5PSSWP6PfNLS
DAZcfxauHMssbPrFUzRNT8DtO2Qeoq9ii5DYyHeon75/X1ZipUDOZJ1PETbm27fu
+rmPNV7aJW2VyB39iqHENHpV8AigCO/riZ0MsdiKGpibAIe8uClF0mn5nbvylcjt
MaAmIidgMeKFWwHYIAxkqfYL1ZpkqIoxxb/pEzxVe4epJYIXJPi7OybBWdorFdOP
J2QxQRlpd8roVL7KsxXNGLPLRcIToilzWZC4FNMPB4hv3VH4NyTmKi1D5fLr7iCB
PgnQaGBgF129jYL9xGM4QGJM8VrEQBIr/aK1v6s6szZBCQVBLYJrwum6DqTgAl5Q
ZMhxclyTn9g8MS5ajFGhi7LU35Rsa1JZoUkVjtwkkeOFXkctvpayfXCYLm7Yx1nk
BW8IolYgF1w2SdfN6pegEIBUKZ6qzb1mJX8LI5KGTwxn9nwRMVclevyqvMnaIcmd
+E7OCMypyPFl3N5fLH0qH9bLIhZpR3B3yQfQsm5YQyoy6sm7jkmgLDIloQZy+/YN
eVX3+a20M+7VqGLfMTXiUEflhrxtt4XGZnM6r3v10hgG6mITGZHogYVZM0J0cOBZ
Rm45IdgheECNgF00gAx0m7v2coQF49Smc9aAGVWFIaVgkZw7PKP6jxzx8AWZUc/G
VZjs9M3UAjPT//ZFHo08NxKaQXdDgnmNMF0M+Xe9hWbLLcLJxMu65aULrlUqf2Tf
XxkDbwkd8v62BrIE/W8X3arPN1iujqnQ6P29r5PpCpNU1CrmmhVUztux8xICGA7f
nCgGKCG5rYMMpc1LWTDOrhwgb+2JQpvuRV9NahPBoG7ZVhdopN1Htqus2QcazIzL
GfF22Ex8DRTF1RuhJ35CyNU6ikjUMBTImbFDN6aN+tjppuUXOQm6DF1twJPZTMos
A4xVOrU+zyY/l1cIKB86boD5x+GX4S+gCcZdlXltynAoQ4DtU3LQ577vkNqciM26
tpV47S9+cF+We+RWcEc9yN0OEgStv7VqGjqNWP1PTDJHOUMQfMQm1M70tMcqrv8W
q6e87szDnS7XfBrajQgna2aemYumOGeZApdoS7S1RO52D+etw6W/ozYLm3R9Eaw9
t9zFqRZxAo+NL9J82TOGLvVBXUqYhTNW21rBYaneWSPuIeNkIWipkpqB+WUoBWYZ
YMk8kaexlwlEYJGOO2caJEHtkdxYNHu0vFNiVpBaLaMSw8019Rx3AB/Nq+JeJk2R
IW2hnApaxlRSty054CV8kSa8pWC4MQR4tvmMKBIHQn1PWpHh3TT33qxFAb2ZGrRo
DFDhDIxjonENseQg08JMG1GxqZb0+b1Z7LM4BKp/xvJaTkdSDX0DgOUBEyNHHRMM
32xSREjzyfillwVao8m3k+EvtcN76OKAv2mCC7Xuzwg8lg0cEGNxa6NY+EIxlvK5
Tshpcc4M86gxMC5gYgnxk4nhJeF1jLE9Q4fAbASKJGObMQXV0X4uIgDAz6BHPRUp
eALVHXrKVK4wl6HuqXZasT0OjHJDdJOh+YNNgeq04Ca7JeNP4wOrJ+Aoki7KzMaH
nXi41CvlC4SowEmbjFrNwNq6xJp4UMmeC2K+J1S76isFx5O87M27Iv4lx1CUmrgo
6lOZAyKMNZigxWJECEBV3uoARfPp9zK8Phm7Ehc4cWUhJwtIzfBDhbXxxTq2cGgc
zTkcgjdEvjI4UVe+z8q096m31C6x56Dt+5CFJMTKQ+8KMbqANfKgH2yqsJ8uRT/U
2XLg39UJeMFBllNndk2qeWQ+0MHu4/Gn77dczy3ae9/HHY3EGVtteeMs+43/Dy1k
GAWwoc35iVDdnJs/J0Y1icuGuP7a6uC463FYXYjqOGxWC2c7rDyCB9z35yMbApcF
UszfXuTxA1MQwMuJMMQWbe38Pzp6NBYSfSZ2UEMXuv27j6plnDK2keR08I6/17bd
70hYoCaENZkkMJTcNl2SrJIR+NYWWJnIdG0YfI61Gk6XAEUc2PSQWJDS7FweR0AN
wcjgyTK5DlFjv9TC0LQxnw4Wd6JPBd6rlHhKY2/NgO9fui+OTCzpLR7wmGhTPsZX
Y0Maxszqpr2bIbA0GG2CZV20QxemRtrAoWdsLbDOr+NemBeiIg9uroZoI9bE1yL2
JllmBFWhBlvrCKCc/MPvQkDhod1gjxAih8Yz3pJsv9tk+WfOiZFhPJp6V58Y2f5V
DAHtM5AGP7VQsw/go5nKcCZgLPl2ZAmqPil44IoHspjunafvMgf+ZoHc49vTXVfn
WhVq3aidXagCIKm2MBV19/iNdhHnQlEhh8WUjM3l/BnoTBO1ntzm2hS96YoU59mv
IqCv+MlIdVTJ8KkniH9Ei48HoJq6iz4GomADFB1oC5Yk7L8vamwhrzjuinf6xRCh
71eWnTKy9EZTB1Ep0zH821xEwCrftyDSJ4FTWZuz+Rc6+fxkuviTUNTboeZLc/Pw
hUSTZENl1OPdFPiw5P1CXEd0JUSq+73BFRBBGTVTu0w/Y04LKVtPLVCCNTJ08fpk
vWiV31qcyMLpAtSajRHVJzom1x2iGcrnbEvPmTsNy/Lym/XfxGLrx0wvUmfp5DuV
HyDUMbvzeZX0Bby0x2+FxbocXQ3NwRWMlicy/hSu/X6Y3MzQsCGxdWgwYjFxokxx
2oFay8czelygLmWSx/1oVrIOD/m2M3XnLOMVPvSHo6TSs4Fp/KjP+3LDM2oe2ehz
1ejcL48XR4kEhOkWf0lRBp2oPj3e2IEzBQpXK6tifmNkQ/0uSJMN9xUvejRWZLrn
biyjpE5l+2x+A3IK+tCGasVW5V/EjJLRREEapq3rqZoWwZbj5BKe/IKJP4Q7lneD
M15tLDsqBza73zSKZhpDNK4JBuHt9iFXP8E3LjbMYcGB7tAVR4FXA4jNsPkOkjzm
wWCt2NI/CB3tW9z9/vQjmZGQpuZseCg91MklCeU7Z8iHih418HKIpxj6iHLFMN7G
0LIspKGbrjoBohN+a1fVVttFKfxAx1ZNaHB/uJnGSev3rhuN5i2uuGwPXMUyjukz
lb5avE+4/2ebHeSgsiVxXrij/bBQQGjgc9ztIUeAfgrCnQ1qjcaU4b/pgOPDKLNU
+35BlS+bI3bSPGaTJvRpbKpa02pCj7ViLjM5C5hJKjk2DiK+U3sRC6vnv4id+uhL
vM9ja/WE5bn4KusoixXu8F8NE5KCJKJCAvxizHMe3JvDB91ZgdK8HuBudbZh0z3P
+IitIg3Rikf9W/FlvfvOLuSF+QqMY3DlkXcaLqy0gK4ggT1MJkm5tfhBQJpz/dmz
qaFGgKWVuxkcILghQI/tifbeDK1LR28dOYS8X9jhx99uSxPaXmFj4UhlRQjANlWt
tlCxAn7KF6VIMrqvwv2CYFGWuEUsPJ0qXtxp+tOvrCzZOgfLRNlvNcFp1LFb663I
tQRfNUhy0reSPuzmVG4+VNGe+DzbLcHwb2V8sjfoUgLB9t124Jj9AC6kJ5gidW+z
NyDYFmFdQ5TkzQX6kojSZuVjewk48wUz76xpyr1ozbYEhu1RDvTZcoaEGZWWybtM
EToqd8/RKTTdH5/C7mJcH4RLBzTmVT1A0xTrb2ZSVvmt0RuRGT/R8F98wcPU8BSk
LJnQ4xhWL0OjxtV2a16IqQCL46ATS+trAPpwFWneq1nlO+YJuSB2M6aEP5bb9aN6
TBcg8Sfnwatwm9/vwo+jk1rHrxY8qjUlrN3J7msaREcD+xPApM9OnUH1O+wjbQpO
HNwto3LDvcgzLtpdKQzCBCJ1eYqlqGhKyB1BMonnhDzDig90hSxCavSPZ/wdwUmD
TJV9NTbKdkoPL+GgXIQUFrt/Z5FRxYYl2zunf7+zDo26i4EkLp3jXwsRC5zfyTQ8
RQMwvaRW0habyPGvCgO6zliPMvZ8AITgxhwVZO+ynNe+rYW+8F+X1fErzV8Y2ewz
StKExGwG2WTp5D4fjojL7PTe6qU2i09qhBOSpkOPvnCovTQGdfUSbIsdRDMxybda
GeHBKl716sDkdm8PUq/ezLCrSveOr6BtOSlkijxeP5YCvz4o+wBPgRtMjJrkBQNz
1d1WazXpAEn1JryJBxZ/l93IU6TlbSMj4t3pZybfQEx6fsaHqaJ+wKpvRwWx5z+b
fBOaTTnUg/fgYLKW2frEsTKk2DY7t9OLxDkNBS43oR++rjjXEGeA54Kpzwv+NuCi
JfXrB66LERNgCJfMtMGtyd97U9O32XT/2OgiBNUchebyWoi2O0oS4tPKIe0B39HQ
LVfxURMWM7iSLHEfxpqwqBJGnJ1Ys4gXqCfA7axHDiVMXTBnTmaQYjcBObCLk8Rc
wwS7Hy7Id8iHYV9SNQ4XGIKqgwJFiz1+GD77PvcVKBribzQXC6vjS17UaXmvW+uN
ZpzVvRYs1b129yPMvyWLMUNVKiK9+hdUNBYPKaBF4GaU622hhubTNxbN6LDMv1mq
FIaJmC2d3xm/jW4CeAgbxuncKzhCxjz7yY6v9ZUuDcNX6+9DuWuXk4wT5Mk+M1wt
l0vMRcXEbWzCpJ5X8gNRxyDhUR7038pS9RKbhgPl1YMdtfnz8k8n+GPB9yWnHuoQ
JO0HwqVFrDlR8W3V8qftqac/dLasbr8A9AeJ3owNZFxMcWZXeJ52xFpGjZKOnzAC
LhjxbpJ9sj+NHdNwrb2Wo+QfXQbUZ+82ARbiCEK0HyeCHu0fhH2T/D78wALO7fkV
yV9myZm1aaLJOsT1tOnvHsNOfcCo7uCagsqBdB9PKl1Bl7w4vNCcE/f4o88Zv4Fl
fBD20qpYCzqDN+PIXHP+6rerE3lUV0N5RcF4x/VYy+SnpvbXmRWDQL+7OCwMjnZz
lijgpbLmfYyVdjfCR2tjM3oLtokkpCIvWoUr/WsEMu0WjZoTd9z+gH3BMMSJww8w
7my+aL9/DwLd6eckM52VNMmbDfnRTBEeyppH1SKLQVi8LgEAeW45PoILPRkegUmU
+21kUlONSnd9io+RFtYvDEJtPbbYdF5ezKBhsv2Ndi5C28osuJ5b+93INWqfdR2C
QL19Vkezr44giIRS2GB9o04QAse77SRSyAczs0Jq9B0hJzVNtH4jLUjB4H2IUM7+
DEETHg+P/KtLZ9ndMwndZvvZ+1fYCjzgdbnqrFxlE5CRctKyOx1C8cbInG1uegaD
NEDQqRMFH0+jJ/yIrvbJOMh5KaxXWWtnUcOR82ZbF8EmthjeKQCW7b/BI2v7NAU1
8Z6G1SVtnZhtshDtAfHZER+FW2fDGhTief6WhtqvaNPZZIz1BDwIS/S4i4O4CqV2
LrIlLj+UVyi28Za+bgAPlygsiddaCUALv7HQ01u5KpH+l1HDQaGZrtcU61arv0rb
f5gZgUsRLnFzPDTGTWTRiRPZAz5Mkg40fEvKwuQ9w3qWkaEtWbg5oAAbWJ5ZwpgI
Hb9nGfyqkRq3fjo8yn9aqmuBTD3nDXC4ebwQNZ4Ql/tBpGeDAFSwEGUsMrZnSZPf
dq/Y1OU67ZDHNs0N/14JJojQHZYOl5EI0jiTJOQvwVwCzi6ZetCJGjbleVE6ShWu
HrMYDF8Ff+HPstr2HugIB0B4l8gItGouz23vgdGupMt7r/QOiuicI3YiU2U6ZvtA
ymad8cD/WzK57c6+xJ0cagOZUZpQRDw0Evpr8csS28+PLxhcvjNLuo6iw3Eo8Gxs
U+WvoygNEYtULWANTlRhRYCSBnR7+Y61jrphLpenSPQrOApsN4p6UmRPv4cx7cAM
KYPDwtLvU6whl/Gp8K20WpHd0m8dsGol6bkdku+bS2dYfWv0y026xrxV7VafRG9U
YWBBzQcOXadnGDuz3VwJyVC0BcqTHTps3xj0dQBkcpSy2euc2tLTbkXlGH6/dQQg
pa0sqydljn7ZbhJc9RDspOl2mlXXhqp5K4aQRjtBDrCXIRhH4WruHJI9gkAAH2tX
0Lou1RdJRWFm3Z9ygJdTjI9D/MgWfc4qxNhmHp7i6bfLgDEF5AtDn8rpjupfHfSG
dImBpDdS1Yy0do4IR4WM4AiIhU6uWm/iV9BowcBuhzvJKX7puBD024mRQsJQuo+H
knjkgds6niYN94T3yZByfRBDH1PyZkpZxx8CVWKI18KP7Tjr78ntjiNXk3Zp/L70
LitmcFz6vpt7PaOcu0B/nvZhDR1Ympw7OiDZUG5GQuUxn4EbYYIqBHqhQD0mXEz4
eaT101jtjmkrCBFk1ux9zqo1BLJ0cHgC0vzIYzahzXYbXdBUpnVq2CQdnAL69VVX
ckH7k5WA8Re1vb4qlEMecaAw6RBsg7Z+dSyvGxMLXTWcHa/KYtJMQRnTMqFrBlmK
3OkaTPMjrepv/DWtdpOWljIwtMO160bunCf28Tx+1+MRwzCY/CAifzcoCs/z1P9V
qfmVcprjUllS8DTP5KDIPnn7A9ZBpos1eFBrAAwV4ABikAS7iSBBl6Fy9vcFmtY4
+AwvSlWh0Oo8DXqkMG8DprwznE18z/uOes/u8Zv3m073oYxb3wzcoAsO5Y14+SBT
Qrcymy03TqTA8QH0XtqxTeozFTzVgzT0EsiCujlXroZ3c09ods6D7TRx9Go0h2SK
qXLAUnaHJNUnUVZyFOnV8BLM/mRKTaPlG2owEccAm5JOjXrtoL6MbTXKyPeFd75s
cwYAtKgSkugmCO/Mm/9KcAWHLIdsaA2vE2fPCyFJRjLA5KCv2A+T9zRXOohTacld
zqxMpyRZASazRt4Txu+dTakG9E7A/+e3L4b4CHC5/qy35x7b1WzSVjj/s0bw2Exl
WJfp0sGK2+bzfEsR8DjX9UDQnLnh5fNl/JuA7vqZWHnz5+BPy57bQfx6JzfB8Mma
ul5HgyK3sUGzPeySaEKrxBwY0G8rbtj0/x9ZyRFXijE/ygtaVCwoLcoGOCkILdVL
WHNvQpEmsGGbWztSTXM6DIaCb4kI/xAH8EMDMLDr9Sz20GE+6vS0mNF3dT2422Dg
98y2Qcxyq7DY0lu3ORe7NGoyxTyz6rmIhVXPyfuMxBa/KA7/UMjBZA3apo7B7FO/
NEu0JboqHBZSmBR65lIcmjRRFbFkLdM/vx93H8VFNKu9QOZ+1Zop7GGkQoaJnbVp
2q4s9cO12HaKk+9ASyhocqgIQeX9JpKVsWl0hKpeBW1h0pCUxIDT11tsHAUkxNgH
XJuphxvGqWtv1nJKmIRv6fvlucX+v5Mziz4ErUQv1ixck0VZCYrfmt57adzgrpmt
nyZJVM5MdjHhmXk53gN4zW93QZ3IZR52FPpgbWSMQaAPbqMW73OeWo1fYAlcJkeW
tuzKDxhdGXrqc+fEuLc2V24ZiZzf6bsRmn6K+F1XskruX1t5XuOGPeYu4jHpMyN8
flEufYcHwdjTVkconS09odxOjJw9M4AOyb5LkZA17EG+kw5b3wP4kxjSziD9U4QW
EsAgBoxhA5CpoqN/VTV95NdNZD832R+mS2e/qIg0nedatq5qDxY6JTTGR7RuOVLv
CMRm1wZgHw4pCgB3HmCBCom2zZJhYjcSR6o6CkoWRMo6XZkFdakrZpQMcD9s6l/d
dSRY+FSAgMeHkjHaUs1YKa3d4456s8QUzuiiPg3xxnCmNeERVnSSPmrIpPMDcwrG
RrI1XqNFu/i/DYHG7j3JQ97yGXMyMW/QHI3wBURAfLkgsklbSmSuJBNwi9l+/K2C
o+kF1yXxDPJgrCGhf1SUGoAXT0QOy7w2I8n4eZ4WSRJZygCOuGlL3VbHTeTA/+ql
LY0jZ2n0keCxchQSu61trS1GIQnpzIJNcNLtz2bfj98yUgfz4LIo6OwHGI6NarjD
5nPLcAR6Hv+vrF/JH7enIkpS8Ve7aGJMJ+iOR/FcaGiJgdkqVweiGv116gAoJkAD
VKj+An6b/7ionU6ffWJX+mJyx9i1PDqKOz63meYO9O/aS/T34W/0YGHOYPnJuPDE
Ts9KajbJkjU2Ahg2adh38j2ExlVSNYzEo6e01DW7rcb9F0biTpOHZN1+3N+faQPP
gebKlfBkJfhEPB4PoIS5cTxgRZ1l3t3OL+WBsZF1MsIy9+PEgOBAeCuRsDnKW4Nv
IHooF7mVV0wu/O4dWZY2YcnZcAWq9sStrW0omOvkmly1u93q1fEIoV+aTDE3XOjx
Wd/uez7X9bc7xa3SJPwxbAD5Gj7ReXyIOxUCGsddpUBvpvYSCAz2ZnxkO+bBcTbS
XmVlULTldrSdlncjtAcMQWsCVHn00FzSG3SN9LQhiVhVWkV8gnHn+1BOGXafAdO+
68fzovQABLhedMUJVhtz+C7p4nAec1Z417Q3oqCyUfofXDOUWEZ7sjtsenjlNXTR
6l+CK7K9yhwIvewm+woGIipsWeVPTGpI89jgkSLhYzAC1B0D+UuGRkrZXCpaEI9f
r4t6NoDlvzHzIgg2WoPCw4Lui91i3N108AsbciGKcmWAA103W74cYms6Mw62qDxZ
W+bFe7WlfDwZgz5Xwlnz19BLMsmtm56mG+rJx352iZnTInfSWa48W6PbBFjskr/u
PRNZpKueeQamgcwsHRRJ3F8kNF6Q+yziV/mXB1zoZioMWtJpcboU6NpatvVti7SW
VbnKo9YY48ZG2vqhBpmWJZx+JPG5wuF2wa61ECisG5W8aNXGjZmLVEu1a4U5axDC
7bch6ExgiqVa+OfjEN0x2ADiiO1Pz8xC/rjqvHVOfpcSRBwTMPFO5P0EmQkJ7Qbm
fkktGIuh/HSJRkzmWL7s3TXXw/stzHeKeBRrKJjtAEd198akOdMwvMGJFd3XMEXt
jBEy5cgfMW/SXUrR1X4WtmTPpqPpYR0er5BgLaaQGjShrWQHrctbL247D4Mvk8wO
Sx0nNUzL7KCgHAIQyyRmtM8e94OdXdOd6XbN8y4k8jS/fZ87yZDjf5a6LMV5wy+e
c30C3REZmJhccJH4gaTVGDXn4sqdEkLF09uu+2P4NGV8YiqwMGxT3b1phucMkt/x
qKlF7JMhjHtnmG4JjFSzgdMUR/VIa4engD+kfkZ2g7jHFLenElBPhygyV23xdzam
C67f93LJFS2unQe1kJUPVOgGRMsI3sGKiYXdx1k9XkIC0UuHBc4FonltOykLkddK
Zdh8HQnmeGq3Hv4N9DPeO3tXF9jPz61OXWmEaz/v7kkNV9ffIyVn6KAGSBnFs9Fx
wSvuNUg9RpgXY+d8fpFaOVDKVuiaBXdj3ioi3koEsIccrAvhbdrsPxrYmKVrvMXa
TN9PFP8rsWVFShnAA579tXg81tYgjju+m9gBEu8kBrjFr3cO032jeCdTrTKNKMtZ
VgvBAs/qN7Xal7pztHWYeVXLk6hszeJJ4br2bangkGFXSeu6RASR2+PuHeVaOdqL
SC6d9cmdQ64szd1pUAwi7tiqlWSJyzvTFC0MDprkzXtw4w6xB7cPxLcuvSbU744G
E6mg/KJ+Lvf0e7zy3Ygj1quC6ow+Efp0Ja7TfpHV6FIJmA9wG/hSSXQu5GcDEAgC
boQ7/St1xAqL7pcwSFxPUGz5cw9X1GdN1KT1AeuE96OTdjBog96dJT7KGBU48KJc
dfXvstged/DqJRm7PlhxyLglLxxc+cjds7irreRnBYLnUhPN4cWTMdepOuM5Cglw
zty7Qg8d26WdHrp2M91FmOgwbDY/W14R2Gfd8xVVDAZIeuFKimhClWe9uuvCo+Wd
lQgwc08oSU6GLJBXYOjlokUFXCwY2HRJC/vuMVSRwQ4awvEaTIgtslr5KMWahwOX
ZWa2lfsZbXceHqvwmR6dLZIe22jZ2GFFCly7ITDWkC+zjS3FDaDtppArXEu/oO7O
B1OOD6jMPskQLaKyTlSbPrX1/k7wH19xkph2HXBv4LBCpfB0ymfEAZUCUtI7umK5
ltryk28iAK6m9JRDyc73TMqaZx5YcU3U+bly1APSoD7Qi9jAfm1a+OZgZ4ztL+fb
LeRvHoDxKKWztv4wWH42kUpZe23KVKLuIMASvf/aRGLqyqDSnCroZc0C7bNWxyOE
zDxwKyRWLFt+l1ogGo71IdSjY07xzyTauWiyOXrVQ8O23spDcx/R75F7qOBZmn0H
OR9IoFbywuFC/fzpfCG3QiH2sh7KWrstyAxv8Logfup5po/dFa4rSOIOzrjJbyEn
S2FyOx0TD6PGvqdB6dKvUMDXPIoSSHwWOXbmeB/D2bO6SQXa/dDOQ26zievzDoRI
g4nOZthsjOxAUD93+jgmtnGkqxybAlLc7M132eSQQ4JLRLgmcZPS2ER/so0JYRan
+DIpB2DwcfOk+bsQLkrW1WxL3l/s1bF50fQMtUj+pu+aHFWogFQr2xryzHy5beTL
QM5JGA5rwBoIKuLwBKqGG6GPrssNmbk0HZae+CfEZhItFjCHamFra2DusK5DDr33
/YN2BiVtTHHE1irXEFlfwQl6rxOfWKTPGh6U7SXl4BaUm/VG1Y2sA7oitMofvljz
vuQheYamgNMohdYTdMaIWvL3u1q0II3iJy7+fD6xZjP8CQd6i9EyKjMPAaawKutm
tdYVbiVJl1w24Eok8EPZ2F1ScptpsDxwA0rvGaO0H5/lUek8Fc/QWzPJZVmNE9op
Fxz+Zy5J0r34CBf9uPsUapfTEKcq1iVtRCe2iTyNl3BQuqe3IlN3F0yUhUYDLOFM
egsZPNNwb0YK+QB6DOrkQACnxYw9NE2zBlNKp1voW1UtUCGHY6hAxxFTPSLSm39y
vH6BPNbecTMbR/U9Kyu5lmWpgedQVdr9OAwKkWyCaWEKuSWsAeARFoCYYc2Vd0p3
GI1toxbYvEQPLbBr+6EWOXc/HzAoyaYBbYO+7zGEIlBeSqMPXlHN89cix5q+og+9
XGfxit8BmSjNif1MlcakDcRm2MnpjT9+adTak5+3Ste3PA8Txv8l/s7FkWSWqhNj
IMUN1DmLWQ4lPoLDiDby7JcfAA5FCCMv8LeSfatMnP9x0ujSDIURNJyXbbexhrLj
xaIsFtzuUeAFEQS3VfNHeONxWICvV1pZLOqJLe7N4ftq50SRvso1Zrre/uWxNSeR
ARy/FklmFC7XLf3c6M6njNwR7LurRqzWWot1+wqGTd9WCwi1qJ2PM9lbva0TGDZb
e3yCFVO2cb8DaIOaHbcECzNUV91EGXNEMuMJGh3ETGNiUPxJiRojFdWjcfb0rj0d
Q0fwQdQK40+riSAV7Ts5VTCvP1iegLjmcA1ECh4GsTxvixKxUODNpX16QTKBUCjt
4gZdHripIn72bHe9J/0prY3VLiA8TLDY1xo57YvuKHMYHnDM840CFAc0eUt4+KWI
V7J8WyKQhujl0WZgZAQc5m7S2yPkSk7fnjAV2qwqs8/GMcwHEnM+0Sj6o4teW5S4
nkiKbp5uk8T8wqYn8+yxK/rmU6L8IvHvDguMW2MhkYRyvYuno5NJuRWbkSJuOW9u
ogZH10m+EGA5DRhhiSBpkSga0uaQ7qmmI9OWjVVaIBqRIUhJCKZoAcOCz8WQV7Z3
k+URAXy0jsn7xLD06YGkmMDfOv5rXXxCvANL90NhbnNwfOjIfsIAPQGW9ZE0Ub+o
xdDwFKaMKhlp5VilbrjDLB6AunDSuTNMgOe3vbzjslFHyXaV+q6cFnTwfkFLV5VC
gg2MBYBNCbqYeNZcC1FFyuX9ExHSVxV/lbMiPNysxx/krqJ7TmMokeRycyota73z
4orFQP7euSpYJadGByT/G0U/f5XxSMKVtD40o1SbaX8fqAvPxvWFw8PqWJ+5JuqJ
qWiwH9dKWcldqPvvX33Ncv0r3RFz3EEvcHbWFUtYhrbAlMpchaWLWh7e3HfkdvI1
gM/Xm0oxgf+d3Dy6nGTjQ3MSV8HrV3hjWMumEZO2QSf0dj3DuZVmhmy081N3kg41
2DDO10fiRTrWpUxIEyC7/ir4+yJgm5VvJVMfkfjEMCu03MRiXQyPN8ilv9dSMcpZ
A7/rzGnZVNSkbW9kdiG2u5z4oRZ5XZDeEWq//QWPqyofM5YfeTN+VxJiZ3oxEBG9
+7trE0ySVp7WajwzW0B/FTaJFJ41ZS4q+QuZpNEDUIzXoXe/xgWnQYAkLHKx4Q1Y
8QpvkKlOfFVfdvTCi1dVOd3A0B1H3bOUc4EhqmaM8hxcekOPq2qSlyG+eImI1KsQ
vIPDDuBpuQ5gMClwkKcjSm4uuv/514ZP9396p4MG76QuY3wquDkt5M2tEzVapDAN
6xrkIRuIDGL34EffUHF1jsXdKfC/2aTyEFxjR9IPGAiAuyALI2XF/JQiBvwKAkfn
UPhYu+qeXPJRo04M3/drwwRIvbPTOBSXhXqmaSKPolPtPzm3uzucBO0BlJHUi/29
AGLqadW0O8NAoCt9rwwbHwMnCK3Td/Ifg99zQTKGuQlyK1u0aIjLIUI3IlGzfhgr
VbanbeXPX8As3qDJ4BRYCYmWZ+SBPm9eLqJ9PkhrF3CiptZ12nuLw5mQmqWpEk3x
oi2fLTOgyPOP74P/EJ/5pmxXwEIS/TNsArbBMji01vOWj0yJOFDnXs7E4944fn+x
4yiKKM1KrqLNMUFHukRoFW4WIezD8/j05ljdwVlR6tzXW7atOY3vN8QlpenB+2vQ
9kuAaBgeLJKsCEEEJtJ3344RUA/1yfNOdI12XWbAcQAd+DqIfgTn5LEqs7ta/haV
PnCdyn7vnVekAMrztHhcnEibg0Gfmuy8Az/c7sRdXZZA6mZrnrSTtg+68g3KFMOv
kNQfAoOy28DtDFSRaxlPah/nB97sonIK07tORbjVwTgcUHU1TZ/xNX1Qg0fvX7TZ
Kr7qdJ6JC/FtJbj1Py3O+JM94XjgeiVhhM5zu3DWCauMWX4F9KuZOkdlRHh2i+ji
cjTrsgFu672a++/qlN6xjpj7XE27lHoi/QtvPoLDI/VLxGnFBLdOe9U4RmX/1HFv
cgemNY5+TQnIB7lE8GYUF/mxiQoKeTLGSKa+gPrXZ04LJa36SUbdLrXd8QTE/NeW
F29gmKBZNKHpfSdttFk1GW7cvXhnZM+oX19z673nsavSPb6iYZX1EgjOJMO4b/Ue
fdP6/ioNj7wOuH9QfvvRjvguHqppptMwquVBksyHYiTVw82RgQsEMvCSqBCv7AuP
lN6guJspzxh97v+j8CaEou9DmT1OvnH1xG9TawXlxkEIhREeM51zis8d+lGRUVFS
wWPm8exPAIHfRLrLKkB11xgCQ/4LwWk5I2XrqpnpfHeUF82pN6e4MT7HZiIysM6P
n3w5zyv10Ko41ewPYRof+Dz5bOEpOYeS5fPz/3onwpm86mHt8fzpFOHF54ZZncJE
TXAGUFFlNExVfCvpk1gYOo36FthWCx3oWHNoJVbgX5Gii3kd3jQ3y+kdHqacon/S
JUZIlXJ8plEXG1n37SPzAGs8xOAGzloSKR6aYkE+yG3xpXI+LtdwSAep3oh452La
zhyyEcWqfLoF+tVroubawZ2hi+lIKEvhlhXQ/XzsA1e2DkAekwRKRX8T80rDTmvT
eSlZnCRGS1ePfBZ7JuqQirfl2MUN8JJsUUxbItLkkK+n0e6lL4DoDtxwz5UHHils
EmSmboayF06/Sq3u7axzrcO+Smi3S7scquG/f1AkwqJfGwilRf+sbWiWxgJ05FCr
//fmFLD4BQLKWFXnf81+v0Ndu3J/rrmnFRe0lsYl3DWiAxyKWjuWksDL1XkYKwYR
kNbSUAxnwzdjf8yrMx37oscOcjCm2Il2FHWEWU8eUoI4SgkXwfIJXmWW4IlwCsil
2p2A18B5l43Xm7+L6JQ/Sznu3l22DxBUxYeWczNMwhqdPu4/K37pq99i3tnA/2N5
vV0fWv38gx6cF+q8mxxBJDJxBc4z+EhzBqDVC59DXI9Zg6bAJyzz/GMFWM/ND1Ue
vCHY6IeSEmXwEWDlhnPG2Q==
`pragma protect end_protected
