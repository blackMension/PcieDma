`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bed5PGmfhMLhRR7yopyaPeq+S9PfUdOIVUVFks2pkl8l5keblO12aOq6lxkAXe8q
SVlVyeP4Y1H65G1S7XvkpIWbmDBY5bCi7WcmjETSUBgrcWAtaaRsNUWvniRIwTMu
CkpZIun3QH0NqHzLtQkdU9CFoR7cIZ9bm5iMcCyfg6Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
4XI3jYoy92G+f1oCeXLaJadOO+GzabeRby75Y4H2dqgi7OuOZMqnBar7vSdkhKDQ
d6kV44lclM+NexUPXw8iL9jwOe2mKyGvmOct1x1+SAKK9avQk4fIJ+X0K6rk/GZa
gT1er5m+pvbru2FEP19HE0iYtMx4+R80Mw40zlP8om7vDWyBrkknZx9IQjaJ43TH
2FXikjPt8kwhcFEgj/oJs4aJaqVVkV7KDsSuegzDg1MymlFpsxlklighlmQ5Mvrp
AVYV7FKbGtjxlYb6oNiPmp7qBXOw1wNk2SUGzlZXuR1AajmkrMi2H7MM4puqdtrN
711af7obYDAQVARPvkwIwqWHkjwdvqOoa45KHPDJnOGbkdchQSmmQTqLRiEYIvM8
/mpz9vqdBg7JsRNPxL3IGczRmi+mwzO5HBfIPD8CyKExE4ToTJlDTVxb+XPz4pz6
HTKS2ANITGLRVDTUKFfN3L4rn7kssDYP+qxYHI4/Y09J05QGfa1z7NgxabptAT2A
cyv2+KgLP+DA3QD84G5bAWXOn5FYolcYUjq69ouMoJ/gMSLttZMQmE0eOfuNvD7M
a87jsjlTYqLZNViGCtv8WGeDSU/SwBj1cUYVzONe1+sbBgynhEHF+QEsRDI0RT+R
BuL1B/GqR1g/6WhoXdC6hekrwgMwZzg5of+dEDGlN3oEoeEi3KAqUNk7irBv/iki
cXczwFtG3klK7ju23GdggLSL3yz0lZcnS+3GGMZBV2yMVRcEjVyXWXlM+v1la05S
1JkFNJxwEkkCp7A9EExhTmZVOt0LLo7I3jXRWdSGxJvjYc2o06okBKFxAVHnn/ZN
JsPs8TEju1a2hP5pskToihNszBkme9p3VnXcKjsdBB6CG/k+/tu4EH7scAFHaqmh
jripujTvzE74Vae2WOjKLc5ctCHvY/LXh7O/aEG/eE0/7IY2chFOvgmeGK3piO8u
M/vRPcL6xUJuLVee8NAZqfs2nYEfSnyazRfPTo+AmdF1nqEidHf166Eg2PwuzSXh
oGkn3Wz0cj3+GuDB5Fby0IGxrPiPOah2B7XEFmLzU5zjHYQuTBSBpHdVo8qQ9Nx0
4+DMn3mMDbAg9acVOBWZWiYnjRKHUdpL1lIl1eBKcs34MwFsJDpTky+FYrd9fZyC
MLfuRsjj5MwxygQyDC/SOUsBxY90vSLsBcWvGaDTDJhITTsMQeauSJnmCGOtTdBD
YPIlGWFgs1IP9H63hSN9sOAtjVLAkKBROMWUw6ZTUqxsIrxNceuzOy+t6zt/S4qQ
M6gECFlK9Bgr1Lv/pSb2SGU3WyF20NI8pZVEo2IYmyH9lIq0Hlw03oaGEiM6OZod
fiBCdACAzVV1gB75hpspheiDNxajyeo3NLyETgWkkuONUQXUA7TzCe/ZaZE/kvgG
niialsHfXE/SrV5dN5zgBELbg7tXe/nuts6Mywlt2/7UUQtCR4Miwa12pfwxqErw
CKZMpQE0ULnDZo520C9hhr7im4GrhqPSSOU+pSYxFPBcj48B97mXmX4LKl1khN44
vJNtmk97ELrEkV2CBh4C9hTgthpq7rO/881ttyaMgIj/9pcZ/IPLApApzSRpw6Po
1GwLJxhaJsmpb+TgkvwgAi42T7T6vZ6NjTmIRmk9op9TM/aX1hpwAKrjwirqvJoU
o0Mhk1WhLZ1L2kiJsbqr+IlaZyRE+fYRXqlRARqiGfSb+plsPpSnm7sZY6jhl/I3
qnz/5vfuSixVEN1jIK9g/BbCVfHFK0oA27wwwhXmSi90L4f5KULbx4oHOhAsdxkW
704aWHKKuVOoIsO3vmbh93NWeOBm9xaLH+l6p3lqudfL48JBUwZl2KVK9LDUTaht
kd5v1R9yFF8tAoJLD7rZhin8YVJa2FFvx6iFB7bb3TJ39j8e0baxE+aja5JQXfxx
7kMm9gwu8TT5EnqvVjDcxfFNPpnRdCzFAqx63Q5nPVJXzPU7bZyILB7IzlDNbNP6
C0YDnrTRgPypY+tzhf9ajOwLgkgxtjjGeQtaDi+WG6dIziPO5WhhqgnH97od1AuB
UDPMH3VvfOy6xXkVHR/E6ZbCZY+Ngru5f2dF9PyTRJcZydU6Um5mnxCOwSbTerB/
oHbbckhrcQvgMDE8/UTg9776XOuEC0VPLoBuTCxyG48uYbazZl4z3Xr4bWs2vKiN
xiZHdB5EINFgwIBw5DRt8io4q3ht/uwzUHsszBg6L/zNmg8K9c2lcfR4pgmEkcqI
naLb5AnJZCt3Nl8I8S4tGKtAqz8YpjlNO+/1fSvBSeVx00/p+HmY7bYS3s5GI7Po
W18Z0XzxzmVYvmJsnhTG98RNYPCPg3gDbJlj5QWiSWOe7+HI8/yaMmyDlO2B+b8n
r5OWn+9yuUd7ZQ/BUhCzvW1xyuZ2Xx1nZCbn71PgakqIVY2lQxex9oTx/bHVRJ/U
MiCUauw104dRmIukdIaZ1uQ/cc0l6x+Su54O4T372E9uTMQ65fgXhBtFPIWzGDeP
ZbYS/zLbJyRAEK1u47F/1IUAFVKzntnef8y3fi/IjzgKZcnsRLbwNOl5mXB431bE
qVtIgd4U+Fsa/xaJOnBF/sX5ay4vp9NrHE5QoaFbRZ/FmSzN9cbLxhXeJcjtTv4Z
05jhxtmk8+L17Yh12vXI+hXvUoiPkODiHZ6ygXKlLvhC9aUfuWi10Ud7TTETlGtO
P09n0eYvszKz5fYaQenobhrBPAmczp0/WPOzqN5z2lSdRGEaek6JDSwSwK2RNl5P
jtLo5etOaJMyeHOJI8swYTHaKeNRUL0F0vy4g+MqA+JgooWO8R7EClESCBRvJO9J
HhlteqMDuoScIZld3IqITuyBnmakVXWanAb/ycgDN0Cun0shSWEHu2eGyjJkmQuG
pHNW616Q8YeDQKjWrnSJ5U9yV2qTABZA/BnV3Qx2P+UHO33TM+eaha9RMqBIwbhv
l4K189Hg6XquZ5TQ5Fg41LoMzzjew/ZyAJzKKOOFZT+TaDFgJF759TriTbF9HlUf
QaDRBA0zRXybwsyl8znL0lFRWbyEQoW7J+zFOtf7OX7DsfC3GSKitwoQOGhzUpMr
YPLBb9MUN6l/j6boKR3Fo8sr1k5aFz+2zjcBiALZfUzHOD5jy/wPIqY2q94w4bwi
YLKqSsZZy+DguKWWU9VAf7QmrqQ6wkMoajFDJy/B9xpJyyzrhoTz41er6gU66fAI
3A2Bl3p5brf07uPz/pu0fMlZHTMlOBWY7sAhyLxkdDDxIRQcUnDKk3PJp/8bOhF6
8dK5HEi1ncUd0IJ3dv2jo01BPu/Kr5q/R6sTjrvWZjZnl/zB867XApsX/omBEuZy
5euxogY5LZvcKgLHGSe7VUkRphFEPOH0fm025K65N/6S0kdvLI2xbJyuf/7N8ly+
Moy71cMuTu0Gri4XbHA9Ajo6IMQmgG2ET1g0zWdJJ5EckRde5BOER7X9isggVO0J
UxC7yx+NqUbjtT7FU5U9cCfFTyjWXBGSetfNzicQ9xBJg8G0NCIlxMffLn2bT/TL
Htuu/+63ajUaCzr/j5O7sHINdPiIJ8wIgLkMDv7Sp16gKmQKmkcE9svnQe/H8T7p
BZpy5yGQvD66BLFXNUjWhpiJuqo9RtrGI8wXjpWp+beYNNYpTmMMAe5DzFY4ioq9
zT/fd/c3P3OAxyFmTAgpfF01+/iUKhy0tqvhHTid0Q9FSvBcwJ61EKtt9zAP2FUI
sOby5/ZERLt+qhKY3Ngi/e+eQZlaeMoCXKlfxv3LKQxSgLt3nksx4RJpNDtUXagB
+MRzehtmyXFaV5k13SvD+4dkLUxkAer/c1OMr/o+q/uaPjDyKhHIziaZkhiN/OBE
6yoY7IQBtGMOcqAfk5y7jwx8BTEQWx28+twpS+mNIwLsF8dwch5HPbGISEFKR0Gn
2RypAA6SoRVugDoIu0ZI4smgwCBb2y8th6ULv8/ojGMFXkQz1CppefR7ZGUQCNm1
149kQay28/9aluyfEHQcBHMLqd4wxQ/YVpL99vZbejCFipUMU7pH1BFjAsLej4ci
sGHG03jw7zP4+CxD2BrsrDitprZChTR9WWkkOxMzKfFCl+X9DBRs+hmzCxvlJyWP
g+gY1HnkLFcishnMSHfzzU3UdastRvRrBRg1/0SWIxh9bMkYw9Upbxk8U592mPvd
OQZcF6I5ZhPa5OebSyboqd4vKci86t1TAButw0wCpQ6lK3V2p7aIWpjQQpRQ4a0D
uI3zA1Fe+KVsM0WXvDRilLF3Jw1fHwzeOC1vdk/073iaG6M5A7vEUgylAZW4bMtl
SqVx/35SX7hxZs5Ow7R9+U++UJN8/cSL4LYzX8LLgcygZiOuHcg2JFTN2XNiCn+0
7+uOJLv0CltzHrfQGeG+p8ySKfMu6wx6+m2LBlON6wqDSSJq4kK9N1hlhgwBq7l/
HwKsLe72s6C05Z9A9JVzKn8jLKUI07KNYvWZjMrQn6BoAqpiXnzLzQPRwysu3Z0b
iKk9pleeDE+tv2iyJKloDTyLTGn+kIPwfmL6bWiRdZutjWwkAyY6+Pe/1zu46mSL
Z1Pf05JHmpEE2uswOzgxIijXU5L1sX5PQ9tQWHUmpeET9mzz/pd0be1biqcQ5GHo
VQnBMb3pQuDJ8xVru8UWGusclBHZD/L6k89R+ZFNj3Ai7dXNMooOIKwQC1+LDF2c
3cwHeevMMV/ms97BJBEItiy956+UIU18J0JAm1c7E8cCUpe90SdEvbVggBtVjv5/
+eyyofKhbChhDOJ5xtEzI5H2cc8Nq+W35naWZOsFQEPu9mLewfXHt1Zs9Eirf5nK
HKA/U7vaOWhmQUFT9NSpvTtEkVztgsC/AitkaAjkbi2EK8+acSmJJDMYvI+kW1Rt
lGPF7EIJSVJGrd9kmM22k2L2OFeP++YmeC5/gR73wUjc0BjrMpxa89sa1hOhDreS
AgWJrLRd0QHnXKHvZjthOUkJYINtrwNOSUGz7nppzvbhMXJ19hzVPv6/TcnYDBw1
7ZlXoHoIUhnD0lZguyuh0jyD+k0ZCtu7yF03ijpBv8q/765oTOgOIxm5AD3npku7
ZMyTKteWto0bNsS/Ku5E0GfMNjvRr3Fp40JX6TGm1XPT0UrOyVWdQaaDCVIwGNM9
jgkIYQdDz80315XhQ/wMZ8L8ShAttGK7H5F0KdlmN1niwQdTNbP6FP/vZd5Dvv9v
5XB0IPQMe68OOysNLGFAr1DjcYRq+92s6I2j56K2A2cfQnQwR0rKVvj3jJ+8M8c9
mO+4iMKR6uMCLBYgdvhTzzx3MQkNfeGlXb6TOun0cZ3ZLYrmm8YNWz7siMWfl/jA
8hlIMO4oQNs7OPyMQM558s4ybvi08Z9J1bMuAuyxKuh6UNFpAip9qdf4a/Ggt63o
x8cWTptmiMb5N2q1EoTr0zaX9C8wcmEeKs6QnlljXtDLEeln6NoBCVw4MC8DR4PK
YX7M+5dzxyUDQUc7K4gM9/7ioiRnIX8Vs3Vt3x9Mfd2/5CJQWgWPbxQJBJCiCjz/
qHP134dQfgAHNQAKn6jtykSWir1cqz1MK8JuEaSMEjNaQdZ9l5xbZTtND/b9HLBN
oEWY8Kq+DtFojilNdAQhHiocejZd77aPhGn9QaZrIEJzhgV0e7pIsctMadYET7Dj
acCd1MbfMu348ZrxS0Ire7vUIayFgPWTa86R0KasC97vAc6RjNYXKKYFnSFOsM2y
8LNLf3luzRU1I3eOSP4M8RA9hTT3QmKB7U8h537yHk1g3O5KCMkSQY26iSg+Hc39
qc93T1ta0t8VOV1KKPtkUP18I3YdEdVLSnbM00sW7PK4jPc3y4dwKjJZqkfyZIH5
mz7q4yG9VC9el0YRAmrkPzkr4D3SWZYyI+TG+U3Le3fwMhJbOaPvj3vNsVbN4bgq
3kpNVHGxAfNtLubqJg7BojXstyqPN3FgZOXLfpdO7ykVvdsXfn/CTZIOKeNGjPCJ
wzIFq4umsR8xQ4XWBh0S03ydgOlqqSeUUJ1pEaarIOWT6FXq43CuOWY3k0pRhILO
//N3e2Xz0wBfMGiSCg95bmO1QCdKnGfTMcmSvvEyaQ1qLlI6RkCbhUmzzvpZCgcL
RQUvbTeUndSTgGULvA//MPbTcjQpHnVHOfMgdbtMPWHqFUpI2wNMFlEBqLV5eovn
5mWzG+2q+06XwyKvL1k291cOLJ9mClIHmYAqBav+Q8OBKRQ5sCAb0maF9MgcspHf
SEOcUnRSjcQxfArRU/zDebyVCWpQ1+N7LDgkIZ9N0hm0b3KgHGaXXXExrWrBnK0N
n6E8eLoEyttDrtQXymRAWMGb5aDKba8FKuGRais66g/V0PiyOUNag7Vl2v1j2ozb
VafY15BuG/HbQmd0j3cHrPu+iXkuxhlu8jBkfX5ywg/wO2BJUyms/rG3lPpORkJA
lWKYUoafaOsGKcAQ9dPlArGiGoCBh5zO5HhEsxb+R/3QsTjjJEqiwIolBWMeBvSD
nuFhFAjvpSAAcud0HVsk+JGc/bQCwO8XbbwFn4cOLdE/h6aBMudVRFborWYqufnS
Psg37ff0FnbWgpcBNzOAQnkDtluLL8X201vdKAcKF3y4YI+VuBFCYTnM8DbDYGkb
iC3765ax53nG1Xo4zp4eAn9Ouq5ReMXU07NsiOVV9u10FT99eLFLoc3OCyzsTv7D
oW24HRTDV83PxanuhZXmU1ykTJPPdzlId0ZglqL1/f58e8F8zR6KgPGBwoioMugS
tQEyx2ZCbyNvz/SBIBF/39TFCrgsh7LmIv5WYtCP86AdadCTU6QKF9yCW9MSt+J7
nYd4O+/7CDNjnAGCKarmFFESUnN/FDVSYFZwKXgr30vJzVdXA2zbacPUxnL5N7HM
DjHD4r2MWwNCjV1BLOQ+EMGgSHMNdFTpGjbcsds1sq4NXldKnPOOVcV9XjK+ywbo
VQpMMXFsfol98PSVCvLBCo7Gp5X+72DwMLkDosLdKBLJFAgxxvOAij3hGsfMNGeZ
KFahiyAPOP/vERca1Hcap6iObu2zhb8T2kqDlSPQsVIETxt1c5Kvc6FF7SH6wg4y
H9LpfAcNAkM77n1N71SjYYq487arLq8JT36w2uiUQ5kvcQPbI56qk+Sw4ztcKNbl
WCiEs2JA7SaRHJ3q/OT2Y4IMQ/PAwNRqNagA+oAxKEJ/Bo0gOGQA+Q6R1i930g9c
M2LH/RxqDRe1Zvc65GgGya3rQGAi/3AdqAP1fXqn6mclESFkEM9cNXU3ERxtm4j0
kQ9iNsk9LAiG6yfSqA0Lw3aAanzL8kiu4cd3wI7visLA9Lw+5WkvaXEsluFIdbvi
OmrQYuou4ZDS6naILC1r4OmQlhol6YqYHJh9Lgf+ShXl97aKGPEFSRyBHUrh85gU
1MOK8/l7VI90z/LBfvWWWwNuBLVFEwpVcvF7SAKxFIwbD5kyvO0bYkdFdYeDqq+2
HSoHHnIU6LXFjH88a4cvNhnePPaRY8T9DHR0H8avi5PlBPS2IxO7ZrBgLaw66ceH
yOisD4jS7lsHIU/T6UJC00DGDPXNnt6eHUx0nuI7aMaV9IG8qAm6n10hetOrsxfB
`pragma protect end_protected
