// lcpll_g3xn.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module lcpll_g3xn #(
		parameter enable_pll_reconfig                                              = 1,
		parameter rcfg_jtag_enable                                                 = 0,
		parameter rcfg_separate_avmm_busy                                          = 0,
		parameter dbg_embedded_debug_enable                                        = 0,
		parameter dbg_capability_reg_enable                                        = 0,
		parameter dbg_user_identifier                                              = 0,
		parameter dbg_stat_soft_logic_enable                                       = 0,
		parameter dbg_ctrl_soft_logic_enable                                       = 0,
		parameter rcfg_emb_strm_enable                                             = 0,
		parameter rcfg_profile_cnt                                                 = 2,
		parameter hssi_pma_lc_refclk_select_mux_powerdown_mode                     = "powerup",
		parameter hssi_pma_lc_refclk_select_mux_refclk_select                      = "ref_iqclk0",
		parameter hssi_pma_lc_refclk_select_mux_silicon_rev                        = "20nm5",
		parameter hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping = "ref_iqclk0",
		parameter hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping = "power_down",
		parameter hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping = "power_down",
		parameter hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping = "power_down",
		parameter hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping = "power_down",
		parameter hssi_refclk_divider_silicon_rev                                  = "20nm5",
		parameter atx_pll_silicon_rev                                              = "20nm5",
		parameter atx_pll_is_cascaded_pll                                          = "false",
		parameter atx_pll_cgb_div                                                  = 1,
		parameter atx_pll_pma_width                                                = 32,
		parameter atx_pll_cp_compensation_enable                                   = "true",
		parameter atx_pll_cp_current_setting                                       = "cp_current_setting26",
		parameter atx_pll_cp_testmode                                              = "cp_normal",
		parameter atx_pll_cp_lf_3rd_pole_freq                                      = "lf_3rd_pole_setting0",
		parameter atx_pll_lf_cbig_size                                             = "lf_cbig_setting4",
		parameter atx_pll_cp_lf_order                                              = "lf_3rd_order",
		parameter atx_pll_lf_resistance                                            = "lf_setting1",
		parameter atx_pll_lf_ripplecap                                             = "lf_ripple_cap_0",
		parameter atx_pll_tank_sel                                                 = "lctank0",
		parameter atx_pll_tank_band                                                = "lc_band3",
		parameter atx_pll_tank_voltage_coarse                                      = "vreg_setting_coarse0",
		parameter atx_pll_tank_voltage_fine                                        = "vreg_setting5",
		parameter atx_pll_output_regulator_supply                                  = "vreg1v_setting0",
		parameter atx_pll_overrange_voltage                                        = "over_setting0",
		parameter atx_pll_underrange_voltage                                       = "under_setting4",
		parameter atx_pll_fb_select                                                = "direct_fb",
		parameter atx_pll_d2a_voltage                                              = "d2a_setting_4",
		parameter atx_pll_dsm_mode                                                 = "dsm_mode_integer",
		parameter atx_pll_dsm_out_sel                                              = "pll_dsm_disable",
		parameter atx_pll_dsm_ecn_bypass                                           = "false",
		parameter atx_pll_dsm_ecn_test_en                                          = "false",
		parameter atx_pll_dsm_fractional_division                                  = "1",
		parameter atx_pll_dsm_fractional_value_ready                               = "pll_k_ready",
		parameter atx_pll_iqclk_mux_sel                                            = "iqtxrxclk0",
		parameter atx_pll_vco_bypass_enable                                        = "false",
		parameter atx_pll_l_counter                                                = 2,
		parameter atx_pll_l_counter_enable                                         = "true",
		parameter atx_pll_cascadeclk_test                                          = "cascadetest_off",
		parameter atx_pll_hclk_divide                                              = 50,
		parameter atx_pll_enable_hclk                                              = "hclk_disabled",
		parameter atx_pll_m_counter                                                = 40,
		parameter atx_pll_ref_clk_div                                              = 1,
		parameter atx_pll_bw_sel                                                   = "high",
		parameter atx_pll_datarate                                                 = "8000000000 bps",
		parameter atx_pll_device_variant                                           = "device1",
		parameter atx_pll_initial_settings                                         = "true",
		parameter atx_pll_lc_mode                                                  = "lccmu_normal",
		parameter atx_pll_output_clock_frequency                                   = "4000000000 Hz",
		parameter atx_pll_powerdown_mode                                           = "powerup",
		parameter atx_pll_prot_mode                                                = "pcie_gen3_tx",
		parameter atx_pll_reference_clock_frequency                                = "100000000 Hz",
		parameter atx_pll_sup_mode                                                 = "user_mode",
		parameter atx_pll_regulator_bypass                                         = "reg_enable",
		parameter atx_pll_vco_freq                                                 = "8000000000 Hz",
		parameter atx_pll_is_otn                                                   = "false",
		parameter atx_pll_is_sdi                                                   = "false",
		parameter atx_pll_primary_use                                              = "hssi_x1",
		parameter atx_pll_fpll_refclk_selection                                    = "select_vco_output",
		parameter atx_pll_lc_to_fpll_l_counter_scratch                             = 1,
		parameter atx_pll_lc_to_fpll_l_counter                                     = "lcounter_setting0",
		parameter atx_pll_pfd_delay_compensation                                   = "normal_delay",
		parameter atx_pll_xcpvco_xchgpmplf_cp_current_boost                        = "normal_setting",
		parameter atx_pll_pfd_pulse_width                                          = "pulse_width_setting0",
		parameter hip_cal_en                                                       = "enable",
		parameter calibration_en                                                   = "enable",
		parameter enable_analog_resets                                             = 0,
		parameter atx_pll_bonding_mode                                             = "cpri_bonding",
		parameter enable_mcgb                                                      = 1,
		parameter enable_mcgb_debug_ports_parameters                               = 0,
		parameter hssi_pma_cgb_master_prot_mode                                    = "pcie_gen3_tx",
		parameter hssi_pma_cgb_master_silicon_rev                                  = "20nm5",
		parameter hssi_pma_cgb_master_x1_div_m_sel                                 = "divbypass",
		parameter hssi_pma_cgb_master_cgb_enable_iqtxrxclk                         = "disable_iqtxrxclk",
		parameter hssi_pma_cgb_master_ser_mode                                     = "thirty_two_bit",
		parameter hssi_pma_cgb_master_datarate                                     = "8000000000 bps",
		parameter hssi_pma_cgb_master_cgb_power_down                               = "normal_cgb",
		parameter hssi_pma_cgb_master_observe_cgb_clocks                           = "observe_nothing",
		parameter hssi_pma_cgb_master_op_mode                                      = "enabled",
		parameter hssi_pma_cgb_master_tx_ucontrol_reset_pcie                       = "pcscorehip_controls_mcgb",
		parameter hssi_pma_cgb_master_vccdreg_output                               = "vccdreg_nominal",
		parameter hssi_pma_cgb_master_input_select                                 = "fpll_top",
		parameter hssi_pma_cgb_master_input_select_gen3                            = "lcpll_top"
	) (
		input  wire        pll_powerdown,         //     pll_powerdown.pll_powerdown
		input  wire        pll_refclk0,           //       pll_refclk0.clk
		output wire        pll_locked,            //        pll_locked.pll_locked
		output wire        pll_pcie_clk,          //      pll_pcie_clk.pll_pcie_clk
		input  wire        reconfig_clk0,         //     reconfig_clk0.clk
		input  wire        reconfig_reset0,       //   reconfig_reset0.reset
		input  wire        reconfig_write0,       //    reconfig_avmm0.write
		input  wire        reconfig_read0,        //                  .read
		input  wire [9:0]  reconfig_address0,     //                  .address
		input  wire [31:0] reconfig_writedata0,   //                  .writedata
		output wire [31:0] reconfig_readdata0,    //                  .readdata
		output wire        reconfig_waitrequest0, //                  .waitrequest
		output wire        pll_cal_busy,          //      pll_cal_busy.pll_cal_busy
		output wire        hip_cal_done,          //      hip_cal_done.hip_cal_done
		input  wire        mcgb_rst,              //          mcgb_rst.mcgb_rst
		input  wire        mcgb_aux_clk0,         //     mcgb_aux_clk0.tx_serial_clk
		output wire [5:0]  tx_bonding_clocks,     // tx_bonding_clocks.clk
		input  wire [1:0]  pcie_sw,               //           pcie_sw.pcie_sw
		output wire [1:0]  pcie_sw_done,          //      pcie_sw_done.pcie_sw_done
		output wire        mcgb_hip_cal_done      // mcgb_hip_cal_done.hip_cal_done
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (enable_pll_reconfig != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_pll_reconfig_check ( .error(1'b1) );
		end
		if (rcfg_jtag_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_jtag_enable_check ( .error(1'b1) );
		end
		if (rcfg_separate_avmm_busy != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_separate_avmm_busy_check ( .error(1'b1) );
		end
		if (dbg_embedded_debug_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_embedded_debug_enable_check ( .error(1'b1) );
		end
		if (dbg_capability_reg_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_capability_reg_enable_check ( .error(1'b1) );
		end
		if (dbg_user_identifier != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_user_identifier_check ( .error(1'b1) );
		end
		if (dbg_stat_soft_logic_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_stat_soft_logic_enable_check ( .error(1'b1) );
		end
		if (dbg_ctrl_soft_logic_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					dbg_ctrl_soft_logic_enable_check ( .error(1'b1) );
		end
		if (rcfg_emb_strm_enable != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_emb_strm_enable_check ( .error(1'b1) );
		end
		if (rcfg_profile_cnt != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					rcfg_profile_cnt_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_powerdown_mode_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_refclk_select != "ref_iqclk0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_refclk_select_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_silicon_rev != "20nm5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping != "ref_iqclk0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping != "power_down")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping != "power_down")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping != "power_down")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping_check ( .error(1'b1) );
		end
		if (hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping != "power_down")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping_check ( .error(1'b1) );
		end
		if (hssi_refclk_divider_silicon_rev != "20nm5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_refclk_divider_silicon_rev_check ( .error(1'b1) );
		end
		if (atx_pll_silicon_rev != "20nm5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_silicon_rev_check ( .error(1'b1) );
		end
		if (atx_pll_is_cascaded_pll != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_is_cascaded_pll_check ( .error(1'b1) );
		end
		if (atx_pll_cgb_div != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cgb_div_check ( .error(1'b1) );
		end
		if (atx_pll_pma_width != 32)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_pma_width_check ( .error(1'b1) );
		end
		if (atx_pll_cp_compensation_enable != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cp_compensation_enable_check ( .error(1'b1) );
		end
		if (atx_pll_cp_current_setting != "cp_current_setting26")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cp_current_setting_check ( .error(1'b1) );
		end
		if (atx_pll_cp_testmode != "cp_normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cp_testmode_check ( .error(1'b1) );
		end
		if (atx_pll_cp_lf_3rd_pole_freq != "lf_3rd_pole_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cp_lf_3rd_pole_freq_check ( .error(1'b1) );
		end
		if (atx_pll_lf_cbig_size != "lf_cbig_setting4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lf_cbig_size_check ( .error(1'b1) );
		end
		if (atx_pll_cp_lf_order != "lf_3rd_order")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cp_lf_order_check ( .error(1'b1) );
		end
		if (atx_pll_lf_resistance != "lf_setting1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lf_resistance_check ( .error(1'b1) );
		end
		if (atx_pll_lf_ripplecap != "lf_ripple_cap_0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lf_ripplecap_check ( .error(1'b1) );
		end
		if (atx_pll_tank_sel != "lctank0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_tank_sel_check ( .error(1'b1) );
		end
		if (atx_pll_tank_band != "lc_band3")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_tank_band_check ( .error(1'b1) );
		end
		if (atx_pll_tank_voltage_coarse != "vreg_setting_coarse0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_tank_voltage_coarse_check ( .error(1'b1) );
		end
		if (atx_pll_tank_voltage_fine != "vreg_setting5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_tank_voltage_fine_check ( .error(1'b1) );
		end
		if (atx_pll_output_regulator_supply != "vreg1v_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_output_regulator_supply_check ( .error(1'b1) );
		end
		if (atx_pll_overrange_voltage != "over_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_overrange_voltage_check ( .error(1'b1) );
		end
		if (atx_pll_underrange_voltage != "under_setting4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_underrange_voltage_check ( .error(1'b1) );
		end
		if (atx_pll_fb_select != "direct_fb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_fb_select_check ( .error(1'b1) );
		end
		if (atx_pll_d2a_voltage != "d2a_setting_4")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_d2a_voltage_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_mode != "dsm_mode_integer")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_mode_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_out_sel != "pll_dsm_disable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_out_sel_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_ecn_bypass != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_ecn_bypass_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_ecn_test_en != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_ecn_test_en_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_fractional_division != "1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_fractional_division_check ( .error(1'b1) );
		end
		if (atx_pll_dsm_fractional_value_ready != "pll_k_ready")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_dsm_fractional_value_ready_check ( .error(1'b1) );
		end
		if (atx_pll_iqclk_mux_sel != "iqtxrxclk0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_iqclk_mux_sel_check ( .error(1'b1) );
		end
		if (atx_pll_vco_bypass_enable != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_vco_bypass_enable_check ( .error(1'b1) );
		end
		if (atx_pll_l_counter != 2)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_l_counter_check ( .error(1'b1) );
		end
		if (atx_pll_l_counter_enable != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_l_counter_enable_check ( .error(1'b1) );
		end
		if (atx_pll_cascadeclk_test != "cascadetest_off")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_cascadeclk_test_check ( .error(1'b1) );
		end
		if (atx_pll_hclk_divide != 50)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_hclk_divide_check ( .error(1'b1) );
		end
		if (atx_pll_enable_hclk != "hclk_disabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_enable_hclk_check ( .error(1'b1) );
		end
		if (atx_pll_m_counter != 40)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_m_counter_check ( .error(1'b1) );
		end
		if (atx_pll_ref_clk_div != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_ref_clk_div_check ( .error(1'b1) );
		end
		if (atx_pll_bw_sel != "high")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_bw_sel_check ( .error(1'b1) );
		end
		if (atx_pll_datarate != "8000000000 bps")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_datarate_check ( .error(1'b1) );
		end
		if (atx_pll_device_variant != "device1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_device_variant_check ( .error(1'b1) );
		end
		if (atx_pll_initial_settings != "true")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_initial_settings_check ( .error(1'b1) );
		end
		if (atx_pll_lc_mode != "lccmu_normal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lc_mode_check ( .error(1'b1) );
		end
		if (atx_pll_output_clock_frequency != "4000000000 Hz")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_output_clock_frequency_check ( .error(1'b1) );
		end
		if (atx_pll_powerdown_mode != "powerup")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_powerdown_mode_check ( .error(1'b1) );
		end
		if (atx_pll_prot_mode != "pcie_gen3_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_prot_mode_check ( .error(1'b1) );
		end
		if (atx_pll_reference_clock_frequency != "100000000 Hz")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_reference_clock_frequency_check ( .error(1'b1) );
		end
		if (atx_pll_sup_mode != "user_mode")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_sup_mode_check ( .error(1'b1) );
		end
		if (atx_pll_regulator_bypass != "reg_enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_regulator_bypass_check ( .error(1'b1) );
		end
		if (atx_pll_vco_freq != "8000000000 Hz")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_vco_freq_check ( .error(1'b1) );
		end
		if (atx_pll_is_otn != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_is_otn_check ( .error(1'b1) );
		end
		if (atx_pll_is_sdi != "false")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_is_sdi_check ( .error(1'b1) );
		end
		if (atx_pll_primary_use != "hssi_x1")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_primary_use_check ( .error(1'b1) );
		end
		if (atx_pll_fpll_refclk_selection != "select_vco_output")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_fpll_refclk_selection_check ( .error(1'b1) );
		end
		if (atx_pll_lc_to_fpll_l_counter_scratch != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lc_to_fpll_l_counter_scratch_check ( .error(1'b1) );
		end
		if (atx_pll_lc_to_fpll_l_counter != "lcounter_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_lc_to_fpll_l_counter_check ( .error(1'b1) );
		end
		if (atx_pll_pfd_delay_compensation != "normal_delay")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_pfd_delay_compensation_check ( .error(1'b1) );
		end
		if (atx_pll_xcpvco_xchgpmplf_cp_current_boost != "normal_setting")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_xcpvco_xchgpmplf_cp_current_boost_check ( .error(1'b1) );
		end
		if (atx_pll_pfd_pulse_width != "pulse_width_setting0")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_pfd_pulse_width_check ( .error(1'b1) );
		end
		if (hip_cal_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hip_cal_en_check ( .error(1'b1) );
		end
		if (calibration_en != "enable")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					calibration_en_check ( .error(1'b1) );
		end
		if (enable_analog_resets != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_analog_resets_check ( .error(1'b1) );
		end
		if (atx_pll_bonding_mode != "cpri_bonding")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					atx_pll_bonding_mode_check ( .error(1'b1) );
		end
		if (enable_mcgb != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_mcgb_check ( .error(1'b1) );
		end
		if (enable_mcgb_debug_ports_parameters != 0)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					enable_mcgb_debug_ports_parameters_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_prot_mode != "pcie_gen3_tx")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_prot_mode_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_silicon_rev != "20nm5")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_silicon_rev_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_x1_div_m_sel != "divbypass")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_x1_div_m_sel_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_cgb_enable_iqtxrxclk != "disable_iqtxrxclk")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_cgb_enable_iqtxrxclk_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_ser_mode != "thirty_two_bit")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_ser_mode_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_datarate != "8000000000 bps")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_datarate_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_cgb_power_down != "normal_cgb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_cgb_power_down_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_observe_cgb_clocks != "observe_nothing")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_observe_cgb_clocks_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_op_mode != "enabled")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_op_mode_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_tx_ucontrol_reset_pcie != "pcscorehip_controls_mcgb")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_tx_ucontrol_reset_pcie_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_vccdreg_output != "vccdreg_nominal")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_vccdreg_output_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_input_select != "fpll_top")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_input_select_check ( .error(1'b1) );
		end
		if (hssi_pma_cgb_master_input_select_gen3 != "lcpll_top")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					hssi_pma_cgb_master_input_select_gen3_check ( .error(1'b1) );
		end
	endgenerate

	ep_g3x8_avmm256_DUT_altera_xcvr_atx_pll_a10_171_pufnv4i #(
		.enable_pll_reconfig                                              (1),
		.rcfg_jtag_enable                                                 (0),
		.rcfg_separate_avmm_busy                                          (0),
		.dbg_embedded_debug_enable                                        (0),
		.dbg_capability_reg_enable                                        (0),
		.dbg_user_identifier                                              (0),
		.dbg_stat_soft_logic_enable                                       (0),
		.dbg_ctrl_soft_logic_enable                                       (0),
		.rcfg_emb_strm_enable                                             (0),
		.rcfg_profile_cnt                                                 (2),
		.hssi_pma_lc_refclk_select_mux_powerdown_mode                     ("powerup"),
		.hssi_pma_lc_refclk_select_mux_refclk_select                      ("ref_iqclk0"),
		.hssi_pma_lc_refclk_select_mux_silicon_rev                        ("20nm5"),
		.hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping ("ref_iqclk0"),
		.hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping ("power_down"),
		.hssi_refclk_divider_silicon_rev                                  ("20nm5"),
		.atx_pll_silicon_rev                                              ("20nm5"),
		.atx_pll_is_cascaded_pll                                          ("false"),
		.atx_pll_cgb_div                                                  (1),
		.atx_pll_pma_width                                                (32),
		.atx_pll_cp_compensation_enable                                   ("true"),
		.atx_pll_cp_current_setting                                       ("cp_current_setting26"),
		.atx_pll_cp_testmode                                              ("cp_normal"),
		.atx_pll_cp_lf_3rd_pole_freq                                      ("lf_3rd_pole_setting0"),
		.atx_pll_lf_cbig_size                                             ("lf_cbig_setting4"),
		.atx_pll_cp_lf_order                                              ("lf_3rd_order"),
		.atx_pll_lf_resistance                                            ("lf_setting1"),
		.atx_pll_lf_ripplecap                                             ("lf_ripple_cap_0"),
		.atx_pll_tank_sel                                                 ("lctank0"),
		.atx_pll_tank_band                                                ("lc_band3"),
		.atx_pll_tank_voltage_coarse                                      ("vreg_setting_coarse0"),
		.atx_pll_tank_voltage_fine                                        ("vreg_setting5"),
		.atx_pll_output_regulator_supply                                  ("vreg1v_setting0"),
		.atx_pll_overrange_voltage                                        ("over_setting0"),
		.atx_pll_underrange_voltage                                       ("under_setting4"),
		.atx_pll_fb_select                                                ("direct_fb"),
		.atx_pll_d2a_voltage                                              ("d2a_setting_4"),
		.atx_pll_dsm_mode                                                 ("dsm_mode_integer"),
		.atx_pll_dsm_out_sel                                              ("pll_dsm_disable"),
		.atx_pll_dsm_ecn_bypass                                           ("false"),
		.atx_pll_dsm_ecn_test_en                                          ("false"),
		.atx_pll_dsm_fractional_division                                  ("1"),
		.atx_pll_dsm_fractional_value_ready                               ("pll_k_ready"),
		.atx_pll_iqclk_mux_sel                                            ("iqtxrxclk0"),
		.atx_pll_vco_bypass_enable                                        ("false"),
		.atx_pll_l_counter                                                (2),
		.atx_pll_l_counter_enable                                         ("true"),
		.atx_pll_cascadeclk_test                                          ("cascadetest_off"),
		.atx_pll_hclk_divide                                              (50),
		.atx_pll_enable_hclk                                              ("hclk_disabled"),
		.atx_pll_m_counter                                                (40),
		.atx_pll_ref_clk_div                                              (1),
		.atx_pll_bw_sel                                                   ("high"),
		.atx_pll_datarate                                                 ("8000000000 bps"),
		.atx_pll_device_variant                                           ("device1"),
		.atx_pll_initial_settings                                         ("true"),
		.atx_pll_lc_mode                                                  ("lccmu_normal"),
		.atx_pll_output_clock_frequency                                   ("4000000000 Hz"),
		.atx_pll_powerdown_mode                                           ("powerup"),
		.atx_pll_prot_mode                                                ("pcie_gen3_tx"),
		.atx_pll_reference_clock_frequency                                ("100000000 Hz"),
		.atx_pll_sup_mode                                                 ("user_mode"),
		.atx_pll_regulator_bypass                                         ("reg_enable"),
		.atx_pll_vco_freq                                                 ("8000000000 Hz"),
		.atx_pll_is_otn                                                   ("false"),
		.atx_pll_is_sdi                                                   ("false"),
		.atx_pll_primary_use                                              ("hssi_x1"),
		.atx_pll_fpll_refclk_selection                                    ("select_vco_output"),
		.atx_pll_lc_to_fpll_l_counter_scratch                             (1),
		.atx_pll_lc_to_fpll_l_counter                                     ("lcounter_setting0"),
		.atx_pll_pfd_delay_compensation                                   ("normal_delay"),
		.atx_pll_xcpvco_xchgpmplf_cp_current_boost                        ("normal_setting"),
		.atx_pll_pfd_pulse_width                                          ("pulse_width_setting0"),
		.hip_cal_en                                                       ("enable"),
		.calibration_en                                                   ("enable"),
		.enable_analog_resets                                             (0),
		.atx_pll_bonding_mode                                             ("cpri_bonding"),
		.enable_mcgb                                                      (1),
		.enable_mcgb_debug_ports_parameters                               (0),
		.hssi_pma_cgb_master_prot_mode                                    ("pcie_gen3_tx"),
		.hssi_pma_cgb_master_silicon_rev                                  ("20nm5"),
		.hssi_pma_cgb_master_x1_div_m_sel                                 ("divbypass"),
		.hssi_pma_cgb_master_cgb_enable_iqtxrxclk                         ("disable_iqtxrxclk"),
		.hssi_pma_cgb_master_ser_mode                                     ("thirty_two_bit"),
		.hssi_pma_cgb_master_datarate                                     ("8000000000 bps"),
		.hssi_pma_cgb_master_cgb_power_down                               ("normal_cgb"),
		.hssi_pma_cgb_master_observe_cgb_clocks                           ("observe_nothing"),
		.hssi_pma_cgb_master_op_mode                                      ("enabled"),
		.hssi_pma_cgb_master_tx_ucontrol_reset_pcie                       ("pcscorehip_controls_mcgb"),
		.hssi_pma_cgb_master_vccdreg_output                               ("vccdreg_nominal"),
		.hssi_pma_cgb_master_input_select                                 ("fpll_top"),
		.hssi_pma_cgb_master_input_select_gen3                            ("lcpll_top")
	) lcpll_g3xn (
		.pll_powerdown           (pll_powerdown),                        //   input,   width = 1,     pll_powerdown.pll_powerdown
		.pll_refclk0             (pll_refclk0),                          //   input,   width = 1,       pll_refclk0.clk
		.pll_locked              (pll_locked),                           //  output,   width = 1,        pll_locked.pll_locked
		.pll_pcie_clk            (pll_pcie_clk),                         //  output,   width = 1,      pll_pcie_clk.pll_pcie_clk
		.reconfig_clk0           (reconfig_clk0),                        //   input,   width = 1,     reconfig_clk0.clk
		.reconfig_reset0         (reconfig_reset0),                      //   input,   width = 1,   reconfig_reset0.reset
		.reconfig_write0         (reconfig_write0),                      //   input,   width = 1,    reconfig_avmm0.write
		.reconfig_read0          (reconfig_read0),                       //   input,   width = 1,                  .read
		.reconfig_address0       (reconfig_address0),                    //   input,  width = 10,                  .address
		.reconfig_writedata0     (reconfig_writedata0),                  //   input,  width = 32,                  .writedata
		.reconfig_readdata0      (reconfig_readdata0),                   //  output,  width = 32,                  .readdata
		.reconfig_waitrequest0   (reconfig_waitrequest0),                //  output,   width = 1,                  .waitrequest
		.pll_cal_busy            (pll_cal_busy),                         //  output,   width = 1,      pll_cal_busy.pll_cal_busy
		.hip_cal_done            (hip_cal_done),                         //  output,   width = 1,      hip_cal_done.hip_cal_done
		.mcgb_rst                (mcgb_rst),                             //   input,   width = 1,          mcgb_rst.mcgb_rst
		.mcgb_aux_clk0           (mcgb_aux_clk0),                        //   input,   width = 1,     mcgb_aux_clk0.tx_serial_clk
		.tx_bonding_clocks       (tx_bonding_clocks),                    //  output,   width = 6, tx_bonding_clocks.clk
		.pcie_sw                 (pcie_sw),                              //   input,   width = 2,           pcie_sw.pcie_sw
		.pcie_sw_done            (pcie_sw_done),                         //  output,   width = 2,      pcie_sw_done.pcie_sw_done
		.mcgb_hip_cal_done       (mcgb_hip_cal_done),                    //  output,   width = 1, mcgb_hip_cal_done.hip_cal_done
		.pll_refclk1             (1'b0),                                 // (terminated),                                
		.pll_refclk2             (1'b0),                                 // (terminated),                                
		.pll_refclk3             (1'b0),                                 // (terminated),                                
		.pll_refclk4             (1'b0),                                 // (terminated),                                
		.tx_serial_clk           (),                                     // (terminated),                                
		.tx_serial_clk_gt        (),                                     // (terminated),                                
		.pll_cascade_clk         (),                                     // (terminated),                                
		.atx_to_fpll_cascade_clk (),                                     // (terminated),                                
		.avmm_busy0              (),                                     // (terminated),                                
		.clklow                  (),                                     // (terminated),                                
		.fref                    (),                                     // (terminated),                                
		.overrange               (),                                     // (terminated),                                
		.underrange              (),                                     // (terminated),                                
		.mcgb_aux_clk1           (1'b0),                                 // (terminated),                                
		.mcgb_aux_clk2           (1'b0),                                 // (terminated),                                
		.mcgb_serial_clk         (),                                     // (terminated),                                
		.reconfig_clk1           (1'b0),                                 // (terminated),                                
		.reconfig_reset1         (1'b0),                                 // (terminated),                                
		.reconfig_write1         (1'b0),                                 // (terminated),                                
		.reconfig_read1          (1'b0),                                 // (terminated),                                
		.reconfig_address1       (10'b0000000000),                       // (terminated),                                
		.reconfig_writedata1     (32'b00000000000000000000000000000000), // (terminated),                                
		.reconfig_readdata1      (),                                     // (terminated),                                
		.reconfig_waitrequest1   (),                                     // (terminated),                                
		.mcgb_cal_busy           ()                                      // (terminated),                                
	);

endmodule
