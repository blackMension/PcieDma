`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fUDkQaRjLTT+y+ObcXEdDkE56RbFkeATDTyXeNMRnJxt7DSdvvjeles0cHYoK/n6
h6rFe91XvxFXV9l9YWEKTKqgV0/m/M67+Pp8jcELumxKSG5DJUlLsNkx0ERAKSQO
/7WcVpI5FJ8y4vzDPuxXMWgrHT2e0RciXq7dOd5jH0A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31728)
PCMRBzf5eb7kIZneonKPfdv7ODgryxBFaV+mp2y7BN97/x6sTyKoS01w270CiYB4
9+QRScCRFvx98yX1z0bAmVdICEqmSXm6PSyqhWEfflE01Kw8a13yd4oWynLmpd/c
R/XWizROazq6HER2AvJ8lZgRMUMgONli6IUcHtnoLLuf6Wx9VU7u0D3eHRBtYFdd
1lBjROO/JRvrfcOR4XN7kP0zMLZAI53JG+0tQaj/0uw5WX/JqzlSeuaLwZc2doLU
PHEJkjKS+WUqbs1KtwS4bmRJDq/j7HrbjgY23/UIvSQ/tk4BURfu3Owt4oOqb4Kd
k2J03APpJHhZRuR+/lA7+fxJoiDWs3BRtBtCPZVL6npUCIzz/y1X49hm3LmLKndM
ulXyirgSh0mEyzjVLb6Iy8NnvN40/RvH4TD5PRkgYPQygP8+AM0lwzyuCswYd3kR
TuvH8B7O2LTrFCNeRjq0+er3BI/WrR6xZQW61EPJLgO+JPyhdqJ4HPc8X04gJlRJ
6M1Fk6c6Kw7Jaq8PZIj+o7g/Zjz250Ap41Z6mXatmMUetfWJi3dwlfCKpJYaCvPI
WuGDjPWklUraI6ABGBQsiOsFBU+4T72Xacr8LI+Q9n5zrfW72HKRwwmfPFwYF49G
L2Rv6ZiPhi0uXmjzwDKwGXb9GdwGW53LpDGnEGMuuxwX7iEAkK4hhKGVpi5QoOXj
PHzgy/FfpuMGlr/alORHyLpLutot4Pa6aosAAgOG5W6IRrU5idDenecoi5FvKBu2
Sa/8afOtrhcXWJRsbAg0WhwrDIv0tnuFe7WzIABtjj+0k7WqymCuj8Qd+G2noOvM
QEWb71/9vKBxWeUGUwyRRAd78ZOaspI2E3+8Vz00YDODrg/CtqHjuZTsN6UeviXk
fMH0wemhUR9NUM+ODojudtCUiZXY8Ll9xQkClSYAb2r4O9IJ1boD89pkda97TdZ5
ZkvbeLLkW5E6xCig3vVmvu7U4jNXbG9lv0rPI5sOossTV71GoDQaQbjIWWiRUZTF
1Ut0Wg+1+0SzRkMheHHOSbW6igZXlNG2jBZpdMtoEMlirarKonJIgd9fXcDDwbwL
a6l2LeaKf7haF+eqd0TeDmA8bpk2Je5G0xONGFi0UFp0xxggECbjLUn5u2nyBB/N
y6VjSfPKroOMFTT4sNABTc48Hoz+ytNJ+CEL32GDo3z7Xj3XKcF8fk7+9wIV+GM6
B9PCcfA0LPj/M4XoBcKuWpf5gKGS/nCFUA+rpfFKUI0I0cAokaQtUdxXNMvDRmFj
Oy6sBOHq0beS5G7Kzz4lfAJ8HBuUxHM35ouUGiOf+t5BVbjFIz84fYkepJ9mgmM5
hQMuPVB0oMLx1b/g3mYxSTucSXU61ejBRcrQTi2idlD55p5A0wOCRH0qgFIfLgNb
XqOBSbJ/2mZrzJ9SNixsbuSWEyfcMJqQrqEUK+YlNU8MhwOuOZNq1GdDszuywLip
Rk9TlEHIf0L2Iroh1mCwTcK4uqrLZo4v7VRWgs101vh623LZokJ775aQqXa6CfSX
T3/bqni0FqN2MjSkrq7tty9lB2Geu4m+Yphtg1Uu17Ky9NdKdF5WfHOWYy1SnFdR
kq9ebvHl31JAoz5HzNWlXC9BsrtYFCWmVDZVUxPFjIvwsniP0X5wi1o/lzPPUUkI
pielS5KQiWXnnEUCoBeqatlwWpF2d2LIZzuGLKeZMe6wBqzFyvkBvYUCRqrWE/Od
plrZCy9WdkepNQxQVZYOqbRSNsXnDwTeHSxxw4jW8JcGO0HRQiLZqLAkPuDwuJIm
9uDBpqjcwrkm5ssZ7hFY/obITMK995mQ79e4KayLAO3u7oiW18JGleLOc+GrKbL9
HZRBvR8pC1ivRzEjmW/qO7B+M/JcfopxwtNaDCVQGvbx4nLLd8Bw03YnXt8EnUiJ
91FnL/QA6NCdeLceQD3ZM33vRPV9mEdbhpP4xwQvpqoWI/OYd/NhJ85ga+x7DgTv
Oi28/LChGZwvOsL8qFyxP0SbN7tRwH5r2W+SR6gpUroxyE5EyUgYn/DnxwTtumLp
1SdCRJ4pdI5nC0MnrvyRAgATehx8yiyfUJK8QEHYEDe4+AADeGwtJUKiPpMkhpd9
ljlUrQEPL1Dz4BMhnCIdh03OaReq0Q0RRCZoXjRDBS4r6HmJUOwyNrzNAMv+yGmF
iSGBZQ/sSudzvBHM9oN1/Y52cTzzGoOzqPYGBg5r4NyF4FpBWzK3pfNMHj+vqYfT
CuEVMbai18jSoztrgpEmteFpUymhGsLTaY6Fp396EUSOiOTeD1nDz8nboAlAz0gX
SAJUcEZpmbZ/NXrsyM74Q8uz2+cdeu4fFKGXn2+yoZo6vbKmtYGJwN+DlqECaYKp
QP7vT9r6BCJMivI0z915bmcP38CRiNC1qjfymws23TsaUMTvK7OMurLxa6QmGCtG
jrz39XIE01gZopRgQpyE405usCukEWbgl51ZmUjmQ3juVcxdSMOVlE+dWEAw2oeI
Asq18YGxUqKPQdf0gqzW94oaN3gySJeJhL5JoZVIP1MYvalpLvbV0i1hSu2JGjl4
DhAfIAM4A7M68fwZ1uIlDu6otB4vN4y0dGQtafzRsklrBYsmdInHMI054gY5zqwQ
6pIiMYBBA5/oZpCxUdZGLCdTAO4ARgEC3poVBCsKGBVX8Z32WJruREF+zdZc9M0Z
Tr+QPksLxIwL68caIjIC2Tf40fXPs14NUTma0S/OoSRG4ZTKNpjXxfRif/sf1zOz
amxPBJJ3aX8ruroWSrzPmTOEjG56pQlnjx1yxF8MOXoq8Vf09a/KRWZH0ls78uwY
CkZ1/WlBozjOPWkttRDiVEqZGkhVdxWtkPzGFdJfEmXNywlbN/Zw+HDUCSsOa8HH
7LtRb9c7eVlNcUQpblUIU32eqR/sAISbcSrkdQpYmzZk6dnIJqiDxUNmwmbVrXVz
k7b0mWN9Qvxj9/yJ+C4w0lmxonsdxcEZTfm77Np0FMgJf8vwFuMnLeJpdE/7XXHQ
Q+d2jbjct+Npncg86G5JzGbsKX+WIY8uc5Lc33bHaqp+7khyIq0IiHmdEmFzylEP
WydYYyvCxZ4qfVe4ei4V4M8BRAuqVmL/7jU7BE6dR4TqnChxb2p8pYKO9a0BeX09
lTTGC9LSgGjPuvu3iAIcim79CGy6jvGTIyBBJPMtSBKb7WigvN2/q3wgxdf6b8Wc
IUJWsEd1lds4HoEGMqPVQOfC4HiySpfJVMXewvfQHmiEKRDJdHKuYj457UM+iS7c
b+ljkIXiOT4Qv1qHtwVX14QkuKYzg17qIBrJrsCCOaaXmxfoOU8tzZKT1HEV/6mA
FVnobtOPleQoIMhk5IDPHYGmS9Bsw7JPdHBiwzdQFF+Zi0gJGR69Z9wy/4JWYp7M
oN4Qy0/Jr6wb00ZWLwJ8dAgYAw1pHVsXYl6caTK6tRiC9JM17cfbjNs+v1LUVEsb
6+4GP+4XXfl+txYBqhdopLKqNQIyili/98aiySMVCICmp+RXL3nyRjLgjOcVDrvl
yjHhXKoVzZRsdeSQ0EirRtVZOdsu4jiG0I5EpHrf/aZz3cLHtnHIbEkNw6SM7lqK
YVwZiA58dXiiFuKhVX86vjKjRjybq5ABHFwNIgcjUroGMxhy6UMZD3DI3duWJq46
2oCbMtBhuM3JIT9SyU7CO0Z6mZeYFIEffgtFJQ970vq/8Lg2sr69hyoJR97TNTpO
1BPxVUeCcKJH6YcsnCA4SYkOFFr7rXON+cJWKWYWr10l3jABzBPSflK4v02Nqlpd
n4203wrh5Z/s2YFkvcCnK13KrfYLF34UXdpgjCs/TG9Dui5DuO9afk+yTAlakZ7F
obKz2rC8KSweZUCfh1WiDS3+1GBbD8sKcFDMdkG1ci5csBr75V0R12aP0Sgu20Fd
UcayNnfSVf0O2KKHDfIEO7Zr0bTO8j4PpApQ6uR7VnpIpCev4xgNiWfM2ayZ1WfW
fEMUAwTxhXK80jgWUBgg4NzCSS2iiLgrPS9H1CbXUat9/hFqem5XyoQLWqkta5KF
BfGPZexOnCAizMOQEPuqvdjigJALYfW7q7eYR6r1gHn6hJCB6S6P0QiF7iWT9ZLI
NlFtFvzrB5QTwkvna22uqe5Tzc2DWu5CkCSXSzC9Nz13ebhDuNWxkRSkFXjo3sh2
EbGQHqisSj64c33woYKt9f8h+SoXtC8FIoQJyXkFjAAWMd4vHly8iGFfB7LnQnJ6
scTheBZa/ceGb/7w5192pHhE4IwOaHCzeeLiLG/FZtUGPtJteOoL7qirCkuHLP3e
YH5yGg/i3geT89517Zm5uZ9UbbYiYpscMzyhfuHcezAXW1yPuJf0YaVGis+kOZt6
dYzoNQi+FFMAEy6PHBX689xH7/hHJAqS/4hQveAbgZPpD3b5roi5nFNo90BaXQmj
EC1bWLFBIuPlMi8KFkmBf9//uIfAGnGSMnQqmSZrZ74L3UsNyBFVVdbm9iMgWZAQ
kCgmucE1e/2xmaI3Dtkl9FcFGQDH6FQeJ8VoXRuONGHDwUmHwFJnuBj+0bhAee1J
/xqhQXzABuZ/Fn4NPUirhWiM0KRWf1/XrXmJ8ANSsFk0QpBNM54VNPkX9oEHmKyP
0eXPu/Q11EeXUzIVnbWdaeH9vBSUsxBNDgi8aIqwzpvaFjabXhJzyWGBiqvUBOS8
CnqomosrRQdYf/Z1/qOpcGqnaLW6BaBTWwWPE7sIBapVveu4NiCMwBex8rLORy3S
WFjjoFn7GEpa+oPvIPe7bHnxcAvsx/I4poYBjbWRY7fghe/joL2gK6vcUnhzUx3S
FpBKKEONRwVJcxyfbC2XsTyiqrmyAc2if4K9a1SjdlhV1hKKb8IMbLrMdtobLviq
ztAhK9TjjjHYqdPH1hzY8FjF1HAq9NN9nmDNz0MyZHcAJp4dRvmKNMpeh9hfxe2x
bsluRwMTHZ9g13kIKvRV6OiKWu2fMyYAZcnWEg3M/lQ2KwSDea5ernaMAXlPlDgd
awwt0L5iizL3kwcx0FbuAwJGz77LyoyKJtTe+FRBK5GQYlg6yzt33H4vTsZExWAS
Yqk/tFDp334g4wYzOimhE6DfdTbF1Ks3fMUwgn244i0VbZNR1XL6frCN71EQ/bOb
/iT9qG0r6tVg0PkKI03OCpv0EhL5FjziAkdSFBVgyjcTsBXkhgtfOGr50FWe6RYE
wYklAcEjlrB/VLGiUxgmwwCEj/8Y5pBQO+wlB+F3Qxsx+t7CkFKuy/BFbz5PQ+TL
gU5rZ4LzhAQx49asTdUbSuYtvO4UCKfLvz2IWJCbh0bTkcwJ+oeg9Qp8y0BLHI4k
ygHYo6RZOyRNGsCD2VCmuDiQTexxTy9d+OJq//bpR9C5sdR5FGWh7r7G73IaFTj5
zaEQsynjIex3DqSFPKkjftOMC+SCTUUPRA7ylQXYQWYrTlZ+yLZeW3rB4VAE4/Y+
GaAvpYIR4B1jBQZPV+FVyU/HTzoPa4g78DdJ91sVmXZLC7c6PdzScLTYyROFWyec
AC1zs3v6IpYblhgGwdG1M44GUv1BTkms0lGhet/PTv6YPRszeS+7fkMB7xEh/TpI
6xit87pWCXmDLsjbKngXcAv5jqMjPw2NtyCEcOH7rfCpW08nLFYIqX5wOQOWutgS
VOPkT+yDTEBOFW02wNrXhFi6IU/hEkyjRXg7misfN7pIlZl8yWs0rRHrl90vx1Zy
5F4+e4L2VjLJpbgPT/CtP65nYpPUlSm7wKwt0BwhK3qJcu50JJ6DSlTj8mVcGCEl
no9rmCHhbEukCr5GFUNDKCzUo7wG1SGtzVhoJXsdz3JLjkuIrvAZNX0PAOwgbnyG
1461o6PxHUsmVbPoUXMwW8PwEZ6+gWNsrCyM8GAr3r71R+w+hJZ9zSdDXrDVqNVr
QnFb37LZ0dYJ+vJPjhL9yIhDb3jd5LzCMxVA13BmxL0mBIu5HvSlSYusiZ09qbQm
5h+YPJoxfaqPnRnIcxo9heXfHjOlVr9BBqh4qNfvpDzlS6nbxv61V7xMc6WkaA03
K4GJa24QZb2ePbkpAlsV8bsvUvnb8LtRWamJfW3sSC+pR3dzNDbuzv+ELvyRO8U8
fAFkBFTyCEsUxQIBYd8tjX7poIX4MZmVg0LIgADIpiCwpgKT1kWz6fHhpJLyykb1
WXo23cBLQAUNe5MmTl3NHzmMbEJccPSJ43Y6O5E5osxOTOIrfh87pR56Hb3Z0EOV
oV3joAzjGEw1SXbMFDzmYEDjJQC0Xo2ZfRSe03p6Rw2VFTXb8y1OxTDhYPz13LdZ
I++G/ixYTLDpSSDKQo9qlKahmwYjO19EucDqcdTH9WHFKVmymwkSzHCYSua8AnHA
1m7Hh8QIP735c+vLuzOqwoWAPq4x54q63ARPUnbha0evmVU1We86ZsNhe6yr0Xnn
yN7s3gko6FjQflHJhmOx1kG8HfZbyUYpQCVxT4VdDSuFmSAMy4AsITPQcfCOLOj2
7UszfpHfri09Nsxw8ZeU4d2sHURBQm3i0LFD3pH4VU69hjTrDbhnMy/Z/kn2f9B+
Pe1Gd2V4r+5J7hwVksldJTN+/ro9hjmGSQnE7B6NzpJF/wVqGqERQjFA6VaB0VkK
5lOJUNZwf6t3jLzNiani7KZvFalY100oHfOrZ1aqPTrbWWH3dFKb9sLimMtSyzel
pUlmBF60YUvjqX5sh0lz1Bt7FRSUVVIH0YJOuAXQsixbloyM71SS2nnkg5wHeXQw
osI4jrQeL+xTny9tgzbtT9xFp9+3kD1kY56MJ2oy1Eqz3j+9gxH5VuRJfJlDueNd
yXetSpaqv5PxkIOfpcTl5+lB1W6UNP27dfFcFJRM8hgwnSVWVgpOLqrKkYNAels/
hf5RKy32qvGpvCm+dZkiKAXII2YIi4hcWi28VFJgopSOmdMqkFVoO2E4UH0/SLjJ
qOVVrtiUVkN9z0At2RkLNWWc3LyE/1LrQWMVdT2W1C3Z627XLibjMCH4LWGxnrUS
WQKso9b6TTyQacs6hual7+EzYduGSNzPGRa2PExSQ3BKMfHTUufNwo+T4EE2hj1f
NL/NVR1iEO4DPwgRoedIR67T7CEZ2tB+/ErKEPFwjO+MsI7HZg/KsjCDhfL27kYB
0pKGw7nHjiXgwlbdnVHJ2Gh+lQD6kjw8P+w1WkMYT38jUVpo0GqotewDLubLN57T
PX8lKiUpP9DjeOxg7y7iG4FNRtd1fiEzgBzNZx3k/kRNhCOvcoWtejjT0eOGM4MN
o+fwY0WDoqL3ULamknq8YWJt3F12YRAQHPUVJvCmSo2vOJPOv9AyZNPTfw2bEFUA
Lbp0O3VBJ5pZ3Dx5yfwH4p0FeNxjF0qP1hjbH7fAK0yLNPMEgy9av33bebxOQE82
c9rBD3H4MdWBtKdxQaUB/HPToTLP91bYh90oViq5u8WzrvpyX6t0pW5FbRaAOU6/
vIGoqvEOKb2rMDGXsFFXAzbHPNZlR5QIcKzf6o+KAESKDITNVd4912PCUPq99Oqt
fo1xIJNPuMEhgH+cTJyLlFDviO8k4x4nu1hiATgUk47rhCGYe7WF99bKd6f4w86/
wO5IXQC3ELag4qf1+DOwTAD5TvGOJ3AwC86XGZm4AQ7+m4VizpmWyHB8w9d8jeub
Lrb0+8GZ3uDQShf2Cr6onXqkzh/ri5xukSwsU+bUo/BxVOkxFnL3TYy0EN8Ze4yJ
E7WqH01+UrFXitSi6G0rNUcGXb9cKArlngv8++asV0QnsufTeuo0fi0kriCzwdl9
8BYFemvXU3/5OJuVzQnye8fv6zpRsw8+jTuItihMbYu/Fg+Fgfu/BPVMxL/inyjl
yjBJ1PCMwLUbtgPSU2XTU98mrX5TDVj1DVUO1AO7CXCaJj5f2MQXm8XR/DNh+h8Z
GRJKK+kMrV7GM0Mt+WEEsVodmEzDljFFte7/OQs+AaZlbm8LqAO3PTtWsZdWtnY2
hp9SBZ81dbVeDPrIxT54+faWQWZ5JyM7Fbbc9yRe9B5QoneSFgNiT4qX3tYu1ZLP
SoEyVfHq8AYphIwetrDnzfZGBX+58eiS6u0KWvFCfFPBkYkhwnbF+wDptSH3/Ku2
mE+efM/+QDwoMaZOVLgnKtZ5+v73/Hfjppz6Ucvs2NXkxVOwrSdWYvSkgL3DLB0z
/y4pC/3VCCRbNAFhO9xJ167O9f7RCRi2GcMFCVyMFpxLVuOkCdC0saf6iImoQM4O
p8M3lqzbAcfhV2KE+S+3k5UQdpCb0iP2J2ZVVcFqVvecApBWlXhhV+Lc4cZ8uL/+
aZp5Wgy+zPlLJ10Bk7RQPanKTr5fdO7YpxmMIUVxsUXyjBD+aVY5YRFbFy9dP/ij
fTfoJaJY0gMcLFBX24w9mrkaF12LuwgJyE5rZ9h5UacE/a43eJASvqlgpVxgGlLa
aRkE0Vr/z23Z28vzSNgYlUCGCQhtcEAzqpu8yDLuE+svRrsFQzRhogddr8kvxK32
bvkHjD1yBJ+jFS5WF9vYI2azJ6nwyjIiwnteOn5n/CTyD4ggegiXbfFG8iH7Gy0Y
AhMLNAF77egCsvrLbj850T3YY4Kzn9cQZ7oaWHjAZMGsKz6Rq+RN1ygAFNJAVfZ8
/k3stXgNZMVT+L2Ie2ajzn2z+o4mJEhiTiqyB/itXdCCQ7v9ZfOdXaA9+hAJhVIY
VrwOxse3F2m4j78m3L3roGB5CIKdMISf05d58H9wr4mZE57zsNd/mK2/DGnRPCaN
6/6i4rP6UVBIZj0GK7gCkOnSgCNr8/3xuVeGKOXUpv5RxKi19BUFHVJfNL9k95qK
llTOHhBrIr/JBZdgYblY2rFloUatsH9cUv9m/lpar1+LFR88rjjzJjT7KX4QJBKD
qtgMGRQdcVIzBhsDcO/WMXiZU/DA/NmI3halhTcMGFfMaOoOZoIzYu9XcS7p/9fz
llF8SIid1B/++ilXKSMoRhHCo3qlyZ2XrHhNqqMAO7e0JZp4nFuzx+0CXX0eZDf6
VRsrdR3EXArI3i1EVu1wFdPUQic4gQM5UkGRtlP5xfAp9RR2WOYZqYrvu9rMGZa0
gqAbbAl81zFgeQyqqrg9CbySrFqARn+DgZw+JV4xQrQq1vLX1Af4bEA75SvwyaYV
ZqNqjDhh4kkU2FGRkIY2fLASXiY3g7VT+7LMkQrBpNvCJhjCWB9nJ930H3yyoZmm
gyBK1pOI5TG+6FojW6mYBh15X5/0Opa3M2vaNkU+RmwiVtoNmXxJDPJsuOEbVl6o
6t91EcE9lSGHT/zYa0wKKl6L4NBw6+tcudyEvqQYhIv2KQs8N5E7kp95jPN/ZZml
4/O4O0iE5J0QqQtrxQYBQU9FQs1p/D5VfohLM6ysE8BhyC626/c+CHzv1z7DM6cO
vXqoictW25vcvZrpbNwg9ofyxZtR4rzjiYKnC5441dLuB4xL8I8CXQGOYZkXP1mQ
uvw/136ts8rT1bDsDB6Wkl97CODj21B7RmP5bWayTtNWaFc++MS6evywgWVmu9lo
/2eqN0Z55UqUjaJAlJNkaNY9HZeTO7aoxeklpXJo+rinXokghLxQHzTu7rzV5nmb
QXr2Dn1qbeqpYUaEnnn5FfdxJdLNpMOpdQNW7FGRpDugTscNtadx1a56XOpKpsIN
AzFgQlnnfOcb2C+o33FJaJ/6OVaJet/qxVdVrluBwFEfiRzby3P1+O5mQY+XU0Cp
WMTLkz6WNkWVv/qzk8za2+EbWjIE/XHI+prFXYwNhd54WtUmnM8gphTlIuglFt1M
bfe9ZJ9jQpG+CoB/Dp/lzQ+tnneWE7YyqApasYLFb9l8eVVISKKkqF1/lEVLKi/y
ryiPOUIghiM0K1mSrGW/pX18sxPnRGWYFD9Urfl9l6ppQYgMDXiCZ035ZBTsIPn1
2MmHylVERzjLmEWSDtDV4QOKVo5fB+i+fRZnYFmZ7Ddh/tSC23wgwEJS0LC0AlEs
+pCFREmhizvXWtvmE2jW1GAZTIWoekOiWx7c7mmB5weFekzEDHBHoebdXJI/a9Lu
ULNcV/EriQURSRSN52J/e8vhlJJHRqtMcePBuObyA8TIJtBNvJViXXRKO5OoNAk0
gPP+VY8naQvm4kGb3ZcZSs8rnZ6xMUUJ/pCbkfKW47TiC1XLU4+VfJnA2O1VExVF
Na7VMI+KWzkG5zxjQXgGMw8GYuQCD3G745n/Jy+KmasE5jKeDMwAkrFx5vpdvwP7
Qo9vO7fP6kwetAjRRfAV4Fo8JUOnkKB0YMgICxp/SqO8KNk5XK52rLT0NUEtKkQV
gkYwfjRnpbye4+UQFw/yAx91Ps/thN6NpMnx49V0BSRRoENWv50tnQiEzFidI6R3
x4CewdabqL8t5w1GLQiBDmVQmMJwjeX9RJltOQK4zF62RNwDFv1inV/GgFmqRE+Q
3NcZyj95vRjRZURAOFNeWOiLj3syqllb2DPQ+zo97VJqNIe1FwER+4x9HniB/PlG
KzJ0+HOnKkw/YFB/m4ts5Va+d3VoeWxoSk3hMJcn91cVx02+y1ItVctM5fidmZya
Sel9x1HzIBMZfJer9y/eitI19OlrJ/4Kam8/YWxgRClyNGcAfcCYcffmJYVbZA5D
aLbUBsS4llgOTSglasBpg8ffPrfoz+ypXBjUyMyVHZIqWEKWz1kCfTgz8EVbxipA
PpdIkJni+H4GhTC4vCle0y2LgZOLZRq0PKwg1q9XlL0wKHgR8hZTRb+9XOECsd1N
H88523dDOhbbHPvDEclDvrQy2T5dV+QWFKzCLQNSqs+sJ2ds/xXW2ow8+9+2neZ9
YWoXMHHeLyQdoJ7GIbcjON4yrJ/+iV8CjHrkHnVTmHxU8slHOkO2S0vd6cUlVq3T
ig70qdml+rAdh/eZLDIBU5U0UWIL9ImMdClhcAXeSEsENGkP/0tDZx4bVQnMjweF
Xc5yksZVW5q2Db3vy+6wKYPnXyv/YVGq/ewHpWBchUvDY7LZFlQivx92lzef0lwA
4v8zjIntQ2uHLBrmnB5mQCo4W0DAsI0nlfE2bzQcuQPH2TwbYROScrmPtsEq+rO6
yB4OHhAwNhZY3sK9cWSZ1wP3PBod1n1/KAqNF8dAmw4zyNu1ETUdAfyYA4VRnqNU
ryuuEwH/DiBzDjC8FJPD0b1/uiVbyhiBLpo+VDyoIWaOjvmiWli3i/VwB98PaOu6
aib6CwvylxnPh2mBx8gGySSReR5gMS7nIPixd2c0ksOO+zpxFjqmLg7qotN8Jt14
AYTMPuFi6x5UW1wxUSdx30yveS9Wv+wvu6uBZU/yk86NjHKaqy187uJ+E9Kw5Wr7
Lo8EEliRonBfIM1GLbP2Q4Wi6FMxwV2nIFzWkP2RB95Dy4+eiYf68hgVdK6iUkUd
pC5pSFoxNlm6fMFDcZstDPG1Yf/nRmtZRg8LWZLR0js/okcTMPEJV+btYvxbVGbt
fT3g8QmTpUoQJxUJK8Z/2EoE0HLyTwUejUfZ3nO5NdXYMyIwBRt1LPL8ybLMFk+l
NytX2QGnjR3gxTrUZB2rfLzT5QkzSQbIUgbvAGVi5bqpKcGKlRLZgcwblD5+AefW
20QAkmhhX+zzZGC4/RsSKy8DfSkhJEtWnAwBeKsfCkJDiTkDCj5t6SVBn/ubfSLJ
zU1HcUrJq2iylKdszK5eZso0Z+TNjJmE0AUPf8uQDpDhYl10dEtkPIMVV4DaGpr2
pELDIDfsgkj+04PhM1gAsznZMlUhqVsvoU/cK5xuuVIISjjOLg6lMX2m+bFcBhml
3HPQ/9fnWIJ/gLBPHMQ1hEXt6BLXgtJMaAXwkMOpyLFtDJFf0wVBMX1wh7nfdak4
lJSpj858EQfzqekTeX/45sutsCbFQiakYeQ4WyoGhrjc3NjG2a4eG9+CQxi5Kmnt
ct1o0reei6NccA8ZkdMHaLNvmjcqZR/Q6sNZe1wAmEdlCBsAyvJtLF8T5teeU5Bw
E9j+SNo5lLj/sK8zmcOgPAdFIWF4h4WLGG3BMQ/0g7p675Z8FkttxDF4GLPBBmmf
agVmCXNWs61EG0MJ3Q6X++XJwSG98boPNCjxAmbdGfg06dClRHhvUkoWQJk1wyi6
sOyclBF/ywMr0dAR+6IuFy306vLICqC0RqK2yka3wIkdp9Se1+JGIYW7qPLGIF/I
ErabnpxPHuL893O6M/+F89Gyo6W8Az1JqwO/18QvMP6P1CGOI2PEd8/2GF9o0loB
jvLneBkCHpz4+4AFjKG2/WasTp27wX6qRMrx/OC67ZV2U3ApFughY6oXd5Td4h30
AbkSJ0kgItzkRAq+2Zy1C73E57WLZThlGYNamlOQ7p42Kd7ZbCIadCfojCcRjJWt
+6R1N30fxOo6EbwAidYSGz2HG8aCJBqTDVvKGYOks9/1m/TIW9ue8sByCvWTJHMg
nhyWFQvv3TS0f5ELsEONrTXP/mxDz9wqVU71PnW+1dmIQ/dYKCgW3SQm542E9H0Z
TGqVR3OuQVewRbNXg5Gn+zf1l8zw/S1I9LNpEH6cDgkNHQ/xxg1YESe3BduyOMa8
0Ydli5InY2LxGOV6aXg7c1kur1pNhNKeIrXA4Ct1+m7Wkpu6Z7DfC1a0OzpY+dTe
e9/75qU/GOK3q8NdNMN+kvGdQ16fRd3vBBggBrU+gFvdfmGXs5+DEYvDbmoooDnT
prhC6ENXh5QG9rhTwMu4pb/bwCRu4Zy07E868fD7mgLE4z+pqIwAAlVNSb2RWOl1
5cWFajQWXm2SkzIPZqKz5GyjeEdLZq9rTUADT5VDRvabPgBtyrQJLT2nt7UmJVBC
QBIVZiL0XyCaxunu84x854LQDU4K5D7kR6n0QohtOOTSl+CvdwpXmpoocSQ+4Qk7
BvQYMcPgc8utKn6LNCBEO2sZp61tYcSTJxXQO/YBwmgLafPVytysHyQDp/wdYWGj
FwSoodjgtgMwBz2jtCT9z8iFJe0nV/DSnsLEFUctXGSc6Rl8e/Ojj3HCtnBT0/y5
OmBIycDyhn/cRy5uujXM9Ih1AlY2qYyNbuXzGAPGqhU49ze0IRqrevfAhlKtUNce
bBnAOv84qJ0TGr6gytmRlwt1vIJFcWBzjEDkaqliE4gfW9m5fb482SlsZTaiZ+w7
8VkdFHSQ+H/u8Y2WYrF1r2Wvb3Tj40WfoFeVC4dgfqscKbNpSTEzUC0xjnSdBRXM
lN7SOSIlSCEyOyULzgiEDW0rZ7iY4ijN+/HmzUe8XDkVFs1SsgndZUmI1i/Ixbpq
J6vdYcne5c56+eYM567jOorKHzOlq2UmLI0qO/KrFnogF6BhNqPBiNQz+erFvXLO
wkvs+kocsnWt+uCgOofPSMTFizN48cA5qzbsiY5a6eyzZm3C3a26StFNJde5i8bL
TTLgy47C8o9fRZdhtZt/OTm2Xpur6+j5fVfQOdFj5zSEZ0QSWrunUEOfmQ2ftiHR
JTUNIGw55s9SU8PKObEYIayMq9CkZGbVoz/1PDtzCsSOeFaP3hzFnSUvZsiy4h2U
/CEhkjQmQ4jc//SHQdEX7KmHecA3AQWyaB5lLJgAPkfmAPRmCJHR6shLdQ7R49Ch
kRhoomllVvU5T8KFyqWIqHMDMMwCs3nqGuarui3AzuWelCTHXzcih7LsxjvlBxSd
7xL1FUsLKPkyUCB3B2/IrxpDpAvTnPjm7VBKyG1+rrRfBIMUz3ycPI/bp7/XKSPD
6UHFIViewDNQZmQEOb0zKgq+Ss0Y2S/sYZBC2VKmYXIEUouAxYMLry96nz/aAEcR
rrCIqubTaL/oYdYDxuMYC/HqwtRnylgsvOx1LYKK63olXhlii0UpZcoPMkl2joUF
j+IbLMeCD5VRW3bWficgDF3psd4K8QfqLnfuSzNjgBbEvSbBZj/VQjNfI80VJXqy
9I3RMo2gAbkIgesiAW8LfpNI0FHwfRNSFsUF0uaj8oQp8+HACuVXKviQOrm1hWI4
0RTa8JHuV3yKdmkBaxgYFBV4gqRbAGLO0MkCnKvBkWT4oeJ7XXwS0ZG/2r1NWdhQ
1wgI+L5oxOT579jLRjmqzFtRyJgH5pi6zWOSX/mDKv5Fw53u4i5dCTDr4mR1Of21
M8OOMaQ2lzceOtmpYKkK11ObiE+dw7cWC5cyXyrQivmY6ATWDU9sNvJgXs4KpVZC
wvT7AM5qO3BgmQsbcs3HGZHwwCktSXxzzEZLdiiufObTfWceTpXpXmn1xHiOxADl
Ah1EgmFkyruFaYTAst2o012GLhqipq2Sol98pVToUfhmo88KsOhKRPUFjhZMZFD7
qk9VIbnabCd/ERgDoHATXmFtGPIIYVCLoY+xmCl5kuXBYLSAf5SaTx6IfuzF7L3k
sgGojMNB8/tm/N3zne7aMUt1YzGrp90zHJ9GfXqeA3CfKp9N4spKeO+OUPS+IGdW
T1Qh8GrqphjjMTOO9sacD2sbeU+rTOEbT3DxqLkMOOOD9b/mGgsu/TsrOgC6ZhM/
oJpOt9AAMnBZzyDiG5UhVCZGdyVH54NT3WRr9aZi6jJEZf2dafkaHDCaeutr2TUr
x1WBenKv4aUNNAXTJSMulgUpubtrQMd6SyxcC9AUGkMKTcnZxnrDAu/f3EtSOkac
HQ2zY6X9DuF1ms5+yagg2cWKGkJZcwDwK0P9rSIFQgIa26yo5ioQfaIoWPvOTZDm
88QthXyud1rN6jc3ccF35ANSBMN22QtWa7134R8IQ+ydzBXX7CETbFqxWama4jJV
lCu4YutUAYzPaRhq9d+bGSR/GDkyk6v6OWmE4bLrnJCS+tdnv5nwr6BPlVrUvfbD
PzK+2zANR10i6TMyToWPb0zDQMsp94M+S9XXcbKKuB0raDaw8qu9jxy2r3YQo87y
+5AwMa16H5O2T8p9qAYvt0sQNrOMnBMMXB4PExaZeodkDBdVkzE1GXktGyYAX4Ps
B763lSglHCo6C4NVkl7FhSaxY8vlJUFJlhfbTW9o0VNsgZRa/hHMYLjIJuERy4D3
kAFA/wxZyL4jeH+IOYUlynOJnkrqDoRREs6SWP8pJQVLNEE3eqKT6p7K0XOx4GLR
fXwlKiPQq8COsTJ4F0SR8YgF+aFfxkL3jqoXbSSFMvDTVG4AKFQgNuaflbtwJs8d
lJMl+kwQs8z9fIfRYgcSGnO66En8lDXBXRQj7q9VrAjUkk0P9CrJOZKXVTZ3V4o9
6UmYvGjtMToqny1SOXUPz/IuMcH72LF9JIahTWSfVNR1MK9u+8TlBemobEoImLte
o+L3qMs3x6UcBOYV2/KZTzjEm59IK0GGfM5wIYmumvv6TfpDD24BwQVqgU2zGDvo
KdAaE2ED5VVGLNlJD6lxECnpMBi3WNyRJOpAuwtuYZsji4Dbtv7BbBNX1bsC2366
IZ891zN2m2YEf4Y3sGkxcZKz7BhiMblDUVBvwM+Z+ZzJkhO/55Nk1N/JA2Sj/MXQ
jcUhMLqSldGpASkRXvtCXY1KAIsgELxY4F3pnhkOkVjGRj+DdZixYbTaeq6eQo4p
RwslYB9ML5Oc5ZRphwf6zQgxjLKXGh02RfTlFYfy5JjOMhSokAWl/JcxJm+629Nm
MsuZ6mc1vA/8YW+R6xveQK9FENKb1wJYN8FzCuIzoF1wAFMWZKA6YuvXSZsyfDpj
qNt0GRbt56C3OY73+zDtp0qTe0CdgXRcaylpSF2OZH3UrF8QiVdsbIxMjme9A6gT
UqhHjxL+fhuh6f8JPvU72EAMC2HNNNeK6bo6lXpSIdj6/VeHyATTnauPPhwighXd
815oTnT+2neUPIxq9OjZ99XgoXjzsJHFe81/77aBiufRgE9Drwa3P88OQqA/3btl
v3bps4ylksDXx64L8GVDpPX8GRfAOECCKvmdw6IBWUyoHtC5khsxicU3vAs2yyr2
L5ymDocZF8YvawYtDUWNJGlfuRUmmhQL19iyZUQdueCnEGVqtDoxaHKR7xVm/Sz+
E2Me9S36W3tN672V0280uOtCB3zF69mnrxFdSfikIDRY8OfUpQChI5DnmQMKqVfn
VCoGciSr/09RH1FPBE8th9a6jUFQZ0dSBmIATIdBVI1DxxXevTRo9tNaOWYmQq9N
znq30jzdjlkXPGTtiXhQT3iJhuS7H5mPRf316AWpcPH9RJDUpeXRTncsaP+c8xuE
QTsAEKzd3iI9dITa2azC+ahFTroGNRV7SsqvnkGG17+M3aS8REAMr+EHsvJIp4Xr
lbot86R3UjV6xzUwDdtYGRbCK5sVhpuNTFMZo9N45RbOdsR1y3VPyW6F/CB0NZ44
DXyZpR0k3jXsjK9lY0jtxMhr2dgbgQabC2e8T/Eiwpkikl4mTmPU15IHMfh8RUpr
sc+XgGrLEYB1idQQVzVahkJS7z5RSk2PNBsMCNcmVrBVVtugPApYYarW6qU9p6i9
8CtcQrIlROrlSbmsSBpoGAG8d3NC7GrUSwJyGRz5YtrLSGEZfgUrp5752HwgNa7l
8jkZhhe4VyIEbQIuhp8KcIF0I4pV/siktrEqqrjyp12c84ZikMmiQveCPnHM3S0g
XwURzkX2XJX69hlFmkkI986v76j0I2ovoEa4QBlDpB3RNuWQtjBeD6MV4UXhTGaX
NSYga1hWUiyvpum7abCU41KxqG7SFrrt0pwABRciSKTdK2VEOGwGaGy/3BFTUpVm
F3mZ2xxZKHJ9vxkObsLKiB3JKx9LBBSO0vPf29g1/MgYPCqjSns7AEIG79C338fn
t0LaCB8gCehqZZYjD+uah9L/LwnuShlxPUsnx5I6mPI70afY81zS+xROG9pF2p2M
nHCCTTJeszIkx8W6zlKuKUwFrHIu6S986g+0GtUFinoEE07ClJl3aAXAJe8QSUOn
fZQujAiSPgleev4Trcxs/weT3qZv7DoaYstpld998AzGwidUdgpjp6PFzA2moWcn
gOC5Jf9GMGx4+QPfa7JqMkA/HtdGB5oo5gsStlYeZ+VE0R9Asd7M5Ge6G4UTK/v2
PMTDONMjt0q4q+LfVXEmZ2mnwccei4ldfq4PrMIZzxyfBBVG6ZcYssYzIToJMB4m
NTKyORX/0Ntg6AYoj5yeKMF/g2VN47LAsN+Zr6eUoYpkJLnIJ2pqCE58ThjxwC3I
YCmmXA15B3asicFqtAGpXPe4Wb+RdiQyahuTiwd5R9dArR6mUptl57BzpSDnjya9
Ou7sfXh/HtbsaaN41qseT7oO8YckzsoprysKNL7UTMiUV1Pkel/UOZpT6Laq1XEA
M8kBoh4xKo2uHyk6g1b122i7WM8XdagaKhjvNinhF58MyOrorcizt1kqTh2vSo+w
yDlddlMCN1mbGWc+aqWw2+bKfT0WraX8g26d5dqkmsvfYRVlpkuAAmcfNk3jPYUo
Hnr9aJrbwLGOKgJ//uEb3fNYiDl55h0Kl3VlBUsJadB8ZNrhxwuQPOvq6pQafkTq
USCStI2APSzrXId0WMgps6IhiagCEJqA8JFVG8V/okMF0AV2lZPRI1lsSeEyU/t3
lYLtkyoxTdGVuXJbO/0c9ppsUixIsM6eJZGN1qhKGlBERoV96FgSkNopRdwg33WM
PA55eCjZcb8JFTgRJDZExlm+uOcBiLIaG/eYlO+JgRRXJb6s5zHv8fOsvR9WbGB2
wvbm+jDKQs6SA7wjLfCcS2uLQKve53yCF169oOJ1zf6AfzDqDSEEUNVIdbwkX7M9
5xYCXHzKT3+TMj4Zunjuc+HhlIMBjOFfjcYHzRZ8WFTAOa5Mgul9uynxPSplofiE
kLdRbRROPwNgXIpTvYB1/EL6e0I2apus/tTQkQzDVj1RMBn7oZoPsOWxgcjmiVZJ
MwDOW+zUkPGWxMzx3SQHzuRzoCA4ZNQMfxzxvSqXaon1Hc3uvYZ9dwdBxLdmawuC
BG1DTQCOt3BJwWXaCsgm1Pp4QVMa5IOUf2GsETUTBfJfXe1vDNW/y+E3r0Hv7HCW
pvKJOmKEzZAncTju3SXyqM3AUYVPlcD9CAXA9H8R7oYjoazqQ0QrUCso0KXEBzIk
qh0SHk9wpi3YfyMTUKOy8DCuaKEeGxpNJbPeHJZekkWq6IaePmNpOKGMMUSN0WvR
3yLyVZIVU5vqG3vAIACWrLCdKiWz5ZLBR8Rx4wtBTWyf+15fiCgjXJ9Z1mbWJvHY
Umj2ZEDbUcEuSOiL3liEgY3btEPJ9eDNOyiQpLyhzd0bRVjtKu+a7Hr8EwlUGoq1
bfEXh6j5lbni2VUMiT09kd502nwEj0dxSwjaQfXlTulO+ebrHxDeBm9NOAlditu5
Wi3gsR94FJdORgYItE94R60YWBVdtR8L+ehun+WSgMpSBwHvuTS2WdiOFBI2hHjD
IFWyScqcooKeAjl1GtHXaectlAyyTATPWPxxQg5GaJdgA3CzzFwxJZJOJ71S9C9Z
DuWRjWJrWIl95azJ+RoC3EUp2Tp3/MNawif89Ei29+q3oqJGK+uS44Hxc2t/VDNE
gLeWKrJkI/gFcl7jlQlnk5Ma/K+1CRsAxnWE8ZdXvi87oTASp6NsWRw8gbxzCysc
p3CsLpbjygIr/uLps3hE+MXDZ6yjiQs64SSkDOxEZCBJnxAPz5MM7OJAE4NNwVyy
aliX6r0u4JwJgYmQoUL1Dk+Fm2wSK3HxSs2VSRsnC/YAOIFx8Us3H0yFeotEmzxu
ITInH3GlhJC/kRIHHBasrkhAveky7sG2JlIU7RW+prKiUyfL3niRALHDpe/30XmY
k4xjU9YLIrDV7Z6NvrImGjtc5pMNxnP/tQrkO7fymbbzqxOCR6+FJeqFBoMenTB6
ZeAtyZoBf7hQHB3myGaY9wz8I2e0sBOxxnzMlkCaLjeqa83ZBCBfitFvOGVBRDJC
V2e6/P7H4Tk15gF0QiToJ3+7IiRwnYjeUX5yddEbjibIL6SGVPHqiSkIEyx0sdzV
3VDAEw3iHfGtD7GnL3hW9q4FQDctMHOM8HJBlN1zGXdteFe8b0tXJ9F6tKHMlmsG
kniDkiDg0ByA9k307xUIxrniMd5Z/OZ4MxEBZYi8noh2U5SRwhVFqcPOUMzHdsG5
+v6K/3Fmy+jpoKPJte8fxGPHyA/epBhPOT3LBPMW59Ln+K11onXK97w8FSFVslKw
e4NlL0v9wHDch4hcTzwdrAigEoXPIbLeDQF93KctUjDzCaJ6kKQ/AI0N4hNDSDu+
OCRr2ECacC9jppWcIYdUVvHGKprWZvP6AP+OKD3jXImNSUtdEwlMdm/p7qrzm2Qk
ldhgu60/90cJzw9ar8gdY2NDagWMfn7xcZKZrQPcVvHFNMGX16HMgyop9rrEnPNg
uW8b6adBmxcQuJbwnRHpCOOTYPnI+mYChrpZJ9Ph/K0cZ7SgI4zUvABxefrBsO7q
tLl4ftZpVwlKymt9WoMCwD9SG+iRDF2QsEkAALg7BmrVrF5qk21Hd9YVB1YcT2Sp
YJDW8wJSbQ+hZmxO+iyQMMd8z3Vhd/C+bPXwzrAQbKJyEN0TY/YkpnW1vahi+oTh
zwEfJCiTgUBhU9qnHLVtCuH5u8O7tXZ2nLxrhwmTwgY3q0lnYFBAZjVhtFnmm0LV
lgDl3gpt6gGGVLrnCZeJnq4O+pAmlz+49+a9NCp+6V0Koy96xVfxKLU6HNY78uLk
KuoXMMAAqp28dgUlZIcsgcpt9uiAMzAc/pgxNgKPhHX//Upc5tGMUGJOEsVMk1HY
GNg+SJ/34HuIfMeARSaGBp5whjWYAjW1YL1nghRdq2C6KvL1ZM2MjSKrPqDAHKTX
i0W2ScrmPLcobkh1zbgwPematEtf5NcWlmiVqpxB7UvbaWi7lEGxmoQriSDjKaPn
QtdYKE4/Yx1xUHDy0NYSLvKghTI6DR/3W/5TaGPfnEzJP5ZVwrJx4yZc7FSe51Qw
eNdlibuYVdmCD9ibMANLVO3xXBP6ciGxE8tythufVcB5iQoTlyiJjFPNTQR5D60f
TL3mPPB4ZUdzDkuMUiFr/KMEOfTmDJabZ3/caJEtszO5u2GOySM8dTveYGtseA3W
QmB2Cb4FlT/GkObzuaPoXGY3NkPRkT6NoIMFTaw/Id01ZZb5y7uAYQV4Y08mLGEb
3zLQRFoCfvT7yuwLKui2qaybatXKicNZXsBGQgpjQ4jV3UVl9MbtFIFjIsH9Tjfe
4hvlJtvWuVLqK4dOiGYp9+2TReFtFLD7OVDWNEGNUchKkERiWtoWFl0VMpNhZnJp
AjTU011IjYID9A3Is4PlYRhgD/OxcZbgwIYlWiSrU0kJ5wo8MN5yFqH1G940h+fs
1aWgmqrEvfretuNITGrVske5lIlAPAsBRHheVhyhGrGmYKPin6lnRQQ7Lu+DyPgB
eQdjOhWlYdXweu4vyn2ENu6t2PIznxRhWvEU4rPWcmNkRESo1W5tc70NKmetj8U5
Ur75CpEtDEl6GPrgJZKgu1hBFEnY6oxA/hT0EjtXBpO1AAmeV6getXYgrTSBx/aj
Bc8FbH5SzR9XiD/sPUo7Q3UHo0YXy4/BlF+TnittROR3nvC8HoJo3bBAPCrAT+MG
4EPD1XvIux0e4PnJdA63mek/4VijFsj55OdLF31GvYRD8cb95JwJt/+HZ5pWZDPW
S5sFiPzJsAmaSfqGdGK0D+LOo/Zz/HBk6mmRs3kJjPf0ZNINTyp5/TWhd1EiiEiL
Gio73DFLE02OD4ECG5fbRbmQYVa2G1VN9DvJnra3DB84SARgf1llfE7LIC0sQx2b
y6b+19+e41f2Iab2vFUNamHlVLulaY4wC4XEVqgF3oBkGY8mNg1KyD6Pal8zUqXr
+nfKJt2917W4zKy2TGoFPuMT10MzDQb4U/YHqIkFSraPY79HCngRtwARnpcE18r+
lbyThxZTdNdNWEEEUsKZP7oRrOEHxNRfaNZeduUeSGaaVV1BYeHNYkqpBeEoDX49
3NPB3H/m3XLeZBKCkcQdb8LiTfibGJty/MhBhnqNeks2KPsG+WTq5nbDJ3/Zjy3v
5hQ1b+jbY0UZMst2tkuZ92J3nOJIzCKwHOgAT7DuXF4V2LyKEZxgXJpLZ262lAFo
IPYW1qaQVbYG4RlHB1SwNxDbu98R4L83V/X3JswzyRJjZxzSEpcIWGsYFaIqM2Lw
mKLz6EqjAS83mF03/FJ+xbV/wQr58bPr/rarkS3EHsUKc+1a1t+Wp2R+JE4xq7V/
npSOWegzjetyxNcEE97rBp1+UK8KuzsD+DwmP8CUVqlbM5s25rhWPaI/0QgBqdNE
ScZKJze0pJQNf1P2agKRIRFpvHS3+o3B1vqRN4sZxiX+u7Opd8FWL2NE+GLGoQAD
cH8qAWsqJ3xCFsUt2H/bknzrpIM9Agp1VTam+n6vuLTzC7nGU+kIvVBU45Isn7xR
248HdJGGP/4d4bEVEN0sSgw5WbO1mIt/J842Zw8J7jQzUWg7XJRm/b8t+SMR3pT9
WilOFqBiDr2oRfL8uvuQ8QW1DPdtAsUgS+qlQKlKSqcJE/MELZsV7c5xp3hw4CpO
KSaw69ZoSDuYfT1NDGD8lG4LDyex7nZ2+G5p+MWvK4amBa5XAxSqf2IHtVo9YzC7
/t6Imm2EUn6RkGb9DFU4ETvp+gR3wNaFkR7z+GXfsDJecX+dntL6sUPXctY9yJ2n
4JabTQcsDrZYtct/kshv09NN7AXYV5DUhDw3pkDNGlkS29J3J/eX1Lm/of+p+7Bv
r0y8bWQ0Ggt6geYq4WscFQ/i53HlXUOw4nr4rw7SfdqE4IgvdJQfnVVEAqQylV+D
akV1NoQttWhAR4SluF1zlRU+rQmDTPgzIZFwuChaRdv8JztjK8EM2A42xiRLITXK
yzkwd8rY7t8q0LXWOcxaEOPervyCwEYkUGKAYzv6LqhYBDkcZjlOh04wDkJhENwB
GiCEDwY0ct6K7ks1XHd+tJMkZt8giC37WiBoFF4wDSYUibfe0rdbO5xEJJ54niaR
c0ol1L/ZBThsWvUqom5vPZth4Wlwp0mTWrNyzWZeH1zgQRuKnwA7gmEkCtUVVqaL
u6xVQmsfXVSMCHqhol077ndbGI0zEDUIuZ2Q9Y23FntrYGJGarVuaztZOGnfR+b+
IikGS+4Mda5f/jYI12XPQ2fl5HCqb9ZJ1CQNz45hgPmCW+2NfH/soIBFpZ59+9P2
YV862OMFIgF33y8Mt9MYpLbsPvSKxK4VkjPGDvjF9ZJKDKaK26o3duW2CjGvsFgS
WsfcqVXBtfeW6POG/i4tMXpsOa+Zl1ph3kyebR3513RBLTcFotRa5r1BZChYJdnE
ka2pfy4HzEH5FSG8BjriRTVLsft5M1/JcpNJtmBuECHSVTniZZOBgAnjgD0q0hRU
IBpjWMrGQ5/3YhCKgssBgwziCfR/51usK9kqPVeJ13F9TpzW7DHE8LfOcHko33rt
QoM8CCGK7+8niGtpx4a9Dw8SmSQkqb+OsBrA7auxn1/R6KKG3NAya4TPlWD/Iv47
fBF12p50MRNoJyEiqfqnKBKOPw4/+0LnakGAgj/J2te9Z4MMJvxV4KAUQ/BzvQDz
BTxLrA/7B65ijj0yU5Cl6xHYITvsPp+N1qBZd1LXELRxx1lgFXIhVRsmCjwUjY7S
cm8kHWdjwmPHL6eKB7BZW+0kiZf9fzym1RFusyN8LERurz6gP7SfS5WapoFkGOlI
5f2MWWKbgP/t76gWT7QR4vMs25G0RmBYlkCeb7iNkb7nWB7CLMmeP7H28GhCFqet
rZlv3eaFIl/U1gKl9bf/zaJz0KQA8HYHcQhNhYyTNko/UDf0nZUeiL/vLDpac67J
VtZ/O4ISvGatwl14L71ngbYar4tvYcA8pSkfYY+3ySL1YussaHWgSSXsxdqRnwVv
2vLulNfoJV9svrWEvTXvh/LgCVEWc9kHQRVj3LR/RQcC3w4i4Ff99tRXTyfVIokv
BQo65Cfq40+3bzpeoQIleeRoqjdRF1easbUaw94Uu2AKAcqlY6MWnjDZV1EIEhdB
XRRmr/fB1ldm9C/ScHILuWo4rYWyvkakv+SUOdKIQtG+rWbv11AkFcBEEqedGnKO
80GWkC7ncjT5Bu9MJr/SjlgxZHNIMhbLUy/W4IRh0wJHX5nHXnTZ0KOYW4XZumRj
NJkUdlkWx/QedkMsF8BXqRwHErXedUGCVmo19l/nMOpBWXD1x8cZtFAR+GXU/Bm9
4xUQpNKBTAKi8hE1srgCJyMj86Zn5wYMTnNwq4QTglyB6LmLMhpOeG4+/cLe+Eiu
CTW65IIZPllNxtnTsnd9WRrCaQcNCKdr5/j9IOWTQ3bA23YbUpdX9s5B/17+yapJ
AnxWjer+zzTMAETeVcEFL5laBcbwNvwOKKQykIaBIebdgbxoGfckFIqfIGOS14qe
p5WqszhCM0ueQ+iRVkc7PKrBzIr35cQSnVAWom4iel3QJaK2qjgE/Yce+CA6SUaw
C9XGZoMJ30dE9OY198dKYg7H1dTd57YY5mbWSM6GuO7qm7/QTfqruG30ru1S3eRe
QFI9HkRG2jQldFpDRtY+rQVXnCPRZzS7WA9JaHEPfCYLUY0hedZ3iCkOC4GGKC0B
cyLRYQCl8ClHtkj+E1ceX4F0QxbWkKtXBAQNcws0M/IGH0YlyGX/7rTY+c6h5Edy
nMxJOBdcOD7B77VEeqv5OC0NEMy5bwkEd0uK5xCB0tMc+n+58DZZJ99r4i6CEGmL
tKlN6tuR8x6qbES1++X5rFTOh8GNsL/yCLqUzYQFgYvRJJXc36twzQSoeTPiUZDa
jvbAYKS58pDYrw6as5RR1KTMHnPCmyoajgL3fduLJCXQiNq+C1U9FoRKOlix3Se8
kMq5aY7RWsAhpwL0J9YBq/Kgj32C8zT8RARkE0Fzm6Xc9Aiq5kaeK+PURFtB310E
eZ4yFwxbh1zuZkEpWGiQxsqs1CUIUalrBV8+oGF+E3TN5OPx6ePZaP1c03wnSQNi
uS4+6gH/l8ghRwJbtbYK9cG8l2wCO85/Pz76bj1f+t0K9GY6mQ2VSncJmE1NDmgF
azB7lMpDA4KIvdFdelaNFPuEsawafA0LhpFvzYcy41FGos/J/pLwZ7p/KX26OJea
q/f+skC3p9HBpz7nSPyZEBbocdh+ae8SLleaMaiNekE21i4Gchl3BrqtIoerzlQi
AIHuk2uUyleFiWTo7h4RGzR2jJdGSYLJ4ujKW9CoFfZczySgsqJgwmQYkiPnWJR+
DwJIb2mz+YUx5S8kGsboJDyK2BdmdCJAD6aKB/HRNVOdvR7ss2Tp61u0v/rLgzsQ
cdgliRlCCCFWpprz2tFRduMNbuoiSqQTACn4WWvDNSanWda5I7RMkmZ6/MeDBWQI
7yUoR9Jtw8rBOMzuaPtwfMAMyj4IDgll5vec/vsCrF/mxbp7ENOJZZCRWuMFe3iZ
FRYTraLu95cvX7AhuFABWEiknLRQKBPiKMoRkd9uNYiqm/brxp3yCYbIj5KcGnB4
64u1mE7n0gQ8UXai1Kz89jD4Rcy6eptX5hpJh4+3rbNJgsr6Ve/p/51ZJcqFEy4K
dVN6a1Phs6HWlqpV1fOCuHs1wrgrgNyZaonzvLmZiLUZh/8MlfoXffs3oIx9/HZk
5zrZesqrPJMALumDyfoAlyaXi5CfYIqLkjlDK4wj9vBYQ4kELQUDnVJ7ePzxZVEi
TvDJEGDV5pjPBYcnydaqbDvdbyeUmJs3n5jARR5JMeFiH1hTqluwJ8dBGQmT99NA
GMAYykTVljPx/63aC/YvRmMDRjpcBA6ef/Ni72KsMByJqusdPoWQyTbN3kpMRuA7
bTJXyrpjZqcQ/g33nDv52Nq1X7xnlTDsDmV8UKzmoDq+AoZm02ZwEnnoE9M9kuGG
kK3hWk4fjRZhbVNs0XXhT2tT4lYjXKAB5EhTFB06eYiykJSX9LXCJe/Uw8ukWRhq
7fvlfesQXeNeZNUlbYDZxA3KSjMHozrhpg9x4crN089rtY8fuc3kylxFKejvns4J
je0GZFjeofamQOAlrMUEZyPOq8QvPaPr2sq8X9TWEIZ+JEWUj9q7jlRMYLY/IHI1
Fve5WsPM5wkAWtWgW1ZTAWu1HMSX6IkJY5kJhFaM+FftcvTrAR+KH/F90mfBWDyV
P/alOfNtOE5lUh2EUzn6Np9W4fmqRxFEQU5SneqmMC19mVOUWG7B7/yT+hkw3tlI
4xzmVUOTkEjKSWC8thBRy/RMu5F0Dzbtna6T212A+m8wnxFmHpOf9Y+xiE4AZM+R
0DCMQOe9N7gTzHiSAPCa2R1p/EvDL8SsIphVleAPH8KUmM7le5Odna7OGvOJcAIi
WirL0/BZL1gbHDN7pC7SyHjP8OPQFyKmPQAqscFEYbyDgdmqGW4T1rgKZdSwaQKR
3R22fME+gmzr7HoiHidpwnM/y2t3Kd9D5KAl/n22H1bQXwnBicNPceWBG8s/qXPb
p+4DOZHDkMFlc4B0G+hxfCkkFfmpgxmKH1bE6mlG4kQo/XD4c79zAwBZBE8PRSZp
1n6x3JFaLTcT8/IX6PTlJ6rYbdLTeL+lDKBXm1C5WzLIKhtSKzVdnbwcoyjdWD6z
Qlm+rteh5TQkqrMh/2Qlp/Cg1JeVWOP9KVM4BIG3lanOsDq7dx2dj+BKc5GRZpw3
RupHHFRwn43H6/iDDAzHLsL2KvKyB1IuA6aK/i8t5o54G0Ho5ofSnJbc35GAYcWU
+iQDfLfm0eDMGw2NAzg4VkRoi1XIUMSizflg4CPheb3I6HyrSW97C0s63OTZQfYb
fiCB+W4LsoRoDiijwXyOrrLO8bijvfycXVlp7q2AAwTr6NFtH01bAgS31E6URJLu
nTi6JBT2jU7RyqeMaulk2acQ4pVTvNtgYBWdwni3f8SWSKo3Y2NhiHKu4+Ad6oLh
mHSYh+Why1+JVWM1Rau4ywLdSwlTBem/2C49XgdL6xMBpGK9cxhEjlQx4t9r0Q1k
4qhpFnjy/8VZEUhQ9pU9o6AhzlX2xD3o9M4m7jq5rfnTXepqSVi4ji0UlCwxbqFY
MmTkwmt5vOXvniRlw6jPrStdNXYMRe3q49uu7R3iQCIZqgdHBUlcheob8IsD81/s
6u+QAwK8tb+mxK4w3OYQQdD19u9GO2t/47W2p2Xdr+FwfnPUDSIP5sN8KPMNGkXc
Usg4U1mwNfv8MOxLPi9Xr8I67BB8IeM+975DNb8rr0vUEeOL6gPNPFJyTzE/JhCd
EBq+98h99N+J6HUuAzu8x7LE9Ng/unL3hKvbMuE5Azgbyyt6EJYR9eYjHGXuzh7f
j34WAnRXcGtnfDjqwK10yJF8kYcq3DSNoWyPGOIuOegq5Gt+L2F7gcEKvbt+RHFV
rQCxyiJO3GkKT5dT49ligpbGJny7SEFsXoSIp8uYopKMVBhHf7pMeWol1schxdjs
ZC77rPcTK3gPWH22ukUDmU/zptT9+kJC989G1B68Hnsa6HnkFBnnqB8RoTolLAnL
pkFE7w98IXrp9jy23K2Z0LUzJB6u+GhOMinZ/cjH+AyqzO8eN2bgEnMF8XrBFGsb
c2kLAVH8BBiRmoy3eJCTbipOzXT5DBALbN/b5PsV/5sUrfaX1iY2a+7/2FN4ldmN
67SNBhMxrsT0LQ/Vrfgu/pQZ9AZ/dX/OWTwscqFuVbnVvUtDQpxZ8JkjPmT2xbkR
xigXx28xT92QCZpmlSqPV1oM/RabqneQZwlVgknNojuYLvAshNB6fIlmQn849kRq
2EfFNB+iZywoEFSjTwbklmEHjEh6UbNgX0joFgWtL4reiU5pGiYis5FjK8vuKuaw
lEwg3hMKMHMhajTwJwWLUQxf7x7FS7aBHvfOVpWJ05mI8vvx7XpW/jUevVhZjREH
b8Ca3B6+2MWn8kugdQ/ZdgvPd8qu2vZuC0otJvDp6FqQ9Pnz21jT2uO6zSTj8+m3
3fSVg8nnHg8oIK5OFYf7PIAAMz7sN5J83tMXKhjhWiN2+c7YGyjvuqExMXFbQHBh
gZ+G5XR+OxL/gKHQa/lrQFl5o4zhPgpo86/x0KwXk8rWarhaX97mPWAii7R8fg8z
2GeR7GWmsfDYSzuUUUVAQrjeG8BmCPvOhBQsJEeh+TFy374dy8qVD9Z3FYx5DRVg
EpohJb/CEE/CpF/7o0EfZC8391BAepUn9vVkPjOYi8R7fNh9Ai9mTj4FaFONvI1i
81DC9GL7Z4dZbmGF3n5dAwsZHyzxTNUyDt62lE+xMqSauJmajNXmqhu/avx5b8Zi
Lopfwq6d9sMaCSa8UqxwtE0AeUJwbbxKueyV/KxblWd4oyi3mhYD1BervnKTj9ja
HGtNw9X4jIg3tdpHHfM7xmIsv9dQHFcBFjeM5d/p+lB6/AKmItTb2lMMBQQITaBK
f42dlgAhfgFmuyLp0gBAFkNRYCdH6+6LlfRABVsh7SmPXLyK1lcwRS2yCEpZnG0w
vs68iHF//A1OgMXDYS1fcNXdhqRVQvc2tzKXMfT+alRWBo0sFEwRRj6WT09oLBxo
8wKArP1bVbJZ64bSYtY5ehBrPm+RNIRS+SDGyP2sMsBTHi0YzQol90UNUS/8Bqso
uiiXTIudUO2lMXiZH7WOQpfV1fgfypMc1ROBqcq3UG2xHLM4T5nJE2iklnsSXYVy
s+kpJtsWoFefkJf1jcie3ABfJlfQdrnlLf8XSbWgybp8oQxBbLLENqLubMVWB+VA
NeFDzeoyuJJJUGjn2prPpYV30LXeO95nH6jGyOtsu5+lHVIWIFu34bdhSr0dIUjl
t4bizEjy4L15jBAuA/oVpo2Fe0JilNQpbVZ4ljaSKX2vbrR9mcpJM0g6KUeluTxT
moVcCkP6yVHeX3Xojs9oKYMOLFmSNvAqbLAvqVvI3XXou8dUfGxoYuYLJqavakHM
8ElsuVA1Athl90lcGYv5U6D/piABto7jCjo/8B76eLvMDdTjNK3yLJp7i/PR68Hf
2rQD4jkKwE9q76OFE8cO34Y2ezjz8KPOvj8QcDCdPBID90/3A2srV0o9/Bbl6EkL
Eb2Sxw1CjjBfpgqwHtIoQYqvjhc9PbklBo5L40mSnV9h/bZRRTgR+JCu2Sv5ubYE
+P6AV1aPy75kziDKHAMFsJHZmw1NHr/TTDnur+rzeKXFMBQYgQiS9taviVs86F41
73lBaB97oco/5Tg+lxUdb1aXhL9uxSCG/fnP0rK6N5BMIksFfNXhR7fAtds2iSNm
Kgt9yZqwjjNKpwy8M/CrZRQRA+bR5a1WIJ1YwE9fPyNLfEKG5L1vFVY0FFLaj1k2
XTbSE4UR29sv6BW/rdl7ZdJbbi7HMQ28hwxvCDaDwHtJ3LHNsM7Gf+HBKEG/PmQL
X+ki+E+/A9ym1439/3a5uakVEiJ8h6GJfnRfnz7el58g2YIo4F8FkGNbVt2rbYyF
oi4Zf+gBxtyzGZhCql2kzgKI/45wF1FDjTCKppqZNmKfH43IOQwRvO0jroZMfPjX
6tRk/lkBgt0rxPkr9/Yt2JZigVkEJXuNAQ5gwOBRYkSHXQ/ntgQzEhT6r55NyxX0
Dgop4e0r0U8SkQttVxOYjyZa2h/SBR1gZOZqmvE4EtUAp4YYsK7FwlS0a8MLhxC4
pw0sQGM3nTm4wXXZ27tAXI+7xIuGJccVfyoymxzNjIaqcPb5x6RCE4uTNm/3Df15
UadxUiBaoztXcdG/NiHEqrM40EitRbL+G+0SN1F+sId77WqHvtzJQGsh5z/peQ7B
K3eBAdOEebIdFpH2Ec2yGgZhIDX/z6aJdTtEWaeC3tpjPaadT8qKfT8Q7QMMJYOG
fRaWGSuSRUxBya7yzacTIGbqM4YFWbRq3DxvaHW9fKp12MYJE762m2AGKMQ4ucv1
GuhwLB+OuAQyYuxhF/WXxw6TlF/ATpDKEBlr18pOFTEABtqzBZG7uTTYSFuq0g7J
5hRGBtFfqfaDZsHgfVUaJsN0EcQeAoaVcnHJDLrR/qBgM7WEYf4rdqgRREg5bmat
/Y5jCGEJRVU6vfBo9PegVqIyYApvc/IuIFvczCv6EpBiKFMrGnYFgqeHFHoxmpfB
3HehOqyMTgcsn4r3+PHGD5KWBDQqigEBlcuHjY0FO3CLHttIynUZTEs793wYgVZz
cSxGhXMRf+QvNrJAzhGd3sNjOQyFdT+3Dgc4VCPvSyH0FHBm7OvMJaRxPBcAHBao
uxb6vod+ezAZJX0dpdq0d07wc/AiGAQojFQQaUerxtZJMuAPh2dIbYjhZ//SV28B
+g0kZpxpzsrI3/L5jkA08+m+KmUCh4u9Tp03jnayDQPrneTyfA7rKLb7Y0wCTwSB
3jeuIaLU4Z0c82cTD89NRwhmL+P3YnLln1FLwKxvFIe8dy5X3wHTUn6jLMIgBmuF
SxpR/sn6f3HbLVUCqaoeAkMwuch+Esd+T41tklSTB9GteY+RhL0zkqRV/nNTwSwo
iX0eZi2Mqi3swUkyXnMHbpxzSrS3BwJP4eofsn3p2aFHwpcw3dlg4I1/MSSoyySx
Gb+WBXXu2DSIrKp4k1ZLAq8A8SZQSmmFis4haAzgGd8d3dN7IsVRGWEU/uBOnMA1
ApNrjb5KC7p9OWrNN4q47Ktx1rQcJQXay1jCPtDqxzAhspA/UFCWf9s0XFREXaPm
c/C0tpfc/7j6QBM8pbOF7aLcmMqnywJ1CCR9x+zO7wgzPZOfQSN2sKWI3MAQbgfJ
zi25ZfLqJZ4S9FNo5mGSUG00pJQiQqsR2qqbCsPT7xJ2Maav9MSqceDrwYRrMaX5
wo91mmzsZi8LP/S+XDpGTH5ovbYYq/rODAPQRHir0k27GBidTTSn53h+C91gKM3Q
mfyMNJ9xRni6GOjNxRcn+NBy5T+YBpcvrFzOdLlnuIRdv6hsSmZVHrnYO3LH7dEo
FMiJDhuWWAdNJLQxPiYXAvGLF+v0tFMba+08SAY+43KY5vUlpvFv46mSsSQvXWjh
Kqu6JtHmohK+QmokSz/yHsSAPPuNZo8/ZyLRPeXQxWRLH4wq7pw9SqCzDTMh8lGP
Wj+Rfbam8g7iO4pl5IGrPlSSR4H6Z39TZNMv5bDaW2LNLDRlfkDLrx/0IjRsuJBO
x3gVWiwrX5L4MfZHvFY6WMLKar4HYQHA9y1rEevDG0an85Bmlig2rQQn6x32BuVN
9Van+lb4HKJNRDz9W9F+iDcQWi4qYADBLqBwyWnkB9yRxxytjSTRHbsSj4zuTqb7
axYPj80JyRGmBJsuYXpzG07x2NVZM6YH0XuHt8b9abwwjTwz0Pzd15dm//5FG87w
oU1SSX3CJhLMs8gzef8BTQ9e9dwG5T951fa9m5HFpxprldbFpXQFiBA6Y6ysJ5s+
9Me2kJtqKUOEgxSeATjIiGqOXUkEjPG+10c1Jh1ICqh89soo59eM1zMeLiM1wGQz
8dEOGshO2dKSRCvQAU95yeLo8I9PGS3zV+pAInCNYHfb5FMeqBA3AehFz6jYPCIG
gizrsAWBG0BxPmMma2++D7Lhq4xTs4iczxXqk1SXM9DGETcJgLfrH/eDkK5P0tny
9/9rXcPEyQ3h7dO08+bsrYwQ0zYNDu2kYfDrf9mXyB8awLV7NOncsi6wiYadw+7q
A8mVZrJotNS0zyCVUc79msWLX3XRsxJ0PVS05xvQbu2MyFc4wfUGeN39GDDQhEMo
O66ZplNSrJhdCUfPDyWczovt6SOpuSifnmTtoL0aDiUBOnnaf+YViZk3w7HJ4fAO
CsKOYF+/M+1KLRu5RTLoHrsxnWO9ecPNkRCZR1Mk4/cUITReETUhjPMLjj59Hf0N
APQzkeq5uaFNZCkacYqr2Z7SmtcjHDHJaZzH4qg22CKAZUZBep9uj8b3TpZL9Vbx
PlOdbMkXVkAzF1rf9rgrf8Hefmh2uAq1W7835lNcljgeGlUH9bHVm3kqR+h7snJc
9vaGd6xnsxRr/JdNSPZ8cv9Wb/OiazfB2HBqSSgHPgRfdZKFynUJcFXXKXZEHuQ9
QFq/pKVZG+QzN5qMFdCKwb43cE0BsrAuDKQpg91vggDfaE+FUbGWmM1o46+L8pm5
+nhnfeW8OcMv4dcDX9YeLrofGR0l4qcrB4rBOj847GWpNPK80XMy4X0sRRR/dZ3N
5T3bu0DoYV2RSW+MnX6nIZy/+7IZpfNinkCOoyl8Qlb9Dx2F6X6kJYtmsW9i5z29
B/YAbIupMCvolomKaD+vwExJ2pHWsXqpncSDiLbCEhg8eQT7Y5QNu85kcTCJNztO
xjO/FEg7cOweQL6B+U+b7mZEgxdY7tPMeH7iYtQHP5FkqZLydWt/Zgx3sDstvLOa
is7YjChN9ryF2IPMtZjQALwervghSBzBuJg207kNqFA/mAkG6rRXzrcKxsIrTQQQ
cQq+F+49z5B/FLUZqceogDYhBOJfZOzhn+dCxYr0QVKoGvk9PUqoYxvtUacIEXzV
46y6+okUwxOp7uIN6SHLArcXeWzoty52QQRN8FIS0BLRl3Yq5lPxIf5PHWz0rXsJ
2cf+SJbOu5m0Vo9syURICjiIFWUAHIlYQtRAMBV0aFYlsxNEkPXhvoTt3w+Qr/ta
RweXPTCn2xXx64q2RsDNOoJEinqx07eyiHPafvZ097/sQwxxXm8baQ4q6SvNAMYs
AZy0FI9ScnGifr9iyBZDCkdfi9nyUsYprFHiLta+E/TWTUYkVCaSgl9mwH/23nE5
AVuwzAMEyHzfTZDyYj/NeMrBUkshViq4gCMG6UzGM9WbIMfwG7YqiCt3/9eAA/za
Jew2QwUFM7PM1qMhUgwQ31jUeYPGs44f4BqMjoD/6lpanbrpYm5rpLSFPjfebVec
1uSl9h4j/tQ+OoUHzQ/ev+wrYqgF80yaUeSixSVhGN3R0o7lGiJ9fr5h5l8F4GhT
vlSHVDzB7UAyO21qheLgIq7h6qMcVnTrH/9FT0hJ2nFdQ6x7QEpUCIYM9QTQ0RA3
3tTsfaOH1j0xnVSCejkVRA+Dth+LFoRIbb1vct/KQdtAThy3+45JZSIqdmT3nwA8
/aHXrDng+Xr1frAq7HYdiJfE8HCBsLsDt8H7ajMTNg6LxAkfTat23RneS0wi2bEv
dnPCq/enlLau3+QuvGwpUp0RI4TDw6y+Y/H/B5BEylx338dtqeh1Z5WqJxa5yuhL
Vg8N1s0NhqsKu1LalYgu0uZfq7pQIAXyN9cWGWNRYzVlP9SuktojGNAtdn9NOzku
Ne4B99X4ND6XS1bEpVbrBgqWB0i+4/5NshR8csdq0TF6rD2nOBJ++DGFhvzdI66V
JgdVIeV02b663tPwI83nAYyjDl1qtHJKxtEgh3FZHD4eFTa5sfwGC2yQag72Cdy7
VgqZ4Mg+OrPZCF2uMMzV6gIyJUt1nmxZFk1i/iBZJ2YsFEgnWsdZ7jT9fT+7Ci6E
ro4e70AgWkwPkk9EyUv6dAQabhTDYDWMCequ4wSvbIUCr8WhoBmGPn6aRGPqc1t4
RSTb8CHLB73U6hIYo+eEEQWNSR2VMeatvGzrrnoIashVdIHQwg8BezIc+sAkKWKR
M4xf8tnZMpA/rS7qxPGBpD6Jd9UuJEgGRYrzHInNps5heemi9CX3evM9pqbVii+Z
Ciu3+6HqCrdasdhNJ+41q/sVK0P8qHsp/q4025VfXfxNtSZo8lcfCWuH13pmZcIj
R2T2/g9IRvuIJMptf4+EWFo9SBvJtY3MrAU0b5n7GifkR4t+JrwXcq77ND2jUh2X
w6JMR40xc4PFBxR+KWRtpkT9Z6+AnneWq7EksSuW/tEMUKtT5FL5yj4ZsvQ6CrwQ
21xDBgxt5W0ymeJlS1am3rIVxUjKGpqn9hSEis47f6g+xlKTo2KjaXZUXAh83srE
KD8RQGOuzVMNNCvyPjSz5754KT4x3mZWjI9Pb6J450kKxhMxUFypV/J+7zOi/x41
kmkqOGX9RPXRLJTTNWpAzNQ3yutpNEfRHXaJv2seUfArcHYJgQtV/BhgkyrYoruf
AuiBe11sRgvmRH7HXNeninr9hybbP7CSUeobqEOIDZf4ilOqGmRq718xoOKGUy9l
g+LucwquAeKmnZQhTAmBHe+cjrQffN+j96fCbQYjFKngIUjbSJrftORwQs2tnRdk
3BpuntsGTSGuwoYCPn+ciliHrTP1WroysD4PCKXb6YbDYKKNKq5+QFF0+ZbqZ7a3
jjqgWpPErY6712QeyYafULlJN2gClIr4p+yw1tMGUGGEyzv0/oO2+4ay8C5Q3aae
Wlxf1QWbWW53tKLqHWKublqx8ypJPDyITYyxLA7D4GZ1nVetZrEd4Dg8655auyEq
GjL6q1nPkYhjy83jrVerT+lVlhLNQF0wl3c/mfq1mEfaZGxJv9Lqy9lqbv76lk0L
uJuVW7r5wdXse7fthRkGyg+gqf1Gif1V43G7HBi/UaieI1cx2Qhja9SjEkcQako+
gAvGnihYgmaMonEJY0p97GN9Zx/+wXtRiFyibzaZ7t0Ra84BQGnjR2JLgydbVaR7
j5tyITPDC2FntSpJ7VdfuhgixrLS6NOBQCHYPKxIR3xZ0ml2LS5S7/BZnkcWr3Fk
4IAH88RoMNkZ8a76En6sKmq3aLb1zr0IlQQk+J6Ltr6di2fJtySQu09z+3QVS7WS
YYHLyjPXBK+jwlwGKt7SSggmufE552xk070i5U3EhzujejWqjxHwf/HUwLv2VavI
DzfLXifTli6dunra+xh7Ep+iQVZ1akjXv1aNNbcmoowG+NGOJ/VCpOSiL0oUTbB1
0vaXVj1ingQJKWEE//5XBvUNZ7UuJSv/UmL+cxAwKD/0YII6CCmWSTh1SHSJ/7Fm
CD5EB4uNdEKj21OE4/K21QvuFaCFj5rcSc+ApDPxUw7OULdLm24QyrRcLkHi+YF+
ZC8OK9/22FtbIAgy9l74OWW90FxzKW+4nLc5QsE8WLkkZgO4HWtWHfevRbF57hkJ
/Be9r7r/uLKan58lei7NhB9bmLBKyw7V2rZQlQhGx6F7eDKFp7rACt+8inh/Bbm3
xDD6rv3sRYUhEfdrgBEl1M1EQLJaWnBqYGSZ9ptqHkE4RnAs9c2nankCKJgcJcNF
Yk4aTqFkc8Pb3amwlQLyHMO6zLK3wDVbZV48Ls6Nti9jeDNLpAlCWujDAB1m4d+t
6fAw0lw/i6J2mS3t55fnJKM89mTfQik3BYXP6PmqAThlQHb+7x/p7z34FFIxKtZL
VZ4/KXLM3Fm0cGrUAFoSdkToGclt0tJHyQwnmYngT0B5k6kLhRBS7vYLA23nqL+0
qTOd1UfqAbZrqHbdXITTI4R9XehEXzKLNQdSVQXFKcWt/7G/3Jmkf7cdso/lDuN2
CssSWBB/tpu2AEptIVBgcu2jw26y6eq1ARG4ugqLDEL93ehKuUclaAMbd/Dte12r
5L558BwVrTG9MoMaSsLCo6BM7ooWc+QVpQv7bWZCFOtZfTFk2K02h+F8W/7Uz9iZ
IP48m3as992Ak9JWGGP8v3jENWus6fr7PI0AwnVaVP+bm2FZHrwjEn7dsX0i45j4
k8GklqT+1KpLWeJW2kM0+WnxbnyRmryxoTZdWU1UnAw3PfPGL7nHm6PsbEk6KhwA
+LZaeg3iKv2gKMbhEqq5+3AydKNRcitgo+XBTKYlY7oB6GFdCijRWaURLdWKOlVC
Ub9pHjI/bPzVrvzD2iwHXaqO2ZVYuQ0HZae4YqP8cQaHWgyJK4p7qtekmx2xGrMo
n0TdsgwKmSWkBE4s10aK1WYThkcoae5I703ShAnLR/6K5/xxsR+DwYCVEtGIv8Oz
tdbDtTsorWTBqypQdgUYVnSa1F8Rs03P2SJbDtuRuzHi3m9dtMKzo/+DhO5rINXq
+29RTKHMxfD+6SJ5bFCqlygJ/4AR8r2aJ/KlxRzVt8mVVOJJGgD0nVIkW/CpF9T0
aq5yzDk6w+1okiLx9HV/UbAYXNUpkG3+jfc3TjEJiShIYz7Mew+Ivt4XNckEJKHD
d/8jtSVbwVp3DW/dO0PHe4ZYcRa78cmCojCHGhoAt8lhJfSGOjSphQuA/L2ogZY8
ilISMw63ZQ8N3b2/u57l/8vEkppsCkIhllRRjaOnzNQesntn53VOrkuXvROgH4SF
3UtvkVc5fw3fhUBOHQkbkPOTFbX0eo/oFtg7NWp+6TMzpgi5wihW0/28LoI9h41y
giivpfaxr12fYSyWudrMKAdYodLNtwBiIWEt9pYRFGsDVZRh045wUe6fi2VbNqs8
xVWSidCXHx6m6pj4QC7qUR/OnxMN9NdhgAJmfFBIIKpWHJX94iX8ijQCs1EyVEZx
BaiaRjYEjIklk42zLubtMoYT83vsoa+t2WOQ69lvUmGFoIOQp3n6hEKbc4Y93bpV
ekDHZ+b+nwHVJ/avwwOGJQCDB1EurlNFa9SLAdWGDhjtGasHKtddfZeFDV+SXBHv
pSpTblZBo3/TGitWtER7PHQiDZYASEBCmVSEALXVvhrLBlI0xTSJNDpasxoYrN52
wMc7SrW0O/zs5LA8V3YthhjV/fhXjbuweVRA6GKCBSgmVLzW5LZHBl8LwkJKncNQ
inapMU0GtnGuEYx/9jNpypClhkfJ/ecHvRcn1PA36uc0v3aESVEZQDZUe25Nlcn4
Z3zVUVSOgG2aw/TwMB+qt+N9VcTE1NR/K3xbe2Og5eVmoYNv4LG85keknsUtDxcU
Osw5607nvy3az9ZPbeacMadmuyupAzof9EOCasJ0GRurU33mg4V6Cf4vQEShCJIH
NiLmKwzr/SeSexy6hal1CxsOoeJNbxx03h8Y24KiAtDi2XU2tcEHr7MyXP/a9Csx
xIFIUg7M+ZNPhwtbV6SAgyTAzIHW6D6W5Ad/z2FTUalaBtiYLHyoqcfIlfBEKpgA
6xk3wsyrH/ol69+UgfXVNqnHLvWE6kp/Au2oQx08p4P1pE4j86WQJOq6euwgqBXV
5/+C18SYWawpy9UBhOps0v1gdbAzXuZFbuovy+kvZbi35GZfADr1ALl2hS4MNBds
MgBLTocxziRj3SwOGAxayzZCEcTdyXCvhzSCK8ysBAZftB/2+2Hwd9KeXWmKWG1+
J7UAuIihHfjgJck0QB4hZVx0eMXnuG9GajVQCq3IpasToPcmLhv3Zzo0timoFdd2
Ux7tybpW7Za/kpDY0VZzysIPAlCr8Qp+aF0BBYq90PfrgBE9TCowl6fCxW66Afk6
6V3omVXWjm9u/kpiluzGa3QEM94U8sKUdiiLB8ziDIHIaUOHUVSoUj2gAsaDfs3Q
qQTGdv8bAcefUpMcq6mROnCEhFYqEzyN1xsqtEKzHVJvxrJEeXqHlChVDms5291b
3zG+GaHnZYn//ziZj1k1xf7b1FXm9W8gxDNjm6G7bMTF5eXvrMhf0AKW46pUUzt8
FHhhbXybMieFd/b8e3ApT2O7vYnkaEDtFmumhjdME/iyK8L0SQNOawJvcKxXXSDd
dcvZr1nszkUUB4kBrRY3VbUyNkx6FuBdptp86nObRLA2ROJ6Ok5lVClALTpBAtdT
N+epUkyt4B104K3piG6/D2PHpTLrR1FyqBomlz7QT/hOEKqLYPfwxFxys49jKSiO
rIxQOIldqXi61XaNRO6egfbWBxHX+Gt8hIx+ggoR/Lxbfx4+6vNrDJX1gJDmL0v8
qzkAc2TteIolhBokkhVpvcxp4+brpSQSdsZWVTeTxn5FPSuXVoxo4F+ZFBxy+PIk
zAS/dx5Xoe7Tu71y9DfsBuueeO5LZN/Xf9d1c7PUc1iiFJH7DIGRuhB6g/E1gJvu
lD3UYEGAAsLqzJIc4Gx4f4nLL6U7BH9TIH/WHGK8M6HNiTa5gpYAEDW3lc5mz7PR
/wNTU4BMsaIBnc+ntL0hm9VWd5PIFI9X789h7voWCqe9iSaUTof0nOj4kR33EcPB
pnBuu2OuznlYz0grgtfdzb0jBid/Pdy0YOWVUfA+9J6MmuKYVGG2PCCkPy7GX0mt
ek/y73RkylCK78gRcY9jb5ieJx80ShDmLRHlmhwR6gwWOMOo7Su0s2WZu6Vl9rzA
5V7/pjob3vyTQVnx5il1AXO3gZmvTObxcLUhKRD9HKvAxtxFxqQHMlqUaodS1T5R
ZQJ21nE67taTbtPpckdhsUbee3RlyzzWFaBgHyVbyQ9twgRxtERapdkqFRcSIE8n
pwI2rksEO5Cckz8R1b1fFoy99T8Z4FUpMK0yZ4BoZswLOG380RBgPEhRG4YXRfE6
rwide3WzVhgj4T9olZzfmfPpJi2bVBPP7IbG6raXVxDq2F7vTyglSMHrlngsvwyq
aEmfhAtZ6+cfbzGBb9cIhZjUhF2yMvz3/D1J91zG4GyTXj3BA1EWTXQuDQCiNsfT
c+t13T1+JK0uQSkn0kodlyx1ukQFJJ/bc68HfWJEyw8QuaA1aG1mJ/UoXKy4c+UR
Kd9BlZCDOHPkYTdBH6EgRktbPnmIAtJYH3vMLAgXKuWH3/sU5oOX6EfnA2tsCR5y
GF9nw73nEW+Dd8CUCuPjfH0iT0r2GaWXdKoP12pBgK3dCyRj7xm6Wm/Sh6yprAQe
j6quS3Br2vx0gGGim3Kb0WE0UuBjkrzQv88oeJc670J13eN0Y9v6w3GoOGXos6w9
nulF3VCI+W+RWGvR7PUi/1qVvP0YxRJjlWi4SgxAhjFKy0cRVqnS2h3EDoxuIClp
bI+Q3aHx2JguGvQNwk+AdVFSThAeAltLGgw3FZ/2VpRiCXeLnB7IXl1Kn/u2tcUH
bFVqIav9aTyF68okbkYyecQiNVX6VAHNzzGt//xQXPi0grbsoK25Vbi3KjpoQqFY
fCx8dL1PO/y+iU7aMY/u1L8Tefl08cawZzxukKMiy7/gD1It2SYUr4QW7UBlf4ZG
hTFogsrd9l58dL1hvg44JYEzWkjYoDcmSFmGUo+OxgiJM9Zkwt9Ai0a88h0TwdgX
YOr/XoRH14pmG/fuCvvRh/6dfRRzChjjeCwqyBG2zKAH9gvR4KbCHmK3H4GeHEWP
yQM6TQRvIP9epvC0fD3+QD9Iq4CALKoGIRcNJFPI1lk/jyaL1UPUIB9aBtFJ6f6C
dQoQPtyMiE6YNJ42ujN1rocsNMcpkE9FRl4XdMbO3aG6n2KI8Tfi04Y+xpP5V8ws
wuyfZq/z0vrfQgx3tJe2s4l1FX6ZGQ2UDHgS/bhI/xrG+80vSB/x/Ug26h/0AMFV
SiGBRt9KbOXZzcP3i2O9sYEIP56/2krU5oKiSIjDu21Do+f7QMXepf5zCt3qkaL6
3gagTlALFhMR0JIsnhGkDhoa38RmZ5qKiSMsgKHVhaTQNuKziNKgbeYeG57exZ5+
KfPTDAA/zvm8W6i9pqjZvARP9Jr34ToCQbnHgbNcIRpEGVWg7nzxxB3rhRxzRvKI
+CgqAByqDPA6S9VzCbATtIHtS1R5uK96HyVe4vl3IEBHTcYZ6mAeK1S4LCQ1B5Ej
CPHmkxoOx9QGLVoN+WA6aKUJZlA5EtNHcb+UVXtdIuSdSsWYUDolbmBZqvdc3C+o
iwbMNByi/H3DtBGQOeRTKgEPPAja5vSQlEIq1tvNX1LnXuZ5mJ/eq8PKVMAUFUIS
JGkLYqQMf3ApdZSF/6MqtmHvNpdQtXCHVD8cHpkGvxITA/RW0ux62jLluDTj2m9K
aqFpIhCiXoMKI4S2TFDUuiy2H1k9Qn+hoESTphwlUSwrU22m7XwttiXYj+f0CkcW
siTjSBGfxAmBvjexCTaxtcf+o6gr3giZ496723WizC2pkSkso0niW6v6Om8T+DdO
WJT8XSRk6JyoUTbDcnliXMdWObm1U+bHcUBTY2CibTTGBnxJ7TNcmU5LNzP/ltiM
LSSjs6ZOWrMxYTJkb9/HJuglLkAaFPrIONhvsj11eXY5yawJYHXJUXBZOb4fPylj
79dRzaUqDT2D4R6j2rXOWuPhlGCmDep60z7Ic13DfKAp/IWtNOWav2WxdrUdM2wo
yY004OjnjTSLC4fblSb6sFM/c+Uo+j0k8nkNfvoV+cNwpDWsBc21c4Ip958yU4fu
Gk7IerbEWkVooZJvg2LxUz4ftsLckqGb7yMALuCTYuPzr6Q9kv471n5AI+2XRvvl
o5ivXV32Pv3Pva9nfMpeCOJQZV9XKTKaihu4NiEZ6bp6S/7gqdXS+E00WoSYEEAR
m7kAvpP/ZaNDDBDs/m3HpoaKCV0UcWkXgczVd34J6NuwllBHUGZvWT8anXmkGphT
o1zF6amdugPGcmgqOwKWPeUXUg9ss9SwXM8j6xGYQR7vqzLi3PjzYO/N+2WjlhOl
f2YNecCZFUUmM3+/29666eio/EM+JxdpV1hxSiWI1xkOZcvG1Aj9OTB8a/C44Qp6
hawB0VYVHP3Uw8rp164eF6jQVvJ087rcs5VRshIGwz/pEkmVM3CfU3745ubm85gz
TfavkJy1LQnHCA1i3CEvxbNynZG2nEqkmvRmHzVEaowuJikqiaTvAcDLac4JER69
hLcWMmGwOkwfUdY0S3bGeqGiF8JhM7zKh9s6gZHYsRqNcJ+rcHnSG6as9JjwlK1U
TdNjFuWhy6x97Xmi5OM+x+pNr0p/fe+9MEANoB5Ssuki4MyvoU2o51LuB4KLfL54
yjhcMPaDr9lzAw5y5DdMr6VMj3qY09pzVQhBPpMgY8KErbkrmC6qIgAyqoYbb3E7
1gYZtWKc9f8w5a9HAO5eIhdW99ajWViaXjohhr/eoy0GbXbEp0rb1oSbOAEOj2ai
67zSgG1eI1UC67+MmRgQoNtHqq7XrcSoBLVpbgOngz3Q/I+kWOGo437xVPMegs2z
1c4EdYJZhxsJ1lz903bmZc8MWU1PzY5wrmqJaiyl2aLsw4X3AIGcn+furIdWQ5aA
PBxqErAKxmvgRlM5/oBPikulvBUKIqvSd8EMwetnjkC58XKTC9v2Ablkcc416LOJ
pJbSQmj0RtzwR3/ubRysjPNxkfJpAOCmbDzT9+GKn5bWUflIPC1tsKbuh42gzbOF
qwBxGwkoGrUJBOJQq5lAFUbeWcjXg/NbFkM1q3AgnDYduJY/V+jKgmuZnT+qhyUA
/zL0ygECczw3wMPevRSkAJxbk1fssEZiYAuPIfFB1Ncgqdnp/0EjkW0jLOo607h4
gXe+JTIJ/FE40/jsWvtwSqUDA0unGoIOEQDlxiQyMcCuIcQ89hDVQFPxKb30Gr51
FDTVYsU2Dp3X/6kTHQXjIFYlPrWoAib2HT+YyQbMw5nOlWivpnMMBWZ5ESlDg0MV
Um3D9ZxNM5ZFtNTYGNFfG4l2CbvXryKOApD2qAztuKzvonhfN8d4tboOreNA2msS
B21r2BR6FeysAAWRCX+cj71QSzj5UMpFFOnAe/ORhc81gRb0jiNfGpWagKgdpHt/
gInvYoymsxqQ1dqXa3kzr8c/7eHEi88ocoS3mz7t9MigZfRKhA/7Vysm18mJ5CDS
W9syixl71O/t55rXAeZY56w2XxN6fTgEREpwNN3PsjpNZVjL+sY8tYgdEqm13VUO
QTsmaNIpQdLQZ7yR1ofQ2mJy5U5VYiUgw61Y0r79wj+SVeVE9jHwm3hiXoHJ55CA
gQxflyjteqcbYMM1Y6UigwXg1wP0qlezrV1KHx+raqTnD1J0fE9A73XaL62M0DL8
y/lF2uCWZ6Hmd5HmezGZ/mMsL8BRK4Gq9eVoeXTKt0D0BupeXw0YwZdCIx3hJjEK
UWw7pPH1epd+QPOrla6Pky7jYpgJYYT8/lEk2b55GutFawM+tGTYgXBul8TRX6fR
AOVhE4A158T7kuveuGXZg3o25Yk40ojF1zmhfTv0DUNc8Ur92OBmb18sDR/L3xqA
GOFM/uBd3CydVv/68EDhjrjc8eTJI0mzJpLBxSL7RlodPehDSImLCrY/jkmvIHNp
/TNJ977m3cK8rlrtZAz2OrpQSiyhn6r966eqX5aNxUuRlK8mOlj/LxxwSgmh192u
SN7APnvmB2cQQUt2kcxnA+ABCvTrDmNoye+Fj+pnueZQYkwxKHyVmXT6CJxbZu4y
bkIZxyvDbNU2+pFamGDb9uw19fuTRE3J3rsn2VKQTeGMDYXdAe13T1vrFTmvyGge
T92F+qTwpKxxm6sf2wa3lg2WhuGJiLR67ptcYvntDGDcwET3B/Qrbbm9Gp6fSjFD
rvQYXLz60BghK/tc8fSEDLduuPKhAfzngAnM6GsyaCGPnwHPaHG9vPnz6N1QWhw0
oUUUjDsD0eJWKfz7Cwqn9jguuSOlzUuBqhzxPWBgVxTbN/fqUPvVU1m+66Vd6iJJ
Q3YSrSIQjKwpeWPP9h0Ybzwnh3oVeIrzEmBMFNE/8GnKqfpt63/nKa/QDkUs9X9M
+ZA/QfsKooxESecLQfMmRjkpqeKI7QxMMdFAawuGFTkky/jOYEKUd4xyc4/35sAE
+H79e/iJ/4D5BG3ueH5bMfBl2lnvNtCQ3v2+vfprBr9OJ6gFow9xla7eW8OiJp61
OlfY6sI5oy6F4nBGHux91ebojKJG7cIBF/XyXKKYuBZ8zDiZPoKUs8qPnDH5d4GS
j4zdiZw9anbL/BXlh/iEfUIejXb4wcLYepuxmXzwNyntz+Hfj5gv+2zthrP7aLu9
+gG+vWiPZHm3ugh04KMMhL0lrc6//u2r6OUp+NeY1f4NnWHB3U+dvHrji6mzBEQf
UvQaW7xoSrab7UW7YxQdOKhgeZUY/vrz4ZO6zeXS8OS0yXYnZqIph2vp1+I/tTJL
enKRk11O/1fOSyDi9jpSPamMBs/3tLowy5BOYp0OZrLA1/GanWfQ6BMkVG8t9iw2
skemmsRJFEtLX5OWTYa+Wsrzg3DcBBM0LkFI6x697EJ5299pPfAzLMkIrLC3FmiS
1ARABIA4GbWDKvpASCyJ+sgPdqy7eWResJkubdIiacgeFHNljRBd9LLGXZaf5GYa
6Xi6nctiYfxFkpwtd3xfX+sSbdpwQvVsv8Os9Fmt/vMwMlTCzkKRHs7PTAJg61IY
TlY5P3W2qm87KH09/qXLNgTEeKUcrUNW311W/2mOGa6rbnULTsihud+YavBBJEwy
6TQ0gy0W9TY0gM14a/QiLORRKwBaG7HiNaCwA71dg10zck7s1Y2vDabBL6YicXRk
wXlkKEerYUJt7QSlkRkgtOKz6CxopIkDU2lZoDrlrBHd6m1MD0V5obLj3p/NaNx7
VLB9e5ZQk/q7QBWuQbmqefYFmSr4Kd6n+qqMW4CmrHipeOnPT6BdYfYQFak2GtsO
vJRGFg2opwEMgvXkQP92GsSI7hNoT1x/aEkxWuTInDD2q7WTiVxfk2rQmgabT9e6
QiCYR7iTOdT+Ns58Ef28uqRmOarRY+d8+pEQknzHU7LoCQv4ThSm67gkiw4EN7nO
gGMiY3s5TTekvG9NeZ/XwRYyMbqE5Bno6FeRrtDqtpwMmpdpyp+f8+oSZs/S54SZ
trgY7VE5NZwhVI4xLwEpxC4ErB1xtW/1zOIY3KkRxSCVJtSINGGR9q/pt5R4AwJT
86hZVoJ5UQGy7LL4q5fddXdtgEWIWy2U2ve6SxgGzwR4GsDjV7HU6Xo+gV9areuA
`pragma protect end_protected
