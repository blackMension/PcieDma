`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EkSWAXjum6+fwr16SeK8StJxeTv0WlyHRUqtUmbyJdzsxwLyWK3F0lkmG+XQdSij
EsxlsjNl4VJLPArXlsF/wiJGPl8h20XCXX4SFJuFw9+ZlAAkbiv2NE9nl1b3pfkJ
00Vncy/gw6lws6ZY8M2H9P3+wpjUDTP/2meOlKCAaG0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70480)
GsK58UR2KoOiNjakUVCSmzQIvKwVUuo/K1wAL5nYGJxQiFYGSBpQ0D0HHBCudoPm
h8XC8b2tmAbXCI6JBW1ugt7zlKgwXM8Qcj4Ue/OKLEwmCZfjd5fp8BS0fjWJHaLV
abMSbruI7BqIzl+P9uw0nu+mU9E0pOrJep/bWbpSRypKD7AmN4DkWnrpXKlG4w7v
n0Yf0O1soDLmncbJw6pf4jWCUIRwoIWLDx7dfAZ/bmwXmUkKXOuurat8qiNK9vnu
hEVNoa43B8kkgwxRM4i2Cz9LNfaOQO6+yg5uxQLAwp6Fc25m3ylFh5QbgxbUdGYF
i+5EfgQK510GG7keuOqQAaSuDAdtVk3nPRf026MbAf/p0ErOYKTC0bq4dSYKL/DH
1BGA0fj5XjVww1wETbgtYSjeqGEztLG3xHauAGD2YUFqX1WuFqs8OoL0pZtL1uKz
RXS2Dk2mz528DaIvw9ETo+Cud02O5wkhQsPHvUpa7ZrnMaoc7/OpeqTGTngvFVJx
B3vhimfPM2sXRQbhjALMglxagwPdmzNzdBZULaDWmAzCqABDi8mmBGMDgQMxETj8
PT7GJ20/azbbTukH5UBaN7N00lDUbli2KCcDyTlgB+Mdrf7Dw9AIdhkJcS+yEvqt
+N8PApE3l8u8CYYSG/hB2zhU4ilGelEJXYRr122sZfHULuRnn6WZRALl1CErf7Ru
/Z2dbzZq10+zWhvB+0VXu8ipNqPiEMxGwDOe/gSkUFC82xDnAYWZycuB+LTJQvhh
us5ZiqLyKohXMxxDGR4Ub8IrEP/moS7qub+0earhmBkBi8PpksbbnOUKV1R8s/Zi
Ybn3c9zq50utsnF5KAiJcVPaUe3aLERkqEis2sS+N81Hv5Lji42X7/XztcOSFuhd
rlLjZ12IjuMY7Q/S9+SehOacZVLv+rvN66QKzX3IbOxB+lh8U9QZdkr1vs7+/avC
GC7zaTy+1wFv6h1slReGWKp0iYZm9FIKN4Bwije/tXOeGoTKvjKsrlArbFDDzxS6
AMhZbP3fB2X/RkxIRz0oXA/pDeNilIJzcSexy9YGZ6CzdTIj6Fw2FhcmrRJ28k/w
pmQ6ImrlR2r3dQficA4YN5gbzCdJYtP3FlrC0dNWz2HnMGvPzbdvj2IecAYOe++2
rq7FLTAmg0CGMAKC/E/rmwnl29CZyiCJwTKjylDx4ze8SEabhRNeHUSkje/2qHLC
2Ext6wmE1ZRIHpOu/nqAcO4r5LsHlM9GecCoESoRah8apmNX0NqeAWdor0CgKv4j
1/EpHqkd1TkvudzpThcekrThzg8TEgvHbj4lZPivkPuRFVZXgYQt5sh89hPEpkpp
RBu5fOsfQW9ta9MgWc8H7ziq7E46mBY1vnYMmDfpGTH1SIEnyA7R5xd2cKVhKM+7
+tcUGGGW9HZBUNAiZLtXh+fJ9CzWlbBkPp/akIDetdr4MwMyr2sNic16BJE57i5n
yO6iuiUP06AAku+ySL3dKIEtCO6HGRCb5qcOWJqf+/4Aj+rQQViDHTRclMGEko7N
B1opCm7kGzaWaFUlqzHF8ISVxqOfBy8nkGZl7Up3yQzn6dDzVU8UIvB2dKSLICpi
YwT9pGPVsOeQWBByHNzhc6dqC8n4GESzo/A+Yd6mfAgTb3ut4qDo+E9vVeaOnIVS
2/QKG/2x7pcn8IxZ98bKGZQxJKrPVePJmJ/NT+EXqmcyXq2Rwx3bePFHaeKJ4qSc
ORs6BzbAZAdoj2iMMmStCmOdIu3fEMqL4QiWnY/hMu45C+jUcmKq0pXRei///vfs
sLw6TpOjmLD/KlL3Jp5V7BcSlW+/pd5MU9TVDRUEZCIHkRv+Qky6cRlyr++8+QiM
X23g8+61iosZFd0O0+KeOrtHPhMDaH118iAUIlEdLKYtT5KQQ0qZWF7Dxou3IXPG
YnBhkAN8AvTJTPB6pOiu+iUNpNI4UVMjoKDM1U60xGd6BwQ2syIlvc4S439x/wFP
R8z4JoQNJFTPCymHzdzNiKPBJ6SQGtidKay8YEweaLt3VVIH3BBVagHwx/mMTgEO
6ch6r/yQfRs3wrvYjKKqdmRA5qgsYufjdZ75+Pd682BiUL4iioippiwt9GLq6hrn
8JaB+2Vl9nBzEtDIPyQY6ysBfWTf++z9Sl6n69VDoOumVE1OsXrfUy6xA5VyE5Yw
nWMtaYZA8VH5255QVocj6DHcg1vjFpEM8vahDsD3RniU+1utQTd6nrViiD1ErQR5
6GHyjKVzpiOQclk8+XyzuHtrWtm4+Qa/frBzjdMi/JIMekRldgf8a91SEdA3J7Oy
ur0tZCshENFwPMAy5tSZ4pNqAPQnsbc51AQsvN+OfEwEzDT0y+PQH9dIQGGY225C
/T68YyvN77O8QYdhjI9rWJAxKnuTJqeDRH8j22Hz3wDWtZ1k0ZbSf0xkFg3tr26l
jPwaWJyadBXtZrdWMPSkS39/9wtWh8t6UzorXtTXs5G20JOw8z59AM/UeA0xOj7W
WZDF+MmJZFVDt8xTxviXMD7OFQfh7Jvz+waZ2mD7n+skFYfxp8mgEqDXlsBnX0PN
1EQOI6j/9JyznfnL2hWkgmhZ2MxH4k1lbdzRIZUuGgacK1CAa6EeyrL2FX5WBAkL
3OWHl7NT+fKbYhAaSbw/sKuTEP5c76yjHrd8EzlStAJGaxmzFLGHm0ghu1k3sciZ
Exes3+0zotvthLaDZhLHRV7X8fFkb/B4G6UHFku3qaK6Aw6uQDx6+cjoj6yEIRiV
yvbVaX8iEHrWqf2k84ZyI/ZKZaTPOToyovXdk3wTSib/XRdlul9m5jLvLCmRfAVC
rPTiGd9GqfuzDVbbmBLLtboPUpBmL6ziUTO/4zgT1AzRGIzOt3z0Jfc3RLLsQOfS
Af4Rtt8foM9uRc28JUVjP3A2ekLACD2Jo9N8CD9Ff5/lS++KO8W1yyjfopNUQ6rx
/Gw3635ZE76ghSm0B6xTOOnCvrYB8orLt0v4wSWkGa2tozuRSmV38Fhn9kEEGFL0
G5yXFfcWfhnIFSrOkDGd/OS/CwuIzGQ7N+RnIo6h/1tc9rtihDZRIWMPdDeiOrfU
oj55+lZK3T7XCEp/lSnWAeZiM9TVw25SH1c8Ccofqo00+3SnVR0JqCjz13svJSn9
jCuM2dX4HVzt65FzhFmIqZdaSdsw9GCFwZNNrXkAme/KZw67NKapIEWm1bmezjnw
M4xwIKmJ88IbiwiRMhKFOEmIdCceMP0okkkjvJnXX6Zodzwfw+x85+qDcTjboen6
GR6ttI1kFQOutwRCMEExUIUJcdLtW4uxVLhHsFFaCbfVM/g8AlTAvsg2q5ladR1t
lvMo6NIlawoMQdhsfViiLfHfEjfO5bcJGWCdHG479AzqV59RXOmKXc/pnja90SMq
MoIv5462ab2iLQ4A2NiuS2DVbUTDMJot/XXzc2b3LmO6OMs7MZDGJTzICdeqIDIu
BNa06ifSJdYkTidqKAzDfJbl8ozaLOVXWEoox+ZlOyif7/a3wTf/FHDkYpAYfDlh
G5tqxCsJiqqkReLuXk+5n8nUJoTxPvLHzbfVpTltDsLXjN5bDiyGlW8YlUQahXwM
hb92ciIqv7vQKtxlRMbwCofeQQxoIV8/1XJjOzM3AjiYgwCvoqNqHjJ4brVOr7Ut
A8PAVIZR8tL21hDITptTnvTrb6V/rZfNc/41gMM0a9yp25rY3cdcHFZJKqKVgMjX
/hUJrYhN+sFkMtm229a/NT1UJzY4oY7riYGPA3RcFcKeMFUEQSvbUeBTGnk6gkDY
s4wfyyvoLLgz3sjZk9vpCGV0OUg26/uanD7gYf6KL7QStEvzjkwoQfzfxsIqBw9J
pL2L/dCeimnRhMpAaGGGCeSHeQuvSuJRbQFGqW/Cio03HTErODjJsQa5zcjco3gG
AO4UYItyUWTyKwyGJMJrAr2m5KZ5uCiqU4WT3nKMhwvSiBaqEtkgxalmVdEX2CQ8
62bvaa8M+f16+Sr311+0BHP8lCz1WPigJUREhVLAdmxvs/GYuci5JgTs1mxSnkT8
ZroDUPI+kG3/dROdqCMXSB5Id9MA5S1C7eBWBxgZoeTkLDtyss34u/NDRK9XpOHY
boR8ZJYZxne2pV/47b/3eqzieI/IPZJEMtS9Lkc/dch3/5fJHbAhW4OGuvCnl45q
auaIjmPE+/9yJoG3wuFJo8fyJiwx50fghFjUCcijLdr+Zm7ZhotkexChrBW4eDOc
F9Vk4DQsaaFH1LlJtLqe2JcoyuxVnBM/DGm6JpebvXw3fZBUuwBLm16f96Q7Weq0
BNCkdDtor27JsbIPdgnqX9mdb40PqCZGlSqqUvWuPmk4/W1ewhKOojsVlipPl33D
M9E8JRGPjDUuasLXPtm5I8wf0WoxH2+0KCT51pN1n2/lIgN5Mik5JYSLemuCgWKM
U+Hr1eoCuP4wFqvfHeF9Uns3t32TmkoWRw7xcpgCd9sF06lkI/PEboEbnXdqDF8z
L9NbY0T1HDMnlFRmHdrT7zxRXITl0XCa3MQCbxT8Idu7B6ioRZ0wqg8cUgOwyVks
PBGhT6D5u+pwIvlgJJfwO3XPQ62Qa1XZPbL0EtcX83nstST1HZqOcqunrhbWCr6i
sttx6WKptCTIhl34/DjnWUuZU5b7kU5DpPmyZENAGJb7v/GJ4XlZD7Ra3ZhSbKX+
hdSbYDyIdkQaAZXEpstVMM+q2lmBLzrB8q1MKc0LOHufYTqczSwcQCCObC8hwKHK
kH+Exm0h3E8cAQv9mwo7MOEYkjc21zk3TrSK7cooJ8UCfi7RiSnFU0AVjhtWe+zW
8txjSIl5Sq/5WHVktPqfFLmxf2ED3ZWnRrjLZETC2ZByR459Eu+HQE4MZ4ISRADA
BsfVh7iHcP58nXXrHeEn/1T/03DxbwZWlbaC02TuyUfv6u4/0b0vh215Cr49odxl
qTGMtLkPOAZ3GCI+TvgGKe787PN086J1fKA5TBsbymvfLn5mhvb1BFTGt6r5bEcX
zpX6YhezN1mn/NS7I0wZw0eXXP84sD0VByJ4XQ8zwBn0feAs5vu+j9XsEci/kuFP
0DyMOItJzWJ7Eotaa+Hlxqh4rXXVU/LXZG3XoElavFKpM/59TW0WwhooVDiJ5jhd
rfODDuxBna4PkLwviFuHOr07Qxpr/vZqTlLdySHLbdie/mEKxdIkndeDXoWOXXLV
U44E6ambsj5HbqAK8O1wjrCrvfTewB+rMA7/7kQHsfrFS7Yolj+RFeYoyqxlFgWc
LabNJy8xZ4bxHZW/kgUd3So+rp8DRYOHe0351uZ9a6hA3VYWI3rbErjFMddigHtO
zim8gjn8a6A7FiJzhIO+BACk0vWM5EwBmLKB08Tv+D/+QJ4xiDjQuaFoTEwDgM05
V/v8Ywr96qO2RSdtViqR8zp/nz/Q8hs/WdG9NvReeLSC57fNwZmldqIFuMhc6SRO
AHJQRAKzQtYhlHdvd6XhSph1ipORXnAVFHb8VSvdoQEI70/xxHQVe3WNIdZ2wEC2
2Qp7543RbVfCB9ovEWUpfVDSOzPYPUPgzcFdQLKC7tLkYcbOEBWWBiCaZSLvJC6i
JOAD0aLOcPEd5SUzjN2E9A6HCmuIi+B3/yitd+LJxZhrZB5GMiSW78P6YBbLo5tG
uhoITWhcJXQXAQLxTMY/lzbkGY0b8DVd4r1UMEM1VMk9u7K44Kt/pLz8WCR3nLGK
Z6rPAuKGSPFnDZEqRtUsLJIuNLGAFzzpUDaNWpDpaDwCPhrHMiEcjz3FLtzSZyiw
x6gS+EPCcxTvqhcDbaGkDsAIokt7WySoL9cUO1nIUXlla5YlNNf0/kKfpNOn7wUE
J3vW628+aiUMks0yPRItkkx52zJh8K3AANadqUfwsxxJxGChLXSb8zktL0VWkicT
UbuEQadD0vb3QAvC/TKhHrX2rOMzQ7I285uXRPz6+EZTu4cFtD7QzuTSwPhdEEUg
0DTss8qTQ1LdHRyxvuILQD0A+wYofCvSDaRAThLl6DpqF8uVrPwv+3bxcZvD1Hm3
n+0Ewn/yvNY5UpsQiM+kilAjJrNF6c3RG3BNdlQhTi3I8looToqQXFSapj3yLKEl
3BmLKe6IGjlnIq3uETX9vYgVqf/gABxzQoFcLSHwtQkPUCevGoHzAG+2gYV+vnfa
5AuttlGNNSJ2OQ/rztWLyOlzY2G60JGuQMUhQc68EAfxyVXvQOIRLxQl5lVR96oE
QVN9tFTPfRkBCYMr4UoSqGNmOUlrXEPrjsiuisYoID8vKRhsvThc14hSJZd8ODQN
XkPeEILzyk3qwzhexdO7/4zwdTAH7XG73gQQKvMyDQwUAe3B5ba+HeQV/6Hb7gHM
vV/mpI1Ua6oUucLsvD2LvuBxtpkqdXL29ayoILEpYm1G8SR+JTAgZ9izIvF6l/Db
8r8Psfd0YjRgWJVJuj+1uKoYZyy8b/aJNubayBcPheFpA7/oEqeKbmUdrVk4PWBz
hTzwUF1gl5w9cjK80U7yLssZqgGWrdBUJajtJSAfgszW5KY99+ZX89Hn0aqMp5P5
JdwU94SqxgRpBA8Mq1y4TzQBRI95XgessL3T8ec6AFtwllaIjFF3IsRjcbBfLvPX
DrBKzzFbSd+byeL8ufT1EafULez4t3X3knc3hLJs5f8I2mUioGOfwEFIAsecpyGp
HpGwYBn4+EuEA3Onh4xIdUdfx+k8vREQXtJ+qWHETc9MHa4j571E+jjKcXSP51ua
9XQpGy8NugbOqoVfsIDUvIpT+FEIGYok12Kcz6rHnw0KygWRJl+jxlLRjOaaSkqK
EPQqQ46kfPqITJ6DP5stbDw46fegRPPBkCx29jVqZA/vT+R0zy27AFacgkodp8mN
e4SuhNBtFi/rNSs6tzFu/0CwB6sm2aKGlK6W2rbs5fkfC1JkgNSAR6hrZndkUdHh
z2waphH+UBPaI7afNv5PtS3nPP0jrSZFqTWGWmoapTpEgA7OnEviRNGHnQNRQRMf
oIJ61GfPdn5k8HQONsOAyUWNmkFQ2KJpfqiaWav2OVs3LBdE7XaHBidUPxs9fkuK
FZmHSjv096+DgOzR1trT3Ls0wRPSaN590f7ZECFHfktIxFTuiYXCvg4y/Ol55oVP
lK/xjrNI4NDVFjSsS2Nc0oQjrjqSCiYtVSnJ47rjdb1axOU/br8C50rKRofEPbvR
ocDUy8707vIRSabOy+7RhMJXgvoQIX0XGwFlF+gv2SO9wnF5KlOrPZF621XEiJ6M
dlu5JcZoAV25w3XxqX9bclr+2Sx39eMDM/uA5Jf3M5s7sNNqvRqs5xQ9lmYIK4hW
1cdV2dAD9OK3Gm6qDyGkR2cV1aP3AJJlI7pXpPMQcrlToRaPY1/zUyv/rXxJG4xN
iSVzolsFyitC61uZBx17My6hN/YtJRUiE86iTyk7IY1vvUQPwH4OMmMZ5FJFxvTX
KTK/5H19mwdDympgdz8QgUBruFn1CUWTtnCS7CRH/CaL5u2ttgnNwhYTGRZP7Ja8
HYDJHlTEWVmfLKyrEq0inAlc0qKBtieZtIJxtFs935TsOlGDrtSf6OGk0zgkDSB1
wYuw85CXyBnUDftL2j2k7RBy0ghmpmbSVCZ3+HcaGPJo9Lfm74uqPjTzUmrTzWN9
imCjJwGQ+dGpCkm4iw0tWT18VZxH4wUwRL02lWjP7eAIpljfvo32IFurpaQ6s86O
YNB3KHIml2rwvVY8RrKOvXmnxfjWdIuKwEtKPz2jG1Kd3TkphC6osZ0Z1X2THqbw
k6Z02ZM7z2MtzQ/ybldLJonWwuScTXfc7xB69zvYpZRkiCc7vuXbIjLF+TwL602Y
C3aNvv6fjrPyIar/Xn9xVCc4rGCIxc0qFtMZE4cNbrbd6Ta/zhvbshsO1goWeYOJ
jbGGeVqJy21R0gt7QPCNL6006unZPkdfS41VmkqW2jJHEKMVTGavNmuNovXve7iK
nADadOow3qSOHdwOTRCvpqHUe+VRW25XHAY8uOU3pcDdhLcDkv+xs54nLhhQ8yFx
gDD3S5oA/xSziByN5kTK4DJeVfhD0ksw1/aDUdtVqmP8oN+E5CT4RXLTbJtfubM+
JRd+ueqTvKzQKUo2TI5nj+fGV+NAieYqgP5WuTz0Hbbn66KMf9BgPjIBfgCpzztZ
CNyBnKiSpjMXui5VOvwF+fet8xNajpa9qnjM+2nLjrZ+s9PB4a66EKBV1B3w6Is7
9617RgE8INjSxhgPP2mh+UUQguLloDuxMBIHQb1L9y1WGXONRGX5BYdbnGl2EOUJ
BrKBdPXaXGUydZNRdB1KibrIuvGcr9OWuIxVOz4/7wWbNTkjeoG3oe7kBLrzZCNU
B3jj+B9RSKSPqM8YpHoH08nUPrsm/pviMtVbV7cki8+TB7N8VzrGr6JikkXiOY+D
gTCr82CDla0G2xmhGoA77+m9F627tUEJhM3Msi2pfAVtFwAwlUj1ETHQXokNIlYm
GJESL8UbaXgGAagDsAmOr3aghoF4CG7rcQI/DNBigZ2VDZfxhVOTOQ6qum/r7UAC
MpBaIyoGth51TdQSUXqighXmtBW/HsWL9bCBf+8BqUOm+B+idH6rcS8a8qUr7mZS
E7zeEQT/qO9CapkrI9GqVZ7mjWCKXQQYAsyxPe0Auo9MxRLaDDtWS7wxjvxMhPbc
RMmtsgfl3jyOvqRU3/FOUc5v0jCuaDyLum+eLzF5Zov3t0FgbGTjy8peDQcHEQSd
GvDXSmrjsVRJDKF2xwEKHWRP1eE5OVDZV5VZD/W+poX0IBhbKRf5jQeB/L5ynD08
TWQojNsfPNP+a2ATAZbP8MNecVs2qTqveL6aZ376c9F+7SB/9SG3QtTANKAUkdVf
IBgzfNBHpjJ69gxJQ7t42FXZHim/ALTiaiSeALSoTMFfJOIQIntmPHvHr9EW8ooQ
MsWnI5qnTSbHBmqOcabLUwy+/Pk1MUL2sHCk4s9DhhogcEgXmcLrOXOuoKI+t9Mv
gv4xTgYN5dVOVKngcpojgqht7feiHZZuJUcPkjRU+UioglmcXZGkiPXw1Jde3nBH
H9veMlyRsnaEZHLZyrnwsuRL128bolLxxfeeZiDh5CbDBL1jk471Is2+pHgbV9oU
gQm86lpLLs8ZQVaaDhnujKwSLwNW4g1XO6z3NB+UBqQEt79M3I/eGXCmy2Tuqdoq
e/ajLVcGVqhUhOihlpNOB1jqcAAFpafIx3+tzQ+K4ewrQ36OBigvEnJHC9DR6qg+
Jdd6PLrALTRv4iGhJmTgGDjeIBA1svmeLN8nVB3zYCTOUVHh7I90UQ2AeLBs5UWf
DKV7qkqSf48Ik0DlNEMBsbAkE65V0MOBxadq4N7sLE8IutF9zHpCRyywhRvNO75+
Ls2hHf1O5Eu2l/Ca6O30KwcpWvThJdXALzjP/H9k2oloVQWfzD0de8drEYB4R2eO
gBTWO/U6STcoSRQyLnQ75Gp3YveFv1aM1iFLTmcjuS26bLpC6VCgFacDSou0iyZb
iyaVmADIqOrzaaQyGR+8/zaWoNc0GQA0H3eYpZKIUbHvfbjAYkfUeR0CeDUrBFp0
JUc5H7iOYMGP74L2CKIOHTlTLXXtLPVRViBL9E4H3UKvOH2Q28zsltICeDycZiIV
0zrsEXM4UD6MvoHB+RpUB71r/CygYrAxyUSvFO0jLpmbahSzzcr7DyEFHbA1prr5
8Xaow9TtS2Oh24fZN6tc6Th/GvuAUZBW9O2AYQO0MHhJKguai8m0zqBbfqPWy993
F2Znd7QWOy28SHPmpNO0HmZ+cBbXGU3mYMk0CZzp+cU2HES0vcDOcEyWxjGrvKZT
poA4u2T7c7p6dAdYVds3HmZbphvCXMztdnZbxyeD5lgyeYK+N9mKcRPEz/Zq6AcL
vjiiWJMcxhU3k1L+w7lY4p9oIj23KFbyFDvtrORnitkpbYOknPgKY9EgaqeCKMFI
kwvUOrnxqWacP82rveVPUG+GcpsTICId2k+h2Xdn9Ro9MmKDvrSsrXHnfkEMxddx
VWxvNFekzagqeyfTw7abKptn8sLrlxj+0r3tiABGRXQzq+9h+f4rTDeqNNjh5/1d
3LFcZ1GGMdPrlYkhvlPAzwoI6uAxL41UX2ZHKKnKKw+9CvHQkme8880C8EU3GI0D
nMVhIPyJHz8CwXRjKuyQXPoTCmkCyvnj7+7EC0cQd61R7iQy391qMId8cV1H3XRE
7bRgTwzH5WbpJbmMng0kIGF3C3f4i3ipZD3/quRwAbPJA3uMZUMXLkQF+CCQgaaN
KseBxBHGqnmsX5yiXJ/zfjjxJV+ZCMnAGKsZcIt5Jj3FiLb+mwplJMf/SSx9D1oe
bdnkHB+f8mmhgKWewnH8hoHQ/DUX9Wun4ppHwxDdqRgEPrtUhLb6lt/6btrQYKGQ
91XTH8TFJDrIjR7nyNdMByyNdOEsVUsVSq8+IT2g7IuUbNDJmHBwwvt1RIMp6DxF
UWBuuXK/gHU+jGEW6Q+9gHe+Kk+KvtVnxW7cksLOY0d2wl3wnCO6t9Cix60TF99r
CEzewIEFGEJkbsPWuNT2F352L50RQJVFS4D9m2dfugxI9v9T/IbhHWZIVvem+3c9
V39dILXA10QfV4mNyx0UNefIY9oyg91dNXrpUSG2bHx1Gwe2Uy4PlnackjQ++nHE
4evkEbrSDuSddivfjhzpFGpsur6ANKLT2865SQFGYBT/doIggfKcxXNnYohw9hIL
agqwH6PnYg3e2mYnk9++e++FVrDVX2vUr1WJNQ3bOrDTlqnwve10qaVoU3hi+aNm
eSaw7oAax9oX6srI88kgBku7wmJGGWfOlEG6gGYVu4EGNWip1CtZkMUDRqhJeLyN
Etz4G5OGYVb2IRwQNGDg2Bvwom/GZdR6FqvT9P+rQBM6sa3S5Y5aRNGdH1jh6aNj
QHM6ynSFcFDRr91UEIk20BU1JG+Av7AbLf2UxyR3TkzG9btXJC101gj1F9/WheqB
+ngaUErMcJNIPBBbZz45iM8v/Qs2s3n3Lec1ilxedk8xVqBXTWNMiQylDh7kuHXu
+BCMQs4f5lLsBNQIvr5GM0vH0NgSg1rnEqmRq/jti4lhqzVuz2/hCP5YqUAt0N+9
vp2Ah5gtKraq0yLv4KgMFCFt9z7yQJmYW7vU0Y/arVEadb/k0BS5Fnz5OTjtdd9K
7wdypi/+SssnIzq5Qe357OJ0hS9IF3UYlUp5FNUzRlVs1ZtpGMWXWqIUwKvln6Qj
anBl01Gs6UccSeAghJv5qiXGXmFz3NRdfvaxztvWAITChQ3pN8keP0eV40CGrPsk
LZKyjhzTiOrMsbZf3LDJ1bA87QonpJpELbiezE/rKqI81aDqntzxj/nsNk5Hrtsv
neEFVaCuL59WsSd1z7ucun1m/AoeBeZMrde3pWvZUanhQ6LAUV5zgMpX+ixN0W+/
rcNXnWi4V/RMsi30ueVzHIoxZ2D6CrsK8Bnsr+iR2eF5aLEPTTK22SWKQUfAaBPf
xPmQRZFXwP+w+TJUJ6ONngmyCBpvKXXHKziIL+GyL4C5d9TVN7n9lEjR8ECcmAo0
o/oJeToPVmTp4dY7PRhEti1SornLZ0E5x0I5AYmoeF3a3xbAhZV4nUF4TcxbjuM4
3Cawi/Ee9PTPnHRt/XVnaJAkezKvaSfEy5HMuihp7oMLGBTCblYoh5DqYy8QUlAk
9f4GHf1mgGCc3K+7QxiB70FRqC3GeLU0zd5KYd/HVBZp+OY2pIsHsLXnBphvulPq
2Newbm+cC5VXfkDWw1J/FFKImUF4czW4eRVS8I1r26PvTZChJz6eZtN0JsNLN63U
/vhA8mIN3B66sOHjlrao++6hQaIgRdGTqpKcTVv8ajICEJoiWNmrV27sgUCez0YM
a54cWNFFiuodsERCEBNuri8/MR5RgEkBVwcXjd2PAnbaBGMU2UESOUMLkLZAUBVZ
Bi9ajf1Ofs20QIq113CBk7299GTHZ2Kc04vhbNncACjJF/rE510RxuS9OAOZfq9J
8dDn0M9o9HRO+OFpJGXvYK0NZtgk1WdqQ7lx4JKT6+0OBLs6hKsGcJMSx1XtdJD/
0VXh5AoeEnnFa25dDTwMv6+E6ANxYmw0WOOGAdsFnK39bXbma3CmarmYyv9ih87j
FWbu2XKkmnJ7in0FQECxa4ASMapp6vgfBawbLrkuK2fEywqxl6IfQpoFP3drKkmE
jIwMG+srJfULGyszNQIuzrFgXavpQyY/pybae8g7EsohAlAeI0dk9Lz71d0PLAmt
rMsr9xCDGokkdeA8021MH8wUsxz5m61a98NZr5TsnehZIdac/OKs/yikiY7VosBp
2Fnh0UOuS8gqbHXMyGO+jLAPUwXnnsOcrUoHOYng7OKuCfwtO2EQbWOLRvVCj3sG
l4IvlKIr3mFAd2v3CFVm89W1gE70oamO5V7kBEOUWk+m2v1bIYeKszvZW6q3g1lO
yiM2J+PQ7EkRNPPHhZ673eMwls76wECnwCuq0TtQ0c8T7te4//JZpcvJL4PrOpRc
5HjyV3/s7ZqFtjIGO5p2q0rL7ZKxI9EiAJmlpNCq9QGo2DWkaXtzgw/OdtVyijCf
0bF1KfOyn0wY+tAjNrYZejOo/LGI4LtQgCkactd8tVP43bgrfgm2iigFzIv90fyI
+YIdwtm7lMhFBZKn84UJX4/9KGcNhs4TeHNTeZMgU2WE0giyEZvcRQeiSVjxsnjz
ZDmVAIqYX/SCkiFMJFAiSo5Ks2nHbcxF7RW6so682UrAHz9cKrwqU9MDg3qLAnZ5
tCviowzYraJPcsRIONSg5EFXUWkr7JEA0Fu7OE6dWleX0oLKRR6kXimC9oGH8ws1
jQbGuQDxB+fQB3FblgQSRV3/BAhGlXLEtfDOm3OY+PlhZxWQnjsIlsMEgLcFXxp5
ljcctMZQRlhLC/8qfNV3yk+qp4nOb7IABPIq6LShvGLNJQbGgdUIkCI6YwW44c9A
4nR5AaPLhS64ZoJZdMIkfKnoCtjIKJWoTAHfc57UfEwf9uzsysGS6YufZZ6W8SuY
/O4CEKGZvop/W3x9pbcnFjKv/r4VRmc58//n+ZRSSygRVpzOLuB8qWSR10++1BAS
tBe8GnsOZL9B5ekrjz1RYbV7x0v3lroaxcFeCJiNCfa10wwgkdkGmzmbVaZIDvcf
RQefTWABLm3hzReZbC5kEkY1m3LJprUtKam6rkwd3YSU4mYs/Bcfln7sFnv6yt9E
UenHUniQ/EnwiWAppzcf+9AQkXb3ATbtecmuzoca0EG5y4IEE8PEPwwVE9ppmEQi
hrNiH4qxlyZpP8OcAV4ZZscQA3uHNsnj+OTRNat+JhmUczCG6+yeaxfwsemnOVqP
X/Cv7/6m+boLp0cmNKOYyWCiDjNKepHcW6ShoSu7mx4TwMk6ODl5yBBIEi3HI9Sk
7ocrgNdbf8RUw5aGXIhfvSAB4T/P4njZhg0nklPWgEoQdvoJSzdkbFgLak6ZoR/7
+tGfTeK4oKEI5oDdPA4XhqHGcqLrh5U3wETJ+XgPxjobi6vzqRFrSLndzBomLdHi
Ux9Fb6fS3YaixCrmRaMzQrCC0yrT1AyoWWdQhgcIRKFJJZ0G0SAxiW+uDrcuG0pT
ZHumGFsEq3vNe/5JEBqgfpyte2EoqUTiHZmZahokwzKzvjWEpLbffVt/gvMXM55s
8hcaT7UZJ0rBknJaYqsF+T206T1/Zrve9ffDnaAX99iolJMJ+d2z/aOdptCrA3OC
L9tebMHUbvqCv7PL6uQsL33pzxBHyyGJASamtwj/10jFxfHuDXn/FNn2sDzsq1OH
8n5clcWuoXY5lmfQZuCk0sIr/UEZaZ6FDof/WgjHUgcRk5khFJOkqZYwoxtKTZjY
Wbzbwd3VF0gppIqQDKG0H8ocgqTLq/KjZAKi0C4mwoloRwUM4nHAnBz2orZFLBOy
MZgiKqTCfmuV5TvC2SiqS5p9nolV2dJgIOX1QiFZJJOUwMVUaVHCa2KZBJlbbzmg
sztum6hbic5yM4PebaOsMFAaFnU71M2ecM9DMmPC01iVfSGMyY8tUcFExVEbNMHd
N5QxGgPQKqX79Xk5v8lJ4Ugu1onVGA0fS5VhD+Swa0IXkDTiPBB6ILY+xVrWjPiF
KkckA/ECK60yTn+cED8Gi6qcNS64W2CeBVtKEnaZhZ6nXiNS5LF4uGa0L7Xw/Eud
fubspeNEZtJQeWDMLkhOiu/BhwEFGjxv0u2DWdi7FySHCdrM5MBF1DyJvDWbiQLQ
hfTfH9Frfmrxm10T6kltdpPeJQHMb7KZHud0pNq5r1F+YasBVPlLk/lQUS8xc5sR
sfNlITB3vkRBzqHKayJ41o1KvkqiyfODzahCCdLWSFyMzYT7Jn3wr50mulSIuUfD
QoHZxRiWpcOVYQYaFwxVftO45GSNpiVkVxsfkR1VHkVE0r0ZmBcysVsrxk/h5XVF
LHUsVUpf9rFM8VNhSyzrHq9Ae03pkc+Ti9h2c/kidTwbSve6PE1sLMrQR0wZXJcy
xttPcficNhJphGDUn0gIhceAn8AU7rjWdj+qWa5arwuueHtUmJp55RLpuhaZwKye
x11SyneM8vOcL+YFVvlWkxoNIJA+xfVE3WPsX4fDcxlAG5lr2HlGHsk3NiTwFzXD
GiUj0T7b93bUrGUxhF7a5rUwRKVvU/j71YxbH3vmU2A61htWnWeo0bq/CCFnigab
ss5vErxqLq+35VT50m5iYXjU8nZVPH/6CMJneiGMBKL9VpN00R0QvH4UFD3C+EVT
XeQAYzKlBszPaGzjsn0ZHOTk48i30G+KiwdGoLNSgPr4Mu0F4teLgeH39GK6rlfN
2UmeRwL2G299ha2Q83KL6UQJsjpzaaFEFQrI5fMf9u5CF9dGjLyg5M9FCXWXdsbK
zPhbFIc8UrqqBxk/BJKv1elvsPOs0hFjIKqPbtkMLu6n7+0+JWmcvTiZ1IxRg1yW
bZsnpYzvXM4RUNCnGPtG0gKn+3mwGLuQPYeCAtNhGPO0guDd7aoGhqCUXj5n8Rmv
d8MMpu2jfjPdYqj/In6VzwBY3qZApeoRPe3tubyljtpNAwTFj6aRWc2yWj6YOtse
6LpW8AFBkNTEU+H6pq9Nc4Ywjx64+RMnQuqzrR3WqZvEuY0dMYLHdUdVJoxNVlwI
nKRn3yDRbRs8y/Tubwg6Xq/mJi5m+7WgGqLEQjt9gk+qtsRZm4CoKyPH3EB/SpdY
+BD3VDCPR/vZyNHUtwd3puxylPOsofhM7/4VJxsMi4NBEtYPPdiz+UkxDyUm6u4C
efrgOffp6JI9Z0TJHm/bilRUeG/xD7+KO+4Ky6zUOAW1pFRAf3bNNXpGSwP6O5sT
4jMWpzcaLwoBiqNhh3eURsqe16Te2Jd1+KcTnFqrqGgPnHg1nN8y45BhdYf0yUvZ
3T0u8fozL0jbedqFsrLPciIY0699xGeDach72PXUquxGIKi1KElmRZBzNt9a18pt
u9IIlNGAFYXUOPl6G65BgDW70Yx4YH24g8GfjrCkVgms62kQNdD2PGbAewQm2uGy
E6KU/FH2DFagVnXCQ0KDX0SE7XgJsRai9G7mMIl8IP5svwuurgXvlpR2SFNBo36r
CcsKtI87FVkczpMW50TGBGbCQDrO2sBVzKTU9Ms3NeuC+rplW3W/zeH3gVYuNAJ+
dpmNeR/gkZK/+hPe+g4SmLH4EwEolY4As/UyJ1ka4GBxFYL4Bd/ztUSmbnvCrTvF
V4qLBXaVOs6FqZlJ6H7ARZTkE9aZxfiHTT+z+7PWt/IWfV2gOjyrN3xLQGA4/lmB
XaD/ZPDPSJ1WcLyuTXxOe6aeyzY+rE4JBsPnRYeltsvuZ7anJDpUA8+Zp74sdqoN
ZPnbFu6s9JzzxB0cxjuH9xoSKGQmWpweYCeFVBJd5U3LSfqyJWIk3G4z4dRW96Hn
DaqambfpXd0/BnvwW5/T7d4dGDPUSnyZOA8syC8n0n58MCdZ6JIZRKua/OFJjkvw
PyzRwabkqhqKL6og5FbBlRR8E/guRotvpDzO0mxXQcjSU6+J9E1OvrY69cz8XqWa
zarvKkwj97WWVrBkIFHQ4trhUCeFl6QQt/7twTNX9LKdN4uaDeh05VYtCIyLZ6AZ
WqSgPlhY9eKs0EHCocxK/HJE+tnBf436f43g6kTpXrkzo+ypcltYcymzS0SZ/k/T
EVDiOAxg6J1VO3vSoLv996ynhgMpw9pMVJLtWL8I9dchDpg8eQr5yfKh6vd5r9iJ
qwl6Ya/W20aZ3SfgRJ6DcvaxaUCUlcvK3KUAHvZNSCagnuoHcrNMVFICtesreheg
9M/juyRnekbFErfHBYRgdJO3sEYndZhtrNxxWqcHwxM5TNU3ZX7pjUJ6C55sapQ0
MdyAP2erzIB0GL0dRktSEb8vXURCCFdZeExXNu0cocuio6PWUe2HLNWXb+gYZqbo
m5vOwWS7dWwSlM7CwElg2s0SYkzcKQS0xVN49of6DtJlBgWJxaTZkLz9VGa+PWxU
AYecy5GHC28TqFfAJspBU2tdjVQzPqSwz9wVF+qWKgqyo9ts0GKB/RHPQxzAQReY
kZdvxHgJ4XG4LHko5Cn/LSpw2LFkm99Lo0YEFqNc3Qy+BkvcShIc/SldKjkiT7fa
SjCQabPbg/oWCgVZmGtF8I9HIfzTFAFbILdIW979dUE1pj8+27pMW2wnkSS9Nr4/
jqMUz9VyfaTFGr49kfu4ijjrzU7gDmT5Ijut1kxKuEnH3F+Mxd5abaalPhn7sXjP
v9zUuLSsD4EgPcRKyW9udZX1hHusb7eIXWa+xBwtXamOuWbeRrDXY4yjThmX9avR
A4wjt4DXEAaHuEuCKxmQFYuNazNqFFQv2cBm6zgb3e+dicVjoL3ZZDdg8CI2mqkC
VR45low/o3Vn74iG6WvJAxg1opV9ePfgsZovl4NmOi9EvDkglDuOUN7d9Lflfq1+
PH1cf6wxvDb+fWN62/pOG2UyYrT+Nowf2Ukd3DgPZqtlSssxxvbkcRQX0E6B0a43
BGdLWgMNLFt5gGk8TS9PDQnD4VRAR+LApbdtCphXgP4CeECe/sevpQBsn1kjsPu5
/ur1nNyhTZBD6fl/XizsrKDB81TxDdwWv9eRp6ArYKUfMa0S5NMoIZUH9MYP8bcj
i5TTiMCI19aenq2PVAAuGUbDp/9+qFj/EEkerYsh1z/8/K+c9hO4cUVwMUyyHC91
Z2vO+JWQSKSFIbW7G8R0iEmaSgNpqvzPFjjoKBTFjjHkyxo305ODj/yTkYo23eeY
nyDMjj+BOcR6bMBkapvbNAAAJGR48r7TLcCwW1XOzho8gVvFv0vuHKadbTIQ7roi
hMA1pEZndQs5GgY/yi2b+wQzY429FPDYXsc6vR1IXp1iDZS/Shqt6LWCD8yJWub7
WISMHI+zgfUjPOPeKfjW/H7P0lPJGUCFXvnr2KM2cdMDIizCcnj63vq9A4YXvGBR
y+UGzh75VkWGLQfBlAW1sOqu8YTmWTe+Vqj7otH2aqI0kXy8eqZ0PjNjut5gLys7
A7v1/ER3etu/qOfT9L+ovjnmCAWuuIoPz3ITGvcNGZHmA4qadklImyY0tPvIi7MD
uNqn/qUB3GO1mHOXVLM3lk5Th/Gr6FzKfVTWxxwBhMlvUikiXp8TWW6ChbPmtTe9
R6bJi2h/iSiPsIOkmvVfuzXj91f/nYSIHl364dNAveX1qXZOtocRQyY202BrBNFO
dGnNfeRms6nuAGKH0TVWw4HvqerSeoIC3CSvRvYGml/Bzn9rdrIRpwj/ufLwYycP
e6Dzg1rsXeVFpZ9+DT/5myyDPUjhJNbO/3O2ZdUSJ4FFCO8iZp8nObn3HgFkS4Xz
Jz/gtFK4oAjhjQ8DpjQE+BEuq1GN3WItMBe0WkXjPQ8YmkzncxCuNl3FlQbWtDtA
YViZ4uwyyZQBa5i5R0gZgdHPCfmPOeBwfg7jzDaPnWAZIPiJFkCdrYIOXLy06zu5
R10uLVckuqbT9bWToPY515IeO1iUhrnA3qJfC/AK+TUhstgLSqyELIAu/5H80fif
KCEd7YgzMMD0iitlH2R1e0pjgTp/FDTjt/Iu6JibDpcNR9iL1zhK+x2dmxQSVliC
iONBDEmhkk1hWhl8OL2xyFGicB8obkm3GMqhxDIwsiVevW+1eU+iIsKnJCeXd8Oz
bmUECi8RqQooccYEjdsJRVsLnEJh50Us34zmULQXYiQa5yLaKQDwPMJcdUVf9+G4
if3Gzf5UY3Mgp8C8G3jvfghyllb+/PELX7f/kosD6WBtezKObV3PcCR8FtIsNiwp
WAZySwXjZ5/PpFk4jyJv04L19c33Y68nDYHxuE5SLI715SEau3XdUutNO1PqTXRA
mosq6l5QxP4w+1OeVEHN4IZLmBKf7jn/1ua738YBHVxQR1x1YUPM0laLDnwh7rqD
nHQB3SYAU3egfw71oDXTvk5sLqWRVdOqFuSieumx4FXZz59wNWmQ4T288FQCxaur
JaUb57VAAxLxGLYwTaZ3ZO+BRoN1LVW4AZYscPyW8vUC0PqblOQ5XfHMbDIfjF+3
C+awLtYltK7YsUNwWgrRkNxOVZSvu6/yk+0YyFzf1cqdbsT1OX0K80y1NZfHZqIm
oDobP/TOFBGAVrg2r4eJwRgXNejCjiW2fvc/10w90QmI4f6MKG6kvzKThjPGN0vJ
Kf9DBdLa8MfjryDGyt/wq7xJoUs6MJziMDZO2QWdoQsmGAZ9ZGCmXMojrhX9Bzv3
eaj+USooUz33cViarqrLQ1y8MWlakowggWm9dasgUW+79b5dl2gg9Kv7JkYSHOEv
hc/rRnCwljPt4tbfhVX5klqxtZPaJ1JAxcoHG0UAk70VzWYNUo9DlixX7ZEQ7Qzj
O6o+1+jFVVliBrp0hjliuMl05eaENWL+0fQeE9oMF5nK5b5veEwB1ck3/M2Jfv6X
c4NSAgazMXDXYhukJu8VWtpuNidNDSwx4JIbKKxN0sM0UC5MKcgN+oM2E86Czp9M
EWJgdOrutw6KE/O7T9azk9Pi9ZSuKPFK6iIxLLdhQxcY4WP8Fh8qDfzFpvB0lGIX
A5pSoTb/i/Ip7m4P2wuPHJ6Ei44CEFmHuguwdWHfdHQmzOXIk0e1xBRIc4yK3joB
ov/0AQ1qqJM9wDIf4WtCqMF0GdJemAGP9EddHKg1bDBRbeAXmHd4H59Sb4Xq4ZNt
2leqOF6E7M1E28CiHwR/8C1QlwI/WcKWTssMq6XwoODLUD+Q3SEbNaVqOPOh7ybm
FEqp4e6fnyQK8dZwJp52CcCRwKUE537Nmmo+QNkyUVlQdHRBOq2/L9ycLUT/bj4k
ZoFSgDMYy58C5M//epundJC4tkhVNHasP88abxCuYZViq0uqa//xA3RmVDYkZUU5
3qFAA9G6rYDkBPWg3T9+OXNrUy/xX3N9H/EAvFjAXyYihqhS1bteyHD4yPFFhCvh
HKHsoua/5UuCA1I44Nn0LT/Toim6teAaN3EubBsKTrst3mFycOIaA6rfyULB59oD
HQi328gEmBBHdxcsBAHFTonY8JX6f8/L2Jx0fpPQPWlmNKESgxapacBap3oqOf84
fpfYCoIC5CzNAFpUbi6lWVH1bEwpKkhxWtkgElmYY8I++i+IiwO/QMT6PinaBheW
deJmM+4w5Di61Z8FK0v/DO6rVdI7Zx/AL5PUZaOTqOd256d+baKox/21422WWF3K
qM5Lrw2kH3VX+uWNjGCPQyL9wlbZZ2Mrzhz2N62PBLC8Ui5qTHdm/gwpVCh9Hp0Z
TphquiNd9oxkFGCLN1g3ofxHewYfOD5Anlxd1kZ/bYbRhIZYpQ4Cfouw9WbsilSM
wETTk6ijIRoxfDR5ItsDwpBJlDenD+8QFqdWlsBDBWwVaYodTWRYvQR+K87rQBNY
Kvf4xMLZag3/io2m80T+eQz6ezQbZaqY4/PAdhlHiZiMNMW4buFHEFVBlPfV+TEC
eccU1YUBaY/jpfbu3Qt5I/hIDlFnFTaJfUXOf5eZwaw4vOth3DE1CH8LzYqQXisM
IfMvIqDel1ZHW7dGSex39kkhV/mLA/CkZv5zLyb3WKQLa8TaKUalCxaOvcUXUT9k
HkvCrSEjasZybEVf3hQziqpq/KPzZ6yfqt5pt9NwZ+0qdr0MpizyPbM2G/C3dRU+
CZiUrfIQDyp+Qd6XJAuysfzi+WOIGAdN7dCTw7vTjAyGnv5dR8tzEh5ThC8OU7vI
ygKUNm2f23iZkFm4kO6Nwhhg/hx3o57mF/gpWWPnK5JEE5CNAZFpA4OILiYSEGja
1N2PFbh+HJHVv5bhuHOFu/+yramUJpBI3rIy5dEhSRT2q96TalZqw6GnOa7M0GZr
DbBei3zzzt1KqXWofjZYo+n0GJqvP7MTfCLip2CJApVclgSz7LGSXuQ6EzvlInB1
j5FkhLpQeksSEpIwIMrU2Ha2Z5Ljj5N2oF3fAXV8qbL6I36VUUh9NpZV/HYgAAOb
d/EDHfWIWhCmNH7Aht+FZVkYGzfeM2tCtS0eZJh7oAofcUUfMZSMLXnUaxj28meO
TUj+llje3KXbt8mH8vzk0Bd+ftmDSJ8JrypmrL11DEBYMlMVtchIKRnwgqpZ8Dpe
TShui67Vq/DYIdTtZxZgUgSn9tFSkmx494brrFWLP1MXbZsfYNPHag9dPn0JbwO7
YPJpPFmvagjsUPgcqJ8+/DFxFG/OHK68XvP8Yn78w8uVsX7h4vPh9WwrWYPhaeNu
ohKKOBKB/QfoCEsyIKGk9E2l7wzTx3/YqtNP+ib2mO3Xg7bIzlyUaNVRIL1RcEHt
7AVIdlmn3B4KnuZqq98ZGwECe2dkdLT2ZQmTIl/uMUyRN6NphYroAS8W6Tsb42sy
ssJgAy23paDzliFlbH8XcYSU7nAPa8MmtBFuGdxCiezl8Lh/CqyD7XEBh4odrBHi
30l6UsH49FgoBxT2mLdaSzudFoUbnfuT+6JEcPztNoKhW+dTkEe9wP+wuG06yX0x
D9ZNmjx7Sd+tbHAaHGJnn/R7gVc7dztVaaYoROfRcm8WpiZcApHuF4DWmPjoxVU/
VhvD3Y2cEh1/Scy1uVfng34viQ9XAQwlY4xO7ep+u8xe5wbN0c6m6o3i1F7pPl82
jaIQaTuEOla2XuSx8pu+nL4BxpDBAEZnEOIBI6qQ44cG699ANuO3c1EORuiHiM9E
lpuydrdJwbw6DOHxW2t6PJszay1xm00EmGPDy9ybnYLECCDc6FfQFXzhrQSBp+76
+XM2HAyLncqgAnfXzW81Yk5HtkRdFQCs4OJrOMOZalXd2z+vKmqmY0jetKAEnxzB
PB9QkurgKp4EiFFVzEcTZPKWRu61XR9t0beq6Ip255ja6+70NVmOZix1wtVo1PRK
8wUnuu7lpGek6Px/kZzgs0wsIQaj33OiO2XHryhqKkKIN5efRzkud57/RbRxkUf4
U3DIn4CavQJnMhbv4rmnFKddtlzGLBNjWS638C6qEt8JnVZQpmVAHWmUcnrtzK/N
DhYizRBb9C4ZX62WimGisuPImEShTeB8498Z8pzzurdokJh0FebgF4gtMlJfVTGG
Z5cLq8jyxMrK/Bfzhp31cENgMGw6ShPMOdxpR1BK8ByrfU5jlm5iT4P11xQjiWTP
uK4vVfDg9aCBaZZLA7EWEv4pmewWYskdaOIpr/v7DBfvGtp8eeKU7QTQrlRMAwp4
oVD0yY13NTScgt2aAqh+pTUut+p/ae3LTDZE8iEXPNSq/3gdOOIFYLHN98pioekq
1uGEMop24I80hrHg8rXgce2OmYQy/K31AWyV7q/L2Lt24Cwljs0TmszGw8QgIZ+k
iFa0lS5yxVxR97fcJlJkfvqNOAnge5N84NMeMTnHWuHRfjjmr03MMBnHCn1TTvuw
5RCzQctsyhtQQYNk25yoHTQaBJIQ/UDb5d/gXLTd38kQFjPJOr0tRLm4t5M2QaTq
f79x1n46z6QqipGMhcxYGoCzV+2jGEhOgWsXERHP+RJfDlpnvYm10YugdMVoqHJv
zGAiNkfonS0PS9KdcaX1/h248dtyiaMFcJLsnpsI0pV/OmPm01oTLlmIC4auEVnV
BXE9deVZVJWBnwYfmm8yOYskOkWq+YfSnjg9zgFy5JeV5iemlQKuxOx9Jac2Tb3S
bbpDwee93FOxSeAdhDpt7UrstPD/OBh/tOHeQRyLnt2tD5mAR6zRSu5AK/FKIgmY
0wnLdEMoIZe0xlJp+7Bzx4c0FOENPdrwKe4HQ9DpUtyolMiFCvVlaiMdRJCNH2vl
Gg1ya02qmFdodXfFJlwq45j8ZGIxAZfon6mqYSq8Q4cl2ziQH6X6V9OAP8DNfKd2
hTyIz+q4lCY3DmEUyR27HVjoz+/4WzgZJ2B9R6qOviaWek4F+veQZb6/tMAPCgxk
aSz1PtAm5lU2BE+6Ny3ThLh63fZCntS+nqusBnLxtxmnoP5RmQe/VvlljXF5KO7e
JOqExPu0HzgjCbwA+EyCZhuniFSClXHdFygVt6iVoQj9aM9Zpn2Kc4nR1hdl/bf7
ExbMUsdzuMoM7STlAqsNFGmhvu3n/dW/lkLiQLV9+85/pdU2PVMf+OO8MNkcNR4q
byZFGaPG/AV74KGs06WRMZG1IXkGMZ9Bj8fR6V9wV7I+F6y0ae2Y4ZZwh9Y+Xza+
v0tIe361sSDToCxWn5NuRJlZ2F07v9NB5/ePaGkkPpMbKtyh19MS3bAJVyQwht+d
aZic2TVldzqCT3KP9caeB1J3xC9EIuE2dQBi9Ce5STE5G8JUTeDdFt5WVVx/PI67
it2e66Nt9c5uDzUv0weowP0bk4Pg8uc1+xjLzWXL/x4MWJ7ZjSjDR2XBToybrOhh
7sLmh5hwQ4QveQx4z3Nj6/r9KDBPd1N5+N/kpuJaGu6sJWzW7OdRrqMag1pXC1W2
J2Qj1pmKcRAKE5VrgXzkLhpImV2RBS2X2XwbFizssFIsxMddQki5fP4cPhSDq2Vi
7Ak1oTypd/05CHyljhQGvL8oAD5HlSEJKEUlrBa7vh60VtOv9WFqyWA54SQMMxor
P2b2dP1NsgywkFXVMu7qFQ3/wlJ9XHNnZ3BXOQMQeRXszF5Lg4ylUkKt2OhBM+l6
MNYcNs43zGiy/Scj1z4aZ9uOQNjvpPBm3MmdRMf+tp0iiL/XHlIZvHSkGSye3lME
AqJ32p3oASdr+4MEcE7oflE16P62JWqwNY8g+kTuQEy+qhsPsKv70d2qTHFA/UIH
Y2Ax0FF4K/Ku9ZT4bNwky06kyk2uyM9+Wk084x1yqxGpdAafYs0og+h3dpwGLj5Y
buEkf3FIKmKjsOrtzbcF7+Xvh4KkS71h7iQSNhspRwZtOBSeWoz4BJoUoCR0pjrj
TRjTn1G/HVh9HMeCf1+BX1NZVolCtZuP+gQ7iAldzTHhiTOHRfo0I1FRXdttmHJ5
jLpbwsWH7wdbm6H53IYH2ljOEBJvq6OW/7HzPu6kbzl8Pt3D65mDixWHLlnFKYjL
j9egfaEMzT555SXuPmeC6NaQL7IZjTKuUjZhmbzAY4sTodXskCRxg/wmWTr4v2D1
o/WMQ7tdGo5FOkLmJA+igk77K83zv2QXqG06m3VU7qYIXF1VYkiOQ5SCnGPz8EOS
IJ4xJiNkNi9R9kaxJ+9QN4ASvZN5xvhD46gxfxBIFkMBUbvsO4x26Aukz+BsMiFR
QSdrMrXcXcMzgdbCXVbHjs6Wtz+Xn9fb0S1FyjLab8NHE+09fspayRFHE0Ez0qqo
stvobXBFy+RrOvKOS1E3VJIyUdYIDZcHEOrt/PKuvy4xchFK5wGVCGh/BfPIlNCR
gLgn0KkM0LiQKi4FeitiS6j6yA0IiqwY1g6CBL7Ty51a8Qq9ZJm7NFOY7maUoKA6
yRvlpdEVoP2DOd1ASb2i4K6eiEWZXJaY14WognfDUZxKtebcPjlqpmmb0PucYzny
dGsOr+4YJERitGkWMC+1Fs3tQMn2nYiMqWwQEfiF/9c+q7qDRoHjmTikeZzzZ95e
8D2BVmGy8R9h6opG6RCPtwk4ORL1wVmhkC5neHzupydICIymxuyWi/bXHV59RFlF
ZI+LOsN4BMxlFZJIPEjeGh8cEhc38KhfuR964QhqDQD9kwh/7Pgxaq7ypkIkju6O
niXlw8k9FDWh2ekF9WVfpx6pgYyJ5oS3SU+wN9Z4VESj1lVaAcsG047lk0i7KlmX
fLpW9LgIM4bnNKt5YsAjHqIFaLOWcI1VGGJiIh7/7SpUSCL6rNBbyZouIxfYNBgb
huIygtT807iMzeH5ipIWHsa1DHNYsxFi3PBciMonu/h0z05idZJ1y2yxpVZgLBsA
zCcNASnkdR0gEk4lNEEWNqZ7Dz31eEYsDxPoVQ+vCK4zfP7IrgOnIZwyDE5gBjas
d1yCnU4HWVlotxD50wHjyhjmbkoD/T2dTKWWi+P7NGDsRY4elZNE6LlRwXsDNPHr
YasD82Pc3zEwkA81HP2T/yjG1rVmxsnzxw4r+eX9lLMdVQru+S+j/vfrpVXNaFG3
6y3TOGzSesU3bOXtnzIy8BRba8gybDNTjXxuJcUvdpXJp68nyJOzh9xjkVbBAclf
VEiwPEY/5mHiDEp4ZAnAVW0U2OYyQPQjB2THu394uccNrmXTlWrGSweJcvX+4pLL
WeqJ/SoZF6EJ1D7VtWnIcmb2PJXnZwVkNgaq4DXeWJPzUkQO+/1c+yhoFlALAXfV
rgq8QWihi39ZGMOsg1ZD8Tif1IkdfgbbG1QQrSW3XuTJpS0cGI6Jw3+21Rn2NX7t
r5+FAG+RSybbeYntjWkQooYyKuOUEfwVjv+2tihaLOQbSZF9bfS5I6YYLTtW1Lhy
NaeNLgWlIonIDd5Jramq16e6oAYlkluVogltMN43MZM0NdOn2DmbZWxyOVYNZJ3e
1tbts7A1Z0BHyPVH4fH/lwy33rTDDTn/vujNCqetj0V9AOV44+NqiboGllou+PY+
gprQKBKjfC6vhjlPiIRSvTLebAY+5eDYcHVDFv6mu74LNmqvbv6FrUgRYdNry6Jv
EvKta5AVw19Pfna7acefCENSKYdyCPAslMkP17KRx4X4paYCrSmYOigtnKP21Tt9
R/MMcV2hX2fr2XnIDcbo1/54H5KXhEXIcTtP3VHohDA4cSPfgC0xnqy/ISQmJgpd
f3EgT5vcMItfSlFYax6i49O2RscdV08NZrfGF1scjE3JFjhM0Bb/ZppYAZ/dQeO7
rnL4ZuPlyBgiLNgdhv3yg4zD/p5aBfETgcndElLVzYCDP+zqOR1PTpNtQbbVoKPB
ukPCzQx1Cxv9H3qwW7rzJ9R4jQeyVEwwbUnolKyYhfhSM9AjKDm8PQFP7YJzyy+f
yPIgt9GxoqEjWifg3z2ic/f6C9cfWh0qWaAppbNgVSIKFS/V7lFcFA6rSYPS5fBr
aDeUYA0kMYY/F8P+qa+vEu9kOTAWWJpvuCKYUY1wj8L04dKRifbTq7SlUYSSieYf
m1cZXluHSd+vXJVPAIAVdMT7ULLlK3rKfWlS8LBnWlqGIwTRJtRqAXpd8MXvRmxC
PX3bmmnEEMoNS4oN4hM+UPgtFaZiGvAlfRPdunIko+9Lbxp4aqhhKmDx8FedJrnf
GcBFxOJJyQ5JckaJnyRx2shZAZtbVngxCrK12S333ysgDmq7YIUyy0r8a0TgRuM2
dX6CwuSv9ZqKfw8bquLqg+MrO/JMvxzaM3gQfoEw0F2MYfrIvASepPvMIKEQMnfy
+Aa9w+1Hapho8KO8JXtDOWa37lT9BTuAcM2rXtIQHiv92rPNCLXZYAOwgHbZZpke
zLdWci7i5pryxWlyym7UzeUJPW7HSSM2lY53RqGXQ5jN+vnwNwjw/20BXPtnYI1r
TpBmJe0fiNHHzRacyiva7Iq4mLBlV2byoUyCmSoz9pTwniXf35UFuc/vm8QMDjJm
g8sb7zHEcWJl9Anmu7t0g9v+T6/6vTGqAzZKdyHcl3+LN8MGFyL5bTN5lu05xjJY
yR2mA8V1VCyauhxbBk2Z6ir0S1t5GYjqIVpmDn3fX+hHKUDiiKSHfZWiXhL00JKM
Gu1dQQqbQ4hpra9MYh4494f/iWjQivy6LoZVs8WzlQNediHm8whZmnNo1cU7YZE8
ExNqG1Y2jKelO4X6SgEFWpOytTin4mpTGEQDU757zuf2SrRJ9jHZtjO2qGfygbBC
KokUTE/F98cBO6b5pOvb1Gd7i15S+OuyFgQob886Dx4se0omFYXLfLInTUtSLakf
D57amIAJArIQpDUc9yRfBCVVTIQDQPkWXQhHI4Gp50M8nSk7EqkxULzHG05LjoPg
cyL8TI93XCWnYpB/5cNT1XShzcPxLXS6PcdvJC/TCzES+Kcsv1s85XS6NwzRdAkK
VzP3On94Fvhx44Akag6MiUL8jHtZ3Hx3yeQcZAfPXJnKU+mbwU0Hvd/I7CraeRyt
n5o65joW2oEDtOd6c4cP7pfRAgW78CYffBgxNZL1GPPY8eFKgRO9qRZexxIn1oAl
doKt4XIxtMZkurMo2g4ee+bkHitR7GsyyDuWsm4Ywtzgqr5kagEldULGVviIU7aH
pa1PksXRWIQCH9/oH5LkXuHJjiTdFTqZ9EFXokPfkEsIJEI3tpcggRmyUxNcJlm6
iAGXoMom9Lgj9J1Ai4iHy9raTkgEBSSjD9K0m62VRBg73XOC/a8XFRha9SHAHQnJ
Cy8KbvUceKPJtG4TGCJJfRbvKjFG1cXu1ZWO4Z/JfZNLpu7mSmROE1aEfe1iXSgg
Q1nlme6YZdqwkGKaljrSUZEC5oOEDuIYzTCdeTrhB5MCcxEfiUDBGQFPLBv0ZrIX
cjcL5xWe9DTK4ne52i/gG8/1PSa0ZWTMuZNS0K8DEPXQ9QK6Hv+rha2Vz+Mv4Z+y
oYeedet/BsDNxpm1aX5kRSyi1HS16Fv79PI4tHhFCLn30CrJWaLuLcgeXn9R2P3q
fSKSpKIppEc6OYpHoqJHwv78zArMAbPNrTMW4WrDAom/i66VG+HZZWUka0doE1g0
yD+M/13txh7HCneFOJaKLzXOPzYjaxcZSK93FPBPCA9FRAWMmoPmCb8EK/Bo8vbz
u47QwbDRO1FoXncS5l/H7HMLH5pfRmnHresn9TGAmr/jHwR7TeuSn7k/WuQz9HT/
E2w81HBMndVIMV9muIR+y9qj3dqAPJbAcn6M5yQ15WkabtshPxmGK96zp/IuMnm/
0j/wFZXVHFJSKdbNEUxPyDMM9SXJFSUl2X1F3BeuOUj3BIFuL4c1ioleUDY8vh6P
3hSN9txGqdGOObokQeI8+OZqBhbmBFTHoaPMFRVJCPmRY/oHh7n1y60ygEsWDHkw
rYqWwEX30To+UmC1C0CpWYSPn9kyNJPxwXakD7bMV8+2UFP3Hk+TFqBxk31YLa4j
ZwCTPBwxz3MD67WqvYS2Rrk0OtotEguMhZXvCdwPWBvL9ZDUV8OAQ7P48jwiPxvz
WY2h89Acc4b6xOE4SiWRhUbbte5Y/rGdJ6GitMwlhrJTomLHHHYMKwdV/5P/aYNQ
Oylupfe62JWvl0Ho9OTxhIlqARozIOUtNZSAhe6F90lLMXTkZo7bshkm1XM5zZxm
nWULJUMHSwmSforOF9CfYG/LGoeXsh55ANKkVcuHlwSqSqVwehmXuYbcy/9zP8kr
X+CpgYceohOmi8MaFd6ZoiOA2HjnFr2qE9Qqzj4NKlWPbf/xZMx6YX3xEzlOIw1Y
x9FIde1v3aSCPp9vFk/f2AcWOcirUa19VxyC++CiONlWNj2kxvnRgxo/txZg9Hpy
4F8hzPelSlcDYWOJ3+vaxXJPc94EOpjPelMMKrdph/zDgY3mgPCi6a+GUviBhgw+
idRams1WD1cy2oIeiEnYHkGNhlm6FTsOxbZzMQESuP1J5j7W4567m4YudznzqG3s
LMnI+nSAOeBQgEtvLAP35ms8IEQkXA7ecXhDegBnYJBDOeyZSXBw8GrBIsVrzbkh
QChjMXvFM//yryoO2euQ2Uh7Vqwl1G2MS7LIk+1yCFM0AlXgisvkuhWShznQQCeq
QQJ23VNUCp6rX+0zbpWHbjyfDcJzSHbke7sAkXkJLhnaUbqLtD4z08DinAQcdxqK
XR0gmR/SD8J3YtbjhrnZPTC8qi2FmZ9kdTx9JrRM5ZLWiJocR+oMUj85v+jz3b0f
nZjNWWj3gj3x5DMGhU54AkBhFxK+25z42cTGNCHi0Vm6JTOnvBZ1zM6ADe9RQunl
+ZEObCSLs+dYXrx6e17JUgOtAxByAeccpfpmYFF1HcWEETaY8cFYr27h1iBm6eDc
TbcPU9pidNRK0qGC73azh/FqQapxSRRN8dPnLTQBiJO+BbnOffIfa0INC6H4schX
2JEc8n5a9pI4wcEtu97NwzV4MIOiCQu4K85hvYDf0wgdORxgeezgm49iOtpf7Ng2
sXi5+oJWM0HEkCuIYGz8kguMwELyzzhFRawh2jTTpSjQtewDHTcQtLrdfvAJNOse
NOWobBcwMYtERNay6ZZpaS8mvckZ5lkBUMzgFvErhXUQAQc2sSz4C2tqBfrNK+1/
tgu+ow0YkMdAz2mMsAi1Ssfe3UKyApwQCZUd+e3K3xVyAEF3DQMRC4IEM0bLyHDK
jrdnC8jkKEJ8u1LZrSTY+DZgdJQtoK4tSIclQRyAfH5Hb/CW7DBNgllRYWT+AVhj
XBwxLF6tNlBs7Hlaf/GImlvOkBIoLIWIhtK/G6qbCZqg16uyF2r1LlAlGoLmk1b/
ZfYUMjDelzUB9KABWsw+FArJuMT64Yjk0GvPNtiShN5SbPFlLAQl4/5rASPoNK3q
IdziwCH4zYZV2U/PIKzM2r+T08CinhidXz2FdrW8NDpunO+nlBAKO8E3jZzEusMU
qAOdK67Ld+C/hGI+p7i5ak3tmnnY9ZlGsMOW10E0TtShnwPIqT8s80eyvd/Db9so
vIhS6bB4yAbWU2Qk78ghLa8zirDu9TBO6jgPECmPSVrZZTlCKHpgC9K0pu+4HYuy
GStmqnt9U61Ey9H3O7CYl2jqBhZfoQk9yuFFJ3mftxNq994jfijx/zBBRIzG+2Hn
0FGFvyM9RVC+lgAYz/OvlUdDZbHoeYtm0lyGB91LIrNCUGwxmuhG6l/p9mYV7YxT
Rc2P6hM/xi4KNEx3rjjtoCi8mDC+yarq2+JKVHwDP5oficR28JCW/eKgIX+09QK5
SPqm6XlthhbkrDS3DB80jgWNmSQQS6cDW2FSVPL2SKW6gyr9cTYHXOd9CJG6aciX
gmlicLwckGd5iCuOs3JVNFHkXbSblrub7Odzjp68azcSjSaQJNHU0urKYAmcY0HA
6xjMJds45lHr/+cfn2knDM9sEZc0IP/rCeJ0uaOuc1H7CFFcQ4Yz5u6ehXMwTZXc
h2lKyv95tvqdoAAC3AMRlmgWQD8irM/PXDNQs9HaiktuB7nWRRRXAv+TDcwEeI0y
d4+kr9CUtAAET6BpbQbPBhWySEgcjuARXvqdsWl/0SaKrVcmwOMzTwiij0ZQebNC
pZhsHpJ+ubegF8Y4+xZChTXsmj0tXhq2vYhZuVl71vxuZYuPTqvcl8NkgUjT5XDr
Ae0uuzniA08ThxdmRPNV0WMA7qcKW+vo+zhP4Nxar9CO/NH9ez4yUKQ0SmDK0WjZ
yaf/vqKwSIlVzhEiwSc8xI7ZfxSIpablTXKsyEuYwIjRdIrRX7X1d7FfLdCquqsV
Ecv1WMv9h1m2qHEgeH4VqPwC2PrwIWqnVFzadDzrlFeX0QxTU56eMPSB4fr6L8ur
Sql3sd6dGSEATF2I0uPudJKfUr5c08G5udk78Adqm5N7ItLzA4vTgfTaCk2m2VqS
7KtJNHeuvj/fY755/0vzpMpmFf7KEKn4ARttSQQRVse12mOih9jevoGI+jYAcZJG
5oEutbWP4msmdivBtqZbhtgzV0R8FEOjwNyHdWbxxIpaj6qvr8/Lm1KrB0ejf5VA
P/2cpGN+MPN/49GJ6vF/cj+OaKcxocqquHSD/vxvfl0XmdqP5nbWCHBaezrLK9a/
Ts8QS+bxsywpJMnA4l9wEnYSBzkAgNdO61Wwe5g7foUK0KMD6IysZ+9+GYEVWzeq
tRTrKLrFkDB3sXo62AanhGaDKTBGn/d3vaBF/kjY7x4nGm0T4n3HXOhLHJhQmxBE
j4oCbNmBlNvbdwIO61uqhP71hJ+IE1675Y29SxW3K6PikZmJKxSF2W6cPk6rIGz+
ZHLSBisWFuw3/gBN1swFmzuu6WrgppFfEsfvGHvYIgOgWEhSMhTg/cKZzQOxb30n
jbHKxLFkpJajvrl4QUD8QNmNp8YRQBMMixCmT4ECPUW5y3v3FrAQZq0wvz6VocHP
MEpyye/Oc+IQVpkmuMVK3BjVF6XCUUTIP7003/JtV1oh0LMb3slGp/UGc87l5P2X
/LGBqktiaCvvVwaWq8GHjRPFF3xzEZFn3CMlZmaXlTcQyjrMcHDvpjFQNdwxAsK8
clA9/Gm6ezTCHYwn4HMzC3TerC/oVYowbXJIZZrlPu3yJv9TscPwYU3OK3bJhkrb
BUOv94Pxs3NNWtVQ76hvjwu4xgmDD4PzZN1snJHDvKAPzx9Vg17DaLgfntm7veGJ
+oYem/iCRgQQnNK1pMwM2KWhtge+JlKXFLpnDe9lGunGWoCOkVgo4jc7SBHrrc3z
XDfUj99BOlSVt9I+/shNEnsFTdli0r4GcIsMGsWl3dUjFYrE2AfU/6/RBQXbnFNN
x0ovEb+hm10flBJuCjC8Df9NXevLQTzBuHP895QYJWnhLIPm90RYYUcuSmC9e4I0
ky3SjQm0xsKJkht68QERFp2mbahGIPD9pU3nTO2tye2ySQ5eA/W4XmcJQepDrcMN
zkkQD/8eEzqbsQU1Y/OBO1B+XaL1qjc+TvNQyexk0IO48f6eddXPwBHhOjfK3SF6
QoWblnXZnib1sHXfQ17QrJqUZZXtVawASCYt57/PHPQfgMV6mMAaMfAeRUgNG3Ip
rxeTRXPmF9IRLZleapKPdbUC3V8Bl9Rl8xS14Tb7z4QfdTGiyxCPd1w7TmZReB86
7E9vwkxENwhHUjpN6CqQsKoyx0kyQFVJlLiflINRDLKcATB5G00jyVa4r70bCe5v
dWOAQns99GjSNhitUXvu+yNYwTfYukOYqEMhCAbgFaoYfDtHfhPuxlZO/EC3tKwW
wNE9EaB6MbL9NKgTGmbFqUqXywYN88zZTpmBnMF3+0auBBcgthCSC35LzrTSqJU3
YgL38RC5NRAxwZBMS+Y+wkE4ZqRTNDgl76jxlP9xl6Ib81Hn7Gol+OqlaD8Wcgr+
gDqQcMFFJQbd6cfQRl5cify/AyjtCl6jYuwvuTr3JkXFoA2d0AFtRObO9LiPkRz/
MWEr072L2Rs1KgrwhTMwERJXCEbmn8kSPmN52SRgfbYyiqB3VXJc26KubJGOlleU
QjCmwV3IQYvg4E99gOjtR0oZlHOS+g5uDGaklZuYEQeL7poqBJd8pjrVM9wYrFrm
5QY/Hp5RRZ4B5OPWGU/oeKvqmKodP5Xn4y7cIRE3tIf+wj/gWxAJGNbJC8l4HE+1
HGemmTCEa8+cU94UQRaN0UJJAe9HbSh+cAvfc83xb5tPK5BnAQQeUp8m+qLjR0SK
X+6HqzfxSnIGrrn5u+cV6+B8tTowpcKHOJIl2pSkaMwwfkZSSICG+hdGcEaQjBEg
9t3As00Y3mW3INgqnY9ZghJHi0r1mfAhnfZKqc8TctY/E+Q//gKt85uoji0zqYRx
lrQTYMu1KRVyVjAvrA8CArr4UiQJILZFaG3bubiTcLTLW4wyHqzv8H5WP3BDve9M
8Q2QOeOHHsJOp474g9LzMxhkc07xSl5SHJaUZdttABx6EJUufvwl2VQRX8XvUh/a
O5GYX3vRJCxeyn1DCrpHGDRgttJX9w+DBv8H93FjPPbrLKuhWZ4wGDS8UXE1Zcm+
i+nneSce843g+uCopUXFGcyCHwZWq8JPhdfzR2mLH0oFPOdF7zRCgDe6LEaSRLo2
HngIGG+xXcStSwGZXq1Coxu5SuIv8LZsQe+lhrLaekK/sMDXaND7hIJGh1q0vmvs
OM75OwiZ+KFxFrlx/nXYmT0HSBMwXfsugO3MaSKDgHelxByBVLMu3QLRDH58XTpJ
VJ9wV3X5apzQjrkxEI2AYOmRTS6GH2ojwt85AyVPMnBnSi7QJcGDfNy34qBUlhMx
/KjzkyNjz4RDAeMJF3sVQEqaBl0+RrlN0o2NAKQP9hSfGfLAZXPSYjpI4lhf6JO4
eYyum8f5hcTET/0992NiY0qMyBePVBg3l02e2RrInnk1snXyPR1zkRK9r+3XxPI0
jP9Ibcu3oAOGTdSip/jrhTT2ZastMJhDCmdNounnOpEVXAiQWPVTWzTgLeSjBZQ5
eK/lhZYt6cU5KnZG5JoZLbV00G6pvzqiWeDnDpAmyPCPFMJRE45qAwpPAx/ygGVR
+Rh2ZMg0QCrwLFVpTZ6FIz+kGsUwv5QO9dagaPERmULi6msfd0of4ATIOCk31vca
MN5J9Hu2jgwe+hnJcsp3qOpfTE0DUYqW89J/JJ3nZU4jOr5G3NvpYlW2sQrnZ+KC
HcGD7RtTZwKM8YuWX70wR+p/Bc7zzip+L4RXho0UnXKjEYMfDA49Ho5WRLz1BVIn
uQp3Z5TCX/exH4LkTbR0Kpki59TyTXhDIv5BTnOSNkbHsgiJR3gTTuxcqHiE6ztE
Hbbxhehfq3tdMAjmovpIv5HY8HuLE/gPxWquhHx+qVDdLbUHqPBSEReTFGjxZxp9
kZoFDquJhDbD6KKCfG3mqBi+0ZNkfRmbAq6JtVabJtAVhCw2Z902p02C/hanPzWz
SkEYrPANE0IhbdeN4WTZ4lty3+uD1gaUAkO4Y0o9pfNFSuF6S81+bgvX/8WGiZHv
eE7DAU31Q0AAwhEDYHmRewhMkyO+A+s1/3+6pWjOLiei6IExxRtoaK4uEQe3HhAu
61i5TT7iygP3+FlR4oc5pl0qm2mikTHnzv64HQrLK/xqXR5WQrTHqLj3zynF+tCH
hR1tH8+s5DowiBgENQnnWS15c9XqB4oGr+RZTKVmqABWKg+6warlUfCcEkroHGaP
aWsqBhgd6lvTVxBYCVa/mmliH8AYuxNsnE/6fzjH8z6SmrHAI8iQqrYNvz6n0Fyy
rTpgqOcNUPhx4qsUSkvckE88k5SHr1sthh7VvKEImqdpIBiD2s18iUV0FKo4l0ZT
tZfu8NGHrVzk7I6LSr5GnJOlIHkFmBu0bTirb5xffE9fmrxDUJfKDGZf09BsjNY8
aVY5OKqKuiJciMG4ASb6j0fGz+lwK4/lDnX/1LQkuYbsy7oP5VvWtSxzzV0J0OCO
uKkXubov5bs8blIZMwt5aXlRuiYnKYU9vlDfpw8Q19i7j0+2OIZBT+f5dgYHt00P
DyGpuAOiI9wNaiMAKSUhWERV50bnr05bikb/8mxH3YVX6e1vAVHn5uc1+m9Di59r
xjeMyCwbhXUhN2otGoZHVn0rCAy8ASnuJ8eRSyqKQxuFtSG3Uh6aoHkcPqKbuFjw
dfpF8P9/jHdbVj5VSusCcPEUm+dXeaNs34Ih/ijkgUkm1OM3IAUSdXP3QzkL64vE
keWm785v0N4YMnhOzhBn9zT+isrNzLr6+JppNyHZ/dpOnLEykZ9cQ4zXXb6/Dn/E
r4a0lPvlrnvJwLT+RZzs+2237XAjtoKX7xa4pnMdUsNOQr9ORLJF4Fq/ZePX9tBw
2BI8r2pZr+DQjzu85ZF1xpilV5TFAMPtkwkM7bqfzG29MY+jKEJ6UfnLdtQnbzOc
hVSkh8wvxZJSQfaGawv+0arZIIzAcWE2oeQJlQaYuY55bfYe8JCDBuKxGezCCze0
RFc2t2MXgPjIlVb0UGB7rkAIupEla5L6tp5uhGo+/9tnPuGydO8y2L20ZxEp9gpo
kHceQrCo0llDhCSAknsr4XqIOTT0KtezU2WcIDZ3TinbwodVffwjQAjDBWG97JKD
t36v5Fj6XR9ucrkHSDmxs935RqjAnPnOJSJkoHqZ37+LqXQwPo5sLLM51XGPb+zx
sC1+Jy4rrY43Cfvb+4a+q53Gu841JEzdlyardBLO9DuYDBBfTqyn3WRvKAIc5Q3E
CC2gf0CW8ugNgejWe52vSvmoPKHgeVNxoYHeTAccXoDnfs0doPxp6wh18YCHArSx
ObcJmA4lnQWombaz3PB3d91Za15rRTU6VWrt3LGMqvl1arqdkX2FsEBjN7b2UdRs
62IfOd4u7omsqRPOIf8ednsYu7ihXkMbmm+oZ9ValUBWnRfEC8XNc70cPYDCyIeF
x+8vmiaEcXUtk5JPMrGzEOZQU4bUVrvZc8nfzg1wffWQJIbCwvcN3k62jtJGiiCq
5Fwoi/9XYRfnzlTU9Q7mCsNQBrTv8McW5W/DsL0uxms4hM0Wgnkf6L2+4GjLdK/z
bqwu9sO5DZ+UwCEp7Vd3MDcPvaBRdXFUZhcUuvRYKZQtFOAz5keIVhDRgvIR+38B
VdW+ntJwO9TA9j7qO8IJWswlOx2sTR//8BgOsbc3uOK9ZhzqQnpYPFB+74eyyoqN
+BT2SDNKwgD1xlBD14yCgxdOoq0k8uNIX2en88Q31O9DRg2Z6GYz+lh+3RZ7bWP4
YCmpsEn1PPQFyW2pz1KlEJzjGWXnQuUpUaTOw4d/qAwLLA9vHBJ5w1WLQBmv5+F/
cetbVZaiyeqFgMbGxJSH873qEy4L6JLTkyKUMQbaUDkj8n7FdfkXCeCtcFcBdUWU
H92cZRrgNb+O+LVvWeuzvKxc2UOstq6dHVQEU1h0zxmBQhWmxxEgn/+PZHStRXsi
eb51gMmtA94YwqKFKMP0Xz68IuVRyiDouOC5btWGoNccu8Uz7moCCcuKv7kvnUVD
UE2S/8vBiyqzCfieBGfmfHnLIuapCa2ZuoWpvDQdKZ+kRKf4TbTasXGu0rshi52h
DSeW/mpYBm+wSNOuI4topgytWuCa8YhIHM/FUzX5GXOENRgmVNHbpZwoxkay9WuO
o68+p1sKNj0YWWB92T37hVsuPgng90M4o6XVjN4AbCtUZAczYj0lnJst7vFA8W77
B3W5imlw0eYaA+QSPvhWxkveZPkrFJgCJOSm1fbpm4VCyVJPZpzxWuxfBGZpFjHc
ikBtjBfaBSoagF2RRc0JlDbSno8Nswji+37jk5ubWHKpsSRTE7pNYp9cvFCZ3eAe
8M1EeawPBzUcnn3S3uf7h3wTP+XniCGs4u0BFt1I2g8cXVesDJZ47Wrc2mH9Zisi
B0STHY+dXGz3mDGm11B6r+Bp02jjHL+0oDi/stEv5T+NBBm2wtuhKDg0tD7vMKm2
CvbgFGSF778l8hdWSBVcJ1ti2NdlTFqMayJm8G1qCuBU6U6x7nU23h+1FYy0eXBD
IKuY7lub3qlerC4RtVJpBGfhv4ZnQrHrJH0X9U7XvZARQUKVf8jSN+69PsxANCBA
IIFSVrV+gimjjdd5cUS5fmtqUFbk3Kj8qhLJFmmUO/8pWXMw03vcw+aNn0sLh0Li
9j8Qq5CKdG76liPwWKMJclUOGXzbVd7KM5r9WMrZXl+hFZ7jaeRokh4VkvbsPVhJ
zgdPO0cCvhJD8w7tmmjWTysaV4dq7gWIHi931lgV6JREtugIVuiINy1jAN1/ZN+v
8ffKoQej/7pFfwDRlt7kWnsS+u9R42dxrS6ri2IyrUIxiIvgx3dqPnyB0BBDKaR3
M27LXziok9AfLP2eUL5nxK/jLWOQYAeD/1fhmMeKYZPsXyB1KStoEHfZXelpyIhk
73xb8qzyaPVPpqlvoXjX3IUmA8SzJxbsgalDXN63MF+pZ2RimUKI1IvwBK3nytpk
Ve2BOHJHnuUDU0ACCZxzFySbxMvqniVGuY2mpuKdoFWijQNxsz1+q242o0Ectzm0
XpSyPdr+RD+Go6nLclvS9C3/pvxbbVY/ylGFDrLpPPCsSsAIFbRRQQcuEpGaToTr
InCa7csjlu9j6N/FK7TE9fLGX1EVGgfNb/A+utv1JWVo8XCKXp3R9tRWYHHhtsVW
fLs/PHmYrGWUU8hHqHdt+obEDQkOlOB7oJDpTw+3VK+qXIrsY+N+Yd7ekVdIVcJ6
LpJN1g5oZQlx6NYiJLXDqzLJhBanSYrg+OW4A21WT/8TzofrYWb9THVRwThpOdQF
2K/Ceq21McvAZNcC26xXGFmGYYritR0NJGRxny3fq2NXTFwiPpdpYGfeQeR8FDZ+
E9UPD2h1feVa5JVTTlHObxY6IpY4xDXr0t4dqdXZnfJqZ2uqjZJi+Yp8wCr6P+JH
w/Flhp4z4eHjkHbKXs5ycXDwVDuCpWb94XQYqqzl89Yl8hJ8E+O8wAC3I8J7Zgqk
k/feeZ6h4brsVIBnrSRzgWBm5ER+aljNaCkdvTPvEAV/b6h/eQ/WkapSdQJ8MOmP
3VuCXyFVnSJamPO7Axpdhz7v0r9b6172jsXo9xrY0GhD1MRF3wMfWIHOxiufbTeW
FD5YJu/vwLIocXxyLtLdt07EK6Il11fiYvyyTIHkM1/J2+NKYDhf0i5JWGqGZrXR
+HWWP6HbAbg+O3ZDUXnVnIsEeT/ZC+Dfxpa4QbVosh0pt4pgo+SEw2R4JCAHL+3j
YE0mudVCWiyc/s9IyB/UJQi7lfBz7Zz6Iv7kDKBp+SPt6fVYlW0x4wbYKmF63m7G
VneqW6F/2Qv+pT7AnZHTno+36SDqR6BntVbSI60vqm1qRc4RRZB//cqf9SKGyMZE
ocoRwqI0BcaSTo3Qp1gxBOr93wcOdhI51iOVDzoyDmorndON5w8StrkQrnS5L5+H
YSFd4NBSv8xtEa1fq9gt1nlMuu2pYIUZdyjfT0ad3rIYHXwRGSsumhCWDbxaEJzi
InbK00VtSGk3QNHFDZHojlyvj95vFmKHpQZzYYM/80MmktgIrZ67V4P+gPOT/Vvx
i/bqeuUInP+lysbb3SpC6lwQzPfYxebfA4CtH9JlwEMna7wEpCx2nCX00i9zN5Ya
RamU5yK61UNJ3xwwcPK3ivEZ1Nu04E9SjOqTlvFsqAevzawS7IZwGisyBaiIUPLY
6tGr8fCDo3WJlbrfF/5Mx/2+5rKu2o6XTPtha7vxuGLV9e9xe79HgaO+rdYNfxrb
OqDiX5rRH6aiTfXegSJZMH8MvMf0A71q5kXFemEloEg+TFPqtju0VMhEIuf8Uz5/
Qbqo66vuyITF/p4dP5YyhN1oF/8q8e20513iIrOZ7Duc2a8FiSHaeLXry0dZybx1
QRuCxJerKfH5cd+6i56vAZASoKwqzfMfpAIGWBptvNsJ0otgIIO+e/8apiIy87fv
uC2JuJATgj2cRm3k0bWlyICkY4L/mPiXlNjsJfvecEOP+g0gALfKToDcLE0+Q/sC
wVqi98OcEX6v1IvoTzlokJnEtNpoIKNgbyAtGUJFcgyY+uI60TJQUvbqdU3yID/y
/daDfd8s7tcIKil0ofjZbojgStZT8Uu8Hx/Dv5sEyvcwTdzHfMDOwJmYch/VXPpD
OfThR1h8O5f4r1kX6QFs4+FGN/9UZjuQ5uOf6hMFJWkJ+oy7mCZ5P6WrFrwyxzSh
+Q3UFVkjAs1Q0MgnSdaFjN+aiyT+bfvuTm8GAaT+ZI0VojkyDMlCcUh/QTz7juEz
KpzbPQAlXXdzr7CkThd72M5SsuHfgpUJ10Q29qCjh9fesCv6ZlXezRWKdRtIqe0H
tSRswcZC3MaD4zcWAEJbK+4dOSr1k8t1oeBSZspfXshWCTvjHG98jiOna1ToUT19
WJv302+nDGI0F1dsebve+kzrmk8+KLqqPRmgc67nTrHerr81B7yqjUNcs7lPxfWL
B3wgl1L+IhbZnQ9xNWbNN4ybkDZZqk90PNE3vYnUn1buAIlMbuSQGa0nrDNJiTKw
T7YcUMTpil+FNunH22rwNgBf6nhI/Bti0nuzzg2I5u5GwTiIGtwSpy61R9fK9+Vm
SqYvX21foquirqRLdRTN1xu0EoJonzGMnf6jsIYMWU7HpHN02G+8b8cQPFy4t9z1
79/IgSttq0izsE444DZLZ49ALgpe0zw32RbO1VRjIJlqwriqgUgDeUD94cL8Joe9
1gWqaYfMbn9aEP3IbGS5HA7qRRzJ8qWu/z9TKZz+ukr4e8fyAnfppiBIgm6+iP8Q
+N8jVYzZzF/bLZ7V19V4RELBQWFxKqNdU5nltfNuDPpnVw1LUMFrTOSXZ0ruNPg2
u66EAF0313gJ/ROCBe3erQW3MrXmB9YniPnAl1VC51y3NIXfeqQl62fiCjsV0YIz
qFjrvsHsk3ZsfAWX4d3PAUnMx5LiWLkbn/fgsIwiHJlaZXUl55sfU8PrhfnhfHcG
p+KLu/4dMhY9/jezSlQQG/nEOletJLpiDdyg41ZAaOAR168pti2P84fnw5IiM2LR
dur+A4cRvPw5HIr1rzY1e1jBhrwtT/uQA8rwciiOF6t6muWW6sKZOeF/f4xtiN6g
CNRodJBXd72yx4DkTGIL6BSRMrUnIvS40y2rwK7H3HlAF7uCrpWjHXDhvbizZrwM
5nDN0g2QvE5TTtxIb97aWXMstzvU54zkrYVkw1ayNtiIWwQpmkvhmGbOmb+JK8tB
AT8bgFrzuGoMRI9mBOvlEOXQweSG6l0GtV1WD4EWo0zxChNyuDe+UupQHeoxU9hr
GCzjbLvyu5miR7JzK/psKfshbFq98QUQ/s0A+Sz3AcuE/fz0s7/45RwBpBkdhSNH
wr/v3XPigoby8WdP7HLPw8m67N5ZyVEAfa9uqsZzwsVoAPBFq2dP7fqVKYs33TYo
6PhQ1KaUeZBIAchy+zq7189SpwdkWnUk2ZA7fbcwuAf44ZzgKoQFU6IDZqylL/QB
GZRDaFTXcQ0xAq4+dvigHJNnH9iM6pMt96Q1FPPYEL3f0Q1/x7EIbYi00bYAKxR0
Lquy2yUsfaFH/omx1azDQENOA0sjfCgx0aJw9PJpWbjvPxSRM+gnhDr7EVRj4dMR
IL9nmMu0thXZU0uw2RQESfDF9hThayaurA3v/sF5PHQFEzhWxTpdgohm05BmIWSf
uym8nLW7bQP6XXJ5ZSUdXLA9YASMzPjn43nALw62lSA/UR+wNi7LPmeQde4ok34i
iGuaMgnt8s4M2lIImR0RcboEYGsS+ke6UgvDfO908/hA0D4WGeRnwNrnPNpIr8jG
iZjb5GQftUn9yILmX5yJqc2L0OG7j8VJQDMC0RLvqwSzs8+qYD4NOTe4KwgCprh7
ODXyrrd3DMp0SCy5yRCrAuM2ObD+5TTDXEdtDPDN/laSPgKtYHWtC/xn/65YB02j
EboDuVo0+IHuvKDV+eaSbw7CDO4FIN/q+Mo4rkdj+6hgdO5JgdLmigQ8u9nlznLv
8keFkUbsHJy8Bp7FQOnvep7LFMM3yxm8GopV9PUceycUbX2plG6tEW24LDz3W3HW
ZpTfFytYWkCcgie4Ot6XoUnaXtpMFaab7aSkZtvsmhkAZA2Mlmlfy5lL4S32fuCS
VTya0KD0xBbSl+iv4bt51Fe9ogHDvpQBpbGfrVS2hSh1GvBfceyEi79ivYzgJhJ/
WnbYrAQ6Kt5B86q7rhnnzTbBfNGsdKuk3CZ077HAmP+RL+IP9i1PKGx3XpQ4Havz
JAfH6fsUWdBJKxF2sH74CdEhk1b8pggp0ssX0d/+9V97tONOTGS0u34goNlyZ+d1
HjvHj41z9JJBG437nRmUEFz3x5D9YpphqeNK0S4OWaKzcMSwVb6WJKmDZX/fgQhF
YLSmLs1ZOjrjx7wLenyXTn23ECd17J3ZB8jGRd7u4v2s8e7X5d7k/duJ4oomk1G/
MEfv2sfzlFAOryOFzwvN+WHoaY0XLIqW6MGEokrfwVOYAHe9xVdUEDp5MhnirnRi
MFLsTdChyBpG1ycJRIQuIAomzOOQO/561QKKbZExjm9ldw28mzHYbqTkSSbIy6YZ
pmg7e99LUydkjTe3hs4GOZdY3otJ3CyKyWKat251NGr9coI0QjJraIHTPi1NrLn6
mRSARAWzXSezcZBJQ2IpJ+w45Y5nuSMrKEh+1sxcrd4bJqaZq8kdjoJqdTyYqN1a
XF5EYlptTYu02EZloFGSX/DwHOvnDHZE2m97zlA2oHxTvFK40ymEdVg9sr3zMawN
G+3t0BKtzl9YROciTYaEqh5Z+asudmEaafR2N9Qc6aQ5jFUznyGy2uzc9BqgGJMB
Hr/wdDS6CgQ7WrxyDmUCWNDv1szuaROZMBq8r+P7QISMeKsR9tYUg9JonZzx5Vud
L+C8mw1zUGgvBGX78hNrZlKfzF50rSFRaKAiUt4aHxnOiyU98oViqVkW3R7m+dfb
cdp8YAEUbqyDMDcxfgfyUAxfeO8HSsO2SEzCGN4S0Giz5wZTar2e7GPmvBN+EA9a
T3zKT+CU+i5sLsbQSxF2D380auV15JTDeufeUOZ/l1Pf5O8gIWJg3WSJ5HGQs8I5
Z6JBiMSlIqgQagFeDXrTnETsUluqpStfLJvtGf3TMvM2ZW4o0dOeGBXTiFh1V8CE
HF5j/a5KAVPkWa1GNphHZ/pQSCGCE/zBNcpY1scSIOR0A37/xnYtflcv3wQgYZzO
sdE3gGbMOs0MvoB9mLjk/Maw+5/NmUrDBHFgTqGVyhHaZ7oMG73GlyLXhaSVHinq
ihTBb8R2BYZv2qpuebRWk9Br2t06byKMN0zl+IBqWE8ais3dofmli0BKs81fBUMl
WEXKpQSRkJLiUux4bZf10z5fDGX6A4gN8QKnhlmL25S9vYHlIn3WGTOFaR+oX39L
RpPGzjpBdMG1KSfu8BfFBGQ3rFdZTE2C0pc13JzF93udkIQ8CEdWtPxvouQLoFM7
LXJq37uf/Jrz7LyO95e6+lIFF8iSVX8ZW5t4v+o7J0qNi8JnlmGmnohTI8rqXXB/
XojsauAoTWxPnI0ocqO/hWXfiwUf/ACTVASEcEmQmjQGlU1YPZYR3kc/YkpGbGDg
FATGG+udP+3y/EF8RhsOck15XJDlyqKlrvDwTmJuij5buuDCZl3Uyz4IhslrMQsq
IqIBR0BVg3rIV/NlrAhQGy3R5x1Y19A/qNdeJYU5OG26YDzsJBj1tkQCQMV1UDtY
XEBJUwWxRfUycXQcTrQr1oGwqpUhWTB4wZmrRDbh+zx2lUFnHzSkXqdjRe/QqcKo
YW685DgsnqCMVnnrM0L8ynDdE18khy5cKT2BfC88RFzPMZhup/j+PaIveubnU/EL
7yAF6Mhu8tIYIRZnZospAiMg+Ih9NbAfMS2rzVMY4uS6PH5BUHC9dHhm5qOIJb1m
sF2Tyr3whFhcouU3bQ/HgB3f3WMtyZjcxOkDtl1YVRjjQz0w1lLqKVYDbFZ5QDwA
WjhwyDAchEVmSmsBJTVobI3Y8A8sUUfGhkknIZAnBTcIVFFB87nQjiwvbahDnT0a
CTNWdvXSDMof+6dIzZkTF9DqV9iLqZ/Ja3E3+rktzNnmWo5I92Hws2r8JrygMX+U
FdgBi+rAUPO8sc6CqYXy0jRUAzpuP7+KV0RX5/CkPUT+u9iQiFOXIkF0N86jbrfM
sNYYPEAJf62SHNO+gOPXmOCo0PpqaAUMpoy7cdk/39RxYSbPUioVm9BGpRUUo9GW
WyluGuepvxWdtIlAmiZh1LD6LXotisiAHom0H0e92TBJ9CnnUOjQldL4TsTQPbw5
w6JrWw6F91ZwgFwqRu9R/IzqLo3pT/e2qpi8fG0glNfgzeZBfixoxUiHQnNc6NqL
AyyVjyb608CG+D+UnBOU6x5iMObfEMUJhJgvMuwfh13lWLSAhdmPvi53AQqyp66C
sXg51Bkdaaz5frj/pZwBTFZi299jnVmEmYKVHkjVRpus/BnZZrvOWE2Z7TcCC/HH
BSnihEdQGufUGYKnV0IyZxojhyGuZJhXV9X26OiJeDSLcpCyGeFnW/2qec+aVJ1V
h5NdF4z9i3RQa0K3vtv/TNQc5QbC7+Y3k8N69hgAnifiLirSEZKmQHC0Plxs9vwL
pqMy2QhX//o7Qf4JJprF2r+7KbQk00/BJ632esgsa8jE8JbzraHAe37tf9D3tu1i
v/EESwuNSNFZBMx9vskZsxOGuXLX7ZmSzmVp2DfF/fFqByEEiHLeVHRKRulwgalf
MmdlDsQzRvjBEB+I3CWkBfm/I/4Wuq+sQjuRqKpW757mgoi3aAn3ywVR3v3owI92
V0X5i7V+sPdmNN0TBwMLRL9Xo9IJuU+y2y/XkJecFm3MPZJ2S5yGCODGqL4AWb/U
0Kj4AspMK2JCdh8UJTbMl+Us0kJITgb6waX7dl+M/1cF9DU/n4F/vvr8wT1dIhJY
aOC9BWXexWneyhDbdpFsDjo4zSdkgfQcsnJTKbm5Z3ZOQtceR+eVMy+U7EU2sLP7
pSKZ3H/YuzKR5GLe6vzD/koCHedXW9SoAgefGCbFkoKMkSw0NQYfgp5wDeE3F7Jq
/HCNfmqGAz0oripnXRc/f4gDXqEj7tIe1X40sllpYDEUZh+TW8mPJZNb3gjzozT6
zicw1Y7HA4oR8r4VTXFVb/82okT0US326dYfJtn6+H5gY1vnz6tmlZwlg10Qpzih
z3kNpLwuITwEvtR2m6mnp5QZR3HHvCZAZZJSwLuckJVKskpR7p6gTwPyzG+AvfUL
2YgERt+fd6SVpvfehcAgQ/zxURMkdju1lxrPCSIexPHEM4+vKbY+8QB6f4E9QhPl
zRAdb3CFXBG36u22hWLuKPcpXktUcFnBqnaHOksdYwfkz+71CzXP7E/Wt1fVtE1R
4d/ALC5UKne+L1ofRbgg+uabJnVuDLHCZgxhGv9C7OPGK4WYThEn0wTqxsZYtzXQ
jG6ieFlgYz57Oa1rxbKuHrnf3qj1pSZTaH+QT/R8a5GlaWg9mKdjSkAnlDc+0v/h
ENm4NrmoiAKz6aTxsZPB3oVI0whnPJ8uzjERokewM2A37pPanlBHgb0EM4vdWsc7
VYMx+Ln/GSRlUfD6UlZuRTy+YWu9H7Z4Wseh4xm1XvCUOxN4o8PagfIVR+Kn2Smq
+7xIL8RrJXKUmlqrI4H3y64SoNTwH8+vo5/+HBAflnIAVHEPf2yX1hD+f1G+l/Ug
KxBzXq/bh8vuNoRilxxWvNHwkSW/IH0b7Nfyc0sDxgDq5z5IJUWP+aLEImOHvJsG
cg8QgYH3deunT95Js0dCm3RnzzF2k8WFWkwasN/IgpZSaukQlE/m4ceKk/08curJ
/W8Y5jU6yCn4bJ5YQ2s/0miBcM4G5J1XGSyBnM2DpbxMDhUKDPONVFuItjFwRgWS
ToA8cs4jE4azJRMpAWKyTOZGdNK043+IPP0SioqUMcYQZZqbrAdKReKSV7nwi488
Jtao+7kLTNAT0gOG5HmcmOcA+ehG7pEMhOZo1L2uLquq1dO5V2Ydcrh+N6MskEd4
IGtyhALcZQ8dYMwL/fXqsbze0qPRE+zOTWAwxeKDKpsLv56tx79o5s+cyKe86P7w
k7T3qZ1JNZu7iV/58izFLfr8ltfsaEi9HR3iViKxvkZmqJ3PYTiYLMPPb8v82bP6
6XO060xgt+z3Um3oDVemBd0dixsOQSbes13DvDouiEsivtREGuCidO8UVuoQtNyr
gg7teH0hTNk2mxPa8ft5fdOjcZ3gZ04c1qoyamXg5C2lxN+g3LCRVbZZoNxEZqOZ
W/4QTTZdBAe8j8nRi42Uek2hCJFE/DoNe6FJDREGYt0/iMHlmfwQCo9HsXLDVMIW
fjrgRbdCle45XUdJnkpqzpLZGDNySDlUEi8XVbkzaHc4uiAyZo0hRRzV0s9sDiAD
aMdzNqsZucySq9+/auASunsC6fEjpM/nvyHWG0XzgaAPUDhgMh0XMVL89V5rdqlK
HrJ0rQSNqmXZ8B9ry0OKhCtWePIi4joGEZt6AKUB4rm/jXAqPhyNcOTcQ1Iq84PS
QvldiIT2qrKscou1n+hPJcpPqmvveqKAhbrcEVIFDrQ8c6XuEetG1uy5mLQNJde+
wf+ScO5f0+SXDnARNi2znHy9gyBc3EavqeaTLKsh74KJF2G1lJqINJQysT8b+CIe
u0X0w0kDojGSiBnUxSIne0NM/5vLniMq22sWScSdF9zqCKmouWXAiaJUgvs9ML5Y
0CbcOpuQ1hAMA4F4E6xBN+omrrxvKbe17D5Q2cZZkBs8KYGCYaxfTDvAd14/3JE3
1SyvnRWCnW9u3VuQq4opsC9/9QpnDjTgvD+ie0h6/mTYnGG3yOXVw/FJa1Vx+APd
wihqI5sXAJinCZSyYUghjMBz3KNX1ce4llg0nndTMkDjTC5HTXqBx/Ip5y4aKbWE
UL5VgGU/jFoQSGxQ/gmXpwSVb29ng1PfwDlcyTGhMyQ0khRrYPF1pCyb7LnC2Vhv
Gv1dq9gl17OfmCzX6rjL2CvZNOwLUHu63/tmCEjfdeJKRDdWWnq5gSL5pCLvT3cL
VWSuITXnP1AeaEMYri9yc8+z3rkjUKY/IlNoMnpF9WMjYpEYRCvuZnFOsvpFGJhm
sUrUMbKoI6WS2SqbT5gN1xMC7IR5wYRTpkUDy7TIvVgPBYbUYqTx6Q/gumOhX8+d
2blLmSPgl8x3ECLnZqDmg1KVNUSjzkDV0ovVC59jf0LpfDWjzjJZtT0gbsskJVz1
qppZoJ5JTPqk0eWE3KVT5+TCpYZUdywXmwg8P3zWU3RmY8jdERVVe46YJx1mS+Yp
ry/wvm5Annm963CtwOUrN1kYQecgYPIe0YdgcBw5jdC6FjiuhVzozdSbbf57lGLc
rfQ3Q9E14Sb8ZfD/e/Jan4iRzqoWylbSSMSuhIuS0EoaM5aitRDr9qMl7ktnAUXP
k1MLm5Q3d4c78GWmNxLzQSyHnCVkkfcNtiaxyPZ4WkMPh0dYdH6Fm9Tgi0HadKvy
jv2fYniedW9cCONX+AWoA3vrCiyh6m1iDTHohUdmnG3eQIi63qbvWUEITCEjXFxD
fzKeofhSjGUXgZ1clUsbsBtXpsebtK0fIO9UVhphKnz93ttuL9zkXgS7+OFk7gev
CaUT/Gf2DnW6Qp2g0cR+KAEBP9RFbO03Yzf8xE9sAraAgT1ZFbGN6so+8X3w5ABQ
UK33MLCLyzCgUi8rCc+oyKJ0lXyXG5XKoFcfw1UREp923K+KTehi/rEjrMPAbFaP
omnjjmBAwopVDPNFXiAdxZIJDidS6fXmUfzzcO6wQQqcZGywy1NzLZhU255V0EaP
a346Yy12XuyButJiD5rP26ofVxdKg/SNKcVki2RLDLioUa8/e02lBJpOSu8sdtNZ
Osqo2GR9e4lAmjLSodeydxANIp79PtJbM/22931u3Lp13d8ewrWGwq9ikTiv+5d/
FX/HsFonOZ77xrOt1z0IVvw0L1AbC9tpKlxKsoOwMmmfK+nmh9hfXJAHm/yN73xo
u0Tt6+5DSirDsX/ABIsHewRtaiI2tNQ7tHZpwsC+V1MF7eBR0S8fJV4khfwnpdrq
VdoY+iBpRVwgUmtzSigk/vrvXSVbpugI6F2FY3k6xZ47m8CIzJXqWqE0IjWdJSrw
0DBXle9/20AM+e59cVYn9gmx1WC2r3QfFTrcUjb+Tc6Cimoo7HMtCFu2dI5BGGye
VVXwm1F6C4D+qXX0CaPIRxV9gC6FtIUipclH81Af4cQMHrXk5VRY6vemvvqLHXf6
8e6f8v9J3bwb6kIbZgdesjejuOUzJ38PJ+cakczaI3KsMUQ/vhR4J5vqJ0vPFdV0
ZlRILuoxPBCqqtTrc1y/Sm249V/suufP6LzBUVtnfMeIRyDZ4qwBlgzT/MZdNDnS
o7k9ir3Ov4uTXkV32g+T9rcjxtGt+Jmg6jOvSOWxzMBkzOg4VRdQjogxKlFHkzh6
SyyBZSqKym3KvvjPP/NEclT/FRCCAJDTpP/XyHHu+5P5F7MlT8PBWEpT/bwLxWyG
cbXmhu5hW8jv9VtSCpmo/qea5hYq5rqFxVWnuHnaQMxdO/LbxcrGC27uN1tt0Kdb
dL4oOpOlHeI6hUrLWSTDXyM3kFEWA7Lzqh0PUOpYOcKup3IbfPMBn0aDkHjIVbz9
McbCl1pcWPR9ugk6FNlZeT83oysdk2Hi9WpCqSm331DXWxtOd1Hb7BlY22N4F82K
gcoZ7NKKJ3TE62yenfTx6IgJyFUbD1VZlClXubonramtuaBk/3Tpe0ySy2XsR152
Q9TNiLsYhemQWvnR4QvBiJZQxvqOUke6RxdTHgmxJdek5Rgtzdbztfv5z2LlNwGi
Vcf+sJZCstM55LYIW75ATnSUCmo/4VbnEueKzEM1427ykM5ZQQp7fbPQfovy2dJt
Phou1YcRp4xBWiS016Ml8H+3yFWHti6WwG5T3SCeX2+1WJbo63+MotnebPUak4mE
W2oOQD22qsblju2MfpwQmvVEZzqsk7Fp9w/e1r36O3NeRWsNAQsG2b+sPxdA/9mm
rXlss0qvMtbQ3/OxDnPRJd7UV/7JmGiagKgu+0e6m3f/7jXV+aCo1QgEmy/U68dy
lt3GBP67IhkAw5QyGmJhn0RvyRgSfpvHmKnl+PZ1QG80IYbxifyi65JF4EkPxiP5
XHjduAnTKIWDPe1lRlmrBkoLSbnD4ENGVH4Ay1xW2UFe8h6LFjJhm5m9VKpk7Xo5
ZM0ix7l1lTG4i1luaFpB6SG9Mor7BuOsrgsWHhbYIZbWE4/aqR4+Hs19Uel/abDG
MU5awIxYR1wh3j2p9wivbo37sEonfJhGQYvsLxT09Yx0+9WqWvBgt/cGB5usfUxb
4DDSj2X2imNpOmtiLnpVuGVgwsFOamCTNSI4jAVOk5NkWvxHMQB0XffrNKu9hcCg
ARjUHMEwsKMT66/JTAjfznw2QXoFof6DZou0C2NLlb/J2KEx8WXdghLzrln4Z6Zx
pB4Kv0kavuvzYbuhc2BdEw0BEanwxIhoIthZD4TEi7v2RKoUkADmTEsYt6AVtavB
1MljWAe78hdoNKQA/Rtyl3TLtapK2hozQyTaudTFkMksagASq9g32EjbIcnpq8pn
1Rwl0bq81hodqjms+W8ABEGzGJdHhQLoW2coEi35s4PSi8ABUenV8GSnrCNq0XIT
lc+1li+Sm2buFTVUHF9T4m0nwARq8VTei2bJtkoOekDraKT+gDdQM8FA56eJROsM
DR0oNuIeXHbnYuV1rXEfEVTbWvgxKdp/PWCh2RZgmr3Vaj6Zl/p/g8sqQ7/u/AXZ
XnetSQjoBIJCsASEwTTb9JNHEa6wGW7FxbSJdo2YEXAKSan5PJLE3jgeobXKkSqD
PJpoOvqC3/Lvy7QbmDN6lvoCE+q2ummKI5WYKLGuyHEOMwE8/fwBFlR13l+NsxOk
X/ThAaVfvvOf3ZwROZl1xmKkK5yfkIdQXFqwjqz+relBIKmVEOnOAEySkoxBH8vQ
mbZzGr8AwmyiVW08DnPh8S8v76dHC7B5szhTEyXZ7qB18wknxT4AEGbjWI+jEC3k
Nj1zcWakOYXVGrpXo4uaA8DPs+t/fIel0yd9AqYJDcnqulEGnZ3A3vWW5lbNLx2u
uNbl0IxhwtkiF5uPgwlp2k+gNFWzhshUTiKmGKNeoo3aQMQqQjAcWarQJXxEYKXN
jekp9dSfrJaRvbjnl0z5PaqW0FJAIyf9FAtuzUMLLydv94XwZ4LdRqUU41E8KRB2
C6hsZd5xqILmFoCfJkGosR2AJ3JFutaBNwR6C5zy1G+xEi5H9K0JgsxAFTlfQrGP
jWO8MqI0YNfE/0aXI3oah+M1lndzA6y/6uVJAxjHxo/DKn67VNbe4DTjQRToU2B1
kdKFO0mkAlELlAGwuizlv6WK56TyHWzzfnSNLUO0ai2VHlhUWZqKInx1GcotdUdj
B4o0JcmopODYTEUu8CkDZAW+sh8beL16DGNi4PGz5MFUJvolhYAavobKxdxj7PVy
U7SpiAfPap24OZkLWtZhnOLoqV4NEjILSqDhw/7f3J8PBQ3s15pHZ0tQeb5Cx87D
+olj9reMyirIc3/XPKsd7Kw4WpSJykX6TzuMNwU7Gva0AoRTDnk3Tr77U4itc/YR
X9SuYzzujdrKCHPfaKfCXZzDlFvzQczKOVAL4Q3dc4enFHQfDCTBv+rIXO1O4dSc
7uBILy6q7XRTwdjK1YgNQTqITbwAUbsVaZex9zeLSORs4eMzdhS+5GoJwom7q1kD
5wjsg7j4i9m4Wwd5jRNVpAKoUUp+IzJgUqY3mwE3iHB94FByzQKzy83sgBAoZvaZ
tNIcO0rHh0TObjMbWykfrPliASLA6nRWToFiX4CBkxkkZsTJKUM1/v4dFfz0dG6w
7GM0NmCMdJbq8iAEg0ZCYbbpInEipnToS5sDY1iH9YqUpP5mY6UovgMke4jkChOq
ynocyc9Rr/SxppapopNQW7BtbI7y7O2VFj6FMNJZhhc5oi5AtMWjeK/yrABxadFi
QzdPBATSTyDih0nhsoO61wB4r8hNBF+mmMdpIVLUSxft6k7lU1F4v2ItpBYFDAiC
+GQTNGXYJlMMRSgGNb5gfOMZqncQ8ctqQ8p8bZ+lNVNuh5jNjmkcgSpSv/7IKwEm
VzfCc5dHByNPdrNzUSqInrNZbYWVppdHjkXn/YnYRZCQ7jTi7NTCBDktS3i6EBs5
6lk4LZZ92tDuKGLqck//DkejjjLnLExgkjKbCFeVFS0xDyWCsqJTA3poWmx+ykj2
v1ATcuoetoxSNKCeF4n3hqv93n4qqUxsdkJhbF82MIlcYYouREHcXY2KU6LYOeTi
0aVxCizW/csdj6Z3YsbVGL8uDrrPnv2ra9tazyHp/DbnIgE6DtW/j7ktaGM0+vKj
8v2J/ARr7C60D8Al1D3dxfEfDiCUVXjrly0cpdLFbH87b+SUb9FcRWCfUpIQAmh9
VoXRaXSMHN3iXQJ5j9ryPeDo6bvsCeFGOYyhTTSHGc+EN1m6/AC2HLtNqWhZTYIA
vHaH6PxQHdYjH3+8g0kQxZ5nPR9G2ZEPExqanVIV4EH0pRg/m8VKW2HjJFcm+5nv
5L1BKkdz4v1S/rRujt64HXufxs3x6A/eh20H9q+mns2iaRLrQc79trmPBUOHmUoV
9cCEY06grDw6u6ep08LN0YSuUOQioRC0uKTqr+ErcN5wqURJXeDmm38PGiMbhX/Z
1Yzz15fKx1xq+eqmGgpeSgDLPYBhEXDU9srzvyUqUvqSiYwrVj9kzol2xmY7l8OR
nv1jdO1PVUtGFFFuJcZAQoxkzomx6TozYOxt55Y02R3XdF3R+TAKNSz0pB4pvrno
lyVMK9ppbDy/opmm+dEX/g2rcoNaK/ovfr4eiiCwrRwG+qUCJrPZLyjE4C9gLRVH
vcg+yBVPo8nZ7Gq8rdVtMaqW3QFuxlsXP7qt7y7OGHnssq63Kha5oVGp1EtzzJ1W
j2uQJzCsL8EshdRye6fG8pDM/73VAGhyjHxJdhPjD8qnStvGZvmMQjyFKyPc5yBs
Y3sw5HxCL2RkJRbvO4lmfnnG1NiQxTkKw3uSEu8sdOyKN25sZSfeKkrkbtj+fM6O
Z7flWfjd14Rj4D3VxGynwbTuyH128xOVu6CXl0r4T7HFCtWeGTSsTVkX8G4X3IdY
BNC09ZlQNm1upf3ShNdWdp+cfsD7ISIpeUS36lb3bqJTq4NvDqI2EYY2JaiYh7eq
3ow6ec8oxK0Bi90THHLUELBAYQ9+jR3Lm3PfYy08FAHSrIqgSkVffdX7MHLW/ZAo
6XlIj/HysNTQecHG2TX+kHoNZab5hG4BRYeLkfulJL795tLAtpiK/Q9LFX1/FZ1a
0qItUlqVgcrfcKfkNNUnb3TjG9emaFMji8v6ex1s1ghlfyDNzpMqWzfgmi7aebo6
sk2mho5XrTKe9PPyJY8ty1BEUmMp7LjKpnUo31wnRceC3xJ+aJ5kwC3SIm/vmI0K
V4RW8VaBVXJwKNeP0VZAZje+FIFb9VvEWy4O0pQ72jUQB4VE7jhpkKhc0CLnUKBP
6AGZZZAOYwkehYwcy7Rn1o+qhfMS8FRrMkjgid9PpXDkCHlr5pBClJmR6xdnajFl
fq8u6+nFhYQ2Fll7gQ2RVf/l0h+l9JXVchlVwd/TdSyc9Sj20NSddFe9SGPhi2NM
v1K8a+fiCRYbbDIpUQxsBH3vlFRBnWGP/o18fjm1PCA6rlUZDLTSx2204x1RM8Ax
jRkgrkd6ER7RI2uX8tWHEBJe2DGyk4u7eb7LopoAE72nAGOTg8N56sFXvP19/QRr
eoC9HqXQhawRzQBlxnBWKBmQjaReJHdEDL4KbEgDsOmVB6WBP4dfsfT2G0o6u5Ia
aKvIQTnW+rCk4ReYJxCNtWri5RXeFTHa7KINdtpHpEqIv1aXi/Hqwa5QcntpUYBK
kGDQgmpJjnvxGtkaV5u+kKACiGnL80gDK/Dk3AOI09avvjEAQOjiS0nlVti7MslL
cKl3PzZEmjlCF1BQkBt9UWBh2znV3xtSEBKoi2iI3UlLhYNlDBvEuVa2Y3Ng67uE
Rcpt5tl5/QqJqGlJ7w6HVcY4sntCXUmvqnYWhbLkBHoXK0DTz08lyPbyvhy8rZZ1
OV5LirO4tlRbXl637zgas4kOFI0GSdsuP3+UGem5i4UuqjmxGLTLkFVSGm+6KpD3
SYMYX2IkKGedIDsGfGN2+YexYV1vnGxV1Nkx2/pJfLgTk8mzSfACUQqHKUOklbOZ
LR6kpD/ExC6aVhM3aTaY4h7chWd6K3K9W0R1djGrOYNRk8fl5IRJSa+QgUj4LM5W
vRc0kxg0enot+yPaVm/xzE7xRZAWcPcQAMTQ7hocffM2PL4int0QSJe36RRmM1aW
2lafL/nmaKJaRaLwDZqYYldqtiT+5Ug7rBxYa5axgFsNYkJF8rXWfMSmyaI5pwO2
xWTxR6sxvbWG3R5WWrR9w/fjNOL9R2lmgaxT8/q6kqYBfIljUxpmbI/RAQpdW8kh
XaWvob4/yl8GzYtARePb1xvoqq/FUSWyuaKK+AaRmjSEw4py4iV9wZatBaJDmDKX
/DWFKASTKrrmeWHdXqCd7gpop1rAh1SJXnN7egwu3fV3ekjwIFjktUL0ObaycKeu
8yEk6tzDEMc6iZ1xdNDEamVyt6S1WsCb93l3nSroef2jIoeepaLvLeDVHrSDhSCt
Ww1D+3Xb1l4MJFPX070WGcPIFRSHqozOGg15G7LY/nGvvbJ0zeVQWZu22ua3NgPF
hz/SgRBa7ng1+PoAcnMxDDew1HSVqPUJBwI9cneyoS13vIUpOBymSR3/QxacgwAD
RWpZ+Ky9/kRL0t59zclDYIvH88ZbJM1Xeb8RDlmkqVUyKENxNUOlm8CdB7ZqpjAd
IgiZUUftvdaULMvKCv+NKJaBtGZ35MrISb5/ew0Vw5eWYtpDigMTPBpHcVxo3uWP
2+b+AOTFTpMKSvuVsv7ZRzMSguMlD8CwXzx9vziLjxSj19QZqmLGXHfieAFNc41z
mHV+FtbKQrPlNU2QRUK1h7rzaCo4KHV1X/HhchOkvq3PIQjp+zoLGD2d5ZLkv77x
+rBEElDHpQ2L30H06Gavv6z+peGRLIQvS8rFXu1oQYLnLu7VcdFlFoVs/LZE1cz0
a+s3/7+kF0TokXrIk1F8yTNvWkhOo/+5IzNwhw3VUAMsTU5PH4sRkoLb/mFMiENa
pko4LslU3x0bo9MuTZkQ+EG9IeOAyxK9JKApNJ+jNXwi2uXaLL6pZ+vXUYPQ8M8J
y+8avkY/EFuah9j++GD5EY+NxQjnLbhhU8OUt/yy00RpWiW1hcoc5irSucz/3E9z
02xYUdjQFhdEBc9nwHTbgx0hYeZ566lxAaxiI4z84t5NJmdm0aaFi5MCFMeMRrAJ
6vcEEZqEAPIzRdGYezt3PtmpAgS7rB6P1WO7ulpcEqL0qh3Wq7zehx/vpM6KIfKm
OEaXdZu/DXBUq49zDhvy/I+mgaFRDVXqiyTT9jasGEBdXhsVb9kM5+pb6zDngvw6
3XNQJkU4fAbEW9o9G+A3SZg9L/A+54jcT482ApdOB4I3AbTI8i/eDbXFsKhoK2ex
WWW2sKi+ci4ZOuWjRbxCyYK0i2nRyfJUfEicFswTaPBofRiu1LpaFF9WM/FUC4Ru
iAxi5eXqyqBiQdrA2npCFM+clAh9zczh/zWSJBR8UJ25xv0ssrghzVLrxaLjSodG
0fuPuKXRIqYIhcYfp5uZsKdk07fkE7UtORG2/NpmH5FTrV+lAWSWvUIz1xYHJc7s
2Ql17vwUtDpyRAY8CNiMdnQ4osUgWC8vZKgcny/8pNbpYvPAn0+uKcWxD+tIxPck
K+ClgJVciEc3NOf4Klv/RflV8sIkNVVY1R6wMLKL3TtlD12SgQ/loP+QrZo5h/UL
Dy7lEbXPgyDVaQm5DiLp6NbLwYpAxJWC3PyUK2eKu27KwVVOXUQcAv5p7crUh19C
9OaiYRefk4dxsVnvNggG7UDJV3f0gW2sPu99iq4Ov3633qphK85mro1fQ3kpltvE
2sJoUECQG2CQnXZwlhHGKQu1mb2HKV6h3m4L4vVRlg4y9T14BqqF1g2YYZNlFoJH
AgBl5gujg+40ulDZRew24YJt+X8DFEqRGJPvSt0PRux99NUcSELU+WD1MBQ5EqMG
40lbxDP1E64wPpTMdS+DGQ6SHKQjMNGfMFJheQc4RjCoXrSBk9WtGBlBJedT3CDF
rwb8Iyl7HjBX+ty6+3bUVWAkkolKd8ExJT0UAMjGsprlikQyPGBDNXsMagxIhLBi
3uTgqcSA+JsunKYgXDqHTXsemw3Bybxpp7w6Z8ieImnNS0RpZuFgnUju/+Sp41sH
A0Z3iDuogEWz758QKlGly9aTYboKi+AVvmy/zzsOFO4XGCfsrL6i5CYhEctLDzPM
hPfgsylivj05MqTwwmP8OQRgHgl8XRbPiK2O1YDS3dmKmWD8sVlRa57Kugl5DoSh
7IVdzAl4Nhr18HAtTH/TrE4dgZZ/jptA90A5L3HASIIetqhSJ+42Bk0aW9BNrSKw
JINSgbG2CsRLvZPHnDafOiN4bnagbK7Wdkam+OZMrhAvZTbBh5HJwr2OgtxFt8Rl
Ag1VwBUfNNJxvt1LCz9Y6A2f0M7f7eHvUNkAm2fHdeOuCRjcMj+yis9NDvmmkDon
VsO67k/rq7VZ4J57o80lJybTZXhRnONXDvppH0fazWnhem/5VPTDmvwGHMIqurpV
shZnvdfJAUg5becuiqnOMGg4+vCnae5GocSva2IIVCDrksvm5mWmJqLj1cvL7P4k
qM2w475ATg6SVz3SavTIpkT2ZUnK19Y7GDYrs8X7jtnv1x0BfQqsW/VZqNv4HpWc
q2v6rWp6TTMoysDZIr0FrzTLN3ptkw3ygbTF5qzFzywzSQNJYWSh1H66/Sz4xjGJ
wZqQDrkSMDXyqub83utDcWsday7W+xo37jq3jXFOpy8p4ZPTLu2XR9PfZQn2ItNW
X8DsqRUEGZaznS98t/QGDIpe3sEtJMYb7QAwKF7Q9dK/gebS9lfHFfbSMrCdbFme
rf90HjdM4iZpj4uBAAjC2WP6mRs6ZmD3GV1cm2PegrEzweCw4LYG6nX0oNlzwk05
ZoixC8kMQV022Hkr5D37KVhucBcjt4gcxs++gBht7XnWj6M6oPNkllBW+7SOqfEg
4YHst9X4Xe96uiPnDyoAFPSL//HCciT+jefJ7Onn5V7d4K13n3SRXLfzoYcLVO5Z
vjHNHonlPizun/3PWW+Eao/gcQf3949nfBOC9QzsW3bzJW3DLJitdIrmmbIaMDwR
KfCNiJgfI4roRTYn5ixPi5x/VLSd0UFW01wC+Pl34lu02gVaPBPtJHf9KxiBqG7K
VawcCzWuWF3HDnWwxTYtzdM0Jw7uJQdZv1nmBB0ETY9HaZIWJ3ei2CqVUGbpdNjQ
w+7jlQaBQ83RMbGdVHW5VDqYnSkYZvLtVg2vQky0PelTpmTbpCTQkPNYVt5Dce3l
4KiGDQnGA0VSdzw/jh5lABx8m36WIW1CZ6jciIZ6S5zfnJe6xTzloo3jWwgXpFtP
z7D4bJP+OLTabHAl3+Aft+v19cFpT7a0c2xQ/jfcLmVPRk8lyuSMbbondQwz8JS2
5+6qxCL98qDgiHi6LDL5PjEIC627K2VX5LZuORa/Sz9fLDzBSgpceHoedUR/mJP2
acrA6CXcsSPP8lZU+rZdY0D0ew3M6srkhXsWqQ9J9XDDM7DrVHthNVQr/pfz3k1F
FWprnSbUJmdB8WVN+aD6SaFKH3RxH8oUWpAqqz0xwNSIP1mXULk+H172JhDGKUpu
LJvGKszCFcMwpRAPGzc6+ggnVkWYt4jpFPG9sM12TOZpm1Kegf25Yns0EgjVyUco
8+bToGLyWu5g+F9FW5Yt6krfUZHYc9ybsTgTxK9pooTpNpcbAW4c5PwhX/rM8PEK
zv/7BfzuimZfWWJkexEqFcBvSbT2zt52Pp+bDFvFAE0sVj2h4VWleTkfLjywlJMY
Dwcud/EiS1clOQLW2MK1bxLVYqNubRHGslA2CGRW1pHahMX+OC2tQ9r+3ZrG2HRI
29Ie7qnILo1bt7wB+O/+koQ9O3Wa9Cexl6kAiOFjg6NypWxEQ30AxOp+205aDZXN
mnHWAl68GfqQEHC8GhwBKNHJRjG2Mz8LMc41oIs5u86FyklGuK2ysFKBlN0vUuI0
LE3351o4K8HLMxXcx4sTClAK5J4mbRUb0ezcmj09qFQjnHsZgykFPBXjDMbNDTWF
LUiEanhicZcKDy3GKOurHzOZFH4qBdw5mKWXl6LkRH4KoEKFKKPm83M7ISUrsqmx
TcDruo+WNMjDKiAWpAlkKl8RmEHfVZ7tDn9hioRP7BBHy5V3xoRqK/NQMHK+m0Oa
g/RS0Qj+6BKdw8nMHwpv1449lONAn7WvwYuIRZFlKQFOraw/MRgtyt89f2KrzYvy
x3wGPjo5uteywcmiwpBhJx9ltpAPqObi7sesrE1m/QNHnhCzK/8vPHu5QOMpMvx2
wG2Uh0QYV8prlsx/gLIKXP+VKZBZOpNeu8jfI2IZvez0QyRSSFWXhxPc2/wmgmel
phh6kz/JrMqTUnKAvXexlFOki8pGc/pFmNSWyyJVE1+EB3lXrlpqAgIiNQOV8vI4
8xllEQzg17uDzExtQ73PGGg5cwvbg4RRXmSa4WDaZJpOeXNvr8DGnkYnP1GeNxXh
JCcBO7CIUYX2n6l1QQnvE8rt2ba2y/PCxl6YFdULPZE85Q5bwDy53bnDmIt3JyKp
wPqhloq8iaM7VswqQZ0cDnLsvGxpM2chQ1r+wDeh3xgydYzChrv0s8FMRJ6Boj1k
7jvYkZpfz2c3+X+tGrmSmPOleNnfqmq8r/b4jXGScU9xhqlu3FVWihKIUgFmPHvQ
XoQTg57RuZadTQd9H/5zsfjL1cjVVa6SJal43d9DnQHilJa+9wge3R1id7GrKFVb
z9DhjBXZjUJq84ZTGWaizHPF1JZa04XUPYEkOUXBKWnDlvzzexcKSr4NFHagzQWp
NOZ3rPZRIQWtIyP7rGFA+Ym+0LIRgR5WHjS6Emd+DJGl7ywizByraljQJEfY8Tdk
cl48lZ91qjaBpU4+cztcw7QR1hyCbMxIHzeAaXIv7xN7cUl8jX2R5fU85fE2qEhh
ycgtIlhw5DECgB3aubg7taEI7nL1ZOldveX7W9nh9ERmTy5Z3Q8jv+KuzG3vJbRt
P4ySu2WE/KsqMc8RNJr2TNBYJIYQ++wTOOJ2wBJUAQR0yCaFeigLDpayiJ9gy7Wk
v8N4XId0h92pk4oU+2JMxC1Fn8zln6kgJWafGYiWEbf+29wQunxqo8k57PnRgM9X
OmRrtLcaxYyMzmqM4oevqLBbyXQdxQRLQQKHJvpRB0Ou3OBgzktZf/K5hgBEVTiw
StRUj4STPy9tjaXpkZv6sfiyoPbwg4DOHBJFIYd+8xaTGloDbTw1bY3f3fKrcyZ6
eHCzlS0U3BsdAWASKwoD+Al8mpx6ym7vCQ9lrV7BDP4xXgucpPzNRF1+LFFo3gNY
0j0Df5v4hFnLefh046Dh1s8sAgBdhsx0hMn4b/qJDplbv5lDko+QrBJpBN4ir9wm
IErgEAHteKalwh9XhFtCfK3Pv+HWFUpqaZWUTvAIHb2T6bxtzAevFzVNXHoLnINp
6PFl7MhV642s3daMPekRPvwCmFSzY8yYNuf0lKFlnL9zn4UcoySd3vsk8/Vb3avL
DOkGXpSqv113r9w1umzxbtVjpwGQwPrlnP8tiLQ48pg6xpp+skIh8VQWu0E36zJr
mwfhmGvyxYMrhR/dLODNMHvJ0yyh84FKiwRR6/q6CELW8WoDQlAbyBBotddmXYCQ
8P0y2a+z/J79CmN+bkHURo6HlbmYGZCtKPrnE0vgUQQfKg/FBJfCnzvnQ1Xijpqv
+mmt9QogVm/FEXQPXIPm+2eXnncM+ZIhIICpSmgX6/hG0iSuGGjoLHSoopGTOMUy
qe1vXbAQszzC3VK1f7BuclWBxI+R3Kf+H1DSMUqhcpXcJRJuphacZMI/SWSmuyjw
o5CqOmW/iTOM9C9Sr7bcQ3yBxuMb2mdBpqrYcnSZb1avrREwObhGhewW/1Mb7as7
XXMr5LALWlMOyjaS+WiMUgn3+joHHbKueE2y52wLQpaoMtVyIv9AHtNUERjVEybx
jYM4QKjNfXCQKIoQNaHMe4HCHgkbtM5eG3zqIMy0pjcj2Y7HUsroYz4JU7HU3um2
YKFB8Z3+BYFtmOECdA8N+H5pIKiOLFXxAOc4sT8XKw/7of1rtUL2O0SI+GOezKLN
9QKnrZQX2CWkL2ZIqF48zZZIUh8DQPG9UKh2UGgeTUnemtihl1ptjdxudd6zu7iB
AUYZhTtDC+iu+HZ0vbL7uvjtCodqfyCg6uMYS/wpnsWRfz89/mdXAfDQHTYzd+rb
ioq6SgJl1NI3cvPt7Qo1UcrhrFEjM91RlJQ/bHsSHvzvX2r6nNjFyNcHI9OA2Io+
ly7vPy48av+KpSWrb0OMlAB7i8HVhNjuJ4N/IttX9ZHuAMFrRjLdoRfJx1vIIYsO
8OkTcoAuesQSBolNu+EN0BgX8tDrI+PBZpn/Ujkz4CaLRMizrPTt//NRbqBajTBJ
NetCW9pH0X48LPih1z6AOkK4Pnoe6Cuj4Abrxiu5TfHviCTszf+siZg2nwgP+A7l
WfEPYDX5frBmdGx9mMKzBayY2lYLG+TIIRJU7uJBAe7AgDNjAqR6Izf97gmhudTK
vTgyyx7K4yuqH4CKBB/cti3T1HjOVVmjcs+uM7Lnc57VYSBcwpRWXpIeDBd0tgDU
pniPEbq4Ybx+89C29FzpRKzGjzAa14us6Ewt9Mh7Hlbcto1mtEmNUDRci3nkMbn0
BCErBlTHhTw5TySHNpbaickEmMzGCsXLKoldFxcdYVOfZWWnPrF2jl0pjSS3FxQp
DlB28Zp3M0QCNpXesBL7VDGUzNX0NEB2F4nvII+/eekKEgHZMSF/63rUUgYO25Rz
0OYkyAAAhkjnq2+XwqyVZB4S8MOVbirpsjK/MAFENH8OziYyAhL1zOhKSDGB/IVi
xFYHoXQ4UpGE35jF3SR35HZTrOuno4pB6NPQMw91dHwBIlgOJLb2mKmYhZjZSKlK
RsNbXWLFMmHyQlvPq/Gz5eywDiCjh6zxsCGcDYmiLGW1R8sREDVAYCMU0oWptM3F
gf8uOt7jrvhtmp7gPNdKHnS0Ry3np25Cdy1LGuxDWVxGcpFg53+fjv1oIiX7uOSF
TIZ+SYFYBN2S8EwObF6MUi06nMlvE2MDc3BXZwbjMUqpEFPnGl4M9DNwdIX8z7vJ
5AgwbLKsjRtWvDrnDl4aL2ozzLd3jiVWd+MfDads4BmdRu2VbpKSg21azhUKAopE
mcIy29tv1OM6WasrXiLGTjkk13RK9zBdv26FAZ35rif6KVriU380ffsOb43dnPOI
cMB3Bd/ehglrZcHuGh69Enbqo1NwkThbmxr6PqyO3MG2voCvxIBZ99b6oDRbvqd1
Gs4DijYLfuYfNvJseGuvqFp1s59Y7yy5F59tl5uqHEzMQrpjI3B+TbFaqyYLO4e0
Zp/57L/Q2v4YIIfmchs+l9ISGYqFgm+UpuSrMDnvpxtuKmzvaxaUePwXqtYvvAyJ
CSWxqKm0qIKx9l/0NJ8htexA95xxWaJEVHH7uRYn3M8nbvd3ivIxBY6mxSo32F8U
JKeBmt8ZqumQ+O1oSmsIBBsrtQz8zKkpI8ezv5fi0UvlPKKSwJ84/ujBv4F5lvr4
6hNdBRMAcNOUyD8SGgYwgWhRci9yAzNJi7K8H8oEBdMSvAVSYzOrkgJo+2wuZqVe
z8W4oAhPuQ+H7HCk8RKo0WFTwucsRAI256mXwa1IBwXsEaPOnjZ9QSpJGtVUpAa2
hb6tNZo8yZ6PInxo0w8AZr2NbLg5umpm6ObO6ukGuTaX/YfzchzNqwOib9D0gtlb
Df7WmQyPRupDTZZ7c8gJbCgxHdsvPxIKIk8p4k9w/g+k5AlwCyfrPHUgRDNFmdrq
YYSmykD/6+bCBKwjBf/j9dtvehi5VepORL8G26NVaaebUT/gEST1rgCL3Ge2WAIh
wuj9XtYs21aHu60Lj9tj540rJnTVUWD0ScPxJnfLgm9wUr4H3E8yZvxDaI45n3XO
j0pXDQfUrFUy5gdbiDEHB6Vmt4LyOCUlZse8EeFulmbx/mFP6NjilHhOTIbZJDm6
XgMAq33h0mLRqAGj9lh8cwscv/MyCiamTrwPrWRk3Ro8cDtkaxlfE/QXRoPHnqx1
tnj+ElWIgRc8VTck/XB1rEZgSCFGLeBRMw6/itJmzRnEN3xKH1ZtwQZBYwlA29Rh
xeYlZ8l8R9W6Zkwu4ozSusTiVU6j3CLSl63McP7k+QaYz1D+LyoqVpt8TD7u+P73
dAE9+uqf1r2ZFrEf51SNeKfoZtDMcG3nxxzGGEPHVVOjXA/3+TmKPsDCPm39ZBTI
fMJeEU0lWhF8vHxdHpULVfGCJ5G2wfN7bDPXYJamUJFOHWJmPs7pGeQQnnAQ1zxN
j72dXVUuyoyzEaqCo7wJ8xe1APYjj3Uybt95yLz54WKak5IXnG86YxeWYk+pBAsc
f+nuh9D03FeMjk08ImZ03MS2pO3FiUlxeS4wFkjeMOLV2Pfae7TLUNhjXPeYwbsG
wv4y9gtZeG+bhyeVnt/kJ8UMhCxQxJygETE/xvQIv8glr9OjRL68O5fc/tWw4yY9
ksZGAhLUPNoAK6UuWmxhHSwqK7wAHwa8gSZuwVdW3Mt9376XjGTZw9GOh3EmbvkS
L11KGkI+f/DkcXj86mP8hleWUQ174nXYLOoxcv/AVrV+pPRiiZqdjxMKxQLfaNzK
m1IFk+VA+F+HyczFNkUcWTnJBD8enWZXWKCzzb3GipzkafLlFUNpJYgkisPJYy+H
KWOgrVvcyh5NaIdW65s/Yp8UiUa4lGUV5bX+epE9xmhy93bxS9jYgbrEFRpimjuy
qzy63nTBixiYSeP3cj+4x5lr4YiuRVDvG21d1PX1+teODcCPaPHITthLmJ/teb0R
oGGv/X7JZoWIIjnkgyQYGTBviO61Lyin3ImjnC7ucEl4/tXSw8CRxn4ie/Xesrmt
xw3560Od1IsmJvi/B2xSgufaenvOGF5wiXoog1gXfMHRUlczQTUELg/RI935g4Jj
n1FSFg2AgaGNosvmw6UG5WDVfJhCAtl/Wej0ys7pEHukkgLeZN0RHXtVtsRTFdU1
Kb4UVTkc8NCleLoIC8Uu98N+lU/+5N5LbeBebwd3Idnr23vhuZL61yI+H2pbv+Fs
2twETkSSJjHy5CSpoCFyR38IUgK7qsAB3q9ln7pPbO7/3D9yZZzKRVML+o6uSUq1
KqHzvAi2vupNXlSAjJ0MPiJBJji/sjXIW32pk/bpPp/gVszglxEo/iwL36JNvIlh
ta7ZKkjTXJvYTBEXJ4Jal06vbuVIpDl7TyP40t4MG7SQAErxn9C68nUz5qAJ94iv
NNNBqxNN98fCJv8TVx8P8aFGqumk/GcjnwQekNXkMH05zx9Zu4jfNYm8EJeL7Js+
34VnDmOQsIk0pDyf6grF80YWTWKiGbBNUTVgzbLsY0nfknTpFjKzic0nIGzS4lC/
S7PqSG93uImr5mXpamHMZsBF7AgGyw7nGljiP7buiQ8V08gOdrMQetyUPY1HkDGQ
IKybfh6Kp9t2v3rsnh5hX+9U12m5LOWp9K9V8ViK2zDwRY4q60c2vMiiRMQr9Llt
yjZSw1JCATFTjmNs2s0nPZ5C0DYM8khnBKyNBjiindGWg+8DyuJIPAUKJUTf1W1r
W8+1SGD5ZkP8+jPUCi4hLrCD7B0VKP5mECDmqiT3hcEbbFym/3MLB0DsVqX8of9a
1TqS97wi5iZnuSr/iYYViJkD09c3mP6CbBpTKv6BhtbvZQN/yI7rj1MGsKhsVWns
Cx174ttK/98bQ6G/lnDEyiQ6KZ86Mmq6n0xGoqee93oWTjSAKzOYcAdsJepRKHCQ
czR7IwJJuaMCIX660aAIU1JxXeI2l9y2ENJXo72QVkhck72EqHCVrd5oiw0xgi3h
GRUCdMSMeILI2cyxkW0kz0CpYCX1vA1Q5KFAZK4432NQdDODbhKxjKWRdH/+q7ZY
aJjvDkZAVejj14psKyB0hM86qDQ8vaMyt8WaW6+JpFVvC7n4RFSoGABAQWfBp0QF
lBDmvDF8kZ5w5AuCfLiAqxvC2QkXf1LjlwjCDxQs4bwvFIg+MI5tijPodVbK4/BJ
B9+Ip62oQCAUpHh0ezB1sHY117/xYowZAUkzaYyGSi0t4Bzb4SrTmnaWrGMzruV3
Iv3KnUDSHZHssmBJXe/Z41HwAsxiE9/fVTzLyvgCCXtfuM+1qcX8nt1IB3b5ta/U
QZK6s+qhpmJBtIEHCQP4XOu8R8YEzNmCmlifL5uySz7oYhLQnNSS7Rh5hUFo9b+3
IPr9/FiETllxTFbsId13WcZbaTQKmOSJ5UPbV8YwhCSfkgv+85IyqD19DYBlt3Wh
jrP5wqFMqhzjEJTcjCWHnCuP9Yp1IVbEwg4ZrzAswuVmSml9tQKam8ksp9n8zr63
Yx6eqBDcLjzLk750mRcSLE4+z7FOcgxf/zWqMzL0n/XQdxzQYCuTDoSqewlNi6hz
EaFQeqsCdSUohtJo/WVZUytPHSCNGc3FeL3uw2xB4fEqQy2cRtLE7Z0tQVRMti5n
dpDZ/YXGhnt84RaMpNMLuT5IKY5fuAhEHenyVMnQvkdtkUnKID5GwjjTdIUjyIEt
9fXYciKHdWxHiZ4n2nPLWvpS+rBlwnDYW4JbhgR4ZNB7rHuVYwFdcVvQiLqwm92S
eR0NzqhzxBB6c45fCANYqte5YCBGEL4yx4lzZxwgHWjuONEkRNnZlQgTkT30o/E4
8ZnjV8MZJs8Eba1v9n4L5bZ1h+hzKqg4dTnT4MQK6NcAayqIQKt2mgFoEJWqh06W
CjrvcWCMCLx5jnPjUNngwn1FqkvJmYIMM7iOL+wJ9hlM+2ZTj/Vd47nQbBDYRAiP
XZtoWC4QrazSFFsG5VYooI0Q3wPj3UAlcEgm2+xcypIzaZDOElEAdF22De97vjJS
AIWIkATIcIy2nZVBsnu9QJ2nAeiU92+bHU/DuGYxS7Y9Xv/aIqUiKxxAiZhv51bY
sSu2qqYF+CfteDz++LFZakeTKP3smY/sHi/vWxOLQ9QaR6omPgSyNNTOXc6jgsZO
llhgeAFYKHOUZ119uZP/Fd4wWFT01+XJml6nfju0IjXlhIUvgAPr/h0WUsH6sx4s
bfRYnMRF0PkXqiglgnjwGerq3xuo4B9Y+yAZuEnrHZG7aBU0TE4hvfitIrF8GQoE
OFEISY1QsEJ8W4bQAl3fPBODZujJL8C4kw8vS2yxtIA5o+E1S7SaMMvuN5Jjy7gn
Cs9X+QmdKUj5XG2ln5vltNSOVGUesOLSELszbHa68xvGm/ZGrbrLoR++X17pF2vV
A2Dy6FycTNdQXiO967C1yDk+RufakBO7PkBwhVEnVzVvE7uvtR+x7MSTf6BankAw
0RbytAGSxPI4jbzF3cJP3jHO4k2QHvsDeh2a5a1yRSdmzR9F9YHU77bIPy0gTQ+M
+/ZVpr6n/IKZrsDCELJfC4Kq/VJT4RPdY+qIuPvkoQipvrKAPtJt8/Q7tk+VgmJo
WYeddwldNaClGSlrS4cN1swqmBBJtAIO/62e7xiRF8Xj07duT5h6+7OsB4FO0jcF
lwi6uaBgA/WxzLADcQsUExOrH2l19gjx3PyD0a1VUTetH+T3W2yKPVJs2cfK1rJ6
mS6SmEadGYC6+p1drfsV6/4SihuL8nMTvmasieq5jFDZcrfSEiVWupBg0V4/vz/4
FV8X5Jb2w6OCfG2H0nvFXu82aH5X7jR0TKmchxEkKVpu6YyNmY4nGHKKbVcyZd5K
s8iAOcMgkPcfMz9BApvhzNuYBm0staUaH+uIyYuuYZh+NANdOs530FrSGsZZBAzF
tp4CkyqkPBXcK2W0kG8wOWK1dkelspCBO8GSFBMXiv1dcnB27RPt52GpKL5Nizaj
Z85w7tcHzU9/BVi4EoMFF1eZFkP9Z82QXGiA6OjVjELraoQWCbDc/S5A6+k8knq/
Q2bHfMswajFI/hFSjTD2XEn3qefaP2VTHGJN5DP7IHeVnvGtH6pK04ZRt/PXQt6O
OvcpFjkWgSHWks/DosVc+1IHbSmKLMMYC+vvwLLb4wjHmFhUS7XKX/OikMRWSzrd
ouJDvo15u5d/ua0KfpfZ6bxwg7CJLQ14U/qg9PMzzAGqixxsgTvIKLr7FOBRA0JX
7+3G0u9+GWanH9Hz2pA802vTk4ZdCd2jKwmcn6WpDSzZxc9iHwnC5hqNuENm6e3B
cltdOqa5MEEPS/I94W49k5349cSbYdUbPiHmOAAzbBGYUuPmHOb/B4/LhwDtbtVL
3b1wh+vY63mj/H2/ZCfk4nnblrlBGDfuck9QnHT2fkZJDFWNqM+LFDshi5zr1QCA
TV4AaAQbGDhTouTkVWK0w0MDd1lXPZycDkQIMcJCJUF2i15LxRdPl3xnIbTNsFih
oDJ/LTroGXtZ7aqOwNbH3o5crCkBkj42kCA/x5DFtcaEd0dkIgiMDyrtq63tt0oM
GKLBHv8WRkofwXK+mbkt4/8bKauOeHPFU9Lkn8loZAJ1qGR2T5a2yTU1lXoB7fDa
6hJEK+j5dzQzoIhQ5vVgdzx2eWY8EHHL8mHnE8YvWqLz9vzJqoS50DOkhT6+WE4H
9oUEKQF7b3qAOkKRYQghbsm7Rm6JDeT1wAL4fuZoLvvPcE6fWKabswUhx/cv8dS6
e9yfh8YNa2Ij5tGL1R8+S7PDaEUGj6gIzju5rMF5RrdBlMvmAyKE88lpzc8DKsIt
5eCieokaIGnpW00SiYcKTqs1PFaed4jR8BNh1sl1eSAY/s5DlA70yqOQi7W935M1
tUo6xLBvjU7/XelckPZBfTosOzlQ9sNkD98egfAogTiisvsvR6cCCt1Ra6Lgk8r5
H6rSX4eJW8RyaJG8+QLDBJMYmGoVhbP/nJjsVVUwSDr9c7Pq9Cxx3OmLl59EeC69
w5I5NbQZixz4E/PzlQJdpCBRHqN1RJ3vzQ8Z1kDd73X3wlb30mFx5nVVz8h/wmID
kiaXkV6bFyHUNGd85dG09/KhIpM9VeGLeVFxjsZ4fhFuT2iSUu4djz3PwOTS5/AW
WnHDaoe5evh9cJCe7mOJZXYYmZFNJV0zUmaOHDz6ebR+gu3LB24c0FJ6tFy2UUX7
/XjQjpogrlGrziVh9SBtmg0R9kiZvO2iaat6Gn2oTUw+rkaC+tjh5PwBF7SCpSwC
42iY/X4V5ZD/nYlKsnOeAMswfdO2rXwa3e6m4ZNxJc8dHk0ClOoeS9pWQcNyNi/5
bYvb8Wf4XSjGIqAEl0uKSBhb2cY4Ued+1xW+sI0wfpIyn8SkZNZYBvqTObedFVak
DcEYG/VRSKSUe+VnITqt8oEtc9Y/I3IC62/WY1YiDa78n3F54R+ZhSj4sGE7vXET
FYXnmyHlLI4miDlFW2z7FlKIg0C9k7niujSG7UEsAYnZ50VaymkaSOc0qVQgAOO7
L5TiJSO5kif3SeJzPRs4BKVOtIm3xoHwZceshmbT+bvenGj0q6eaYaly2RJ/CPg3
Nq4JFwALkpVpEzpbBhRkzw5FkmvTkqoUSnN+KACbJ5JjCxn8Q0CqXELz/pJsNwLE
R1NhSiB2KWUgWsW0Iq9ItuqGWTKI3tELnqAiMgfy0wcAgjqd+hsn0CJG3T0abpyj
59kE5w8Q0v9Zjsiin6jui1BhUjL09rc+ayQwSJs+G0hzkDP5GvcTAMi5tho8KuB/
76o8F/1grnAU5ZhPZg6f7YEN9YnZbdk3mkGVvl31WumBgMb7leWW7trxW6GFmFes
kI4S8kXQ83oGBeKQuLHs1QCT5tcP1IYrz+Lr2RxXXCtp6nka0GpJubN49MEYxLWi
Xo7LCDRQdxixFjOleuYsFBV7mgI4rWMPpIta8tA6vZocSKgAeNpz/JjRkh2gSRVf
3uRKW3veu1ZQDR11G0qxSyqTjs0GIgYgJey82hvW+9b5jmtRWaqQhcj6H6NCLJlX
WcoyHYs8fIY1iFSkCU97s6ly2sOqa2+j2nrOeqSJr7kKY8W+M3wdL8x2iUz71oap
YvfXPqDP1pBkrIoKF1RIxHqXYjP89oPXaHQRqQQXLGqMctdmdu91cXEmSisY6WI3
G9+jMUeOiFXLtoqWEi2JQDV7NNffOhwBXw7Ie8MMk9lWjxkCYyxJB2H2YP0GGh1t
/ijmm+WZsQB6pBmcRr/Szf93uPHlJn8SwZ504Q9FMk9yBXrBxXhJMlJaI7Me9I3J
enC8gxKlzKA4sBAwPL34x+sfZt7w7pVtId2cqcvjoOTaeGecxsyY9ev+AE/kW+CN
QnbyK3wPOhY6W9sCpBomXKKbIuxhfPUz6ug4CQMlbdqMCYKz+sMmW5MiWy8mrdkI
RbwJ/bxRrzev8JG3jio0kS1Bo7ZK0nZ++ez2JB1AvOOzB7FSOwRk7i5ynfJGtdNe
eUwJi1MQ6ywOWh0NRPc2D0SHabQeH3dDY/GDHIN4bSRp1j814XU49R5HfiC2woTn
sZH72LATG4ciYEHJ0Pue2VcWFyUmwfy0hW6dmvD/Tak3AOTlHFVk2KWW211lnNPE
GlYqUgM/lc2BG35jajtLs4NnCTtpfAX8pi3Dk4vg+99LAvexUnOrCtf3kFg0S6eH
5uRiSTdzPKqVc7oBnC5bItdVGCFcgkr0kjpjFe8uHRllJ6mQ/ioEdPFdzLIG1wUu
vRTisflsWVTi73fxCVusTxsGNxXTfMTu5SdzYY20Gq5hBiLaYl9k+vcr2FUofYYf
ckSeCRZg3ljrmcfmQF41oTaJ6M4eHjm4Fnzeq6KDjczhC1EbnRN9Pt3FDIu15ByE
/vHXVDvZJnDtGO8pG1Er9Sw58Q7xHhWMphbX4/HS+wrPaKynseNtwWN3W3XQ0FDU
VXZEPkI3MWug7A5T6Tlpkg8uwJueD2wHxQYn8Daev9Bns7+oF9/tszo3PelsPh90
HVO3st3/UZVWfInLFnjK6gZWAMMLYTuwiBbX05vuTegVniLFAHQOjap+ddTyFIMR
ift4sR2ujp7BA3GLggQPA7SvRH9cm2gtJ+PtVJMDfpHn6GoJRDYkHYA/pu+4UvsH
IpbGdOwDoAP63SzOFkPBPprjB8SrwiDt1lviqvD0pMBVB4pO6jzJa7yTuC0U8JrM
gl8K5XqC2eHJrUrKu57FMqa6FyaBp/zQO7njUiqaUDoZL72mUZ5A70H4tqqmqiwF
VRPPTztpTjYxeg038q8qRQmI/nbi3SRHeP9cXQdo+vjyKf1ZiIjwat3VFi5va+pn
taAgSA9jGe48vbOvGM9W1GahhQoWBuNH3rrZvlKrhj67K/wAFJtoed/isgurl2FG
Pqv4jBA5m9uuvbGJHu1NjZnhFD/f7Ins4F0eTb7cwKu4yvIwqek99cV8KW0EY/eT
SNbNDehRYuq1kzxiH+FqeA3YmzNlkFMlYzqkw/jqMAsi0AF3FdZB2RVSKqXO0cWV
lMg5RaH5SdZuLitORiVHyiZHc+4QgUHs+NuEmh/4zL5T4xHeoK4zuh3UhkxdPEj0
IKxsYPmW/uoBZWvJo/jzhzjgERif7gMD0IieofFCUM7ASG4uLZEbvXSuKm5h0IMO
MUTXUh5weyPHKtfPtO8yEqsYHvRSmAjp/Ww5ITqvE4ujuVz3TaUYY0BNOl+hn/EO
WIf/dHaJcq5Z+UL7u+y6rNK9QJrnj8kWJXAI2OR54xGjxCfvoUSrgTNRm2gj37Y5
AsDWhgmo0ZPqr4Wl2HKuUXRQSD3BDmtnmEfZQpm4auXssr/1p8EhT28J55Sm6rW/
8cHJ1nmCBmbF6mECu7RCg1Pzup53PWYJjX+JHOHWbdnFxFdeGgeHn5ESGnT6JN2c
ZUOb+Ao1OdZ+QnOaYnkJeW/nDTzSB5b8eQ8+hpDh5Zb8yCVICiYcnk+Eqg7wb2qa
Lc4Sy909aH+UqOEaxywre1gi0Bx7/pCYdbiq6k8OEV1UiEyj5Ky3E93w9Z39glwi
kHiSR6YvvX1XA7YvzuJotms9VHI2yGbNxYrebtc/dAnn7lsN8ZHhPlpLoKA6JFIC
eFgf2KnAdivYWVvQ5E/B/WzhW/FI/0oF2v82r0WwTl20LYj/lH+1cqwC5q9GUGY+
KAtC2/gEfZuf9oMXuhLRFbovXJYzpjgZ1OygtGg7TgI1KHL7qQOpnNqrhqCAVXcP
uZftuWAlJP8KYoHLavgJQNyvf1Go9gNOYc7iFn2Jv+/WPnHkpbaJlsZZq1aafwas
os4+Sv2eZ0yPtXGSg/lilemIbbrFAQCrQuHpsrc58h2nFeXUtx2wKQ6cWxg3k8Pe
eQ1PtwlYqiBFisDJ53CWSv/Myjvy7U3TKg0RIgYV34mQVELRilLzSnlD+qM7XGK3
5qt7I09XI2NKMimZhMUfzVgCV5gLjH2lLJMkkC0DB4TgyDvHPlO/VFE0G4Zh7JqY
CVvU4R/w4zY66hRYAUIi84IASfw396A/sp03YroZFPB0v25r/iS9L+zI/0VT+nOY
2jMpkjnyPj9zFjnbynCRYD6BHeaLnI1dIW0i4ucovKn5wBovUHTadZBYOGiWwuyR
meR23mpLxnRM0ImwQPJ+tAQecIUOPZaa0Y64g1oYwL5G0IBaz+x//RfotzKEyZCo
Y+37p7nr2dkXLLVCQVBN7ULnflchMYerDv+BRJDRlz4x3BE93dIKVNTrXKObRcEi
g+VQqETLpySYVQ3LHknmjjp9EXlmUSodjRMVRFckf0AO37oRQJfgqhmrUMDXArzl
SrsveKPOdBNk41qhbQiuQqh5sEkNrn1aCEbj5174CcV6XZSTFJFGqCw7iQeYrJK5
gj8rY2XPPaJYdWz/MofpRXcRnpXTDXPvmPUsuOx053tgFal3hnPOF1Ub72SPieB/
LXIDkJAjYqYlsAYNsvsSYp3BaImTYTBSm/W9/Vxh6gPMcOtiJLoXaM9feBJJq4cs
dAmEKFrdbIV7yzFxwWebDWuVbbISf7sk6oY3P+MIw6Ew1m4F5F/M1KxX60QITOTe
j3rIsZPHMuNMSImRzE1jc/RJLyHp4TCffJDrZro8x4spfhRu2cGLn1VdvY12tiD4
EfYqUlplQInAAoDI5nlKdy6ISaoSZRRWceHCoeAZjZ52MCptzCnMNeEG4GBDhTA7
hhSlqvi4zzrrkSR0eJZ6jd24ggmqGwE+C4KuI73UWi5NmpoVJ4JLH0axkebJnkkp
BXsB29yGHwswc7E7LH0Z+JIE+K+HiGdKP2XtSogTC+YKhS3VcHmfddn4g/OLcC70
fws84muEeNXmOKKztE9OvQf8h+ci1cY+szkbg60S2GpySJH2bmKKgGsbHTI1rUgZ
ho/LjMk6O/CtkAcylhVZEsSeGT3Fis+IDfYAF7Wdp9YzjL5TsqSHGStZWuzZ1sjO
5zx9x4rssLO9EmLD+ptkA/Clx68QuWdrSzfVJ27Vvv2jKWN/HsKta4JY2uAmSlfs
zuT+uABidCV2idhU5662NiqV37D3J1hRuTzMeH+q2CCtw7xBfVXsh87ECT8hBgjA
ZCJeGEMWrDpY6EKkm59U7Hb7y2nigdQhLXsdu0xXCH95FKTBSieYSqnp9r3lwNX+
k58Kdz4bx5ZeqVwaPX2noNIBRkYnGMzllezDXo15kVVyMCwN8ciMnE8KJr7byAvR
5hQ+hcIZalB2aqPvLpyDuVNPRHM7tE452O3rQnU8wr6m/os/VronvLU8xXD/aLcO
18R7AtlOtOdi2zfFSMqLc0lRhvi2mRiMDL7KPu8/NTVcRM17DP0ANd+ldH+9bFb2
bK1tpu8U2f459LvGMvUo32VJv8c5zYCtLa/UW2ZdpKgEEx+DHPxxzYX5dDSdxfo5
qw1pBoQm3clWsPpgJRy60oFSmQd4arbsSvobOYkvhbCggMOvbYEGYsU/vn22D3WZ
smSpb1PJVFm62A6cAnOAIpu3KTVGz5QtYV9hEVeNzeOd1b+Sq+pjHaKQ1ucr0qdw
S8c5iPEdJ8FVWpErHUDF8nkbfTFW/77mTr4cO7qLYHd0Djq04G4Q5S4dtwOHJj0I
hTfKaKy1WH5n3hZJqenF9hkoeROJ6fsiEjUN2WWkmX5wTBErnXQG7bDacpdfHxKu
ep2xmZGF0EINYqJImgSYPlh76vXmMYEWY+7Rc17WTu37jeSvl8MRGIrEz+Y1NGEp
nZdICXPM/+Xe97bM6AY+yr8YI8srUO5m0GefsHEVbRiEVKudvVfvnOdkYnOq55Js
joh+nJndgS+mwEyS/KRd7dv6eeVtdH3r3oBImdAOkmUp2OR7oNqTsL6IOcNmILrd
bqyOD7Ei9nyi9uv2t2uFBFCjKpmADOKWifdYnZRUe9SPKJrPiEjbIM2mukrbH3qw
B9Zox2tMTNfT5wTdSD45XRQjbTXtPgWiD1m6ey0vBN6q0XkN+gjrPbLwa+JUCu5a
HjYUwYrKQjV60wxORYY3IeJupfp0SCpVXBVQ3NDeC3g3CddKu6d3R9kp/zk5mi+t
29lao0sp52o9tgc/7062JOu2khMv3Bn4TC/lY5tb/t3uMiXHgZEC4m1FbW84/pjz
U3vnjgYkCk8zsIzzmCriirSIibKsuupWYrvyDdIp2IuErWjSbf5d3Dbso7BJjTzn
qEGVb0D9fd8DTG67TaTak+CZT7+YLi22EGEuis4QDpnw10oX7BpUhgL19UwwU1VM
jYGK0nTavNAmzul63JTIrwYuC8rS7OBqlrdiW5bNQ+9BKY5WKPSQWsP9JI5rZHc9
JnCfU8InC0WRGWm+JXC5AdmTL2QT5TvUa5fhLZxng4Nj/a7WXJX79IAWOfLRZpMB
7FcEv21cjztl5TXT0VJsu65b0X4Bc2X+EE4YIvvIdJDRlDwpmYI9MC2v4bRCsmW7
xQoWcvIlR0GLwjYaR3TyWjLwQjz1IytXsTBpaI065gE9XuuBWcKU0v40UZCegRfU
4OOudaEcJjPCNAgDcatTN/e+uNhQLN11M0xNetoFX79c4GHYKZT29fMwxcx6PdtC
stGIn801hLjRBqtqo/hYSWHGFTOlULmyiJ1t/O6DHfQMZWG5rCoC1A+zfeJ0KKw+
YPnWJEj54FvTgypjKXXE+RDbA4nseVoWSNuLkhtrW8DFRq1jjtPl1GepJZikGRC9
jJtCsQ8PBcyb3zvLnzUgAI4C9ENRYLagufVVxWlDdi2oKq33xz9jd8gIfmJZiual
GqHfKZPH1jtSeCzjtRQXFTv+hXDhBG6RQ41CgrDVByA2zSGH/Ie4oRMh/agT3Z9U
atFiuZrdGz9PCs4KfXwu5By4e9WP/MLdjRu3n5G4cBOehwahXqZaJZq5yvYJaGPj
Q9MQMfxA9rlhlET/H3ZkKX7/wSuTOQVp8+Na5ljbAD2cg0EWt2KdutZ64KfUU/UT
H8DM7J780x1WHNEIitgK1RKtB2BK3H0zhxMff9sh+aFAN2Nzc3tpM59v6ubIDaPZ
oTisgWACDS4MQRSN2dw48boRUkUybIaZjrfkT3yd6HmDESXFcW0Vu2dZXXhbi22e
Rcjn39MkqR7q8RCJGczg7e3bzblD3kT+1CEynuEqWWm48fBPFOPrUcnZG/2kY/qf
v367JV76m5zGtKxF2CJsuxZ2neHBe1ccMs1d/Sc2j86ZMh3N6mF5xUuoNIWdWT4Z
WIYyyN/WBENQPHaSESc4kLhO84nBJhTopn3RxQrtD8A2+JkIoDT7RktR0Fl/CcvL
MvpgleHg+24p0Oftlqveug8CUNPTXNjx/7lw8irdTnVSczAFzAZlY/Hg0d1gRA55
fhffash2j6UoH4YBBSkMQitxcuKyjwqRh60J07U+nhWbvhllrYZVa/Q/o/P0Udgq
IVIuH9tfiXTG/FeN3nx5cWHtWtbNCkvnxrkR8slu/2G1wcxE8PguoQANk8KW3u0M
YLn9JZf7EHNkBOmFg911I4V0qUZGndN3qw0OUCWaADPHiZXIHobnSxsrQojKFDYt
Lprsk7uIbGx8xSKvSK8UPCE6qKNfZfWmiJR6FJ3AjnYBMqSFyaLLbt/LKBXlLybk
nXeFMHH984jhv5g7+88RmMBRjAaZ4pmavZwhJSVEJtS5iwodp/rPWRzrC12PJ6WC
0scNslN4HyINS6PYz+eZesISf/5S1mmFcf898GTdXjyIzjSGDCzE2IjcO/mBl6P+
KwNuvv2Iw1Zt3DJGjhxPc2H74EjchPy5kpdoMW8bmxUDnPmtpfj5uPrRbARw09Zz
IgUT32BgJwEgpj9NWd+bX3GLeLZMFJCd7LKwEQqc4psdHKnxi+tqe5MBOs5AgD2J
LjDo9jh8rsSK4ZArr8x34Ai91FS59nZ42VgPptw9V9wRYBZx6GZmw86xwA3BTUVf
6WAuOZf9bzvbF0V8oC1/jCLr/Vd5SbMB7F9EIy/4Jr5jUPa3mdRlEIfK2esfJ6Nc
aj81amjagjW7l4CTe2n5jyCu+X9GVccesaAZzwF9U1KWWX5vH3ft9XYBgd9lv0g4
cYDRhXwSPyIdHpISQor8MeTzTZABNSyf1GmGMCoog2tI+sg5jAeqMPVxGaq1IdzE
M2/5/x7oqPjiJY4H7ZIsI9p/RNG9eY/W+MUOVzcDXoRHPdVbJS2Vy1wy7Ko1Fcp/
SvB8fk5AOgVQetsdqaDni8NSBCJT8wUcryPGTVVka9iScs/UEJt7jb0+vZafX47W
df41doZ67he8pFoflS0IP/0bIEf8S3lpDndtwyjhfvm0+n2QeV1zVTRZqojCOhEu
I1WinjiO7/4W9+qPM4+faX5wMY3vg+fQdRXPwkIlT2qs7MYCz/JxiVn22Gy+4m16
Sz5LQOWncgQXvMBH7y6n/nB4M8clSBQmMRFvOGhPNQ/eCTZq5maYR3IPr/ollkko
d6Zq7vQDVcJ0JVvnVNLWl3EBlpsk9lc1nqdd9r/orv8VYdUtiogiH5+PxDRjoxQj
0dA1LtqlQ3Yx5CNowUailn9KXEB19oAdhdTnJxaWZfZ0erQZ0TWDvG2V+lEYqyJA
SUfQAh5ZgAjCku3XyL+LFXBlMbXJ2ps2eixGPvjtm//p+7iF+mwR69lbG079Ex4a
3noLU4tCyE699qT2puCff12nl61fbSSly3Q0G3NngENJj0BqtIwYxCSyWfERa5Fo
m/3x/JCONonI4L3ccl19MA9COCmLz1UwbKHXuCAIxO13CXmwWlIMScWOQLr6fzHm
4qn1gvTJf/JEofmagQ0wWli+OspyFXnQPpx1v7n+BxGlAAxwpA1YaAbFj9WYNRNx
4B8sXrAtny4D3YMqQUQHZ+ZUZO8FF4CszC63Ig2eDBYzutlb78xVvrqKuPzR3Cz0
YUU5b+R8AcA33DyAIOECvHVfFLwl1NRfUZyV8stfqwd0qu7iY80lI1kWjhlaEPkh
6Ox4zvZNBSC7IaAvulfyvENeDhB7dMbfc7AOpzRdi3vLHhrS8T5bN9ll+2B4Cw13
9lDt7ybs2zltZfqipCE/LZmqf6pXp5QGgAzjMVRZ61JLau+0zGtlsLUKZG91Kgby
oPKc9URDPn9kbMOQTWAls0ToRzsmQInasFD5cS9eWoFBV1NOpUgxqeds3jYVEfwp
igNLGioOGy6/QHVp0t0+MZllNFGcYBfJ9YhFhCSIQrK6Dy1kYKLbo7Y7fDffAegu
HWs8VtBpiR5hgPCpiKjnv6hYWY6s4AbpvDf7zpV22zwKNXh4H0Uw+ePKxR4wZfB+
xH2l4F3fz/+zpq7hhZ0DPpihCmfh/P8LbglsSeTtucDRSEV2emGidegjrUa0VOhJ
TQMcOtgdAUsbrn2//UXLyCwcMj/sj6Z1XXnnzI6PxE3cYxBsEy/T6XOWRMP+1Le+
NI6sot8SclbzVzDl3mVdX9siprAMjWTaFTkIKf4bPqKuz7jScb3G+IcqUsR9D6P/
e52wIm0JFLTYJWMSPJs02iBbbZyU2AUcr1libRHyWx5UQ+oSjxV9w4BfekB/rrGG
ke9ZdvNjfFuJFPoYPWDxsG1KQGE8ZgiFNUs4Kcx3XCcjmQrpQN3yagWShfz4k0Z5
7uYdZRzwjR0uVqxrhTLRFA22Vh9YoXYWeHcx9kEZpnupfgMQjLTxLl3tvThIl8YE
JOd8fwenQLt7gLOSDjZXSji1Pzy0vuk9yhHTjNNOwdtGXUaztEo4BCGMOogEsUUC
Tz9qKOyF0HOndpQVFiyKR6NM9ntVzlW8Ya7d6d7ey7vALSV4zkAdTLBcSZIxHu6e
cYPZHpugdh7pZMZnSd3tq0Iu0Xf/TYfmCdWWvkXqSURez98CsKSdekjezrXR05h7
N7NpFj6KaWw0KVNBZhpOsxVs0oWZzgCqzA9kmpY+1Oimsm5NE6XkkgKyen1mRVLo
NHqD9DKGCe2eZmFmEaqaUNHMeHY9p/ARSDeKKqujh41MNiRwPcCp+vGFoDVNaI6J
40LnAiSuBCHnX3+CLcpHNUxtFiGpWNotSGFVB6DrNff3S0b8Il8m5sxRHq/OTdvw
YyMWf8QQANIyToTnHaVVjOC1xvNEkms6jOOqc92gVZoUzOwzeP8r71VPkss0roxz
6feAdCzLdw0oI2JARvFnaQASdm8pZJ/aOwjK3vrkQ2hWWW91ekV5qmNGcz4bApbH
hm/8DwkgRUmlXxo2cu15WuXccCjTkNAaWd9r0dOm/EAAh72g6XLTCWx8hKPfboIB
6AYacnVCuwjbbighb4fidnsRdFxvR8ZEJ6tRhoEu1i1aMREJYF5PK1miE+K8/SXO
4ZAbBmZGZRtEtHQLGhnYeBbM0ZqvlLOSVfL6OPLpASfCKQo6oC8exEYAm9Iw27+J
JbSxsxm9JMQXqpxfNRiWzzHWNlC6xa8G8YWQ9FGWRW/2qpBCH+OeiQ8sfE+Oa9Ee
tLXbsqO2ggiaAbUye5ULIYBcuiRoKWqzxS73OAxgEIOJcAN722FSKUs39FR6BQbI
GTQb9lbdOmVMICaz2n8pDtzUKPPyHgLJU+BCh1BxbJ/8Ecn9Vm4zE8smBV+OqlFY
tP39JJLKSxsb/A/yJitxNYb3XLvvA4gRCcxurs5AueKOCxWx7CkPsNdWpMXZFO3p
acIqtUTese2nse94n2/JTCMHZfSlQKKscLTf0nafulxVS8C15lWMLQs2ffd9woNR
CaZWkszPQZ0osWK1C5YU5tTv7BM2eAYXFmYDdoe5r7x1GmkxvzlP8S16q1xdeJfW
xpttcs1oJ1kLiJx4WAYS8To8hg9GEzZ4z1rmAm1AA6nM832wEwXmvdRDtMb22XB/
0g6trDahwme+HBqxTOLdZ7+clqQqfDlvDFYaAjn3ccdJj8D1U9qQd97aEvglCdzY
IolnDrG+weDbTjRtQuaC0gY+W0PELqFFLrvtyUPEZAB0QRuqGvdXiRZfoj/Xru0m
PzYXQTmvRLk1yJm3IJMiDgH0oWYY4hASeoMlTW1+aLSKF7NUaoZb2UKkkQQ3Ut/v
BRGRDQGHXDjpuSqraK7/rdo7CjaDi7JI5ZmJL9mN4SrTEPztR2MVmC9MO9daGNE1
pqUSMH/4USNrxiF4KIk+vrHgt7UnyrRk5rJDdxgHJWBhgppufqJLW6snPEFIeAf0
rrP2ZrwWQTme5XpsfiQrkJv98YnXeO6d6hu/JZV07Rr9jdzj24Qu/ZrvuJfInM0e
/bDqmuAo1R4jsvd976ATHJPtZersvf2hiE9x37Sk8MNEJO9bd4yjCN04kZ8yHQJF
zYFmfTXjBOcpFRTI7tPdlaXMirD9WFOVSYyW9KPy29sCJA1CJPnMSJ+QYlYQtiqG
3DEI6qxnkvbL6bS0oV8al5tj6HJ9Z03wjkH7zDHQ4eVxGSc8hDsf8/0JzyS/CtY/
sKHB0uCONB7w5vvFy39GaOwqwmoULyHOzZTyIehqD7iWlSNytCz17nE/xN6XsX3e
0802bN35xGZivChnPlGeZ+sG/9GWMCdVlw/FAEu9gBQfF75Qyf3+bpohGM7evfdp
ts/NzS1xmqpAshmOmdbbDekeWAUjgU4KP4q/ZHVmPgxKQDhBeWZPAwymw3/AJwQ7
URRkJ3d6oXF2pz09UZWBazTYMmpp3Z9RMpjJkFSsC6ZaqTkfECXyz+4ybBtUrUiB
fYOHdXTk1zXvvAz6ukMG8a3mor1S0ZHgsKqTK3bYH1iqZHAHH1lvUPR5ldw7kxky
swlsMjce4R/PZE3GGiziiv5HK43rwkOGSqVbo0An7AYQqriPp/gQIYfmyuRAkUB0
bsYUYwFTcULPunHEUuZHIeMPdbGoEjpS4ON47+2OR2NVqVVn50suJhh5IJltNddZ
RMr2Q+/Py668vvIi2F/LMUNhTUt/13sRO5aK0tbTPVe6veOZ6YA2eFv2UsrXJb9z
XpELrdNP10LXCpNaJS+F6T9x1BBY6i9uBn+20fsxqdWI09w7Gc32y9SQhaatC4ob
G6PaFrHPl0cm6QkakNOFSV6wUsI5cpiFAyIgL5f4svfOBeHMQ+TUlxEisWoZ2OBC
mJdF7n/Iepc7bAlwLOMx57G6fNLV2y609Hkf0hZ/MIBLDWhXysKePNsddPFAeFLX
kAmWbsDce2O1N/z5MGACqaQyqlzCqlrLmx/4Dd/xVrSgHaA++Atqn2RZTd28+6s1
QML9jXU1yxiZyz/UkAm1TYWQQVzMzDuHiH9iYAAKc0Wtn53vr0TN+RT0qIHknjsN
RZo7NlpCiYworggcSQkLe72Qj1kfflhIzhq3Hpyl8XSl1fxMovPi30Yyv8RRnE7Y
umKWdZJMyFMoQOiig/BHtZ260VbsER82AP/U6KNQdh0Ej1SE5+7haeyo7Ycdgv/p
lW5WWbTUGiFbfuk7YSw43ZgNVe9fThWmN0ie+MbJz/xukVGB/FW8l+m4LYfcmO3l
NVuZ2IP+FB9SCansSKjBPmYRZIzY23H2DN9bEUkLpQmZ8QH3KYIElqK/EEyLLbQ/
D5Iz6ZpppEczED0BULWpDcjWHE9tRisDpReKhpvdJW6ZEbsoZKmPxqSKqi4AA/z/
j1jC3yfDTnAsFEef9tyZsJVgdIiXKQP4YKbL82rBPv1gpm0Z3uBvSjQE0glcHI4U
Pl+Pk+Pf8cXvtAwpNTeOveMyEfMCJjralpMwOoSb+NcBc1kVpekPSyMuotUSAsbL
sPKYJgfkQ8xF44gHGS7P//qInkbj7Q6tiJG3/8oZgJVjUWuel0CGWchW4ssr0Wmd
cx4aomLo4eEz8jGtyVNGkK3R/uwbaWXDCakuVd8c7mjFR4c35ZBsm6K0vGDNJkAD
q64t81Mhx2nLMS/KRYww9VN3Ugtr68C42UqumHeyuS3iwg4uV/Nyv2UK3zT0HPBc
r+uMijPdxO/E3db65H4j9ZNFRx7qUDv+cp6XAu0Oo1phK13P5Yxybx43ODooKg/9
pqrLks3JGTdfrFmCAQ2u6dE1k3GuXWw/z+YxFMPh4K6PX1C5bOzfSSNoF4YIpv0D
aVvgExsq69LrW6xH/PPjggRiiaoabTZCYhEQ7DWbCuFmm61SBkrbXgVT7D2CePKR
zJTaCvDBzTVL3u8gdFyxRBiwk6O+TAjjxMTvzzpL2UazSINHAMUKS7Uojxu77EVm
Ym7RFZdcbtgVEAEM5rMv/O4WrU2VAkm4qeM03cDTAopBYBB+Sen3rji7iKE1kK4o
nj3zdygt2VZHJUKcWJVAS5wIj78V8pv8Jo3AJZR6fx5Pn75dhb2Pe8EMD66WAHiz
eNIm3/5wZxLZuZlHuFqW1znAPq4Sde0+TothDRLyHf+Q8PnEIacg1ps0D00JNuVN
oIhGjFqEf9q9HQRxrQTKTCgfntPYt0+mRO7fPyTUjWyNb2KxTgl1aDxWN1cZAz7D
e3jBD8n7g0GutcCXnfZ9H7eTP5qz76BTLh3eKBryedHRqVZzISyjb5FYUm1tHtjY
t3B+LVQGhTdk3T1/qSi19MTmUSgfUwq1t7iQw+L8FwSUNYJ/gn/1UxHG04TWkUAg
BWQs4kfIbmp7FR7Nf1p4TRzkaB+e4ToKj1diodBwHKYA0GZAHohau2k82P27mbUm
e4SDPeRLsjfnVCxLmfX4AVE1ZwhWCXzPWBx5rKJkOohcNOg2evttfCpTtziNt1s/
33jtN20tzBTTXil5X5eeY2LR8LE8CSVpKdOfT+r1iJBRElIFJtU5WZq9BO2ThglA
gDKVwxCsCQo9cuwwXaCtd7UZ+P7Fx/JAUa8JJKlNmRVPMqzFpq3363+JmRf4hD1+
j08lGzJiv3Lq1z1T2QGBRx6iD045t9IlbTr59TaY5yJ2MhKWQq3bd2F8mHNhmk7o
/qgWfY34i3rUlakN/zqUPeMdgasqSQPXqHzqc5pY1rJ2Ufp85GL67wXA6j5V6fSr
Ats/PH+QnzfaQFRDL+HyMmREKUhYZZ74QXQOhH9FuR4MFcpIsSozd5S5EFfXC3th
8kKhIGd3G7vdnBlp6D0Fu9mM4xrOo/uNZl0UOAg9CJBGShzpMbKM+5PgQ29bQdFV
643MAQZ5gMGn3S61bbFEojmlIn9EBEAdIK6Bi+mnChTdtIHUSYEahUKi2VVSOKVg
iplH/CwNO+APKMnw+thH2FgTt4t/48GPmjQxj0ToCvJan1bDarhEeMSaZLcNucuK
Skp4E9ufZ2ovRmo+mZAs/C8j/fkhzEkTxtT3Szzqr3JUD1aQRo20RZO4PlDwtuHi
bMaZuHKCxArV56nFdoLR2UOzL/zxztsdeGSpYRLZX+EblJr5lQ0hIF9mEvVmCyWl
syv6V0ZXOl/cBO2cv4NdTPw40InOGp561fM5u3qBbBG+KdQnxL60aAgI+waXQV5L
85FGrxr2fpcti0hPfbg9hWfKGh97eUBni2EyhE7ViKxmCG/L5rALZ48HYNUuslUy
zy5d/TXWwt2FekC7vi0jPAO1+W3woAglukiD1IGXQLi2c2DFELqO7xHhxTvflKNM
+r233j4q+M/35JNd3WpLmtR0xmtITDF8m65H2FqKPIQOlS/pHFIwgKnzTfDTTTE0
BrKp1N+ARGEVR4Y4rA9qCEyq2F3IA4M7SwDgIDyapFyS1KZLdtENu2fntMLBWvGs
YUNJA8as9pEpb2Bt76Tz0xaLDvFKrHOmsjelKOt0ogYdnlpiPiSFkqxKjZSO+lEN
2xg68ZTO3Papvzsk7ICRfX+Q0LtYcX12FYZPrAONwhABITy/skQ8tw6G+KWwXeix
tYweW32pMKj+1zlxfttM6ddPfdaAmiO4wJl6lyoWmVIvoV88Ae0+ya5sReZogSp/
6nvjuLlnangNcFy8+AffULbpKCElfB1FX5KeSD/KUaVy5rCGf0JPj0QjegQUWaRF
gMByLTUJ+n74lRFPsmpcf44buyYWHU+FoQWqHG1Lq6UvNDvIcW9wv0Xlmbln/SyU
o3XlTNkOlIKzs59+NuiecIYbhhe4upn/Yp0aRqXZsGt6zEtJqeDpBjXIFdhPv8jC
Ay80HnOWCwB3DtEaxEjkMywT7Uxv6sxAxwsoCUPDaPNcsAfxVJ03oMbvho1MH4Sb
wE+wxQrP86vlOPDcSmLyUhWH/wURgZaDrK9DbEyomA5PKa/w3ueeQtvDRJhGF58i
ZQ6IQwpezO3OXxztBiXdy07/Dnd/E9+X6CuUkrXbPYnX/gtS7qLc8Lqw5Wqhx20y
eXjDtG2FqO2t1qpicoMunY076oy+zpm7kRQItdEh8aRgN+Y9DvE31x1sV4mqviDD
D3XwLTT4kcQrbUTpT/DFTc2Vn9/uN6Z9WDkBNUizyD4ZCFHQ4jbYJt/avP2wGDOj
z+pJILCRa1+R1jYFElsvSEuo/vvIgdNsoEjx354Z/Oo2n+dhFaxmSALQWnmbLV50
bm/JTvysuIXVlprvKDvZNeJXg1vaXOwuLIeo44RATO/VNIhg+bVwbimDy2qeDlw3
TOMwXJ9PcSp/Dr3eAXcNA67qRhEktot7vZau9fTz7f6MFWA/ORNAa68XfhoTr2hX
KxrIdx6vEXO6lemOG6VWwRJ5YUHb0mZXXsNhFSt+BCnB8Wtqc2lR6WBdw7APd94e
lpFK8tz0DwCoZeLxSqw55ta8RFR5Dsqw/Z+xPvNWZsN5eMhlw1grSYFOO4dU5Aau
RHJaBk1D2MQCuCNP8m1UEL8KrlPLzc8a5ndqDxfTl2pZ870YX9LBJfib2pZrfTNY
avrUOcMt92ie2gGwShgNS6RvG27mBOpn02FrojqAyLyoE9c/7j66L44lhGaFxnlH
W95E6XCS+C/PbknYwJIon/yqtv7ubyRgXgOkyE7MG0VjrRv8SqYmmww9bgBiCuyl
6uFb/wsq66fxObdkUq8sk+zypxtTt7E9T+g77NUdjXIAVDn1tdteljD4H5PGbS0f
VJ30y7VRHet3oPKAhyPJM4zucSxrzfgmEZQh7ku3cNappRoJy8dYKWS2mV8YhxCI
Tc5/yki/V4PCFTthXsIn7RWf64GRrGl+lzAEldqmefmMAuu55LkcGlr9cM5XqdKF
Be+G01VI/OgYJGJmx6zNaocXyr5uUoKlQNO37K+2SKiLYcTVS0GTECUs2PMG+jYH
TG5aPqGEc7l7mBTHapRhQblgz75X+822H/Bb5O7Jj3UV1HJDwrBDTw+eiE6TtPFO
CCx98Yd6JrCmMo6cizN0esnkjxNVyfWzjSLEryo4QpVxqXjEnP89qHJWj6OjxHQB
X+dbfEuW4cvsZy5V8psHUV+lWgsNtj4UFu4DiFDmeXOyRUX+gHT04qaex0aTi8gG
f4WxgfcoIyMBA8poFhVMYIdzfb3t86Oi4pHpQ3n8g+yZHcQ60/1wu+2/UIqMlXSb
uzrI0SzCNy9G5o+V9UH3h4TvDgK61nN+tmLNskHE77ThN8yTgap4anGuH1s9XmOU
/47Ohb+tmKxR84AgcjalbCJWSoOe8A3MB2TKVOGVPIam4gkBhJ+UdXXqEVkw9dzb
NL38ElVICWXFKL0LmnusacglobaO0eKGzjMGC2593B/ZM/JIsuRk4BJMhpozbdid
J6BfF/nmiM8PWA3zXqKVU1QjBbdURb5g8tWCZwBLgI8eqMaeopJw+69yc5dAztse
ueq+CZAvNDABhBrRoOX3ycYHyK7Z2Iv8PgQfvYWR6izuqGCTeR3lNHuqMEFWaQMF
dTKaRVYQtZG8KYoq1skxop0s/hHLyS2m1CaRnG3Y/Xtatoct0xyu8oKoGX+CjaQB
dDLouYyPOfVgsWMnyxMQ4U5ITVkqhfSrfsow46dKbdKH9Y/hm1GM82wuXiV6t8+U
rnojpDDjCzF7P5fzIbBy/7TBd33CJawymSL2/gepfe/ludpKqy18jh6vxtIuZikT
qDkkEhHiSKWyw4EATxXGqOKv5EZ6i29ykTv7Ezqyzb61A7HKn3SmRSjl+fEfRZi8
l84n7W7lSkXrvlYCHFAZzniI/pHB9sj55KRAOWetG7K+H4EMTJPBixKhy5VoU80e
J64ZvVsSOPE+pgGltVo2n1ji0mOveXCgxG+D1SsUIP+aLrxy/ykk01cpiWVtm+Ds
CkbLGBH2wgC+B3hqg9TpanbeG4BihXQGkBqceJxhrqGLVRBitflav6teS9p5T6q6
uMwzX1CTCQ2lVouyMdvVbQ8s95bGuUWPkeY4A2V9q7SaUihziV28FA173sFKvAeu
ZIgWCRVauQlQxcmfDOwU0XaHKIbDmyc708e0R0tGkCWrYWWcN1qIvcy3i0k59wMY
M16RIKuLaxTTLzx42/qYXAYyJEOODSRMJXd0LV4p8p7r+nECVswKerHh5N77AUUx
K4K+uF5pRtgd26XzSUsPPKbSUCkcZz7TrLlILtYf8FoB1SYjDVE/dlSfA6lAipus
+4jCHlfoeWn6r9RLPVCAKd66ny6R9z80dpdkyDVjjon3uQ5vPryd/neLnVYPF2/F
0YUZSL+9MRQrJU9qQFFvT90ORbUevkYnXLp8cyctAiXNYQafzzq6fnChhw8/vMwQ
DFChXg6VNXZcY+iV67NYur/mlZFVcFEBz1nrhJpG4BzieQmlp/9DwNAbvdalnTh7
TguFU1l8mGSANoz7xa/T9aKCDcbLvWnX8YCiykDKDvX2A2r5Tsqj7UIj101AFH+W
rqc2I2hppuaNlCtUoVG1xOF8otUR1FjoiW3GOVJXki3AktxzTz3SYU52ZiPKqcIh
NY14bgFcQ9orAYZbqR1J81qDR/dwTTeNa8tkNGxNyyiw2b/BJOEtIOiGMoM4/OWC
i1gza9Nh7cxlUh30pLGjhWrWWL0DBpHAsyzpLa+FUCJQQ/yB4M9d3JihmwWz5QUc
HSEd6AcFsxVizXqXFMCKAzxSaoWdMYzENeN1gFMYSihg7yHQDz2GfVzTrms0gRD1
yUrTOQkPSBHpcU4dAlGOqQ6xLyGtto5gJuhAF6J1JStHCKqqyR6OOMiMmNwAK50L
Au7DKdmf21WcW2a/NJyoqc3AeDGfkoMx0aeBQ+Piukm9rrT3Rtoal8E5snsOZHrc
7TqTWr5+qX1ev6mltR+8Xitgln7018Dm71LaVZog9bFDm81Iy/A8MAqLZ8EbZvL7
JBeCDZMXBdF08HNOTOFUQ9Id7Uc3VfUPOwGL2Gv1YRAOrC+pANUmcEwipVLuc6FZ
/H0pRIOxFwjDpSJC6cJOIpAahrOpscxPNTNXqaNg27cgKzA+gj3feSEwho9eVwE5
BctUTYblOZVQ6po1QRE/CI9zggwk+/RkM1V5ZHgHGWbgCoS9FvP079dMnY5vQiVW
ZnqUdp34hRgqmr75cntgaF1ZZ5gpEVPDNLvh4wHkLnKc9EZOUnYvWw7B2MyC3f6P
Nt6OO062UhNV181PnEfdF1Gpat8RMz78Ay0MJ3eiz0h0ya5ezxRhj4VpVn3+BSO2
Pb6x4+uvysVQzMDd59Jr2M2wkeId/xXLU0i/tykLtS3VIr6yokQxGSE4D2rTUcDp
oNYMHQAmxKg+Jw1MwEmUBuGA9Az0N4YdaIeimFq8NSux2396OxNXd8ePkyGudiMp
qMTAGSeDpydebZm2TKN8lydlFOoeyjp3fQOoV3jryuUAnBbVbUzJYVReOJG6PvQB
ezd2iGBw6jwv/wXC85UMOksTXcU2HqzaGpX3SqoJJetxlm8MF1wGg6Nw9Nsbyu1a
6VR1rjBmF+w/7nToOGtGWyulQ18IViY80F2ji1wB4oTEnRt215RuYAfB9IVRZiFC
glwjfapMj5fJc08gnOmiFfSobQ00RrTG67zE3UD/P8Y+xtO5liNfCPWAXBPWGlje
DkI7xipZszysWTj9vdi/QMhQ+uh+tHpt5HxIKqQo/W6MtmFsW3Z2qaEmAn97NiwO
o5vFYqdeGBoyhIEpo5RCFq/FbXavbZ5RB7TksFoWmziHS+1diOetFMIFtIWMZdOs
4Mbb0OlOhSYoU48FjcbF0iALVZZWTkd34iNDfjZKF8kwU9p4hBYiTaVVZv7Wdope
XGtQKrzun9wI5FIncqTDVd/UPzCxq8OZc8g+THxGm2IojBdsneGJ6KE8jkglHER8
kRRejuP+ZqAZU+UUbckBk1pRghOjEwB4ppr5/pKwVNT6ZpNE3lSD6SVzDMBKB77H
GfWZEImWmeyPGAsSvlFTjFI12UOJm3modJNOFWziiiPWiwKjRknAtAy48jIaQtDm
Ml07ECClGKJ0Dc1L1fMnXdoBOVJS0qiCeVIQ6EyGhsENgnql7w4S2CrKN4VdXPAn
qYXlIkrvYVdBlPO7H6ApqaS34MRBqdAwlaFQs64XF/VStQiTrtNzDaqoikx76TQF
WwOyTQuHDIjeu3Pq81boyzXDa1XP5MMkrhGSg11dXoFHlmYT0mOxun1hn/7me4t+
IOKCDTtZBwYvnNj5m5jSaIpWJugTFQoZEjVZUbCeZLoi4etBpV9H8bee9OyQ0YrX
a3yQSJnfUKkWkGTUpmidk3CClZ1GCr1e5DDwOnbQwsXf312bfNNV3rOgkt3JzL2R
hk2xf7o6LqKLW2C2aGqRAcKN+Q446z3mP7gcP6ChgXzgESp02eCEqIvCu8Rxmzaq
taLMOZbR/A5rype3tOPQ1Oarf5jqIHBAVAzl9S7bDMGFGxdy/4g/a2TOEQnDeXGJ
xSAhTluJKKa1FlWqR+65Ays6w/4R64+nhkOgJE1AKH6W6dt31xVRFkNjx8kAG9WB
vRs/cFX/Q0gQmkTxgR9HGxXClIoy9GOETy9Dpcx0rS7Jhtz8WzxdJ8B/aLPpMk6E
tV4PpyBmfzJbr1Y90YpYD2Dngp7Ahyd30JXv2bEpiQK+gq8Y5Pf4RI3Tnv4LS2cG
kFR7+U6gvPSrE0q6z1+ICunCsJmGUivxojMBNknlMCNF5GOtPq9HnAVVzyfW52bZ
pfolpjv47XwZXG7tc0cbEXEXrO58VEzqFDWu67d+N4bJ7fZPMv5YRsAe91pk2/iF
jIWCLN3JzMfnqO/cvx3gLdlf30DVjngwmcH50mJwK0cXeEFLpIfj7KhzKfWV1Wi5
mrfvsio8ZLkxEpJl4fCbSZnsax+VVhoBlyZPfnii8vSxW+Ec03JPnjGkKtzO1V1E
zmp9CX2tK3AFA4jXjnUYvgB3KRx3QdO+nEi0X/89rKWU6yS+EKd1ZiLR4v/r6BCk
VOLm8LgACMOMyxkKxJw2xJK/S9Azk+2r/MPpafjyGkgPoE43p1cJcplOgxU16MJX
bToHpANqVs9/p8hKrI67sHCPg0cromYtFT8LbFH51hdGh618aLE/w0778ppqRAdM
E+qEybBnsdCdTcsM1hvW9rmjO1OknUvxgxJbjUR+15HtqP0Ns9ue0wjCJWRZswCA
5RKu3iyO30qsIdLezZG/q48NSUhFIzmhFic83Wj/UQdCP32dnqamUsR/pGm+M+O8
Gp6gdig8bXiVws38uSC8YuSG0wcnPdeaZkxGdJGZgfQ3Fbo/8Wz/rUddyIwLyIhf
popA7fsNsBbHomofBMu8wUod3AmAKEpfGwD5DDdgYCxs47shFjpQUkysW6+/7uKY
TdkfOypa9J8x7qbEcRI+uNi+gXq8Lin0n+rW/z/IsnR2w8NjrWQagMJaKmUINu6f
Hny+ZMGw105aEXlU8E+8ywoOD5/jZgu3Hvs69wfiAQWaqLN40+m7wphEzyFi+GuE
n3u6vulzXbCRT9sdMr85r/7CxQChoPiKt+vkoR+HFJbBHsLCOqUM+6NVad3XWpBb
L4LcbbGg+O2n4qFgK/ek3zGFh1NutIFax0VAz/C4bFL6IrTCh1ktnkOa6GGx5Zqm
AX1immOL7/KH2Il0ZNar2ZYW3Lr83hB/cQcoYjdZRY9our8OONrb4K69kUyGp8hw
vGmLEdHcOYzzSUwVekgRAarmAXFTUEUOdcvP1EG/Qf5pTz+HOk3RqQLEgIpyIJmn
qG7S+76VLF3FpPtfi05Yclo//Rzcv4x6b5Dl+ellnIf5cG5/XFMhcnHWrg/MjZrr
YCxO1PPDLjGcSqrpEFwbYxx5r40igQ0k3nFucbcOjUDcj/Ejq8nTegNKQSOysvgE
nyDT+GLG//TQY8ke90Dlt0avHane9FeV72tzOrfQD2PfMI1GZMFNHFL9kotxr8KF
lkCph3e6OhCY2LIOR8yo2HP4Cf/gz9+MwPkMvuCrF8r7pfYCBvyYZ2jtVeAvxgA0
bZrW87UuTDpyG0nwdiaTLNIElDRJGZ/mjU3KMGlH0t9fOAumSwZZCvKzk69Juyon
lQq/cIQXntK3Zpio3Lc0XoH9vIte7sGaETmuMHjsPGaNVEvP1vKrQ/TE32TnUdoi
U6ahS88Y4UpUFB0mHdjJ8b4sIwkYOVT2X6ByY2QiVG51MLyiJ5qgTSp1h5y1wdUG
El1vuvWxYtWbJZe7Vq9wx/Opf3NSWxd2ph1HHNMKR/Bd7D3+awR/jW8TYGd9ByRI
MTN/hj24ga+ckyLBZzotOC98AMrQroVMnPU4oXJapwAdWWHrqMAR/FFjPlvDUoXD
IliZ/ZkLqut1osm0QGiiCiBn/6+BQpfc9TfI7/klvg4gq8wmXO4D4cpG+abVT28L
tvalVUUHRbYqGIwa2Xc3sIbOWWJ4h73Dubeo7Cb4u67UQBeWnp/2tABCL6t9zPJY
Cq+2NVrYAJD0lr3kKylloQrdW5qy67pFBnkOH07lArEQakvFBS5h7qoFg7BqmTZG
CT5gvDWS3G3dq35y1Es8tXsvSfi+d+oMzQBOPq+HnPm6Uz5+qgsE++JJp/CzyRfV
AziXcK5eSKU2EDQcuDjWcsZEL29BrLe8LIjUuG/FM97VSJzImDfSxV4bEiFdoIBa
1olcPG8HxNzY62NZnpZ8tENLxRqJV39Jk5thdgyc7DWFV2AmeYuWRWIensoYDTQ3
YQyTR6uwX/Z5VuvDWWol+iQusVdaPmWc8nUlhq3l2bf+ajTV/0/9yT/l884YO4GW
gU5rUYRoTGMCTVipKAoqnWXQDGyIYusxEwJbPJNp4Wn0lyLALg+cLUGOuYpZSxZh
LCgLvu3elTUtLfd2dmZa4/dhyohuWOho3/bvti4J7hTMur4Y41Cwl1l+25sjrvv1
No8LDLKWgimG9e6LUIYRa/Qe49O2dtgKHr0PrMp3v7bzYGB+l3L6vsGmXfGm7KUc
RSW6h1Np8sLjgUJo/847shCehUKC9hHMROUHBbbKM1fKUJr139tziA+u+nVsU4Gx
r2AsU58j3KP4bUHaa1099+GUdaq3tB+8ZtkKFLOXsrtuYCuoSX5x1VHE5QTzvltD
0fqS3juMbc9djm087KZ+uvCIgk4RXY2BQe/p1grRvK/sf3/H1BGSvnS14AScvWRV
8Ef7L6K19Sr9DbLmjKs+0TYYEQeof8scyFYcmTG3EpnRB8U8UpRZgsL21IIbq3Ce
XJ9jcGqtcQZZiA54ug3gFz+lIEr1nHNR2+5FUXqlyGpDcER+/WzDeqfGJPCf9v2h
WaOQYwgBxRK4zfBjpAwiNUIi4iC1wKDy++Izv90qAOyXpI34Hdh27wcs3VaqHBVF
cVl1XRyItVTdLrZ7yvugD5vJ7R73GhIP6fCZCNFeMIzaNxQ8F7ITfaNq/UlIBi92
vR4IBorDbHvAedrpU1soDX9Kx/YwYt84iJeR2oLoGUBzOduTkCUN+mv5KJUvncbw
19w79e3Bqj/Y9f6nNjhuTx9afQ2B/1u7Uz83P4jKZevZdbSU3qM5W7xqSZso+kO0
fWCsJ/wdv88EHLvkZw99IY2bmesCk+eT29WMDujKd6KPNYVMGBZgQ6mxUq7R8Naq
YIs/osV6R/0D1NYOnyBKRZzj3kO/cywUukU3R26FpBDsqjZtVJFQ0lN1KdF5IwFe
9P179Zr/jCU/13UNB2JbvKP8IyUCTTAdjT4K9y/zoSK26ub3tSKabp5ofAdJ/vbu
mT/fqq2t9vIRPGFT/x+PDggi30EKiQkfCVfpaOgsCqHzpPHGlUbUVKcIpOuWn24s
XEthSP3JCfklTjTZ/AcMFEbwGWXi5kehIuPFLC6njWR9PfPb6teHd3a5qFhkIjwu
0v7GH5b68PqoeGpTztBfkbR2tkolfY62RlvDu5d8R0r6r1+sG1XBAjaFmRpatpYz
6GeJn6ySmE222812Wa7RxgBls+0/7/KYdZkWFdsueFkqtLeLgYNtojZRDlsowuE/
BBELESDQfvWebT8V3VV/Rr3nhEC5JaLuolQPUUm7hAnkLfSXbtrueZtCHq+icpMZ
OibQF032PxI92hCV3qbfndLDvvyql96R048hY+ZCDbPauY9aVpQds4GdFncMovr8
1ov63WbaO1I56tJbrQhrkj0PJFQk9NA6kYMMBEquTzJWtAPKuP+6UF+K55//0UKl
my9NmwuciS3Hk/TZgnhqJvt6BG+61X5s6uQXcxitpFW8UfnDI7flZtOdAjg1A+VJ
6bIYHjC9shGsvHydN/cw3/pI32aXUHKoQorc4n4bFjJY61W3mMmQrfm0odJzQAdf
0p90hEQpYMZIoLFRGrWyYx6LYw9TrREsZIxVI7AZVAPV/Ief/i7WmA0x0zL+z8HF
eYWSu0ZqPq/eh9rbYXIDvG9J5I7h71mzPqDSR4qNA/uJhCbwkEwF6UaBJKLNbPYC
gV8J7MvgepKx5aXqkYkNab4F4JFHfRT01/OONBGqGrhKfOkn4tFyDcYBCBcm1CRt
Ej5Nyld18d/5QRUJuIZUpnDNi6KK1oLpDgXsbodKnfr3m32pDgqaR8WXObzKfVXG
agPPegX9A4o1BQUR9sUQ22ZgfceymbDtvP1YGdYgYhbpdzXbLz9WbgcRQaTPnbMN
l5LZkTqpE/BH8y7KVBm30x8wAZnO4mFOSUmIDTrTZyAk6TAYJLSZhDte68CLpV9+
myxSWLzVubmEZs+b7xdGvzGvQIuUTD9z2WBaKML4q2SEDEMOovB4zUISOVgtz03j
RlmMHJ3Pev/wWEYlaRR1xrk7368ZV1mmiNt3q33b0RNUtfbTNjvKUPDH4VqctdED
tvEndjl3jTcX/n1xdtfSg3V0OPF4+Glh3M1OqL4Js0boH9wkPX8O3DeSJHKr/tZ1
iadU2oZlHFGqZaOGiFmJxO6s9bB/6OfyYr7tFqlepXGTWU5Vtm8B3dPoRjyaK5JP
XrNa4svzl9l16wRo/ZAsIXEudVZh7/AykZQ70FC7vtY1g7EP7hmg6bqQutOtDXgy
jekIWqX3RYwc7b/ipVwmSdtQ8G/q4xmfMPWxmILCYggUWjui89tH0ZriNl7K3Ljl
6C86TBvDVBFrUjl83MN1noUVFiokizEgDKSu3lbcChZD/L5TxZCh68HCupk74EUk
wpnhm2pY8mJ03i9gP2OdMRUjO0Jrugak935jdH6U3oEHYDGjjHTJgeHRnmmqHb/4
ONcYIl28xnM+qCm/t1axNlui1LbMuIgbZTeVOZFbRq1TbFRjJh/mCTbPcsfI/J2J
jvSZP7BpQ2XO8I+ZcZe+pe20XYMGN1kDq3ubfT53dATfyuu9YXXShY1c+J7dknWd
w36/OUAp3auxQCzS9Dkh8sHWme45goFBqr51i3Rh0JXkltEhMnZNHE+cXMlNZem3
TqVzSIBGDayrAgCCnNerH12KYmrCj8tZD+/h1Vw/TeSx6l3NpMx1dYdLLskWnrn7
nvUCXhP/Z+A58qab08SdRX2liYY5RMLxmqb2jLXfPmb0/dkkOK2DVBzFXqxIO16x
PxrIb4aLMelfXqKrVnRkZBn9YMLtK6MletGtCwi2bfjaPrvth0ED7djbi1emjtFX
L+guAJGE3odEj2q9LzDPitKr/axXMXr7kblMkH0jKXdc1NgNXSe75iWVs1233Hq9
rf5iDulB65mdPzGKTs2jnp1CDDYYzH9ZnFpL5zMMjkGbxf3hhev5uGmZQsilUDwz
VY+V74cfQVmclxYYH5l0gsQpjH+g+AmMgRAPp1cCj7HU+89i3hmwmGAMh2ADwxQf
082KrA/RjeBn3LlhAADsadrCFWqFclgu5GdIoUzWepLQq/7iOxRX+fz2eSVMTyl8
LMXaPp3ZQNMMHUkMre4QBq2ZtsCg5y5ianVToLEMUG1WzxruWN2P6lHVOsb+5n8V
vCy+SxxslpHLAVLhDY9XqBs6i9MeIdO4Ua9EzGdfp6KGZImdNaWK1tUkZ2K9UQ/8
Rr5SzUVhYNfiZPKyRRciAQnzdNpVKl+InYiWKToA/3AqohIfZIk9pvMN0ZPKGY1/
6waYWfpHlprAAEo7A1SFcgrCgbyEbRyf3XScm1w8OVzgAO/d8cFmD63FczBKmQEt
g2WX4xEtwPa2rjJ0Q/ymzocXkDaHXhCs9uo9HiTAGG3MHjNdYh+K7OLcsbXNw1Q3
6q87xQVORHjh+L0cXvzLrQnJIYGiI0xOrRTr+0T08UHdPSv08drP2MTwLgqmNNOM
bVdNip5+whALjyF0jmSXhXin1+7B0WWlF290DHozI8XeSBoVm1gxjl/+g4R+Ii0q
cvkI9P+ANhngEkEFyM4JKP7ZzMa+hC3WgFZfmRemHc7azVy0u4ZLqea1Q0k/NlDo
7KmGdnxYRlDLvoPx4UTln89ukb+pQjCJqS9L58oEnZKA+4Y+80ZriLm83HTJ6qHy
5b87oXkm9Da6OwtItMRbT6184Id6Il6Rk8fhH0ZcZJzquzWhWPtgUu8eE4zHm1y1
KTPGyAhAriKslV3rSJ/pzFe9it6i1czT8PBq3csuSj6tUY+n/ikTiBxF+jWBbRVR
FOL2OGr4HaCd7A1gEDjmnyNOW6wjsETFemN/LFYEa6oOCUAYFpnQsuas54MRcS8G
SP+OFiDzCl/mkWpNsdtXGIKf+Z4AN/Tzb70RStrG6D/fE3LAyR91mCfx181EPKnt
00UqrWhcEeR2Mbi7y2UyAJGGq+9PIiOor46iawOviY2MprDpPb3kUqXZ8KCEsJy6
93jhZ5lVAvhvYhXYeKUmDYMqnHHn12C9T3LjDyJ9HVxxf+2K/+/bD/y9cXdmivxa
UjFfGk+M34XLK8tYrLz5CsNWIsqWaoCCQWcrst+N4NPLoXKmJlaIqkuEd5QWe2b+
Xz7xPsi/44upiURCg729pafqmjXB4LtRSSvxQBdIRGfb7FHAt0OpRxSu7l60b28O
OQKf3EFwF/rKjUUypcw1ElahAyOIxbOuoTAtBNYhoNdMFE0jcjvwdIvRxWiKO9TS
0sSjKsfHjHBd0mfVr6hfduhn8jGWx0PBuNgjD4HJj33VFWykhgtT6nvcfypxwYDT
wUPdhRHkQ5Deo91YZLGY6+U5cROuUfsIWOyB7KRY1aWL7kuQ9hU7mO80bQM4KcfP
p7ls1GtPalssnNllkvdvuOBMXdFtn2nEw9N+YH3Fpk4ahuNchOVXmmurM1JX4bsJ
56zcRGqTfeVmnR4XN8U0e//ZSWcf4HDwrzy5vVjB2NSUTqclCMcXglmtK/SVJBkr
sE4XoPxJX08A3+9pKPTw4PqrrO1/z31S+OgLmADjHlhUSpPybOKkk3AHyp3FI4YD
NVWZ/1ii5rNEEB7+sCCPiu5YxZVlEl0vAp9cKMCn8Iic+55xuRqf6A1+1XeC9c4/
PFa8Ww7NE2COfejGVck5obX4pNm8NDbAoEzHwPly7+Z90Kod+vrqylqu6z1XbNFd
EBdwEJoUWvUi9WpUVHdyV0SRFsrEzGtBjfdQmPVHwoeWn6q+RQQvcBrpQjDJ6Kbv
kVs4n9z3qee66bjPP0EBESnRikuzj1J2EGxx991LknJBkvSgXP379jjjz2LiRmmY
zQ4uFk8OwGykS/UhRaTanpSi72K1R/+PMnHzAmBdrexqQbWoSKhRLOF/vgY8flyK
J926D33UunbWuZfDvHDyjxIrIcgZm3haDmm1UxSI02Z9lRkPlMA/t33Vzn2CIr86
SYPujr3NFveMyERQJtWG3OmLzDZigAUsUK16TOMbzwztmUfC+GNtTQVkJP1Ieexl
0yMGwBLJaHnI7iOPMvSMh3XaoZMwrraeGGBmdGSrIzb6fSjlMfwlGeYm5AZRjCyU
VjqCvKDpCukh5mZBiSY+uigM/IAazgjSQOgfyFasvmbBnB+vIbuTy+kIKOPomVJo
pCezM1mlCiaZaBpxLTwybn/gH6rJD6hRopleAPoIsk4FQdaoJ1NSgSJQ6eUoI6DI
ahYXlYg9DpRmSR7Vju36ZBYGQkJ7IvKbG/JbU356ygDcjyYE3rCySc+m1LC/LNd8
PEBpcpysYDJ3bLKWR+/GwxZeWxddAeOU+s5+Et6S4djB9ahnS5x7UWCOAns6LFVk
P1kPPKaicKbK7hUvWyeQTUdrwgqJZxWr+RP2HLmN/nJbp+ZocNPDytnxc0spSyxv
8V33HGAsOyuCxBz0eYPif+bfSwnaH0uBNYNvHpXTnbFNfpiUgb4e4Peg9kS16Sog
0kAQTcUJRsq6fqnQn/Yra++ZGiltSZpKg/hRg6Qw/AnJ4sB77vkglZybO3EybdJM
IAixPtCJpXHjabWDqrBPeHKDPt5sHJUtTXMk6AnazcebhKPZZAQrVe5vgZxMEAgU
p4qpxv5y00CpKEAc9kMmOLiUJdF5btsNXCju2aVktWRstoAU0HcuwE9h5MJqWyHg
4Qrf7byN9QOa/AaBRf644Co8UHQ+G/3PtZ0mg3xXgfduFKjtVFdu+1dfBdartQPI
d3SW3bP4tidbATQ5HnGhk0GGHNA4Ikql/mR8uglGOtDOzs1cInyL7h5DwU7CAS9/
ljxO1+rhXx+B53Ij2mZeHS6Q8EAFhh0FllddDRJV6hKgLqVoj3qrLJ4H8Vsa+LaC
kb0C3gvqBnLWiLtfOV8GN9oIEA1i/YMsEpaL3QBhNLTYqabCqWALr0s9IgzVxhlx
bLYMQM9Sn2o5MaDOloCCw4tcrOuTQeAQpdweAN8uoKmbfKo+b+pWTjQS3iXiVb6W
MeHytoCLGaDdY2lPxc0fEohYY6q+JhlJCImjY5xrJw24mr7odWUP6/ty+Axms0T6
LepdwW9US0saTsbZ5+uR5GDtp3vyl2pvGMTJkgdGYOADc7GOSznpgJBmkxZCfes6
CzBX4GbPYOQrHCilr8ovbWv9WLmbKG63JrYsbEy2KCzlq5RrNoa5+g02b8rnsIpw
M1M0C725ySgpZPTbb8arWTrLvSMQtMeFpaqosayEt85EJ3x7nyf906MvX1fhRe/M
9+2JFaYtevuSpfFOTnxlPmXvLwW3VmINCLkTYs+Kzre88mXVpAMm6l2s2J93rKHh
O4HoI3TvMMCy0KglRRRLc1EJ7WDZU383T6CTSRkCcvbmIKxaijxyNL7fGy6FgH32
sCw9xPl154CYOUhBjtHqgIuJQVHcnp+a7kp9GBMJ1r2F44T6ylC/SQqvxlHd5vSE
h63IOjEVUdmi8NCyukqTstCdpO0S88mmUe3cCKyy+nRxfu/LGzGPk5bjk97bNI4I
gWS0mTxeCf2lF0m7R2/Ad6VCn8zxUjNoFzbdvNk+hPRz/CeVRSWsw43/Zc9M5+o3
6MXEzk/4yY6ZgcwzQ3ZVSFmy7Y3mHrJzyZ3GTiLhn/XLtd+SIhJ9DyuIZNgItcMb
PhD7hTNFueBW4iv/x1H24txoVeO658wAW2PRCqZpP4pAquliE+YUbbrh0+jUurjI
fZPiP3kFdBAhrcdSnRyQ+wybIZKp/2Igvj0YMOrcOk7bXV2Y2MAiaVqh19m6Xm9p
/YHI6777cAyDlh/rCN7eDuE5QpLmyykDqrKH46oUVO4DknPzLfmTiV2Bsm/S+kWY
Aw6CuTZlOF8cviyL7rHsOoPwiHmW1mo9VHbQFikY91S2lTvnAlknEm80ysyeDvz4
sdM5nYSigXRdw3TNLiuyLB3AgD+Hz9H1KSWcyU2eAaQVwVMZkvGdT0itN1k5IfX3
6V/+mcvJ6MD2zP7AlBR7VdyqtIFS4imaRPgiKyKlehC5cPBe57PDSgTp/mhDBtJE
YcufZx5LG+Lb90nU4VG0gayMx0oFuRF+lCqBmiTqOiqD8lHJebWNtlNEzPrC16HA
ni/AdqH69LR2NMzmzkxM663ilxxw1Nsl/DUvwZ2hR51EdtMaUpCWiJis480hgs/Y
T2KfQf5rd6svQeVNeje+ivjML/a248QiTaF+GTqOA5oWg3XtNW2ykafuV1xqJpeF
mk8p+hnv9vDz9pDZOEEEDP8ZJ40uCzVLoIj4bMQBubJc1fRiF3quoLWuy7hNXVVz
aao7XNs050n8bBKKwsJhP8G9nz4tjSeFVUFchFVHLcG8zjosIgNcGbXX6LWmwk8A
JURAJb07GOdYfOQj1kivoAKcvdLGbLaQto8fyWyDlyGLIvhyREgeRqnDNmLj6pOO
kIijkQW3FMOgxTU/u7ylVvOhlUWWZ0djgEhDp8fMUzNPRAPsxUlEwPXqHh879boc
kVMXQIP8YiVx/757nM34jIeliSkdefnbQ68aW1+pHijM1MWSTCy5YwhoISz/ugH9
MfxbK/CitKCWyocztavmUlIAI1m6HFgzMyYFut5D1bE731c4dDYTWM2UB/rMXFi1
eUkngaLMj09pzIGefQhN6UjYdw0O5gYk/IwAeAn4MHuHrRVY3EbAhqgTh1mWrb1w
HLDVt/jLm9kPWPD+qPV9JVxDOp4kKTCiKEPafbs0yCMV3LR/SfEnQ4nMNIrIyJuv
lpz1WNDF1Ezqx/PmNPkVzSic50KWBtB2wjM5TCMkj21ckeYXEiQjR9VZAvKZ9Uvt
hEGHYLGZf/gfFDHDtOK5cP4d9gEhCo3g1rqYeM4N6W47buuKadQr2LX0PPnIliGi
dy8p7xwTEbAiyoXjrpdn6g6/zTGeIQSfg963qUa5k3qvPpevF2+EijjF6IJpns2j
LGWLSO24+caaVluhBgbHwI01HvSQ6ZRsi+6PEI3EdmuizRQzm8xbyP0RZDW16OJ8
3P2DU1HtCHlrOI+/zZ7ohHA5id/BtezFv7pUG6AWH3pdq6xoHFcUT54oVdTznORm
4fTwDoeMP6JnqEieXlSeAHPOS588eah6iihA6FbSjZDUAbiTv3qy6bm2o50NvzSa
7xEYwM/PeXuQBvtKrYmhWC7yKprSWXA4Tn8KzAT3BTYUUpn51i3wAvWJJAYUKlIu
lij8gumlKnQWz813vBbgA/bdI4w1EkidB1yhgutK1eIFrwNyKH8/MJKNNmArHusl
o+6/uYjQsr2/+3GCs38FRp+rBJ+u5JrfHIEQjy3vJJ9CuTDhP70eqp9ubfjVLzmw
pMLSgDGVUWMb3tORnf3GnaSpojLS/Nt4JXUGOY40Keg6I/tr/wS5eSgLeRGeEi0n
C4N+mY3JT/LlIlqLXyue3coifAGjng82hhz/46XObDHEQ8ryQj8xDAo5f9ogZf9f
fFqQlPRM33yZg4rRyjIt51mm3X/5bvU8DHV4Q+6mVj5FrhSdOOLCno58K3FBYfS7
JwCrQ2lSstFTWc4bDQU+qhuoyWjw50hP1xB5P0qjeCj7+9EYRigEJLga1mojMvqm
qzP6qTeeLyCqhVi+DprHx2Sq23xPplThz38ryzMXzGh1kgFqp8C4nMRpbPVJ+g+B
WvOcedyHlqp1FMLC3bJvZEsmKwjg/73dB83+wDt38aXE1sHAZzZcy7+OAyK50GDY
IEs5a61j+q0shVZh85LRQSUUhCBGMFitGZckE7C0CrKf3S5aWT7Y7+2YR6FKgWhb
ZNWVIwEfA88BCeOC96tvUPCNQ9B82V4qEbIlP1aaDHpzsIjIk59/eEY+TmPzs/TO
lksWa5hfy66tK1Vo468f+v2P9pp9tVUDUMvvnkbsZi2cVxjznX5ZsUC6ec2w6Pvh
PheDR3Ngyt/emhV5EmzAvP6OZ5vyj8onIFrKT+or9e4hURLLewAHUOH++4bF2a6g
4y6mPFVVVVapwBSbHio6s9ShVCWZgkGbrZ9EjGdEzoY8kx3WQR+9sIE/JwjKIKvp
a30K7PyG5VRWK06+f3Un+yBBLFUusFisJZ8SKQH2OE5yXJxY3YSDdtwKQFqNeZbb
gP97w47UPEuothlBWQ0iPzTHikeoxvlnIhVSBLY+QSfBWxbPvBN03dQzv04YOIzx
EcB0Wrtf2f+i3iNRLKNvR5AChF6Yw8hQX+W38F1KaZpv0PYxF1+NHhHPW+zTQzEd
FhXshjU1Vzh9zi2Ha5IePB+kYKEHa4kunMC0B+ObbusF+RIiSQOYE5S4Yx88LtNl
f/rkLGcoN5hatRGmCcvOwA==
`pragma protect end_protected
